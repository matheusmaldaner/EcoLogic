library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(5119 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(5119 downto 0);
    signal layer1_outputs : std_logic_vector(5119 downto 0);
    signal layer2_outputs : std_logic_vector(5119 downto 0);
    signal layer3_outputs : std_logic_vector(5119 downto 0);
    signal layer4_outputs : std_logic_vector(5119 downto 0);
    signal layer5_outputs : std_logic_vector(5119 downto 0);
    signal layer6_outputs : std_logic_vector(5119 downto 0);
    signal layer7_outputs : std_logic_vector(5119 downto 0);
    signal layer8_outputs : std_logic_vector(5119 downto 0);

begin

    layer0_outputs(0) <= '1';
    layer0_outputs(1) <= '1';
    layer0_outputs(2) <= not((inputs(134)) and (inputs(68)));
    layer0_outputs(3) <= '0';
    layer0_outputs(4) <= not((inputs(32)) or (inputs(62)));
    layer0_outputs(5) <= '1';
    layer0_outputs(6) <= (inputs(138)) or (inputs(232));
    layer0_outputs(7) <= (inputs(100)) and not (inputs(253));
    layer0_outputs(8) <= '0';
    layer0_outputs(9) <= (inputs(2)) or (inputs(110));
    layer0_outputs(10) <= not((inputs(205)) and (inputs(31)));
    layer0_outputs(11) <= inputs(197);
    layer0_outputs(12) <= not(inputs(78)) or (inputs(38));
    layer0_outputs(13) <= '1';
    layer0_outputs(14) <= (inputs(86)) or (inputs(115));
    layer0_outputs(15) <= (inputs(141)) or (inputs(15));
    layer0_outputs(16) <= (inputs(63)) xor (inputs(189));
    layer0_outputs(17) <= inputs(20);
    layer0_outputs(18) <= (inputs(132)) or (inputs(149));
    layer0_outputs(19) <= inputs(39);
    layer0_outputs(20) <= not(inputs(118));
    layer0_outputs(21) <= not(inputs(237)) or (inputs(61));
    layer0_outputs(22) <= not(inputs(23)) or (inputs(240));
    layer0_outputs(23) <= '0';
    layer0_outputs(24) <= '1';
    layer0_outputs(25) <= not((inputs(161)) and (inputs(230)));
    layer0_outputs(26) <= '0';
    layer0_outputs(27) <= '0';
    layer0_outputs(28) <= '0';
    layer0_outputs(29) <= (inputs(193)) and not (inputs(195));
    layer0_outputs(30) <= inputs(76);
    layer0_outputs(31) <= not((inputs(61)) or (inputs(224)));
    layer0_outputs(32) <= inputs(184);
    layer0_outputs(33) <= not((inputs(176)) and (inputs(134)));
    layer0_outputs(34) <= (inputs(5)) and (inputs(108));
    layer0_outputs(35) <= (inputs(235)) and not (inputs(245));
    layer0_outputs(36) <= not(inputs(14)) or (inputs(137));
    layer0_outputs(37) <= '0';
    layer0_outputs(38) <= (inputs(68)) and not (inputs(229));
    layer0_outputs(39) <= '1';
    layer0_outputs(40) <= inputs(56);
    layer0_outputs(41) <= (inputs(201)) and (inputs(180));
    layer0_outputs(42) <= '0';
    layer0_outputs(43) <= not(inputs(85)) or (inputs(204));
    layer0_outputs(44) <= '0';
    layer0_outputs(45) <= inputs(123);
    layer0_outputs(46) <= (inputs(113)) and not (inputs(27));
    layer0_outputs(47) <= inputs(192);
    layer0_outputs(48) <= (inputs(189)) and not (inputs(101));
    layer0_outputs(49) <= not(inputs(21));
    layer0_outputs(50) <= not((inputs(254)) and (inputs(72)));
    layer0_outputs(51) <= not((inputs(15)) xor (inputs(116)));
    layer0_outputs(52) <= '0';
    layer0_outputs(53) <= '0';
    layer0_outputs(54) <= not(inputs(53)) or (inputs(150));
    layer0_outputs(55) <= (inputs(12)) and not (inputs(253));
    layer0_outputs(56) <= (inputs(27)) and (inputs(253));
    layer0_outputs(57) <= '0';
    layer0_outputs(58) <= (inputs(237)) xor (inputs(122));
    layer0_outputs(59) <= '1';
    layer0_outputs(60) <= '1';
    layer0_outputs(61) <= (inputs(12)) and not (inputs(93));
    layer0_outputs(62) <= not(inputs(110)) or (inputs(248));
    layer0_outputs(63) <= '0';
    layer0_outputs(64) <= inputs(162);
    layer0_outputs(65) <= inputs(29);
    layer0_outputs(66) <= '0';
    layer0_outputs(67) <= not(inputs(52));
    layer0_outputs(68) <= not(inputs(183)) or (inputs(4));
    layer0_outputs(69) <= (inputs(151)) xor (inputs(98));
    layer0_outputs(70) <= '1';
    layer0_outputs(71) <= inputs(119);
    layer0_outputs(72) <= not(inputs(93));
    layer0_outputs(73) <= '0';
    layer0_outputs(74) <= inputs(36);
    layer0_outputs(75) <= '1';
    layer0_outputs(76) <= inputs(162);
    layer0_outputs(77) <= (inputs(13)) or (inputs(76));
    layer0_outputs(78) <= not(inputs(253));
    layer0_outputs(79) <= not(inputs(181));
    layer0_outputs(80) <= not(inputs(200)) or (inputs(190));
    layer0_outputs(81) <= inputs(104);
    layer0_outputs(82) <= inputs(108);
    layer0_outputs(83) <= not((inputs(198)) or (inputs(194)));
    layer0_outputs(84) <= not(inputs(199)) or (inputs(17));
    layer0_outputs(85) <= (inputs(43)) and (inputs(10));
    layer0_outputs(86) <= not((inputs(95)) and (inputs(117)));
    layer0_outputs(87) <= '0';
    layer0_outputs(88) <= not(inputs(247));
    layer0_outputs(89) <= '0';
    layer0_outputs(90) <= not(inputs(212));
    layer0_outputs(91) <= not(inputs(2));
    layer0_outputs(92) <= (inputs(241)) or (inputs(210));
    layer0_outputs(93) <= not(inputs(210));
    layer0_outputs(94) <= inputs(210);
    layer0_outputs(95) <= (inputs(23)) or (inputs(64));
    layer0_outputs(96) <= (inputs(223)) and not (inputs(82));
    layer0_outputs(97) <= not((inputs(184)) or (inputs(165)));
    layer0_outputs(98) <= (inputs(139)) and (inputs(184));
    layer0_outputs(99) <= not(inputs(201));
    layer0_outputs(100) <= (inputs(182)) and not (inputs(183));
    layer0_outputs(101) <= not((inputs(104)) or (inputs(231)));
    layer0_outputs(102) <= not(inputs(54)) or (inputs(44));
    layer0_outputs(103) <= '0';
    layer0_outputs(104) <= '0';
    layer0_outputs(105) <= '1';
    layer0_outputs(106) <= (inputs(29)) and not (inputs(235));
    layer0_outputs(107) <= '1';
    layer0_outputs(108) <= not(inputs(143));
    layer0_outputs(109) <= (inputs(42)) and not (inputs(28));
    layer0_outputs(110) <= not(inputs(28));
    layer0_outputs(111) <= not(inputs(135)) or (inputs(117));
    layer0_outputs(112) <= '1';
    layer0_outputs(113) <= not(inputs(201));
    layer0_outputs(114) <= not((inputs(185)) and (inputs(92)));
    layer0_outputs(115) <= inputs(227);
    layer0_outputs(116) <= '1';
    layer0_outputs(117) <= not(inputs(230)) or (inputs(219));
    layer0_outputs(118) <= (inputs(169)) and (inputs(137));
    layer0_outputs(119) <= not(inputs(203)) or (inputs(111));
    layer0_outputs(120) <= not(inputs(197)) or (inputs(83));
    layer0_outputs(121) <= not(inputs(255)) or (inputs(63));
    layer0_outputs(122) <= (inputs(146)) xor (inputs(113));
    layer0_outputs(123) <= '1';
    layer0_outputs(124) <= not(inputs(187));
    layer0_outputs(125) <= (inputs(31)) or (inputs(205));
    layer0_outputs(126) <= (inputs(140)) and not (inputs(41));
    layer0_outputs(127) <= (inputs(61)) or (inputs(95));
    layer0_outputs(128) <= (inputs(105)) and (inputs(38));
    layer0_outputs(129) <= '0';
    layer0_outputs(130) <= not(inputs(246));
    layer0_outputs(131) <= not(inputs(146));
    layer0_outputs(132) <= '0';
    layer0_outputs(133) <= (inputs(194)) or (inputs(108));
    layer0_outputs(134) <= inputs(1);
    layer0_outputs(135) <= not(inputs(61)) or (inputs(178));
    layer0_outputs(136) <= inputs(183);
    layer0_outputs(137) <= '0';
    layer0_outputs(138) <= '0';
    layer0_outputs(139) <= inputs(139);
    layer0_outputs(140) <= not(inputs(71)) or (inputs(34));
    layer0_outputs(141) <= '1';
    layer0_outputs(142) <= not(inputs(7));
    layer0_outputs(143) <= '0';
    layer0_outputs(144) <= not((inputs(181)) and (inputs(142)));
    layer0_outputs(145) <= '0';
    layer0_outputs(146) <= not(inputs(136));
    layer0_outputs(147) <= (inputs(54)) or (inputs(127));
    layer0_outputs(148) <= (inputs(104)) and (inputs(181));
    layer0_outputs(149) <= not(inputs(141)) or (inputs(126));
    layer0_outputs(150) <= '1';
    layer0_outputs(151) <= '1';
    layer0_outputs(152) <= not((inputs(95)) and (inputs(156)));
    layer0_outputs(153) <= '0';
    layer0_outputs(154) <= not((inputs(141)) or (inputs(29)));
    layer0_outputs(155) <= inputs(148);
    layer0_outputs(156) <= not(inputs(63)) or (inputs(67));
    layer0_outputs(157) <= (inputs(240)) and (inputs(152));
    layer0_outputs(158) <= '0';
    layer0_outputs(159) <= (inputs(36)) and not (inputs(51));
    layer0_outputs(160) <= '0';
    layer0_outputs(161) <= inputs(127);
    layer0_outputs(162) <= inputs(210);
    layer0_outputs(163) <= not((inputs(144)) and (inputs(61)));
    layer0_outputs(164) <= (inputs(170)) xor (inputs(168));
    layer0_outputs(165) <= (inputs(224)) and (inputs(12));
    layer0_outputs(166) <= not((inputs(112)) and (inputs(55)));
    layer0_outputs(167) <= (inputs(126)) or (inputs(197));
    layer0_outputs(168) <= not(inputs(14));
    layer0_outputs(169) <= (inputs(27)) and not (inputs(84));
    layer0_outputs(170) <= inputs(101);
    layer0_outputs(171) <= '1';
    layer0_outputs(172) <= (inputs(46)) xor (inputs(121));
    layer0_outputs(173) <= not(inputs(140));
    layer0_outputs(174) <= not(inputs(0));
    layer0_outputs(175) <= not((inputs(138)) and (inputs(190)));
    layer0_outputs(176) <= (inputs(180)) or (inputs(238));
    layer0_outputs(177) <= '1';
    layer0_outputs(178) <= '0';
    layer0_outputs(179) <= '0';
    layer0_outputs(180) <= not((inputs(19)) or (inputs(143)));
    layer0_outputs(181) <= (inputs(64)) and not (inputs(209));
    layer0_outputs(182) <= inputs(48);
    layer0_outputs(183) <= (inputs(127)) or (inputs(245));
    layer0_outputs(184) <= (inputs(246)) and not (inputs(67));
    layer0_outputs(185) <= not(inputs(85)) or (inputs(251));
    layer0_outputs(186) <= not(inputs(248)) or (inputs(238));
    layer0_outputs(187) <= '0';
    layer0_outputs(188) <= '0';
    layer0_outputs(189) <= not(inputs(18)) or (inputs(30));
    layer0_outputs(190) <= '1';
    layer0_outputs(191) <= '1';
    layer0_outputs(192) <= inputs(177);
    layer0_outputs(193) <= not((inputs(157)) or (inputs(150)));
    layer0_outputs(194) <= (inputs(31)) or (inputs(125));
    layer0_outputs(195) <= not(inputs(96));
    layer0_outputs(196) <= (inputs(137)) and not (inputs(199));
    layer0_outputs(197) <= (inputs(231)) or (inputs(71));
    layer0_outputs(198) <= (inputs(88)) and not (inputs(112));
    layer0_outputs(199) <= not(inputs(186)) or (inputs(109));
    layer0_outputs(200) <= (inputs(94)) and (inputs(30));
    layer0_outputs(201) <= inputs(110);
    layer0_outputs(202) <= inputs(236);
    layer0_outputs(203) <= '1';
    layer0_outputs(204) <= not(inputs(21));
    layer0_outputs(205) <= (inputs(235)) and not (inputs(101));
    layer0_outputs(206) <= not(inputs(211)) or (inputs(150));
    layer0_outputs(207) <= '0';
    layer0_outputs(208) <= '1';
    layer0_outputs(209) <= '1';
    layer0_outputs(210) <= inputs(210);
    layer0_outputs(211) <= (inputs(61)) and not (inputs(154));
    layer0_outputs(212) <= not(inputs(1)) or (inputs(193));
    layer0_outputs(213) <= not(inputs(217));
    layer0_outputs(214) <= not(inputs(96));
    layer0_outputs(215) <= inputs(101);
    layer0_outputs(216) <= (inputs(151)) and not (inputs(5));
    layer0_outputs(217) <= not((inputs(141)) and (inputs(214)));
    layer0_outputs(218) <= '1';
    layer0_outputs(219) <= '1';
    layer0_outputs(220) <= not(inputs(255)) or (inputs(68));
    layer0_outputs(221) <= inputs(110);
    layer0_outputs(222) <= not((inputs(141)) xor (inputs(172)));
    layer0_outputs(223) <= (inputs(233)) or (inputs(255));
    layer0_outputs(224) <= inputs(194);
    layer0_outputs(225) <= not(inputs(18));
    layer0_outputs(226) <= not(inputs(49));
    layer0_outputs(227) <= not(inputs(95));
    layer0_outputs(228) <= inputs(62);
    layer0_outputs(229) <= not(inputs(94)) or (inputs(17));
    layer0_outputs(230) <= (inputs(127)) and (inputs(221));
    layer0_outputs(231) <= '0';
    layer0_outputs(232) <= not((inputs(95)) and (inputs(5)));
    layer0_outputs(233) <= not(inputs(221));
    layer0_outputs(234) <= (inputs(143)) and not (inputs(57));
    layer0_outputs(235) <= '1';
    layer0_outputs(236) <= '1';
    layer0_outputs(237) <= not((inputs(110)) and (inputs(39)));
    layer0_outputs(238) <= (inputs(103)) or (inputs(1));
    layer0_outputs(239) <= (inputs(115)) xor (inputs(70));
    layer0_outputs(240) <= inputs(255);
    layer0_outputs(241) <= '0';
    layer0_outputs(242) <= (inputs(10)) and not (inputs(13));
    layer0_outputs(243) <= '0';
    layer0_outputs(244) <= '1';
    layer0_outputs(245) <= inputs(75);
    layer0_outputs(246) <= (inputs(105)) and not (inputs(178));
    layer0_outputs(247) <= inputs(48);
    layer0_outputs(248) <= (inputs(113)) and not (inputs(92));
    layer0_outputs(249) <= inputs(119);
    layer0_outputs(250) <= (inputs(166)) and not (inputs(174));
    layer0_outputs(251) <= inputs(30);
    layer0_outputs(252) <= not(inputs(13)) or (inputs(39));
    layer0_outputs(253) <= '0';
    layer0_outputs(254) <= '0';
    layer0_outputs(255) <= '0';
    layer0_outputs(256) <= not(inputs(248));
    layer0_outputs(257) <= '1';
    layer0_outputs(258) <= (inputs(23)) and not (inputs(209));
    layer0_outputs(259) <= inputs(160);
    layer0_outputs(260) <= not(inputs(142));
    layer0_outputs(261) <= not(inputs(150)) or (inputs(63));
    layer0_outputs(262) <= inputs(12);
    layer0_outputs(263) <= not((inputs(229)) and (inputs(147)));
    layer0_outputs(264) <= inputs(63);
    layer0_outputs(265) <= inputs(253);
    layer0_outputs(266) <= inputs(202);
    layer0_outputs(267) <= not(inputs(201));
    layer0_outputs(268) <= '0';
    layer0_outputs(269) <= '0';
    layer0_outputs(270) <= (inputs(249)) and not (inputs(188));
    layer0_outputs(271) <= not(inputs(4));
    layer0_outputs(272) <= (inputs(65)) or (inputs(133));
    layer0_outputs(273) <= (inputs(169)) or (inputs(232));
    layer0_outputs(274) <= (inputs(33)) or (inputs(223));
    layer0_outputs(275) <= (inputs(155)) and not (inputs(255));
    layer0_outputs(276) <= inputs(34);
    layer0_outputs(277) <= (inputs(6)) and (inputs(216));
    layer0_outputs(278) <= not((inputs(161)) or (inputs(246)));
    layer0_outputs(279) <= not(inputs(202)) or (inputs(173));
    layer0_outputs(280) <= inputs(150);
    layer0_outputs(281) <= (inputs(62)) or (inputs(22));
    layer0_outputs(282) <= not((inputs(241)) and (inputs(4)));
    layer0_outputs(283) <= '1';
    layer0_outputs(284) <= inputs(161);
    layer0_outputs(285) <= '0';
    layer0_outputs(286) <= (inputs(114)) xor (inputs(84));
    layer0_outputs(287) <= not((inputs(209)) or (inputs(229)));
    layer0_outputs(288) <= inputs(94);
    layer0_outputs(289) <= not((inputs(133)) xor (inputs(193)));
    layer0_outputs(290) <= not((inputs(21)) or (inputs(173)));
    layer0_outputs(291) <= not(inputs(246)) or (inputs(220));
    layer0_outputs(292) <= (inputs(169)) and not (inputs(20));
    layer0_outputs(293) <= (inputs(183)) and (inputs(169));
    layer0_outputs(294) <= not((inputs(7)) and (inputs(100)));
    layer0_outputs(295) <= '1';
    layer0_outputs(296) <= not(inputs(69)) or (inputs(118));
    layer0_outputs(297) <= (inputs(49)) and not (inputs(91));
    layer0_outputs(298) <= (inputs(214)) and not (inputs(119));
    layer0_outputs(299) <= (inputs(192)) and (inputs(55));
    layer0_outputs(300) <= '1';
    layer0_outputs(301) <= (inputs(56)) or (inputs(73));
    layer0_outputs(302) <= inputs(154);
    layer0_outputs(303) <= inputs(252);
    layer0_outputs(304) <= '1';
    layer0_outputs(305) <= '1';
    layer0_outputs(306) <= (inputs(35)) and not (inputs(54));
    layer0_outputs(307) <= (inputs(2)) or (inputs(255));
    layer0_outputs(308) <= inputs(175);
    layer0_outputs(309) <= not((inputs(69)) and (inputs(118)));
    layer0_outputs(310) <= (inputs(216)) and not (inputs(52));
    layer0_outputs(311) <= not((inputs(44)) and (inputs(185)));
    layer0_outputs(312) <= not(inputs(253)) or (inputs(61));
    layer0_outputs(313) <= '1';
    layer0_outputs(314) <= inputs(122);
    layer0_outputs(315) <= not((inputs(0)) and (inputs(119)));
    layer0_outputs(316) <= inputs(112);
    layer0_outputs(317) <= '1';
    layer0_outputs(318) <= '0';
    layer0_outputs(319) <= (inputs(31)) or (inputs(127));
    layer0_outputs(320) <= inputs(232);
    layer0_outputs(321) <= not(inputs(186));
    layer0_outputs(322) <= not(inputs(78));
    layer0_outputs(323) <= not(inputs(193)) or (inputs(48));
    layer0_outputs(324) <= not((inputs(45)) and (inputs(7)));
    layer0_outputs(325) <= '0';
    layer0_outputs(326) <= not((inputs(94)) and (inputs(175)));
    layer0_outputs(327) <= '0';
    layer0_outputs(328) <= not((inputs(81)) and (inputs(165)));
    layer0_outputs(329) <= (inputs(184)) or (inputs(134));
    layer0_outputs(330) <= inputs(221);
    layer0_outputs(331) <= (inputs(121)) xor (inputs(73));
    layer0_outputs(332) <= (inputs(70)) and (inputs(146));
    layer0_outputs(333) <= (inputs(89)) and (inputs(205));
    layer0_outputs(334) <= not((inputs(101)) or (inputs(221)));
    layer0_outputs(335) <= (inputs(43)) or (inputs(229));
    layer0_outputs(336) <= not((inputs(42)) and (inputs(254)));
    layer0_outputs(337) <= inputs(151);
    layer0_outputs(338) <= (inputs(163)) or (inputs(141));
    layer0_outputs(339) <= '0';
    layer0_outputs(340) <= inputs(15);
    layer0_outputs(341) <= (inputs(107)) and not (inputs(167));
    layer0_outputs(342) <= '1';
    layer0_outputs(343) <= '0';
    layer0_outputs(344) <= not(inputs(143));
    layer0_outputs(345) <= (inputs(176)) and not (inputs(203));
    layer0_outputs(346) <= not(inputs(3));
    layer0_outputs(347) <= not((inputs(28)) and (inputs(130)));
    layer0_outputs(348) <= (inputs(218)) or (inputs(234));
    layer0_outputs(349) <= not(inputs(43));
    layer0_outputs(350) <= (inputs(203)) and (inputs(45));
    layer0_outputs(351) <= inputs(255);
    layer0_outputs(352) <= not((inputs(124)) or (inputs(116)));
    layer0_outputs(353) <= inputs(138);
    layer0_outputs(354) <= inputs(6);
    layer0_outputs(355) <= not((inputs(157)) or (inputs(47)));
    layer0_outputs(356) <= not(inputs(168));
    layer0_outputs(357) <= (inputs(71)) and (inputs(22));
    layer0_outputs(358) <= not(inputs(85));
    layer0_outputs(359) <= '1';
    layer0_outputs(360) <= (inputs(219)) or (inputs(172));
    layer0_outputs(361) <= not((inputs(224)) or (inputs(33)));
    layer0_outputs(362) <= '0';
    layer0_outputs(363) <= not(inputs(184));
    layer0_outputs(364) <= inputs(39);
    layer0_outputs(365) <= '0';
    layer0_outputs(366) <= not((inputs(153)) or (inputs(215)));
    layer0_outputs(367) <= '1';
    layer0_outputs(368) <= not(inputs(88)) or (inputs(10));
    layer0_outputs(369) <= inputs(2);
    layer0_outputs(370) <= (inputs(242)) and not (inputs(23));
    layer0_outputs(371) <= '0';
    layer0_outputs(372) <= (inputs(156)) and (inputs(191));
    layer0_outputs(373) <= '0';
    layer0_outputs(374) <= not((inputs(232)) or (inputs(225)));
    layer0_outputs(375) <= (inputs(12)) and not (inputs(184));
    layer0_outputs(376) <= inputs(1);
    layer0_outputs(377) <= not(inputs(105)) or (inputs(189));
    layer0_outputs(378) <= '0';
    layer0_outputs(379) <= '1';
    layer0_outputs(380) <= (inputs(159)) and not (inputs(79));
    layer0_outputs(381) <= inputs(252);
    layer0_outputs(382) <= not(inputs(174));
    layer0_outputs(383) <= '0';
    layer0_outputs(384) <= not((inputs(236)) and (inputs(138)));
    layer0_outputs(385) <= '1';
    layer0_outputs(386) <= inputs(18);
    layer0_outputs(387) <= '1';
    layer0_outputs(388) <= not((inputs(247)) and (inputs(196)));
    layer0_outputs(389) <= '1';
    layer0_outputs(390) <= not((inputs(89)) or (inputs(41)));
    layer0_outputs(391) <= '0';
    layer0_outputs(392) <= not((inputs(41)) xor (inputs(87)));
    layer0_outputs(393) <= (inputs(103)) or (inputs(163));
    layer0_outputs(394) <= not(inputs(196));
    layer0_outputs(395) <= not((inputs(65)) or (inputs(208)));
    layer0_outputs(396) <= '0';
    layer0_outputs(397) <= '0';
    layer0_outputs(398) <= not(inputs(99)) or (inputs(226));
    layer0_outputs(399) <= '0';
    layer0_outputs(400) <= '1';
    layer0_outputs(401) <= (inputs(0)) and not (inputs(178));
    layer0_outputs(402) <= not(inputs(211)) or (inputs(2));
    layer0_outputs(403) <= not(inputs(145));
    layer0_outputs(404) <= (inputs(77)) xor (inputs(4));
    layer0_outputs(405) <= '0';
    layer0_outputs(406) <= (inputs(14)) and not (inputs(122));
    layer0_outputs(407) <= inputs(76);
    layer0_outputs(408) <= inputs(162);
    layer0_outputs(409) <= not(inputs(106));
    layer0_outputs(410) <= '1';
    layer0_outputs(411) <= '1';
    layer0_outputs(412) <= '1';
    layer0_outputs(413) <= inputs(239);
    layer0_outputs(414) <= not(inputs(57)) or (inputs(191));
    layer0_outputs(415) <= '1';
    layer0_outputs(416) <= (inputs(145)) and not (inputs(81));
    layer0_outputs(417) <= not(inputs(170)) or (inputs(187));
    layer0_outputs(418) <= not(inputs(81));
    layer0_outputs(419) <= not((inputs(178)) and (inputs(216)));
    layer0_outputs(420) <= not(inputs(96));
    layer0_outputs(421) <= inputs(128);
    layer0_outputs(422) <= not(inputs(160));
    layer0_outputs(423) <= (inputs(49)) or (inputs(22));
    layer0_outputs(424) <= not(inputs(125));
    layer0_outputs(425) <= (inputs(176)) or (inputs(241));
    layer0_outputs(426) <= (inputs(170)) or (inputs(110));
    layer0_outputs(427) <= '1';
    layer0_outputs(428) <= '1';
    layer0_outputs(429) <= not(inputs(12));
    layer0_outputs(430) <= '1';
    layer0_outputs(431) <= not(inputs(159));
    layer0_outputs(432) <= (inputs(2)) and not (inputs(209));
    layer0_outputs(433) <= not(inputs(148)) or (inputs(152));
    layer0_outputs(434) <= not(inputs(130));
    layer0_outputs(435) <= not(inputs(82));
    layer0_outputs(436) <= (inputs(99)) and not (inputs(124));
    layer0_outputs(437) <= '1';
    layer0_outputs(438) <= not(inputs(59));
    layer0_outputs(439) <= not((inputs(46)) and (inputs(213)));
    layer0_outputs(440) <= '1';
    layer0_outputs(441) <= not((inputs(3)) and (inputs(252)));
    layer0_outputs(442) <= not((inputs(9)) and (inputs(135)));
    layer0_outputs(443) <= '1';
    layer0_outputs(444) <= inputs(129);
    layer0_outputs(445) <= '0';
    layer0_outputs(446) <= not(inputs(63));
    layer0_outputs(447) <= not(inputs(41)) or (inputs(31));
    layer0_outputs(448) <= (inputs(132)) or (inputs(200));
    layer0_outputs(449) <= '0';
    layer0_outputs(450) <= (inputs(211)) and (inputs(12));
    layer0_outputs(451) <= '0';
    layer0_outputs(452) <= not((inputs(119)) and (inputs(126)));
    layer0_outputs(453) <= (inputs(87)) and not (inputs(89));
    layer0_outputs(454) <= (inputs(56)) and (inputs(18));
    layer0_outputs(455) <= not((inputs(176)) or (inputs(199)));
    layer0_outputs(456) <= (inputs(131)) or (inputs(85));
    layer0_outputs(457) <= (inputs(6)) xor (inputs(158));
    layer0_outputs(458) <= not((inputs(235)) or (inputs(171)));
    layer0_outputs(459) <= inputs(254);
    layer0_outputs(460) <= '0';
    layer0_outputs(461) <= '1';
    layer0_outputs(462) <= not(inputs(205));
    layer0_outputs(463) <= not((inputs(159)) and (inputs(196)));
    layer0_outputs(464) <= (inputs(146)) or (inputs(196));
    layer0_outputs(465) <= (inputs(156)) and not (inputs(172));
    layer0_outputs(466) <= inputs(95);
    layer0_outputs(467) <= '1';
    layer0_outputs(468) <= not(inputs(104)) or (inputs(40));
    layer0_outputs(469) <= not(inputs(16));
    layer0_outputs(470) <= inputs(158);
    layer0_outputs(471) <= inputs(227);
    layer0_outputs(472) <= inputs(169);
    layer0_outputs(473) <= inputs(94);
    layer0_outputs(474) <= '0';
    layer0_outputs(475) <= '0';
    layer0_outputs(476) <= not(inputs(47));
    layer0_outputs(477) <= not((inputs(159)) and (inputs(230)));
    layer0_outputs(478) <= not((inputs(85)) and (inputs(79)));
    layer0_outputs(479) <= inputs(134);
    layer0_outputs(480) <= not(inputs(72));
    layer0_outputs(481) <= '1';
    layer0_outputs(482) <= '0';
    layer0_outputs(483) <= (inputs(112)) or (inputs(110));
    layer0_outputs(484) <= inputs(26);
    layer0_outputs(485) <= inputs(239);
    layer0_outputs(486) <= not((inputs(230)) or (inputs(212)));
    layer0_outputs(487) <= inputs(225);
    layer0_outputs(488) <= '1';
    layer0_outputs(489) <= inputs(77);
    layer0_outputs(490) <= '0';
    layer0_outputs(491) <= not(inputs(165));
    layer0_outputs(492) <= (inputs(65)) or (inputs(101));
    layer0_outputs(493) <= not(inputs(21));
    layer0_outputs(494) <= (inputs(54)) and (inputs(232));
    layer0_outputs(495) <= not(inputs(34));
    layer0_outputs(496) <= inputs(57);
    layer0_outputs(497) <= inputs(206);
    layer0_outputs(498) <= '1';
    layer0_outputs(499) <= '1';
    layer0_outputs(500) <= inputs(150);
    layer0_outputs(501) <= not(inputs(178));
    layer0_outputs(502) <= (inputs(133)) or (inputs(67));
    layer0_outputs(503) <= not(inputs(59));
    layer0_outputs(504) <= '1';
    layer0_outputs(505) <= not((inputs(127)) or (inputs(92)));
    layer0_outputs(506) <= (inputs(69)) and not (inputs(89));
    layer0_outputs(507) <= '1';
    layer0_outputs(508) <= not((inputs(105)) and (inputs(96)));
    layer0_outputs(509) <= '1';
    layer0_outputs(510) <= inputs(15);
    layer0_outputs(511) <= '0';
    layer0_outputs(512) <= not((inputs(231)) and (inputs(219)));
    layer0_outputs(513) <= not(inputs(162));
    layer0_outputs(514) <= not(inputs(20));
    layer0_outputs(515) <= (inputs(161)) or (inputs(252));
    layer0_outputs(516) <= not(inputs(251));
    layer0_outputs(517) <= '0';
    layer0_outputs(518) <= not(inputs(7)) or (inputs(116));
    layer0_outputs(519) <= not(inputs(72));
    layer0_outputs(520) <= not((inputs(201)) xor (inputs(200)));
    layer0_outputs(521) <= inputs(121);
    layer0_outputs(522) <= inputs(51);
    layer0_outputs(523) <= (inputs(106)) xor (inputs(79));
    layer0_outputs(524) <= not((inputs(63)) and (inputs(217)));
    layer0_outputs(525) <= (inputs(78)) and not (inputs(24));
    layer0_outputs(526) <= '0';
    layer0_outputs(527) <= not(inputs(103));
    layer0_outputs(528) <= (inputs(160)) and not (inputs(187));
    layer0_outputs(529) <= (inputs(133)) and not (inputs(213));
    layer0_outputs(530) <= (inputs(65)) and not (inputs(31));
    layer0_outputs(531) <= (inputs(154)) and not (inputs(221));
    layer0_outputs(532) <= inputs(18);
    layer0_outputs(533) <= not((inputs(173)) and (inputs(227)));
    layer0_outputs(534) <= '0';
    layer0_outputs(535) <= not((inputs(220)) xor (inputs(112)));
    layer0_outputs(536) <= (inputs(206)) or (inputs(32));
    layer0_outputs(537) <= '0';
    layer0_outputs(538) <= (inputs(84)) and not (inputs(0));
    layer0_outputs(539) <= inputs(120);
    layer0_outputs(540) <= '1';
    layer0_outputs(541) <= inputs(73);
    layer0_outputs(542) <= inputs(244);
    layer0_outputs(543) <= not(inputs(236)) or (inputs(103));
    layer0_outputs(544) <= (inputs(145)) and not (inputs(95));
    layer0_outputs(545) <= (inputs(93)) xor (inputs(33));
    layer0_outputs(546) <= (inputs(252)) or (inputs(91));
    layer0_outputs(547) <= '1';
    layer0_outputs(548) <= inputs(224);
    layer0_outputs(549) <= not((inputs(67)) and (inputs(181)));
    layer0_outputs(550) <= not((inputs(168)) or (inputs(182)));
    layer0_outputs(551) <= not((inputs(159)) and (inputs(59)));
    layer0_outputs(552) <= not(inputs(47));
    layer0_outputs(553) <= not(inputs(131)) or (inputs(216));
    layer0_outputs(554) <= (inputs(138)) and (inputs(45));
    layer0_outputs(555) <= inputs(33);
    layer0_outputs(556) <= (inputs(247)) or (inputs(97));
    layer0_outputs(557) <= not(inputs(129));
    layer0_outputs(558) <= '0';
    layer0_outputs(559) <= not((inputs(37)) and (inputs(130)));
    layer0_outputs(560) <= not(inputs(195));
    layer0_outputs(561) <= '0';
    layer0_outputs(562) <= '0';
    layer0_outputs(563) <= not(inputs(46));
    layer0_outputs(564) <= inputs(25);
    layer0_outputs(565) <= inputs(135);
    layer0_outputs(566) <= inputs(185);
    layer0_outputs(567) <= '1';
    layer0_outputs(568) <= not(inputs(165)) or (inputs(117));
    layer0_outputs(569) <= (inputs(208)) xor (inputs(37));
    layer0_outputs(570) <= not(inputs(24));
    layer0_outputs(571) <= not((inputs(67)) xor (inputs(67)));
    layer0_outputs(572) <= '0';
    layer0_outputs(573) <= (inputs(243)) and not (inputs(0));
    layer0_outputs(574) <= inputs(5);
    layer0_outputs(575) <= (inputs(87)) or (inputs(231));
    layer0_outputs(576) <= inputs(27);
    layer0_outputs(577) <= (inputs(68)) and (inputs(74));
    layer0_outputs(578) <= (inputs(214)) and (inputs(217));
    layer0_outputs(579) <= (inputs(233)) or (inputs(238));
    layer0_outputs(580) <= not(inputs(137));
    layer0_outputs(581) <= inputs(131);
    layer0_outputs(582) <= (inputs(202)) and not (inputs(65));
    layer0_outputs(583) <= '1';
    layer0_outputs(584) <= '0';
    layer0_outputs(585) <= (inputs(93)) and not (inputs(167));
    layer0_outputs(586) <= (inputs(146)) or (inputs(56));
    layer0_outputs(587) <= '0';
    layer0_outputs(588) <= not(inputs(203)) or (inputs(110));
    layer0_outputs(589) <= '0';
    layer0_outputs(590) <= not(inputs(31));
    layer0_outputs(591) <= '1';
    layer0_outputs(592) <= (inputs(135)) and not (inputs(233));
    layer0_outputs(593) <= not((inputs(155)) or (inputs(78)));
    layer0_outputs(594) <= (inputs(1)) or (inputs(219));
    layer0_outputs(595) <= '1';
    layer0_outputs(596) <= not(inputs(126)) or (inputs(51));
    layer0_outputs(597) <= not(inputs(99));
    layer0_outputs(598) <= inputs(64);
    layer0_outputs(599) <= not(inputs(186));
    layer0_outputs(600) <= not(inputs(61));
    layer0_outputs(601) <= not(inputs(103));
    layer0_outputs(602) <= not(inputs(190)) or (inputs(9));
    layer0_outputs(603) <= (inputs(68)) or (inputs(58));
    layer0_outputs(604) <= (inputs(197)) xor (inputs(163));
    layer0_outputs(605) <= not(inputs(121));
    layer0_outputs(606) <= (inputs(87)) and not (inputs(66));
    layer0_outputs(607) <= inputs(109);
    layer0_outputs(608) <= '1';
    layer0_outputs(609) <= '0';
    layer0_outputs(610) <= '1';
    layer0_outputs(611) <= not(inputs(10));
    layer0_outputs(612) <= not((inputs(63)) or (inputs(220)));
    layer0_outputs(613) <= (inputs(32)) and not (inputs(41));
    layer0_outputs(614) <= not(inputs(0));
    layer0_outputs(615) <= (inputs(229)) xor (inputs(243));
    layer0_outputs(616) <= inputs(70);
    layer0_outputs(617) <= not((inputs(13)) and (inputs(231)));
    layer0_outputs(618) <= not(inputs(76));
    layer0_outputs(619) <= not((inputs(5)) and (inputs(52)));
    layer0_outputs(620) <= '1';
    layer0_outputs(621) <= inputs(121);
    layer0_outputs(622) <= '1';
    layer0_outputs(623) <= (inputs(36)) and not (inputs(127));
    layer0_outputs(624) <= inputs(190);
    layer0_outputs(625) <= not((inputs(155)) or (inputs(230)));
    layer0_outputs(626) <= '0';
    layer0_outputs(627) <= not(inputs(145)) or (inputs(154));
    layer0_outputs(628) <= not((inputs(140)) or (inputs(127)));
    layer0_outputs(629) <= (inputs(39)) xor (inputs(32));
    layer0_outputs(630) <= '1';
    layer0_outputs(631) <= not(inputs(49));
    layer0_outputs(632) <= inputs(150);
    layer0_outputs(633) <= not(inputs(94));
    layer0_outputs(634) <= not(inputs(103)) or (inputs(9));
    layer0_outputs(635) <= inputs(127);
    layer0_outputs(636) <= (inputs(142)) and (inputs(206));
    layer0_outputs(637) <= (inputs(223)) and not (inputs(94));
    layer0_outputs(638) <= not(inputs(59));
    layer0_outputs(639) <= not(inputs(204));
    layer0_outputs(640) <= inputs(234);
    layer0_outputs(641) <= (inputs(28)) or (inputs(83));
    layer0_outputs(642) <= (inputs(254)) and not (inputs(124));
    layer0_outputs(643) <= inputs(242);
    layer0_outputs(644) <= not((inputs(173)) and (inputs(52)));
    layer0_outputs(645) <= not(inputs(161)) or (inputs(130));
    layer0_outputs(646) <= (inputs(66)) and not (inputs(90));
    layer0_outputs(647) <= (inputs(215)) and not (inputs(65));
    layer0_outputs(648) <= (inputs(162)) and (inputs(169));
    layer0_outputs(649) <= (inputs(173)) and (inputs(222));
    layer0_outputs(650) <= (inputs(3)) and not (inputs(96));
    layer0_outputs(651) <= not((inputs(227)) xor (inputs(88)));
    layer0_outputs(652) <= '1';
    layer0_outputs(653) <= (inputs(136)) and not (inputs(26));
    layer0_outputs(654) <= not(inputs(246)) or (inputs(67));
    layer0_outputs(655) <= inputs(110);
    layer0_outputs(656) <= (inputs(87)) and not (inputs(6));
    layer0_outputs(657) <= not(inputs(0)) or (inputs(46));
    layer0_outputs(658) <= '0';
    layer0_outputs(659) <= inputs(145);
    layer0_outputs(660) <= '1';
    layer0_outputs(661) <= '0';
    layer0_outputs(662) <= inputs(142);
    layer0_outputs(663) <= '1';
    layer0_outputs(664) <= not(inputs(12));
    layer0_outputs(665) <= '0';
    layer0_outputs(666) <= inputs(107);
    layer0_outputs(667) <= not((inputs(37)) and (inputs(252)));
    layer0_outputs(668) <= (inputs(50)) or (inputs(219));
    layer0_outputs(669) <= '0';
    layer0_outputs(670) <= (inputs(192)) or (inputs(244));
    layer0_outputs(671) <= '1';
    layer0_outputs(672) <= (inputs(0)) and not (inputs(197));
    layer0_outputs(673) <= (inputs(251)) xor (inputs(110));
    layer0_outputs(674) <= not((inputs(138)) xor (inputs(33)));
    layer0_outputs(675) <= not((inputs(142)) and (inputs(253)));
    layer0_outputs(676) <= not(inputs(119)) or (inputs(153));
    layer0_outputs(677) <= (inputs(1)) or (inputs(130));
    layer0_outputs(678) <= not((inputs(48)) or (inputs(152)));
    layer0_outputs(679) <= '0';
    layer0_outputs(680) <= (inputs(36)) and not (inputs(97));
    layer0_outputs(681) <= not(inputs(101));
    layer0_outputs(682) <= '1';
    layer0_outputs(683) <= '0';
    layer0_outputs(684) <= not((inputs(191)) or (inputs(142)));
    layer0_outputs(685) <= (inputs(57)) and (inputs(67));
    layer0_outputs(686) <= (inputs(239)) and (inputs(85));
    layer0_outputs(687) <= (inputs(223)) and not (inputs(20));
    layer0_outputs(688) <= inputs(124);
    layer0_outputs(689) <= inputs(81);
    layer0_outputs(690) <= inputs(208);
    layer0_outputs(691) <= (inputs(35)) xor (inputs(97));
    layer0_outputs(692) <= (inputs(165)) and not (inputs(80));
    layer0_outputs(693) <= (inputs(216)) or (inputs(53));
    layer0_outputs(694) <= '0';
    layer0_outputs(695) <= (inputs(80)) and not (inputs(93));
    layer0_outputs(696) <= inputs(161);
    layer0_outputs(697) <= (inputs(67)) and (inputs(152));
    layer0_outputs(698) <= not((inputs(78)) and (inputs(170)));
    layer0_outputs(699) <= (inputs(82)) and not (inputs(135));
    layer0_outputs(700) <= inputs(179);
    layer0_outputs(701) <= inputs(38);
    layer0_outputs(702) <= inputs(68);
    layer0_outputs(703) <= '0';
    layer0_outputs(704) <= not((inputs(89)) or (inputs(16)));
    layer0_outputs(705) <= not(inputs(193)) or (inputs(68));
    layer0_outputs(706) <= not(inputs(120));
    layer0_outputs(707) <= not(inputs(77));
    layer0_outputs(708) <= not(inputs(194)) or (inputs(111));
    layer0_outputs(709) <= not((inputs(57)) xor (inputs(117)));
    layer0_outputs(710) <= (inputs(84)) and not (inputs(178));
    layer0_outputs(711) <= '1';
    layer0_outputs(712) <= not(inputs(81));
    layer0_outputs(713) <= not(inputs(235)) or (inputs(67));
    layer0_outputs(714) <= not((inputs(22)) or (inputs(62)));
    layer0_outputs(715) <= not((inputs(235)) or (inputs(204)));
    layer0_outputs(716) <= '1';
    layer0_outputs(717) <= not((inputs(185)) or (inputs(157)));
    layer0_outputs(718) <= not((inputs(81)) and (inputs(23)));
    layer0_outputs(719) <= inputs(67);
    layer0_outputs(720) <= not(inputs(142));
    layer0_outputs(721) <= inputs(141);
    layer0_outputs(722) <= not((inputs(86)) xor (inputs(102)));
    layer0_outputs(723) <= inputs(250);
    layer0_outputs(724) <= not(inputs(159));
    layer0_outputs(725) <= (inputs(68)) and not (inputs(102));
    layer0_outputs(726) <= '1';
    layer0_outputs(727) <= (inputs(242)) and (inputs(90));
    layer0_outputs(728) <= '1';
    layer0_outputs(729) <= (inputs(107)) or (inputs(106));
    layer0_outputs(730) <= '0';
    layer0_outputs(731) <= '0';
    layer0_outputs(732) <= inputs(7);
    layer0_outputs(733) <= '1';
    layer0_outputs(734) <= '0';
    layer0_outputs(735) <= '0';
    layer0_outputs(736) <= '0';
    layer0_outputs(737) <= '1';
    layer0_outputs(738) <= '1';
    layer0_outputs(739) <= '0';
    layer0_outputs(740) <= not(inputs(120)) or (inputs(176));
    layer0_outputs(741) <= not(inputs(245)) or (inputs(81));
    layer0_outputs(742) <= '1';
    layer0_outputs(743) <= inputs(202);
    layer0_outputs(744) <= inputs(112);
    layer0_outputs(745) <= '0';
    layer0_outputs(746) <= (inputs(174)) or (inputs(192));
    layer0_outputs(747) <= inputs(161);
    layer0_outputs(748) <= not((inputs(225)) or (inputs(20)));
    layer0_outputs(749) <= not(inputs(255));
    layer0_outputs(750) <= '0';
    layer0_outputs(751) <= not(inputs(203));
    layer0_outputs(752) <= (inputs(42)) and not (inputs(231));
    layer0_outputs(753) <= (inputs(147)) xor (inputs(169));
    layer0_outputs(754) <= not((inputs(59)) xor (inputs(225)));
    layer0_outputs(755) <= (inputs(101)) and (inputs(33));
    layer0_outputs(756) <= (inputs(67)) and not (inputs(67));
    layer0_outputs(757) <= '0';
    layer0_outputs(758) <= (inputs(122)) xor (inputs(154));
    layer0_outputs(759) <= '0';
    layer0_outputs(760) <= not((inputs(153)) or (inputs(168)));
    layer0_outputs(761) <= '1';
    layer0_outputs(762) <= inputs(116);
    layer0_outputs(763) <= (inputs(226)) and not (inputs(100));
    layer0_outputs(764) <= inputs(147);
    layer0_outputs(765) <= not((inputs(249)) and (inputs(65)));
    layer0_outputs(766) <= not(inputs(168)) or (inputs(86));
    layer0_outputs(767) <= '1';
    layer0_outputs(768) <= not((inputs(63)) and (inputs(15)));
    layer0_outputs(769) <= (inputs(227)) and not (inputs(185));
    layer0_outputs(770) <= '0';
    layer0_outputs(771) <= (inputs(132)) and not (inputs(71));
    layer0_outputs(772) <= (inputs(133)) and (inputs(75));
    layer0_outputs(773) <= '1';
    layer0_outputs(774) <= '1';
    layer0_outputs(775) <= '1';
    layer0_outputs(776) <= not(inputs(222));
    layer0_outputs(777) <= not((inputs(79)) xor (inputs(175)));
    layer0_outputs(778) <= '0';
    layer0_outputs(779) <= '0';
    layer0_outputs(780) <= '0';
    layer0_outputs(781) <= not(inputs(111));
    layer0_outputs(782) <= (inputs(35)) and not (inputs(219));
    layer0_outputs(783) <= (inputs(45)) and (inputs(53));
    layer0_outputs(784) <= '1';
    layer0_outputs(785) <= not(inputs(118));
    layer0_outputs(786) <= (inputs(63)) and not (inputs(243));
    layer0_outputs(787) <= not(inputs(180)) or (inputs(141));
    layer0_outputs(788) <= not(inputs(67)) or (inputs(207));
    layer0_outputs(789) <= inputs(23);
    layer0_outputs(790) <= not(inputs(210)) or (inputs(10));
    layer0_outputs(791) <= (inputs(197)) and (inputs(165));
    layer0_outputs(792) <= '0';
    layer0_outputs(793) <= '0';
    layer0_outputs(794) <= (inputs(206)) and not (inputs(105));
    layer0_outputs(795) <= not((inputs(202)) and (inputs(32)));
    layer0_outputs(796) <= (inputs(249)) and not (inputs(158));
    layer0_outputs(797) <= not(inputs(232));
    layer0_outputs(798) <= not((inputs(132)) xor (inputs(71)));
    layer0_outputs(799) <= inputs(220);
    layer0_outputs(800) <= '1';
    layer0_outputs(801) <= not(inputs(141));
    layer0_outputs(802) <= (inputs(174)) and not (inputs(140));
    layer0_outputs(803) <= not((inputs(104)) and (inputs(84)));
    layer0_outputs(804) <= not(inputs(122));
    layer0_outputs(805) <= not(inputs(12));
    layer0_outputs(806) <= (inputs(142)) and not (inputs(19));
    layer0_outputs(807) <= inputs(138);
    layer0_outputs(808) <= '0';
    layer0_outputs(809) <= '0';
    layer0_outputs(810) <= '1';
    layer0_outputs(811) <= not(inputs(222));
    layer0_outputs(812) <= (inputs(224)) and not (inputs(169));
    layer0_outputs(813) <= (inputs(0)) xor (inputs(75));
    layer0_outputs(814) <= not(inputs(165)) or (inputs(85));
    layer0_outputs(815) <= (inputs(219)) or (inputs(63));
    layer0_outputs(816) <= not(inputs(106)) or (inputs(113));
    layer0_outputs(817) <= inputs(77);
    layer0_outputs(818) <= '0';
    layer0_outputs(819) <= '1';
    layer0_outputs(820) <= not(inputs(93)) or (inputs(210));
    layer0_outputs(821) <= (inputs(86)) or (inputs(115));
    layer0_outputs(822) <= (inputs(149)) xor (inputs(190));
    layer0_outputs(823) <= inputs(151);
    layer0_outputs(824) <= not(inputs(133));
    layer0_outputs(825) <= not(inputs(120)) or (inputs(69));
    layer0_outputs(826) <= not(inputs(167));
    layer0_outputs(827) <= '0';
    layer0_outputs(828) <= not((inputs(206)) and (inputs(50)));
    layer0_outputs(829) <= not((inputs(178)) or (inputs(248)));
    layer0_outputs(830) <= (inputs(137)) and (inputs(51));
    layer0_outputs(831) <= inputs(177);
    layer0_outputs(832) <= (inputs(32)) and not (inputs(248));
    layer0_outputs(833) <= '0';
    layer0_outputs(834) <= (inputs(215)) and (inputs(195));
    layer0_outputs(835) <= not((inputs(206)) and (inputs(87)));
    layer0_outputs(836) <= not((inputs(237)) and (inputs(127)));
    layer0_outputs(837) <= inputs(191);
    layer0_outputs(838) <= (inputs(61)) xor (inputs(47));
    layer0_outputs(839) <= inputs(240);
    layer0_outputs(840) <= '0';
    layer0_outputs(841) <= not((inputs(98)) or (inputs(149)));
    layer0_outputs(842) <= '1';
    layer0_outputs(843) <= '1';
    layer0_outputs(844) <= (inputs(125)) and (inputs(50));
    layer0_outputs(845) <= not(inputs(212)) or (inputs(27));
    layer0_outputs(846) <= not(inputs(104)) or (inputs(129));
    layer0_outputs(847) <= '0';
    layer0_outputs(848) <= '0';
    layer0_outputs(849) <= '0';
    layer0_outputs(850) <= inputs(25);
    layer0_outputs(851) <= not(inputs(241)) or (inputs(27));
    layer0_outputs(852) <= '1';
    layer0_outputs(853) <= not(inputs(201)) or (inputs(229));
    layer0_outputs(854) <= '1';
    layer0_outputs(855) <= not(inputs(25));
    layer0_outputs(856) <= (inputs(214)) and not (inputs(24));
    layer0_outputs(857) <= not((inputs(148)) and (inputs(207)));
    layer0_outputs(858) <= '1';
    layer0_outputs(859) <= not((inputs(142)) or (inputs(237)));
    layer0_outputs(860) <= not((inputs(152)) and (inputs(241)));
    layer0_outputs(861) <= inputs(140);
    layer0_outputs(862) <= '0';
    layer0_outputs(863) <= (inputs(204)) or (inputs(71));
    layer0_outputs(864) <= not(inputs(145));
    layer0_outputs(865) <= (inputs(0)) and not (inputs(175));
    layer0_outputs(866) <= not((inputs(1)) and (inputs(40)));
    layer0_outputs(867) <= '1';
    layer0_outputs(868) <= not((inputs(178)) and (inputs(12)));
    layer0_outputs(869) <= '0';
    layer0_outputs(870) <= not((inputs(234)) and (inputs(251)));
    layer0_outputs(871) <= not(inputs(31)) or (inputs(77));
    layer0_outputs(872) <= (inputs(184)) and not (inputs(197));
    layer0_outputs(873) <= (inputs(85)) and (inputs(32));
    layer0_outputs(874) <= inputs(222);
    layer0_outputs(875) <= (inputs(180)) or (inputs(148));
    layer0_outputs(876) <= not(inputs(131));
    layer0_outputs(877) <= not((inputs(93)) and (inputs(108)));
    layer0_outputs(878) <= '1';
    layer0_outputs(879) <= not((inputs(189)) and (inputs(255)));
    layer0_outputs(880) <= (inputs(247)) and not (inputs(222));
    layer0_outputs(881) <= not((inputs(43)) and (inputs(70)));
    layer0_outputs(882) <= '0';
    layer0_outputs(883) <= '1';
    layer0_outputs(884) <= inputs(164);
    layer0_outputs(885) <= not(inputs(159)) or (inputs(19));
    layer0_outputs(886) <= inputs(73);
    layer0_outputs(887) <= inputs(182);
    layer0_outputs(888) <= inputs(47);
    layer0_outputs(889) <= '0';
    layer0_outputs(890) <= '1';
    layer0_outputs(891) <= not(inputs(132)) or (inputs(230));
    layer0_outputs(892) <= inputs(245);
    layer0_outputs(893) <= '1';
    layer0_outputs(894) <= not((inputs(52)) or (inputs(155)));
    layer0_outputs(895) <= not(inputs(180));
    layer0_outputs(896) <= not((inputs(18)) and (inputs(55)));
    layer0_outputs(897) <= inputs(230);
    layer0_outputs(898) <= not(inputs(171));
    layer0_outputs(899) <= (inputs(218)) and not (inputs(58));
    layer0_outputs(900) <= (inputs(77)) or (inputs(90));
    layer0_outputs(901) <= not(inputs(214)) or (inputs(236));
    layer0_outputs(902) <= (inputs(149)) or (inputs(34));
    layer0_outputs(903) <= not(inputs(123));
    layer0_outputs(904) <= not(inputs(160));
    layer0_outputs(905) <= '0';
    layer0_outputs(906) <= (inputs(176)) and not (inputs(130));
    layer0_outputs(907) <= not(inputs(241)) or (inputs(153));
    layer0_outputs(908) <= not(inputs(233));
    layer0_outputs(909) <= '1';
    layer0_outputs(910) <= not(inputs(192));
    layer0_outputs(911) <= not(inputs(238));
    layer0_outputs(912) <= not(inputs(197));
    layer0_outputs(913) <= (inputs(211)) or (inputs(107));
    layer0_outputs(914) <= (inputs(217)) or (inputs(219));
    layer0_outputs(915) <= not((inputs(65)) or (inputs(22)));
    layer0_outputs(916) <= not(inputs(191)) or (inputs(1));
    layer0_outputs(917) <= (inputs(165)) xor (inputs(194));
    layer0_outputs(918) <= '0';
    layer0_outputs(919) <= inputs(53);
    layer0_outputs(920) <= not((inputs(21)) and (inputs(251)));
    layer0_outputs(921) <= '0';
    layer0_outputs(922) <= (inputs(154)) and (inputs(195));
    layer0_outputs(923) <= not(inputs(67));
    layer0_outputs(924) <= (inputs(33)) and not (inputs(100));
    layer0_outputs(925) <= (inputs(78)) and not (inputs(31));
    layer0_outputs(926) <= inputs(36);
    layer0_outputs(927) <= (inputs(102)) and (inputs(64));
    layer0_outputs(928) <= not(inputs(234));
    layer0_outputs(929) <= '0';
    layer0_outputs(930) <= not(inputs(229));
    layer0_outputs(931) <= '1';
    layer0_outputs(932) <= '0';
    layer0_outputs(933) <= not((inputs(77)) and (inputs(171)));
    layer0_outputs(934) <= not((inputs(147)) and (inputs(227)));
    layer0_outputs(935) <= not(inputs(251));
    layer0_outputs(936) <= not((inputs(34)) and (inputs(47)));
    layer0_outputs(937) <= inputs(18);
    layer0_outputs(938) <= inputs(228);
    layer0_outputs(939) <= (inputs(175)) and not (inputs(166));
    layer0_outputs(940) <= not(inputs(163)) or (inputs(174));
    layer0_outputs(941) <= '1';
    layer0_outputs(942) <= (inputs(194)) xor (inputs(37));
    layer0_outputs(943) <= not(inputs(176));
    layer0_outputs(944) <= not((inputs(120)) or (inputs(63)));
    layer0_outputs(945) <= '0';
    layer0_outputs(946) <= '0';
    layer0_outputs(947) <= not((inputs(87)) and (inputs(168)));
    layer0_outputs(948) <= '0';
    layer0_outputs(949) <= '1';
    layer0_outputs(950) <= inputs(22);
    layer0_outputs(951) <= not(inputs(95)) or (inputs(98));
    layer0_outputs(952) <= not((inputs(199)) and (inputs(38)));
    layer0_outputs(953) <= '1';
    layer0_outputs(954) <= inputs(140);
    layer0_outputs(955) <= (inputs(185)) and (inputs(16));
    layer0_outputs(956) <= '1';
    layer0_outputs(957) <= inputs(191);
    layer0_outputs(958) <= not((inputs(76)) or (inputs(66)));
    layer0_outputs(959) <= '0';
    layer0_outputs(960) <= '1';
    layer0_outputs(961) <= inputs(29);
    layer0_outputs(962) <= (inputs(35)) and not (inputs(230));
    layer0_outputs(963) <= not((inputs(146)) or (inputs(212)));
    layer0_outputs(964) <= '1';
    layer0_outputs(965) <= (inputs(252)) and not (inputs(54));
    layer0_outputs(966) <= '0';
    layer0_outputs(967) <= '1';
    layer0_outputs(968) <= '1';
    layer0_outputs(969) <= (inputs(79)) and (inputs(125));
    layer0_outputs(970) <= not(inputs(64));
    layer0_outputs(971) <= not(inputs(161));
    layer0_outputs(972) <= not((inputs(132)) and (inputs(93)));
    layer0_outputs(973) <= inputs(43);
    layer0_outputs(974) <= not(inputs(104));
    layer0_outputs(975) <= not((inputs(102)) or (inputs(255)));
    layer0_outputs(976) <= not(inputs(198)) or (inputs(234));
    layer0_outputs(977) <= not(inputs(60)) or (inputs(2));
    layer0_outputs(978) <= (inputs(32)) and not (inputs(157));
    layer0_outputs(979) <= not((inputs(148)) xor (inputs(255)));
    layer0_outputs(980) <= (inputs(120)) or (inputs(206));
    layer0_outputs(981) <= not(inputs(92)) or (inputs(58));
    layer0_outputs(982) <= '0';
    layer0_outputs(983) <= (inputs(16)) and (inputs(200));
    layer0_outputs(984) <= '1';
    layer0_outputs(985) <= not(inputs(193)) or (inputs(4));
    layer0_outputs(986) <= (inputs(176)) or (inputs(246));
    layer0_outputs(987) <= '1';
    layer0_outputs(988) <= not(inputs(94));
    layer0_outputs(989) <= '0';
    layer0_outputs(990) <= not(inputs(210)) or (inputs(215));
    layer0_outputs(991) <= inputs(96);
    layer0_outputs(992) <= '1';
    layer0_outputs(993) <= inputs(94);
    layer0_outputs(994) <= not((inputs(96)) or (inputs(162)));
    layer0_outputs(995) <= not((inputs(47)) xor (inputs(253)));
    layer0_outputs(996) <= inputs(228);
    layer0_outputs(997) <= not(inputs(90));
    layer0_outputs(998) <= inputs(158);
    layer0_outputs(999) <= not(inputs(161)) or (inputs(249));
    layer0_outputs(1000) <= inputs(6);
    layer0_outputs(1001) <= '1';
    layer0_outputs(1002) <= not(inputs(240));
    layer0_outputs(1003) <= (inputs(239)) and not (inputs(229));
    layer0_outputs(1004) <= (inputs(241)) and (inputs(74));
    layer0_outputs(1005) <= not((inputs(51)) or (inputs(169)));
    layer0_outputs(1006) <= '0';
    layer0_outputs(1007) <= not(inputs(179)) or (inputs(151));
    layer0_outputs(1008) <= not(inputs(209)) or (inputs(121));
    layer0_outputs(1009) <= not(inputs(173));
    layer0_outputs(1010) <= '1';
    layer0_outputs(1011) <= not((inputs(222)) and (inputs(208)));
    layer0_outputs(1012) <= '0';
    layer0_outputs(1013) <= (inputs(6)) and not (inputs(54));
    layer0_outputs(1014) <= (inputs(124)) or (inputs(111));
    layer0_outputs(1015) <= not(inputs(175)) or (inputs(158));
    layer0_outputs(1016) <= (inputs(125)) xor (inputs(90));
    layer0_outputs(1017) <= not(inputs(97));
    layer0_outputs(1018) <= inputs(100);
    layer0_outputs(1019) <= (inputs(73)) and (inputs(112));
    layer0_outputs(1020) <= not((inputs(50)) and (inputs(160)));
    layer0_outputs(1021) <= '1';
    layer0_outputs(1022) <= not((inputs(0)) or (inputs(123)));
    layer0_outputs(1023) <= not((inputs(110)) or (inputs(229)));
    layer0_outputs(1024) <= '1';
    layer0_outputs(1025) <= '1';
    layer0_outputs(1026) <= not(inputs(13)) or (inputs(53));
    layer0_outputs(1027) <= not((inputs(96)) or (inputs(101)));
    layer0_outputs(1028) <= (inputs(235)) and (inputs(66));
    layer0_outputs(1029) <= '1';
    layer0_outputs(1030) <= (inputs(77)) or (inputs(106));
    layer0_outputs(1031) <= inputs(43);
    layer0_outputs(1032) <= '1';
    layer0_outputs(1033) <= (inputs(24)) and (inputs(75));
    layer0_outputs(1034) <= not(inputs(44)) or (inputs(115));
    layer0_outputs(1035) <= not(inputs(112));
    layer0_outputs(1036) <= inputs(114);
    layer0_outputs(1037) <= (inputs(118)) or (inputs(222));
    layer0_outputs(1038) <= (inputs(27)) and not (inputs(168));
    layer0_outputs(1039) <= '1';
    layer0_outputs(1040) <= '1';
    layer0_outputs(1041) <= inputs(111);
    layer0_outputs(1042) <= not(inputs(111)) or (inputs(240));
    layer0_outputs(1043) <= '0';
    layer0_outputs(1044) <= not(inputs(48)) or (inputs(101));
    layer0_outputs(1045) <= inputs(8);
    layer0_outputs(1046) <= not((inputs(12)) and (inputs(107)));
    layer0_outputs(1047) <= not(inputs(170)) or (inputs(48));
    layer0_outputs(1048) <= inputs(142);
    layer0_outputs(1049) <= (inputs(1)) or (inputs(144));
    layer0_outputs(1050) <= inputs(239);
    layer0_outputs(1051) <= not(inputs(33));
    layer0_outputs(1052) <= not(inputs(230)) or (inputs(143));
    layer0_outputs(1053) <= not(inputs(81));
    layer0_outputs(1054) <= not((inputs(18)) or (inputs(124)));
    layer0_outputs(1055) <= '1';
    layer0_outputs(1056) <= '1';
    layer0_outputs(1057) <= '0';
    layer0_outputs(1058) <= (inputs(13)) xor (inputs(250));
    layer0_outputs(1059) <= not(inputs(129)) or (inputs(28));
    layer0_outputs(1060) <= not((inputs(162)) or (inputs(122)));
    layer0_outputs(1061) <= inputs(163);
    layer0_outputs(1062) <= not((inputs(140)) and (inputs(244)));
    layer0_outputs(1063) <= (inputs(58)) and not (inputs(127));
    layer0_outputs(1064) <= (inputs(166)) or (inputs(237));
    layer0_outputs(1065) <= '0';
    layer0_outputs(1066) <= (inputs(157)) and not (inputs(18));
    layer0_outputs(1067) <= not(inputs(161)) or (inputs(139));
    layer0_outputs(1068) <= not(inputs(172));
    layer0_outputs(1069) <= '0';
    layer0_outputs(1070) <= '0';
    layer0_outputs(1071) <= not((inputs(206)) and (inputs(7)));
    layer0_outputs(1072) <= inputs(230);
    layer0_outputs(1073) <= inputs(150);
    layer0_outputs(1074) <= not(inputs(221));
    layer0_outputs(1075) <= '1';
    layer0_outputs(1076) <= (inputs(91)) and (inputs(159));
    layer0_outputs(1077) <= '0';
    layer0_outputs(1078) <= (inputs(122)) or (inputs(78));
    layer0_outputs(1079) <= '0';
    layer0_outputs(1080) <= '0';
    layer0_outputs(1081) <= '0';
    layer0_outputs(1082) <= (inputs(192)) or (inputs(211));
    layer0_outputs(1083) <= '1';
    layer0_outputs(1084) <= (inputs(180)) and (inputs(109));
    layer0_outputs(1085) <= (inputs(227)) or (inputs(9));
    layer0_outputs(1086) <= not(inputs(230));
    layer0_outputs(1087) <= (inputs(127)) and not (inputs(230));
    layer0_outputs(1088) <= not(inputs(125));
    layer0_outputs(1089) <= inputs(116);
    layer0_outputs(1090) <= '0';
    layer0_outputs(1091) <= inputs(160);
    layer0_outputs(1092) <= not((inputs(158)) or (inputs(240)));
    layer0_outputs(1093) <= (inputs(104)) and not (inputs(240));
    layer0_outputs(1094) <= (inputs(188)) xor (inputs(50));
    layer0_outputs(1095) <= (inputs(200)) xor (inputs(185));
    layer0_outputs(1096) <= '1';
    layer0_outputs(1097) <= not((inputs(207)) and (inputs(203)));
    layer0_outputs(1098) <= (inputs(66)) xor (inputs(146));
    layer0_outputs(1099) <= '1';
    layer0_outputs(1100) <= '0';
    layer0_outputs(1101) <= '0';
    layer0_outputs(1102) <= inputs(147);
    layer0_outputs(1103) <= '1';
    layer0_outputs(1104) <= '0';
    layer0_outputs(1105) <= (inputs(145)) and (inputs(56));
    layer0_outputs(1106) <= (inputs(33)) xor (inputs(146));
    layer0_outputs(1107) <= not(inputs(51)) or (inputs(203));
    layer0_outputs(1108) <= (inputs(58)) and not (inputs(135));
    layer0_outputs(1109) <= inputs(143);
    layer0_outputs(1110) <= '1';
    layer0_outputs(1111) <= not((inputs(74)) and (inputs(147)));
    layer0_outputs(1112) <= not(inputs(123)) or (inputs(55));
    layer0_outputs(1113) <= (inputs(156)) or (inputs(189));
    layer0_outputs(1114) <= not((inputs(0)) or (inputs(90)));
    layer0_outputs(1115) <= not(inputs(43));
    layer0_outputs(1116) <= '0';
    layer0_outputs(1117) <= inputs(95);
    layer0_outputs(1118) <= (inputs(83)) or (inputs(94));
    layer0_outputs(1119) <= '0';
    layer0_outputs(1120) <= not((inputs(243)) and (inputs(44)));
    layer0_outputs(1121) <= '0';
    layer0_outputs(1122) <= not((inputs(75)) or (inputs(132)));
    layer0_outputs(1123) <= not((inputs(15)) or (inputs(85)));
    layer0_outputs(1124) <= '0';
    layer0_outputs(1125) <= inputs(219);
    layer0_outputs(1126) <= inputs(99);
    layer0_outputs(1127) <= inputs(18);
    layer0_outputs(1128) <= inputs(130);
    layer0_outputs(1129) <= not(inputs(113)) or (inputs(13));
    layer0_outputs(1130) <= (inputs(87)) and not (inputs(221));
    layer0_outputs(1131) <= (inputs(69)) and not (inputs(167));
    layer0_outputs(1132) <= inputs(236);
    layer0_outputs(1133) <= '0';
    layer0_outputs(1134) <= not(inputs(103)) or (inputs(50));
    layer0_outputs(1135) <= not(inputs(178));
    layer0_outputs(1136) <= not(inputs(211)) or (inputs(42));
    layer0_outputs(1137) <= not((inputs(76)) and (inputs(43)));
    layer0_outputs(1138) <= '0';
    layer0_outputs(1139) <= not((inputs(26)) or (inputs(47)));
    layer0_outputs(1140) <= not((inputs(62)) or (inputs(96)));
    layer0_outputs(1141) <= inputs(9);
    layer0_outputs(1142) <= not(inputs(194));
    layer0_outputs(1143) <= '0';
    layer0_outputs(1144) <= (inputs(94)) and not (inputs(183));
    layer0_outputs(1145) <= inputs(254);
    layer0_outputs(1146) <= '1';
    layer0_outputs(1147) <= (inputs(35)) or (inputs(2));
    layer0_outputs(1148) <= '1';
    layer0_outputs(1149) <= (inputs(146)) xor (inputs(28));
    layer0_outputs(1150) <= inputs(77);
    layer0_outputs(1151) <= not(inputs(192));
    layer0_outputs(1152) <= (inputs(207)) and not (inputs(72));
    layer0_outputs(1153) <= '0';
    layer0_outputs(1154) <= not(inputs(15));
    layer0_outputs(1155) <= (inputs(74)) and not (inputs(188));
    layer0_outputs(1156) <= (inputs(58)) xor (inputs(218));
    layer0_outputs(1157) <= not(inputs(188)) or (inputs(198));
    layer0_outputs(1158) <= '1';
    layer0_outputs(1159) <= not(inputs(45)) or (inputs(75));
    layer0_outputs(1160) <= '0';
    layer0_outputs(1161) <= not(inputs(45));
    layer0_outputs(1162) <= '1';
    layer0_outputs(1163) <= not(inputs(34));
    layer0_outputs(1164) <= '0';
    layer0_outputs(1165) <= '1';
    layer0_outputs(1166) <= (inputs(80)) or (inputs(75));
    layer0_outputs(1167) <= '1';
    layer0_outputs(1168) <= not(inputs(216));
    layer0_outputs(1169) <= '1';
    layer0_outputs(1170) <= inputs(20);
    layer0_outputs(1171) <= '1';
    layer0_outputs(1172) <= (inputs(133)) and not (inputs(30));
    layer0_outputs(1173) <= not((inputs(74)) and (inputs(241)));
    layer0_outputs(1174) <= (inputs(70)) xor (inputs(102));
    layer0_outputs(1175) <= not(inputs(153));
    layer0_outputs(1176) <= (inputs(19)) and not (inputs(119));
    layer0_outputs(1177) <= not(inputs(8));
    layer0_outputs(1178) <= '1';
    layer0_outputs(1179) <= (inputs(143)) or (inputs(18));
    layer0_outputs(1180) <= not(inputs(173));
    layer0_outputs(1181) <= not((inputs(188)) xor (inputs(178)));
    layer0_outputs(1182) <= inputs(176);
    layer0_outputs(1183) <= '0';
    layer0_outputs(1184) <= not(inputs(121));
    layer0_outputs(1185) <= '1';
    layer0_outputs(1186) <= not(inputs(30));
    layer0_outputs(1187) <= inputs(220);
    layer0_outputs(1188) <= not((inputs(19)) and (inputs(24)));
    layer0_outputs(1189) <= not(inputs(212));
    layer0_outputs(1190) <= '1';
    layer0_outputs(1191) <= not((inputs(166)) or (inputs(121)));
    layer0_outputs(1192) <= not(inputs(204)) or (inputs(98));
    layer0_outputs(1193) <= '0';
    layer0_outputs(1194) <= (inputs(176)) or (inputs(76));
    layer0_outputs(1195) <= '1';
    layer0_outputs(1196) <= '1';
    layer0_outputs(1197) <= inputs(112);
    layer0_outputs(1198) <= (inputs(69)) and (inputs(210));
    layer0_outputs(1199) <= inputs(34);
    layer0_outputs(1200) <= not((inputs(227)) or (inputs(231)));
    layer0_outputs(1201) <= not((inputs(26)) or (inputs(10)));
    layer0_outputs(1202) <= not((inputs(200)) and (inputs(174)));
    layer0_outputs(1203) <= not(inputs(192)) or (inputs(12));
    layer0_outputs(1204) <= inputs(241);
    layer0_outputs(1205) <= not((inputs(172)) and (inputs(167)));
    layer0_outputs(1206) <= inputs(65);
    layer0_outputs(1207) <= '1';
    layer0_outputs(1208) <= not(inputs(234));
    layer0_outputs(1209) <= not(inputs(190));
    layer0_outputs(1210) <= not(inputs(29)) or (inputs(134));
    layer0_outputs(1211) <= not(inputs(30));
    layer0_outputs(1212) <= '1';
    layer0_outputs(1213) <= inputs(241);
    layer0_outputs(1214) <= '0';
    layer0_outputs(1215) <= not(inputs(191)) or (inputs(39));
    layer0_outputs(1216) <= (inputs(225)) and (inputs(53));
    layer0_outputs(1217) <= (inputs(152)) and not (inputs(136));
    layer0_outputs(1218) <= '0';
    layer0_outputs(1219) <= '1';
    layer0_outputs(1220) <= (inputs(101)) or (inputs(87));
    layer0_outputs(1221) <= not(inputs(24));
    layer0_outputs(1222) <= (inputs(241)) and not (inputs(153));
    layer0_outputs(1223) <= '0';
    layer0_outputs(1224) <= inputs(39);
    layer0_outputs(1225) <= '1';
    layer0_outputs(1226) <= '1';
    layer0_outputs(1227) <= not((inputs(238)) and (inputs(236)));
    layer0_outputs(1228) <= '0';
    layer0_outputs(1229) <= inputs(122);
    layer0_outputs(1230) <= inputs(110);
    layer0_outputs(1231) <= not(inputs(5));
    layer0_outputs(1232) <= '1';
    layer0_outputs(1233) <= (inputs(151)) and not (inputs(154));
    layer0_outputs(1234) <= inputs(207);
    layer0_outputs(1235) <= inputs(78);
    layer0_outputs(1236) <= '0';
    layer0_outputs(1237) <= '1';
    layer0_outputs(1238) <= (inputs(249)) and not (inputs(182));
    layer0_outputs(1239) <= (inputs(4)) and not (inputs(2));
    layer0_outputs(1240) <= inputs(180);
    layer0_outputs(1241) <= '1';
    layer0_outputs(1242) <= not(inputs(52)) or (inputs(171));
    layer0_outputs(1243) <= (inputs(200)) and (inputs(160));
    layer0_outputs(1244) <= (inputs(86)) and not (inputs(230));
    layer0_outputs(1245) <= not((inputs(249)) or (inputs(229)));
    layer0_outputs(1246) <= not(inputs(31));
    layer0_outputs(1247) <= (inputs(102)) or (inputs(84));
    layer0_outputs(1248) <= not((inputs(101)) and (inputs(201)));
    layer0_outputs(1249) <= not((inputs(18)) and (inputs(183)));
    layer0_outputs(1250) <= '1';
    layer0_outputs(1251) <= inputs(180);
    layer0_outputs(1252) <= not(inputs(166)) or (inputs(100));
    layer0_outputs(1253) <= not((inputs(217)) or (inputs(37)));
    layer0_outputs(1254) <= not(inputs(155)) or (inputs(113));
    layer0_outputs(1255) <= (inputs(147)) and (inputs(245));
    layer0_outputs(1256) <= inputs(60);
    layer0_outputs(1257) <= not((inputs(225)) or (inputs(127)));
    layer0_outputs(1258) <= '0';
    layer0_outputs(1259) <= (inputs(183)) and not (inputs(157));
    layer0_outputs(1260) <= inputs(63);
    layer0_outputs(1261) <= inputs(14);
    layer0_outputs(1262) <= inputs(91);
    layer0_outputs(1263) <= inputs(84);
    layer0_outputs(1264) <= inputs(213);
    layer0_outputs(1265) <= '0';
    layer0_outputs(1266) <= inputs(77);
    layer0_outputs(1267) <= not(inputs(81)) or (inputs(99));
    layer0_outputs(1268) <= (inputs(143)) or (inputs(208));
    layer0_outputs(1269) <= (inputs(12)) and not (inputs(189));
    layer0_outputs(1270) <= (inputs(7)) or (inputs(107));
    layer0_outputs(1271) <= (inputs(106)) or (inputs(241));
    layer0_outputs(1272) <= not(inputs(70)) or (inputs(151));
    layer0_outputs(1273) <= not(inputs(247)) or (inputs(68));
    layer0_outputs(1274) <= '0';
    layer0_outputs(1275) <= (inputs(15)) and (inputs(201));
    layer0_outputs(1276) <= '1';
    layer0_outputs(1277) <= not((inputs(48)) or (inputs(114)));
    layer0_outputs(1278) <= not(inputs(221)) or (inputs(50));
    layer0_outputs(1279) <= (inputs(80)) and not (inputs(142));
    layer0_outputs(1280) <= not(inputs(227)) or (inputs(39));
    layer0_outputs(1281) <= '1';
    layer0_outputs(1282) <= inputs(112);
    layer0_outputs(1283) <= '0';
    layer0_outputs(1284) <= inputs(20);
    layer0_outputs(1285) <= not((inputs(113)) xor (inputs(146)));
    layer0_outputs(1286) <= '0';
    layer0_outputs(1287) <= (inputs(111)) or (inputs(77));
    layer0_outputs(1288) <= not((inputs(84)) or (inputs(164)));
    layer0_outputs(1289) <= '0';
    layer0_outputs(1290) <= not((inputs(119)) and (inputs(176)));
    layer0_outputs(1291) <= not((inputs(184)) and (inputs(84)));
    layer0_outputs(1292) <= (inputs(132)) or (inputs(193));
    layer0_outputs(1293) <= (inputs(3)) and not (inputs(242));
    layer0_outputs(1294) <= not(inputs(71));
    layer0_outputs(1295) <= '0';
    layer0_outputs(1296) <= not(inputs(170)) or (inputs(106));
    layer0_outputs(1297) <= '0';
    layer0_outputs(1298) <= not(inputs(140)) or (inputs(122));
    layer0_outputs(1299) <= (inputs(0)) and (inputs(151));
    layer0_outputs(1300) <= not((inputs(167)) or (inputs(15)));
    layer0_outputs(1301) <= (inputs(250)) and (inputs(61));
    layer0_outputs(1302) <= (inputs(125)) and not (inputs(131));
    layer0_outputs(1303) <= inputs(84);
    layer0_outputs(1304) <= inputs(208);
    layer0_outputs(1305) <= not(inputs(217)) or (inputs(82));
    layer0_outputs(1306) <= not(inputs(33));
    layer0_outputs(1307) <= not(inputs(255));
    layer0_outputs(1308) <= '1';
    layer0_outputs(1309) <= not((inputs(188)) or (inputs(215)));
    layer0_outputs(1310) <= (inputs(72)) xor (inputs(204));
    layer0_outputs(1311) <= not(inputs(52)) or (inputs(108));
    layer0_outputs(1312) <= '0';
    layer0_outputs(1313) <= '1';
    layer0_outputs(1314) <= inputs(191);
    layer0_outputs(1315) <= (inputs(205)) and not (inputs(215));
    layer0_outputs(1316) <= (inputs(0)) and not (inputs(100));
    layer0_outputs(1317) <= '1';
    layer0_outputs(1318) <= not((inputs(88)) and (inputs(71)));
    layer0_outputs(1319) <= not(inputs(195)) or (inputs(132));
    layer0_outputs(1320) <= not((inputs(159)) and (inputs(249)));
    layer0_outputs(1321) <= not(inputs(23)) or (inputs(220));
    layer0_outputs(1322) <= (inputs(223)) and not (inputs(214));
    layer0_outputs(1323) <= not((inputs(21)) xor (inputs(65)));
    layer0_outputs(1324) <= not(inputs(189));
    layer0_outputs(1325) <= not((inputs(70)) xor (inputs(85)));
    layer0_outputs(1326) <= '1';
    layer0_outputs(1327) <= not((inputs(126)) or (inputs(103)));
    layer0_outputs(1328) <= not((inputs(3)) and (inputs(195)));
    layer0_outputs(1329) <= not(inputs(118));
    layer0_outputs(1330) <= not(inputs(193));
    layer0_outputs(1331) <= '1';
    layer0_outputs(1332) <= (inputs(139)) and not (inputs(142));
    layer0_outputs(1333) <= inputs(62);
    layer0_outputs(1334) <= (inputs(147)) and (inputs(104));
    layer0_outputs(1335) <= '1';
    layer0_outputs(1336) <= not(inputs(4)) or (inputs(173));
    layer0_outputs(1337) <= inputs(125);
    layer0_outputs(1338) <= '0';
    layer0_outputs(1339) <= not((inputs(221)) or (inputs(204)));
    layer0_outputs(1340) <= (inputs(88)) and not (inputs(45));
    layer0_outputs(1341) <= not((inputs(175)) xor (inputs(219)));
    layer0_outputs(1342) <= '0';
    layer0_outputs(1343) <= not(inputs(198)) or (inputs(254));
    layer0_outputs(1344) <= not((inputs(233)) or (inputs(187)));
    layer0_outputs(1345) <= inputs(190);
    layer0_outputs(1346) <= not(inputs(241));
    layer0_outputs(1347) <= not(inputs(137)) or (inputs(8));
    layer0_outputs(1348) <= '0';
    layer0_outputs(1349) <= not((inputs(55)) xor (inputs(192)));
    layer0_outputs(1350) <= (inputs(78)) and (inputs(30));
    layer0_outputs(1351) <= '0';
    layer0_outputs(1352) <= '1';
    layer0_outputs(1353) <= (inputs(116)) and not (inputs(228));
    layer0_outputs(1354) <= (inputs(214)) and not (inputs(201));
    layer0_outputs(1355) <= inputs(184);
    layer0_outputs(1356) <= (inputs(162)) and (inputs(202));
    layer0_outputs(1357) <= '0';
    layer0_outputs(1358) <= '1';
    layer0_outputs(1359) <= (inputs(77)) and (inputs(213));
    layer0_outputs(1360) <= not((inputs(194)) xor (inputs(44)));
    layer0_outputs(1361) <= inputs(128);
    layer0_outputs(1362) <= '1';
    layer0_outputs(1363) <= not(inputs(65)) or (inputs(0));
    layer0_outputs(1364) <= not((inputs(67)) and (inputs(123)));
    layer0_outputs(1365) <= (inputs(195)) and (inputs(79));
    layer0_outputs(1366) <= not(inputs(50)) or (inputs(177));
    layer0_outputs(1367) <= not((inputs(91)) or (inputs(38)));
    layer0_outputs(1368) <= (inputs(232)) and not (inputs(114));
    layer0_outputs(1369) <= not((inputs(2)) and (inputs(133)));
    layer0_outputs(1370) <= not(inputs(253)) or (inputs(115));
    layer0_outputs(1371) <= not((inputs(83)) or (inputs(223)));
    layer0_outputs(1372) <= not((inputs(133)) and (inputs(245)));
    layer0_outputs(1373) <= '1';
    layer0_outputs(1374) <= (inputs(146)) or (inputs(147));
    layer0_outputs(1375) <= inputs(75);
    layer0_outputs(1376) <= not(inputs(245));
    layer0_outputs(1377) <= inputs(17);
    layer0_outputs(1378) <= (inputs(6)) and not (inputs(164));
    layer0_outputs(1379) <= not((inputs(31)) xor (inputs(80)));
    layer0_outputs(1380) <= (inputs(29)) xor (inputs(229));
    layer0_outputs(1381) <= '1';
    layer0_outputs(1382) <= not((inputs(163)) or (inputs(173)));
    layer0_outputs(1383) <= (inputs(56)) and not (inputs(243));
    layer0_outputs(1384) <= not((inputs(209)) or (inputs(165)));
    layer0_outputs(1385) <= not(inputs(151));
    layer0_outputs(1386) <= inputs(158);
    layer0_outputs(1387) <= '1';
    layer0_outputs(1388) <= '1';
    layer0_outputs(1389) <= not((inputs(49)) and (inputs(161)));
    layer0_outputs(1390) <= not(inputs(228)) or (inputs(190));
    layer0_outputs(1391) <= '0';
    layer0_outputs(1392) <= '1';
    layer0_outputs(1393) <= not(inputs(41));
    layer0_outputs(1394) <= '1';
    layer0_outputs(1395) <= '1';
    layer0_outputs(1396) <= not((inputs(214)) or (inputs(234)));
    layer0_outputs(1397) <= (inputs(0)) and not (inputs(72));
    layer0_outputs(1398) <= '1';
    layer0_outputs(1399) <= '1';
    layer0_outputs(1400) <= (inputs(129)) and (inputs(31));
    layer0_outputs(1401) <= not(inputs(171));
    layer0_outputs(1402) <= not(inputs(91)) or (inputs(202));
    layer0_outputs(1403) <= '0';
    layer0_outputs(1404) <= '1';
    layer0_outputs(1405) <= inputs(20);
    layer0_outputs(1406) <= not(inputs(79));
    layer0_outputs(1407) <= (inputs(26)) and not (inputs(24));
    layer0_outputs(1408) <= inputs(3);
    layer0_outputs(1409) <= (inputs(157)) or (inputs(177));
    layer0_outputs(1410) <= not(inputs(97)) or (inputs(75));
    layer0_outputs(1411) <= inputs(222);
    layer0_outputs(1412) <= not(inputs(43)) or (inputs(41));
    layer0_outputs(1413) <= not(inputs(210));
    layer0_outputs(1414) <= (inputs(79)) xor (inputs(29));
    layer0_outputs(1415) <= inputs(223);
    layer0_outputs(1416) <= not((inputs(255)) or (inputs(117)));
    layer0_outputs(1417) <= (inputs(226)) and (inputs(191));
    layer0_outputs(1418) <= not((inputs(224)) and (inputs(44)));
    layer0_outputs(1419) <= not((inputs(6)) xor (inputs(41)));
    layer0_outputs(1420) <= '1';
    layer0_outputs(1421) <= not((inputs(36)) xor (inputs(239)));
    layer0_outputs(1422) <= inputs(60);
    layer0_outputs(1423) <= not(inputs(4)) or (inputs(97));
    layer0_outputs(1424) <= '0';
    layer0_outputs(1425) <= inputs(137);
    layer0_outputs(1426) <= '1';
    layer0_outputs(1427) <= not(inputs(204)) or (inputs(132));
    layer0_outputs(1428) <= (inputs(143)) and not (inputs(181));
    layer0_outputs(1429) <= not((inputs(193)) and (inputs(239)));
    layer0_outputs(1430) <= not((inputs(29)) and (inputs(172)));
    layer0_outputs(1431) <= not(inputs(188)) or (inputs(75));
    layer0_outputs(1432) <= '1';
    layer0_outputs(1433) <= '1';
    layer0_outputs(1434) <= (inputs(161)) and not (inputs(243));
    layer0_outputs(1435) <= inputs(177);
    layer0_outputs(1436) <= not(inputs(84));
    layer0_outputs(1437) <= not(inputs(119));
    layer0_outputs(1438) <= (inputs(204)) and not (inputs(202));
    layer0_outputs(1439) <= not((inputs(238)) and (inputs(125)));
    layer0_outputs(1440) <= inputs(239);
    layer0_outputs(1441) <= (inputs(117)) and (inputs(170));
    layer0_outputs(1442) <= not(inputs(59));
    layer0_outputs(1443) <= not(inputs(111)) or (inputs(131));
    layer0_outputs(1444) <= '1';
    layer0_outputs(1445) <= (inputs(98)) and not (inputs(163));
    layer0_outputs(1446) <= not((inputs(132)) or (inputs(130)));
    layer0_outputs(1447) <= (inputs(108)) or (inputs(214));
    layer0_outputs(1448) <= not((inputs(198)) or (inputs(177)));
    layer0_outputs(1449) <= not((inputs(23)) and (inputs(176)));
    layer0_outputs(1450) <= (inputs(252)) and (inputs(139));
    layer0_outputs(1451) <= '1';
    layer0_outputs(1452) <= (inputs(153)) and (inputs(134));
    layer0_outputs(1453) <= not(inputs(127)) or (inputs(219));
    layer0_outputs(1454) <= (inputs(65)) or (inputs(134));
    layer0_outputs(1455) <= '1';
    layer0_outputs(1456) <= '0';
    layer0_outputs(1457) <= not((inputs(246)) xor (inputs(224)));
    layer0_outputs(1458) <= not(inputs(163)) or (inputs(90));
    layer0_outputs(1459) <= (inputs(181)) and (inputs(98));
    layer0_outputs(1460) <= '1';
    layer0_outputs(1461) <= not(inputs(69)) or (inputs(238));
    layer0_outputs(1462) <= not(inputs(21)) or (inputs(212));
    layer0_outputs(1463) <= (inputs(194)) and (inputs(195));
    layer0_outputs(1464) <= inputs(247);
    layer0_outputs(1465) <= (inputs(238)) and (inputs(151));
    layer0_outputs(1466) <= (inputs(196)) and not (inputs(74));
    layer0_outputs(1467) <= '0';
    layer0_outputs(1468) <= '0';
    layer0_outputs(1469) <= inputs(62);
    layer0_outputs(1470) <= (inputs(0)) and not (inputs(171));
    layer0_outputs(1471) <= (inputs(147)) and (inputs(15));
    layer0_outputs(1472) <= (inputs(91)) and not (inputs(67));
    layer0_outputs(1473) <= (inputs(174)) and not (inputs(8));
    layer0_outputs(1474) <= not(inputs(0));
    layer0_outputs(1475) <= (inputs(112)) or (inputs(10));
    layer0_outputs(1476) <= not(inputs(75));
    layer0_outputs(1477) <= '0';
    layer0_outputs(1478) <= (inputs(192)) and not (inputs(177));
    layer0_outputs(1479) <= (inputs(123)) and not (inputs(231));
    layer0_outputs(1480) <= '0';
    layer0_outputs(1481) <= '0';
    layer0_outputs(1482) <= '0';
    layer0_outputs(1483) <= not((inputs(10)) or (inputs(162)));
    layer0_outputs(1484) <= not(inputs(98));
    layer0_outputs(1485) <= '1';
    layer0_outputs(1486) <= (inputs(211)) and not (inputs(162));
    layer0_outputs(1487) <= not((inputs(186)) or (inputs(153)));
    layer0_outputs(1488) <= (inputs(231)) and not (inputs(147));
    layer0_outputs(1489) <= not(inputs(205)) or (inputs(138));
    layer0_outputs(1490) <= (inputs(233)) and not (inputs(98));
    layer0_outputs(1491) <= inputs(194);
    layer0_outputs(1492) <= inputs(97);
    layer0_outputs(1493) <= (inputs(108)) xor (inputs(121));
    layer0_outputs(1494) <= not((inputs(22)) or (inputs(187)));
    layer0_outputs(1495) <= (inputs(239)) or (inputs(35));
    layer0_outputs(1496) <= not((inputs(92)) or (inputs(77)));
    layer0_outputs(1497) <= inputs(162);
    layer0_outputs(1498) <= (inputs(159)) and not (inputs(212));
    layer0_outputs(1499) <= '0';
    layer0_outputs(1500) <= not(inputs(65)) or (inputs(46));
    layer0_outputs(1501) <= not(inputs(144)) or (inputs(255));
    layer0_outputs(1502) <= not(inputs(124)) or (inputs(73));
    layer0_outputs(1503) <= (inputs(250)) or (inputs(33));
    layer0_outputs(1504) <= (inputs(90)) xor (inputs(47));
    layer0_outputs(1505) <= (inputs(0)) and (inputs(97));
    layer0_outputs(1506) <= '0';
    layer0_outputs(1507) <= '1';
    layer0_outputs(1508) <= (inputs(31)) and not (inputs(77));
    layer0_outputs(1509) <= not(inputs(127)) or (inputs(48));
    layer0_outputs(1510) <= (inputs(51)) or (inputs(134));
    layer0_outputs(1511) <= not((inputs(93)) and (inputs(208)));
    layer0_outputs(1512) <= not(inputs(208)) or (inputs(110));
    layer0_outputs(1513) <= not(inputs(60)) or (inputs(197));
    layer0_outputs(1514) <= not(inputs(142));
    layer0_outputs(1515) <= (inputs(60)) and not (inputs(46));
    layer0_outputs(1516) <= '0';
    layer0_outputs(1517) <= inputs(139);
    layer0_outputs(1518) <= not(inputs(47));
    layer0_outputs(1519) <= '0';
    layer0_outputs(1520) <= not(inputs(115));
    layer0_outputs(1521) <= not((inputs(136)) and (inputs(128)));
    layer0_outputs(1522) <= not((inputs(83)) or (inputs(42)));
    layer0_outputs(1523) <= not((inputs(138)) or (inputs(234)));
    layer0_outputs(1524) <= '0';
    layer0_outputs(1525) <= (inputs(91)) and not (inputs(173));
    layer0_outputs(1526) <= not(inputs(167));
    layer0_outputs(1527) <= (inputs(213)) and not (inputs(220));
    layer0_outputs(1528) <= not(inputs(237)) or (inputs(162));
    layer0_outputs(1529) <= '0';
    layer0_outputs(1530) <= (inputs(205)) and (inputs(71));
    layer0_outputs(1531) <= (inputs(117)) or (inputs(205));
    layer0_outputs(1532) <= inputs(220);
    layer0_outputs(1533) <= '1';
    layer0_outputs(1534) <= '0';
    layer0_outputs(1535) <= not((inputs(223)) and (inputs(135)));
    layer0_outputs(1536) <= not(inputs(191));
    layer0_outputs(1537) <= inputs(119);
    layer0_outputs(1538) <= not(inputs(101)) or (inputs(5));
    layer0_outputs(1539) <= not(inputs(4)) or (inputs(24));
    layer0_outputs(1540) <= inputs(16);
    layer0_outputs(1541) <= '0';
    layer0_outputs(1542) <= (inputs(251)) and (inputs(50));
    layer0_outputs(1543) <= (inputs(183)) or (inputs(45));
    layer0_outputs(1544) <= '0';
    layer0_outputs(1545) <= not((inputs(254)) xor (inputs(82)));
    layer0_outputs(1546) <= not((inputs(21)) xor (inputs(238)));
    layer0_outputs(1547) <= not(inputs(102)) or (inputs(160));
    layer0_outputs(1548) <= '1';
    layer0_outputs(1549) <= inputs(171);
    layer0_outputs(1550) <= (inputs(136)) and (inputs(209));
    layer0_outputs(1551) <= (inputs(205)) and not (inputs(52));
    layer0_outputs(1552) <= '1';
    layer0_outputs(1553) <= not((inputs(134)) and (inputs(161)));
    layer0_outputs(1554) <= not(inputs(117));
    layer0_outputs(1555) <= '1';
    layer0_outputs(1556) <= (inputs(13)) and (inputs(130));
    layer0_outputs(1557) <= (inputs(181)) and not (inputs(11));
    layer0_outputs(1558) <= (inputs(140)) and not (inputs(216));
    layer0_outputs(1559) <= (inputs(255)) and (inputs(1));
    layer0_outputs(1560) <= not(inputs(117)) or (inputs(15));
    layer0_outputs(1561) <= '1';
    layer0_outputs(1562) <= not((inputs(38)) or (inputs(158)));
    layer0_outputs(1563) <= (inputs(120)) and not (inputs(14));
    layer0_outputs(1564) <= not(inputs(74)) or (inputs(231));
    layer0_outputs(1565) <= not((inputs(141)) xor (inputs(79)));
    layer0_outputs(1566) <= (inputs(39)) or (inputs(197));
    layer0_outputs(1567) <= '0';
    layer0_outputs(1568) <= '0';
    layer0_outputs(1569) <= not(inputs(86));
    layer0_outputs(1570) <= '1';
    layer0_outputs(1571) <= inputs(221);
    layer0_outputs(1572) <= '0';
    layer0_outputs(1573) <= '0';
    layer0_outputs(1574) <= '1';
    layer0_outputs(1575) <= not((inputs(95)) and (inputs(91)));
    layer0_outputs(1576) <= not(inputs(233));
    layer0_outputs(1577) <= not(inputs(117)) or (inputs(187));
    layer0_outputs(1578) <= (inputs(234)) and not (inputs(58));
    layer0_outputs(1579) <= '0';
    layer0_outputs(1580) <= (inputs(7)) and (inputs(127));
    layer0_outputs(1581) <= '0';
    layer0_outputs(1582) <= '0';
    layer0_outputs(1583) <= '0';
    layer0_outputs(1584) <= not((inputs(162)) or (inputs(126)));
    layer0_outputs(1585) <= inputs(143);
    layer0_outputs(1586) <= '0';
    layer0_outputs(1587) <= not(inputs(162)) or (inputs(171));
    layer0_outputs(1588) <= '0';
    layer0_outputs(1589) <= inputs(37);
    layer0_outputs(1590) <= not(inputs(132)) or (inputs(42));
    layer0_outputs(1591) <= inputs(114);
    layer0_outputs(1592) <= not((inputs(126)) or (inputs(129)));
    layer0_outputs(1593) <= not(inputs(167)) or (inputs(113));
    layer0_outputs(1594) <= not(inputs(175)) or (inputs(59));
    layer0_outputs(1595) <= not(inputs(126));
    layer0_outputs(1596) <= inputs(30);
    layer0_outputs(1597) <= inputs(144);
    layer0_outputs(1598) <= not(inputs(23)) or (inputs(194));
    layer0_outputs(1599) <= '1';
    layer0_outputs(1600) <= '0';
    layer0_outputs(1601) <= not(inputs(19));
    layer0_outputs(1602) <= inputs(253);
    layer0_outputs(1603) <= not(inputs(127)) or (inputs(237));
    layer0_outputs(1604) <= not(inputs(33));
    layer0_outputs(1605) <= '0';
    layer0_outputs(1606) <= '0';
    layer0_outputs(1607) <= (inputs(150)) and not (inputs(7));
    layer0_outputs(1608) <= '1';
    layer0_outputs(1609) <= not(inputs(247)) or (inputs(19));
    layer0_outputs(1610) <= (inputs(21)) or (inputs(11));
    layer0_outputs(1611) <= not((inputs(158)) and (inputs(158)));
    layer0_outputs(1612) <= '0';
    layer0_outputs(1613) <= not((inputs(59)) and (inputs(100)));
    layer0_outputs(1614) <= not(inputs(79)) or (inputs(144));
    layer0_outputs(1615) <= not((inputs(236)) and (inputs(215)));
    layer0_outputs(1616) <= '0';
    layer0_outputs(1617) <= not(inputs(113));
    layer0_outputs(1618) <= '0';
    layer0_outputs(1619) <= not(inputs(88)) or (inputs(64));
    layer0_outputs(1620) <= not(inputs(149)) or (inputs(221));
    layer0_outputs(1621) <= (inputs(180)) or (inputs(117));
    layer0_outputs(1622) <= (inputs(56)) and not (inputs(188));
    layer0_outputs(1623) <= (inputs(215)) and not (inputs(183));
    layer0_outputs(1624) <= (inputs(106)) and not (inputs(82));
    layer0_outputs(1625) <= not((inputs(86)) xor (inputs(161)));
    layer0_outputs(1626) <= not(inputs(255));
    layer0_outputs(1627) <= not(inputs(53)) or (inputs(210));
    layer0_outputs(1628) <= '1';
    layer0_outputs(1629) <= '1';
    layer0_outputs(1630) <= not(inputs(106));
    layer0_outputs(1631) <= not(inputs(130));
    layer0_outputs(1632) <= not(inputs(229));
    layer0_outputs(1633) <= inputs(110);
    layer0_outputs(1634) <= '1';
    layer0_outputs(1635) <= not((inputs(181)) and (inputs(222)));
    layer0_outputs(1636) <= not(inputs(139)) or (inputs(220));
    layer0_outputs(1637) <= (inputs(115)) and not (inputs(19));
    layer0_outputs(1638) <= '1';
    layer0_outputs(1639) <= not(inputs(43)) or (inputs(223));
    layer0_outputs(1640) <= (inputs(121)) and not (inputs(24));
    layer0_outputs(1641) <= (inputs(22)) and (inputs(87));
    layer0_outputs(1642) <= inputs(185);
    layer0_outputs(1643) <= not((inputs(27)) or (inputs(115)));
    layer0_outputs(1644) <= (inputs(14)) and not (inputs(125));
    layer0_outputs(1645) <= not(inputs(163)) or (inputs(191));
    layer0_outputs(1646) <= not(inputs(114));
    layer0_outputs(1647) <= (inputs(61)) and (inputs(75));
    layer0_outputs(1648) <= not(inputs(112)) or (inputs(139));
    layer0_outputs(1649) <= (inputs(168)) or (inputs(56));
    layer0_outputs(1650) <= (inputs(50)) and not (inputs(125));
    layer0_outputs(1651) <= (inputs(71)) and not (inputs(201));
    layer0_outputs(1652) <= '1';
    layer0_outputs(1653) <= not((inputs(209)) and (inputs(209)));
    layer0_outputs(1654) <= '1';
    layer0_outputs(1655) <= not((inputs(80)) and (inputs(187)));
    layer0_outputs(1656) <= '0';
    layer0_outputs(1657) <= '1';
    layer0_outputs(1658) <= not(inputs(118));
    layer0_outputs(1659) <= (inputs(225)) and not (inputs(220));
    layer0_outputs(1660) <= not(inputs(153));
    layer0_outputs(1661) <= not((inputs(188)) and (inputs(75)));
    layer0_outputs(1662) <= inputs(50);
    layer0_outputs(1663) <= not(inputs(140)) or (inputs(20));
    layer0_outputs(1664) <= not(inputs(47)) or (inputs(89));
    layer0_outputs(1665) <= not((inputs(224)) or (inputs(114)));
    layer0_outputs(1666) <= '0';
    layer0_outputs(1667) <= not((inputs(113)) or (inputs(112)));
    layer0_outputs(1668) <= not((inputs(104)) or (inputs(84)));
    layer0_outputs(1669) <= not(inputs(119));
    layer0_outputs(1670) <= not(inputs(238)) or (inputs(205));
    layer0_outputs(1671) <= inputs(101);
    layer0_outputs(1672) <= inputs(149);
    layer0_outputs(1673) <= '1';
    layer0_outputs(1674) <= (inputs(179)) and (inputs(25));
    layer0_outputs(1675) <= '0';
    layer0_outputs(1676) <= not((inputs(194)) xor (inputs(207)));
    layer0_outputs(1677) <= (inputs(150)) or (inputs(57));
    layer0_outputs(1678) <= '0';
    layer0_outputs(1679) <= not((inputs(120)) and (inputs(241)));
    layer0_outputs(1680) <= not(inputs(64)) or (inputs(50));
    layer0_outputs(1681) <= '1';
    layer0_outputs(1682) <= inputs(208);
    layer0_outputs(1683) <= not((inputs(160)) and (inputs(252)));
    layer0_outputs(1684) <= (inputs(205)) and not (inputs(191));
    layer0_outputs(1685) <= '1';
    layer0_outputs(1686) <= inputs(217);
    layer0_outputs(1687) <= (inputs(72)) or (inputs(121));
    layer0_outputs(1688) <= '0';
    layer0_outputs(1689) <= inputs(29);
    layer0_outputs(1690) <= '1';
    layer0_outputs(1691) <= not(inputs(224)) or (inputs(164));
    layer0_outputs(1692) <= not(inputs(55)) or (inputs(29));
    layer0_outputs(1693) <= inputs(228);
    layer0_outputs(1694) <= '0';
    layer0_outputs(1695) <= '1';
    layer0_outputs(1696) <= inputs(130);
    layer0_outputs(1697) <= inputs(78);
    layer0_outputs(1698) <= (inputs(93)) and not (inputs(107));
    layer0_outputs(1699) <= (inputs(161)) and not (inputs(139));
    layer0_outputs(1700) <= not(inputs(35)) or (inputs(37));
    layer0_outputs(1701) <= not((inputs(92)) and (inputs(116)));
    layer0_outputs(1702) <= not(inputs(49));
    layer0_outputs(1703) <= (inputs(32)) and not (inputs(154));
    layer0_outputs(1704) <= (inputs(80)) and not (inputs(115));
    layer0_outputs(1705) <= '0';
    layer0_outputs(1706) <= not(inputs(45));
    layer0_outputs(1707) <= (inputs(168)) xor (inputs(79));
    layer0_outputs(1708) <= (inputs(246)) and not (inputs(58));
    layer0_outputs(1709) <= (inputs(144)) or (inputs(151));
    layer0_outputs(1710) <= (inputs(54)) and not (inputs(206));
    layer0_outputs(1711) <= not(inputs(66));
    layer0_outputs(1712) <= not(inputs(112));
    layer0_outputs(1713) <= '0';
    layer0_outputs(1714) <= (inputs(27)) and (inputs(68));
    layer0_outputs(1715) <= inputs(25);
    layer0_outputs(1716) <= '0';
    layer0_outputs(1717) <= '1';
    layer0_outputs(1718) <= not(inputs(197));
    layer0_outputs(1719) <= '0';
    layer0_outputs(1720) <= '1';
    layer0_outputs(1721) <= not(inputs(179));
    layer0_outputs(1722) <= not(inputs(149)) or (inputs(192));
    layer0_outputs(1723) <= not(inputs(133));
    layer0_outputs(1724) <= not((inputs(242)) and (inputs(121)));
    layer0_outputs(1725) <= (inputs(198)) or (inputs(233));
    layer0_outputs(1726) <= '1';
    layer0_outputs(1727) <= not(inputs(65));
    layer0_outputs(1728) <= '1';
    layer0_outputs(1729) <= inputs(85);
    layer0_outputs(1730) <= (inputs(153)) and not (inputs(242));
    layer0_outputs(1731) <= '0';
    layer0_outputs(1732) <= '0';
    layer0_outputs(1733) <= inputs(231);
    layer0_outputs(1734) <= not(inputs(111)) or (inputs(140));
    layer0_outputs(1735) <= (inputs(219)) and (inputs(46));
    layer0_outputs(1736) <= '1';
    layer0_outputs(1737) <= '1';
    layer0_outputs(1738) <= not(inputs(213)) or (inputs(50));
    layer0_outputs(1739) <= inputs(216);
    layer0_outputs(1740) <= (inputs(224)) or (inputs(225));
    layer0_outputs(1741) <= '0';
    layer0_outputs(1742) <= not(inputs(113));
    layer0_outputs(1743) <= (inputs(104)) and not (inputs(75));
    layer0_outputs(1744) <= inputs(48);
    layer0_outputs(1745) <= inputs(135);
    layer0_outputs(1746) <= '1';
    layer0_outputs(1747) <= '0';
    layer0_outputs(1748) <= '1';
    layer0_outputs(1749) <= (inputs(70)) or (inputs(53));
    layer0_outputs(1750) <= '1';
    layer0_outputs(1751) <= inputs(18);
    layer0_outputs(1752) <= not(inputs(190)) or (inputs(72));
    layer0_outputs(1753) <= not(inputs(103));
    layer0_outputs(1754) <= not(inputs(78)) or (inputs(15));
    layer0_outputs(1755) <= inputs(3);
    layer0_outputs(1756) <= '0';
    layer0_outputs(1757) <= '0';
    layer0_outputs(1758) <= not((inputs(100)) and (inputs(92)));
    layer0_outputs(1759) <= not(inputs(148));
    layer0_outputs(1760) <= (inputs(199)) and (inputs(218));
    layer0_outputs(1761) <= not(inputs(77));
    layer0_outputs(1762) <= not(inputs(178)) or (inputs(205));
    layer0_outputs(1763) <= not((inputs(38)) or (inputs(104)));
    layer0_outputs(1764) <= '1';
    layer0_outputs(1765) <= not((inputs(99)) and (inputs(238)));
    layer0_outputs(1766) <= not(inputs(234)) or (inputs(24));
    layer0_outputs(1767) <= not(inputs(111)) or (inputs(110));
    layer0_outputs(1768) <= not(inputs(117));
    layer0_outputs(1769) <= '1';
    layer0_outputs(1770) <= (inputs(40)) xor (inputs(9));
    layer0_outputs(1771) <= (inputs(149)) and not (inputs(133));
    layer0_outputs(1772) <= not(inputs(132)) or (inputs(21));
    layer0_outputs(1773) <= not(inputs(45)) or (inputs(211));
    layer0_outputs(1774) <= not(inputs(191));
    layer0_outputs(1775) <= not(inputs(223));
    layer0_outputs(1776) <= '1';
    layer0_outputs(1777) <= '1';
    layer0_outputs(1778) <= (inputs(226)) and (inputs(126));
    layer0_outputs(1779) <= not(inputs(57));
    layer0_outputs(1780) <= inputs(71);
    layer0_outputs(1781) <= inputs(1);
    layer0_outputs(1782) <= not(inputs(144));
    layer0_outputs(1783) <= (inputs(15)) or (inputs(99));
    layer0_outputs(1784) <= inputs(1);
    layer0_outputs(1785) <= (inputs(168)) or (inputs(163));
    layer0_outputs(1786) <= (inputs(1)) and not (inputs(249));
    layer0_outputs(1787) <= '0';
    layer0_outputs(1788) <= not(inputs(152)) or (inputs(225));
    layer0_outputs(1789) <= '1';
    layer0_outputs(1790) <= not(inputs(128));
    layer0_outputs(1791) <= not((inputs(94)) and (inputs(251)));
    layer0_outputs(1792) <= '1';
    layer0_outputs(1793) <= not(inputs(53));
    layer0_outputs(1794) <= '1';
    layer0_outputs(1795) <= inputs(52);
    layer0_outputs(1796) <= not(inputs(92));
    layer0_outputs(1797) <= (inputs(114)) and not (inputs(248));
    layer0_outputs(1798) <= (inputs(205)) or (inputs(16));
    layer0_outputs(1799) <= inputs(98);
    layer0_outputs(1800) <= inputs(3);
    layer0_outputs(1801) <= (inputs(43)) or (inputs(36));
    layer0_outputs(1802) <= inputs(179);
    layer0_outputs(1803) <= not(inputs(153));
    layer0_outputs(1804) <= '1';
    layer0_outputs(1805) <= '1';
    layer0_outputs(1806) <= '0';
    layer0_outputs(1807) <= inputs(56);
    layer0_outputs(1808) <= not(inputs(63));
    layer0_outputs(1809) <= '1';
    layer0_outputs(1810) <= (inputs(109)) and (inputs(239));
    layer0_outputs(1811) <= (inputs(219)) or (inputs(160));
    layer0_outputs(1812) <= not(inputs(59)) or (inputs(117));
    layer0_outputs(1813) <= '1';
    layer0_outputs(1814) <= '0';
    layer0_outputs(1815) <= not(inputs(26)) or (inputs(90));
    layer0_outputs(1816) <= not(inputs(239));
    layer0_outputs(1817) <= (inputs(138)) and not (inputs(241));
    layer0_outputs(1818) <= not(inputs(239));
    layer0_outputs(1819) <= not(inputs(218));
    layer0_outputs(1820) <= not((inputs(38)) and (inputs(240)));
    layer0_outputs(1821) <= not((inputs(85)) and (inputs(134)));
    layer0_outputs(1822) <= inputs(164);
    layer0_outputs(1823) <= not((inputs(211)) and (inputs(45)));
    layer0_outputs(1824) <= '0';
    layer0_outputs(1825) <= not(inputs(198));
    layer0_outputs(1826) <= not(inputs(167));
    layer0_outputs(1827) <= not(inputs(99));
    layer0_outputs(1828) <= not(inputs(242));
    layer0_outputs(1829) <= (inputs(120)) and (inputs(8));
    layer0_outputs(1830) <= '1';
    layer0_outputs(1831) <= inputs(113);
    layer0_outputs(1832) <= not((inputs(248)) or (inputs(41)));
    layer0_outputs(1833) <= '0';
    layer0_outputs(1834) <= not(inputs(33)) or (inputs(155));
    layer0_outputs(1835) <= (inputs(113)) and not (inputs(202));
    layer0_outputs(1836) <= (inputs(100)) and (inputs(153));
    layer0_outputs(1837) <= (inputs(63)) or (inputs(237));
    layer0_outputs(1838) <= inputs(191);
    layer0_outputs(1839) <= not(inputs(200));
    layer0_outputs(1840) <= inputs(160);
    layer0_outputs(1841) <= (inputs(253)) or (inputs(238));
    layer0_outputs(1842) <= '1';
    layer0_outputs(1843) <= (inputs(120)) and (inputs(70));
    layer0_outputs(1844) <= not(inputs(28)) or (inputs(171));
    layer0_outputs(1845) <= not(inputs(238)) or (inputs(167));
    layer0_outputs(1846) <= '0';
    layer0_outputs(1847) <= '0';
    layer0_outputs(1848) <= inputs(228);
    layer0_outputs(1849) <= (inputs(22)) and not (inputs(247));
    layer0_outputs(1850) <= not(inputs(75));
    layer0_outputs(1851) <= '0';
    layer0_outputs(1852) <= '1';
    layer0_outputs(1853) <= '0';
    layer0_outputs(1854) <= '1';
    layer0_outputs(1855) <= inputs(219);
    layer0_outputs(1856) <= '1';
    layer0_outputs(1857) <= not((inputs(141)) and (inputs(69)));
    layer0_outputs(1858) <= '1';
    layer0_outputs(1859) <= not(inputs(56));
    layer0_outputs(1860) <= not(inputs(159));
    layer0_outputs(1861) <= not(inputs(69)) or (inputs(22));
    layer0_outputs(1862) <= not(inputs(201));
    layer0_outputs(1863) <= (inputs(148)) and not (inputs(227));
    layer0_outputs(1864) <= inputs(164);
    layer0_outputs(1865) <= inputs(190);
    layer0_outputs(1866) <= inputs(182);
    layer0_outputs(1867) <= not(inputs(103)) or (inputs(175));
    layer0_outputs(1868) <= not(inputs(198)) or (inputs(121));
    layer0_outputs(1869) <= inputs(54);
    layer0_outputs(1870) <= (inputs(125)) and (inputs(199));
    layer0_outputs(1871) <= inputs(80);
    layer0_outputs(1872) <= '1';
    layer0_outputs(1873) <= '1';
    layer0_outputs(1874) <= not(inputs(142)) or (inputs(219));
    layer0_outputs(1875) <= not((inputs(65)) and (inputs(14)));
    layer0_outputs(1876) <= inputs(20);
    layer0_outputs(1877) <= not(inputs(35)) or (inputs(55));
    layer0_outputs(1878) <= inputs(146);
    layer0_outputs(1879) <= '1';
    layer0_outputs(1880) <= (inputs(39)) and not (inputs(203));
    layer0_outputs(1881) <= (inputs(102)) or (inputs(212));
    layer0_outputs(1882) <= not(inputs(69));
    layer0_outputs(1883) <= not(inputs(12)) or (inputs(133));
    layer0_outputs(1884) <= not((inputs(3)) or (inputs(135)));
    layer0_outputs(1885) <= not((inputs(10)) or (inputs(114)));
    layer0_outputs(1886) <= not(inputs(110)) or (inputs(125));
    layer0_outputs(1887) <= (inputs(14)) or (inputs(123));
    layer0_outputs(1888) <= '1';
    layer0_outputs(1889) <= (inputs(249)) and not (inputs(74));
    layer0_outputs(1890) <= inputs(117);
    layer0_outputs(1891) <= '0';
    layer0_outputs(1892) <= '0';
    layer0_outputs(1893) <= not(inputs(174)) or (inputs(11));
    layer0_outputs(1894) <= '0';
    layer0_outputs(1895) <= not(inputs(11));
    layer0_outputs(1896) <= (inputs(106)) and not (inputs(245));
    layer0_outputs(1897) <= inputs(11);
    layer0_outputs(1898) <= inputs(119);
    layer0_outputs(1899) <= '0';
    layer0_outputs(1900) <= inputs(226);
    layer0_outputs(1901) <= '1';
    layer0_outputs(1902) <= not(inputs(182));
    layer0_outputs(1903) <= '0';
    layer0_outputs(1904) <= (inputs(133)) and not (inputs(190));
    layer0_outputs(1905) <= not(inputs(145)) or (inputs(190));
    layer0_outputs(1906) <= inputs(123);
    layer0_outputs(1907) <= not(inputs(112));
    layer0_outputs(1908) <= '1';
    layer0_outputs(1909) <= '1';
    layer0_outputs(1910) <= '0';
    layer0_outputs(1911) <= inputs(161);
    layer0_outputs(1912) <= (inputs(113)) or (inputs(98));
    layer0_outputs(1913) <= (inputs(107)) or (inputs(55));
    layer0_outputs(1914) <= (inputs(22)) and not (inputs(3));
    layer0_outputs(1915) <= '1';
    layer0_outputs(1916) <= '1';
    layer0_outputs(1917) <= not(inputs(212));
    layer0_outputs(1918) <= not((inputs(204)) and (inputs(28)));
    layer0_outputs(1919) <= (inputs(7)) and (inputs(141));
    layer0_outputs(1920) <= not(inputs(33)) or (inputs(111));
    layer0_outputs(1921) <= not(inputs(176)) or (inputs(3));
    layer0_outputs(1922) <= '0';
    layer0_outputs(1923) <= not((inputs(43)) and (inputs(234)));
    layer0_outputs(1924) <= '1';
    layer0_outputs(1925) <= (inputs(208)) and not (inputs(11));
    layer0_outputs(1926) <= '0';
    layer0_outputs(1927) <= (inputs(49)) and not (inputs(159));
    layer0_outputs(1928) <= inputs(232);
    layer0_outputs(1929) <= not((inputs(111)) xor (inputs(241)));
    layer0_outputs(1930) <= not((inputs(86)) or (inputs(177)));
    layer0_outputs(1931) <= '1';
    layer0_outputs(1932) <= inputs(79);
    layer0_outputs(1933) <= inputs(101);
    layer0_outputs(1934) <= (inputs(34)) and not (inputs(73));
    layer0_outputs(1935) <= '1';
    layer0_outputs(1936) <= '1';
    layer0_outputs(1937) <= not(inputs(121));
    layer0_outputs(1938) <= inputs(177);
    layer0_outputs(1939) <= (inputs(236)) and not (inputs(154));
    layer0_outputs(1940) <= '0';
    layer0_outputs(1941) <= not((inputs(63)) or (inputs(229)));
    layer0_outputs(1942) <= '1';
    layer0_outputs(1943) <= not(inputs(76));
    layer0_outputs(1944) <= not((inputs(155)) or (inputs(7)));
    layer0_outputs(1945) <= not(inputs(244));
    layer0_outputs(1946) <= '0';
    layer0_outputs(1947) <= inputs(116);
    layer0_outputs(1948) <= not(inputs(120));
    layer0_outputs(1949) <= (inputs(178)) and not (inputs(228));
    layer0_outputs(1950) <= (inputs(45)) and not (inputs(137));
    layer0_outputs(1951) <= '1';
    layer0_outputs(1952) <= '0';
    layer0_outputs(1953) <= not((inputs(114)) or (inputs(40)));
    layer0_outputs(1954) <= inputs(115);
    layer0_outputs(1955) <= inputs(19);
    layer0_outputs(1956) <= (inputs(163)) xor (inputs(95));
    layer0_outputs(1957) <= inputs(176);
    layer0_outputs(1958) <= (inputs(167)) and (inputs(19));
    layer0_outputs(1959) <= not(inputs(98));
    layer0_outputs(1960) <= '0';
    layer0_outputs(1961) <= not((inputs(48)) xor (inputs(235)));
    layer0_outputs(1962) <= '0';
    layer0_outputs(1963) <= '0';
    layer0_outputs(1964) <= (inputs(173)) and not (inputs(4));
    layer0_outputs(1965) <= inputs(220);
    layer0_outputs(1966) <= (inputs(57)) or (inputs(231));
    layer0_outputs(1967) <= not(inputs(21)) or (inputs(137));
    layer0_outputs(1968) <= (inputs(82)) and (inputs(237));
    layer0_outputs(1969) <= '0';
    layer0_outputs(1970) <= inputs(249);
    layer0_outputs(1971) <= inputs(40);
    layer0_outputs(1972) <= not((inputs(160)) and (inputs(128)));
    layer0_outputs(1973) <= not(inputs(14)) or (inputs(26));
    layer0_outputs(1974) <= (inputs(173)) and (inputs(251));
    layer0_outputs(1975) <= inputs(130);
    layer0_outputs(1976) <= (inputs(232)) and not (inputs(96));
    layer0_outputs(1977) <= not(inputs(148));
    layer0_outputs(1978) <= '1';
    layer0_outputs(1979) <= '0';
    layer0_outputs(1980) <= not(inputs(78)) or (inputs(210));
    layer0_outputs(1981) <= inputs(234);
    layer0_outputs(1982) <= not((inputs(98)) and (inputs(57)));
    layer0_outputs(1983) <= (inputs(207)) and (inputs(241));
    layer0_outputs(1984) <= not((inputs(239)) and (inputs(111)));
    layer0_outputs(1985) <= inputs(179);
    layer0_outputs(1986) <= not(inputs(96)) or (inputs(108));
    layer0_outputs(1987) <= '0';
    layer0_outputs(1988) <= not(inputs(146));
    layer0_outputs(1989) <= (inputs(57)) and not (inputs(199));
    layer0_outputs(1990) <= not((inputs(22)) or (inputs(225)));
    layer0_outputs(1991) <= '1';
    layer0_outputs(1992) <= (inputs(254)) and (inputs(155));
    layer0_outputs(1993) <= '1';
    layer0_outputs(1994) <= '0';
    layer0_outputs(1995) <= (inputs(86)) and not (inputs(217));
    layer0_outputs(1996) <= not(inputs(254));
    layer0_outputs(1997) <= not((inputs(36)) and (inputs(124)));
    layer0_outputs(1998) <= not(inputs(250));
    layer0_outputs(1999) <= '0';
    layer0_outputs(2000) <= not((inputs(218)) and (inputs(189)));
    layer0_outputs(2001) <= inputs(185);
    layer0_outputs(2002) <= not(inputs(58));
    layer0_outputs(2003) <= not((inputs(116)) or (inputs(42)));
    layer0_outputs(2004) <= '0';
    layer0_outputs(2005) <= not((inputs(112)) xor (inputs(82)));
    layer0_outputs(2006) <= not(inputs(175)) or (inputs(110));
    layer0_outputs(2007) <= '0';
    layer0_outputs(2008) <= inputs(9);
    layer0_outputs(2009) <= '1';
    layer0_outputs(2010) <= '1';
    layer0_outputs(2011) <= '0';
    layer0_outputs(2012) <= (inputs(228)) and not (inputs(203));
    layer0_outputs(2013) <= not(inputs(28));
    layer0_outputs(2014) <= not(inputs(154));
    layer0_outputs(2015) <= '1';
    layer0_outputs(2016) <= (inputs(100)) or (inputs(21));
    layer0_outputs(2017) <= (inputs(23)) and not (inputs(174));
    layer0_outputs(2018) <= '1';
    layer0_outputs(2019) <= '0';
    layer0_outputs(2020) <= not((inputs(175)) or (inputs(224)));
    layer0_outputs(2021) <= not((inputs(212)) or (inputs(95)));
    layer0_outputs(2022) <= inputs(182);
    layer0_outputs(2023) <= '1';
    layer0_outputs(2024) <= (inputs(156)) and (inputs(48));
    layer0_outputs(2025) <= '0';
    layer0_outputs(2026) <= not((inputs(225)) or (inputs(227)));
    layer0_outputs(2027) <= '1';
    layer0_outputs(2028) <= not(inputs(80));
    layer0_outputs(2029) <= (inputs(21)) and (inputs(26));
    layer0_outputs(2030) <= '0';
    layer0_outputs(2031) <= not(inputs(152)) or (inputs(193));
    layer0_outputs(2032) <= '0';
    layer0_outputs(2033) <= (inputs(255)) and not (inputs(209));
    layer0_outputs(2034) <= '0';
    layer0_outputs(2035) <= '1';
    layer0_outputs(2036) <= '1';
    layer0_outputs(2037) <= not(inputs(8)) or (inputs(97));
    layer0_outputs(2038) <= '1';
    layer0_outputs(2039) <= (inputs(89)) or (inputs(241));
    layer0_outputs(2040) <= not(inputs(52));
    layer0_outputs(2041) <= (inputs(69)) and (inputs(240));
    layer0_outputs(2042) <= not(inputs(255));
    layer0_outputs(2043) <= inputs(234);
    layer0_outputs(2044) <= inputs(90);
    layer0_outputs(2045) <= (inputs(81)) and not (inputs(182));
    layer0_outputs(2046) <= not(inputs(213));
    layer0_outputs(2047) <= '0';
    layer0_outputs(2048) <= not(inputs(107)) or (inputs(251));
    layer0_outputs(2049) <= '0';
    layer0_outputs(2050) <= (inputs(21)) or (inputs(142));
    layer0_outputs(2051) <= (inputs(148)) and not (inputs(150));
    layer0_outputs(2052) <= not((inputs(79)) and (inputs(4)));
    layer0_outputs(2053) <= '1';
    layer0_outputs(2054) <= (inputs(78)) or (inputs(114));
    layer0_outputs(2055) <= not((inputs(43)) and (inputs(13)));
    layer0_outputs(2056) <= not(inputs(0));
    layer0_outputs(2057) <= inputs(34);
    layer0_outputs(2058) <= '1';
    layer0_outputs(2059) <= '0';
    layer0_outputs(2060) <= inputs(78);
    layer0_outputs(2061) <= not(inputs(59)) or (inputs(73));
    layer0_outputs(2062) <= not(inputs(65));
    layer0_outputs(2063) <= (inputs(47)) or (inputs(44));
    layer0_outputs(2064) <= '0';
    layer0_outputs(2065) <= (inputs(98)) or (inputs(131));
    layer0_outputs(2066) <= '1';
    layer0_outputs(2067) <= not(inputs(183));
    layer0_outputs(2068) <= not(inputs(231)) or (inputs(240));
    layer0_outputs(2069) <= '1';
    layer0_outputs(2070) <= '0';
    layer0_outputs(2071) <= inputs(146);
    layer0_outputs(2072) <= '0';
    layer0_outputs(2073) <= (inputs(20)) and not (inputs(97));
    layer0_outputs(2074) <= not((inputs(250)) or (inputs(132)));
    layer0_outputs(2075) <= inputs(82);
    layer0_outputs(2076) <= not(inputs(3));
    layer0_outputs(2077) <= inputs(88);
    layer0_outputs(2078) <= not(inputs(9)) or (inputs(31));
    layer0_outputs(2079) <= not(inputs(126)) or (inputs(165));
    layer0_outputs(2080) <= (inputs(58)) and (inputs(26));
    layer0_outputs(2081) <= (inputs(3)) and not (inputs(244));
    layer0_outputs(2082) <= '0';
    layer0_outputs(2083) <= inputs(35);
    layer0_outputs(2084) <= inputs(158);
    layer0_outputs(2085) <= '0';
    layer0_outputs(2086) <= not((inputs(43)) and (inputs(93)));
    layer0_outputs(2087) <= not((inputs(112)) or (inputs(116)));
    layer0_outputs(2088) <= (inputs(149)) and not (inputs(56));
    layer0_outputs(2089) <= '0';
    layer0_outputs(2090) <= (inputs(31)) and (inputs(248));
    layer0_outputs(2091) <= '1';
    layer0_outputs(2092) <= '0';
    layer0_outputs(2093) <= not(inputs(121)) or (inputs(9));
    layer0_outputs(2094) <= inputs(230);
    layer0_outputs(2095) <= not(inputs(102));
    layer0_outputs(2096) <= (inputs(121)) or (inputs(31));
    layer0_outputs(2097) <= (inputs(95)) and (inputs(250));
    layer0_outputs(2098) <= '1';
    layer0_outputs(2099) <= not((inputs(88)) and (inputs(121)));
    layer0_outputs(2100) <= '0';
    layer0_outputs(2101) <= (inputs(148)) and not (inputs(245));
    layer0_outputs(2102) <= '0';
    layer0_outputs(2103) <= not(inputs(244)) or (inputs(163));
    layer0_outputs(2104) <= (inputs(5)) or (inputs(189));
    layer0_outputs(2105) <= not(inputs(62)) or (inputs(18));
    layer0_outputs(2106) <= not(inputs(20));
    layer0_outputs(2107) <= inputs(157);
    layer0_outputs(2108) <= (inputs(176)) and (inputs(2));
    layer0_outputs(2109) <= (inputs(19)) and not (inputs(213));
    layer0_outputs(2110) <= inputs(174);
    layer0_outputs(2111) <= not(inputs(90)) or (inputs(223));
    layer0_outputs(2112) <= not(inputs(41));
    layer0_outputs(2113) <= (inputs(59)) or (inputs(4));
    layer0_outputs(2114) <= inputs(66);
    layer0_outputs(2115) <= not(inputs(175)) or (inputs(115));
    layer0_outputs(2116) <= (inputs(26)) xor (inputs(72));
    layer0_outputs(2117) <= (inputs(130)) and not (inputs(122));
    layer0_outputs(2118) <= (inputs(78)) or (inputs(111));
    layer0_outputs(2119) <= inputs(184);
    layer0_outputs(2120) <= not((inputs(212)) or (inputs(177)));
    layer0_outputs(2121) <= (inputs(127)) and not (inputs(13));
    layer0_outputs(2122) <= inputs(21);
    layer0_outputs(2123) <= '0';
    layer0_outputs(2124) <= (inputs(38)) and (inputs(241));
    layer0_outputs(2125) <= inputs(45);
    layer0_outputs(2126) <= not(inputs(89));
    layer0_outputs(2127) <= '1';
    layer0_outputs(2128) <= not(inputs(226));
    layer0_outputs(2129) <= not((inputs(100)) or (inputs(120)));
    layer0_outputs(2130) <= '1';
    layer0_outputs(2131) <= '0';
    layer0_outputs(2132) <= not(inputs(195));
    layer0_outputs(2133) <= inputs(122);
    layer0_outputs(2134) <= (inputs(22)) and not (inputs(136));
    layer0_outputs(2135) <= not(inputs(128));
    layer0_outputs(2136) <= not(inputs(22));
    layer0_outputs(2137) <= not((inputs(136)) or (inputs(138)));
    layer0_outputs(2138) <= not(inputs(87));
    layer0_outputs(2139) <= not((inputs(33)) and (inputs(110)));
    layer0_outputs(2140) <= (inputs(71)) and not (inputs(222));
    layer0_outputs(2141) <= (inputs(255)) xor (inputs(36));
    layer0_outputs(2142) <= (inputs(167)) and (inputs(245));
    layer0_outputs(2143) <= inputs(111);
    layer0_outputs(2144) <= (inputs(203)) and not (inputs(137));
    layer0_outputs(2145) <= (inputs(235)) and not (inputs(209));
    layer0_outputs(2146) <= not(inputs(228));
    layer0_outputs(2147) <= not(inputs(196));
    layer0_outputs(2148) <= '0';
    layer0_outputs(2149) <= (inputs(106)) and not (inputs(165));
    layer0_outputs(2150) <= '0';
    layer0_outputs(2151) <= (inputs(180)) and not (inputs(90));
    layer0_outputs(2152) <= inputs(233);
    layer0_outputs(2153) <= not((inputs(86)) xor (inputs(144)));
    layer0_outputs(2154) <= not(inputs(62));
    layer0_outputs(2155) <= '1';
    layer0_outputs(2156) <= '1';
    layer0_outputs(2157) <= (inputs(41)) or (inputs(2));
    layer0_outputs(2158) <= (inputs(35)) and not (inputs(46));
    layer0_outputs(2159) <= (inputs(27)) and not (inputs(243));
    layer0_outputs(2160) <= '1';
    layer0_outputs(2161) <= '1';
    layer0_outputs(2162) <= not(inputs(180));
    layer0_outputs(2163) <= '1';
    layer0_outputs(2164) <= (inputs(26)) and (inputs(205));
    layer0_outputs(2165) <= not(inputs(18));
    layer0_outputs(2166) <= not((inputs(118)) or (inputs(224)));
    layer0_outputs(2167) <= '1';
    layer0_outputs(2168) <= inputs(247);
    layer0_outputs(2169) <= inputs(133);
    layer0_outputs(2170) <= not(inputs(140)) or (inputs(36));
    layer0_outputs(2171) <= '1';
    layer0_outputs(2172) <= (inputs(245)) and (inputs(226));
    layer0_outputs(2173) <= not(inputs(75)) or (inputs(47));
    layer0_outputs(2174) <= (inputs(18)) or (inputs(208));
    layer0_outputs(2175) <= inputs(128);
    layer0_outputs(2176) <= '0';
    layer0_outputs(2177) <= inputs(160);
    layer0_outputs(2178) <= (inputs(136)) and not (inputs(249));
    layer0_outputs(2179) <= '0';
    layer0_outputs(2180) <= '0';
    layer0_outputs(2181) <= (inputs(30)) and not (inputs(217));
    layer0_outputs(2182) <= '1';
    layer0_outputs(2183) <= (inputs(45)) and not (inputs(105));
    layer0_outputs(2184) <= '1';
    layer0_outputs(2185) <= (inputs(51)) xor (inputs(207));
    layer0_outputs(2186) <= not(inputs(188));
    layer0_outputs(2187) <= '1';
    layer0_outputs(2188) <= '0';
    layer0_outputs(2189) <= '1';
    layer0_outputs(2190) <= not(inputs(255));
    layer0_outputs(2191) <= inputs(153);
    layer0_outputs(2192) <= inputs(163);
    layer0_outputs(2193) <= not(inputs(225));
    layer0_outputs(2194) <= '1';
    layer0_outputs(2195) <= '1';
    layer0_outputs(2196) <= '0';
    layer0_outputs(2197) <= '0';
    layer0_outputs(2198) <= not(inputs(146));
    layer0_outputs(2199) <= '1';
    layer0_outputs(2200) <= not(inputs(187)) or (inputs(147));
    layer0_outputs(2201) <= '1';
    layer0_outputs(2202) <= not(inputs(96));
    layer0_outputs(2203) <= (inputs(206)) and (inputs(176));
    layer0_outputs(2204) <= '0';
    layer0_outputs(2205) <= inputs(15);
    layer0_outputs(2206) <= '1';
    layer0_outputs(2207) <= not(inputs(233)) or (inputs(88));
    layer0_outputs(2208) <= inputs(157);
    layer0_outputs(2209) <= (inputs(42)) and (inputs(160));
    layer0_outputs(2210) <= not(inputs(2)) or (inputs(62));
    layer0_outputs(2211) <= (inputs(58)) or (inputs(219));
    layer0_outputs(2212) <= inputs(145);
    layer0_outputs(2213) <= (inputs(199)) and (inputs(169));
    layer0_outputs(2214) <= not((inputs(114)) and (inputs(6)));
    layer0_outputs(2215) <= '0';
    layer0_outputs(2216) <= inputs(35);
    layer0_outputs(2217) <= '1';
    layer0_outputs(2218) <= not(inputs(166));
    layer0_outputs(2219) <= not(inputs(141));
    layer0_outputs(2220) <= (inputs(130)) and not (inputs(227));
    layer0_outputs(2221) <= not(inputs(104)) or (inputs(81));
    layer0_outputs(2222) <= not((inputs(56)) and (inputs(171)));
    layer0_outputs(2223) <= not(inputs(153));
    layer0_outputs(2224) <= not((inputs(223)) and (inputs(246)));
    layer0_outputs(2225) <= '1';
    layer0_outputs(2226) <= not(inputs(73));
    layer0_outputs(2227) <= '1';
    layer0_outputs(2228) <= (inputs(69)) and not (inputs(206));
    layer0_outputs(2229) <= '0';
    layer0_outputs(2230) <= not((inputs(227)) or (inputs(239)));
    layer0_outputs(2231) <= not((inputs(87)) or (inputs(136)));
    layer0_outputs(2232) <= '1';
    layer0_outputs(2233) <= not((inputs(152)) or (inputs(168)));
    layer0_outputs(2234) <= inputs(195);
    layer0_outputs(2235) <= '1';
    layer0_outputs(2236) <= '1';
    layer0_outputs(2237) <= (inputs(64)) or (inputs(97));
    layer0_outputs(2238) <= '0';
    layer0_outputs(2239) <= '1';
    layer0_outputs(2240) <= '0';
    layer0_outputs(2241) <= (inputs(246)) xor (inputs(199));
    layer0_outputs(2242) <= not(inputs(187)) or (inputs(68));
    layer0_outputs(2243) <= inputs(152);
    layer0_outputs(2244) <= not(inputs(79));
    layer0_outputs(2245) <= not(inputs(116));
    layer0_outputs(2246) <= not(inputs(76));
    layer0_outputs(2247) <= '1';
    layer0_outputs(2248) <= '1';
    layer0_outputs(2249) <= '0';
    layer0_outputs(2250) <= inputs(11);
    layer0_outputs(2251) <= (inputs(142)) and not (inputs(166));
    layer0_outputs(2252) <= not((inputs(206)) and (inputs(226)));
    layer0_outputs(2253) <= (inputs(136)) and not (inputs(34));
    layer0_outputs(2254) <= inputs(72);
    layer0_outputs(2255) <= '0';
    layer0_outputs(2256) <= (inputs(218)) or (inputs(219));
    layer0_outputs(2257) <= (inputs(169)) and (inputs(28));
    layer0_outputs(2258) <= (inputs(9)) and not (inputs(161));
    layer0_outputs(2259) <= not(inputs(6));
    layer0_outputs(2260) <= not((inputs(120)) and (inputs(17)));
    layer0_outputs(2261) <= not(inputs(209));
    layer0_outputs(2262) <= not(inputs(53)) or (inputs(38));
    layer0_outputs(2263) <= '0';
    layer0_outputs(2264) <= '1';
    layer0_outputs(2265) <= not(inputs(179));
    layer0_outputs(2266) <= not(inputs(179));
    layer0_outputs(2267) <= inputs(154);
    layer0_outputs(2268) <= not(inputs(235));
    layer0_outputs(2269) <= not(inputs(59)) or (inputs(105));
    layer0_outputs(2270) <= not((inputs(189)) and (inputs(130)));
    layer0_outputs(2271) <= inputs(0);
    layer0_outputs(2272) <= inputs(85);
    layer0_outputs(2273) <= (inputs(26)) and not (inputs(14));
    layer0_outputs(2274) <= not((inputs(127)) or (inputs(144)));
    layer0_outputs(2275) <= not(inputs(226));
    layer0_outputs(2276) <= not(inputs(1));
    layer0_outputs(2277) <= not(inputs(8)) or (inputs(229));
    layer0_outputs(2278) <= '1';
    layer0_outputs(2279) <= '1';
    layer0_outputs(2280) <= '1';
    layer0_outputs(2281) <= not(inputs(187));
    layer0_outputs(2282) <= (inputs(206)) xor (inputs(61));
    layer0_outputs(2283) <= '0';
    layer0_outputs(2284) <= not(inputs(161));
    layer0_outputs(2285) <= not(inputs(83)) or (inputs(190));
    layer0_outputs(2286) <= '0';
    layer0_outputs(2287) <= not(inputs(207)) or (inputs(66));
    layer0_outputs(2288) <= '1';
    layer0_outputs(2289) <= not(inputs(157)) or (inputs(149));
    layer0_outputs(2290) <= (inputs(160)) or (inputs(177));
    layer0_outputs(2291) <= not((inputs(149)) and (inputs(9)));
    layer0_outputs(2292) <= (inputs(26)) and not (inputs(203));
    layer0_outputs(2293) <= '1';
    layer0_outputs(2294) <= not((inputs(170)) or (inputs(253)));
    layer0_outputs(2295) <= (inputs(186)) xor (inputs(120));
    layer0_outputs(2296) <= (inputs(168)) xor (inputs(182));
    layer0_outputs(2297) <= '0';
    layer0_outputs(2298) <= '1';
    layer0_outputs(2299) <= '1';
    layer0_outputs(2300) <= (inputs(208)) and not (inputs(215));
    layer0_outputs(2301) <= not(inputs(98));
    layer0_outputs(2302) <= '0';
    layer0_outputs(2303) <= inputs(93);
    layer0_outputs(2304) <= not(inputs(47)) or (inputs(242));
    layer0_outputs(2305) <= not((inputs(165)) or (inputs(48)));
    layer0_outputs(2306) <= not(inputs(141)) or (inputs(167));
    layer0_outputs(2307) <= '0';
    layer0_outputs(2308) <= '0';
    layer0_outputs(2309) <= '0';
    layer0_outputs(2310) <= '0';
    layer0_outputs(2311) <= not((inputs(91)) and (inputs(127)));
    layer0_outputs(2312) <= inputs(54);
    layer0_outputs(2313) <= '0';
    layer0_outputs(2314) <= not(inputs(233)) or (inputs(233));
    layer0_outputs(2315) <= '1';
    layer0_outputs(2316) <= (inputs(247)) or (inputs(112));
    layer0_outputs(2317) <= (inputs(38)) and not (inputs(85));
    layer0_outputs(2318) <= not((inputs(74)) or (inputs(58)));
    layer0_outputs(2319) <= '1';
    layer0_outputs(2320) <= (inputs(157)) or (inputs(25));
    layer0_outputs(2321) <= inputs(54);
    layer0_outputs(2322) <= not((inputs(80)) and (inputs(251)));
    layer0_outputs(2323) <= inputs(205);
    layer0_outputs(2324) <= not(inputs(29));
    layer0_outputs(2325) <= not((inputs(191)) xor (inputs(132)));
    layer0_outputs(2326) <= (inputs(64)) and (inputs(94));
    layer0_outputs(2327) <= not(inputs(207)) or (inputs(181));
    layer0_outputs(2328) <= '1';
    layer0_outputs(2329) <= (inputs(29)) and (inputs(251));
    layer0_outputs(2330) <= not(inputs(109)) or (inputs(147));
    layer0_outputs(2331) <= inputs(38);
    layer0_outputs(2332) <= '1';
    layer0_outputs(2333) <= not(inputs(170)) or (inputs(215));
    layer0_outputs(2334) <= not((inputs(110)) xor (inputs(174)));
    layer0_outputs(2335) <= not(inputs(29)) or (inputs(85));
    layer0_outputs(2336) <= not(inputs(103));
    layer0_outputs(2337) <= '1';
    layer0_outputs(2338) <= not(inputs(35));
    layer0_outputs(2339) <= '0';
    layer0_outputs(2340) <= not(inputs(77));
    layer0_outputs(2341) <= not(inputs(178));
    layer0_outputs(2342) <= '1';
    layer0_outputs(2343) <= inputs(118);
    layer0_outputs(2344) <= (inputs(172)) or (inputs(157));
    layer0_outputs(2345) <= inputs(158);
    layer0_outputs(2346) <= not(inputs(9));
    layer0_outputs(2347) <= inputs(213);
    layer0_outputs(2348) <= '0';
    layer0_outputs(2349) <= not((inputs(4)) or (inputs(229)));
    layer0_outputs(2350) <= not(inputs(68));
    layer0_outputs(2351) <= inputs(134);
    layer0_outputs(2352) <= inputs(215);
    layer0_outputs(2353) <= inputs(121);
    layer0_outputs(2354) <= (inputs(44)) and (inputs(118));
    layer0_outputs(2355) <= not(inputs(107)) or (inputs(213));
    layer0_outputs(2356) <= not(inputs(24));
    layer0_outputs(2357) <= '1';
    layer0_outputs(2358) <= (inputs(245)) and (inputs(246));
    layer0_outputs(2359) <= not((inputs(148)) or (inputs(182)));
    layer0_outputs(2360) <= not(inputs(172));
    layer0_outputs(2361) <= not((inputs(139)) or (inputs(152)));
    layer0_outputs(2362) <= not((inputs(145)) xor (inputs(239)));
    layer0_outputs(2363) <= '1';
    layer0_outputs(2364) <= '0';
    layer0_outputs(2365) <= (inputs(31)) and not (inputs(105));
    layer0_outputs(2366) <= not(inputs(168));
    layer0_outputs(2367) <= inputs(106);
    layer0_outputs(2368) <= (inputs(122)) or (inputs(255));
    layer0_outputs(2369) <= not((inputs(240)) and (inputs(244)));
    layer0_outputs(2370) <= '1';
    layer0_outputs(2371) <= (inputs(193)) and not (inputs(23));
    layer0_outputs(2372) <= not(inputs(198)) or (inputs(94));
    layer0_outputs(2373) <= not(inputs(130)) or (inputs(178));
    layer0_outputs(2374) <= (inputs(109)) xor (inputs(23));
    layer0_outputs(2375) <= inputs(96);
    layer0_outputs(2376) <= (inputs(175)) and (inputs(196));
    layer0_outputs(2377) <= '0';
    layer0_outputs(2378) <= not(inputs(165));
    layer0_outputs(2379) <= '0';
    layer0_outputs(2380) <= not((inputs(74)) and (inputs(190)));
    layer0_outputs(2381) <= (inputs(27)) and not (inputs(244));
    layer0_outputs(2382) <= (inputs(125)) and (inputs(169));
    layer0_outputs(2383) <= not(inputs(163));
    layer0_outputs(2384) <= '0';
    layer0_outputs(2385) <= not(inputs(1)) or (inputs(41));
    layer0_outputs(2386) <= (inputs(27)) and not (inputs(91));
    layer0_outputs(2387) <= not(inputs(144));
    layer0_outputs(2388) <= (inputs(24)) and (inputs(84));
    layer0_outputs(2389) <= (inputs(4)) and not (inputs(133));
    layer0_outputs(2390) <= not(inputs(235));
    layer0_outputs(2391) <= inputs(120);
    layer0_outputs(2392) <= '1';
    layer0_outputs(2393) <= not((inputs(85)) and (inputs(75)));
    layer0_outputs(2394) <= (inputs(70)) or (inputs(147));
    layer0_outputs(2395) <= not((inputs(183)) and (inputs(57)));
    layer0_outputs(2396) <= not((inputs(155)) or (inputs(3)));
    layer0_outputs(2397) <= not(inputs(39)) or (inputs(36));
    layer0_outputs(2398) <= (inputs(140)) and (inputs(16));
    layer0_outputs(2399) <= not(inputs(152));
    layer0_outputs(2400) <= (inputs(223)) and (inputs(65));
    layer0_outputs(2401) <= (inputs(207)) and (inputs(39));
    layer0_outputs(2402) <= '0';
    layer0_outputs(2403) <= not((inputs(96)) xor (inputs(211)));
    layer0_outputs(2404) <= '1';
    layer0_outputs(2405) <= not(inputs(179)) or (inputs(49));
    layer0_outputs(2406) <= '0';
    layer0_outputs(2407) <= not(inputs(96)) or (inputs(136));
    layer0_outputs(2408) <= (inputs(46)) and (inputs(121));
    layer0_outputs(2409) <= '1';
    layer0_outputs(2410) <= not((inputs(86)) or (inputs(108)));
    layer0_outputs(2411) <= not(inputs(172));
    layer0_outputs(2412) <= inputs(179);
    layer0_outputs(2413) <= not(inputs(252)) or (inputs(202));
    layer0_outputs(2414) <= not((inputs(51)) or (inputs(147)));
    layer0_outputs(2415) <= not(inputs(7));
    layer0_outputs(2416) <= not(inputs(160));
    layer0_outputs(2417) <= '1';
    layer0_outputs(2418) <= not((inputs(45)) and (inputs(143)));
    layer0_outputs(2419) <= not(inputs(145));
    layer0_outputs(2420) <= (inputs(247)) and (inputs(113));
    layer0_outputs(2421) <= inputs(103);
    layer0_outputs(2422) <= '1';
    layer0_outputs(2423) <= (inputs(196)) and not (inputs(115));
    layer0_outputs(2424) <= '1';
    layer0_outputs(2425) <= '1';
    layer0_outputs(2426) <= not(inputs(128));
    layer0_outputs(2427) <= not((inputs(59)) or (inputs(43)));
    layer0_outputs(2428) <= '0';
    layer0_outputs(2429) <= inputs(108);
    layer0_outputs(2430) <= not(inputs(141)) or (inputs(254));
    layer0_outputs(2431) <= (inputs(184)) and (inputs(196));
    layer0_outputs(2432) <= inputs(114);
    layer0_outputs(2433) <= inputs(8);
    layer0_outputs(2434) <= '1';
    layer0_outputs(2435) <= (inputs(0)) and not (inputs(194));
    layer0_outputs(2436) <= '1';
    layer0_outputs(2437) <= '0';
    layer0_outputs(2438) <= not(inputs(4)) or (inputs(215));
    layer0_outputs(2439) <= '0';
    layer0_outputs(2440) <= not(inputs(82)) or (inputs(181));
    layer0_outputs(2441) <= inputs(144);
    layer0_outputs(2442) <= not((inputs(45)) and (inputs(95)));
    layer0_outputs(2443) <= not(inputs(3)) or (inputs(226));
    layer0_outputs(2444) <= not((inputs(203)) or (inputs(26)));
    layer0_outputs(2445) <= not(inputs(189));
    layer0_outputs(2446) <= not(inputs(161));
    layer0_outputs(2447) <= (inputs(179)) or (inputs(254));
    layer0_outputs(2448) <= inputs(29);
    layer0_outputs(2449) <= not(inputs(209)) or (inputs(155));
    layer0_outputs(2450) <= not((inputs(181)) and (inputs(202)));
    layer0_outputs(2451) <= '0';
    layer0_outputs(2452) <= '0';
    layer0_outputs(2453) <= inputs(196);
    layer0_outputs(2454) <= not(inputs(90)) or (inputs(37));
    layer0_outputs(2455) <= not((inputs(29)) or (inputs(224)));
    layer0_outputs(2456) <= not(inputs(41));
    layer0_outputs(2457) <= '1';
    layer0_outputs(2458) <= not(inputs(75)) or (inputs(191));
    layer0_outputs(2459) <= not((inputs(245)) xor (inputs(133)));
    layer0_outputs(2460) <= not(inputs(157));
    layer0_outputs(2461) <= '1';
    layer0_outputs(2462) <= '1';
    layer0_outputs(2463) <= not(inputs(163));
    layer0_outputs(2464) <= '0';
    layer0_outputs(2465) <= '0';
    layer0_outputs(2466) <= (inputs(41)) or (inputs(80));
    layer0_outputs(2467) <= '0';
    layer0_outputs(2468) <= not(inputs(165));
    layer0_outputs(2469) <= (inputs(168)) and not (inputs(69));
    layer0_outputs(2470) <= not(inputs(200));
    layer0_outputs(2471) <= (inputs(243)) or (inputs(30));
    layer0_outputs(2472) <= inputs(4);
    layer0_outputs(2473) <= inputs(183);
    layer0_outputs(2474) <= '0';
    layer0_outputs(2475) <= (inputs(225)) and not (inputs(69));
    layer0_outputs(2476) <= '0';
    layer0_outputs(2477) <= '1';
    layer0_outputs(2478) <= (inputs(2)) and (inputs(233));
    layer0_outputs(2479) <= '0';
    layer0_outputs(2480) <= not(inputs(80));
    layer0_outputs(2481) <= '1';
    layer0_outputs(2482) <= not(inputs(52)) or (inputs(3));
    layer0_outputs(2483) <= not(inputs(167));
    layer0_outputs(2484) <= '1';
    layer0_outputs(2485) <= (inputs(19)) and not (inputs(109));
    layer0_outputs(2486) <= (inputs(129)) or (inputs(195));
    layer0_outputs(2487) <= not(inputs(225));
    layer0_outputs(2488) <= inputs(44);
    layer0_outputs(2489) <= not(inputs(171)) or (inputs(26));
    layer0_outputs(2490) <= inputs(155);
    layer0_outputs(2491) <= not(inputs(253));
    layer0_outputs(2492) <= (inputs(189)) and not (inputs(204));
    layer0_outputs(2493) <= inputs(78);
    layer0_outputs(2494) <= '0';
    layer0_outputs(2495) <= (inputs(191)) or (inputs(25));
    layer0_outputs(2496) <= not((inputs(90)) and (inputs(117)));
    layer0_outputs(2497) <= not((inputs(138)) or (inputs(113)));
    layer0_outputs(2498) <= (inputs(48)) and (inputs(54));
    layer0_outputs(2499) <= inputs(39);
    layer0_outputs(2500) <= '0';
    layer0_outputs(2501) <= (inputs(70)) and not (inputs(132));
    layer0_outputs(2502) <= (inputs(53)) or (inputs(131));
    layer0_outputs(2503) <= not((inputs(27)) or (inputs(88)));
    layer0_outputs(2504) <= not(inputs(181)) or (inputs(166));
    layer0_outputs(2505) <= not((inputs(207)) xor (inputs(149)));
    layer0_outputs(2506) <= not((inputs(250)) and (inputs(32)));
    layer0_outputs(2507) <= inputs(17);
    layer0_outputs(2508) <= '1';
    layer0_outputs(2509) <= (inputs(250)) and not (inputs(200));
    layer0_outputs(2510) <= not((inputs(255)) xor (inputs(88)));
    layer0_outputs(2511) <= '0';
    layer0_outputs(2512) <= not((inputs(29)) or (inputs(103)));
    layer0_outputs(2513) <= inputs(97);
    layer0_outputs(2514) <= '1';
    layer0_outputs(2515) <= (inputs(228)) and not (inputs(103));
    layer0_outputs(2516) <= (inputs(7)) or (inputs(68));
    layer0_outputs(2517) <= '0';
    layer0_outputs(2518) <= not(inputs(99));
    layer0_outputs(2519) <= inputs(82);
    layer0_outputs(2520) <= '0';
    layer0_outputs(2521) <= inputs(66);
    layer0_outputs(2522) <= not(inputs(186)) or (inputs(71));
    layer0_outputs(2523) <= not(inputs(252));
    layer0_outputs(2524) <= not((inputs(61)) and (inputs(53)));
    layer0_outputs(2525) <= (inputs(144)) and not (inputs(13));
    layer0_outputs(2526) <= inputs(148);
    layer0_outputs(2527) <= not((inputs(143)) and (inputs(241)));
    layer0_outputs(2528) <= '0';
    layer0_outputs(2529) <= not((inputs(115)) or (inputs(238)));
    layer0_outputs(2530) <= not(inputs(243)) or (inputs(180));
    layer0_outputs(2531) <= inputs(17);
    layer0_outputs(2532) <= '1';
    layer0_outputs(2533) <= '0';
    layer0_outputs(2534) <= (inputs(218)) and (inputs(124));
    layer0_outputs(2535) <= '0';
    layer0_outputs(2536) <= '1';
    layer0_outputs(2537) <= (inputs(89)) or (inputs(245));
    layer0_outputs(2538) <= inputs(76);
    layer0_outputs(2539) <= not(inputs(69)) or (inputs(225));
    layer0_outputs(2540) <= (inputs(187)) or (inputs(207));
    layer0_outputs(2541) <= inputs(211);
    layer0_outputs(2542) <= not((inputs(102)) and (inputs(55)));
    layer0_outputs(2543) <= '0';
    layer0_outputs(2544) <= not(inputs(104)) or (inputs(28));
    layer0_outputs(2545) <= '0';
    layer0_outputs(2546) <= not(inputs(93));
    layer0_outputs(2547) <= inputs(148);
    layer0_outputs(2548) <= not(inputs(246));
    layer0_outputs(2549) <= not((inputs(52)) or (inputs(128)));
    layer0_outputs(2550) <= '0';
    layer0_outputs(2551) <= inputs(233);
    layer0_outputs(2552) <= inputs(199);
    layer0_outputs(2553) <= '0';
    layer0_outputs(2554) <= inputs(49);
    layer0_outputs(2555) <= '1';
    layer0_outputs(2556) <= not((inputs(120)) and (inputs(5)));
    layer0_outputs(2557) <= inputs(70);
    layer0_outputs(2558) <= not(inputs(205));
    layer0_outputs(2559) <= not(inputs(97)) or (inputs(16));
    layer0_outputs(2560) <= (inputs(21)) and not (inputs(154));
    layer0_outputs(2561) <= not((inputs(96)) or (inputs(160)));
    layer0_outputs(2562) <= (inputs(192)) or (inputs(193));
    layer0_outputs(2563) <= not(inputs(178)) or (inputs(70));
    layer0_outputs(2564) <= '1';
    layer0_outputs(2565) <= '0';
    layer0_outputs(2566) <= not(inputs(96));
    layer0_outputs(2567) <= (inputs(109)) and not (inputs(251));
    layer0_outputs(2568) <= not(inputs(64));
    layer0_outputs(2569) <= not(inputs(255));
    layer0_outputs(2570) <= not(inputs(234)) or (inputs(12));
    layer0_outputs(2571) <= inputs(105);
    layer0_outputs(2572) <= inputs(168);
    layer0_outputs(2573) <= not((inputs(237)) or (inputs(196)));
    layer0_outputs(2574) <= not(inputs(145)) or (inputs(79));
    layer0_outputs(2575) <= '0';
    layer0_outputs(2576) <= '1';
    layer0_outputs(2577) <= (inputs(178)) or (inputs(176));
    layer0_outputs(2578) <= inputs(17);
    layer0_outputs(2579) <= '0';
    layer0_outputs(2580) <= '1';
    layer0_outputs(2581) <= not(inputs(193)) or (inputs(228));
    layer0_outputs(2582) <= (inputs(113)) and (inputs(30));
    layer0_outputs(2583) <= (inputs(224)) and not (inputs(123));
    layer0_outputs(2584) <= (inputs(228)) or (inputs(112));
    layer0_outputs(2585) <= not(inputs(236)) or (inputs(32));
    layer0_outputs(2586) <= not(inputs(240));
    layer0_outputs(2587) <= (inputs(12)) and not (inputs(132));
    layer0_outputs(2588) <= (inputs(193)) xor (inputs(215));
    layer0_outputs(2589) <= '0';
    layer0_outputs(2590) <= not(inputs(38));
    layer0_outputs(2591) <= (inputs(66)) and not (inputs(176));
    layer0_outputs(2592) <= (inputs(206)) or (inputs(222));
    layer0_outputs(2593) <= '1';
    layer0_outputs(2594) <= not((inputs(27)) or (inputs(7)));
    layer0_outputs(2595) <= inputs(106);
    layer0_outputs(2596) <= (inputs(79)) and not (inputs(122));
    layer0_outputs(2597) <= not((inputs(226)) and (inputs(143)));
    layer0_outputs(2598) <= (inputs(93)) and not (inputs(35));
    layer0_outputs(2599) <= (inputs(19)) or (inputs(119));
    layer0_outputs(2600) <= inputs(33);
    layer0_outputs(2601) <= not(inputs(214));
    layer0_outputs(2602) <= not(inputs(48)) or (inputs(16));
    layer0_outputs(2603) <= not((inputs(237)) or (inputs(122)));
    layer0_outputs(2604) <= not((inputs(134)) and (inputs(142)));
    layer0_outputs(2605) <= inputs(142);
    layer0_outputs(2606) <= '0';
    layer0_outputs(2607) <= not(inputs(130));
    layer0_outputs(2608) <= inputs(143);
    layer0_outputs(2609) <= inputs(206);
    layer0_outputs(2610) <= inputs(168);
    layer0_outputs(2611) <= not((inputs(124)) xor (inputs(155)));
    layer0_outputs(2612) <= not((inputs(218)) and (inputs(68)));
    layer0_outputs(2613) <= '0';
    layer0_outputs(2614) <= (inputs(156)) and (inputs(133));
    layer0_outputs(2615) <= (inputs(159)) or (inputs(78));
    layer0_outputs(2616) <= (inputs(230)) and not (inputs(230));
    layer0_outputs(2617) <= (inputs(206)) xor (inputs(48));
    layer0_outputs(2618) <= not(inputs(57));
    layer0_outputs(2619) <= inputs(118);
    layer0_outputs(2620) <= not(inputs(164));
    layer0_outputs(2621) <= not(inputs(99)) or (inputs(233));
    layer0_outputs(2622) <= not(inputs(210)) or (inputs(123));
    layer0_outputs(2623) <= (inputs(30)) xor (inputs(79));
    layer0_outputs(2624) <= (inputs(65)) and not (inputs(55));
    layer0_outputs(2625) <= not((inputs(113)) and (inputs(97)));
    layer0_outputs(2626) <= not(inputs(112));
    layer0_outputs(2627) <= '0';
    layer0_outputs(2628) <= not(inputs(79));
    layer0_outputs(2629) <= (inputs(56)) and not (inputs(56));
    layer0_outputs(2630) <= not(inputs(201)) or (inputs(208));
    layer0_outputs(2631) <= not((inputs(34)) or (inputs(61)));
    layer0_outputs(2632) <= not(inputs(64)) or (inputs(112));
    layer0_outputs(2633) <= (inputs(247)) or (inputs(72));
    layer0_outputs(2634) <= not((inputs(72)) xor (inputs(72)));
    layer0_outputs(2635) <= (inputs(9)) and not (inputs(91));
    layer0_outputs(2636) <= not(inputs(105));
    layer0_outputs(2637) <= not((inputs(95)) and (inputs(159)));
    layer0_outputs(2638) <= not((inputs(173)) or (inputs(181)));
    layer0_outputs(2639) <= (inputs(51)) xor (inputs(252));
    layer0_outputs(2640) <= '0';
    layer0_outputs(2641) <= '1';
    layer0_outputs(2642) <= (inputs(63)) and not (inputs(163));
    layer0_outputs(2643) <= '0';
    layer0_outputs(2644) <= '1';
    layer0_outputs(2645) <= not(inputs(30));
    layer0_outputs(2646) <= inputs(247);
    layer0_outputs(2647) <= not(inputs(108));
    layer0_outputs(2648) <= not(inputs(181));
    layer0_outputs(2649) <= inputs(34);
    layer0_outputs(2650) <= (inputs(114)) or (inputs(131));
    layer0_outputs(2651) <= not(inputs(82));
    layer0_outputs(2652) <= not(inputs(70));
    layer0_outputs(2653) <= not(inputs(103)) or (inputs(227));
    layer0_outputs(2654) <= not(inputs(92));
    layer0_outputs(2655) <= '0';
    layer0_outputs(2656) <= '0';
    layer0_outputs(2657) <= not(inputs(91)) or (inputs(128));
    layer0_outputs(2658) <= (inputs(47)) and (inputs(121));
    layer0_outputs(2659) <= inputs(85);
    layer0_outputs(2660) <= not((inputs(37)) and (inputs(73)));
    layer0_outputs(2661) <= (inputs(31)) and (inputs(0));
    layer0_outputs(2662) <= (inputs(200)) xor (inputs(66));
    layer0_outputs(2663) <= not(inputs(64));
    layer0_outputs(2664) <= '0';
    layer0_outputs(2665) <= not((inputs(5)) or (inputs(24)));
    layer0_outputs(2666) <= inputs(23);
    layer0_outputs(2667) <= '1';
    layer0_outputs(2668) <= (inputs(159)) or (inputs(43));
    layer0_outputs(2669) <= not(inputs(192));
    layer0_outputs(2670) <= '0';
    layer0_outputs(2671) <= (inputs(67)) and not (inputs(131));
    layer0_outputs(2672) <= '1';
    layer0_outputs(2673) <= not(inputs(60));
    layer0_outputs(2674) <= not(inputs(55));
    layer0_outputs(2675) <= (inputs(240)) and (inputs(207));
    layer0_outputs(2676) <= not(inputs(203));
    layer0_outputs(2677) <= '0';
    layer0_outputs(2678) <= not(inputs(145));
    layer0_outputs(2679) <= not(inputs(206)) or (inputs(80));
    layer0_outputs(2680) <= not((inputs(159)) or (inputs(111)));
    layer0_outputs(2681) <= inputs(201);
    layer0_outputs(2682) <= (inputs(176)) and (inputs(161));
    layer0_outputs(2683) <= inputs(50);
    layer0_outputs(2684) <= (inputs(83)) and not (inputs(220));
    layer0_outputs(2685) <= '1';
    layer0_outputs(2686) <= not(inputs(53));
    layer0_outputs(2687) <= (inputs(124)) xor (inputs(170));
    layer0_outputs(2688) <= (inputs(143)) and not (inputs(118));
    layer0_outputs(2689) <= '0';
    layer0_outputs(2690) <= '1';
    layer0_outputs(2691) <= (inputs(43)) and not (inputs(29));
    layer0_outputs(2692) <= '0';
    layer0_outputs(2693) <= '0';
    layer0_outputs(2694) <= not(inputs(218));
    layer0_outputs(2695) <= (inputs(108)) or (inputs(188));
    layer0_outputs(2696) <= not(inputs(179)) or (inputs(137));
    layer0_outputs(2697) <= (inputs(239)) and not (inputs(236));
    layer0_outputs(2698) <= (inputs(40)) and not (inputs(240));
    layer0_outputs(2699) <= '0';
    layer0_outputs(2700) <= (inputs(173)) and not (inputs(232));
    layer0_outputs(2701) <= '0';
    layer0_outputs(2702) <= '0';
    layer0_outputs(2703) <= (inputs(36)) or (inputs(109));
    layer0_outputs(2704) <= inputs(167);
    layer0_outputs(2705) <= not((inputs(47)) and (inputs(94)));
    layer0_outputs(2706) <= '1';
    layer0_outputs(2707) <= (inputs(100)) and not (inputs(99));
    layer0_outputs(2708) <= '0';
    layer0_outputs(2709) <= not((inputs(225)) and (inputs(32)));
    layer0_outputs(2710) <= inputs(11);
    layer0_outputs(2711) <= not(inputs(198)) or (inputs(168));
    layer0_outputs(2712) <= '1';
    layer0_outputs(2713) <= inputs(126);
    layer0_outputs(2714) <= (inputs(209)) and not (inputs(98));
    layer0_outputs(2715) <= (inputs(3)) and not (inputs(234));
    layer0_outputs(2716) <= not((inputs(85)) or (inputs(71)));
    layer0_outputs(2717) <= not(inputs(196)) or (inputs(38));
    layer0_outputs(2718) <= inputs(248);
    layer0_outputs(2719) <= (inputs(110)) and not (inputs(76));
    layer0_outputs(2720) <= (inputs(176)) and (inputs(228));
    layer0_outputs(2721) <= (inputs(155)) and (inputs(41));
    layer0_outputs(2722) <= '1';
    layer0_outputs(2723) <= inputs(47);
    layer0_outputs(2724) <= '1';
    layer0_outputs(2725) <= not(inputs(200));
    layer0_outputs(2726) <= not(inputs(236)) or (inputs(105));
    layer0_outputs(2727) <= not(inputs(47));
    layer0_outputs(2728) <= inputs(2);
    layer0_outputs(2729) <= inputs(61);
    layer0_outputs(2730) <= '1';
    layer0_outputs(2731) <= '1';
    layer0_outputs(2732) <= (inputs(243)) and not (inputs(163));
    layer0_outputs(2733) <= (inputs(111)) or (inputs(85));
    layer0_outputs(2734) <= not(inputs(41)) or (inputs(0));
    layer0_outputs(2735) <= not(inputs(171)) or (inputs(250));
    layer0_outputs(2736) <= not(inputs(171));
    layer0_outputs(2737) <= (inputs(65)) and not (inputs(221));
    layer0_outputs(2738) <= (inputs(36)) xor (inputs(88));
    layer0_outputs(2739) <= not(inputs(236)) or (inputs(5));
    layer0_outputs(2740) <= (inputs(238)) and (inputs(143));
    layer0_outputs(2741) <= not(inputs(167)) or (inputs(72));
    layer0_outputs(2742) <= '1';
    layer0_outputs(2743) <= not((inputs(200)) and (inputs(146)));
    layer0_outputs(2744) <= (inputs(220)) and not (inputs(125));
    layer0_outputs(2745) <= '1';
    layer0_outputs(2746) <= not(inputs(197)) or (inputs(43));
    layer0_outputs(2747) <= (inputs(222)) and not (inputs(27));
    layer0_outputs(2748) <= not(inputs(253)) or (inputs(228));
    layer0_outputs(2749) <= inputs(82);
    layer0_outputs(2750) <= (inputs(188)) and (inputs(1));
    layer0_outputs(2751) <= '1';
    layer0_outputs(2752) <= '0';
    layer0_outputs(2753) <= '1';
    layer0_outputs(2754) <= (inputs(123)) and not (inputs(213));
    layer0_outputs(2755) <= not(inputs(69)) or (inputs(211));
    layer0_outputs(2756) <= inputs(48);
    layer0_outputs(2757) <= not(inputs(78)) or (inputs(129));
    layer0_outputs(2758) <= (inputs(239)) and not (inputs(38));
    layer0_outputs(2759) <= not(inputs(253));
    layer0_outputs(2760) <= (inputs(190)) and not (inputs(165));
    layer0_outputs(2761) <= not((inputs(74)) or (inputs(94)));
    layer0_outputs(2762) <= not((inputs(137)) and (inputs(146)));
    layer0_outputs(2763) <= (inputs(239)) or (inputs(252));
    layer0_outputs(2764) <= inputs(10);
    layer0_outputs(2765) <= '0';
    layer0_outputs(2766) <= (inputs(12)) and not (inputs(176));
    layer0_outputs(2767) <= '0';
    layer0_outputs(2768) <= '1';
    layer0_outputs(2769) <= not(inputs(33));
    layer0_outputs(2770) <= inputs(198);
    layer0_outputs(2771) <= not(inputs(247)) or (inputs(105));
    layer0_outputs(2772) <= '1';
    layer0_outputs(2773) <= not(inputs(65)) or (inputs(215));
    layer0_outputs(2774) <= not(inputs(252));
    layer0_outputs(2775) <= inputs(139);
    layer0_outputs(2776) <= '0';
    layer0_outputs(2777) <= not(inputs(238));
    layer0_outputs(2778) <= (inputs(251)) and not (inputs(3));
    layer0_outputs(2779) <= (inputs(172)) and not (inputs(116));
    layer0_outputs(2780) <= not(inputs(233)) or (inputs(164));
    layer0_outputs(2781) <= not((inputs(188)) and (inputs(163)));
    layer0_outputs(2782) <= '1';
    layer0_outputs(2783) <= not(inputs(96));
    layer0_outputs(2784) <= (inputs(248)) and (inputs(17));
    layer0_outputs(2785) <= '0';
    layer0_outputs(2786) <= not(inputs(180)) or (inputs(75));
    layer0_outputs(2787) <= '1';
    layer0_outputs(2788) <= '1';
    layer0_outputs(2789) <= not((inputs(255)) or (inputs(49)));
    layer0_outputs(2790) <= '1';
    layer0_outputs(2791) <= (inputs(23)) xor (inputs(71));
    layer0_outputs(2792) <= '1';
    layer0_outputs(2793) <= (inputs(249)) or (inputs(31));
    layer0_outputs(2794) <= '0';
    layer0_outputs(2795) <= not((inputs(26)) or (inputs(60)));
    layer0_outputs(2796) <= (inputs(207)) and not (inputs(164));
    layer0_outputs(2797) <= '1';
    layer0_outputs(2798) <= '0';
    layer0_outputs(2799) <= not((inputs(80)) xor (inputs(79)));
    layer0_outputs(2800) <= (inputs(42)) and not (inputs(154));
    layer0_outputs(2801) <= not((inputs(25)) or (inputs(35)));
    layer0_outputs(2802) <= not(inputs(133)) or (inputs(96));
    layer0_outputs(2803) <= not(inputs(157)) or (inputs(74));
    layer0_outputs(2804) <= not((inputs(69)) and (inputs(189)));
    layer0_outputs(2805) <= not(inputs(29));
    layer0_outputs(2806) <= (inputs(84)) and (inputs(185));
    layer0_outputs(2807) <= not(inputs(154));
    layer0_outputs(2808) <= not((inputs(125)) or (inputs(219)));
    layer0_outputs(2809) <= (inputs(197)) and not (inputs(63));
    layer0_outputs(2810) <= '0';
    layer0_outputs(2811) <= inputs(232);
    layer0_outputs(2812) <= not((inputs(219)) or (inputs(248)));
    layer0_outputs(2813) <= (inputs(248)) and not (inputs(233));
    layer0_outputs(2814) <= not((inputs(159)) and (inputs(217)));
    layer0_outputs(2815) <= inputs(165);
    layer0_outputs(2816) <= '0';
    layer0_outputs(2817) <= '1';
    layer0_outputs(2818) <= '0';
    layer0_outputs(2819) <= '1';
    layer0_outputs(2820) <= (inputs(50)) and not (inputs(74));
    layer0_outputs(2821) <= (inputs(155)) and not (inputs(86));
    layer0_outputs(2822) <= (inputs(79)) and (inputs(137));
    layer0_outputs(2823) <= (inputs(196)) and not (inputs(227));
    layer0_outputs(2824) <= (inputs(102)) and (inputs(249));
    layer0_outputs(2825) <= '0';
    layer0_outputs(2826) <= '1';
    layer0_outputs(2827) <= not(inputs(233));
    layer0_outputs(2828) <= '0';
    layer0_outputs(2829) <= '1';
    layer0_outputs(2830) <= '1';
    layer0_outputs(2831) <= '0';
    layer0_outputs(2832) <= not(inputs(212));
    layer0_outputs(2833) <= not((inputs(188)) and (inputs(106)));
    layer0_outputs(2834) <= not(inputs(9));
    layer0_outputs(2835) <= not((inputs(135)) or (inputs(88)));
    layer0_outputs(2836) <= (inputs(201)) and not (inputs(248));
    layer0_outputs(2837) <= (inputs(82)) or (inputs(20));
    layer0_outputs(2838) <= (inputs(124)) and (inputs(85));
    layer0_outputs(2839) <= not(inputs(211));
    layer0_outputs(2840) <= not(inputs(67)) or (inputs(147));
    layer0_outputs(2841) <= (inputs(30)) and not (inputs(167));
    layer0_outputs(2842) <= not((inputs(222)) and (inputs(25)));
    layer0_outputs(2843) <= '1';
    layer0_outputs(2844) <= (inputs(193)) and not (inputs(71));
    layer0_outputs(2845) <= inputs(216);
    layer0_outputs(2846) <= not(inputs(4)) or (inputs(219));
    layer0_outputs(2847) <= not((inputs(139)) and (inputs(179)));
    layer0_outputs(2848) <= '0';
    layer0_outputs(2849) <= inputs(167);
    layer0_outputs(2850) <= '1';
    layer0_outputs(2851) <= inputs(243);
    layer0_outputs(2852) <= not(inputs(13));
    layer0_outputs(2853) <= (inputs(214)) and (inputs(166));
    layer0_outputs(2854) <= inputs(198);
    layer0_outputs(2855) <= not((inputs(66)) or (inputs(75)));
    layer0_outputs(2856) <= '0';
    layer0_outputs(2857) <= '0';
    layer0_outputs(2858) <= (inputs(180)) xor (inputs(207));
    layer0_outputs(2859) <= '0';
    layer0_outputs(2860) <= '0';
    layer0_outputs(2861) <= (inputs(85)) and (inputs(212));
    layer0_outputs(2862) <= (inputs(129)) and (inputs(40));
    layer0_outputs(2863) <= (inputs(248)) and (inputs(153));
    layer0_outputs(2864) <= not((inputs(127)) and (inputs(205)));
    layer0_outputs(2865) <= (inputs(56)) and (inputs(187));
    layer0_outputs(2866) <= not(inputs(220)) or (inputs(93));
    layer0_outputs(2867) <= not(inputs(6)) or (inputs(211));
    layer0_outputs(2868) <= (inputs(144)) and (inputs(154));
    layer0_outputs(2869) <= inputs(239);
    layer0_outputs(2870) <= not(inputs(123)) or (inputs(101));
    layer0_outputs(2871) <= '1';
    layer0_outputs(2872) <= '0';
    layer0_outputs(2873) <= '0';
    layer0_outputs(2874) <= not((inputs(237)) or (inputs(239)));
    layer0_outputs(2875) <= not(inputs(61)) or (inputs(27));
    layer0_outputs(2876) <= (inputs(24)) and (inputs(73));
    layer0_outputs(2877) <= not((inputs(104)) and (inputs(62)));
    layer0_outputs(2878) <= not(inputs(160)) or (inputs(111));
    layer0_outputs(2879) <= '0';
    layer0_outputs(2880) <= '0';
    layer0_outputs(2881) <= inputs(237);
    layer0_outputs(2882) <= inputs(130);
    layer0_outputs(2883) <= not((inputs(92)) or (inputs(109)));
    layer0_outputs(2884) <= '1';
    layer0_outputs(2885) <= '1';
    layer0_outputs(2886) <= not(inputs(126));
    layer0_outputs(2887) <= inputs(222);
    layer0_outputs(2888) <= '0';
    layer0_outputs(2889) <= not(inputs(162));
    layer0_outputs(2890) <= '0';
    layer0_outputs(2891) <= '1';
    layer0_outputs(2892) <= (inputs(25)) and not (inputs(40));
    layer0_outputs(2893) <= not(inputs(122));
    layer0_outputs(2894) <= (inputs(161)) and not (inputs(86));
    layer0_outputs(2895) <= not((inputs(237)) or (inputs(150)));
    layer0_outputs(2896) <= '1';
    layer0_outputs(2897) <= (inputs(187)) or (inputs(239));
    layer0_outputs(2898) <= not(inputs(178));
    layer0_outputs(2899) <= not((inputs(51)) and (inputs(46)));
    layer0_outputs(2900) <= not(inputs(242)) or (inputs(135));
    layer0_outputs(2901) <= (inputs(115)) and not (inputs(255));
    layer0_outputs(2902) <= (inputs(213)) and (inputs(232));
    layer0_outputs(2903) <= not(inputs(157));
    layer0_outputs(2904) <= not(inputs(8));
    layer0_outputs(2905) <= '1';
    layer0_outputs(2906) <= '0';
    layer0_outputs(2907) <= (inputs(184)) and not (inputs(145));
    layer0_outputs(2908) <= not(inputs(64));
    layer0_outputs(2909) <= (inputs(140)) and not (inputs(38));
    layer0_outputs(2910) <= '0';
    layer0_outputs(2911) <= (inputs(119)) and (inputs(107));
    layer0_outputs(2912) <= (inputs(190)) and not (inputs(25));
    layer0_outputs(2913) <= (inputs(63)) or (inputs(152));
    layer0_outputs(2914) <= not((inputs(136)) or (inputs(102)));
    layer0_outputs(2915) <= '1';
    layer0_outputs(2916) <= not((inputs(90)) and (inputs(11)));
    layer0_outputs(2917) <= not((inputs(50)) or (inputs(152)));
    layer0_outputs(2918) <= '0';
    layer0_outputs(2919) <= '0';
    layer0_outputs(2920) <= inputs(117);
    layer0_outputs(2921) <= not(inputs(191));
    layer0_outputs(2922) <= inputs(190);
    layer0_outputs(2923) <= not(inputs(63));
    layer0_outputs(2924) <= '1';
    layer0_outputs(2925) <= '0';
    layer0_outputs(2926) <= '1';
    layer0_outputs(2927) <= (inputs(71)) and not (inputs(1));
    layer0_outputs(2928) <= (inputs(190)) and not (inputs(199));
    layer0_outputs(2929) <= (inputs(44)) and not (inputs(243));
    layer0_outputs(2930) <= '0';
    layer0_outputs(2931) <= not(inputs(150));
    layer0_outputs(2932) <= '0';
    layer0_outputs(2933) <= inputs(79);
    layer0_outputs(2934) <= inputs(169);
    layer0_outputs(2935) <= not(inputs(107));
    layer0_outputs(2936) <= '1';
    layer0_outputs(2937) <= not((inputs(18)) or (inputs(222)));
    layer0_outputs(2938) <= not(inputs(24));
    layer0_outputs(2939) <= '1';
    layer0_outputs(2940) <= '1';
    layer0_outputs(2941) <= (inputs(152)) and not (inputs(92));
    layer0_outputs(2942) <= '0';
    layer0_outputs(2943) <= not(inputs(37)) or (inputs(131));
    layer0_outputs(2944) <= (inputs(177)) and (inputs(114));
    layer0_outputs(2945) <= '1';
    layer0_outputs(2946) <= inputs(15);
    layer0_outputs(2947) <= not((inputs(172)) and (inputs(112)));
    layer0_outputs(2948) <= not(inputs(220));
    layer0_outputs(2949) <= '1';
    layer0_outputs(2950) <= inputs(32);
    layer0_outputs(2951) <= (inputs(115)) and (inputs(112));
    layer0_outputs(2952) <= inputs(247);
    layer0_outputs(2953) <= not(inputs(143));
    layer0_outputs(2954) <= inputs(203);
    layer0_outputs(2955) <= (inputs(174)) or (inputs(72));
    layer0_outputs(2956) <= '1';
    layer0_outputs(2957) <= not((inputs(166)) and (inputs(107)));
    layer0_outputs(2958) <= (inputs(189)) and not (inputs(49));
    layer0_outputs(2959) <= (inputs(97)) or (inputs(251));
    layer0_outputs(2960) <= (inputs(70)) and not (inputs(17));
    layer0_outputs(2961) <= '1';
    layer0_outputs(2962) <= (inputs(92)) and (inputs(215));
    layer0_outputs(2963) <= not(inputs(178));
    layer0_outputs(2964) <= not((inputs(237)) xor (inputs(20)));
    layer0_outputs(2965) <= (inputs(200)) or (inputs(152));
    layer0_outputs(2966) <= not(inputs(96));
    layer0_outputs(2967) <= (inputs(128)) or (inputs(75));
    layer0_outputs(2968) <= '0';
    layer0_outputs(2969) <= '0';
    layer0_outputs(2970) <= (inputs(100)) and (inputs(244));
    layer0_outputs(2971) <= '1';
    layer0_outputs(2972) <= not((inputs(209)) or (inputs(115)));
    layer0_outputs(2973) <= inputs(48);
    layer0_outputs(2974) <= inputs(111);
    layer0_outputs(2975) <= (inputs(193)) and (inputs(220));
    layer0_outputs(2976) <= (inputs(84)) or (inputs(15));
    layer0_outputs(2977) <= '0';
    layer0_outputs(2978) <= (inputs(205)) and not (inputs(114));
    layer0_outputs(2979) <= not(inputs(2));
    layer0_outputs(2980) <= not(inputs(26));
    layer0_outputs(2981) <= '1';
    layer0_outputs(2982) <= '0';
    layer0_outputs(2983) <= '0';
    layer0_outputs(2984) <= (inputs(255)) and not (inputs(197));
    layer0_outputs(2985) <= '1';
    layer0_outputs(2986) <= inputs(93);
    layer0_outputs(2987) <= (inputs(164)) and not (inputs(7));
    layer0_outputs(2988) <= '0';
    layer0_outputs(2989) <= '0';
    layer0_outputs(2990) <= '1';
    layer0_outputs(2991) <= (inputs(211)) or (inputs(218));
    layer0_outputs(2992) <= not((inputs(5)) and (inputs(216)));
    layer0_outputs(2993) <= inputs(139);
    layer0_outputs(2994) <= (inputs(124)) and not (inputs(231));
    layer0_outputs(2995) <= (inputs(92)) or (inputs(66));
    layer0_outputs(2996) <= not(inputs(236));
    layer0_outputs(2997) <= inputs(48);
    layer0_outputs(2998) <= (inputs(74)) and not (inputs(250));
    layer0_outputs(2999) <= (inputs(196)) and not (inputs(68));
    layer0_outputs(3000) <= not(inputs(193));
    layer0_outputs(3001) <= (inputs(13)) and (inputs(246));
    layer0_outputs(3002) <= (inputs(33)) and not (inputs(40));
    layer0_outputs(3003) <= '1';
    layer0_outputs(3004) <= '1';
    layer0_outputs(3005) <= '1';
    layer0_outputs(3006) <= (inputs(100)) and not (inputs(206));
    layer0_outputs(3007) <= not(inputs(142)) or (inputs(214));
    layer0_outputs(3008) <= (inputs(250)) and (inputs(177));
    layer0_outputs(3009) <= not(inputs(39)) or (inputs(75));
    layer0_outputs(3010) <= '1';
    layer0_outputs(3011) <= not((inputs(140)) xor (inputs(1)));
    layer0_outputs(3012) <= '1';
    layer0_outputs(3013) <= '0';
    layer0_outputs(3014) <= inputs(167);
    layer0_outputs(3015) <= inputs(109);
    layer0_outputs(3016) <= (inputs(82)) and not (inputs(43));
    layer0_outputs(3017) <= '1';
    layer0_outputs(3018) <= (inputs(213)) or (inputs(175));
    layer0_outputs(3019) <= '1';
    layer0_outputs(3020) <= not((inputs(7)) or (inputs(121)));
    layer0_outputs(3021) <= inputs(115);
    layer0_outputs(3022) <= (inputs(83)) or (inputs(171));
    layer0_outputs(3023) <= (inputs(88)) or (inputs(22));
    layer0_outputs(3024) <= not(inputs(24));
    layer0_outputs(3025) <= (inputs(174)) or (inputs(202));
    layer0_outputs(3026) <= (inputs(204)) and not (inputs(20));
    layer0_outputs(3027) <= not(inputs(195)) or (inputs(29));
    layer0_outputs(3028) <= '0';
    layer0_outputs(3029) <= '0';
    layer0_outputs(3030) <= (inputs(23)) and not (inputs(146));
    layer0_outputs(3031) <= (inputs(164)) and not (inputs(45));
    layer0_outputs(3032) <= not(inputs(52)) or (inputs(67));
    layer0_outputs(3033) <= '0';
    layer0_outputs(3034) <= not(inputs(34)) or (inputs(26));
    layer0_outputs(3035) <= (inputs(181)) and not (inputs(195));
    layer0_outputs(3036) <= inputs(178);
    layer0_outputs(3037) <= '0';
    layer0_outputs(3038) <= not(inputs(49));
    layer0_outputs(3039) <= inputs(164);
    layer0_outputs(3040) <= not(inputs(146));
    layer0_outputs(3041) <= '0';
    layer0_outputs(3042) <= not(inputs(195)) or (inputs(247));
    layer0_outputs(3043) <= (inputs(6)) and not (inputs(200));
    layer0_outputs(3044) <= '0';
    layer0_outputs(3045) <= '0';
    layer0_outputs(3046) <= not(inputs(234)) or (inputs(225));
    layer0_outputs(3047) <= (inputs(111)) and (inputs(175));
    layer0_outputs(3048) <= inputs(169);
    layer0_outputs(3049) <= not(inputs(13)) or (inputs(201));
    layer0_outputs(3050) <= inputs(80);
    layer0_outputs(3051) <= inputs(121);
    layer0_outputs(3052) <= '1';
    layer0_outputs(3053) <= '0';
    layer0_outputs(3054) <= (inputs(55)) and not (inputs(133));
    layer0_outputs(3055) <= not(inputs(9)) or (inputs(176));
    layer0_outputs(3056) <= '1';
    layer0_outputs(3057) <= '1';
    layer0_outputs(3058) <= not((inputs(49)) and (inputs(216)));
    layer0_outputs(3059) <= '0';
    layer0_outputs(3060) <= not(inputs(113)) or (inputs(150));
    layer0_outputs(3061) <= not(inputs(208)) or (inputs(8));
    layer0_outputs(3062) <= inputs(101);
    layer0_outputs(3063) <= not(inputs(110));
    layer0_outputs(3064) <= not((inputs(214)) and (inputs(146)));
    layer0_outputs(3065) <= (inputs(73)) and not (inputs(149));
    layer0_outputs(3066) <= not(inputs(97));
    layer0_outputs(3067) <= not((inputs(111)) xor (inputs(238)));
    layer0_outputs(3068) <= (inputs(201)) and (inputs(145));
    layer0_outputs(3069) <= (inputs(94)) or (inputs(195));
    layer0_outputs(3070) <= not(inputs(133));
    layer0_outputs(3071) <= '0';
    layer0_outputs(3072) <= not(inputs(87));
    layer0_outputs(3073) <= not(inputs(112));
    layer0_outputs(3074) <= not((inputs(85)) and (inputs(9)));
    layer0_outputs(3075) <= '1';
    layer0_outputs(3076) <= inputs(68);
    layer0_outputs(3077) <= not((inputs(235)) or (inputs(125)));
    layer0_outputs(3078) <= not((inputs(45)) or (inputs(23)));
    layer0_outputs(3079) <= (inputs(238)) and not (inputs(217));
    layer0_outputs(3080) <= not((inputs(245)) and (inputs(15)));
    layer0_outputs(3081) <= (inputs(213)) and not (inputs(119));
    layer0_outputs(3082) <= (inputs(248)) or (inputs(208));
    layer0_outputs(3083) <= not((inputs(43)) xor (inputs(134)));
    layer0_outputs(3084) <= '0';
    layer0_outputs(3085) <= not(inputs(231));
    layer0_outputs(3086) <= not(inputs(39)) or (inputs(36));
    layer0_outputs(3087) <= not((inputs(18)) and (inputs(228)));
    layer0_outputs(3088) <= inputs(142);
    layer0_outputs(3089) <= (inputs(48)) or (inputs(107));
    layer0_outputs(3090) <= '0';
    layer0_outputs(3091) <= not(inputs(143));
    layer0_outputs(3092) <= '0';
    layer0_outputs(3093) <= '1';
    layer0_outputs(3094) <= not(inputs(24));
    layer0_outputs(3095) <= '1';
    layer0_outputs(3096) <= not((inputs(37)) or (inputs(235)));
    layer0_outputs(3097) <= (inputs(165)) and not (inputs(32));
    layer0_outputs(3098) <= not((inputs(19)) or (inputs(169)));
    layer0_outputs(3099) <= '0';
    layer0_outputs(3100) <= '1';
    layer0_outputs(3101) <= not(inputs(187)) or (inputs(149));
    layer0_outputs(3102) <= inputs(228);
    layer0_outputs(3103) <= '1';
    layer0_outputs(3104) <= inputs(166);
    layer0_outputs(3105) <= not((inputs(218)) or (inputs(177)));
    layer0_outputs(3106) <= (inputs(6)) and not (inputs(2));
    layer0_outputs(3107) <= (inputs(28)) and (inputs(13));
    layer0_outputs(3108) <= not(inputs(60)) or (inputs(48));
    layer0_outputs(3109) <= '1';
    layer0_outputs(3110) <= inputs(55);
    layer0_outputs(3111) <= '1';
    layer0_outputs(3112) <= (inputs(162)) xor (inputs(119));
    layer0_outputs(3113) <= (inputs(48)) or (inputs(210));
    layer0_outputs(3114) <= inputs(172);
    layer0_outputs(3115) <= '0';
    layer0_outputs(3116) <= inputs(179);
    layer0_outputs(3117) <= inputs(143);
    layer0_outputs(3118) <= (inputs(71)) and not (inputs(174));
    layer0_outputs(3119) <= '1';
    layer0_outputs(3120) <= (inputs(167)) or (inputs(58));
    layer0_outputs(3121) <= (inputs(124)) and (inputs(50));
    layer0_outputs(3122) <= not(inputs(202)) or (inputs(225));
    layer0_outputs(3123) <= not((inputs(233)) xor (inputs(161)));
    layer0_outputs(3124) <= not(inputs(214));
    layer0_outputs(3125) <= (inputs(126)) or (inputs(91));
    layer0_outputs(3126) <= not(inputs(21));
    layer0_outputs(3127) <= '1';
    layer0_outputs(3128) <= (inputs(23)) xor (inputs(55));
    layer0_outputs(3129) <= (inputs(182)) and not (inputs(127));
    layer0_outputs(3130) <= '0';
    layer0_outputs(3131) <= (inputs(47)) and not (inputs(20));
    layer0_outputs(3132) <= '0';
    layer0_outputs(3133) <= not((inputs(227)) or (inputs(211)));
    layer0_outputs(3134) <= '1';
    layer0_outputs(3135) <= not(inputs(14));
    layer0_outputs(3136) <= inputs(249);
    layer0_outputs(3137) <= (inputs(53)) or (inputs(81));
    layer0_outputs(3138) <= (inputs(223)) or (inputs(79));
    layer0_outputs(3139) <= '1';
    layer0_outputs(3140) <= not(inputs(216)) or (inputs(140));
    layer0_outputs(3141) <= '0';
    layer0_outputs(3142) <= not(inputs(140)) or (inputs(50));
    layer0_outputs(3143) <= '0';
    layer0_outputs(3144) <= not((inputs(253)) or (inputs(32)));
    layer0_outputs(3145) <= (inputs(28)) and not (inputs(146));
    layer0_outputs(3146) <= inputs(137);
    layer0_outputs(3147) <= not((inputs(220)) and (inputs(148)));
    layer0_outputs(3148) <= (inputs(90)) and (inputs(42));
    layer0_outputs(3149) <= '0';
    layer0_outputs(3150) <= '0';
    layer0_outputs(3151) <= (inputs(25)) or (inputs(222));
    layer0_outputs(3152) <= not(inputs(62)) or (inputs(234));
    layer0_outputs(3153) <= not((inputs(179)) and (inputs(253)));
    layer0_outputs(3154) <= (inputs(152)) and not (inputs(196));
    layer0_outputs(3155) <= (inputs(71)) and not (inputs(214));
    layer0_outputs(3156) <= inputs(63);
    layer0_outputs(3157) <= not(inputs(110));
    layer0_outputs(3158) <= inputs(161);
    layer0_outputs(3159) <= '0';
    layer0_outputs(3160) <= '0';
    layer0_outputs(3161) <= (inputs(177)) or (inputs(182));
    layer0_outputs(3162) <= '0';
    layer0_outputs(3163) <= '1';
    layer0_outputs(3164) <= not(inputs(223));
    layer0_outputs(3165) <= not(inputs(79)) or (inputs(83));
    layer0_outputs(3166) <= not((inputs(204)) and (inputs(150)));
    layer0_outputs(3167) <= not(inputs(39));
    layer0_outputs(3168) <= not((inputs(102)) and (inputs(49)));
    layer0_outputs(3169) <= (inputs(124)) and (inputs(193));
    layer0_outputs(3170) <= not(inputs(187)) or (inputs(209));
    layer0_outputs(3171) <= not((inputs(252)) or (inputs(203)));
    layer0_outputs(3172) <= not((inputs(29)) and (inputs(159)));
    layer0_outputs(3173) <= not(inputs(197));
    layer0_outputs(3174) <= not(inputs(125));
    layer0_outputs(3175) <= not((inputs(181)) and (inputs(228)));
    layer0_outputs(3176) <= not(inputs(84)) or (inputs(87));
    layer0_outputs(3177) <= (inputs(220)) xor (inputs(62));
    layer0_outputs(3178) <= '1';
    layer0_outputs(3179) <= not(inputs(236)) or (inputs(126));
    layer0_outputs(3180) <= '1';
    layer0_outputs(3181) <= not(inputs(17));
    layer0_outputs(3182) <= not(inputs(151)) or (inputs(142));
    layer0_outputs(3183) <= (inputs(33)) and (inputs(93));
    layer0_outputs(3184) <= not(inputs(233)) or (inputs(23));
    layer0_outputs(3185) <= inputs(152);
    layer0_outputs(3186) <= not((inputs(192)) or (inputs(132)));
    layer0_outputs(3187) <= '0';
    layer0_outputs(3188) <= '0';
    layer0_outputs(3189) <= (inputs(147)) and not (inputs(65));
    layer0_outputs(3190) <= (inputs(69)) or (inputs(163));
    layer0_outputs(3191) <= (inputs(155)) and not (inputs(84));
    layer0_outputs(3192) <= '1';
    layer0_outputs(3193) <= not(inputs(239)) or (inputs(198));
    layer0_outputs(3194) <= (inputs(97)) and (inputs(84));
    layer0_outputs(3195) <= (inputs(204)) or (inputs(120));
    layer0_outputs(3196) <= not((inputs(202)) or (inputs(100)));
    layer0_outputs(3197) <= (inputs(158)) or (inputs(218));
    layer0_outputs(3198) <= not(inputs(26));
    layer0_outputs(3199) <= '1';
    layer0_outputs(3200) <= inputs(247);
    layer0_outputs(3201) <= not(inputs(237));
    layer0_outputs(3202) <= '0';
    layer0_outputs(3203) <= not(inputs(71));
    layer0_outputs(3204) <= (inputs(223)) xor (inputs(105));
    layer0_outputs(3205) <= not(inputs(211)) or (inputs(143));
    layer0_outputs(3206) <= '0';
    layer0_outputs(3207) <= (inputs(192)) or (inputs(135));
    layer0_outputs(3208) <= '1';
    layer0_outputs(3209) <= (inputs(165)) and not (inputs(72));
    layer0_outputs(3210) <= not((inputs(175)) or (inputs(81)));
    layer0_outputs(3211) <= not((inputs(49)) and (inputs(176)));
    layer0_outputs(3212) <= '0';
    layer0_outputs(3213) <= (inputs(9)) and not (inputs(161));
    layer0_outputs(3214) <= '1';
    layer0_outputs(3215) <= '0';
    layer0_outputs(3216) <= not(inputs(138));
    layer0_outputs(3217) <= not(inputs(99));
    layer0_outputs(3218) <= (inputs(58)) and (inputs(187));
    layer0_outputs(3219) <= (inputs(176)) and not (inputs(244));
    layer0_outputs(3220) <= '0';
    layer0_outputs(3221) <= not(inputs(64)) or (inputs(103));
    layer0_outputs(3222) <= not(inputs(188)) or (inputs(103));
    layer0_outputs(3223) <= not(inputs(207));
    layer0_outputs(3224) <= not(inputs(248));
    layer0_outputs(3225) <= inputs(100);
    layer0_outputs(3226) <= '0';
    layer0_outputs(3227) <= '0';
    layer0_outputs(3228) <= not((inputs(148)) or (inputs(220)));
    layer0_outputs(3229) <= '1';
    layer0_outputs(3230) <= '0';
    layer0_outputs(3231) <= not(inputs(199)) or (inputs(187));
    layer0_outputs(3232) <= '0';
    layer0_outputs(3233) <= '1';
    layer0_outputs(3234) <= '0';
    layer0_outputs(3235) <= (inputs(169)) or (inputs(223));
    layer0_outputs(3236) <= (inputs(185)) and (inputs(205));
    layer0_outputs(3237) <= '0';
    layer0_outputs(3238) <= '1';
    layer0_outputs(3239) <= not((inputs(20)) and (inputs(108)));
    layer0_outputs(3240) <= '1';
    layer0_outputs(3241) <= (inputs(245)) or (inputs(158));
    layer0_outputs(3242) <= not(inputs(151));
    layer0_outputs(3243) <= (inputs(87)) and not (inputs(251));
    layer0_outputs(3244) <= '1';
    layer0_outputs(3245) <= not((inputs(9)) and (inputs(169)));
    layer0_outputs(3246) <= (inputs(112)) and (inputs(209));
    layer0_outputs(3247) <= (inputs(252)) and not (inputs(191));
    layer0_outputs(3248) <= not((inputs(157)) and (inputs(163)));
    layer0_outputs(3249) <= not(inputs(106));
    layer0_outputs(3250) <= '1';
    layer0_outputs(3251) <= inputs(17);
    layer0_outputs(3252) <= not(inputs(100));
    layer0_outputs(3253) <= inputs(255);
    layer0_outputs(3254) <= inputs(209);
    layer0_outputs(3255) <= inputs(95);
    layer0_outputs(3256) <= not((inputs(77)) or (inputs(177)));
    layer0_outputs(3257) <= not(inputs(44)) or (inputs(7));
    layer0_outputs(3258) <= '0';
    layer0_outputs(3259) <= (inputs(218)) or (inputs(181));
    layer0_outputs(3260) <= (inputs(164)) or (inputs(108));
    layer0_outputs(3261) <= inputs(187);
    layer0_outputs(3262) <= inputs(147);
    layer0_outputs(3263) <= inputs(57);
    layer0_outputs(3264) <= (inputs(200)) or (inputs(160));
    layer0_outputs(3265) <= inputs(94);
    layer0_outputs(3266) <= (inputs(19)) and not (inputs(144));
    layer0_outputs(3267) <= not(inputs(150));
    layer0_outputs(3268) <= not((inputs(145)) or (inputs(28)));
    layer0_outputs(3269) <= (inputs(180)) or (inputs(179));
    layer0_outputs(3270) <= '1';
    layer0_outputs(3271) <= not((inputs(250)) or (inputs(204)));
    layer0_outputs(3272) <= '0';
    layer0_outputs(3273) <= inputs(16);
    layer0_outputs(3274) <= (inputs(201)) and not (inputs(2));
    layer0_outputs(3275) <= '0';
    layer0_outputs(3276) <= inputs(212);
    layer0_outputs(3277) <= not(inputs(119)) or (inputs(67));
    layer0_outputs(3278) <= (inputs(21)) and (inputs(84));
    layer0_outputs(3279) <= inputs(221);
    layer0_outputs(3280) <= '0';
    layer0_outputs(3281) <= not(inputs(83)) or (inputs(62));
    layer0_outputs(3282) <= not(inputs(152));
    layer0_outputs(3283) <= (inputs(128)) and not (inputs(163));
    layer0_outputs(3284) <= not(inputs(223)) or (inputs(244));
    layer0_outputs(3285) <= not((inputs(150)) and (inputs(38)));
    layer0_outputs(3286) <= not(inputs(171));
    layer0_outputs(3287) <= '0';
    layer0_outputs(3288) <= '1';
    layer0_outputs(3289) <= not(inputs(137));
    layer0_outputs(3290) <= not((inputs(219)) and (inputs(141)));
    layer0_outputs(3291) <= (inputs(202)) or (inputs(60));
    layer0_outputs(3292) <= (inputs(255)) and not (inputs(181));
    layer0_outputs(3293) <= '1';
    layer0_outputs(3294) <= (inputs(231)) xor (inputs(213));
    layer0_outputs(3295) <= not((inputs(81)) or (inputs(179)));
    layer0_outputs(3296) <= not(inputs(72)) or (inputs(17));
    layer0_outputs(3297) <= not((inputs(74)) xor (inputs(78)));
    layer0_outputs(3298) <= not(inputs(21));
    layer0_outputs(3299) <= (inputs(92)) and (inputs(182));
    layer0_outputs(3300) <= inputs(15);
    layer0_outputs(3301) <= not(inputs(37));
    layer0_outputs(3302) <= (inputs(60)) or (inputs(146));
    layer0_outputs(3303) <= (inputs(94)) and (inputs(20));
    layer0_outputs(3304) <= not(inputs(89)) or (inputs(20));
    layer0_outputs(3305) <= not(inputs(74)) or (inputs(151));
    layer0_outputs(3306) <= inputs(218);
    layer0_outputs(3307) <= inputs(102);
    layer0_outputs(3308) <= (inputs(89)) or (inputs(137));
    layer0_outputs(3309) <= '0';
    layer0_outputs(3310) <= '1';
    layer0_outputs(3311) <= (inputs(169)) and (inputs(79));
    layer0_outputs(3312) <= '0';
    layer0_outputs(3313) <= (inputs(168)) and not (inputs(236));
    layer0_outputs(3314) <= not(inputs(94));
    layer0_outputs(3315) <= not(inputs(116));
    layer0_outputs(3316) <= not(inputs(236));
    layer0_outputs(3317) <= not(inputs(165)) or (inputs(5));
    layer0_outputs(3318) <= not(inputs(180));
    layer0_outputs(3319) <= inputs(13);
    layer0_outputs(3320) <= (inputs(116)) or (inputs(66));
    layer0_outputs(3321) <= '0';
    layer0_outputs(3322) <= '0';
    layer0_outputs(3323) <= not(inputs(194));
    layer0_outputs(3324) <= '0';
    layer0_outputs(3325) <= (inputs(240)) and not (inputs(54));
    layer0_outputs(3326) <= not(inputs(1));
    layer0_outputs(3327) <= not(inputs(91)) or (inputs(177));
    layer0_outputs(3328) <= (inputs(111)) and (inputs(186));
    layer0_outputs(3329) <= '0';
    layer0_outputs(3330) <= inputs(122);
    layer0_outputs(3331) <= '0';
    layer0_outputs(3332) <= inputs(232);
    layer0_outputs(3333) <= '0';
    layer0_outputs(3334) <= not(inputs(25));
    layer0_outputs(3335) <= not((inputs(139)) and (inputs(93)));
    layer0_outputs(3336) <= not(inputs(46)) or (inputs(123));
    layer0_outputs(3337) <= (inputs(48)) and (inputs(96));
    layer0_outputs(3338) <= '1';
    layer0_outputs(3339) <= '0';
    layer0_outputs(3340) <= '0';
    layer0_outputs(3341) <= (inputs(5)) and (inputs(44));
    layer0_outputs(3342) <= not(inputs(104));
    layer0_outputs(3343) <= '1';
    layer0_outputs(3344) <= (inputs(29)) and (inputs(102));
    layer0_outputs(3345) <= '0';
    layer0_outputs(3346) <= (inputs(115)) or (inputs(82));
    layer0_outputs(3347) <= (inputs(227)) and (inputs(169));
    layer0_outputs(3348) <= (inputs(210)) xor (inputs(95));
    layer0_outputs(3349) <= '0';
    layer0_outputs(3350) <= inputs(24);
    layer0_outputs(3351) <= '0';
    layer0_outputs(3352) <= inputs(134);
    layer0_outputs(3353) <= (inputs(61)) or (inputs(32));
    layer0_outputs(3354) <= not(inputs(84));
    layer0_outputs(3355) <= not(inputs(2)) or (inputs(197));
    layer0_outputs(3356) <= not(inputs(64));
    layer0_outputs(3357) <= (inputs(174)) and (inputs(42));
    layer0_outputs(3358) <= (inputs(220)) and (inputs(191));
    layer0_outputs(3359) <= '0';
    layer0_outputs(3360) <= inputs(37);
    layer0_outputs(3361) <= not(inputs(75));
    layer0_outputs(3362) <= inputs(108);
    layer0_outputs(3363) <= (inputs(142)) and (inputs(112));
    layer0_outputs(3364) <= (inputs(78)) and (inputs(239));
    layer0_outputs(3365) <= inputs(195);
    layer0_outputs(3366) <= '0';
    layer0_outputs(3367) <= not((inputs(160)) and (inputs(71)));
    layer0_outputs(3368) <= '0';
    layer0_outputs(3369) <= '1';
    layer0_outputs(3370) <= (inputs(59)) and not (inputs(24));
    layer0_outputs(3371) <= inputs(172);
    layer0_outputs(3372) <= not((inputs(54)) or (inputs(246)));
    layer0_outputs(3373) <= inputs(162);
    layer0_outputs(3374) <= (inputs(232)) and not (inputs(52));
    layer0_outputs(3375) <= '0';
    layer0_outputs(3376) <= not((inputs(232)) or (inputs(42)));
    layer0_outputs(3377) <= '0';
    layer0_outputs(3378) <= inputs(40);
    layer0_outputs(3379) <= not(inputs(123)) or (inputs(142));
    layer0_outputs(3380) <= (inputs(20)) or (inputs(5));
    layer0_outputs(3381) <= not(inputs(36)) or (inputs(117));
    layer0_outputs(3382) <= (inputs(22)) and not (inputs(249));
    layer0_outputs(3383) <= '1';
    layer0_outputs(3384) <= not((inputs(253)) or (inputs(35)));
    layer0_outputs(3385) <= not(inputs(139)) or (inputs(91));
    layer0_outputs(3386) <= (inputs(7)) or (inputs(207));
    layer0_outputs(3387) <= not((inputs(16)) or (inputs(138)));
    layer0_outputs(3388) <= (inputs(0)) or (inputs(107));
    layer0_outputs(3389) <= (inputs(206)) and (inputs(216));
    layer0_outputs(3390) <= '0';
    layer0_outputs(3391) <= not(inputs(182));
    layer0_outputs(3392) <= inputs(218);
    layer0_outputs(3393) <= not(inputs(114));
    layer0_outputs(3394) <= not((inputs(39)) or (inputs(43)));
    layer0_outputs(3395) <= not((inputs(138)) or (inputs(190)));
    layer0_outputs(3396) <= (inputs(132)) or (inputs(162));
    layer0_outputs(3397) <= not(inputs(145)) or (inputs(62));
    layer0_outputs(3398) <= '0';
    layer0_outputs(3399) <= not((inputs(207)) or (inputs(107)));
    layer0_outputs(3400) <= (inputs(153)) and (inputs(226));
    layer0_outputs(3401) <= not(inputs(64)) or (inputs(106));
    layer0_outputs(3402) <= inputs(164);
    layer0_outputs(3403) <= '0';
    layer0_outputs(3404) <= not(inputs(77));
    layer0_outputs(3405) <= not(inputs(227)) or (inputs(39));
    layer0_outputs(3406) <= not((inputs(61)) or (inputs(57)));
    layer0_outputs(3407) <= '1';
    layer0_outputs(3408) <= (inputs(131)) and not (inputs(199));
    layer0_outputs(3409) <= not(inputs(82));
    layer0_outputs(3410) <= (inputs(19)) and not (inputs(244));
    layer0_outputs(3411) <= inputs(164);
    layer0_outputs(3412) <= '1';
    layer0_outputs(3413) <= '0';
    layer0_outputs(3414) <= '0';
    layer0_outputs(3415) <= '1';
    layer0_outputs(3416) <= inputs(252);
    layer0_outputs(3417) <= not(inputs(140)) or (inputs(31));
    layer0_outputs(3418) <= (inputs(209)) or (inputs(192));
    layer0_outputs(3419) <= not(inputs(35));
    layer0_outputs(3420) <= (inputs(157)) or (inputs(45));
    layer0_outputs(3421) <= not(inputs(246)) or (inputs(58));
    layer0_outputs(3422) <= not(inputs(37));
    layer0_outputs(3423) <= not(inputs(226));
    layer0_outputs(3424) <= (inputs(2)) and not (inputs(194));
    layer0_outputs(3425) <= not(inputs(245)) or (inputs(197));
    layer0_outputs(3426) <= not((inputs(76)) or (inputs(187)));
    layer0_outputs(3427) <= not(inputs(41)) or (inputs(90));
    layer0_outputs(3428) <= '0';
    layer0_outputs(3429) <= '1';
    layer0_outputs(3430) <= not(inputs(239)) or (inputs(56));
    layer0_outputs(3431) <= not(inputs(182)) or (inputs(145));
    layer0_outputs(3432) <= (inputs(249)) or (inputs(176));
    layer0_outputs(3433) <= '1';
    layer0_outputs(3434) <= not(inputs(229)) or (inputs(181));
    layer0_outputs(3435) <= not(inputs(80));
    layer0_outputs(3436) <= '0';
    layer0_outputs(3437) <= not((inputs(141)) and (inputs(119)));
    layer0_outputs(3438) <= not(inputs(235));
    layer0_outputs(3439) <= inputs(196);
    layer0_outputs(3440) <= (inputs(192)) and not (inputs(173));
    layer0_outputs(3441) <= not(inputs(7));
    layer0_outputs(3442) <= not((inputs(97)) xor (inputs(3)));
    layer0_outputs(3443) <= '0';
    layer0_outputs(3444) <= '1';
    layer0_outputs(3445) <= (inputs(85)) and not (inputs(33));
    layer0_outputs(3446) <= '0';
    layer0_outputs(3447) <= '1';
    layer0_outputs(3448) <= '1';
    layer0_outputs(3449) <= (inputs(149)) or (inputs(106));
    layer0_outputs(3450) <= '1';
    layer0_outputs(3451) <= not(inputs(120));
    layer0_outputs(3452) <= '0';
    layer0_outputs(3453) <= (inputs(157)) and not (inputs(49));
    layer0_outputs(3454) <= not(inputs(60));
    layer0_outputs(3455) <= (inputs(102)) or (inputs(132));
    layer0_outputs(3456) <= not((inputs(165)) or (inputs(149)));
    layer0_outputs(3457) <= '1';
    layer0_outputs(3458) <= not((inputs(87)) and (inputs(13)));
    layer0_outputs(3459) <= inputs(178);
    layer0_outputs(3460) <= not((inputs(209)) and (inputs(76)));
    layer0_outputs(3461) <= not(inputs(107));
    layer0_outputs(3462) <= (inputs(21)) or (inputs(226));
    layer0_outputs(3463) <= (inputs(108)) and (inputs(220));
    layer0_outputs(3464) <= '0';
    layer0_outputs(3465) <= (inputs(232)) and not (inputs(103));
    layer0_outputs(3466) <= (inputs(144)) and not (inputs(151));
    layer0_outputs(3467) <= (inputs(242)) and not (inputs(163));
    layer0_outputs(3468) <= not(inputs(82)) or (inputs(152));
    layer0_outputs(3469) <= inputs(82);
    layer0_outputs(3470) <= '0';
    layer0_outputs(3471) <= not(inputs(155)) or (inputs(17));
    layer0_outputs(3472) <= '0';
    layer0_outputs(3473) <= not(inputs(210)) or (inputs(220));
    layer0_outputs(3474) <= (inputs(172)) and (inputs(65));
    layer0_outputs(3475) <= not(inputs(113)) or (inputs(83));
    layer0_outputs(3476) <= not((inputs(106)) or (inputs(217)));
    layer0_outputs(3477) <= not(inputs(114)) or (inputs(57));
    layer0_outputs(3478) <= (inputs(27)) and not (inputs(156));
    layer0_outputs(3479) <= inputs(228);
    layer0_outputs(3480) <= not(inputs(223));
    layer0_outputs(3481) <= inputs(237);
    layer0_outputs(3482) <= inputs(109);
    layer0_outputs(3483) <= (inputs(69)) and not (inputs(216));
    layer0_outputs(3484) <= not((inputs(144)) and (inputs(207)));
    layer0_outputs(3485) <= '0';
    layer0_outputs(3486) <= '0';
    layer0_outputs(3487) <= (inputs(232)) and not (inputs(234));
    layer0_outputs(3488) <= '0';
    layer0_outputs(3489) <= inputs(134);
    layer0_outputs(3490) <= '0';
    layer0_outputs(3491) <= '0';
    layer0_outputs(3492) <= '0';
    layer0_outputs(3493) <= '0';
    layer0_outputs(3494) <= (inputs(219)) and not (inputs(140));
    layer0_outputs(3495) <= not(inputs(6));
    layer0_outputs(3496) <= '1';
    layer0_outputs(3497) <= '1';
    layer0_outputs(3498) <= '1';
    layer0_outputs(3499) <= not(inputs(116));
    layer0_outputs(3500) <= not((inputs(218)) or (inputs(118)));
    layer0_outputs(3501) <= not(inputs(174)) or (inputs(113));
    layer0_outputs(3502) <= '1';
    layer0_outputs(3503) <= not(inputs(29)) or (inputs(10));
    layer0_outputs(3504) <= (inputs(146)) and not (inputs(192));
    layer0_outputs(3505) <= not(inputs(193));
    layer0_outputs(3506) <= (inputs(59)) and not (inputs(14));
    layer0_outputs(3507) <= '1';
    layer0_outputs(3508) <= not(inputs(10));
    layer0_outputs(3509) <= '1';
    layer0_outputs(3510) <= inputs(162);
    layer0_outputs(3511) <= '0';
    layer0_outputs(3512) <= (inputs(83)) and not (inputs(77));
    layer0_outputs(3513) <= '1';
    layer0_outputs(3514) <= (inputs(254)) or (inputs(114));
    layer0_outputs(3515) <= '1';
    layer0_outputs(3516) <= '1';
    layer0_outputs(3517) <= not(inputs(251)) or (inputs(13));
    layer0_outputs(3518) <= '0';
    layer0_outputs(3519) <= not((inputs(107)) and (inputs(204)));
    layer0_outputs(3520) <= (inputs(127)) and not (inputs(91));
    layer0_outputs(3521) <= not((inputs(156)) and (inputs(189)));
    layer0_outputs(3522) <= (inputs(44)) and (inputs(14));
    layer0_outputs(3523) <= not(inputs(188));
    layer0_outputs(3524) <= not(inputs(97));
    layer0_outputs(3525) <= (inputs(99)) and (inputs(64));
    layer0_outputs(3526) <= '1';
    layer0_outputs(3527) <= (inputs(168)) and not (inputs(142));
    layer0_outputs(3528) <= not((inputs(132)) xor (inputs(166)));
    layer0_outputs(3529) <= inputs(214);
    layer0_outputs(3530) <= not(inputs(195));
    layer0_outputs(3531) <= not((inputs(148)) and (inputs(113)));
    layer0_outputs(3532) <= '0';
    layer0_outputs(3533) <= not(inputs(201)) or (inputs(92));
    layer0_outputs(3534) <= inputs(206);
    layer0_outputs(3535) <= (inputs(189)) and (inputs(125));
    layer0_outputs(3536) <= (inputs(181)) and (inputs(228));
    layer0_outputs(3537) <= not(inputs(1)) or (inputs(164));
    layer0_outputs(3538) <= not(inputs(162));
    layer0_outputs(3539) <= not((inputs(88)) xor (inputs(20)));
    layer0_outputs(3540) <= '1';
    layer0_outputs(3541) <= not((inputs(255)) and (inputs(60)));
    layer0_outputs(3542) <= (inputs(112)) or (inputs(147));
    layer0_outputs(3543) <= (inputs(126)) or (inputs(101));
    layer0_outputs(3544) <= (inputs(200)) xor (inputs(248));
    layer0_outputs(3545) <= '1';
    layer0_outputs(3546) <= '0';
    layer0_outputs(3547) <= inputs(74);
    layer0_outputs(3548) <= not(inputs(36)) or (inputs(37));
    layer0_outputs(3549) <= not(inputs(46));
    layer0_outputs(3550) <= (inputs(117)) or (inputs(67));
    layer0_outputs(3551) <= (inputs(147)) or (inputs(187));
    layer0_outputs(3552) <= (inputs(82)) and not (inputs(225));
    layer0_outputs(3553) <= not(inputs(139)) or (inputs(27));
    layer0_outputs(3554) <= not(inputs(92));
    layer0_outputs(3555) <= not(inputs(112));
    layer0_outputs(3556) <= '1';
    layer0_outputs(3557) <= '0';
    layer0_outputs(3558) <= '0';
    layer0_outputs(3559) <= inputs(81);
    layer0_outputs(3560) <= (inputs(158)) or (inputs(18));
    layer0_outputs(3561) <= not(inputs(83)) or (inputs(1));
    layer0_outputs(3562) <= not(inputs(128)) or (inputs(186));
    layer0_outputs(3563) <= '1';
    layer0_outputs(3564) <= '0';
    layer0_outputs(3565) <= (inputs(16)) and not (inputs(248));
    layer0_outputs(3566) <= not((inputs(238)) or (inputs(227)));
    layer0_outputs(3567) <= not(inputs(82));
    layer0_outputs(3568) <= not(inputs(81)) or (inputs(6));
    layer0_outputs(3569) <= not((inputs(25)) or (inputs(95)));
    layer0_outputs(3570) <= not(inputs(182));
    layer0_outputs(3571) <= not(inputs(83));
    layer0_outputs(3572) <= not(inputs(48));
    layer0_outputs(3573) <= (inputs(240)) and (inputs(59));
    layer0_outputs(3574) <= (inputs(166)) and (inputs(7));
    layer0_outputs(3575) <= '1';
    layer0_outputs(3576) <= not((inputs(244)) xor (inputs(232)));
    layer0_outputs(3577) <= not(inputs(147));
    layer0_outputs(3578) <= (inputs(131)) and not (inputs(134));
    layer0_outputs(3579) <= inputs(0);
    layer0_outputs(3580) <= inputs(58);
    layer0_outputs(3581) <= not(inputs(189)) or (inputs(233));
    layer0_outputs(3582) <= not(inputs(134));
    layer0_outputs(3583) <= (inputs(103)) or (inputs(27));
    layer0_outputs(3584) <= (inputs(149)) or (inputs(24));
    layer0_outputs(3585) <= not(inputs(103));
    layer0_outputs(3586) <= not(inputs(221)) or (inputs(221));
    layer0_outputs(3587) <= '1';
    layer0_outputs(3588) <= '0';
    layer0_outputs(3589) <= not((inputs(240)) and (inputs(178)));
    layer0_outputs(3590) <= '1';
    layer0_outputs(3591) <= '0';
    layer0_outputs(3592) <= '1';
    layer0_outputs(3593) <= '1';
    layer0_outputs(3594) <= not(inputs(108));
    layer0_outputs(3595) <= '0';
    layer0_outputs(3596) <= not(inputs(171));
    layer0_outputs(3597) <= '1';
    layer0_outputs(3598) <= inputs(111);
    layer0_outputs(3599) <= not(inputs(25)) or (inputs(230));
    layer0_outputs(3600) <= not(inputs(122));
    layer0_outputs(3601) <= (inputs(92)) and (inputs(66));
    layer0_outputs(3602) <= (inputs(61)) and not (inputs(91));
    layer0_outputs(3603) <= '1';
    layer0_outputs(3604) <= (inputs(71)) and (inputs(29));
    layer0_outputs(3605) <= not(inputs(203)) or (inputs(83));
    layer0_outputs(3606) <= not(inputs(213));
    layer0_outputs(3607) <= '1';
    layer0_outputs(3608) <= not(inputs(204));
    layer0_outputs(3609) <= inputs(16);
    layer0_outputs(3610) <= not(inputs(182)) or (inputs(104));
    layer0_outputs(3611) <= not(inputs(229));
    layer0_outputs(3612) <= (inputs(158)) xor (inputs(222));
    layer0_outputs(3613) <= (inputs(77)) and not (inputs(31));
    layer0_outputs(3614) <= not((inputs(229)) and (inputs(112)));
    layer0_outputs(3615) <= not((inputs(98)) and (inputs(174)));
    layer0_outputs(3616) <= not((inputs(123)) and (inputs(89)));
    layer0_outputs(3617) <= '0';
    layer0_outputs(3618) <= not(inputs(49)) or (inputs(7));
    layer0_outputs(3619) <= not(inputs(61)) or (inputs(167));
    layer0_outputs(3620) <= (inputs(33)) and not (inputs(80));
    layer0_outputs(3621) <= inputs(104);
    layer0_outputs(3622) <= inputs(128);
    layer0_outputs(3623) <= not(inputs(24));
    layer0_outputs(3624) <= '0';
    layer0_outputs(3625) <= '1';
    layer0_outputs(3626) <= (inputs(24)) and not (inputs(236));
    layer0_outputs(3627) <= inputs(69);
    layer0_outputs(3628) <= inputs(232);
    layer0_outputs(3629) <= not(inputs(18)) or (inputs(232));
    layer0_outputs(3630) <= not((inputs(127)) and (inputs(105)));
    layer0_outputs(3631) <= (inputs(136)) and not (inputs(87));
    layer0_outputs(3632) <= '0';
    layer0_outputs(3633) <= not(inputs(188));
    layer0_outputs(3634) <= '0';
    layer0_outputs(3635) <= (inputs(55)) or (inputs(30));
    layer0_outputs(3636) <= '1';
    layer0_outputs(3637) <= '1';
    layer0_outputs(3638) <= '1';
    layer0_outputs(3639) <= (inputs(57)) or (inputs(190));
    layer0_outputs(3640) <= inputs(27);
    layer0_outputs(3641) <= not(inputs(80));
    layer0_outputs(3642) <= not(inputs(101));
    layer0_outputs(3643) <= not((inputs(48)) or (inputs(105)));
    layer0_outputs(3644) <= inputs(223);
    layer0_outputs(3645) <= not(inputs(147));
    layer0_outputs(3646) <= '0';
    layer0_outputs(3647) <= inputs(209);
    layer0_outputs(3648) <= not(inputs(102));
    layer0_outputs(3649) <= not(inputs(226));
    layer0_outputs(3650) <= not(inputs(198)) or (inputs(75));
    layer0_outputs(3651) <= not(inputs(154)) or (inputs(108));
    layer0_outputs(3652) <= '1';
    layer0_outputs(3653) <= not((inputs(231)) xor (inputs(83)));
    layer0_outputs(3654) <= (inputs(231)) and (inputs(120));
    layer0_outputs(3655) <= not(inputs(11)) or (inputs(52));
    layer0_outputs(3656) <= '1';
    layer0_outputs(3657) <= not(inputs(108)) or (inputs(137));
    layer0_outputs(3658) <= '1';
    layer0_outputs(3659) <= not(inputs(124));
    layer0_outputs(3660) <= inputs(17);
    layer0_outputs(3661) <= (inputs(242)) or (inputs(212));
    layer0_outputs(3662) <= inputs(128);
    layer0_outputs(3663) <= inputs(29);
    layer0_outputs(3664) <= inputs(74);
    layer0_outputs(3665) <= '1';
    layer0_outputs(3666) <= (inputs(129)) and not (inputs(68));
    layer0_outputs(3667) <= not(inputs(168));
    layer0_outputs(3668) <= not((inputs(158)) or (inputs(131)));
    layer0_outputs(3669) <= '1';
    layer0_outputs(3670) <= (inputs(33)) and not (inputs(116));
    layer0_outputs(3671) <= (inputs(231)) or (inputs(224));
    layer0_outputs(3672) <= (inputs(195)) and not (inputs(100));
    layer0_outputs(3673) <= inputs(140);
    layer0_outputs(3674) <= not((inputs(218)) or (inputs(138)));
    layer0_outputs(3675) <= not((inputs(235)) and (inputs(54)));
    layer0_outputs(3676) <= (inputs(242)) and (inputs(186));
    layer0_outputs(3677) <= '1';
    layer0_outputs(3678) <= '0';
    layer0_outputs(3679) <= (inputs(144)) xor (inputs(84));
    layer0_outputs(3680) <= not((inputs(227)) and (inputs(183)));
    layer0_outputs(3681) <= not(inputs(194)) or (inputs(112));
    layer0_outputs(3682) <= (inputs(115)) and not (inputs(244));
    layer0_outputs(3683) <= not(inputs(76));
    layer0_outputs(3684) <= (inputs(156)) and (inputs(87));
    layer0_outputs(3685) <= not(inputs(26)) or (inputs(211));
    layer0_outputs(3686) <= '0';
    layer0_outputs(3687) <= (inputs(129)) or (inputs(225));
    layer0_outputs(3688) <= (inputs(92)) or (inputs(171));
    layer0_outputs(3689) <= '1';
    layer0_outputs(3690) <= (inputs(8)) and not (inputs(170));
    layer0_outputs(3691) <= (inputs(251)) or (inputs(188));
    layer0_outputs(3692) <= (inputs(236)) and (inputs(119));
    layer0_outputs(3693) <= '0';
    layer0_outputs(3694) <= inputs(182);
    layer0_outputs(3695) <= not((inputs(93)) or (inputs(24)));
    layer0_outputs(3696) <= (inputs(14)) and not (inputs(240));
    layer0_outputs(3697) <= inputs(23);
    layer0_outputs(3698) <= not(inputs(244));
    layer0_outputs(3699) <= '0';
    layer0_outputs(3700) <= inputs(189);
    layer0_outputs(3701) <= not(inputs(161)) or (inputs(134));
    layer0_outputs(3702) <= not(inputs(2));
    layer0_outputs(3703) <= '1';
    layer0_outputs(3704) <= (inputs(61)) and (inputs(192));
    layer0_outputs(3705) <= '1';
    layer0_outputs(3706) <= inputs(65);
    layer0_outputs(3707) <= '1';
    layer0_outputs(3708) <= '1';
    layer0_outputs(3709) <= inputs(27);
    layer0_outputs(3710) <= not(inputs(81)) or (inputs(129));
    layer0_outputs(3711) <= not(inputs(129));
    layer0_outputs(3712) <= not((inputs(245)) and (inputs(81)));
    layer0_outputs(3713) <= (inputs(204)) and not (inputs(134));
    layer0_outputs(3714) <= inputs(25);
    layer0_outputs(3715) <= (inputs(141)) and not (inputs(169));
    layer0_outputs(3716) <= not(inputs(57)) or (inputs(30));
    layer0_outputs(3717) <= not(inputs(187)) or (inputs(39));
    layer0_outputs(3718) <= '0';
    layer0_outputs(3719) <= inputs(49);
    layer0_outputs(3720) <= '0';
    layer0_outputs(3721) <= (inputs(66)) or (inputs(254));
    layer0_outputs(3722) <= '1';
    layer0_outputs(3723) <= '0';
    layer0_outputs(3724) <= '0';
    layer0_outputs(3725) <= (inputs(78)) and not (inputs(244));
    layer0_outputs(3726) <= (inputs(17)) and (inputs(250));
    layer0_outputs(3727) <= (inputs(28)) and (inputs(235));
    layer0_outputs(3728) <= not(inputs(5)) or (inputs(109));
    layer0_outputs(3729) <= inputs(215);
    layer0_outputs(3730) <= not((inputs(77)) or (inputs(151)));
    layer0_outputs(3731) <= '0';
    layer0_outputs(3732) <= not((inputs(138)) and (inputs(35)));
    layer0_outputs(3733) <= inputs(19);
    layer0_outputs(3734) <= inputs(80);
    layer0_outputs(3735) <= '1';
    layer0_outputs(3736) <= '0';
    layer0_outputs(3737) <= inputs(229);
    layer0_outputs(3738) <= not((inputs(103)) or (inputs(161)));
    layer0_outputs(3739) <= not(inputs(222)) or (inputs(52));
    layer0_outputs(3740) <= not(inputs(149));
    layer0_outputs(3741) <= '1';
    layer0_outputs(3742) <= not(inputs(115));
    layer0_outputs(3743) <= '0';
    layer0_outputs(3744) <= inputs(161);
    layer0_outputs(3745) <= '1';
    layer0_outputs(3746) <= '0';
    layer0_outputs(3747) <= not(inputs(151)) or (inputs(94));
    layer0_outputs(3748) <= not((inputs(35)) and (inputs(199)));
    layer0_outputs(3749) <= (inputs(173)) or (inputs(240));
    layer0_outputs(3750) <= '1';
    layer0_outputs(3751) <= not(inputs(236)) or (inputs(112));
    layer0_outputs(3752) <= '0';
    layer0_outputs(3753) <= '0';
    layer0_outputs(3754) <= (inputs(37)) and (inputs(123));
    layer0_outputs(3755) <= not((inputs(210)) xor (inputs(242)));
    layer0_outputs(3756) <= not(inputs(47)) or (inputs(117));
    layer0_outputs(3757) <= (inputs(124)) and not (inputs(76));
    layer0_outputs(3758) <= (inputs(75)) and (inputs(46));
    layer0_outputs(3759) <= '0';
    layer0_outputs(3760) <= not(inputs(108)) or (inputs(67));
    layer0_outputs(3761) <= not((inputs(52)) and (inputs(188)));
    layer0_outputs(3762) <= (inputs(122)) or (inputs(129));
    layer0_outputs(3763) <= not(inputs(203));
    layer0_outputs(3764) <= not((inputs(113)) or (inputs(170)));
    layer0_outputs(3765) <= '0';
    layer0_outputs(3766) <= '1';
    layer0_outputs(3767) <= not(inputs(222));
    layer0_outputs(3768) <= '0';
    layer0_outputs(3769) <= not(inputs(59)) or (inputs(224));
    layer0_outputs(3770) <= not(inputs(15));
    layer0_outputs(3771) <= (inputs(32)) and not (inputs(189));
    layer0_outputs(3772) <= (inputs(173)) and not (inputs(14));
    layer0_outputs(3773) <= inputs(61);
    layer0_outputs(3774) <= not((inputs(123)) or (inputs(33)));
    layer0_outputs(3775) <= (inputs(114)) and not (inputs(156));
    layer0_outputs(3776) <= (inputs(104)) and not (inputs(170));
    layer0_outputs(3777) <= not(inputs(67)) or (inputs(224));
    layer0_outputs(3778) <= '1';
    layer0_outputs(3779) <= '1';
    layer0_outputs(3780) <= not((inputs(15)) and (inputs(49)));
    layer0_outputs(3781) <= not(inputs(164)) or (inputs(43));
    layer0_outputs(3782) <= not(inputs(27));
    layer0_outputs(3783) <= not(inputs(72)) or (inputs(123));
    layer0_outputs(3784) <= not(inputs(87)) or (inputs(172));
    layer0_outputs(3785) <= not((inputs(161)) xor (inputs(133)));
    layer0_outputs(3786) <= (inputs(83)) or (inputs(142));
    layer0_outputs(3787) <= inputs(98);
    layer0_outputs(3788) <= (inputs(66)) and (inputs(66));
    layer0_outputs(3789) <= '0';
    layer0_outputs(3790) <= not((inputs(153)) or (inputs(227)));
    layer0_outputs(3791) <= not(inputs(216));
    layer0_outputs(3792) <= '0';
    layer0_outputs(3793) <= inputs(76);
    layer0_outputs(3794) <= '0';
    layer0_outputs(3795) <= not(inputs(223)) or (inputs(55));
    layer0_outputs(3796) <= '0';
    layer0_outputs(3797) <= (inputs(68)) and not (inputs(153));
    layer0_outputs(3798) <= not(inputs(178)) or (inputs(28));
    layer0_outputs(3799) <= not(inputs(71));
    layer0_outputs(3800) <= not((inputs(130)) xor (inputs(1)));
    layer0_outputs(3801) <= (inputs(116)) xor (inputs(81));
    layer0_outputs(3802) <= inputs(83);
    layer0_outputs(3803) <= (inputs(79)) and not (inputs(110));
    layer0_outputs(3804) <= not(inputs(134));
    layer0_outputs(3805) <= not((inputs(126)) and (inputs(138)));
    layer0_outputs(3806) <= '0';
    layer0_outputs(3807) <= '0';
    layer0_outputs(3808) <= not((inputs(41)) and (inputs(145)));
    layer0_outputs(3809) <= inputs(162);
    layer0_outputs(3810) <= inputs(76);
    layer0_outputs(3811) <= '0';
    layer0_outputs(3812) <= not(inputs(198));
    layer0_outputs(3813) <= (inputs(198)) and not (inputs(154));
    layer0_outputs(3814) <= (inputs(120)) or (inputs(153));
    layer0_outputs(3815) <= inputs(132);
    layer0_outputs(3816) <= '1';
    layer0_outputs(3817) <= (inputs(253)) and not (inputs(4));
    layer0_outputs(3818) <= '0';
    layer0_outputs(3819) <= '1';
    layer0_outputs(3820) <= '0';
    layer0_outputs(3821) <= not((inputs(211)) or (inputs(193)));
    layer0_outputs(3822) <= inputs(113);
    layer0_outputs(3823) <= (inputs(239)) and (inputs(6));
    layer0_outputs(3824) <= inputs(228);
    layer0_outputs(3825) <= not(inputs(1)) or (inputs(82));
    layer0_outputs(3826) <= (inputs(155)) and not (inputs(184));
    layer0_outputs(3827) <= inputs(81);
    layer0_outputs(3828) <= '1';
    layer0_outputs(3829) <= '1';
    layer0_outputs(3830) <= '1';
    layer0_outputs(3831) <= not(inputs(206));
    layer0_outputs(3832) <= '1';
    layer0_outputs(3833) <= '0';
    layer0_outputs(3834) <= not(inputs(104)) or (inputs(0));
    layer0_outputs(3835) <= (inputs(129)) or (inputs(63));
    layer0_outputs(3836) <= '1';
    layer0_outputs(3837) <= '0';
    layer0_outputs(3838) <= (inputs(194)) or (inputs(103));
    layer0_outputs(3839) <= (inputs(83)) or (inputs(113));
    layer0_outputs(3840) <= '0';
    layer0_outputs(3841) <= inputs(148);
    layer0_outputs(3842) <= inputs(89);
    layer0_outputs(3843) <= not((inputs(231)) and (inputs(217)));
    layer0_outputs(3844) <= not((inputs(64)) xor (inputs(2)));
    layer0_outputs(3845) <= inputs(18);
    layer0_outputs(3846) <= not((inputs(217)) and (inputs(90)));
    layer0_outputs(3847) <= not(inputs(13));
    layer0_outputs(3848) <= not(inputs(208));
    layer0_outputs(3849) <= not((inputs(184)) and (inputs(43)));
    layer0_outputs(3850) <= not(inputs(29)) or (inputs(22));
    layer0_outputs(3851) <= not(inputs(140)) or (inputs(246));
    layer0_outputs(3852) <= '1';
    layer0_outputs(3853) <= not((inputs(205)) and (inputs(54)));
    layer0_outputs(3854) <= not(inputs(32));
    layer0_outputs(3855) <= '1';
    layer0_outputs(3856) <= '0';
    layer0_outputs(3857) <= (inputs(166)) and not (inputs(132));
    layer0_outputs(3858) <= (inputs(22)) and not (inputs(231));
    layer0_outputs(3859) <= not(inputs(75)) or (inputs(61));
    layer0_outputs(3860) <= '1';
    layer0_outputs(3861) <= not((inputs(201)) and (inputs(220)));
    layer0_outputs(3862) <= not((inputs(148)) or (inputs(181)));
    layer0_outputs(3863) <= not(inputs(105)) or (inputs(170));
    layer0_outputs(3864) <= not((inputs(197)) and (inputs(187)));
    layer0_outputs(3865) <= (inputs(146)) xor (inputs(255));
    layer0_outputs(3866) <= '1';
    layer0_outputs(3867) <= not((inputs(224)) and (inputs(218)));
    layer0_outputs(3868) <= not(inputs(79)) or (inputs(217));
    layer0_outputs(3869) <= (inputs(145)) and (inputs(54));
    layer0_outputs(3870) <= (inputs(135)) and not (inputs(233));
    layer0_outputs(3871) <= not(inputs(139)) or (inputs(53));
    layer0_outputs(3872) <= not(inputs(250)) or (inputs(29));
    layer0_outputs(3873) <= '0';
    layer0_outputs(3874) <= '0';
    layer0_outputs(3875) <= inputs(129);
    layer0_outputs(3876) <= '1';
    layer0_outputs(3877) <= (inputs(39)) or (inputs(32));
    layer0_outputs(3878) <= not(inputs(49));
    layer0_outputs(3879) <= not((inputs(27)) and (inputs(55)));
    layer0_outputs(3880) <= not(inputs(142));
    layer0_outputs(3881) <= not((inputs(136)) xor (inputs(105)));
    layer0_outputs(3882) <= not(inputs(4)) or (inputs(94));
    layer0_outputs(3883) <= not(inputs(189)) or (inputs(167));
    layer0_outputs(3884) <= inputs(193);
    layer0_outputs(3885) <= '0';
    layer0_outputs(3886) <= not((inputs(35)) or (inputs(76)));
    layer0_outputs(3887) <= '1';
    layer0_outputs(3888) <= not((inputs(105)) or (inputs(51)));
    layer0_outputs(3889) <= (inputs(87)) and not (inputs(41));
    layer0_outputs(3890) <= '1';
    layer0_outputs(3891) <= '1';
    layer0_outputs(3892) <= '0';
    layer0_outputs(3893) <= inputs(254);
    layer0_outputs(3894) <= (inputs(157)) or (inputs(73));
    layer0_outputs(3895) <= not(inputs(188)) or (inputs(117));
    layer0_outputs(3896) <= (inputs(131)) or (inputs(130));
    layer0_outputs(3897) <= '1';
    layer0_outputs(3898) <= (inputs(8)) and (inputs(187));
    layer0_outputs(3899) <= inputs(93);
    layer0_outputs(3900) <= (inputs(108)) and (inputs(66));
    layer0_outputs(3901) <= not(inputs(100));
    layer0_outputs(3902) <= '1';
    layer0_outputs(3903) <= not(inputs(53));
    layer0_outputs(3904) <= not((inputs(52)) or (inputs(30)));
    layer0_outputs(3905) <= '1';
    layer0_outputs(3906) <= not(inputs(230));
    layer0_outputs(3907) <= not((inputs(209)) xor (inputs(74)));
    layer0_outputs(3908) <= not(inputs(193)) or (inputs(86));
    layer0_outputs(3909) <= not(inputs(17));
    layer0_outputs(3910) <= inputs(232);
    layer0_outputs(3911) <= not((inputs(168)) and (inputs(147)));
    layer0_outputs(3912) <= (inputs(111)) and (inputs(233));
    layer0_outputs(3913) <= not(inputs(178)) or (inputs(101));
    layer0_outputs(3914) <= (inputs(216)) and not (inputs(49));
    layer0_outputs(3915) <= '1';
    layer0_outputs(3916) <= '1';
    layer0_outputs(3917) <= '1';
    layer0_outputs(3918) <= '0';
    layer0_outputs(3919) <= not(inputs(74));
    layer0_outputs(3920) <= not(inputs(66)) or (inputs(151));
    layer0_outputs(3921) <= (inputs(130)) or (inputs(88));
    layer0_outputs(3922) <= (inputs(120)) and (inputs(114));
    layer0_outputs(3923) <= not(inputs(84));
    layer0_outputs(3924) <= '1';
    layer0_outputs(3925) <= inputs(157);
    layer0_outputs(3926) <= not((inputs(158)) xor (inputs(31)));
    layer0_outputs(3927) <= not((inputs(144)) or (inputs(179)));
    layer0_outputs(3928) <= (inputs(64)) and (inputs(83));
    layer0_outputs(3929) <= not(inputs(146)) or (inputs(148));
    layer0_outputs(3930) <= '1';
    layer0_outputs(3931) <= inputs(71);
    layer0_outputs(3932) <= '0';
    layer0_outputs(3933) <= '1';
    layer0_outputs(3934) <= '1';
    layer0_outputs(3935) <= (inputs(17)) and not (inputs(185));
    layer0_outputs(3936) <= not((inputs(88)) and (inputs(56)));
    layer0_outputs(3937) <= (inputs(85)) and not (inputs(129));
    layer0_outputs(3938) <= (inputs(17)) and not (inputs(235));
    layer0_outputs(3939) <= (inputs(116)) and (inputs(70));
    layer0_outputs(3940) <= '1';
    layer0_outputs(3941) <= (inputs(193)) and not (inputs(158));
    layer0_outputs(3942) <= not(inputs(247));
    layer0_outputs(3943) <= '1';
    layer0_outputs(3944) <= inputs(144);
    layer0_outputs(3945) <= '0';
    layer0_outputs(3946) <= not(inputs(121));
    layer0_outputs(3947) <= not(inputs(128));
    layer0_outputs(3948) <= not(inputs(172));
    layer0_outputs(3949) <= '0';
    layer0_outputs(3950) <= (inputs(117)) and not (inputs(54));
    layer0_outputs(3951) <= (inputs(99)) and not (inputs(76));
    layer0_outputs(3952) <= (inputs(91)) xor (inputs(63));
    layer0_outputs(3953) <= not(inputs(115)) or (inputs(100));
    layer0_outputs(3954) <= not((inputs(156)) and (inputs(33)));
    layer0_outputs(3955) <= (inputs(154)) and (inputs(235));
    layer0_outputs(3956) <= not((inputs(171)) or (inputs(158)));
    layer0_outputs(3957) <= '1';
    layer0_outputs(3958) <= (inputs(153)) and not (inputs(119));
    layer0_outputs(3959) <= inputs(174);
    layer0_outputs(3960) <= not(inputs(9)) or (inputs(146));
    layer0_outputs(3961) <= not(inputs(216));
    layer0_outputs(3962) <= (inputs(132)) and (inputs(81));
    layer0_outputs(3963) <= (inputs(213)) and not (inputs(223));
    layer0_outputs(3964) <= (inputs(123)) or (inputs(127));
    layer0_outputs(3965) <= (inputs(200)) or (inputs(152));
    layer0_outputs(3966) <= (inputs(187)) and (inputs(133));
    layer0_outputs(3967) <= not((inputs(121)) and (inputs(108)));
    layer0_outputs(3968) <= (inputs(98)) or (inputs(183));
    layer0_outputs(3969) <= not((inputs(95)) or (inputs(212)));
    layer0_outputs(3970) <= (inputs(44)) and not (inputs(141));
    layer0_outputs(3971) <= not(inputs(179));
    layer0_outputs(3972) <= '0';
    layer0_outputs(3973) <= inputs(165);
    layer0_outputs(3974) <= inputs(152);
    layer0_outputs(3975) <= not(inputs(228));
    layer0_outputs(3976) <= '1';
    layer0_outputs(3977) <= '0';
    layer0_outputs(3978) <= (inputs(127)) and not (inputs(247));
    layer0_outputs(3979) <= not((inputs(8)) and (inputs(236)));
    layer0_outputs(3980) <= '1';
    layer0_outputs(3981) <= (inputs(201)) and not (inputs(124));
    layer0_outputs(3982) <= not(inputs(27));
    layer0_outputs(3983) <= not(inputs(110));
    layer0_outputs(3984) <= '1';
    layer0_outputs(3985) <= '0';
    layer0_outputs(3986) <= '0';
    layer0_outputs(3987) <= not(inputs(42)) or (inputs(206));
    layer0_outputs(3988) <= not((inputs(73)) or (inputs(218)));
    layer0_outputs(3989) <= '1';
    layer0_outputs(3990) <= '1';
    layer0_outputs(3991) <= inputs(9);
    layer0_outputs(3992) <= not(inputs(95)) or (inputs(166));
    layer0_outputs(3993) <= '1';
    layer0_outputs(3994) <= '1';
    layer0_outputs(3995) <= inputs(130);
    layer0_outputs(3996) <= (inputs(67)) xor (inputs(160));
    layer0_outputs(3997) <= not(inputs(77));
    layer0_outputs(3998) <= (inputs(89)) and not (inputs(77));
    layer0_outputs(3999) <= (inputs(53)) and (inputs(63));
    layer0_outputs(4000) <= not((inputs(192)) or (inputs(204)));
    layer0_outputs(4001) <= not((inputs(219)) and (inputs(245)));
    layer0_outputs(4002) <= '1';
    layer0_outputs(4003) <= not((inputs(70)) and (inputs(95)));
    layer0_outputs(4004) <= '0';
    layer0_outputs(4005) <= (inputs(228)) or (inputs(131));
    layer0_outputs(4006) <= (inputs(36)) or (inputs(243));
    layer0_outputs(4007) <= '1';
    layer0_outputs(4008) <= (inputs(122)) and not (inputs(14));
    layer0_outputs(4009) <= not((inputs(86)) xor (inputs(42)));
    layer0_outputs(4010) <= (inputs(110)) and not (inputs(120));
    layer0_outputs(4011) <= (inputs(234)) and not (inputs(219));
    layer0_outputs(4012) <= not(inputs(167)) or (inputs(165));
    layer0_outputs(4013) <= '1';
    layer0_outputs(4014) <= inputs(3);
    layer0_outputs(4015) <= (inputs(82)) and (inputs(223));
    layer0_outputs(4016) <= not((inputs(127)) and (inputs(46)));
    layer0_outputs(4017) <= not((inputs(47)) xor (inputs(151)));
    layer0_outputs(4018) <= '0';
    layer0_outputs(4019) <= inputs(34);
    layer0_outputs(4020) <= (inputs(143)) and not (inputs(120));
    layer0_outputs(4021) <= '0';
    layer0_outputs(4022) <= (inputs(92)) and not (inputs(224));
    layer0_outputs(4023) <= (inputs(128)) and (inputs(233));
    layer0_outputs(4024) <= not(inputs(54)) or (inputs(74));
    layer0_outputs(4025) <= '1';
    layer0_outputs(4026) <= '1';
    layer0_outputs(4027) <= not((inputs(23)) or (inputs(66)));
    layer0_outputs(4028) <= '0';
    layer0_outputs(4029) <= not(inputs(48)) or (inputs(135));
    layer0_outputs(4030) <= '1';
    layer0_outputs(4031) <= not((inputs(136)) or (inputs(148)));
    layer0_outputs(4032) <= (inputs(204)) or (inputs(227));
    layer0_outputs(4033) <= (inputs(221)) or (inputs(205));
    layer0_outputs(4034) <= (inputs(206)) and not (inputs(15));
    layer0_outputs(4035) <= not(inputs(23)) or (inputs(158));
    layer0_outputs(4036) <= not(inputs(102));
    layer0_outputs(4037) <= (inputs(46)) and not (inputs(95));
    layer0_outputs(4038) <= not((inputs(241)) xor (inputs(224)));
    layer0_outputs(4039) <= (inputs(42)) and (inputs(45));
    layer0_outputs(4040) <= not((inputs(227)) and (inputs(172)));
    layer0_outputs(4041) <= not((inputs(86)) and (inputs(32)));
    layer0_outputs(4042) <= (inputs(172)) or (inputs(188));
    layer0_outputs(4043) <= not(inputs(176));
    layer0_outputs(4044) <= not(inputs(122));
    layer0_outputs(4045) <= (inputs(56)) and (inputs(249));
    layer0_outputs(4046) <= inputs(1);
    layer0_outputs(4047) <= '1';
    layer0_outputs(4048) <= not((inputs(20)) or (inputs(44)));
    layer0_outputs(4049) <= '0';
    layer0_outputs(4050) <= (inputs(134)) xor (inputs(105));
    layer0_outputs(4051) <= not((inputs(214)) or (inputs(25)));
    layer0_outputs(4052) <= not(inputs(10)) or (inputs(159));
    layer0_outputs(4053) <= (inputs(38)) and not (inputs(23));
    layer0_outputs(4054) <= not((inputs(73)) and (inputs(104)));
    layer0_outputs(4055) <= inputs(60);
    layer0_outputs(4056) <= '1';
    layer0_outputs(4057) <= (inputs(181)) and (inputs(251));
    layer0_outputs(4058) <= not(inputs(215));
    layer0_outputs(4059) <= inputs(84);
    layer0_outputs(4060) <= not((inputs(16)) xor (inputs(109)));
    layer0_outputs(4061) <= (inputs(163)) or (inputs(197));
    layer0_outputs(4062) <= '1';
    layer0_outputs(4063) <= (inputs(187)) and not (inputs(100));
    layer0_outputs(4064) <= '1';
    layer0_outputs(4065) <= '0';
    layer0_outputs(4066) <= '0';
    layer0_outputs(4067) <= not(inputs(237)) or (inputs(30));
    layer0_outputs(4068) <= inputs(252);
    layer0_outputs(4069) <= '1';
    layer0_outputs(4070) <= (inputs(188)) or (inputs(236));
    layer0_outputs(4071) <= not((inputs(242)) and (inputs(68)));
    layer0_outputs(4072) <= not(inputs(151));
    layer0_outputs(4073) <= not(inputs(6)) or (inputs(83));
    layer0_outputs(4074) <= inputs(66);
    layer0_outputs(4075) <= not(inputs(32)) or (inputs(38));
    layer0_outputs(4076) <= '1';
    layer0_outputs(4077) <= not(inputs(62));
    layer0_outputs(4078) <= not(inputs(94));
    layer0_outputs(4079) <= (inputs(63)) and not (inputs(110));
    layer0_outputs(4080) <= inputs(185);
    layer0_outputs(4081) <= not((inputs(182)) and (inputs(174)));
    layer0_outputs(4082) <= not(inputs(142));
    layer0_outputs(4083) <= not(inputs(233));
    layer0_outputs(4084) <= inputs(107);
    layer0_outputs(4085) <= '0';
    layer0_outputs(4086) <= inputs(212);
    layer0_outputs(4087) <= not((inputs(208)) or (inputs(82)));
    layer0_outputs(4088) <= not(inputs(239)) or (inputs(50));
    layer0_outputs(4089) <= inputs(100);
    layer0_outputs(4090) <= '1';
    layer0_outputs(4091) <= '1';
    layer0_outputs(4092) <= not(inputs(59));
    layer0_outputs(4093) <= '0';
    layer0_outputs(4094) <= not(inputs(110));
    layer0_outputs(4095) <= (inputs(232)) and not (inputs(224));
    layer0_outputs(4096) <= '1';
    layer0_outputs(4097) <= not(inputs(87));
    layer0_outputs(4098) <= (inputs(45)) and (inputs(34));
    layer0_outputs(4099) <= not(inputs(191)) or (inputs(21));
    layer0_outputs(4100) <= (inputs(56)) and not (inputs(111));
    layer0_outputs(4101) <= not((inputs(229)) and (inputs(150)));
    layer0_outputs(4102) <= not((inputs(19)) or (inputs(224)));
    layer0_outputs(4103) <= '0';
    layer0_outputs(4104) <= (inputs(139)) or (inputs(191));
    layer0_outputs(4105) <= '0';
    layer0_outputs(4106) <= inputs(254);
    layer0_outputs(4107) <= not(inputs(95));
    layer0_outputs(4108) <= not((inputs(243)) and (inputs(128)));
    layer0_outputs(4109) <= (inputs(108)) and (inputs(59));
    layer0_outputs(4110) <= inputs(253);
    layer0_outputs(4111) <= '1';
    layer0_outputs(4112) <= '1';
    layer0_outputs(4113) <= '0';
    layer0_outputs(4114) <= not(inputs(236));
    layer0_outputs(4115) <= not((inputs(32)) and (inputs(122)));
    layer0_outputs(4116) <= not((inputs(106)) xor (inputs(124)));
    layer0_outputs(4117) <= not((inputs(254)) or (inputs(176)));
    layer0_outputs(4118) <= '1';
    layer0_outputs(4119) <= not((inputs(183)) and (inputs(212)));
    layer0_outputs(4120) <= '1';
    layer0_outputs(4121) <= (inputs(127)) or (inputs(207));
    layer0_outputs(4122) <= '0';
    layer0_outputs(4123) <= inputs(255);
    layer0_outputs(4124) <= '0';
    layer0_outputs(4125) <= not(inputs(230)) or (inputs(72));
    layer0_outputs(4126) <= not(inputs(189));
    layer0_outputs(4127) <= not(inputs(202));
    layer0_outputs(4128) <= not(inputs(114));
    layer0_outputs(4129) <= inputs(207);
    layer0_outputs(4130) <= '1';
    layer0_outputs(4131) <= inputs(6);
    layer0_outputs(4132) <= '1';
    layer0_outputs(4133) <= '1';
    layer0_outputs(4134) <= not((inputs(72)) and (inputs(199)));
    layer0_outputs(4135) <= not(inputs(112));
    layer0_outputs(4136) <= not((inputs(97)) and (inputs(233)));
    layer0_outputs(4137) <= inputs(70);
    layer0_outputs(4138) <= not(inputs(103));
    layer0_outputs(4139) <= not((inputs(230)) and (inputs(170)));
    layer0_outputs(4140) <= not(inputs(21)) or (inputs(142));
    layer0_outputs(4141) <= not(inputs(220));
    layer0_outputs(4142) <= (inputs(18)) or (inputs(211));
    layer0_outputs(4143) <= (inputs(145)) and not (inputs(11));
    layer0_outputs(4144) <= '1';
    layer0_outputs(4145) <= '0';
    layer0_outputs(4146) <= not(inputs(44));
    layer0_outputs(4147) <= not(inputs(98)) or (inputs(171));
    layer0_outputs(4148) <= '1';
    layer0_outputs(4149) <= (inputs(73)) and (inputs(51));
    layer0_outputs(4150) <= '1';
    layer0_outputs(4151) <= (inputs(177)) and not (inputs(148));
    layer0_outputs(4152) <= not(inputs(5));
    layer0_outputs(4153) <= '0';
    layer0_outputs(4154) <= not(inputs(213)) or (inputs(77));
    layer0_outputs(4155) <= not(inputs(179)) or (inputs(105));
    layer0_outputs(4156) <= not((inputs(205)) xor (inputs(214)));
    layer0_outputs(4157) <= not(inputs(89)) or (inputs(253));
    layer0_outputs(4158) <= not(inputs(69));
    layer0_outputs(4159) <= not(inputs(198));
    layer0_outputs(4160) <= '0';
    layer0_outputs(4161) <= not(inputs(56));
    layer0_outputs(4162) <= not(inputs(93));
    layer0_outputs(4163) <= inputs(223);
    layer0_outputs(4164) <= not(inputs(235));
    layer0_outputs(4165) <= '0';
    layer0_outputs(4166) <= '0';
    layer0_outputs(4167) <= (inputs(99)) and not (inputs(93));
    layer0_outputs(4168) <= (inputs(2)) and not (inputs(2));
    layer0_outputs(4169) <= not((inputs(189)) and (inputs(211)));
    layer0_outputs(4170) <= (inputs(236)) and (inputs(213));
    layer0_outputs(4171) <= '0';
    layer0_outputs(4172) <= not(inputs(6));
    layer0_outputs(4173) <= (inputs(197)) and (inputs(191));
    layer0_outputs(4174) <= '1';
    layer0_outputs(4175) <= '1';
    layer0_outputs(4176) <= (inputs(143)) and not (inputs(86));
    layer0_outputs(4177) <= '0';
    layer0_outputs(4178) <= (inputs(8)) or (inputs(240));
    layer0_outputs(4179) <= '1';
    layer0_outputs(4180) <= not(inputs(201));
    layer0_outputs(4181) <= (inputs(9)) and not (inputs(169));
    layer0_outputs(4182) <= not(inputs(207)) or (inputs(210));
    layer0_outputs(4183) <= inputs(95);
    layer0_outputs(4184) <= not(inputs(185)) or (inputs(97));
    layer0_outputs(4185) <= not(inputs(238));
    layer0_outputs(4186) <= not(inputs(159)) or (inputs(183));
    layer0_outputs(4187) <= inputs(244);
    layer0_outputs(4188) <= not(inputs(245)) or (inputs(73));
    layer0_outputs(4189) <= not(inputs(70)) or (inputs(15));
    layer0_outputs(4190) <= '0';
    layer0_outputs(4191) <= '1';
    layer0_outputs(4192) <= (inputs(235)) and (inputs(9));
    layer0_outputs(4193) <= (inputs(167)) or (inputs(225));
    layer0_outputs(4194) <= '1';
    layer0_outputs(4195) <= inputs(38);
    layer0_outputs(4196) <= '0';
    layer0_outputs(4197) <= not((inputs(250)) or (inputs(227)));
    layer0_outputs(4198) <= '0';
    layer0_outputs(4199) <= inputs(28);
    layer0_outputs(4200) <= '1';
    layer0_outputs(4201) <= (inputs(99)) and not (inputs(174));
    layer0_outputs(4202) <= (inputs(194)) and (inputs(5));
    layer0_outputs(4203) <= (inputs(62)) or (inputs(116));
    layer0_outputs(4204) <= inputs(67);
    layer0_outputs(4205) <= not(inputs(24)) or (inputs(110));
    layer0_outputs(4206) <= inputs(16);
    layer0_outputs(4207) <= '1';
    layer0_outputs(4208) <= inputs(114);
    layer0_outputs(4209) <= (inputs(185)) or (inputs(236));
    layer0_outputs(4210) <= (inputs(49)) and (inputs(90));
    layer0_outputs(4211) <= not(inputs(126));
    layer0_outputs(4212) <= '1';
    layer0_outputs(4213) <= inputs(21);
    layer0_outputs(4214) <= '1';
    layer0_outputs(4215) <= '0';
    layer0_outputs(4216) <= not((inputs(172)) and (inputs(153)));
    layer0_outputs(4217) <= inputs(236);
    layer0_outputs(4218) <= '0';
    layer0_outputs(4219) <= not(inputs(8));
    layer0_outputs(4220) <= (inputs(104)) and (inputs(245));
    layer0_outputs(4221) <= not(inputs(226));
    layer0_outputs(4222) <= (inputs(230)) and (inputs(182));
    layer0_outputs(4223) <= inputs(184);
    layer0_outputs(4224) <= not(inputs(150)) or (inputs(57));
    layer0_outputs(4225) <= not((inputs(109)) or (inputs(126)));
    layer0_outputs(4226) <= (inputs(109)) and (inputs(127));
    layer0_outputs(4227) <= not((inputs(177)) or (inputs(251)));
    layer0_outputs(4228) <= '1';
    layer0_outputs(4229) <= (inputs(60)) or (inputs(158));
    layer0_outputs(4230) <= '1';
    layer0_outputs(4231) <= '1';
    layer0_outputs(4232) <= '0';
    layer0_outputs(4233) <= not(inputs(35)) or (inputs(113));
    layer0_outputs(4234) <= '1';
    layer0_outputs(4235) <= '0';
    layer0_outputs(4236) <= inputs(4);
    layer0_outputs(4237) <= (inputs(44)) and (inputs(5));
    layer0_outputs(4238) <= (inputs(86)) or (inputs(206));
    layer0_outputs(4239) <= not(inputs(24)) or (inputs(212));
    layer0_outputs(4240) <= '0';
    layer0_outputs(4241) <= inputs(47);
    layer0_outputs(4242) <= '0';
    layer0_outputs(4243) <= '1';
    layer0_outputs(4244) <= not(inputs(188));
    layer0_outputs(4245) <= '0';
    layer0_outputs(4246) <= (inputs(230)) and (inputs(149));
    layer0_outputs(4247) <= not(inputs(96));
    layer0_outputs(4248) <= '0';
    layer0_outputs(4249) <= '1';
    layer0_outputs(4250) <= '1';
    layer0_outputs(4251) <= '1';
    layer0_outputs(4252) <= (inputs(40)) and not (inputs(211));
    layer0_outputs(4253) <= not(inputs(226)) or (inputs(70));
    layer0_outputs(4254) <= (inputs(21)) and not (inputs(217));
    layer0_outputs(4255) <= not(inputs(3));
    layer0_outputs(4256) <= (inputs(52)) and not (inputs(225));
    layer0_outputs(4257) <= '1';
    layer0_outputs(4258) <= not((inputs(144)) or (inputs(36)));
    layer0_outputs(4259) <= not(inputs(34)) or (inputs(82));
    layer0_outputs(4260) <= not((inputs(245)) or (inputs(148)));
    layer0_outputs(4261) <= not((inputs(230)) and (inputs(151)));
    layer0_outputs(4262) <= (inputs(167)) and not (inputs(133));
    layer0_outputs(4263) <= (inputs(16)) and not (inputs(108));
    layer0_outputs(4264) <= not(inputs(238)) or (inputs(139));
    layer0_outputs(4265) <= inputs(234);
    layer0_outputs(4266) <= not(inputs(2)) or (inputs(164));
    layer0_outputs(4267) <= '0';
    layer0_outputs(4268) <= (inputs(186)) and not (inputs(21));
    layer0_outputs(4269) <= '0';
    layer0_outputs(4270) <= (inputs(87)) and not (inputs(76));
    layer0_outputs(4271) <= not((inputs(252)) and (inputs(5)));
    layer0_outputs(4272) <= (inputs(164)) and not (inputs(73));
    layer0_outputs(4273) <= not(inputs(4));
    layer0_outputs(4274) <= (inputs(168)) and (inputs(68));
    layer0_outputs(4275) <= '1';
    layer0_outputs(4276) <= not((inputs(17)) xor (inputs(232)));
    layer0_outputs(4277) <= not(inputs(226));
    layer0_outputs(4278) <= '1';
    layer0_outputs(4279) <= inputs(176);
    layer0_outputs(4280) <= (inputs(100)) and not (inputs(211));
    layer0_outputs(4281) <= '0';
    layer0_outputs(4282) <= '0';
    layer0_outputs(4283) <= not((inputs(251)) or (inputs(169)));
    layer0_outputs(4284) <= (inputs(85)) and not (inputs(209));
    layer0_outputs(4285) <= not(inputs(170));
    layer0_outputs(4286) <= '0';
    layer0_outputs(4287) <= not((inputs(63)) or (inputs(137)));
    layer0_outputs(4288) <= '1';
    layer0_outputs(4289) <= inputs(133);
    layer0_outputs(4290) <= not(inputs(224));
    layer0_outputs(4291) <= not(inputs(1)) or (inputs(238));
    layer0_outputs(4292) <= inputs(252);
    layer0_outputs(4293) <= not(inputs(199)) or (inputs(48));
    layer0_outputs(4294) <= inputs(122);
    layer0_outputs(4295) <= (inputs(190)) xor (inputs(164));
    layer0_outputs(4296) <= not((inputs(38)) and (inputs(2)));
    layer0_outputs(4297) <= (inputs(194)) or (inputs(210));
    layer0_outputs(4298) <= (inputs(44)) xor (inputs(83));
    layer0_outputs(4299) <= not((inputs(28)) and (inputs(189)));
    layer0_outputs(4300) <= (inputs(50)) and (inputs(1));
    layer0_outputs(4301) <= inputs(70);
    layer0_outputs(4302) <= not((inputs(249)) or (inputs(80)));
    layer0_outputs(4303) <= '0';
    layer0_outputs(4304) <= not(inputs(117));
    layer0_outputs(4305) <= '1';
    layer0_outputs(4306) <= (inputs(135)) and not (inputs(203));
    layer0_outputs(4307) <= inputs(139);
    layer0_outputs(4308) <= '0';
    layer0_outputs(4309) <= inputs(42);
    layer0_outputs(4310) <= (inputs(150)) and not (inputs(87));
    layer0_outputs(4311) <= not((inputs(164)) or (inputs(229)));
    layer0_outputs(4312) <= (inputs(154)) and (inputs(220));
    layer0_outputs(4313) <= '1';
    layer0_outputs(4314) <= (inputs(116)) or (inputs(214));
    layer0_outputs(4315) <= '1';
    layer0_outputs(4316) <= not(inputs(245));
    layer0_outputs(4317) <= '0';
    layer0_outputs(4318) <= not(inputs(191)) or (inputs(100));
    layer0_outputs(4319) <= not(inputs(86)) or (inputs(192));
    layer0_outputs(4320) <= '1';
    layer0_outputs(4321) <= (inputs(46)) or (inputs(119));
    layer0_outputs(4322) <= '0';
    layer0_outputs(4323) <= not(inputs(206)) or (inputs(103));
    layer0_outputs(4324) <= inputs(18);
    layer0_outputs(4325) <= inputs(247);
    layer0_outputs(4326) <= (inputs(202)) or (inputs(110));
    layer0_outputs(4327) <= inputs(164);
    layer0_outputs(4328) <= '0';
    layer0_outputs(4329) <= (inputs(179)) or (inputs(226));
    layer0_outputs(4330) <= (inputs(59)) or (inputs(187));
    layer0_outputs(4331) <= not(inputs(115)) or (inputs(17));
    layer0_outputs(4332) <= (inputs(154)) and not (inputs(160));
    layer0_outputs(4333) <= not(inputs(205)) or (inputs(130));
    layer0_outputs(4334) <= not(inputs(108));
    layer0_outputs(4335) <= not((inputs(109)) or (inputs(146)));
    layer0_outputs(4336) <= '0';
    layer0_outputs(4337) <= not((inputs(151)) xor (inputs(144)));
    layer0_outputs(4338) <= '1';
    layer0_outputs(4339) <= inputs(216);
    layer0_outputs(4340) <= inputs(177);
    layer0_outputs(4341) <= not(inputs(207)) or (inputs(231));
    layer0_outputs(4342) <= not(inputs(211)) or (inputs(104));
    layer0_outputs(4343) <= not(inputs(9)) or (inputs(246));
    layer0_outputs(4344) <= '0';
    layer0_outputs(4345) <= not((inputs(58)) and (inputs(238)));
    layer0_outputs(4346) <= inputs(233);
    layer0_outputs(4347) <= (inputs(255)) and not (inputs(22));
    layer0_outputs(4348) <= (inputs(3)) and (inputs(143));
    layer0_outputs(4349) <= inputs(64);
    layer0_outputs(4350) <= '1';
    layer0_outputs(4351) <= (inputs(27)) and not (inputs(236));
    layer0_outputs(4352) <= not(inputs(36)) or (inputs(222));
    layer0_outputs(4353) <= (inputs(94)) and (inputs(240));
    layer0_outputs(4354) <= '1';
    layer0_outputs(4355) <= not((inputs(155)) or (inputs(250)));
    layer0_outputs(4356) <= '0';
    layer0_outputs(4357) <= not((inputs(120)) or (inputs(104)));
    layer0_outputs(4358) <= (inputs(175)) and (inputs(63));
    layer0_outputs(4359) <= inputs(160);
    layer0_outputs(4360) <= '0';
    layer0_outputs(4361) <= (inputs(228)) or (inputs(190));
    layer0_outputs(4362) <= not(inputs(175));
    layer0_outputs(4363) <= '0';
    layer0_outputs(4364) <= '0';
    layer0_outputs(4365) <= '0';
    layer0_outputs(4366) <= '1';
    layer0_outputs(4367) <= not(inputs(47));
    layer0_outputs(4368) <= (inputs(80)) and not (inputs(178));
    layer0_outputs(4369) <= not(inputs(131)) or (inputs(26));
    layer0_outputs(4370) <= '0';
    layer0_outputs(4371) <= inputs(192);
    layer0_outputs(4372) <= not(inputs(184));
    layer0_outputs(4373) <= '1';
    layer0_outputs(4374) <= not((inputs(234)) or (inputs(27)));
    layer0_outputs(4375) <= (inputs(140)) or (inputs(34));
    layer0_outputs(4376) <= '1';
    layer0_outputs(4377) <= not(inputs(126)) or (inputs(15));
    layer0_outputs(4378) <= not((inputs(86)) and (inputs(34)));
    layer0_outputs(4379) <= '0';
    layer0_outputs(4380) <= inputs(223);
    layer0_outputs(4381) <= inputs(18);
    layer0_outputs(4382) <= '0';
    layer0_outputs(4383) <= '1';
    layer0_outputs(4384) <= inputs(144);
    layer0_outputs(4385) <= (inputs(7)) and not (inputs(55));
    layer0_outputs(4386) <= '0';
    layer0_outputs(4387) <= not(inputs(100));
    layer0_outputs(4388) <= not(inputs(62)) or (inputs(251));
    layer0_outputs(4389) <= (inputs(229)) and (inputs(228));
    layer0_outputs(4390) <= (inputs(187)) and (inputs(153));
    layer0_outputs(4391) <= (inputs(135)) and not (inputs(235));
    layer0_outputs(4392) <= '1';
    layer0_outputs(4393) <= '1';
    layer0_outputs(4394) <= not((inputs(126)) xor (inputs(84)));
    layer0_outputs(4395) <= '1';
    layer0_outputs(4396) <= '1';
    layer0_outputs(4397) <= not((inputs(120)) and (inputs(204)));
    layer0_outputs(4398) <= '0';
    layer0_outputs(4399) <= (inputs(117)) and not (inputs(19));
    layer0_outputs(4400) <= '1';
    layer0_outputs(4401) <= not(inputs(181)) or (inputs(7));
    layer0_outputs(4402) <= inputs(25);
    layer0_outputs(4403) <= '1';
    layer0_outputs(4404) <= not(inputs(4)) or (inputs(49));
    layer0_outputs(4405) <= (inputs(160)) or (inputs(229));
    layer0_outputs(4406) <= not(inputs(241)) or (inputs(199));
    layer0_outputs(4407) <= inputs(177);
    layer0_outputs(4408) <= '0';
    layer0_outputs(4409) <= '1';
    layer0_outputs(4410) <= (inputs(24)) and not (inputs(6));
    layer0_outputs(4411) <= (inputs(135)) and not (inputs(105));
    layer0_outputs(4412) <= (inputs(193)) or (inputs(108));
    layer0_outputs(4413) <= inputs(21);
    layer0_outputs(4414) <= (inputs(94)) and not (inputs(137));
    layer0_outputs(4415) <= not(inputs(9));
    layer0_outputs(4416) <= '0';
    layer0_outputs(4417) <= '0';
    layer0_outputs(4418) <= '1';
    layer0_outputs(4419) <= '1';
    layer0_outputs(4420) <= '1';
    layer0_outputs(4421) <= '1';
    layer0_outputs(4422) <= not(inputs(228)) or (inputs(134));
    layer0_outputs(4423) <= inputs(121);
    layer0_outputs(4424) <= '0';
    layer0_outputs(4425) <= not((inputs(69)) and (inputs(49)));
    layer0_outputs(4426) <= inputs(203);
    layer0_outputs(4427) <= not(inputs(34)) or (inputs(41));
    layer0_outputs(4428) <= not((inputs(212)) and (inputs(92)));
    layer0_outputs(4429) <= not(inputs(152)) or (inputs(54));
    layer0_outputs(4430) <= not(inputs(134)) or (inputs(235));
    layer0_outputs(4431) <= '1';
    layer0_outputs(4432) <= (inputs(19)) and not (inputs(208));
    layer0_outputs(4433) <= (inputs(3)) and not (inputs(237));
    layer0_outputs(4434) <= '1';
    layer0_outputs(4435) <= not((inputs(126)) and (inputs(206)));
    layer0_outputs(4436) <= not(inputs(42)) or (inputs(74));
    layer0_outputs(4437) <= (inputs(237)) and (inputs(27));
    layer0_outputs(4438) <= '1';
    layer0_outputs(4439) <= '0';
    layer0_outputs(4440) <= not((inputs(96)) and (inputs(211)));
    layer0_outputs(4441) <= inputs(211);
    layer0_outputs(4442) <= not((inputs(132)) or (inputs(251)));
    layer0_outputs(4443) <= inputs(180);
    layer0_outputs(4444) <= '0';
    layer0_outputs(4445) <= inputs(11);
    layer0_outputs(4446) <= not(inputs(247));
    layer0_outputs(4447) <= (inputs(52)) and not (inputs(89));
    layer0_outputs(4448) <= not(inputs(157)) or (inputs(185));
    layer0_outputs(4449) <= (inputs(204)) or (inputs(155));
    layer0_outputs(4450) <= not(inputs(75));
    layer0_outputs(4451) <= (inputs(91)) xor (inputs(95));
    layer0_outputs(4452) <= not(inputs(140)) or (inputs(116));
    layer0_outputs(4453) <= not(inputs(46));
    layer0_outputs(4454) <= not(inputs(97));
    layer0_outputs(4455) <= not(inputs(207)) or (inputs(147));
    layer0_outputs(4456) <= inputs(197);
    layer0_outputs(4457) <= (inputs(210)) xor (inputs(219));
    layer0_outputs(4458) <= not(inputs(78));
    layer0_outputs(4459) <= inputs(155);
    layer0_outputs(4460) <= not(inputs(14));
    layer0_outputs(4461) <= (inputs(59)) or (inputs(11));
    layer0_outputs(4462) <= not(inputs(154));
    layer0_outputs(4463) <= (inputs(145)) or (inputs(239));
    layer0_outputs(4464) <= (inputs(76)) and not (inputs(54));
    layer0_outputs(4465) <= '0';
    layer0_outputs(4466) <= (inputs(222)) and not (inputs(144));
    layer0_outputs(4467) <= '1';
    layer0_outputs(4468) <= '0';
    layer0_outputs(4469) <= '0';
    layer0_outputs(4470) <= '1';
    layer0_outputs(4471) <= inputs(162);
    layer0_outputs(4472) <= (inputs(60)) and (inputs(80));
    layer0_outputs(4473) <= inputs(80);
    layer0_outputs(4474) <= not((inputs(113)) or (inputs(12)));
    layer0_outputs(4475) <= not(inputs(58)) or (inputs(94));
    layer0_outputs(4476) <= (inputs(4)) and not (inputs(158));
    layer0_outputs(4477) <= (inputs(230)) and not (inputs(215));
    layer0_outputs(4478) <= not(inputs(28)) or (inputs(68));
    layer0_outputs(4479) <= (inputs(143)) and not (inputs(232));
    layer0_outputs(4480) <= not(inputs(102));
    layer0_outputs(4481) <= '0';
    layer0_outputs(4482) <= not(inputs(96)) or (inputs(130));
    layer0_outputs(4483) <= '0';
    layer0_outputs(4484) <= (inputs(126)) or (inputs(228));
    layer0_outputs(4485) <= not(inputs(135));
    layer0_outputs(4486) <= not(inputs(102)) or (inputs(205));
    layer0_outputs(4487) <= not(inputs(81));
    layer0_outputs(4488) <= '0';
    layer0_outputs(4489) <= not(inputs(193));
    layer0_outputs(4490) <= (inputs(3)) and (inputs(125));
    layer0_outputs(4491) <= '0';
    layer0_outputs(4492) <= not(inputs(44));
    layer0_outputs(4493) <= '0';
    layer0_outputs(4494) <= '1';
    layer0_outputs(4495) <= not((inputs(203)) or (inputs(115)));
    layer0_outputs(4496) <= not(inputs(174));
    layer0_outputs(4497) <= (inputs(53)) or (inputs(129));
    layer0_outputs(4498) <= inputs(14);
    layer0_outputs(4499) <= '0';
    layer0_outputs(4500) <= '1';
    layer0_outputs(4501) <= '1';
    layer0_outputs(4502) <= '0';
    layer0_outputs(4503) <= '1';
    layer0_outputs(4504) <= inputs(118);
    layer0_outputs(4505) <= not((inputs(132)) or (inputs(229)));
    layer0_outputs(4506) <= not(inputs(226)) or (inputs(0));
    layer0_outputs(4507) <= '1';
    layer0_outputs(4508) <= '1';
    layer0_outputs(4509) <= '0';
    layer0_outputs(4510) <= '0';
    layer0_outputs(4511) <= '1';
    layer0_outputs(4512) <= not(inputs(241)) or (inputs(47));
    layer0_outputs(4513) <= inputs(113);
    layer0_outputs(4514) <= '1';
    layer0_outputs(4515) <= (inputs(6)) and (inputs(85));
    layer0_outputs(4516) <= inputs(12);
    layer0_outputs(4517) <= '0';
    layer0_outputs(4518) <= not(inputs(72)) or (inputs(244));
    layer0_outputs(4519) <= '0';
    layer0_outputs(4520) <= not(inputs(88)) or (inputs(155));
    layer0_outputs(4521) <= '0';
    layer0_outputs(4522) <= (inputs(164)) xor (inputs(135));
    layer0_outputs(4523) <= not(inputs(62)) or (inputs(15));
    layer0_outputs(4524) <= not(inputs(172)) or (inputs(33));
    layer0_outputs(4525) <= inputs(69);
    layer0_outputs(4526) <= '1';
    layer0_outputs(4527) <= (inputs(20)) and not (inputs(143));
    layer0_outputs(4528) <= '1';
    layer0_outputs(4529) <= not(inputs(22));
    layer0_outputs(4530) <= '1';
    layer0_outputs(4531) <= '0';
    layer0_outputs(4532) <= '0';
    layer0_outputs(4533) <= (inputs(116)) and not (inputs(191));
    layer0_outputs(4534) <= not((inputs(175)) and (inputs(175)));
    layer0_outputs(4535) <= (inputs(107)) and not (inputs(55));
    layer0_outputs(4536) <= '0';
    layer0_outputs(4537) <= not(inputs(176));
    layer0_outputs(4538) <= not(inputs(158));
    layer0_outputs(4539) <= (inputs(224)) or (inputs(17));
    layer0_outputs(4540) <= (inputs(160)) and (inputs(8));
    layer0_outputs(4541) <= not(inputs(248));
    layer0_outputs(4542) <= '0';
    layer0_outputs(4543) <= not(inputs(130));
    layer0_outputs(4544) <= not(inputs(232));
    layer0_outputs(4545) <= not(inputs(95));
    layer0_outputs(4546) <= '1';
    layer0_outputs(4547) <= not(inputs(159));
    layer0_outputs(4548) <= '0';
    layer0_outputs(4549) <= '0';
    layer0_outputs(4550) <= (inputs(25)) and (inputs(0));
    layer0_outputs(4551) <= not((inputs(71)) or (inputs(148)));
    layer0_outputs(4552) <= not(inputs(77)) or (inputs(173));
    layer0_outputs(4553) <= (inputs(46)) and not (inputs(57));
    layer0_outputs(4554) <= not((inputs(128)) or (inputs(173)));
    layer0_outputs(4555) <= '1';
    layer0_outputs(4556) <= not(inputs(18)) or (inputs(226));
    layer0_outputs(4557) <= not((inputs(79)) and (inputs(18)));
    layer0_outputs(4558) <= inputs(45);
    layer0_outputs(4559) <= (inputs(215)) or (inputs(88));
    layer0_outputs(4560) <= not((inputs(105)) xor (inputs(111)));
    layer0_outputs(4561) <= (inputs(89)) and not (inputs(93));
    layer0_outputs(4562) <= (inputs(176)) and not (inputs(247));
    layer0_outputs(4563) <= inputs(237);
    layer0_outputs(4564) <= '1';
    layer0_outputs(4565) <= (inputs(221)) and not (inputs(155));
    layer0_outputs(4566) <= (inputs(194)) or (inputs(69));
    layer0_outputs(4567) <= '1';
    layer0_outputs(4568) <= not(inputs(28)) or (inputs(65));
    layer0_outputs(4569) <= inputs(193);
    layer0_outputs(4570) <= inputs(218);
    layer0_outputs(4571) <= not(inputs(89)) or (inputs(76));
    layer0_outputs(4572) <= '1';
    layer0_outputs(4573) <= (inputs(172)) and (inputs(190));
    layer0_outputs(4574) <= (inputs(11)) and not (inputs(43));
    layer0_outputs(4575) <= (inputs(125)) and not (inputs(226));
    layer0_outputs(4576) <= not((inputs(166)) and (inputs(28)));
    layer0_outputs(4577) <= (inputs(244)) or (inputs(110));
    layer0_outputs(4578) <= '1';
    layer0_outputs(4579) <= inputs(151);
    layer0_outputs(4580) <= not(inputs(123));
    layer0_outputs(4581) <= (inputs(220)) or (inputs(126));
    layer0_outputs(4582) <= (inputs(193)) and not (inputs(165));
    layer0_outputs(4583) <= inputs(13);
    layer0_outputs(4584) <= not((inputs(213)) or (inputs(154)));
    layer0_outputs(4585) <= not(inputs(68));
    layer0_outputs(4586) <= '0';
    layer0_outputs(4587) <= (inputs(247)) and not (inputs(53));
    layer0_outputs(4588) <= not(inputs(137));
    layer0_outputs(4589) <= (inputs(126)) and not (inputs(143));
    layer0_outputs(4590) <= inputs(166);
    layer0_outputs(4591) <= '1';
    layer0_outputs(4592) <= (inputs(1)) and (inputs(192));
    layer0_outputs(4593) <= not((inputs(16)) and (inputs(53)));
    layer0_outputs(4594) <= inputs(151);
    layer0_outputs(4595) <= '0';
    layer0_outputs(4596) <= '0';
    layer0_outputs(4597) <= not(inputs(57));
    layer0_outputs(4598) <= not(inputs(226)) or (inputs(114));
    layer0_outputs(4599) <= inputs(30);
    layer0_outputs(4600) <= not(inputs(136));
    layer0_outputs(4601) <= (inputs(225)) and not (inputs(91));
    layer0_outputs(4602) <= '1';
    layer0_outputs(4603) <= not(inputs(175));
    layer0_outputs(4604) <= inputs(254);
    layer0_outputs(4605) <= (inputs(80)) and not (inputs(220));
    layer0_outputs(4606) <= not(inputs(242));
    layer0_outputs(4607) <= (inputs(72)) and not (inputs(249));
    layer0_outputs(4608) <= (inputs(14)) or (inputs(51));
    layer0_outputs(4609) <= '0';
    layer0_outputs(4610) <= '0';
    layer0_outputs(4611) <= '1';
    layer0_outputs(4612) <= not((inputs(128)) and (inputs(0)));
    layer0_outputs(4613) <= not(inputs(90)) or (inputs(208));
    layer0_outputs(4614) <= '0';
    layer0_outputs(4615) <= '1';
    layer0_outputs(4616) <= inputs(34);
    layer0_outputs(4617) <= not(inputs(65));
    layer0_outputs(4618) <= '0';
    layer0_outputs(4619) <= (inputs(191)) or (inputs(210));
    layer0_outputs(4620) <= not((inputs(249)) and (inputs(241)));
    layer0_outputs(4621) <= not(inputs(148)) or (inputs(226));
    layer0_outputs(4622) <= '0';
    layer0_outputs(4623) <= '0';
    layer0_outputs(4624) <= inputs(117);
    layer0_outputs(4625) <= not(inputs(106));
    layer0_outputs(4626) <= (inputs(212)) xor (inputs(234));
    layer0_outputs(4627) <= '1';
    layer0_outputs(4628) <= not(inputs(4)) or (inputs(189));
    layer0_outputs(4629) <= not(inputs(167));
    layer0_outputs(4630) <= not((inputs(243)) and (inputs(254)));
    layer0_outputs(4631) <= (inputs(70)) and not (inputs(201));
    layer0_outputs(4632) <= '1';
    layer0_outputs(4633) <= not(inputs(220)) or (inputs(206));
    layer0_outputs(4634) <= not(inputs(127)) or (inputs(194));
    layer0_outputs(4635) <= '0';
    layer0_outputs(4636) <= not((inputs(52)) and (inputs(9)));
    layer0_outputs(4637) <= not(inputs(244));
    layer0_outputs(4638) <= not(inputs(52));
    layer0_outputs(4639) <= inputs(113);
    layer0_outputs(4640) <= not((inputs(81)) or (inputs(197)));
    layer0_outputs(4641) <= '0';
    layer0_outputs(4642) <= '0';
    layer0_outputs(4643) <= '1';
    layer0_outputs(4644) <= not(inputs(244)) or (inputs(147));
    layer0_outputs(4645) <= (inputs(180)) and (inputs(173));
    layer0_outputs(4646) <= (inputs(3)) xor (inputs(204));
    layer0_outputs(4647) <= not(inputs(198)) or (inputs(61));
    layer0_outputs(4648) <= '1';
    layer0_outputs(4649) <= not(inputs(18)) or (inputs(93));
    layer0_outputs(4650) <= not((inputs(204)) or (inputs(157)));
    layer0_outputs(4651) <= '1';
    layer0_outputs(4652) <= (inputs(19)) or (inputs(43));
    layer0_outputs(4653) <= '0';
    layer0_outputs(4654) <= not(inputs(228)) or (inputs(254));
    layer0_outputs(4655) <= not(inputs(19));
    layer0_outputs(4656) <= not(inputs(170)) or (inputs(22));
    layer0_outputs(4657) <= not(inputs(80)) or (inputs(13));
    layer0_outputs(4658) <= (inputs(9)) and not (inputs(143));
    layer0_outputs(4659) <= inputs(142);
    layer0_outputs(4660) <= inputs(86);
    layer0_outputs(4661) <= not((inputs(91)) and (inputs(96)));
    layer0_outputs(4662) <= not(inputs(158));
    layer0_outputs(4663) <= '1';
    layer0_outputs(4664) <= '1';
    layer0_outputs(4665) <= '0';
    layer0_outputs(4666) <= (inputs(80)) xor (inputs(170));
    layer0_outputs(4667) <= '1';
    layer0_outputs(4668) <= (inputs(159)) and not (inputs(174));
    layer0_outputs(4669) <= (inputs(32)) and not (inputs(137));
    layer0_outputs(4670) <= not(inputs(131)) or (inputs(119));
    layer0_outputs(4671) <= (inputs(152)) and (inputs(148));
    layer0_outputs(4672) <= not(inputs(77));
    layer0_outputs(4673) <= not(inputs(161)) or (inputs(163));
    layer0_outputs(4674) <= not((inputs(227)) and (inputs(58)));
    layer0_outputs(4675) <= not((inputs(207)) xor (inputs(180)));
    layer0_outputs(4676) <= '0';
    layer0_outputs(4677) <= (inputs(132)) and not (inputs(56));
    layer0_outputs(4678) <= not((inputs(60)) and (inputs(179)));
    layer0_outputs(4679) <= inputs(7);
    layer0_outputs(4680) <= not(inputs(177));
    layer0_outputs(4681) <= '1';
    layer0_outputs(4682) <= '0';
    layer0_outputs(4683) <= '1';
    layer0_outputs(4684) <= '1';
    layer0_outputs(4685) <= not((inputs(129)) and (inputs(119)));
    layer0_outputs(4686) <= not(inputs(140)) or (inputs(124));
    layer0_outputs(4687) <= not((inputs(4)) xor (inputs(254)));
    layer0_outputs(4688) <= not(inputs(183));
    layer0_outputs(4689) <= not(inputs(59));
    layer0_outputs(4690) <= '0';
    layer0_outputs(4691) <= not(inputs(232)) or (inputs(162));
    layer0_outputs(4692) <= not((inputs(221)) xor (inputs(208)));
    layer0_outputs(4693) <= not(inputs(72)) or (inputs(101));
    layer0_outputs(4694) <= inputs(44);
    layer0_outputs(4695) <= not(inputs(154));
    layer0_outputs(4696) <= not(inputs(166));
    layer0_outputs(4697) <= inputs(24);
    layer0_outputs(4698) <= not((inputs(139)) xor (inputs(248)));
    layer0_outputs(4699) <= inputs(153);
    layer0_outputs(4700) <= (inputs(242)) and not (inputs(254));
    layer0_outputs(4701) <= not(inputs(10)) or (inputs(134));
    layer0_outputs(4702) <= '1';
    layer0_outputs(4703) <= not(inputs(231)) or (inputs(254));
    layer0_outputs(4704) <= not(inputs(207));
    layer0_outputs(4705) <= not((inputs(238)) and (inputs(254)));
    layer0_outputs(4706) <= '1';
    layer0_outputs(4707) <= inputs(25);
    layer0_outputs(4708) <= not(inputs(25)) or (inputs(157));
    layer0_outputs(4709) <= not(inputs(144));
    layer0_outputs(4710) <= not((inputs(247)) xor (inputs(43)));
    layer0_outputs(4711) <= not(inputs(112));
    layer0_outputs(4712) <= inputs(167);
    layer0_outputs(4713) <= (inputs(228)) and not (inputs(113));
    layer0_outputs(4714) <= not((inputs(46)) or (inputs(22)));
    layer0_outputs(4715) <= not((inputs(207)) and (inputs(6)));
    layer0_outputs(4716) <= (inputs(159)) and (inputs(21));
    layer0_outputs(4717) <= '1';
    layer0_outputs(4718) <= inputs(86);
    layer0_outputs(4719) <= (inputs(224)) and not (inputs(219));
    layer0_outputs(4720) <= not(inputs(253)) or (inputs(59));
    layer0_outputs(4721) <= not(inputs(80));
    layer0_outputs(4722) <= inputs(44);
    layer0_outputs(4723) <= '1';
    layer0_outputs(4724) <= inputs(243);
    layer0_outputs(4725) <= not(inputs(45));
    layer0_outputs(4726) <= not(inputs(38)) or (inputs(145));
    layer0_outputs(4727) <= not((inputs(162)) or (inputs(93)));
    layer0_outputs(4728) <= (inputs(129)) xor (inputs(163));
    layer0_outputs(4729) <= inputs(202);
    layer0_outputs(4730) <= not((inputs(125)) and (inputs(180)));
    layer0_outputs(4731) <= inputs(144);
    layer0_outputs(4732) <= not(inputs(102)) or (inputs(119));
    layer0_outputs(4733) <= (inputs(200)) and (inputs(115));
    layer0_outputs(4734) <= '1';
    layer0_outputs(4735) <= inputs(163);
    layer0_outputs(4736) <= (inputs(75)) and not (inputs(53));
    layer0_outputs(4737) <= not(inputs(147)) or (inputs(200));
    layer0_outputs(4738) <= (inputs(158)) and (inputs(172));
    layer0_outputs(4739) <= '1';
    layer0_outputs(4740) <= '1';
    layer0_outputs(4741) <= '0';
    layer0_outputs(4742) <= (inputs(9)) and (inputs(17));
    layer0_outputs(4743) <= (inputs(99)) or (inputs(225));
    layer0_outputs(4744) <= '0';
    layer0_outputs(4745) <= '1';
    layer0_outputs(4746) <= not((inputs(48)) or (inputs(175)));
    layer0_outputs(4747) <= not(inputs(156));
    layer0_outputs(4748) <= not((inputs(227)) and (inputs(50)));
    layer0_outputs(4749) <= not(inputs(194));
    layer0_outputs(4750) <= not(inputs(93));
    layer0_outputs(4751) <= not(inputs(240));
    layer0_outputs(4752) <= (inputs(82)) and (inputs(47));
    layer0_outputs(4753) <= (inputs(242)) and not (inputs(185));
    layer0_outputs(4754) <= not(inputs(199)) or (inputs(34));
    layer0_outputs(4755) <= not(inputs(88)) or (inputs(31));
    layer0_outputs(4756) <= not((inputs(116)) or (inputs(248)));
    layer0_outputs(4757) <= not(inputs(136)) or (inputs(202));
    layer0_outputs(4758) <= (inputs(242)) or (inputs(154));
    layer0_outputs(4759) <= '0';
    layer0_outputs(4760) <= '1';
    layer0_outputs(4761) <= '0';
    layer0_outputs(4762) <= (inputs(210)) or (inputs(40));
    layer0_outputs(4763) <= inputs(62);
    layer0_outputs(4764) <= not(inputs(92));
    layer0_outputs(4765) <= not(inputs(109)) or (inputs(147));
    layer0_outputs(4766) <= (inputs(127)) and not (inputs(154));
    layer0_outputs(4767) <= not(inputs(144)) or (inputs(58));
    layer0_outputs(4768) <= not((inputs(223)) and (inputs(110)));
    layer0_outputs(4769) <= (inputs(181)) and not (inputs(106));
    layer0_outputs(4770) <= '0';
    layer0_outputs(4771) <= (inputs(185)) and (inputs(205));
    layer0_outputs(4772) <= not(inputs(154)) or (inputs(115));
    layer0_outputs(4773) <= '0';
    layer0_outputs(4774) <= not((inputs(138)) and (inputs(175)));
    layer0_outputs(4775) <= '1';
    layer0_outputs(4776) <= not(inputs(133)) or (inputs(149));
    layer0_outputs(4777) <= '0';
    layer0_outputs(4778) <= '0';
    layer0_outputs(4779) <= inputs(136);
    layer0_outputs(4780) <= '1';
    layer0_outputs(4781) <= '0';
    layer0_outputs(4782) <= (inputs(82)) or (inputs(126));
    layer0_outputs(4783) <= not(inputs(130));
    layer0_outputs(4784) <= inputs(158);
    layer0_outputs(4785) <= (inputs(210)) or (inputs(149));
    layer0_outputs(4786) <= (inputs(117)) and not (inputs(11));
    layer0_outputs(4787) <= not((inputs(233)) and (inputs(88)));
    layer0_outputs(4788) <= (inputs(232)) and not (inputs(111));
    layer0_outputs(4789) <= (inputs(17)) and not (inputs(182));
    layer0_outputs(4790) <= '0';
    layer0_outputs(4791) <= (inputs(16)) and (inputs(205));
    layer0_outputs(4792) <= (inputs(168)) and not (inputs(214));
    layer0_outputs(4793) <= (inputs(202)) and not (inputs(110));
    layer0_outputs(4794) <= not((inputs(217)) and (inputs(225)));
    layer0_outputs(4795) <= not((inputs(164)) or (inputs(133)));
    layer0_outputs(4796) <= (inputs(212)) and (inputs(135));
    layer0_outputs(4797) <= not(inputs(29));
    layer0_outputs(4798) <= '0';
    layer0_outputs(4799) <= (inputs(215)) and (inputs(111));
    layer0_outputs(4800) <= (inputs(31)) and not (inputs(56));
    layer0_outputs(4801) <= '1';
    layer0_outputs(4802) <= not(inputs(254));
    layer0_outputs(4803) <= not(inputs(89)) or (inputs(156));
    layer0_outputs(4804) <= '1';
    layer0_outputs(4805) <= '0';
    layer0_outputs(4806) <= (inputs(187)) and not (inputs(41));
    layer0_outputs(4807) <= '1';
    layer0_outputs(4808) <= not((inputs(56)) or (inputs(37)));
    layer0_outputs(4809) <= inputs(238);
    layer0_outputs(4810) <= inputs(44);
    layer0_outputs(4811) <= not((inputs(66)) and (inputs(106)));
    layer0_outputs(4812) <= (inputs(131)) and not (inputs(120));
    layer0_outputs(4813) <= '0';
    layer0_outputs(4814) <= not(inputs(34));
    layer0_outputs(4815) <= inputs(60);
    layer0_outputs(4816) <= '1';
    layer0_outputs(4817) <= (inputs(68)) and (inputs(92));
    layer0_outputs(4818) <= '0';
    layer0_outputs(4819) <= not(inputs(20)) or (inputs(72));
    layer0_outputs(4820) <= not((inputs(126)) and (inputs(226)));
    layer0_outputs(4821) <= '1';
    layer0_outputs(4822) <= not((inputs(221)) or (inputs(158)));
    layer0_outputs(4823) <= (inputs(219)) or (inputs(220));
    layer0_outputs(4824) <= not((inputs(249)) and (inputs(234)));
    layer0_outputs(4825) <= (inputs(67)) or (inputs(15));
    layer0_outputs(4826) <= not(inputs(234));
    layer0_outputs(4827) <= not((inputs(212)) and (inputs(56)));
    layer0_outputs(4828) <= (inputs(128)) and not (inputs(146));
    layer0_outputs(4829) <= '0';
    layer0_outputs(4830) <= '1';
    layer0_outputs(4831) <= '0';
    layer0_outputs(4832) <= not(inputs(108));
    layer0_outputs(4833) <= '0';
    layer0_outputs(4834) <= '0';
    layer0_outputs(4835) <= not(inputs(65)) or (inputs(86));
    layer0_outputs(4836) <= not(inputs(22)) or (inputs(58));
    layer0_outputs(4837) <= '0';
    layer0_outputs(4838) <= not((inputs(200)) and (inputs(21)));
    layer0_outputs(4839) <= not(inputs(157)) or (inputs(168));
    layer0_outputs(4840) <= not(inputs(65)) or (inputs(245));
    layer0_outputs(4841) <= not((inputs(223)) or (inputs(198)));
    layer0_outputs(4842) <= inputs(254);
    layer0_outputs(4843) <= not(inputs(14)) or (inputs(169));
    layer0_outputs(4844) <= '1';
    layer0_outputs(4845) <= not(inputs(7)) or (inputs(98));
    layer0_outputs(4846) <= '0';
    layer0_outputs(4847) <= not((inputs(101)) xor (inputs(131)));
    layer0_outputs(4848) <= (inputs(0)) and not (inputs(137));
    layer0_outputs(4849) <= not(inputs(194));
    layer0_outputs(4850) <= not(inputs(15)) or (inputs(35));
    layer0_outputs(4851) <= not(inputs(121)) or (inputs(236));
    layer0_outputs(4852) <= not((inputs(173)) and (inputs(168)));
    layer0_outputs(4853) <= '0';
    layer0_outputs(4854) <= '0';
    layer0_outputs(4855) <= not(inputs(84)) or (inputs(239));
    layer0_outputs(4856) <= inputs(1);
    layer0_outputs(4857) <= '1';
    layer0_outputs(4858) <= not(inputs(41));
    layer0_outputs(4859) <= not(inputs(111)) or (inputs(136));
    layer0_outputs(4860) <= (inputs(191)) and not (inputs(34));
    layer0_outputs(4861) <= inputs(130);
    layer0_outputs(4862) <= (inputs(177)) and not (inputs(207));
    layer0_outputs(4863) <= (inputs(163)) and (inputs(22));
    layer0_outputs(4864) <= (inputs(198)) and not (inputs(235));
    layer0_outputs(4865) <= not(inputs(237));
    layer0_outputs(4866) <= inputs(90);
    layer0_outputs(4867) <= not((inputs(55)) and (inputs(247)));
    layer0_outputs(4868) <= (inputs(59)) and not (inputs(169));
    layer0_outputs(4869) <= not((inputs(89)) or (inputs(205)));
    layer0_outputs(4870) <= inputs(92);
    layer0_outputs(4871) <= (inputs(92)) and (inputs(52));
    layer0_outputs(4872) <= '0';
    layer0_outputs(4873) <= (inputs(25)) or (inputs(221));
    layer0_outputs(4874) <= inputs(198);
    layer0_outputs(4875) <= '0';
    layer0_outputs(4876) <= (inputs(218)) and not (inputs(182));
    layer0_outputs(4877) <= not(inputs(107)) or (inputs(43));
    layer0_outputs(4878) <= '1';
    layer0_outputs(4879) <= '0';
    layer0_outputs(4880) <= not((inputs(175)) xor (inputs(102)));
    layer0_outputs(4881) <= not((inputs(216)) and (inputs(114)));
    layer0_outputs(4882) <= not((inputs(60)) or (inputs(83)));
    layer0_outputs(4883) <= not(inputs(240));
    layer0_outputs(4884) <= '0';
    layer0_outputs(4885) <= not(inputs(113));
    layer0_outputs(4886) <= '1';
    layer0_outputs(4887) <= '1';
    layer0_outputs(4888) <= not((inputs(207)) xor (inputs(29)));
    layer0_outputs(4889) <= not(inputs(252)) or (inputs(178));
    layer0_outputs(4890) <= (inputs(229)) and not (inputs(248));
    layer0_outputs(4891) <= '0';
    layer0_outputs(4892) <= (inputs(158)) xor (inputs(175));
    layer0_outputs(4893) <= not(inputs(128));
    layer0_outputs(4894) <= (inputs(53)) and (inputs(0));
    layer0_outputs(4895) <= (inputs(16)) xor (inputs(136));
    layer0_outputs(4896) <= not(inputs(144));
    layer0_outputs(4897) <= '1';
    layer0_outputs(4898) <= (inputs(9)) and not (inputs(178));
    layer0_outputs(4899) <= (inputs(213)) and not (inputs(195));
    layer0_outputs(4900) <= inputs(124);
    layer0_outputs(4901) <= not(inputs(176));
    layer0_outputs(4902) <= not((inputs(15)) and (inputs(98)));
    layer0_outputs(4903) <= '0';
    layer0_outputs(4904) <= not(inputs(165));
    layer0_outputs(4905) <= not(inputs(223)) or (inputs(164));
    layer0_outputs(4906) <= not(inputs(156)) or (inputs(8));
    layer0_outputs(4907) <= (inputs(63)) and not (inputs(28));
    layer0_outputs(4908) <= not(inputs(241));
    layer0_outputs(4909) <= '0';
    layer0_outputs(4910) <= not(inputs(189)) or (inputs(33));
    layer0_outputs(4911) <= (inputs(189)) and not (inputs(142));
    layer0_outputs(4912) <= '0';
    layer0_outputs(4913) <= inputs(218);
    layer0_outputs(4914) <= (inputs(120)) and not (inputs(176));
    layer0_outputs(4915) <= inputs(87);
    layer0_outputs(4916) <= not(inputs(209)) or (inputs(91));
    layer0_outputs(4917) <= (inputs(15)) and not (inputs(197));
    layer0_outputs(4918) <= '0';
    layer0_outputs(4919) <= '1';
    layer0_outputs(4920) <= '0';
    layer0_outputs(4921) <= '1';
    layer0_outputs(4922) <= not(inputs(194));
    layer0_outputs(4923) <= (inputs(8)) and not (inputs(192));
    layer0_outputs(4924) <= not((inputs(203)) or (inputs(115)));
    layer0_outputs(4925) <= (inputs(233)) and (inputs(98));
    layer0_outputs(4926) <= '1';
    layer0_outputs(4927) <= '1';
    layer0_outputs(4928) <= not(inputs(160)) or (inputs(172));
    layer0_outputs(4929) <= '0';
    layer0_outputs(4930) <= not(inputs(38));
    layer0_outputs(4931) <= not((inputs(250)) and (inputs(23)));
    layer0_outputs(4932) <= '1';
    layer0_outputs(4933) <= not(inputs(146));
    layer0_outputs(4934) <= '1';
    layer0_outputs(4935) <= not((inputs(68)) or (inputs(214)));
    layer0_outputs(4936) <= not(inputs(68));
    layer0_outputs(4937) <= not((inputs(67)) and (inputs(90)));
    layer0_outputs(4938) <= '0';
    layer0_outputs(4939) <= '1';
    layer0_outputs(4940) <= inputs(104);
    layer0_outputs(4941) <= (inputs(215)) and not (inputs(216));
    layer0_outputs(4942) <= (inputs(21)) and not (inputs(238));
    layer0_outputs(4943) <= inputs(2);
    layer0_outputs(4944) <= (inputs(13)) xor (inputs(174));
    layer0_outputs(4945) <= not(inputs(166)) or (inputs(128));
    layer0_outputs(4946) <= '1';
    layer0_outputs(4947) <= not(inputs(227)) or (inputs(129));
    layer0_outputs(4948) <= inputs(125);
    layer0_outputs(4949) <= not(inputs(94));
    layer0_outputs(4950) <= inputs(115);
    layer0_outputs(4951) <= '0';
    layer0_outputs(4952) <= not(inputs(185));
    layer0_outputs(4953) <= '1';
    layer0_outputs(4954) <= not(inputs(97));
    layer0_outputs(4955) <= inputs(168);
    layer0_outputs(4956) <= '0';
    layer0_outputs(4957) <= (inputs(35)) and (inputs(196));
    layer0_outputs(4958) <= '1';
    layer0_outputs(4959) <= '1';
    layer0_outputs(4960) <= '0';
    layer0_outputs(4961) <= not(inputs(17)) or (inputs(221));
    layer0_outputs(4962) <= not(inputs(78)) or (inputs(164));
    layer0_outputs(4963) <= '0';
    layer0_outputs(4964) <= (inputs(254)) and not (inputs(226));
    layer0_outputs(4965) <= not(inputs(223));
    layer0_outputs(4966) <= not((inputs(135)) and (inputs(254)));
    layer0_outputs(4967) <= not(inputs(108));
    layer0_outputs(4968) <= (inputs(140)) or (inputs(74));
    layer0_outputs(4969) <= '0';
    layer0_outputs(4970) <= '0';
    layer0_outputs(4971) <= '0';
    layer0_outputs(4972) <= (inputs(123)) and not (inputs(7));
    layer0_outputs(4973) <= (inputs(193)) and not (inputs(125));
    layer0_outputs(4974) <= inputs(97);
    layer0_outputs(4975) <= not((inputs(166)) and (inputs(127)));
    layer0_outputs(4976) <= inputs(141);
    layer0_outputs(4977) <= '1';
    layer0_outputs(4978) <= '0';
    layer0_outputs(4979) <= not(inputs(66)) or (inputs(89));
    layer0_outputs(4980) <= '1';
    layer0_outputs(4981) <= (inputs(93)) and not (inputs(185));
    layer0_outputs(4982) <= inputs(108);
    layer0_outputs(4983) <= '0';
    layer0_outputs(4984) <= inputs(23);
    layer0_outputs(4985) <= (inputs(11)) or (inputs(121));
    layer0_outputs(4986) <= '0';
    layer0_outputs(4987) <= not(inputs(115)) or (inputs(182));
    layer0_outputs(4988) <= not(inputs(52));
    layer0_outputs(4989) <= (inputs(19)) and not (inputs(240));
    layer0_outputs(4990) <= '1';
    layer0_outputs(4991) <= '1';
    layer0_outputs(4992) <= (inputs(46)) and (inputs(2));
    layer0_outputs(4993) <= '0';
    layer0_outputs(4994) <= (inputs(229)) xor (inputs(45));
    layer0_outputs(4995) <= '0';
    layer0_outputs(4996) <= not((inputs(43)) and (inputs(14)));
    layer0_outputs(4997) <= '1';
    layer0_outputs(4998) <= '1';
    layer0_outputs(4999) <= (inputs(130)) and (inputs(82));
    layer0_outputs(5000) <= '0';
    layer0_outputs(5001) <= '1';
    layer0_outputs(5002) <= (inputs(95)) xor (inputs(24));
    layer0_outputs(5003) <= not(inputs(237)) or (inputs(1));
    layer0_outputs(5004) <= '0';
    layer0_outputs(5005) <= '1';
    layer0_outputs(5006) <= not((inputs(61)) or (inputs(32)));
    layer0_outputs(5007) <= (inputs(181)) and (inputs(58));
    layer0_outputs(5008) <= (inputs(126)) and not (inputs(117));
    layer0_outputs(5009) <= not((inputs(253)) and (inputs(255)));
    layer0_outputs(5010) <= not((inputs(130)) or (inputs(140)));
    layer0_outputs(5011) <= (inputs(192)) or (inputs(40));
    layer0_outputs(5012) <= inputs(222);
    layer0_outputs(5013) <= '0';
    layer0_outputs(5014) <= not(inputs(236));
    layer0_outputs(5015) <= (inputs(64)) xor (inputs(144));
    layer0_outputs(5016) <= not(inputs(90)) or (inputs(128));
    layer0_outputs(5017) <= inputs(107);
    layer0_outputs(5018) <= '0';
    layer0_outputs(5019) <= '0';
    layer0_outputs(5020) <= not((inputs(35)) or (inputs(178)));
    layer0_outputs(5021) <= (inputs(201)) or (inputs(161));
    layer0_outputs(5022) <= not(inputs(127)) or (inputs(58));
    layer0_outputs(5023) <= inputs(8);
    layer0_outputs(5024) <= '0';
    layer0_outputs(5025) <= '1';
    layer0_outputs(5026) <= inputs(254);
    layer0_outputs(5027) <= (inputs(28)) and (inputs(9));
    layer0_outputs(5028) <= not(inputs(149)) or (inputs(31));
    layer0_outputs(5029) <= not(inputs(173)) or (inputs(44));
    layer0_outputs(5030) <= (inputs(26)) xor (inputs(236));
    layer0_outputs(5031) <= not(inputs(44));
    layer0_outputs(5032) <= inputs(187);
    layer0_outputs(5033) <= (inputs(25)) and not (inputs(149));
    layer0_outputs(5034) <= not((inputs(164)) xor (inputs(242)));
    layer0_outputs(5035) <= '1';
    layer0_outputs(5036) <= '0';
    layer0_outputs(5037) <= (inputs(64)) and not (inputs(134));
    layer0_outputs(5038) <= inputs(62);
    layer0_outputs(5039) <= '0';
    layer0_outputs(5040) <= not((inputs(46)) or (inputs(76)));
    layer0_outputs(5041) <= (inputs(202)) and not (inputs(118));
    layer0_outputs(5042) <= not(inputs(83)) or (inputs(227));
    layer0_outputs(5043) <= (inputs(179)) and not (inputs(32));
    layer0_outputs(5044) <= not((inputs(60)) or (inputs(175)));
    layer0_outputs(5045) <= not((inputs(13)) and (inputs(73)));
    layer0_outputs(5046) <= '1';
    layer0_outputs(5047) <= not(inputs(156));
    layer0_outputs(5048) <= inputs(239);
    layer0_outputs(5049) <= (inputs(62)) and (inputs(130));
    layer0_outputs(5050) <= (inputs(211)) and not (inputs(149));
    layer0_outputs(5051) <= '1';
    layer0_outputs(5052) <= inputs(57);
    layer0_outputs(5053) <= not((inputs(65)) xor (inputs(1)));
    layer0_outputs(5054) <= '0';
    layer0_outputs(5055) <= not(inputs(128)) or (inputs(63));
    layer0_outputs(5056) <= not(inputs(223)) or (inputs(37));
    layer0_outputs(5057) <= inputs(246);
    layer0_outputs(5058) <= (inputs(173)) and not (inputs(155));
    layer0_outputs(5059) <= (inputs(69)) or (inputs(234));
    layer0_outputs(5060) <= (inputs(193)) or (inputs(165));
    layer0_outputs(5061) <= inputs(106);
    layer0_outputs(5062) <= not(inputs(162)) or (inputs(180));
    layer0_outputs(5063) <= '0';
    layer0_outputs(5064) <= '0';
    layer0_outputs(5065) <= inputs(117);
    layer0_outputs(5066) <= not(inputs(193)) or (inputs(162));
    layer0_outputs(5067) <= inputs(251);
    layer0_outputs(5068) <= (inputs(139)) or (inputs(153));
    layer0_outputs(5069) <= '1';
    layer0_outputs(5070) <= (inputs(206)) and (inputs(132));
    layer0_outputs(5071) <= '0';
    layer0_outputs(5072) <= '1';
    layer0_outputs(5073) <= not(inputs(6)) or (inputs(200));
    layer0_outputs(5074) <= not(inputs(232));
    layer0_outputs(5075) <= not((inputs(245)) or (inputs(70)));
    layer0_outputs(5076) <= not(inputs(163));
    layer0_outputs(5077) <= '1';
    layer0_outputs(5078) <= not(inputs(63));
    layer0_outputs(5079) <= '0';
    layer0_outputs(5080) <= not((inputs(138)) or (inputs(145)));
    layer0_outputs(5081) <= not((inputs(156)) or (inputs(108)));
    layer0_outputs(5082) <= not(inputs(165));
    layer0_outputs(5083) <= (inputs(41)) or (inputs(208));
    layer0_outputs(5084) <= '1';
    layer0_outputs(5085) <= not(inputs(223));
    layer0_outputs(5086) <= not(inputs(242));
    layer0_outputs(5087) <= (inputs(28)) and not (inputs(136));
    layer0_outputs(5088) <= (inputs(186)) or (inputs(191));
    layer0_outputs(5089) <= not(inputs(149)) or (inputs(158));
    layer0_outputs(5090) <= '0';
    layer0_outputs(5091) <= not(inputs(194)) or (inputs(40));
    layer0_outputs(5092) <= inputs(251);
    layer0_outputs(5093) <= not(inputs(124)) or (inputs(92));
    layer0_outputs(5094) <= '0';
    layer0_outputs(5095) <= '1';
    layer0_outputs(5096) <= not(inputs(164)) or (inputs(83));
    layer0_outputs(5097) <= '1';
    layer0_outputs(5098) <= not((inputs(129)) or (inputs(213)));
    layer0_outputs(5099) <= inputs(202);
    layer0_outputs(5100) <= not(inputs(158));
    layer0_outputs(5101) <= '1';
    layer0_outputs(5102) <= not(inputs(120));
    layer0_outputs(5103) <= (inputs(192)) and (inputs(106));
    layer0_outputs(5104) <= '0';
    layer0_outputs(5105) <= not(inputs(16));
    layer0_outputs(5106) <= not(inputs(86));
    layer0_outputs(5107) <= not(inputs(96));
    layer0_outputs(5108) <= (inputs(138)) or (inputs(125));
    layer0_outputs(5109) <= '1';
    layer0_outputs(5110) <= not(inputs(144)) or (inputs(42));
    layer0_outputs(5111) <= inputs(187);
    layer0_outputs(5112) <= not(inputs(94)) or (inputs(234));
    layer0_outputs(5113) <= '1';
    layer0_outputs(5114) <= not(inputs(252));
    layer0_outputs(5115) <= '0';
    layer0_outputs(5116) <= not(inputs(204)) or (inputs(129));
    layer0_outputs(5117) <= not((inputs(217)) and (inputs(181)));
    layer0_outputs(5118) <= not(inputs(253));
    layer0_outputs(5119) <= inputs(241);
    layer1_outputs(0) <= layer0_outputs(3228);
    layer1_outputs(1) <= not((layer0_outputs(585)) or (layer0_outputs(36)));
    layer1_outputs(2) <= not(layer0_outputs(471));
    layer1_outputs(3) <= '1';
    layer1_outputs(4) <= '1';
    layer1_outputs(5) <= not(layer0_outputs(1694));
    layer1_outputs(6) <= (layer0_outputs(3751)) and not (layer0_outputs(680));
    layer1_outputs(7) <= '0';
    layer1_outputs(8) <= not((layer0_outputs(907)) xor (layer0_outputs(1031)));
    layer1_outputs(9) <= '1';
    layer1_outputs(10) <= not((layer0_outputs(3599)) and (layer0_outputs(2384)));
    layer1_outputs(11) <= layer0_outputs(4006);
    layer1_outputs(12) <= not(layer0_outputs(2270)) or (layer0_outputs(4820));
    layer1_outputs(13) <= not((layer0_outputs(3919)) and (layer0_outputs(3613)));
    layer1_outputs(14) <= '1';
    layer1_outputs(15) <= '0';
    layer1_outputs(16) <= (layer0_outputs(1535)) and not (layer0_outputs(3018));
    layer1_outputs(17) <= '1';
    layer1_outputs(18) <= '1';
    layer1_outputs(19) <= (layer0_outputs(2922)) and not (layer0_outputs(4571));
    layer1_outputs(20) <= (layer0_outputs(4650)) and (layer0_outputs(2856));
    layer1_outputs(21) <= '1';
    layer1_outputs(22) <= not(layer0_outputs(3848));
    layer1_outputs(23) <= not(layer0_outputs(1855)) or (layer0_outputs(2320));
    layer1_outputs(24) <= (layer0_outputs(4150)) or (layer0_outputs(814));
    layer1_outputs(25) <= '1';
    layer1_outputs(26) <= not(layer0_outputs(4183));
    layer1_outputs(27) <= layer0_outputs(1689);
    layer1_outputs(28) <= not((layer0_outputs(1069)) and (layer0_outputs(2989)));
    layer1_outputs(29) <= (layer0_outputs(4213)) and not (layer0_outputs(3224));
    layer1_outputs(30) <= '0';
    layer1_outputs(31) <= (layer0_outputs(3913)) and not (layer0_outputs(162));
    layer1_outputs(32) <= '0';
    layer1_outputs(33) <= not(layer0_outputs(3579)) or (layer0_outputs(2446));
    layer1_outputs(34) <= '0';
    layer1_outputs(35) <= (layer0_outputs(514)) and not (layer0_outputs(4702));
    layer1_outputs(36) <= (layer0_outputs(3598)) or (layer0_outputs(1347));
    layer1_outputs(37) <= not((layer0_outputs(3611)) and (layer0_outputs(3253)));
    layer1_outputs(38) <= not(layer0_outputs(2253)) or (layer0_outputs(4745));
    layer1_outputs(39) <= not(layer0_outputs(1077)) or (layer0_outputs(1973));
    layer1_outputs(40) <= not(layer0_outputs(1230));
    layer1_outputs(41) <= (layer0_outputs(1564)) or (layer0_outputs(3021));
    layer1_outputs(42) <= (layer0_outputs(483)) or (layer0_outputs(1887));
    layer1_outputs(43) <= not(layer0_outputs(2274)) or (layer0_outputs(57));
    layer1_outputs(44) <= layer0_outputs(3770);
    layer1_outputs(45) <= not(layer0_outputs(4895)) or (layer0_outputs(2609));
    layer1_outputs(46) <= '1';
    layer1_outputs(47) <= '0';
    layer1_outputs(48) <= '0';
    layer1_outputs(49) <= not(layer0_outputs(4072)) or (layer0_outputs(3345));
    layer1_outputs(50) <= '0';
    layer1_outputs(51) <= layer0_outputs(4699);
    layer1_outputs(52) <= not((layer0_outputs(4459)) or (layer0_outputs(3187)));
    layer1_outputs(53) <= not((layer0_outputs(2410)) or (layer0_outputs(4952)));
    layer1_outputs(54) <= layer0_outputs(3586);
    layer1_outputs(55) <= layer0_outputs(1443);
    layer1_outputs(56) <= '1';
    layer1_outputs(57) <= (layer0_outputs(4784)) or (layer0_outputs(3573));
    layer1_outputs(58) <= '1';
    layer1_outputs(59) <= not(layer0_outputs(4919));
    layer1_outputs(60) <= not(layer0_outputs(3406)) or (layer0_outputs(4652));
    layer1_outputs(61) <= (layer0_outputs(2043)) or (layer0_outputs(2891));
    layer1_outputs(62) <= '1';
    layer1_outputs(63) <= not(layer0_outputs(1453));
    layer1_outputs(64) <= (layer0_outputs(1113)) or (layer0_outputs(837));
    layer1_outputs(65) <= layer0_outputs(5055);
    layer1_outputs(66) <= not(layer0_outputs(4679));
    layer1_outputs(67) <= (layer0_outputs(3351)) and not (layer0_outputs(4717));
    layer1_outputs(68) <= not(layer0_outputs(2658));
    layer1_outputs(69) <= not(layer0_outputs(3917)) or (layer0_outputs(3615));
    layer1_outputs(70) <= not(layer0_outputs(1860)) or (layer0_outputs(2897));
    layer1_outputs(71) <= layer0_outputs(3236);
    layer1_outputs(72) <= (layer0_outputs(2096)) and not (layer0_outputs(4712));
    layer1_outputs(73) <= (layer0_outputs(444)) and (layer0_outputs(1881));
    layer1_outputs(74) <= (layer0_outputs(1100)) and (layer0_outputs(1997));
    layer1_outputs(75) <= not(layer0_outputs(845)) or (layer0_outputs(2023));
    layer1_outputs(76) <= (layer0_outputs(4117)) and not (layer0_outputs(3541));
    layer1_outputs(77) <= '1';
    layer1_outputs(78) <= (layer0_outputs(576)) or (layer0_outputs(2587));
    layer1_outputs(79) <= (layer0_outputs(3394)) and (layer0_outputs(3623));
    layer1_outputs(80) <= '1';
    layer1_outputs(81) <= not((layer0_outputs(1364)) or (layer0_outputs(2882)));
    layer1_outputs(82) <= layer0_outputs(2835);
    layer1_outputs(83) <= not((layer0_outputs(3556)) or (layer0_outputs(2392)));
    layer1_outputs(84) <= not((layer0_outputs(3707)) or (layer0_outputs(792)));
    layer1_outputs(85) <= not(layer0_outputs(3987));
    layer1_outputs(86) <= not((layer0_outputs(3539)) or (layer0_outputs(1590)));
    layer1_outputs(87) <= '0';
    layer1_outputs(88) <= '1';
    layer1_outputs(89) <= layer0_outputs(2881);
    layer1_outputs(90) <= '1';
    layer1_outputs(91) <= layer0_outputs(1336);
    layer1_outputs(92) <= '1';
    layer1_outputs(93) <= '0';
    layer1_outputs(94) <= not(layer0_outputs(2868)) or (layer0_outputs(2006));
    layer1_outputs(95) <= '0';
    layer1_outputs(96) <= (layer0_outputs(1885)) and (layer0_outputs(3313));
    layer1_outputs(97) <= (layer0_outputs(1174)) and not (layer0_outputs(3979));
    layer1_outputs(98) <= (layer0_outputs(3216)) and not (layer0_outputs(1532));
    layer1_outputs(99) <= not(layer0_outputs(3884)) or (layer0_outputs(1695));
    layer1_outputs(100) <= (layer0_outputs(4496)) or (layer0_outputs(1923));
    layer1_outputs(101) <= '1';
    layer1_outputs(102) <= '1';
    layer1_outputs(103) <= '0';
    layer1_outputs(104) <= not((layer0_outputs(2510)) or (layer0_outputs(3402)));
    layer1_outputs(105) <= (layer0_outputs(2144)) and (layer0_outputs(2183));
    layer1_outputs(106) <= '0';
    layer1_outputs(107) <= not((layer0_outputs(2954)) or (layer0_outputs(4864)));
    layer1_outputs(108) <= (layer0_outputs(4977)) or (layer0_outputs(2404));
    layer1_outputs(109) <= layer0_outputs(453);
    layer1_outputs(110) <= layer0_outputs(4647);
    layer1_outputs(111) <= '1';
    layer1_outputs(112) <= (layer0_outputs(587)) and (layer0_outputs(2174));
    layer1_outputs(113) <= '1';
    layer1_outputs(114) <= (layer0_outputs(1880)) and (layer0_outputs(3900));
    layer1_outputs(115) <= '0';
    layer1_outputs(116) <= not(layer0_outputs(2273));
    layer1_outputs(117) <= (layer0_outputs(2723)) and not (layer0_outputs(4447));
    layer1_outputs(118) <= not((layer0_outputs(3240)) xor (layer0_outputs(1322)));
    layer1_outputs(119) <= (layer0_outputs(3653)) or (layer0_outputs(4141));
    layer1_outputs(120) <= not(layer0_outputs(3479));
    layer1_outputs(121) <= (layer0_outputs(3124)) and not (layer0_outputs(3599));
    layer1_outputs(122) <= '1';
    layer1_outputs(123) <= not((layer0_outputs(5033)) xor (layer0_outputs(4060)));
    layer1_outputs(124) <= (layer0_outputs(5022)) or (layer0_outputs(4720));
    layer1_outputs(125) <= (layer0_outputs(4395)) and not (layer0_outputs(4409));
    layer1_outputs(126) <= (layer0_outputs(3216)) and not (layer0_outputs(4901));
    layer1_outputs(127) <= (layer0_outputs(2807)) or (layer0_outputs(4597));
    layer1_outputs(128) <= not(layer0_outputs(5082)) or (layer0_outputs(524));
    layer1_outputs(129) <= layer0_outputs(2396);
    layer1_outputs(130) <= (layer0_outputs(1520)) and not (layer0_outputs(1261));
    layer1_outputs(131) <= not(layer0_outputs(677)) or (layer0_outputs(4722));
    layer1_outputs(132) <= not(layer0_outputs(1298)) or (layer0_outputs(2523));
    layer1_outputs(133) <= not(layer0_outputs(3072)) or (layer0_outputs(5067));
    layer1_outputs(134) <= '0';
    layer1_outputs(135) <= (layer0_outputs(2787)) or (layer0_outputs(1673));
    layer1_outputs(136) <= not(layer0_outputs(2021)) or (layer0_outputs(400));
    layer1_outputs(137) <= (layer0_outputs(3021)) and not (layer0_outputs(4129));
    layer1_outputs(138) <= not(layer0_outputs(1497));
    layer1_outputs(139) <= (layer0_outputs(1542)) and (layer0_outputs(155));
    layer1_outputs(140) <= (layer0_outputs(4726)) and not (layer0_outputs(724));
    layer1_outputs(141) <= '1';
    layer1_outputs(142) <= layer0_outputs(979);
    layer1_outputs(143) <= '1';
    layer1_outputs(144) <= '0';
    layer1_outputs(145) <= '1';
    layer1_outputs(146) <= (layer0_outputs(3836)) or (layer0_outputs(3902));
    layer1_outputs(147) <= layer0_outputs(3838);
    layer1_outputs(148) <= (layer0_outputs(3207)) or (layer0_outputs(5101));
    layer1_outputs(149) <= (layer0_outputs(3045)) and (layer0_outputs(3811));
    layer1_outputs(150) <= (layer0_outputs(4159)) and (layer0_outputs(1842));
    layer1_outputs(151) <= (layer0_outputs(4502)) and (layer0_outputs(1219));
    layer1_outputs(152) <= (layer0_outputs(188)) and not (layer0_outputs(1856));
    layer1_outputs(153) <= layer0_outputs(3622);
    layer1_outputs(154) <= not((layer0_outputs(780)) and (layer0_outputs(2804)));
    layer1_outputs(155) <= (layer0_outputs(4719)) or (layer0_outputs(4247));
    layer1_outputs(156) <= (layer0_outputs(4161)) or (layer0_outputs(296));
    layer1_outputs(157) <= not(layer0_outputs(3661));
    layer1_outputs(158) <= '1';
    layer1_outputs(159) <= layer0_outputs(1930);
    layer1_outputs(160) <= '1';
    layer1_outputs(161) <= (layer0_outputs(3104)) and not (layer0_outputs(2435));
    layer1_outputs(162) <= not(layer0_outputs(2788));
    layer1_outputs(163) <= not(layer0_outputs(2709));
    layer1_outputs(164) <= not(layer0_outputs(4324));
    layer1_outputs(165) <= '1';
    layer1_outputs(166) <= not((layer0_outputs(3445)) xor (layer0_outputs(2966)));
    layer1_outputs(167) <= not(layer0_outputs(1500)) or (layer0_outputs(1714));
    layer1_outputs(168) <= (layer0_outputs(2531)) and (layer0_outputs(3700));
    layer1_outputs(169) <= layer0_outputs(4520);
    layer1_outputs(170) <= layer0_outputs(1296);
    layer1_outputs(171) <= not(layer0_outputs(441));
    layer1_outputs(172) <= '1';
    layer1_outputs(173) <= '0';
    layer1_outputs(174) <= not(layer0_outputs(3218)) or (layer0_outputs(4916));
    layer1_outputs(175) <= not((layer0_outputs(470)) or (layer0_outputs(1247)));
    layer1_outputs(176) <= (layer0_outputs(4620)) and (layer0_outputs(4114));
    layer1_outputs(177) <= '0';
    layer1_outputs(178) <= not((layer0_outputs(1808)) and (layer0_outputs(2684)));
    layer1_outputs(179) <= '0';
    layer1_outputs(180) <= not(layer0_outputs(638));
    layer1_outputs(181) <= (layer0_outputs(4791)) and not (layer0_outputs(5053));
    layer1_outputs(182) <= not((layer0_outputs(4515)) and (layer0_outputs(3568)));
    layer1_outputs(183) <= layer0_outputs(1878);
    layer1_outputs(184) <= layer0_outputs(772);
    layer1_outputs(185) <= layer0_outputs(3415);
    layer1_outputs(186) <= not(layer0_outputs(3249));
    layer1_outputs(187) <= not(layer0_outputs(3651));
    layer1_outputs(188) <= layer0_outputs(2338);
    layer1_outputs(189) <= not(layer0_outputs(1282));
    layer1_outputs(190) <= not((layer0_outputs(2140)) xor (layer0_outputs(5028)));
    layer1_outputs(191) <= (layer0_outputs(2288)) or (layer0_outputs(3048));
    layer1_outputs(192) <= '1';
    layer1_outputs(193) <= '0';
    layer1_outputs(194) <= '0';
    layer1_outputs(195) <= '0';
    layer1_outputs(196) <= layer0_outputs(2106);
    layer1_outputs(197) <= (layer0_outputs(1012)) and not (layer0_outputs(2524));
    layer1_outputs(198) <= '1';
    layer1_outputs(199) <= '0';
    layer1_outputs(200) <= not(layer0_outputs(2213));
    layer1_outputs(201) <= not(layer0_outputs(402));
    layer1_outputs(202) <= not(layer0_outputs(1868)) or (layer0_outputs(2855));
    layer1_outputs(203) <= '0';
    layer1_outputs(204) <= not((layer0_outputs(2143)) or (layer0_outputs(236)));
    layer1_outputs(205) <= (layer0_outputs(5065)) and not (layer0_outputs(1970));
    layer1_outputs(206) <= not(layer0_outputs(2271)) or (layer0_outputs(3346));
    layer1_outputs(207) <= layer0_outputs(673);
    layer1_outputs(208) <= '1';
    layer1_outputs(209) <= not((layer0_outputs(2071)) xor (layer0_outputs(1679)));
    layer1_outputs(210) <= layer0_outputs(1022);
    layer1_outputs(211) <= (layer0_outputs(4926)) or (layer0_outputs(3603));
    layer1_outputs(212) <= not((layer0_outputs(2843)) or (layer0_outputs(1915)));
    layer1_outputs(213) <= not((layer0_outputs(3453)) xor (layer0_outputs(76)));
    layer1_outputs(214) <= (layer0_outputs(682)) and (layer0_outputs(450));
    layer1_outputs(215) <= not(layer0_outputs(937)) or (layer0_outputs(1656));
    layer1_outputs(216) <= (layer0_outputs(4669)) or (layer0_outputs(4331));
    layer1_outputs(217) <= not(layer0_outputs(3823)) or (layer0_outputs(1402));
    layer1_outputs(218) <= layer0_outputs(4293);
    layer1_outputs(219) <= '0';
    layer1_outputs(220) <= not(layer0_outputs(5032)) or (layer0_outputs(2581));
    layer1_outputs(221) <= (layer0_outputs(373)) and not (layer0_outputs(2541));
    layer1_outputs(222) <= '0';
    layer1_outputs(223) <= (layer0_outputs(1880)) and not (layer0_outputs(1107));
    layer1_outputs(224) <= layer0_outputs(2946);
    layer1_outputs(225) <= not(layer0_outputs(4566)) or (layer0_outputs(2757));
    layer1_outputs(226) <= (layer0_outputs(283)) or (layer0_outputs(4312));
    layer1_outputs(227) <= '0';
    layer1_outputs(228) <= not(layer0_outputs(527)) or (layer0_outputs(3027));
    layer1_outputs(229) <= not((layer0_outputs(4051)) and (layer0_outputs(2732)));
    layer1_outputs(230) <= (layer0_outputs(2253)) and (layer0_outputs(1706));
    layer1_outputs(231) <= not(layer0_outputs(2472));
    layer1_outputs(232) <= '1';
    layer1_outputs(233) <= not((layer0_outputs(1782)) and (layer0_outputs(2607)));
    layer1_outputs(234) <= not(layer0_outputs(3289));
    layer1_outputs(235) <= '1';
    layer1_outputs(236) <= '1';
    layer1_outputs(237) <= (layer0_outputs(492)) and not (layer0_outputs(4219));
    layer1_outputs(238) <= (layer0_outputs(2694)) and not (layer0_outputs(338));
    layer1_outputs(239) <= not(layer0_outputs(4423)) or (layer0_outputs(4750));
    layer1_outputs(240) <= not((layer0_outputs(588)) or (layer0_outputs(2126)));
    layer1_outputs(241) <= not(layer0_outputs(991)) or (layer0_outputs(3301));
    layer1_outputs(242) <= '1';
    layer1_outputs(243) <= not(layer0_outputs(4471));
    layer1_outputs(244) <= (layer0_outputs(2466)) and (layer0_outputs(2005));
    layer1_outputs(245) <= not((layer0_outputs(3783)) and (layer0_outputs(3858)));
    layer1_outputs(246) <= '1';
    layer1_outputs(247) <= '1';
    layer1_outputs(248) <= not(layer0_outputs(3316));
    layer1_outputs(249) <= (layer0_outputs(2328)) and (layer0_outputs(3841));
    layer1_outputs(250) <= '1';
    layer1_outputs(251) <= not(layer0_outputs(3039)) or (layer0_outputs(1296));
    layer1_outputs(252) <= not(layer0_outputs(4233));
    layer1_outputs(253) <= layer0_outputs(357);
    layer1_outputs(254) <= '0';
    layer1_outputs(255) <= not((layer0_outputs(381)) and (layer0_outputs(1332)));
    layer1_outputs(256) <= not(layer0_outputs(4059));
    layer1_outputs(257) <= not(layer0_outputs(1754));
    layer1_outputs(258) <= not(layer0_outputs(2300));
    layer1_outputs(259) <= not(layer0_outputs(4387));
    layer1_outputs(260) <= '1';
    layer1_outputs(261) <= (layer0_outputs(544)) and not (layer0_outputs(4033));
    layer1_outputs(262) <= '1';
    layer1_outputs(263) <= layer0_outputs(603);
    layer1_outputs(264) <= (layer0_outputs(461)) or (layer0_outputs(3814));
    layer1_outputs(265) <= (layer0_outputs(4295)) and not (layer0_outputs(3646));
    layer1_outputs(266) <= not((layer0_outputs(1429)) or (layer0_outputs(960)));
    layer1_outputs(267) <= (layer0_outputs(996)) and not (layer0_outputs(3156));
    layer1_outputs(268) <= '0';
    layer1_outputs(269) <= '1';
    layer1_outputs(270) <= not(layer0_outputs(5011));
    layer1_outputs(271) <= not(layer0_outputs(988));
    layer1_outputs(272) <= (layer0_outputs(4830)) or (layer0_outputs(2156));
    layer1_outputs(273) <= (layer0_outputs(4484)) and not (layer0_outputs(1632));
    layer1_outputs(274) <= '1';
    layer1_outputs(275) <= (layer0_outputs(2684)) or (layer0_outputs(1259));
    layer1_outputs(276) <= not((layer0_outputs(55)) or (layer0_outputs(160)));
    layer1_outputs(277) <= not(layer0_outputs(4346));
    layer1_outputs(278) <= '1';
    layer1_outputs(279) <= layer0_outputs(3651);
    layer1_outputs(280) <= not(layer0_outputs(1726)) or (layer0_outputs(3211));
    layer1_outputs(281) <= '0';
    layer1_outputs(282) <= '1';
    layer1_outputs(283) <= layer0_outputs(4462);
    layer1_outputs(284) <= (layer0_outputs(2970)) and not (layer0_outputs(4000));
    layer1_outputs(285) <= (layer0_outputs(2977)) and not (layer0_outputs(4683));
    layer1_outputs(286) <= not((layer0_outputs(1006)) and (layer0_outputs(2642)));
    layer1_outputs(287) <= layer0_outputs(3318);
    layer1_outputs(288) <= layer0_outputs(3857);
    layer1_outputs(289) <= not((layer0_outputs(3011)) and (layer0_outputs(3118)));
    layer1_outputs(290) <= not(layer0_outputs(1718)) or (layer0_outputs(1552));
    layer1_outputs(291) <= (layer0_outputs(5020)) and (layer0_outputs(4216));
    layer1_outputs(292) <= '1';
    layer1_outputs(293) <= not(layer0_outputs(152));
    layer1_outputs(294) <= '0';
    layer1_outputs(295) <= '1';
    layer1_outputs(296) <= '0';
    layer1_outputs(297) <= not(layer0_outputs(118)) or (layer0_outputs(1856));
    layer1_outputs(298) <= layer0_outputs(483);
    layer1_outputs(299) <= not(layer0_outputs(1180)) or (layer0_outputs(3644));
    layer1_outputs(300) <= not(layer0_outputs(2349));
    layer1_outputs(301) <= '0';
    layer1_outputs(302) <= (layer0_outputs(604)) or (layer0_outputs(4142));
    layer1_outputs(303) <= '0';
    layer1_outputs(304) <= not(layer0_outputs(4675));
    layer1_outputs(305) <= not(layer0_outputs(85)) or (layer0_outputs(1977));
    layer1_outputs(306) <= not(layer0_outputs(4942));
    layer1_outputs(307) <= not(layer0_outputs(189));
    layer1_outputs(308) <= not((layer0_outputs(2969)) and (layer0_outputs(4481)));
    layer1_outputs(309) <= (layer0_outputs(206)) and not (layer0_outputs(1369));
    layer1_outputs(310) <= (layer0_outputs(3079)) and not (layer0_outputs(3178));
    layer1_outputs(311) <= (layer0_outputs(611)) and not (layer0_outputs(754));
    layer1_outputs(312) <= not(layer0_outputs(4355));
    layer1_outputs(313) <= not((layer0_outputs(2946)) xor (layer0_outputs(15)));
    layer1_outputs(314) <= (layer0_outputs(4906)) and (layer0_outputs(2182));
    layer1_outputs(315) <= not(layer0_outputs(3194)) or (layer0_outputs(3638));
    layer1_outputs(316) <= not(layer0_outputs(2493)) or (layer0_outputs(1483));
    layer1_outputs(317) <= (layer0_outputs(1705)) and not (layer0_outputs(4957));
    layer1_outputs(318) <= (layer0_outputs(3447)) or (layer0_outputs(112));
    layer1_outputs(319) <= (layer0_outputs(500)) and not (layer0_outputs(4527));
    layer1_outputs(320) <= '1';
    layer1_outputs(321) <= '0';
    layer1_outputs(322) <= '1';
    layer1_outputs(323) <= (layer0_outputs(2084)) and not (layer0_outputs(1355));
    layer1_outputs(324) <= (layer0_outputs(838)) and not (layer0_outputs(629));
    layer1_outputs(325) <= layer0_outputs(1234);
    layer1_outputs(326) <= not(layer0_outputs(1982));
    layer1_outputs(327) <= layer0_outputs(1674);
    layer1_outputs(328) <= (layer0_outputs(1583)) and not (layer0_outputs(1761));
    layer1_outputs(329) <= not(layer0_outputs(1957));
    layer1_outputs(330) <= '1';
    layer1_outputs(331) <= layer0_outputs(3899);
    layer1_outputs(332) <= (layer0_outputs(1111)) and not (layer0_outputs(586));
    layer1_outputs(333) <= not(layer0_outputs(3960)) or (layer0_outputs(1439));
    layer1_outputs(334) <= (layer0_outputs(2564)) and not (layer0_outputs(344));
    layer1_outputs(335) <= '0';
    layer1_outputs(336) <= '0';
    layer1_outputs(337) <= not(layer0_outputs(1085)) or (layer0_outputs(3039));
    layer1_outputs(338) <= layer0_outputs(2246);
    layer1_outputs(339) <= (layer0_outputs(326)) or (layer0_outputs(5095));
    layer1_outputs(340) <= (layer0_outputs(189)) or (layer0_outputs(1960));
    layer1_outputs(341) <= not(layer0_outputs(1877));
    layer1_outputs(342) <= (layer0_outputs(2222)) or (layer0_outputs(1894));
    layer1_outputs(343) <= layer0_outputs(2256);
    layer1_outputs(344) <= '0';
    layer1_outputs(345) <= not((layer0_outputs(3784)) or (layer0_outputs(2207)));
    layer1_outputs(346) <= not(layer0_outputs(4959));
    layer1_outputs(347) <= '1';
    layer1_outputs(348) <= not(layer0_outputs(1780)) or (layer0_outputs(3594));
    layer1_outputs(349) <= (layer0_outputs(3034)) and not (layer0_outputs(2244));
    layer1_outputs(350) <= '0';
    layer1_outputs(351) <= '1';
    layer1_outputs(352) <= layer0_outputs(3716);
    layer1_outputs(353) <= (layer0_outputs(2422)) and not (layer0_outputs(4406));
    layer1_outputs(354) <= not((layer0_outputs(3296)) or (layer0_outputs(4520)));
    layer1_outputs(355) <= '0';
    layer1_outputs(356) <= '0';
    layer1_outputs(357) <= not((layer0_outputs(192)) and (layer0_outputs(4111)));
    layer1_outputs(358) <= not(layer0_outputs(2472));
    layer1_outputs(359) <= not(layer0_outputs(4959)) or (layer0_outputs(4843));
    layer1_outputs(360) <= not((layer0_outputs(1250)) or (layer0_outputs(1695)));
    layer1_outputs(361) <= '1';
    layer1_outputs(362) <= '0';
    layer1_outputs(363) <= not((layer0_outputs(96)) and (layer0_outputs(4532)));
    layer1_outputs(364) <= not(layer0_outputs(825)) or (layer0_outputs(3434));
    layer1_outputs(365) <= not(layer0_outputs(649));
    layer1_outputs(366) <= layer0_outputs(2710);
    layer1_outputs(367) <= not((layer0_outputs(4319)) or (layer0_outputs(2306)));
    layer1_outputs(368) <= '1';
    layer1_outputs(369) <= layer0_outputs(3909);
    layer1_outputs(370) <= not(layer0_outputs(458)) or (layer0_outputs(115));
    layer1_outputs(371) <= not(layer0_outputs(4063));
    layer1_outputs(372) <= (layer0_outputs(228)) and not (layer0_outputs(3449));
    layer1_outputs(373) <= not(layer0_outputs(2387));
    layer1_outputs(374) <= not((layer0_outputs(523)) xor (layer0_outputs(2761)));
    layer1_outputs(375) <= '1';
    layer1_outputs(376) <= (layer0_outputs(1949)) and not (layer0_outputs(2949));
    layer1_outputs(377) <= not((layer0_outputs(2301)) or (layer0_outputs(736)));
    layer1_outputs(378) <= (layer0_outputs(3513)) and (layer0_outputs(5111));
    layer1_outputs(379) <= not(layer0_outputs(751)) or (layer0_outputs(4209));
    layer1_outputs(380) <= not((layer0_outputs(2010)) or (layer0_outputs(3513)));
    layer1_outputs(381) <= (layer0_outputs(4354)) or (layer0_outputs(1201));
    layer1_outputs(382) <= not(layer0_outputs(1036)) or (layer0_outputs(2887));
    layer1_outputs(383) <= not((layer0_outputs(2769)) or (layer0_outputs(3880)));
    layer1_outputs(384) <= layer0_outputs(1655);
    layer1_outputs(385) <= not(layer0_outputs(2750)) or (layer0_outputs(1587));
    layer1_outputs(386) <= (layer0_outputs(2749)) xor (layer0_outputs(2976));
    layer1_outputs(387) <= not(layer0_outputs(1062));
    layer1_outputs(388) <= '0';
    layer1_outputs(389) <= not(layer0_outputs(4418)) or (layer0_outputs(277));
    layer1_outputs(390) <= not((layer0_outputs(4560)) or (layer0_outputs(4)));
    layer1_outputs(391) <= (layer0_outputs(1739)) and not (layer0_outputs(3838));
    layer1_outputs(392) <= (layer0_outputs(2129)) xor (layer0_outputs(203));
    layer1_outputs(393) <= (layer0_outputs(3219)) and not (layer0_outputs(1099));
    layer1_outputs(394) <= '1';
    layer1_outputs(395) <= '1';
    layer1_outputs(396) <= not((layer0_outputs(3707)) or (layer0_outputs(519)));
    layer1_outputs(397) <= (layer0_outputs(2570)) or (layer0_outputs(4125));
    layer1_outputs(398) <= not(layer0_outputs(969));
    layer1_outputs(399) <= not(layer0_outputs(321));
    layer1_outputs(400) <= not(layer0_outputs(3201));
    layer1_outputs(401) <= not((layer0_outputs(4191)) or (layer0_outputs(1998)));
    layer1_outputs(402) <= (layer0_outputs(3159)) and (layer0_outputs(1806));
    layer1_outputs(403) <= layer0_outputs(916);
    layer1_outputs(404) <= (layer0_outputs(719)) and (layer0_outputs(2834));
    layer1_outputs(405) <= (layer0_outputs(4227)) and (layer0_outputs(1082));
    layer1_outputs(406) <= not(layer0_outputs(1665)) or (layer0_outputs(3665));
    layer1_outputs(407) <= '1';
    layer1_outputs(408) <= not((layer0_outputs(3660)) and (layer0_outputs(656)));
    layer1_outputs(409) <= (layer0_outputs(3027)) and not (layer0_outputs(2503));
    layer1_outputs(410) <= (layer0_outputs(5104)) or (layer0_outputs(2549));
    layer1_outputs(411) <= layer0_outputs(3167);
    layer1_outputs(412) <= not(layer0_outputs(2517)) or (layer0_outputs(3967));
    layer1_outputs(413) <= not(layer0_outputs(1937));
    layer1_outputs(414) <= not((layer0_outputs(2431)) and (layer0_outputs(2725)));
    layer1_outputs(415) <= (layer0_outputs(3666)) and not (layer0_outputs(4144));
    layer1_outputs(416) <= not(layer0_outputs(4378)) or (layer0_outputs(883));
    layer1_outputs(417) <= '1';
    layer1_outputs(418) <= '0';
    layer1_outputs(419) <= not((layer0_outputs(1182)) xor (layer0_outputs(548)));
    layer1_outputs(420) <= not((layer0_outputs(983)) or (layer0_outputs(4250)));
    layer1_outputs(421) <= '0';
    layer1_outputs(422) <= (layer0_outputs(3553)) xor (layer0_outputs(1145));
    layer1_outputs(423) <= layer0_outputs(1475);
    layer1_outputs(424) <= '1';
    layer1_outputs(425) <= not(layer0_outputs(217));
    layer1_outputs(426) <= (layer0_outputs(577)) or (layer0_outputs(2869));
    layer1_outputs(427) <= (layer0_outputs(4407)) or (layer0_outputs(2707));
    layer1_outputs(428) <= layer0_outputs(2889);
    layer1_outputs(429) <= layer0_outputs(4766);
    layer1_outputs(430) <= not(layer0_outputs(4798));
    layer1_outputs(431) <= not((layer0_outputs(993)) or (layer0_outputs(2373)));
    layer1_outputs(432) <= (layer0_outputs(2793)) and not (layer0_outputs(768));
    layer1_outputs(433) <= '1';
    layer1_outputs(434) <= '0';
    layer1_outputs(435) <= (layer0_outputs(4389)) and (layer0_outputs(1484));
    layer1_outputs(436) <= not(layer0_outputs(2547)) or (layer0_outputs(2847));
    layer1_outputs(437) <= not(layer0_outputs(3550));
    layer1_outputs(438) <= layer0_outputs(741);
    layer1_outputs(439) <= (layer0_outputs(1011)) and not (layer0_outputs(4170));
    layer1_outputs(440) <= not(layer0_outputs(2656)) or (layer0_outputs(2623));
    layer1_outputs(441) <= (layer0_outputs(231)) and (layer0_outputs(4771));
    layer1_outputs(442) <= layer0_outputs(5050);
    layer1_outputs(443) <= '1';
    layer1_outputs(444) <= layer0_outputs(3655);
    layer1_outputs(445) <= not(layer0_outputs(1463));
    layer1_outputs(446) <= '0';
    layer1_outputs(447) <= (layer0_outputs(4806)) and not (layer0_outputs(726));
    layer1_outputs(448) <= not(layer0_outputs(673));
    layer1_outputs(449) <= (layer0_outputs(590)) and not (layer0_outputs(4539));
    layer1_outputs(450) <= '0';
    layer1_outputs(451) <= not((layer0_outputs(3153)) xor (layer0_outputs(5098)));
    layer1_outputs(452) <= not(layer0_outputs(4963));
    layer1_outputs(453) <= '0';
    layer1_outputs(454) <= (layer0_outputs(1476)) and (layer0_outputs(1267));
    layer1_outputs(455) <= '1';
    layer1_outputs(456) <= (layer0_outputs(3315)) and (layer0_outputs(102));
    layer1_outputs(457) <= '1';
    layer1_outputs(458) <= not(layer0_outputs(4341)) or (layer0_outputs(1631));
    layer1_outputs(459) <= not(layer0_outputs(100));
    layer1_outputs(460) <= not(layer0_outputs(4763)) or (layer0_outputs(1652));
    layer1_outputs(461) <= (layer0_outputs(884)) and (layer0_outputs(2255));
    layer1_outputs(462) <= (layer0_outputs(4658)) and not (layer0_outputs(1947));
    layer1_outputs(463) <= not(layer0_outputs(4828)) or (layer0_outputs(3804));
    layer1_outputs(464) <= not((layer0_outputs(2460)) xor (layer0_outputs(348)));
    layer1_outputs(465) <= '1';
    layer1_outputs(466) <= not(layer0_outputs(2632));
    layer1_outputs(467) <= (layer0_outputs(2888)) and not (layer0_outputs(127));
    layer1_outputs(468) <= not((layer0_outputs(3318)) and (layer0_outputs(2738)));
    layer1_outputs(469) <= (layer0_outputs(3050)) and not (layer0_outputs(4199));
    layer1_outputs(470) <= not(layer0_outputs(2633)) or (layer0_outputs(3514));
    layer1_outputs(471) <= not((layer0_outputs(4841)) xor (layer0_outputs(5060)));
    layer1_outputs(472) <= '1';
    layer1_outputs(473) <= (layer0_outputs(1671)) and not (layer0_outputs(2426));
    layer1_outputs(474) <= (layer0_outputs(196)) and not (layer0_outputs(3915));
    layer1_outputs(475) <= (layer0_outputs(135)) and (layer0_outputs(89));
    layer1_outputs(476) <= not((layer0_outputs(4473)) or (layer0_outputs(1745)));
    layer1_outputs(477) <= not(layer0_outputs(1900));
    layer1_outputs(478) <= '0';
    layer1_outputs(479) <= not((layer0_outputs(3582)) and (layer0_outputs(2674)));
    layer1_outputs(480) <= '1';
    layer1_outputs(481) <= not(layer0_outputs(1742));
    layer1_outputs(482) <= '0';
    layer1_outputs(483) <= (layer0_outputs(685)) or (layer0_outputs(4135));
    layer1_outputs(484) <= layer0_outputs(1252);
    layer1_outputs(485) <= not(layer0_outputs(4716)) or (layer0_outputs(845));
    layer1_outputs(486) <= layer0_outputs(1438);
    layer1_outputs(487) <= '1';
    layer1_outputs(488) <= not(layer0_outputs(1738)) or (layer0_outputs(1194));
    layer1_outputs(489) <= '1';
    layer1_outputs(490) <= not(layer0_outputs(3903));
    layer1_outputs(491) <= not(layer0_outputs(4321));
    layer1_outputs(492) <= '0';
    layer1_outputs(493) <= not((layer0_outputs(2418)) and (layer0_outputs(1203)));
    layer1_outputs(494) <= layer0_outputs(3705);
    layer1_outputs(495) <= not(layer0_outputs(3165)) or (layer0_outputs(1978));
    layer1_outputs(496) <= (layer0_outputs(3054)) xor (layer0_outputs(2528));
    layer1_outputs(497) <= '1';
    layer1_outputs(498) <= '1';
    layer1_outputs(499) <= not(layer0_outputs(2342));
    layer1_outputs(500) <= (layer0_outputs(4241)) and not (layer0_outputs(1818));
    layer1_outputs(501) <= not(layer0_outputs(81));
    layer1_outputs(502) <= (layer0_outputs(3376)) and not (layer0_outputs(3614));
    layer1_outputs(503) <= layer0_outputs(3403);
    layer1_outputs(504) <= not(layer0_outputs(3422)) or (layer0_outputs(3280));
    layer1_outputs(505) <= not(layer0_outputs(2760)) or (layer0_outputs(2269));
    layer1_outputs(506) <= not(layer0_outputs(4158)) or (layer0_outputs(1435));
    layer1_outputs(507) <= not(layer0_outputs(4713));
    layer1_outputs(508) <= '0';
    layer1_outputs(509) <= (layer0_outputs(1649)) and not (layer0_outputs(2914));
    layer1_outputs(510) <= '0';
    layer1_outputs(511) <= layer0_outputs(407);
    layer1_outputs(512) <= (layer0_outputs(2536)) and (layer0_outputs(4272));
    layer1_outputs(513) <= '0';
    layer1_outputs(514) <= (layer0_outputs(1316)) and not (layer0_outputs(1072));
    layer1_outputs(515) <= not(layer0_outputs(3572)) or (layer0_outputs(124));
    layer1_outputs(516) <= not(layer0_outputs(148)) or (layer0_outputs(3285));
    layer1_outputs(517) <= '1';
    layer1_outputs(518) <= (layer0_outputs(4328)) and not (layer0_outputs(2186));
    layer1_outputs(519) <= (layer0_outputs(2332)) and not (layer0_outputs(1229));
    layer1_outputs(520) <= not((layer0_outputs(4220)) or (layer0_outputs(4462)));
    layer1_outputs(521) <= '0';
    layer1_outputs(522) <= '0';
    layer1_outputs(523) <= (layer0_outputs(2319)) and not (layer0_outputs(632));
    layer1_outputs(524) <= not(layer0_outputs(991)) or (layer0_outputs(4276));
    layer1_outputs(525) <= (layer0_outputs(3503)) and not (layer0_outputs(3060));
    layer1_outputs(526) <= (layer0_outputs(4269)) and not (layer0_outputs(4234));
    layer1_outputs(527) <= not(layer0_outputs(1493)) or (layer0_outputs(2416));
    layer1_outputs(528) <= (layer0_outputs(4412)) and not (layer0_outputs(924));
    layer1_outputs(529) <= (layer0_outputs(140)) and not (layer0_outputs(3958));
    layer1_outputs(530) <= layer0_outputs(462);
    layer1_outputs(531) <= not((layer0_outputs(445)) or (layer0_outputs(2198)));
    layer1_outputs(532) <= '1';
    layer1_outputs(533) <= layer0_outputs(4793);
    layer1_outputs(534) <= not((layer0_outputs(494)) and (layer0_outputs(414)));
    layer1_outputs(535) <= not((layer0_outputs(416)) or (layer0_outputs(5074)));
    layer1_outputs(536) <= not((layer0_outputs(1359)) or (layer0_outputs(1539)));
    layer1_outputs(537) <= layer0_outputs(615);
    layer1_outputs(538) <= (layer0_outputs(2613)) and not (layer0_outputs(1639));
    layer1_outputs(539) <= '0';
    layer1_outputs(540) <= (layer0_outputs(3064)) xor (layer0_outputs(3654));
    layer1_outputs(541) <= not((layer0_outputs(1468)) and (layer0_outputs(4619)));
    layer1_outputs(542) <= '1';
    layer1_outputs(543) <= (layer0_outputs(1890)) xor (layer0_outputs(784));
    layer1_outputs(544) <= layer0_outputs(343);
    layer1_outputs(545) <= layer0_outputs(4699);
    layer1_outputs(546) <= (layer0_outputs(11)) and (layer0_outputs(3176));
    layer1_outputs(547) <= '1';
    layer1_outputs(548) <= (layer0_outputs(233)) or (layer0_outputs(2557));
    layer1_outputs(549) <= (layer0_outputs(3676)) and (layer0_outputs(2471));
    layer1_outputs(550) <= '0';
    layer1_outputs(551) <= '1';
    layer1_outputs(552) <= (layer0_outputs(1412)) or (layer0_outputs(2035));
    layer1_outputs(553) <= not((layer0_outputs(4787)) and (layer0_outputs(4301)));
    layer1_outputs(554) <= layer0_outputs(3875);
    layer1_outputs(555) <= not((layer0_outputs(2500)) and (layer0_outputs(4491)));
    layer1_outputs(556) <= '0';
    layer1_outputs(557) <= not((layer0_outputs(2838)) and (layer0_outputs(381)));
    layer1_outputs(558) <= (layer0_outputs(848)) and not (layer0_outputs(120));
    layer1_outputs(559) <= layer0_outputs(4697);
    layer1_outputs(560) <= '1';
    layer1_outputs(561) <= layer0_outputs(171);
    layer1_outputs(562) <= '1';
    layer1_outputs(563) <= not(layer0_outputs(4097));
    layer1_outputs(564) <= (layer0_outputs(3268)) and not (layer0_outputs(4396));
    layer1_outputs(565) <= '0';
    layer1_outputs(566) <= (layer0_outputs(1258)) or (layer0_outputs(429));
    layer1_outputs(567) <= (layer0_outputs(3811)) and not (layer0_outputs(3126));
    layer1_outputs(568) <= (layer0_outputs(3396)) and not (layer0_outputs(1368));
    layer1_outputs(569) <= (layer0_outputs(602)) and (layer0_outputs(3725));
    layer1_outputs(570) <= layer0_outputs(1699);
    layer1_outputs(571) <= not((layer0_outputs(2013)) or (layer0_outputs(1812)));
    layer1_outputs(572) <= not((layer0_outputs(727)) and (layer0_outputs(122)));
    layer1_outputs(573) <= '0';
    layer1_outputs(574) <= not(layer0_outputs(1070)) or (layer0_outputs(3477));
    layer1_outputs(575) <= (layer0_outputs(4684)) and not (layer0_outputs(3993));
    layer1_outputs(576) <= not((layer0_outputs(215)) and (layer0_outputs(3612)));
    layer1_outputs(577) <= not(layer0_outputs(2756)) or (layer0_outputs(3122));
    layer1_outputs(578) <= not(layer0_outputs(1850)) or (layer0_outputs(4966));
    layer1_outputs(579) <= not(layer0_outputs(1253));
    layer1_outputs(580) <= (layer0_outputs(179)) and not (layer0_outputs(4182));
    layer1_outputs(581) <= '1';
    layer1_outputs(582) <= '0';
    layer1_outputs(583) <= not(layer0_outputs(5036)) or (layer0_outputs(4280));
    layer1_outputs(584) <= not(layer0_outputs(607));
    layer1_outputs(585) <= (layer0_outputs(3941)) or (layer0_outputs(3738));
    layer1_outputs(586) <= (layer0_outputs(4268)) and not (layer0_outputs(926));
    layer1_outputs(587) <= not(layer0_outputs(2629)) or (layer0_outputs(2082));
    layer1_outputs(588) <= layer0_outputs(3259);
    layer1_outputs(589) <= '1';
    layer1_outputs(590) <= layer0_outputs(546);
    layer1_outputs(591) <= (layer0_outputs(4627)) and not (layer0_outputs(2014));
    layer1_outputs(592) <= '0';
    layer1_outputs(593) <= (layer0_outputs(5109)) and not (layer0_outputs(420));
    layer1_outputs(594) <= layer0_outputs(3714);
    layer1_outputs(595) <= (layer0_outputs(228)) and (layer0_outputs(1052));
    layer1_outputs(596) <= not((layer0_outputs(273)) and (layer0_outputs(4724)));
    layer1_outputs(597) <= not(layer0_outputs(623));
    layer1_outputs(598) <= (layer0_outputs(1738)) and (layer0_outputs(3576));
    layer1_outputs(599) <= not(layer0_outputs(4136)) or (layer0_outputs(737));
    layer1_outputs(600) <= (layer0_outputs(256)) and not (layer0_outputs(769));
    layer1_outputs(601) <= not((layer0_outputs(2841)) or (layer0_outputs(4067)));
    layer1_outputs(602) <= '1';
    layer1_outputs(603) <= layer0_outputs(2935);
    layer1_outputs(604) <= (layer0_outputs(1904)) or (layer0_outputs(2745));
    layer1_outputs(605) <= '1';
    layer1_outputs(606) <= not(layer0_outputs(1251));
    layer1_outputs(607) <= not(layer0_outputs(4423)) or (layer0_outputs(1609));
    layer1_outputs(608) <= (layer0_outputs(2251)) and (layer0_outputs(1704));
    layer1_outputs(609) <= (layer0_outputs(2603)) and not (layer0_outputs(198));
    layer1_outputs(610) <= not(layer0_outputs(4178));
    layer1_outputs(611) <= layer0_outputs(4443);
    layer1_outputs(612) <= not(layer0_outputs(172)) or (layer0_outputs(111));
    layer1_outputs(613) <= (layer0_outputs(4971)) and not (layer0_outputs(4733));
    layer1_outputs(614) <= '1';
    layer1_outputs(615) <= not(layer0_outputs(1715));
    layer1_outputs(616) <= not((layer0_outputs(3737)) or (layer0_outputs(3168)));
    layer1_outputs(617) <= '0';
    layer1_outputs(618) <= not(layer0_outputs(1836)) or (layer0_outputs(4855));
    layer1_outputs(619) <= not(layer0_outputs(684)) or (layer0_outputs(4404));
    layer1_outputs(620) <= (layer0_outputs(3920)) and not (layer0_outputs(3347));
    layer1_outputs(621) <= not((layer0_outputs(525)) or (layer0_outputs(2138)));
    layer1_outputs(622) <= not((layer0_outputs(2201)) or (layer0_outputs(1051)));
    layer1_outputs(623) <= (layer0_outputs(2127)) and not (layer0_outputs(4603));
    layer1_outputs(624) <= '0';
    layer1_outputs(625) <= not(layer0_outputs(2937));
    layer1_outputs(626) <= (layer0_outputs(551)) and (layer0_outputs(2849));
    layer1_outputs(627) <= not(layer0_outputs(1244));
    layer1_outputs(628) <= not(layer0_outputs(416)) or (layer0_outputs(3985));
    layer1_outputs(629) <= (layer0_outputs(339)) and (layer0_outputs(779));
    layer1_outputs(630) <= (layer0_outputs(1857)) or (layer0_outputs(442));
    layer1_outputs(631) <= (layer0_outputs(3846)) and (layer0_outputs(651));
    layer1_outputs(632) <= not(layer0_outputs(1125));
    layer1_outputs(633) <= '0';
    layer1_outputs(634) <= (layer0_outputs(2973)) or (layer0_outputs(1876));
    layer1_outputs(635) <= (layer0_outputs(4441)) and not (layer0_outputs(3701));
    layer1_outputs(636) <= not(layer0_outputs(3969));
    layer1_outputs(637) <= '0';
    layer1_outputs(638) <= not(layer0_outputs(3720));
    layer1_outputs(639) <= not((layer0_outputs(3797)) and (layer0_outputs(962)));
    layer1_outputs(640) <= '0';
    layer1_outputs(641) <= '0';
    layer1_outputs(642) <= (layer0_outputs(4854)) and not (layer0_outputs(2262));
    layer1_outputs(643) <= (layer0_outputs(3275)) and (layer0_outputs(506));
    layer1_outputs(644) <= not((layer0_outputs(2341)) or (layer0_outputs(2056)));
    layer1_outputs(645) <= not((layer0_outputs(129)) or (layer0_outputs(2514)));
    layer1_outputs(646) <= layer0_outputs(2713);
    layer1_outputs(647) <= '0';
    layer1_outputs(648) <= '1';
    layer1_outputs(649) <= '1';
    layer1_outputs(650) <= layer0_outputs(4830);
    layer1_outputs(651) <= not(layer0_outputs(2596)) or (layer0_outputs(300));
    layer1_outputs(652) <= (layer0_outputs(2913)) and not (layer0_outputs(3117));
    layer1_outputs(653) <= layer0_outputs(3380);
    layer1_outputs(654) <= not(layer0_outputs(2346));
    layer1_outputs(655) <= not((layer0_outputs(856)) and (layer0_outputs(4126)));
    layer1_outputs(656) <= not(layer0_outputs(5035));
    layer1_outputs(657) <= '0';
    layer1_outputs(658) <= layer0_outputs(3271);
    layer1_outputs(659) <= not(layer0_outputs(3663)) or (layer0_outputs(3648));
    layer1_outputs(660) <= '0';
    layer1_outputs(661) <= '1';
    layer1_outputs(662) <= (layer0_outputs(4797)) or (layer0_outputs(4203));
    layer1_outputs(663) <= (layer0_outputs(1089)) and (layer0_outputs(3798));
    layer1_outputs(664) <= not((layer0_outputs(662)) and (layer0_outputs(4574)));
    layer1_outputs(665) <= '0';
    layer1_outputs(666) <= not((layer0_outputs(2815)) and (layer0_outputs(1073)));
    layer1_outputs(667) <= not(layer0_outputs(1232)) or (layer0_outputs(4414));
    layer1_outputs(668) <= '0';
    layer1_outputs(669) <= not(layer0_outputs(4583)) or (layer0_outputs(570));
    layer1_outputs(670) <= '0';
    layer1_outputs(671) <= not((layer0_outputs(4662)) and (layer0_outputs(724)));
    layer1_outputs(672) <= layer0_outputs(1680);
    layer1_outputs(673) <= not(layer0_outputs(1821));
    layer1_outputs(674) <= not((layer0_outputs(4789)) and (layer0_outputs(3197)));
    layer1_outputs(675) <= layer0_outputs(4988);
    layer1_outputs(676) <= '1';
    layer1_outputs(677) <= '1';
    layer1_outputs(678) <= not((layer0_outputs(4223)) or (layer0_outputs(75)));
    layer1_outputs(679) <= '0';
    layer1_outputs(680) <= not(layer0_outputs(892));
    layer1_outputs(681) <= '1';
    layer1_outputs(682) <= (layer0_outputs(5011)) and not (layer0_outputs(2504));
    layer1_outputs(683) <= not(layer0_outputs(3813)) or (layer0_outputs(4626));
    layer1_outputs(684) <= (layer0_outputs(3239)) and not (layer0_outputs(713));
    layer1_outputs(685) <= not(layer0_outputs(2709));
    layer1_outputs(686) <= (layer0_outputs(4365)) and not (layer0_outputs(4646));
    layer1_outputs(687) <= not(layer0_outputs(1117)) or (layer0_outputs(2633));
    layer1_outputs(688) <= layer0_outputs(3810);
    layer1_outputs(689) <= not((layer0_outputs(18)) or (layer0_outputs(3399)));
    layer1_outputs(690) <= not(layer0_outputs(3254));
    layer1_outputs(691) <= '1';
    layer1_outputs(692) <= '1';
    layer1_outputs(693) <= not(layer0_outputs(4608)) or (layer0_outputs(1516));
    layer1_outputs(694) <= not(layer0_outputs(4335));
    layer1_outputs(695) <= not(layer0_outputs(2290)) or (layer0_outputs(4222));
    layer1_outputs(696) <= not(layer0_outputs(370)) or (layer0_outputs(3441));
    layer1_outputs(697) <= (layer0_outputs(455)) and not (layer0_outputs(2361));
    layer1_outputs(698) <= '0';
    layer1_outputs(699) <= not(layer0_outputs(3077)) or (layer0_outputs(598));
    layer1_outputs(700) <= not((layer0_outputs(3105)) and (layer0_outputs(2984)));
    layer1_outputs(701) <= '1';
    layer1_outputs(702) <= (layer0_outputs(3113)) and not (layer0_outputs(4676));
    layer1_outputs(703) <= (layer0_outputs(1719)) and not (layer0_outputs(1379));
    layer1_outputs(704) <= not(layer0_outputs(4923)) or (layer0_outputs(1626));
    layer1_outputs(705) <= not(layer0_outputs(2125));
    layer1_outputs(706) <= '1';
    layer1_outputs(707) <= layer0_outputs(3190);
    layer1_outputs(708) <= not(layer0_outputs(3106)) or (layer0_outputs(2722));
    layer1_outputs(709) <= '0';
    layer1_outputs(710) <= not(layer0_outputs(3369)) or (layer0_outputs(3404));
    layer1_outputs(711) <= layer0_outputs(618);
    layer1_outputs(712) <= not(layer0_outputs(3112)) or (layer0_outputs(1445));
    layer1_outputs(713) <= (layer0_outputs(995)) or (layer0_outputs(3548));
    layer1_outputs(714) <= not(layer0_outputs(371)) or (layer0_outputs(1313));
    layer1_outputs(715) <= not((layer0_outputs(3920)) or (layer0_outputs(922)));
    layer1_outputs(716) <= layer0_outputs(3431);
    layer1_outputs(717) <= (layer0_outputs(1872)) or (layer0_outputs(2227));
    layer1_outputs(718) <= not(layer0_outputs(4202)) or (layer0_outputs(1349));
    layer1_outputs(719) <= not(layer0_outputs(4728)) or (layer0_outputs(182));
    layer1_outputs(720) <= (layer0_outputs(3245)) or (layer0_outputs(2076));
    layer1_outputs(721) <= '0';
    layer1_outputs(722) <= '0';
    layer1_outputs(723) <= not((layer0_outputs(261)) or (layer0_outputs(4320)));
    layer1_outputs(724) <= not((layer0_outputs(4722)) or (layer0_outputs(362)));
    layer1_outputs(725) <= '1';
    layer1_outputs(726) <= layer0_outputs(2640);
    layer1_outputs(727) <= '1';
    layer1_outputs(728) <= not(layer0_outputs(264)) or (layer0_outputs(4131));
    layer1_outputs(729) <= not(layer0_outputs(760));
    layer1_outputs(730) <= not(layer0_outputs(2335));
    layer1_outputs(731) <= not(layer0_outputs(2575)) or (layer0_outputs(3681));
    layer1_outputs(732) <= not((layer0_outputs(3215)) and (layer0_outputs(2047)));
    layer1_outputs(733) <= '0';
    layer1_outputs(734) <= not((layer0_outputs(2366)) and (layer0_outputs(318)));
    layer1_outputs(735) <= '0';
    layer1_outputs(736) <= (layer0_outputs(3144)) and not (layer0_outputs(539));
    layer1_outputs(737) <= (layer0_outputs(3088)) and not (layer0_outputs(2443));
    layer1_outputs(738) <= '0';
    layer1_outputs(739) <= (layer0_outputs(1616)) or (layer0_outputs(4654));
    layer1_outputs(740) <= '1';
    layer1_outputs(741) <= '1';
    layer1_outputs(742) <= layer0_outputs(2364);
    layer1_outputs(743) <= (layer0_outputs(2573)) and not (layer0_outputs(2766));
    layer1_outputs(744) <= '0';
    layer1_outputs(745) <= '0';
    layer1_outputs(746) <= not((layer0_outputs(2210)) or (layer0_outputs(1346)));
    layer1_outputs(747) <= (layer0_outputs(4612)) and (layer0_outputs(3158));
    layer1_outputs(748) <= (layer0_outputs(1638)) and not (layer0_outputs(2966));
    layer1_outputs(749) <= (layer0_outputs(1531)) xor (layer0_outputs(1373));
    layer1_outputs(750) <= (layer0_outputs(4246)) and (layer0_outputs(4942));
    layer1_outputs(751) <= not(layer0_outputs(1670));
    layer1_outputs(752) <= not(layer0_outputs(2636));
    layer1_outputs(753) <= '1';
    layer1_outputs(754) <= (layer0_outputs(3536)) and not (layer0_outputs(2987));
    layer1_outputs(755) <= '0';
    layer1_outputs(756) <= '1';
    layer1_outputs(757) <= '0';
    layer1_outputs(758) <= not(layer0_outputs(3374));
    layer1_outputs(759) <= '1';
    layer1_outputs(760) <= layer0_outputs(3839);
    layer1_outputs(761) <= not((layer0_outputs(3333)) xor (layer0_outputs(880)));
    layer1_outputs(762) <= '1';
    layer1_outputs(763) <= not(layer0_outputs(4296)) or (layer0_outputs(3067));
    layer1_outputs(764) <= not((layer0_outputs(1225)) or (layer0_outputs(3013)));
    layer1_outputs(765) <= layer0_outputs(612);
    layer1_outputs(766) <= '0';
    layer1_outputs(767) <= '0';
    layer1_outputs(768) <= (layer0_outputs(4982)) and (layer0_outputs(4671));
    layer1_outputs(769) <= not((layer0_outputs(5034)) or (layer0_outputs(1249)));
    layer1_outputs(770) <= (layer0_outputs(2680)) and (layer0_outputs(3835));
    layer1_outputs(771) <= '1';
    layer1_outputs(772) <= '0';
    layer1_outputs(773) <= (layer0_outputs(634)) or (layer0_outputs(2771));
    layer1_outputs(774) <= (layer0_outputs(4218)) and (layer0_outputs(2421));
    layer1_outputs(775) <= layer0_outputs(3727);
    layer1_outputs(776) <= not((layer0_outputs(3230)) and (layer0_outputs(4848)));
    layer1_outputs(777) <= layer0_outputs(2296);
    layer1_outputs(778) <= not((layer0_outputs(4203)) xor (layer0_outputs(1041)));
    layer1_outputs(779) <= (layer0_outputs(3817)) and (layer0_outputs(161));
    layer1_outputs(780) <= (layer0_outputs(3886)) or (layer0_outputs(4136));
    layer1_outputs(781) <= not(layer0_outputs(1312)) or (layer0_outputs(3119));
    layer1_outputs(782) <= not((layer0_outputs(1527)) and (layer0_outputs(3035)));
    layer1_outputs(783) <= not((layer0_outputs(3913)) and (layer0_outputs(170)));
    layer1_outputs(784) <= (layer0_outputs(670)) or (layer0_outputs(3031));
    layer1_outputs(785) <= not(layer0_outputs(1753));
    layer1_outputs(786) <= not((layer0_outputs(4863)) and (layer0_outputs(5114)));
    layer1_outputs(787) <= (layer0_outputs(4258)) and not (layer0_outputs(668));
    layer1_outputs(788) <= not((layer0_outputs(3846)) and (layer0_outputs(1233)));
    layer1_outputs(789) <= '1';
    layer1_outputs(790) <= (layer0_outputs(1027)) and not (layer0_outputs(3444));
    layer1_outputs(791) <= (layer0_outputs(4238)) and not (layer0_outputs(5089));
    layer1_outputs(792) <= '1';
    layer1_outputs(793) <= not(layer0_outputs(1000)) or (layer0_outputs(4831));
    layer1_outputs(794) <= '1';
    layer1_outputs(795) <= (layer0_outputs(4416)) or (layer0_outputs(1791));
    layer1_outputs(796) <= (layer0_outputs(4838)) and (layer0_outputs(4767));
    layer1_outputs(797) <= '0';
    layer1_outputs(798) <= not(layer0_outputs(4289)) or (layer0_outputs(2728));
    layer1_outputs(799) <= not((layer0_outputs(1868)) or (layer0_outputs(1763)));
    layer1_outputs(800) <= (layer0_outputs(812)) and not (layer0_outputs(828));
    layer1_outputs(801) <= not((layer0_outputs(2639)) or (layer0_outputs(3279)));
    layer1_outputs(802) <= (layer0_outputs(2116)) or (layer0_outputs(1845));
    layer1_outputs(803) <= layer0_outputs(176);
    layer1_outputs(804) <= not(layer0_outputs(2625));
    layer1_outputs(805) <= '0';
    layer1_outputs(806) <= not(layer0_outputs(3744)) or (layer0_outputs(1215));
    layer1_outputs(807) <= layer0_outputs(2967);
    layer1_outputs(808) <= not((layer0_outputs(4180)) or (layer0_outputs(4256)));
    layer1_outputs(809) <= not((layer0_outputs(4670)) or (layer0_outputs(245)));
    layer1_outputs(810) <= '0';
    layer1_outputs(811) <= (layer0_outputs(3851)) or (layer0_outputs(3704));
    layer1_outputs(812) <= not(layer0_outputs(1841));
    layer1_outputs(813) <= layer0_outputs(491);
    layer1_outputs(814) <= (layer0_outputs(572)) and not (layer0_outputs(1039));
    layer1_outputs(815) <= '1';
    layer1_outputs(816) <= layer0_outputs(2058);
    layer1_outputs(817) <= not(layer0_outputs(4397));
    layer1_outputs(818) <= not((layer0_outputs(1024)) and (layer0_outputs(2600)));
    layer1_outputs(819) <= '1';
    layer1_outputs(820) <= (layer0_outputs(841)) and not (layer0_outputs(3284));
    layer1_outputs(821) <= '0';
    layer1_outputs(822) <= (layer0_outputs(2616)) and not (layer0_outputs(4092));
    layer1_outputs(823) <= '1';
    layer1_outputs(824) <= (layer0_outputs(4073)) and not (layer0_outputs(867));
    layer1_outputs(825) <= '0';
    layer1_outputs(826) <= not((layer0_outputs(5072)) or (layer0_outputs(4116)));
    layer1_outputs(827) <= '1';
    layer1_outputs(828) <= '1';
    layer1_outputs(829) <= not(layer0_outputs(2450));
    layer1_outputs(830) <= '1';
    layer1_outputs(831) <= not(layer0_outputs(2574));
    layer1_outputs(832) <= layer0_outputs(2898);
    layer1_outputs(833) <= not((layer0_outputs(841)) and (layer0_outputs(1501)));
    layer1_outputs(834) <= '0';
    layer1_outputs(835) <= not((layer0_outputs(5087)) or (layer0_outputs(4748)));
    layer1_outputs(836) <= layer0_outputs(2809);
    layer1_outputs(837) <= not((layer0_outputs(2525)) or (layer0_outputs(218)));
    layer1_outputs(838) <= (layer0_outputs(3126)) and (layer0_outputs(3492));
    layer1_outputs(839) <= not(layer0_outputs(2912));
    layer1_outputs(840) <= '1';
    layer1_outputs(841) <= not(layer0_outputs(4137)) or (layer0_outputs(4568));
    layer1_outputs(842) <= (layer0_outputs(1276)) or (layer0_outputs(3338));
    layer1_outputs(843) <= (layer0_outputs(4937)) and not (layer0_outputs(2628));
    layer1_outputs(844) <= (layer0_outputs(4915)) and not (layer0_outputs(3138));
    layer1_outputs(845) <= '0';
    layer1_outputs(846) <= not((layer0_outputs(1773)) and (layer0_outputs(4941)));
    layer1_outputs(847) <= (layer0_outputs(1721)) and (layer0_outputs(3757));
    layer1_outputs(848) <= not(layer0_outputs(3613)) or (layer0_outputs(4232));
    layer1_outputs(849) <= not(layer0_outputs(1081));
    layer1_outputs(850) <= layer0_outputs(4842);
    layer1_outputs(851) <= layer0_outputs(3975);
    layer1_outputs(852) <= '1';
    layer1_outputs(853) <= '0';
    layer1_outputs(854) <= layer0_outputs(1217);
    layer1_outputs(855) <= '1';
    layer1_outputs(856) <= layer0_outputs(22);
    layer1_outputs(857) <= (layer0_outputs(185)) or (layer0_outputs(2625));
    layer1_outputs(858) <= layer0_outputs(3822);
    layer1_outputs(859) <= '1';
    layer1_outputs(860) <= (layer0_outputs(3082)) and (layer0_outputs(1008));
    layer1_outputs(861) <= '0';
    layer1_outputs(862) <= (layer0_outputs(2526)) and not (layer0_outputs(2801));
    layer1_outputs(863) <= '1';
    layer1_outputs(864) <= not(layer0_outputs(3154));
    layer1_outputs(865) <= layer0_outputs(4782);
    layer1_outputs(866) <= '1';
    layer1_outputs(867) <= '0';
    layer1_outputs(868) <= not(layer0_outputs(1922)) or (layer0_outputs(2604));
    layer1_outputs(869) <= not(layer0_outputs(980)) or (layer0_outputs(4338));
    layer1_outputs(870) <= layer0_outputs(271);
    layer1_outputs(871) <= layer0_outputs(898);
    layer1_outputs(872) <= not((layer0_outputs(1374)) and (layer0_outputs(4248)));
    layer1_outputs(873) <= not(layer0_outputs(1139));
    layer1_outputs(874) <= (layer0_outputs(4656)) or (layer0_outputs(430));
    layer1_outputs(875) <= (layer0_outputs(3753)) and not (layer0_outputs(1250));
    layer1_outputs(876) <= not(layer0_outputs(1088));
    layer1_outputs(877) <= '1';
    layer1_outputs(878) <= '1';
    layer1_outputs(879) <= not((layer0_outputs(9)) and (layer0_outputs(981)));
    layer1_outputs(880) <= (layer0_outputs(2136)) and not (layer0_outputs(454));
    layer1_outputs(881) <= not(layer0_outputs(1072));
    layer1_outputs(882) <= not((layer0_outputs(466)) and (layer0_outputs(4751)));
    layer1_outputs(883) <= '1';
    layer1_outputs(884) <= not(layer0_outputs(4954)) or (layer0_outputs(1009));
    layer1_outputs(885) <= not(layer0_outputs(1592));
    layer1_outputs(886) <= (layer0_outputs(1666)) and (layer0_outputs(3511));
    layer1_outputs(887) <= (layer0_outputs(5004)) and not (layer0_outputs(1654));
    layer1_outputs(888) <= layer0_outputs(4460);
    layer1_outputs(889) <= (layer0_outputs(3329)) xor (layer0_outputs(2429));
    layer1_outputs(890) <= layer0_outputs(1788);
    layer1_outputs(891) <= '1';
    layer1_outputs(892) <= not((layer0_outputs(328)) or (layer0_outputs(3867)));
    layer1_outputs(893) <= not(layer0_outputs(1819));
    layer1_outputs(894) <= not(layer0_outputs(2067)) or (layer0_outputs(574));
    layer1_outputs(895) <= not(layer0_outputs(509));
    layer1_outputs(896) <= '1';
    layer1_outputs(897) <= layer0_outputs(3776);
    layer1_outputs(898) <= layer0_outputs(986);
    layer1_outputs(899) <= '1';
    layer1_outputs(900) <= not(layer0_outputs(2847));
    layer1_outputs(901) <= (layer0_outputs(5049)) and not (layer0_outputs(5079));
    layer1_outputs(902) <= (layer0_outputs(3926)) and not (layer0_outputs(237));
    layer1_outputs(903) <= not(layer0_outputs(3004)) or (layer0_outputs(233));
    layer1_outputs(904) <= (layer0_outputs(1280)) and (layer0_outputs(691));
    layer1_outputs(905) <= layer0_outputs(2054);
    layer1_outputs(906) <= (layer0_outputs(192)) or (layer0_outputs(1616));
    layer1_outputs(907) <= not(layer0_outputs(4563)) or (layer0_outputs(3674));
    layer1_outputs(908) <= '0';
    layer1_outputs(909) <= not((layer0_outputs(3341)) and (layer0_outputs(1895)));
    layer1_outputs(910) <= (layer0_outputs(1724)) and not (layer0_outputs(2350));
    layer1_outputs(911) <= (layer0_outputs(2022)) or (layer0_outputs(2391));
    layer1_outputs(912) <= '0';
    layer1_outputs(913) <= not(layer0_outputs(3506));
    layer1_outputs(914) <= not(layer0_outputs(544));
    layer1_outputs(915) <= '1';
    layer1_outputs(916) <= '1';
    layer1_outputs(917) <= '0';
    layer1_outputs(918) <= '0';
    layer1_outputs(919) <= (layer0_outputs(3728)) and not (layer0_outputs(4224));
    layer1_outputs(920) <= (layer0_outputs(1947)) and not (layer0_outputs(1390));
    layer1_outputs(921) <= '1';
    layer1_outputs(922) <= '0';
    layer1_outputs(923) <= (layer0_outputs(1132)) or (layer0_outputs(1589));
    layer1_outputs(924) <= '0';
    layer1_outputs(925) <= '1';
    layer1_outputs(926) <= '1';
    layer1_outputs(927) <= not(layer0_outputs(4034));
    layer1_outputs(928) <= not((layer0_outputs(5090)) and (layer0_outputs(474)));
    layer1_outputs(929) <= not(layer0_outputs(2476)) or (layer0_outputs(4278));
    layer1_outputs(930) <= not(layer0_outputs(4413));
    layer1_outputs(931) <= not((layer0_outputs(2448)) and (layer0_outputs(4691)));
    layer1_outputs(932) <= (layer0_outputs(2082)) and not (layer0_outputs(1942));
    layer1_outputs(933) <= '0';
    layer1_outputs(934) <= (layer0_outputs(4710)) and not (layer0_outputs(572));
    layer1_outputs(935) <= '0';
    layer1_outputs(936) <= layer0_outputs(4727);
    layer1_outputs(937) <= layer0_outputs(4127);
    layer1_outputs(938) <= (layer0_outputs(2927)) and (layer0_outputs(2177));
    layer1_outputs(939) <= not(layer0_outputs(2266));
    layer1_outputs(940) <= not(layer0_outputs(1936)) or (layer0_outputs(1604));
    layer1_outputs(941) <= not(layer0_outputs(3005));
    layer1_outputs(942) <= (layer0_outputs(1235)) and (layer0_outputs(3994));
    layer1_outputs(943) <= '1';
    layer1_outputs(944) <= not(layer0_outputs(1154));
    layer1_outputs(945) <= (layer0_outputs(1265)) and not (layer0_outputs(4362));
    layer1_outputs(946) <= (layer0_outputs(3904)) and (layer0_outputs(4587));
    layer1_outputs(947) <= not(layer0_outputs(2018)) or (layer0_outputs(1035));
    layer1_outputs(948) <= not((layer0_outputs(1996)) or (layer0_outputs(1198)));
    layer1_outputs(949) <= '0';
    layer1_outputs(950) <= not(layer0_outputs(3135)) or (layer0_outputs(1153));
    layer1_outputs(951) <= layer0_outputs(247);
    layer1_outputs(952) <= '0';
    layer1_outputs(953) <= layer0_outputs(3844);
    layer1_outputs(954) <= '0';
    layer1_outputs(955) <= (layer0_outputs(2363)) or (layer0_outputs(13));
    layer1_outputs(956) <= '1';
    layer1_outputs(957) <= (layer0_outputs(72)) xor (layer0_outputs(4989));
    layer1_outputs(958) <= not(layer0_outputs(3956));
    layer1_outputs(959) <= (layer0_outputs(1783)) or (layer0_outputs(3591));
    layer1_outputs(960) <= not((layer0_outputs(3636)) or (layer0_outputs(1165)));
    layer1_outputs(961) <= not((layer0_outputs(2254)) and (layer0_outputs(1512)));
    layer1_outputs(962) <= '0';
    layer1_outputs(963) <= not(layer0_outputs(4487));
    layer1_outputs(964) <= layer0_outputs(1955);
    layer1_outputs(965) <= (layer0_outputs(2654)) or (layer0_outputs(1204));
    layer1_outputs(966) <= not(layer0_outputs(1747)) or (layer0_outputs(3067));
    layer1_outputs(967) <= layer0_outputs(5116);
    layer1_outputs(968) <= '0';
    layer1_outputs(969) <= not(layer0_outputs(3304));
    layer1_outputs(970) <= not((layer0_outputs(4070)) or (layer0_outputs(3165)));
    layer1_outputs(971) <= '0';
    layer1_outputs(972) <= not(layer0_outputs(2204)) or (layer0_outputs(4325));
    layer1_outputs(973) <= '0';
    layer1_outputs(974) <= not(layer0_outputs(1504)) or (layer0_outputs(2408));
    layer1_outputs(975) <= not(layer0_outputs(3344)) or (layer0_outputs(4075));
    layer1_outputs(976) <= (layer0_outputs(3361)) or (layer0_outputs(2858));
    layer1_outputs(977) <= (layer0_outputs(3592)) or (layer0_outputs(2229));
    layer1_outputs(978) <= (layer0_outputs(4137)) and not (layer0_outputs(2733));
    layer1_outputs(979) <= '0';
    layer1_outputs(980) <= not((layer0_outputs(1672)) xor (layer0_outputs(1848)));
    layer1_outputs(981) <= (layer0_outputs(1677)) xor (layer0_outputs(2276));
    layer1_outputs(982) <= not(layer0_outputs(3387)) or (layer0_outputs(3924));
    layer1_outputs(983) <= not(layer0_outputs(3833)) or (layer0_outputs(3429));
    layer1_outputs(984) <= '0';
    layer1_outputs(985) <= '1';
    layer1_outputs(986) <= layer0_outputs(2523);
    layer1_outputs(987) <= (layer0_outputs(4778)) and not (layer0_outputs(620));
    layer1_outputs(988) <= (layer0_outputs(2631)) or (layer0_outputs(3212));
    layer1_outputs(989) <= (layer0_outputs(2973)) and (layer0_outputs(433));
    layer1_outputs(990) <= '0';
    layer1_outputs(991) <= (layer0_outputs(4945)) xor (layer0_outputs(2303));
    layer1_outputs(992) <= not((layer0_outputs(1744)) xor (layer0_outputs(307)));
    layer1_outputs(993) <= '1';
    layer1_outputs(994) <= '0';
    layer1_outputs(995) <= (layer0_outputs(510)) and not (layer0_outputs(4847));
    layer1_outputs(996) <= '0';
    layer1_outputs(997) <= not((layer0_outputs(3487)) and (layer0_outputs(3299)));
    layer1_outputs(998) <= not((layer0_outputs(688)) and (layer0_outputs(3573)));
    layer1_outputs(999) <= '1';
    layer1_outputs(1000) <= '1';
    layer1_outputs(1001) <= (layer0_outputs(4883)) or (layer0_outputs(2037));
    layer1_outputs(1002) <= '1';
    layer1_outputs(1003) <= layer0_outputs(1238);
    layer1_outputs(1004) <= not((layer0_outputs(4119)) and (layer0_outputs(3117)));
    layer1_outputs(1005) <= '0';
    layer1_outputs(1006) <= (layer0_outputs(4540)) and not (layer0_outputs(1462));
    layer1_outputs(1007) <= (layer0_outputs(526)) and (layer0_outputs(474));
    layer1_outputs(1008) <= not(layer0_outputs(2775)) or (layer0_outputs(2081));
    layer1_outputs(1009) <= (layer0_outputs(4564)) and not (layer0_outputs(4772));
    layer1_outputs(1010) <= (layer0_outputs(3803)) and not (layer0_outputs(4570));
    layer1_outputs(1011) <= (layer0_outputs(5080)) and not (layer0_outputs(1054));
    layer1_outputs(1012) <= not(layer0_outputs(2034)) or (layer0_outputs(2438));
    layer1_outputs(1013) <= layer0_outputs(4090);
    layer1_outputs(1014) <= not((layer0_outputs(4615)) and (layer0_outputs(512)));
    layer1_outputs(1015) <= '0';
    layer1_outputs(1016) <= not((layer0_outputs(3350)) or (layer0_outputs(2150)));
    layer1_outputs(1017) <= not(layer0_outputs(2131)) or (layer0_outputs(4096));
    layer1_outputs(1018) <= not(layer0_outputs(2589)) or (layer0_outputs(844));
    layer1_outputs(1019) <= not(layer0_outputs(3209)) or (layer0_outputs(2056));
    layer1_outputs(1020) <= '0';
    layer1_outputs(1021) <= (layer0_outputs(1840)) and not (layer0_outputs(3853));
    layer1_outputs(1022) <= not(layer0_outputs(47)) or (layer0_outputs(1578));
    layer1_outputs(1023) <= '1';
    layer1_outputs(1024) <= '1';
    layer1_outputs(1025) <= '0';
    layer1_outputs(1026) <= not(layer0_outputs(1017)) or (layer0_outputs(395));
    layer1_outputs(1027) <= not(layer0_outputs(870)) or (layer0_outputs(2493));
    layer1_outputs(1028) <= '1';
    layer1_outputs(1029) <= layer0_outputs(4031);
    layer1_outputs(1030) <= (layer0_outputs(882)) and (layer0_outputs(554));
    layer1_outputs(1031) <= not(layer0_outputs(3477));
    layer1_outputs(1032) <= '1';
    layer1_outputs(1033) <= (layer0_outputs(1392)) or (layer0_outputs(2000));
    layer1_outputs(1034) <= not(layer0_outputs(2386));
    layer1_outputs(1035) <= (layer0_outputs(3196)) and not (layer0_outputs(3679));
    layer1_outputs(1036) <= '0';
    layer1_outputs(1037) <= not((layer0_outputs(1979)) and (layer0_outputs(3970)));
    layer1_outputs(1038) <= '0';
    layer1_outputs(1039) <= (layer0_outputs(4763)) or (layer0_outputs(2073));
    layer1_outputs(1040) <= not(layer0_outputs(365)) or (layer0_outputs(152));
    layer1_outputs(1041) <= not((layer0_outputs(3380)) and (layer0_outputs(2077)));
    layer1_outputs(1042) <= not(layer0_outputs(217)) or (layer0_outputs(1067));
    layer1_outputs(1043) <= '0';
    layer1_outputs(1044) <= '0';
    layer1_outputs(1045) <= (layer0_outputs(3608)) and (layer0_outputs(2020));
    layer1_outputs(1046) <= '1';
    layer1_outputs(1047) <= not(layer0_outputs(2907)) or (layer0_outputs(795));
    layer1_outputs(1048) <= '1';
    layer1_outputs(1049) <= '0';
    layer1_outputs(1050) <= '1';
    layer1_outputs(1051) <= not((layer0_outputs(5025)) or (layer0_outputs(1661)));
    layer1_outputs(1052) <= layer0_outputs(3433);
    layer1_outputs(1053) <= not((layer0_outputs(399)) and (layer0_outputs(350)));
    layer1_outputs(1054) <= layer0_outputs(4162);
    layer1_outputs(1055) <= '0';
    layer1_outputs(1056) <= layer0_outputs(4367);
    layer1_outputs(1057) <= '1';
    layer1_outputs(1058) <= (layer0_outputs(4529)) and (layer0_outputs(3551));
    layer1_outputs(1059) <= not(layer0_outputs(4028)) or (layer0_outputs(3198));
    layer1_outputs(1060) <= '0';
    layer1_outputs(1061) <= (layer0_outputs(4274)) and not (layer0_outputs(2866));
    layer1_outputs(1062) <= not(layer0_outputs(3486)) or (layer0_outputs(3086));
    layer1_outputs(1063) <= (layer0_outputs(2450)) or (layer0_outputs(2895));
    layer1_outputs(1064) <= not(layer0_outputs(3505)) or (layer0_outputs(1696));
    layer1_outputs(1065) <= layer0_outputs(5113);
    layer1_outputs(1066) <= (layer0_outputs(1693)) and not (layer0_outputs(2193));
    layer1_outputs(1067) <= not((layer0_outputs(1102)) and (layer0_outputs(2028)));
    layer1_outputs(1068) <= (layer0_outputs(1334)) and not (layer0_outputs(1061));
    layer1_outputs(1069) <= '1';
    layer1_outputs(1070) <= '1';
    layer1_outputs(1071) <= not(layer0_outputs(844)) or (layer0_outputs(947));
    layer1_outputs(1072) <= '1';
    layer1_outputs(1073) <= '0';
    layer1_outputs(1074) <= layer0_outputs(4277);
    layer1_outputs(1075) <= '0';
    layer1_outputs(1076) <= (layer0_outputs(2877)) and not (layer0_outputs(77));
    layer1_outputs(1077) <= not(layer0_outputs(404)) or (layer0_outputs(4200));
    layer1_outputs(1078) <= layer0_outputs(580);
    layer1_outputs(1079) <= '0';
    layer1_outputs(1080) <= not(layer0_outputs(441)) or (layer0_outputs(2585));
    layer1_outputs(1081) <= not(layer0_outputs(2485));
    layer1_outputs(1082) <= not((layer0_outputs(3057)) xor (layer0_outputs(2166)));
    layer1_outputs(1083) <= not((layer0_outputs(1528)) or (layer0_outputs(4116)));
    layer1_outputs(1084) <= (layer0_outputs(1445)) and not (layer0_outputs(5089));
    layer1_outputs(1085) <= (layer0_outputs(3159)) and (layer0_outputs(4695));
    layer1_outputs(1086) <= not(layer0_outputs(2753));
    layer1_outputs(1087) <= not((layer0_outputs(1013)) xor (layer0_outputs(894)));
    layer1_outputs(1088) <= layer0_outputs(2068);
    layer1_outputs(1089) <= layer0_outputs(2366);
    layer1_outputs(1090) <= (layer0_outputs(1939)) or (layer0_outputs(17));
    layer1_outputs(1091) <= not((layer0_outputs(4138)) and (layer0_outputs(2885)));
    layer1_outputs(1092) <= not(layer0_outputs(3125));
    layer1_outputs(1093) <= '1';
    layer1_outputs(1094) <= (layer0_outputs(1103)) and not (layer0_outputs(3152));
    layer1_outputs(1095) <= '0';
    layer1_outputs(1096) <= '0';
    layer1_outputs(1097) <= '0';
    layer1_outputs(1098) <= layer0_outputs(503);
    layer1_outputs(1099) <= not(layer0_outputs(224));
    layer1_outputs(1100) <= '1';
    layer1_outputs(1101) <= not(layer0_outputs(680)) or (layer0_outputs(4025));
    layer1_outputs(1102) <= '1';
    layer1_outputs(1103) <= (layer0_outputs(4391)) and not (layer0_outputs(1619));
    layer1_outputs(1104) <= not(layer0_outputs(625)) or (layer0_outputs(91));
    layer1_outputs(1105) <= '0';
    layer1_outputs(1106) <= not(layer0_outputs(4522)) or (layer0_outputs(1208));
    layer1_outputs(1107) <= '1';
    layer1_outputs(1108) <= not(layer0_outputs(426)) or (layer0_outputs(4870));
    layer1_outputs(1109) <= layer0_outputs(290);
    layer1_outputs(1110) <= (layer0_outputs(4721)) or (layer0_outputs(4350));
    layer1_outputs(1111) <= not(layer0_outputs(2483));
    layer1_outputs(1112) <= not((layer0_outputs(4145)) or (layer0_outputs(3456)));
    layer1_outputs(1113) <= '0';
    layer1_outputs(1114) <= not(layer0_outputs(455)) or (layer0_outputs(657));
    layer1_outputs(1115) <= (layer0_outputs(3391)) and not (layer0_outputs(1206));
    layer1_outputs(1116) <= '1';
    layer1_outputs(1117) <= '0';
    layer1_outputs(1118) <= layer0_outputs(900);
    layer1_outputs(1119) <= (layer0_outputs(490)) and not (layer0_outputs(1653));
    layer1_outputs(1120) <= not((layer0_outputs(2690)) or (layer0_outputs(4748)));
    layer1_outputs(1121) <= layer0_outputs(2931);
    layer1_outputs(1122) <= not(layer0_outputs(3439)) or (layer0_outputs(2622));
    layer1_outputs(1123) <= '0';
    layer1_outputs(1124) <= '0';
    layer1_outputs(1125) <= not(layer0_outputs(4635)) or (layer0_outputs(859));
    layer1_outputs(1126) <= layer0_outputs(214);
    layer1_outputs(1127) <= (layer0_outputs(1705)) and (layer0_outputs(4405));
    layer1_outputs(1128) <= '1';
    layer1_outputs(1129) <= not(layer0_outputs(4786)) or (layer0_outputs(4980));
    layer1_outputs(1130) <= (layer0_outputs(716)) and not (layer0_outputs(2765));
    layer1_outputs(1131) <= layer0_outputs(1443);
    layer1_outputs(1132) <= not(layer0_outputs(1591));
    layer1_outputs(1133) <= not(layer0_outputs(2412)) or (layer0_outputs(4197));
    layer1_outputs(1134) <= not(layer0_outputs(4052));
    layer1_outputs(1135) <= not((layer0_outputs(3351)) or (layer0_outputs(1646)));
    layer1_outputs(1136) <= not((layer0_outputs(1386)) and (layer0_outputs(975)));
    layer1_outputs(1137) <= not((layer0_outputs(776)) and (layer0_outputs(153)));
    layer1_outputs(1138) <= not(layer0_outputs(4558)) or (layer0_outputs(2233));
    layer1_outputs(1139) <= (layer0_outputs(4636)) and not (layer0_outputs(3653));
    layer1_outputs(1140) <= not(layer0_outputs(2893)) or (layer0_outputs(139));
    layer1_outputs(1141) <= (layer0_outputs(886)) and not (layer0_outputs(1611));
    layer1_outputs(1142) <= not(layer0_outputs(4809));
    layer1_outputs(1143) <= '0';
    layer1_outputs(1144) <= not((layer0_outputs(4663)) or (layer0_outputs(516)));
    layer1_outputs(1145) <= '0';
    layer1_outputs(1146) <= '0';
    layer1_outputs(1147) <= layer0_outputs(1003);
    layer1_outputs(1148) <= (layer0_outputs(3239)) and not (layer0_outputs(520));
    layer1_outputs(1149) <= (layer0_outputs(3868)) and not (layer0_outputs(3213));
    layer1_outputs(1150) <= not((layer0_outputs(2002)) or (layer0_outputs(2726)));
    layer1_outputs(1151) <= layer0_outputs(3713);
    layer1_outputs(1152) <= not((layer0_outputs(3337)) xor (layer0_outputs(792)));
    layer1_outputs(1153) <= (layer0_outputs(2387)) and (layer0_outputs(681));
    layer1_outputs(1154) <= (layer0_outputs(5101)) and not (layer0_outputs(310));
    layer1_outputs(1155) <= layer0_outputs(3128);
    layer1_outputs(1156) <= '1';
    layer1_outputs(1157) <= (layer0_outputs(419)) or (layer0_outputs(3244));
    layer1_outputs(1158) <= not(layer0_outputs(3146));
    layer1_outputs(1159) <= not(layer0_outputs(3610));
    layer1_outputs(1160) <= not(layer0_outputs(3400));
    layer1_outputs(1161) <= not((layer0_outputs(4048)) or (layer0_outputs(4932)));
    layer1_outputs(1162) <= not(layer0_outputs(2566));
    layer1_outputs(1163) <= not(layer0_outputs(785)) or (layer0_outputs(3543));
    layer1_outputs(1164) <= not((layer0_outputs(4408)) and (layer0_outputs(4598)));
    layer1_outputs(1165) <= '0';
    layer1_outputs(1166) <= layer0_outputs(3371);
    layer1_outputs(1167) <= not(layer0_outputs(636)) or (layer0_outputs(1683));
    layer1_outputs(1168) <= (layer0_outputs(2586)) or (layer0_outputs(2505));
    layer1_outputs(1169) <= not(layer0_outputs(3879));
    layer1_outputs(1170) <= (layer0_outputs(3988)) and not (layer0_outputs(738));
    layer1_outputs(1171) <= (layer0_outputs(383)) and not (layer0_outputs(2214));
    layer1_outputs(1172) <= '0';
    layer1_outputs(1173) <= not((layer0_outputs(1711)) or (layer0_outputs(4590)));
    layer1_outputs(1174) <= layer0_outputs(3553);
    layer1_outputs(1175) <= '1';
    layer1_outputs(1176) <= layer0_outputs(3297);
    layer1_outputs(1177) <= layer0_outputs(4854);
    layer1_outputs(1178) <= '0';
    layer1_outputs(1179) <= not(layer0_outputs(3296));
    layer1_outputs(1180) <= layer0_outputs(3576);
    layer1_outputs(1181) <= not(layer0_outputs(4570)) or (layer0_outputs(4869));
    layer1_outputs(1182) <= not(layer0_outputs(4920)) or (layer0_outputs(1533));
    layer1_outputs(1183) <= '1';
    layer1_outputs(1184) <= not((layer0_outputs(1734)) or (layer0_outputs(3519)));
    layer1_outputs(1185) <= not(layer0_outputs(4094)) or (layer0_outputs(4770));
    layer1_outputs(1186) <= not((layer0_outputs(4745)) and (layer0_outputs(2979)));
    layer1_outputs(1187) <= layer0_outputs(4104);
    layer1_outputs(1188) <= layer0_outputs(213);
    layer1_outputs(1189) <= not(layer0_outputs(2772)) or (layer0_outputs(4835));
    layer1_outputs(1190) <= layer0_outputs(320);
    layer1_outputs(1191) <= (layer0_outputs(2994)) or (layer0_outputs(4737));
    layer1_outputs(1192) <= not(layer0_outputs(3348));
    layer1_outputs(1193) <= '0';
    layer1_outputs(1194) <= '0';
    layer1_outputs(1195) <= (layer0_outputs(3499)) and not (layer0_outputs(606));
    layer1_outputs(1196) <= not(layer0_outputs(1797));
    layer1_outputs(1197) <= '0';
    layer1_outputs(1198) <= layer0_outputs(958);
    layer1_outputs(1199) <= layer0_outputs(2577);
    layer1_outputs(1200) <= '1';
    layer1_outputs(1201) <= layer0_outputs(2039);
    layer1_outputs(1202) <= (layer0_outputs(4714)) and (layer0_outputs(4981));
    layer1_outputs(1203) <= '0';
    layer1_outputs(1204) <= '0';
    layer1_outputs(1205) <= layer0_outputs(2101);
    layer1_outputs(1206) <= not((layer0_outputs(380)) and (layer0_outputs(5004)));
    layer1_outputs(1207) <= (layer0_outputs(1934)) and not (layer0_outputs(3942));
    layer1_outputs(1208) <= not((layer0_outputs(32)) and (layer0_outputs(1523)));
    layer1_outputs(1209) <= '1';
    layer1_outputs(1210) <= not(layer0_outputs(4193));
    layer1_outputs(1211) <= layer0_outputs(1664);
    layer1_outputs(1212) <= not(layer0_outputs(2747)) or (layer0_outputs(2963));
    layer1_outputs(1213) <= layer0_outputs(4210);
    layer1_outputs(1214) <= '1';
    layer1_outputs(1215) <= (layer0_outputs(3937)) and not (layer0_outputs(992));
    layer1_outputs(1216) <= layer0_outputs(3363);
    layer1_outputs(1217) <= '1';
    layer1_outputs(1218) <= not((layer0_outputs(713)) or (layer0_outputs(2532)));
    layer1_outputs(1219) <= not(layer0_outputs(1304)) or (layer0_outputs(279));
    layer1_outputs(1220) <= not(layer0_outputs(4504));
    layer1_outputs(1221) <= layer0_outputs(1758);
    layer1_outputs(1222) <= '1';
    layer1_outputs(1223) <= layer0_outputs(556);
    layer1_outputs(1224) <= layer0_outputs(3442);
    layer1_outputs(1225) <= not((layer0_outputs(3327)) and (layer0_outputs(5058)));
    layer1_outputs(1226) <= not(layer0_outputs(2017)) or (layer0_outputs(3968));
    layer1_outputs(1227) <= '1';
    layer1_outputs(1228) <= (layer0_outputs(2911)) and not (layer0_outputs(4033));
    layer1_outputs(1229) <= not(layer0_outputs(4641)) or (layer0_outputs(4762));
    layer1_outputs(1230) <= not(layer0_outputs(669)) or (layer0_outputs(2184));
    layer1_outputs(1231) <= not((layer0_outputs(3729)) or (layer0_outputs(2351)));
    layer1_outputs(1232) <= (layer0_outputs(55)) or (layer0_outputs(1426));
    layer1_outputs(1233) <= '0';
    layer1_outputs(1234) <= not(layer0_outputs(4819)) or (layer0_outputs(2646));
    layer1_outputs(1235) <= not(layer0_outputs(3783));
    layer1_outputs(1236) <= '1';
    layer1_outputs(1237) <= not((layer0_outputs(2358)) and (layer0_outputs(429)));
    layer1_outputs(1238) <= (layer0_outputs(3631)) and not (layer0_outputs(451));
    layer1_outputs(1239) <= not(layer0_outputs(2710)) or (layer0_outputs(2712));
    layer1_outputs(1240) <= layer0_outputs(1092);
    layer1_outputs(1241) <= not(layer0_outputs(1650)) or (layer0_outputs(411));
    layer1_outputs(1242) <= (layer0_outputs(3202)) and not (layer0_outputs(435));
    layer1_outputs(1243) <= not(layer0_outputs(681)) or (layer0_outputs(2687));
    layer1_outputs(1244) <= not((layer0_outputs(431)) or (layer0_outputs(3458)));
    layer1_outputs(1245) <= layer0_outputs(1988);
    layer1_outputs(1246) <= '1';
    layer1_outputs(1247) <= (layer0_outputs(2990)) or (layer0_outputs(395));
    layer1_outputs(1248) <= not(layer0_outputs(1772)) or (layer0_outputs(1303));
    layer1_outputs(1249) <= (layer0_outputs(4452)) and (layer0_outputs(125));
    layer1_outputs(1250) <= (layer0_outputs(1721)) and not (layer0_outputs(2896));
    layer1_outputs(1251) <= (layer0_outputs(846)) or (layer0_outputs(195));
    layer1_outputs(1252) <= not(layer0_outputs(401)) or (layer0_outputs(4732));
    layer1_outputs(1253) <= '0';
    layer1_outputs(1254) <= (layer0_outputs(2553)) and not (layer0_outputs(4638));
    layer1_outputs(1255) <= (layer0_outputs(4477)) and not (layer0_outputs(4744));
    layer1_outputs(1256) <= (layer0_outputs(2891)) and not (layer0_outputs(1243));
    layer1_outputs(1257) <= '1';
    layer1_outputs(1258) <= not((layer0_outputs(2612)) or (layer0_outputs(1575)));
    layer1_outputs(1259) <= not(layer0_outputs(303)) or (layer0_outputs(187));
    layer1_outputs(1260) <= (layer0_outputs(1127)) and not (layer0_outputs(1785));
    layer1_outputs(1261) <= not((layer0_outputs(1712)) or (layer0_outputs(1136)));
    layer1_outputs(1262) <= '1';
    layer1_outputs(1263) <= '1';
    layer1_outputs(1264) <= not((layer0_outputs(564)) and (layer0_outputs(1923)));
    layer1_outputs(1265) <= '0';
    layer1_outputs(1266) <= not(layer0_outputs(1440)) or (layer0_outputs(269));
    layer1_outputs(1267) <= '0';
    layer1_outputs(1268) <= not((layer0_outputs(3870)) or (layer0_outputs(2799)));
    layer1_outputs(1269) <= not(layer0_outputs(3757)) or (layer0_outputs(2237));
    layer1_outputs(1270) <= (layer0_outputs(2836)) and (layer0_outputs(1521));
    layer1_outputs(1271) <= (layer0_outputs(1473)) xor (layer0_outputs(546));
    layer1_outputs(1272) <= layer0_outputs(4782);
    layer1_outputs(1273) <= not((layer0_outputs(3896)) or (layer0_outputs(1172)));
    layer1_outputs(1274) <= (layer0_outputs(4160)) and not (layer0_outputs(2884));
    layer1_outputs(1275) <= layer0_outputs(2874);
    layer1_outputs(1276) <= (layer0_outputs(2910)) and not (layer0_outputs(4555));
    layer1_outputs(1277) <= (layer0_outputs(352)) and not (layer0_outputs(5003));
    layer1_outputs(1278) <= '0';
    layer1_outputs(1279) <= not(layer0_outputs(3618));
    layer1_outputs(1280) <= (layer0_outputs(4998)) and (layer0_outputs(1464));
    layer1_outputs(1281) <= not((layer0_outputs(2802)) and (layer0_outputs(1550)));
    layer1_outputs(1282) <= (layer0_outputs(4700)) and not (layer0_outputs(12));
    layer1_outputs(1283) <= (layer0_outputs(4711)) and not (layer0_outputs(2042));
    layer1_outputs(1284) <= '1';
    layer1_outputs(1285) <= layer0_outputs(3612);
    layer1_outputs(1286) <= (layer0_outputs(1201)) and not (layer0_outputs(1758));
    layer1_outputs(1287) <= not(layer0_outputs(5002)) or (layer0_outputs(3712));
    layer1_outputs(1288) <= not(layer0_outputs(3858));
    layer1_outputs(1289) <= not(layer0_outputs(1077)) or (layer0_outputs(5001));
    layer1_outputs(1290) <= (layer0_outputs(1146)) or (layer0_outputs(1506));
    layer1_outputs(1291) <= not(layer0_outputs(2626));
    layer1_outputs(1292) <= (layer0_outputs(3085)) and not (layer0_outputs(3223));
    layer1_outputs(1293) <= '1';
    layer1_outputs(1294) <= not(layer0_outputs(2482)) or (layer0_outputs(1549));
    layer1_outputs(1295) <= not(layer0_outputs(3742)) or (layer0_outputs(3772));
    layer1_outputs(1296) <= (layer0_outputs(1795)) and not (layer0_outputs(3402));
    layer1_outputs(1297) <= not((layer0_outputs(477)) and (layer0_outputs(3156)));
    layer1_outputs(1298) <= '0';
    layer1_outputs(1299) <= not((layer0_outputs(1112)) and (layer0_outputs(4279)));
    layer1_outputs(1300) <= not(layer0_outputs(3686)) or (layer0_outputs(410));
    layer1_outputs(1301) <= (layer0_outputs(2550)) and not (layer0_outputs(1024));
    layer1_outputs(1302) <= not(layer0_outputs(1488));
    layer1_outputs(1303) <= not((layer0_outputs(3857)) or (layer0_outputs(2383)));
    layer1_outputs(1304) <= not((layer0_outputs(5008)) and (layer0_outputs(223)));
    layer1_outputs(1305) <= layer0_outputs(1466);
    layer1_outputs(1306) <= not(layer0_outputs(2962)) or (layer0_outputs(3405));
    layer1_outputs(1307) <= not(layer0_outputs(2243));
    layer1_outputs(1308) <= (layer0_outputs(733)) or (layer0_outputs(3567));
    layer1_outputs(1309) <= '0';
    layer1_outputs(1310) <= '0';
    layer1_outputs(1311) <= not(layer0_outputs(3267));
    layer1_outputs(1312) <= (layer0_outputs(2108)) and (layer0_outputs(1542));
    layer1_outputs(1313) <= '0';
    layer1_outputs(1314) <= (layer0_outputs(4003)) or (layer0_outputs(3251));
    layer1_outputs(1315) <= (layer0_outputs(1925)) and (layer0_outputs(868));
    layer1_outputs(1316) <= not(layer0_outputs(3737));
    layer1_outputs(1317) <= (layer0_outputs(1577)) or (layer0_outputs(822));
    layer1_outputs(1318) <= (layer0_outputs(3779)) or (layer0_outputs(2184));
    layer1_outputs(1319) <= layer0_outputs(134);
    layer1_outputs(1320) <= not(layer0_outputs(2789));
    layer1_outputs(1321) <= not(layer0_outputs(4785));
    layer1_outputs(1322) <= not(layer0_outputs(382));
    layer1_outputs(1323) <= not((layer0_outputs(1788)) or (layer0_outputs(3934)));
    layer1_outputs(1324) <= '1';
    layer1_outputs(1325) <= layer0_outputs(4399);
    layer1_outputs(1326) <= (layer0_outputs(1681)) or (layer0_outputs(630));
    layer1_outputs(1327) <= '0';
    layer1_outputs(1328) <= not(layer0_outputs(3995));
    layer1_outputs(1329) <= not((layer0_outputs(3155)) or (layer0_outputs(1432)));
    layer1_outputs(1330) <= (layer0_outputs(2070)) and not (layer0_outputs(4133));
    layer1_outputs(1331) <= not(layer0_outputs(4107));
    layer1_outputs(1332) <= layer0_outputs(46);
    layer1_outputs(1333) <= layer0_outputs(1694);
    layer1_outputs(1334) <= (layer0_outputs(1046)) or (layer0_outputs(2833));
    layer1_outputs(1335) <= '0';
    layer1_outputs(1336) <= '0';
    layer1_outputs(1337) <= not((layer0_outputs(2012)) and (layer0_outputs(1567)));
    layer1_outputs(1338) <= not((layer0_outputs(267)) and (layer0_outputs(2687)));
    layer1_outputs(1339) <= '1';
    layer1_outputs(1340) <= '1';
    layer1_outputs(1341) <= layer0_outputs(2323);
    layer1_outputs(1342) <= '1';
    layer1_outputs(1343) <= layer0_outputs(3024);
    layer1_outputs(1344) <= layer0_outputs(2680);
    layer1_outputs(1345) <= (layer0_outputs(4217)) or (layer0_outputs(895));
    layer1_outputs(1346) <= not(layer0_outputs(2142)) or (layer0_outputs(2221));
    layer1_outputs(1347) <= '1';
    layer1_outputs(1348) <= '0';
    layer1_outputs(1349) <= (layer0_outputs(1442)) and not (layer0_outputs(489));
    layer1_outputs(1350) <= (layer0_outputs(4912)) and (layer0_outputs(3981));
    layer1_outputs(1351) <= '0';
    layer1_outputs(1352) <= (layer0_outputs(4092)) and not (layer0_outputs(2829));
    layer1_outputs(1353) <= '1';
    layer1_outputs(1354) <= '0';
    layer1_outputs(1355) <= (layer0_outputs(3900)) or (layer0_outputs(2572));
    layer1_outputs(1356) <= '1';
    layer1_outputs(1357) <= not(layer0_outputs(1607)) or (layer0_outputs(173));
    layer1_outputs(1358) <= not((layer0_outputs(3389)) or (layer0_outputs(3066)));
    layer1_outputs(1359) <= (layer0_outputs(4401)) and not (layer0_outputs(611));
    layer1_outputs(1360) <= not((layer0_outputs(1123)) or (layer0_outputs(679)));
    layer1_outputs(1361) <= layer0_outputs(323);
    layer1_outputs(1362) <= layer0_outputs(3951);
    layer1_outputs(1363) <= (layer0_outputs(2805)) and not (layer0_outputs(2110));
    layer1_outputs(1364) <= layer0_outputs(519);
    layer1_outputs(1365) <= (layer0_outputs(12)) and not (layer0_outputs(2360));
    layer1_outputs(1366) <= not(layer0_outputs(4120)) or (layer0_outputs(3805));
    layer1_outputs(1367) <= '1';
    layer1_outputs(1368) <= (layer0_outputs(1228)) and not (layer0_outputs(909));
    layer1_outputs(1369) <= not(layer0_outputs(384)) or (layer0_outputs(337));
    layer1_outputs(1370) <= layer0_outputs(1324);
    layer1_outputs(1371) <= layer0_outputs(624);
    layer1_outputs(1372) <= (layer0_outputs(2617)) and not (layer0_outputs(1989));
    layer1_outputs(1373) <= '1';
    layer1_outputs(1374) <= layer0_outputs(1114);
    layer1_outputs(1375) <= (layer0_outputs(145)) and not (layer0_outputs(1215));
    layer1_outputs(1376) <= layer0_outputs(1512);
    layer1_outputs(1377) <= (layer0_outputs(554)) and not (layer0_outputs(4861));
    layer1_outputs(1378) <= '1';
    layer1_outputs(1379) <= not((layer0_outputs(286)) and (layer0_outputs(3498)));
    layer1_outputs(1380) <= not(layer0_outputs(3671)) or (layer0_outputs(2236));
    layer1_outputs(1381) <= '0';
    layer1_outputs(1382) <= not((layer0_outputs(1010)) or (layer0_outputs(4300)));
    layer1_outputs(1383) <= (layer0_outputs(2237)) and not (layer0_outputs(4376));
    layer1_outputs(1384) <= (layer0_outputs(2901)) and not (layer0_outputs(3148));
    layer1_outputs(1385) <= not((layer0_outputs(1010)) or (layer0_outputs(1099)));
    layer1_outputs(1386) <= layer0_outputs(3224);
    layer1_outputs(1387) <= not(layer0_outputs(248)) or (layer0_outputs(2742));
    layer1_outputs(1388) <= (layer0_outputs(1188)) or (layer0_outputs(4480));
    layer1_outputs(1389) <= layer0_outputs(3507);
    layer1_outputs(1390) <= not(layer0_outputs(1989)) or (layer0_outputs(2811));
    layer1_outputs(1391) <= '1';
    layer1_outputs(1392) <= (layer0_outputs(3488)) and not (layer0_outputs(3144));
    layer1_outputs(1393) <= (layer0_outputs(3582)) and not (layer0_outputs(1135));
    layer1_outputs(1394) <= not((layer0_outputs(2281)) and (layer0_outputs(3469)));
    layer1_outputs(1395) <= '1';
    layer1_outputs(1396) <= (layer0_outputs(1311)) and not (layer0_outputs(2397));
    layer1_outputs(1397) <= layer0_outputs(4644);
    layer1_outputs(1398) <= '1';
    layer1_outputs(1399) <= '1';
    layer1_outputs(1400) <= '1';
    layer1_outputs(1401) <= not((layer0_outputs(385)) or (layer0_outputs(2039)));
    layer1_outputs(1402) <= not(layer0_outputs(4572)) or (layer0_outputs(418));
    layer1_outputs(1403) <= (layer0_outputs(4526)) or (layer0_outputs(690));
    layer1_outputs(1404) <= '0';
    layer1_outputs(1405) <= not(layer0_outputs(3254));
    layer1_outputs(1406) <= not((layer0_outputs(4185)) or (layer0_outputs(795)));
    layer1_outputs(1407) <= (layer0_outputs(1396)) and not (layer0_outputs(2786));
    layer1_outputs(1408) <= '0';
    layer1_outputs(1409) <= '1';
    layer1_outputs(1410) <= (layer0_outputs(4974)) and not (layer0_outputs(4077));
    layer1_outputs(1411) <= layer0_outputs(4138);
    layer1_outputs(1412) <= (layer0_outputs(317)) and not (layer0_outputs(2757));
    layer1_outputs(1413) <= (layer0_outputs(3962)) or (layer0_outputs(4454));
    layer1_outputs(1414) <= (layer0_outputs(1715)) or (layer0_outputs(5052));
    layer1_outputs(1415) <= (layer0_outputs(2016)) and not (layer0_outputs(2264));
    layer1_outputs(1416) <= not(layer0_outputs(2694));
    layer1_outputs(1417) <= '0';
    layer1_outputs(1418) <= layer0_outputs(3460);
    layer1_outputs(1419) <= '1';
    layer1_outputs(1420) <= not((layer0_outputs(263)) and (layer0_outputs(976)));
    layer1_outputs(1421) <= not(layer0_outputs(1332)) or (layer0_outputs(2375));
    layer1_outputs(1422) <= not(layer0_outputs(4226));
    layer1_outputs(1423) <= '0';
    layer1_outputs(1424) <= '1';
    layer1_outputs(1425) <= '1';
    layer1_outputs(1426) <= layer0_outputs(4106);
    layer1_outputs(1427) <= not(layer0_outputs(693)) or (layer0_outputs(5014));
    layer1_outputs(1428) <= (layer0_outputs(3311)) and not (layer0_outputs(564));
    layer1_outputs(1429) <= not(layer0_outputs(1160)) or (layer0_outputs(4467));
    layer1_outputs(1430) <= (layer0_outputs(4591)) or (layer0_outputs(3540));
    layer1_outputs(1431) <= '0';
    layer1_outputs(1432) <= (layer0_outputs(3280)) and (layer0_outputs(435));
    layer1_outputs(1433) <= not(layer0_outputs(4381)) or (layer0_outputs(2826));
    layer1_outputs(1434) <= '1';
    layer1_outputs(1435) <= not((layer0_outputs(2895)) or (layer0_outputs(3131)));
    layer1_outputs(1436) <= '0';
    layer1_outputs(1437) <= (layer0_outputs(2134)) or (layer0_outputs(2875));
    layer1_outputs(1438) <= layer0_outputs(3063);
    layer1_outputs(1439) <= '1';
    layer1_outputs(1440) <= '1';
    layer1_outputs(1441) <= (layer0_outputs(2964)) and (layer0_outputs(1314));
    layer1_outputs(1442) <= (layer0_outputs(3952)) and not (layer0_outputs(2160));
    layer1_outputs(1443) <= (layer0_outputs(3763)) and (layer0_outputs(1309));
    layer1_outputs(1444) <= '1';
    layer1_outputs(1445) <= not(layer0_outputs(1272));
    layer1_outputs(1446) <= (layer0_outputs(278)) or (layer0_outputs(1620));
    layer1_outputs(1447) <= '0';
    layer1_outputs(1448) <= (layer0_outputs(3171)) and not (layer0_outputs(2423));
    layer1_outputs(1449) <= (layer0_outputs(2650)) and not (layer0_outputs(1170));
    layer1_outputs(1450) <= (layer0_outputs(2358)) and not (layer0_outputs(2806));
    layer1_outputs(1451) <= '0';
    layer1_outputs(1452) <= '0';
    layer1_outputs(1453) <= (layer0_outputs(3089)) and (layer0_outputs(2791));
    layer1_outputs(1454) <= (layer0_outputs(3450)) or (layer0_outputs(4751));
    layer1_outputs(1455) <= (layer0_outputs(1645)) and (layer0_outputs(4445));
    layer1_outputs(1456) <= (layer0_outputs(2915)) and not (layer0_outputs(601));
    layer1_outputs(1457) <= '1';
    layer1_outputs(1458) <= (layer0_outputs(553)) and (layer0_outputs(4079));
    layer1_outputs(1459) <= not(layer0_outputs(364)) or (layer0_outputs(1954));
    layer1_outputs(1460) <= not((layer0_outputs(3747)) and (layer0_outputs(4900)));
    layer1_outputs(1461) <= not((layer0_outputs(4102)) and (layer0_outputs(155)));
    layer1_outputs(1462) <= (layer0_outputs(1019)) and (layer0_outputs(4349));
    layer1_outputs(1463) <= not((layer0_outputs(3262)) and (layer0_outputs(3878)));
    layer1_outputs(1464) <= (layer0_outputs(242)) or (layer0_outputs(708));
    layer1_outputs(1465) <= '0';
    layer1_outputs(1466) <= (layer0_outputs(332)) and not (layer0_outputs(559));
    layer1_outputs(1467) <= layer0_outputs(3911);
    layer1_outputs(1468) <= (layer0_outputs(1623)) and not (layer0_outputs(4060));
    layer1_outputs(1469) <= not(layer0_outputs(2767)) or (layer0_outputs(4473));
    layer1_outputs(1470) <= (layer0_outputs(4159)) xor (layer0_outputs(3171));
    layer1_outputs(1471) <= not((layer0_outputs(1171)) or (layer0_outputs(4429)));
    layer1_outputs(1472) <= not(layer0_outputs(1245)) or (layer0_outputs(2499));
    layer1_outputs(1473) <= not((layer0_outputs(2588)) or (layer0_outputs(4207)));
    layer1_outputs(1474) <= not(layer0_outputs(4847));
    layer1_outputs(1475) <= (layer0_outputs(985)) or (layer0_outputs(476));
    layer1_outputs(1476) <= not((layer0_outputs(3266)) or (layer0_outputs(1328)));
    layer1_outputs(1477) <= (layer0_outputs(4357)) and not (layer0_outputs(3209));
    layer1_outputs(1478) <= (layer0_outputs(1118)) and not (layer0_outputs(3680));
    layer1_outputs(1479) <= not(layer0_outputs(3133));
    layer1_outputs(1480) <= '1';
    layer1_outputs(1481) <= layer0_outputs(4677);
    layer1_outputs(1482) <= (layer0_outputs(482)) and not (layer0_outputs(2776));
    layer1_outputs(1483) <= layer0_outputs(2652);
    layer1_outputs(1484) <= '0';
    layer1_outputs(1485) <= '0';
    layer1_outputs(1486) <= (layer0_outputs(3912)) and not (layer0_outputs(2730));
    layer1_outputs(1487) <= (layer0_outputs(3084)) or (layer0_outputs(2079));
    layer1_outputs(1488) <= not(layer0_outputs(475)) or (layer0_outputs(3214));
    layer1_outputs(1489) <= (layer0_outputs(4653)) and not (layer0_outputs(3708));
    layer1_outputs(1490) <= not(layer0_outputs(3667));
    layer1_outputs(1491) <= (layer0_outputs(593)) and not (layer0_outputs(559));
    layer1_outputs(1492) <= not((layer0_outputs(2518)) and (layer0_outputs(2040)));
    layer1_outputs(1493) <= (layer0_outputs(2641)) or (layer0_outputs(2402));
    layer1_outputs(1494) <= (layer0_outputs(1452)) and not (layer0_outputs(2899));
    layer1_outputs(1495) <= not(layer0_outputs(513));
    layer1_outputs(1496) <= (layer0_outputs(1277)) and (layer0_outputs(3809));
    layer1_outputs(1497) <= '1';
    layer1_outputs(1498) <= not(layer0_outputs(2959)) or (layer0_outputs(1560));
    layer1_outputs(1499) <= '0';
    layer1_outputs(1500) <= '1';
    layer1_outputs(1501) <= (layer0_outputs(4196)) and not (layer0_outputs(4958));
    layer1_outputs(1502) <= not(layer0_outputs(3569)) or (layer0_outputs(3972));
    layer1_outputs(1503) <= '0';
    layer1_outputs(1504) <= not((layer0_outputs(1938)) and (layer0_outputs(718)));
    layer1_outputs(1505) <= '0';
    layer1_outputs(1506) <= layer0_outputs(2072);
    layer1_outputs(1507) <= layer0_outputs(1647);
    layer1_outputs(1508) <= not(layer0_outputs(3424)) or (layer0_outputs(1825));
    layer1_outputs(1509) <= layer0_outputs(1591);
    layer1_outputs(1510) <= (layer0_outputs(4010)) and not (layer0_outputs(4189));
    layer1_outputs(1511) <= '0';
    layer1_outputs(1512) <= (layer0_outputs(1294)) xor (layer0_outputs(1513));
    layer1_outputs(1513) <= layer0_outputs(4656);
    layer1_outputs(1514) <= not((layer0_outputs(3182)) and (layer0_outputs(1091)));
    layer1_outputs(1515) <= layer0_outputs(1838);
    layer1_outputs(1516) <= '0';
    layer1_outputs(1517) <= (layer0_outputs(4621)) and (layer0_outputs(1346));
    layer1_outputs(1518) <= (layer0_outputs(3953)) and not (layer0_outputs(4767));
    layer1_outputs(1519) <= not((layer0_outputs(48)) and (layer0_outputs(1199)));
    layer1_outputs(1520) <= (layer0_outputs(2311)) or (layer0_outputs(1875));
    layer1_outputs(1521) <= not((layer0_outputs(3533)) and (layer0_outputs(2718)));
    layer1_outputs(1522) <= '0';
    layer1_outputs(1523) <= not((layer0_outputs(1274)) or (layer0_outputs(74)));
    layer1_outputs(1524) <= layer0_outputs(274);
    layer1_outputs(1525) <= (layer0_outputs(2254)) and not (layer0_outputs(2521));
    layer1_outputs(1526) <= '1';
    layer1_outputs(1527) <= layer0_outputs(1571);
    layer1_outputs(1528) <= '1';
    layer1_outputs(1529) <= not(layer0_outputs(2947));
    layer1_outputs(1530) <= not(layer0_outputs(2510)) or (layer0_outputs(3625));
    layer1_outputs(1531) <= '1';
    layer1_outputs(1532) <= layer0_outputs(850);
    layer1_outputs(1533) <= '1';
    layer1_outputs(1534) <= not((layer0_outputs(3922)) and (layer0_outputs(1068)));
    layer1_outputs(1535) <= not(layer0_outputs(1096)) or (layer0_outputs(2419));
    layer1_outputs(1536) <= layer0_outputs(1569);
    layer1_outputs(1537) <= not(layer0_outputs(1494));
    layer1_outputs(1538) <= (layer0_outputs(4975)) and not (layer0_outputs(573));
    layer1_outputs(1539) <= '1';
    layer1_outputs(1540) <= not((layer0_outputs(1474)) and (layer0_outputs(2388)));
    layer1_outputs(1541) <= not((layer0_outputs(2115)) or (layer0_outputs(2647)));
    layer1_outputs(1542) <= '0';
    layer1_outputs(1543) <= (layer0_outputs(2969)) and not (layer0_outputs(59));
    layer1_outputs(1544) <= (layer0_outputs(2568)) xor (layer0_outputs(923));
    layer1_outputs(1545) <= not(layer0_outputs(103));
    layer1_outputs(1546) <= (layer0_outputs(4135)) or (layer0_outputs(1804));
    layer1_outputs(1547) <= '1';
    layer1_outputs(1548) <= (layer0_outputs(5026)) and (layer0_outputs(4311));
    layer1_outputs(1549) <= not((layer0_outputs(1125)) or (layer0_outputs(2608)));
    layer1_outputs(1550) <= not((layer0_outputs(3153)) and (layer0_outputs(3621)));
    layer1_outputs(1551) <= not((layer0_outputs(580)) or (layer0_outputs(3100)));
    layer1_outputs(1552) <= '1';
    layer1_outputs(1553) <= '1';
    layer1_outputs(1554) <= layer0_outputs(3375);
    layer1_outputs(1555) <= '1';
    layer1_outputs(1556) <= '0';
    layer1_outputs(1557) <= not((layer0_outputs(4366)) or (layer0_outputs(4056)));
    layer1_outputs(1558) <= not((layer0_outputs(2125)) and (layer0_outputs(3520)));
    layer1_outputs(1559) <= (layer0_outputs(2044)) and not (layer0_outputs(4788));
    layer1_outputs(1560) <= (layer0_outputs(4382)) and not (layer0_outputs(3625));
    layer1_outputs(1561) <= not((layer0_outputs(2614)) or (layer0_outputs(1323)));
    layer1_outputs(1562) <= '0';
    layer1_outputs(1563) <= '1';
    layer1_outputs(1564) <= '1';
    layer1_outputs(1565) <= layer0_outputs(434);
    layer1_outputs(1566) <= not(layer0_outputs(472));
    layer1_outputs(1567) <= (layer0_outputs(641)) and not (layer0_outputs(262));
    layer1_outputs(1568) <= not((layer0_outputs(1574)) and (layer0_outputs(4210)));
    layer1_outputs(1569) <= '1';
    layer1_outputs(1570) <= '0';
    layer1_outputs(1571) <= (layer0_outputs(368)) and not (layer0_outputs(315));
    layer1_outputs(1572) <= '0';
    layer1_outputs(1573) <= '0';
    layer1_outputs(1574) <= '0';
    layer1_outputs(1575) <= (layer0_outputs(5076)) and (layer0_outputs(4896));
    layer1_outputs(1576) <= not((layer0_outputs(4024)) or (layer0_outputs(3815)));
    layer1_outputs(1577) <= not(layer0_outputs(302)) or (layer0_outputs(3186));
    layer1_outputs(1578) <= layer0_outputs(2800);
    layer1_outputs(1579) <= '1';
    layer1_outputs(1580) <= '0';
    layer1_outputs(1581) <= not(layer0_outputs(4357));
    layer1_outputs(1582) <= '1';
    layer1_outputs(1583) <= not(layer0_outputs(661));
    layer1_outputs(1584) <= not(layer0_outputs(1691)) or (layer0_outputs(4781));
    layer1_outputs(1585) <= not((layer0_outputs(3734)) and (layer0_outputs(4048)));
    layer1_outputs(1586) <= not(layer0_outputs(3454)) or (layer0_outputs(1059));
    layer1_outputs(1587) <= not(layer0_outputs(4065)) or (layer0_outputs(703));
    layer1_outputs(1588) <= (layer0_outputs(3997)) or (layer0_outputs(4901));
    layer1_outputs(1589) <= not(layer0_outputs(699)) or (layer0_outputs(1748));
    layer1_outputs(1590) <= layer0_outputs(4444);
    layer1_outputs(1591) <= not(layer0_outputs(4695)) or (layer0_outputs(4807));
    layer1_outputs(1592) <= not((layer0_outputs(2402)) and (layer0_outputs(727)));
    layer1_outputs(1593) <= (layer0_outputs(3831)) or (layer0_outputs(2234));
    layer1_outputs(1594) <= not(layer0_outputs(1531));
    layer1_outputs(1595) <= not((layer0_outputs(2514)) or (layer0_outputs(4564)));
    layer1_outputs(1596) <= not(layer0_outputs(87)) or (layer0_outputs(1389));
    layer1_outputs(1597) <= '0';
    layer1_outputs(1598) <= (layer0_outputs(2233)) or (layer0_outputs(1517));
    layer1_outputs(1599) <= '0';
    layer1_outputs(1600) <= (layer0_outputs(4419)) or (layer0_outputs(1455));
    layer1_outputs(1601) <= '1';
    layer1_outputs(1602) <= not(layer0_outputs(2504)) or (layer0_outputs(2208));
    layer1_outputs(1603) <= not((layer0_outputs(3430)) and (layer0_outputs(1981)));
    layer1_outputs(1604) <= not((layer0_outputs(1306)) or (layer0_outputs(3030)));
    layer1_outputs(1605) <= (layer0_outputs(764)) and not (layer0_outputs(919));
    layer1_outputs(1606) <= not((layer0_outputs(4511)) and (layer0_outputs(1994)));
    layer1_outputs(1607) <= not(layer0_outputs(2618)) or (layer0_outputs(2980));
    layer1_outputs(1608) <= not((layer0_outputs(3552)) xor (layer0_outputs(4371)));
    layer1_outputs(1609) <= (layer0_outputs(4225)) and not (layer0_outputs(2367));
    layer1_outputs(1610) <= '1';
    layer1_outputs(1611) <= '0';
    layer1_outputs(1612) <= (layer0_outputs(1348)) and (layer0_outputs(3520));
    layer1_outputs(1613) <= (layer0_outputs(3033)) and not (layer0_outputs(4076));
    layer1_outputs(1614) <= '0';
    layer1_outputs(1615) <= '1';
    layer1_outputs(1616) <= not((layer0_outputs(3143)) and (layer0_outputs(3368)));
    layer1_outputs(1617) <= layer0_outputs(963);
    layer1_outputs(1618) <= not((layer0_outputs(4742)) and (layer0_outputs(5014)));
    layer1_outputs(1619) <= not(layer0_outputs(2901));
    layer1_outputs(1620) <= '0';
    layer1_outputs(1621) <= '1';
    layer1_outputs(1622) <= layer0_outputs(143);
    layer1_outputs(1623) <= '0';
    layer1_outputs(1624) <= '0';
    layer1_outputs(1625) <= '0';
    layer1_outputs(1626) <= not((layer0_outputs(356)) or (layer0_outputs(4904)));
    layer1_outputs(1627) <= '0';
    layer1_outputs(1628) <= '1';
    layer1_outputs(1629) <= (layer0_outputs(1507)) and (layer0_outputs(3410));
    layer1_outputs(1630) <= not((layer0_outputs(4965)) or (layer0_outputs(4212)));
    layer1_outputs(1631) <= (layer0_outputs(4177)) and not (layer0_outputs(3270));
    layer1_outputs(1632) <= not((layer0_outputs(530)) or (layer0_outputs(2157)));
    layer1_outputs(1633) <= '1';
    layer1_outputs(1634) <= layer0_outputs(1423);
    layer1_outputs(1635) <= (layer0_outputs(3966)) and not (layer0_outputs(4544));
    layer1_outputs(1636) <= layer0_outputs(2611);
    layer1_outputs(1637) <= layer0_outputs(4163);
    layer1_outputs(1638) <= not(layer0_outputs(817)) or (layer0_outputs(5081));
    layer1_outputs(1639) <= layer0_outputs(3107);
    layer1_outputs(1640) <= '0';
    layer1_outputs(1641) <= not((layer0_outputs(2097)) or (layer0_outputs(402)));
    layer1_outputs(1642) <= (layer0_outputs(3281)) and (layer0_outputs(3703));
    layer1_outputs(1643) <= (layer0_outputs(3342)) and not (layer0_outputs(2808));
    layer1_outputs(1644) <= '1';
    layer1_outputs(1645) <= not(layer0_outputs(266)) or (layer0_outputs(1883));
    layer1_outputs(1646) <= '1';
    layer1_outputs(1647) <= not((layer0_outputs(1288)) and (layer0_outputs(403)));
    layer1_outputs(1648) <= (layer0_outputs(3991)) and not (layer0_outputs(1425));
    layer1_outputs(1649) <= (layer0_outputs(581)) and (layer0_outputs(3534));
    layer1_outputs(1650) <= layer0_outputs(537);
    layer1_outputs(1651) <= '1';
    layer1_outputs(1652) <= '1';
    layer1_outputs(1653) <= (layer0_outputs(4978)) and (layer0_outputs(421));
    layer1_outputs(1654) <= (layer0_outputs(4685)) or (layer0_outputs(1767));
    layer1_outputs(1655) <= not(layer0_outputs(1227)) or (layer0_outputs(4541));
    layer1_outputs(1656) <= not((layer0_outputs(3063)) or (layer0_outputs(3134)));
    layer1_outputs(1657) <= not(layer0_outputs(136));
    layer1_outputs(1658) <= layer0_outputs(2673);
    layer1_outputs(1659) <= '1';
    layer1_outputs(1660) <= '0';
    layer1_outputs(1661) <= (layer0_outputs(4649)) and not (layer0_outputs(4795));
    layer1_outputs(1662) <= not(layer0_outputs(776)) or (layer0_outputs(904));
    layer1_outputs(1663) <= not(layer0_outputs(2128)) or (layer0_outputs(2051));
    layer1_outputs(1664) <= not(layer0_outputs(2535)) or (layer0_outputs(2338));
    layer1_outputs(1665) <= (layer0_outputs(2970)) and not (layer0_outputs(1615));
    layer1_outputs(1666) <= not(layer0_outputs(2197));
    layer1_outputs(1667) <= (layer0_outputs(3981)) xor (layer0_outputs(687));
    layer1_outputs(1668) <= (layer0_outputs(2971)) and not (layer0_outputs(1626));
    layer1_outputs(1669) <= (layer0_outputs(710)) and (layer0_outputs(1317));
    layer1_outputs(1670) <= (layer0_outputs(617)) or (layer0_outputs(3589));
    layer1_outputs(1671) <= not(layer0_outputs(2816)) or (layer0_outputs(2834));
    layer1_outputs(1672) <= not(layer0_outputs(4369));
    layer1_outputs(1673) <= layer0_outputs(4544);
    layer1_outputs(1674) <= not((layer0_outputs(4715)) and (layer0_outputs(369)));
    layer1_outputs(1675) <= not(layer0_outputs(812)) or (layer0_outputs(3092));
    layer1_outputs(1676) <= not((layer0_outputs(3609)) or (layer0_outputs(3395)));
    layer1_outputs(1677) <= '0';
    layer1_outputs(1678) <= not(layer0_outputs(3242));
    layer1_outputs(1679) <= (layer0_outputs(2685)) and not (layer0_outputs(2061));
    layer1_outputs(1680) <= not((layer0_outputs(529)) or (layer0_outputs(4657)));
    layer1_outputs(1681) <= '1';
    layer1_outputs(1682) <= layer0_outputs(1957);
    layer1_outputs(1683) <= '1';
    layer1_outputs(1684) <= not(layer0_outputs(729)) or (layer0_outputs(4426));
    layer1_outputs(1685) <= not(layer0_outputs(506)) or (layer0_outputs(2926));
    layer1_outputs(1686) <= layer0_outputs(620);
    layer1_outputs(1687) <= (layer0_outputs(4533)) and (layer0_outputs(1760));
    layer1_outputs(1688) <= '0';
    layer1_outputs(1689) <= '1';
    layer1_outputs(1690) <= not(layer0_outputs(826)) or (layer0_outputs(5078));
    layer1_outputs(1691) <= not(layer0_outputs(4558)) or (layer0_outputs(3112));
    layer1_outputs(1692) <= layer0_outputs(3100);
    layer1_outputs(1693) <= '0';
    layer1_outputs(1694) <= layer0_outputs(4045);
    layer1_outputs(1695) <= '1';
    layer1_outputs(1696) <= '0';
    layer1_outputs(1697) <= '0';
    layer1_outputs(1698) <= layer0_outputs(4894);
    layer1_outputs(1699) <= layer0_outputs(4047);
    layer1_outputs(1700) <= not((layer0_outputs(4844)) and (layer0_outputs(397)));
    layer1_outputs(1701) <= '0';
    layer1_outputs(1702) <= '1';
    layer1_outputs(1703) <= (layer0_outputs(4972)) or (layer0_outputs(4617));
    layer1_outputs(1704) <= '1';
    layer1_outputs(1705) <= '1';
    layer1_outputs(1706) <= '0';
    layer1_outputs(1707) <= (layer0_outputs(3812)) or (layer0_outputs(3428));
    layer1_outputs(1708) <= '0';
    layer1_outputs(1709) <= '0';
    layer1_outputs(1710) <= not(layer0_outputs(48));
    layer1_outputs(1711) <= not((layer0_outputs(2188)) or (layer0_outputs(427)));
    layer1_outputs(1712) <= (layer0_outputs(136)) and not (layer0_outputs(1794));
    layer1_outputs(1713) <= not(layer0_outputs(3538)) or (layer0_outputs(1866));
    layer1_outputs(1714) <= not(layer0_outputs(422));
    layer1_outputs(1715) <= not(layer0_outputs(2816)) or (layer0_outputs(2597));
    layer1_outputs(1716) <= (layer0_outputs(3984)) and not (layer0_outputs(2292));
    layer1_outputs(1717) <= '0';
    layer1_outputs(1718) <= '1';
    layer1_outputs(1719) <= not(layer0_outputs(4542)) or (layer0_outputs(4470));
    layer1_outputs(1720) <= '1';
    layer1_outputs(1721) <= '0';
    layer1_outputs(1722) <= not((layer0_outputs(3933)) and (layer0_outputs(2785)));
    layer1_outputs(1723) <= not((layer0_outputs(4273)) or (layer0_outputs(2542)));
    layer1_outputs(1724) <= (layer0_outputs(2411)) and not (layer0_outputs(3740));
    layer1_outputs(1725) <= '1';
    layer1_outputs(1726) <= not((layer0_outputs(4934)) or (layer0_outputs(289)));
    layer1_outputs(1727) <= not(layer0_outputs(4446));
    layer1_outputs(1728) <= '0';
    layer1_outputs(1729) <= '1';
    layer1_outputs(1730) <= (layer0_outputs(4868)) and not (layer0_outputs(931));
    layer1_outputs(1731) <= '0';
    layer1_outputs(1732) <= not(layer0_outputs(17));
    layer1_outputs(1733) <= '0';
    layer1_outputs(1734) <= not((layer0_outputs(246)) or (layer0_outputs(4726)));
    layer1_outputs(1735) <= '1';
    layer1_outputs(1736) <= not(layer0_outputs(4753)) or (layer0_outputs(197));
    layer1_outputs(1737) <= (layer0_outputs(1480)) and not (layer0_outputs(567));
    layer1_outputs(1738) <= (layer0_outputs(266)) and (layer0_outputs(3074));
    layer1_outputs(1739) <= layer0_outputs(4680);
    layer1_outputs(1740) <= layer0_outputs(1502);
    layer1_outputs(1741) <= (layer0_outputs(2441)) and (layer0_outputs(3745));
    layer1_outputs(1742) <= not(layer0_outputs(1284));
    layer1_outputs(1743) <= not((layer0_outputs(4559)) and (layer0_outputs(1624)));
    layer1_outputs(1744) <= '0';
    layer1_outputs(1745) <= not(layer0_outputs(4513));
    layer1_outputs(1746) <= not((layer0_outputs(633)) and (layer0_outputs(3230)));
    layer1_outputs(1747) <= '1';
    layer1_outputs(1748) <= not(layer0_outputs(314));
    layer1_outputs(1749) <= not(layer0_outputs(2179)) or (layer0_outputs(2099));
    layer1_outputs(1750) <= not(layer0_outputs(659));
    layer1_outputs(1751) <= (layer0_outputs(1907)) or (layer0_outputs(5045));
    layer1_outputs(1752) <= '0';
    layer1_outputs(1753) <= not(layer0_outputs(3164)) or (layer0_outputs(4483));
    layer1_outputs(1754) <= '0';
    layer1_outputs(1755) <= not(layer0_outputs(4465)) or (layer0_outputs(3343));
    layer1_outputs(1756) <= (layer0_outputs(1066)) or (layer0_outputs(4295));
    layer1_outputs(1757) <= (layer0_outputs(1953)) and not (layer0_outputs(1176));
    layer1_outputs(1758) <= not(layer0_outputs(2268)) or (layer0_outputs(3197));
    layer1_outputs(1759) <= '0';
    layer1_outputs(1760) <= layer0_outputs(1898);
    layer1_outputs(1761) <= not(layer0_outputs(3720));
    layer1_outputs(1762) <= layer0_outputs(329);
    layer1_outputs(1763) <= not((layer0_outputs(907)) or (layer0_outputs(1909)));
    layer1_outputs(1764) <= (layer0_outputs(1540)) and (layer0_outputs(599));
    layer1_outputs(1765) <= layer0_outputs(25);
    layer1_outputs(1766) <= '1';
    layer1_outputs(1767) <= not((layer0_outputs(2691)) xor (layer0_outputs(1262)));
    layer1_outputs(1768) <= (layer0_outputs(1095)) and not (layer0_outputs(2063));
    layer1_outputs(1769) <= '1';
    layer1_outputs(1770) <= not(layer0_outputs(1534)) or (layer0_outputs(199));
    layer1_outputs(1771) <= not((layer0_outputs(3927)) and (layer0_outputs(5098)));
    layer1_outputs(1772) <= not(layer0_outputs(1006)) or (layer0_outputs(2194));
    layer1_outputs(1773) <= '1';
    layer1_outputs(1774) <= '0';
    layer1_outputs(1775) <= '0';
    layer1_outputs(1776) <= not((layer0_outputs(2644)) or (layer0_outputs(731)));
    layer1_outputs(1777) <= not(layer0_outputs(188)) or (layer0_outputs(2052));
    layer1_outputs(1778) <= (layer0_outputs(1666)) and (layer0_outputs(4833));
    layer1_outputs(1779) <= not((layer0_outputs(583)) or (layer0_outputs(3005)));
    layer1_outputs(1780) <= '1';
    layer1_outputs(1781) <= '1';
    layer1_outputs(1782) <= not((layer0_outputs(3277)) or (layer0_outputs(2529)));
    layer1_outputs(1783) <= not(layer0_outputs(1308)) or (layer0_outputs(4235));
    layer1_outputs(1784) <= '0';
    layer1_outputs(1785) <= '1';
    layer1_outputs(1786) <= (layer0_outputs(4425)) and not (layer0_outputs(4629));
    layer1_outputs(1787) <= layer0_outputs(2638);
    layer1_outputs(1788) <= not((layer0_outputs(942)) or (layer0_outputs(970)));
    layer1_outputs(1789) <= (layer0_outputs(3089)) and not (layer0_outputs(1074));
    layer1_outputs(1790) <= not(layer0_outputs(1263));
    layer1_outputs(1791) <= '0';
    layer1_outputs(1792) <= not(layer0_outputs(3292)) or (layer0_outputs(4552));
    layer1_outputs(1793) <= (layer0_outputs(777)) and not (layer0_outputs(3195));
    layer1_outputs(1794) <= '0';
    layer1_outputs(1795) <= (layer0_outputs(4855)) and (layer0_outputs(1617));
    layer1_outputs(1796) <= '0';
    layer1_outputs(1797) <= '1';
    layer1_outputs(1798) <= '1';
    layer1_outputs(1799) <= layer0_outputs(563);
    layer1_outputs(1800) <= (layer0_outputs(4498)) and not (layer0_outputs(686));
    layer1_outputs(1801) <= not(layer0_outputs(3910));
    layer1_outputs(1802) <= '1';
    layer1_outputs(1803) <= (layer0_outputs(4320)) and (layer0_outputs(865));
    layer1_outputs(1804) <= layer0_outputs(2704);
    layer1_outputs(1805) <= '0';
    layer1_outputs(1806) <= (layer0_outputs(3327)) and (layer0_outputs(2147));
    layer1_outputs(1807) <= not((layer0_outputs(2951)) or (layer0_outputs(3108)));
    layer1_outputs(1808) <= not(layer0_outputs(2824));
    layer1_outputs(1809) <= (layer0_outputs(1238)) and not (layer0_outputs(3170));
    layer1_outputs(1810) <= '1';
    layer1_outputs(1811) <= (layer0_outputs(353)) or (layer0_outputs(4258));
    layer1_outputs(1812) <= '1';
    layer1_outputs(1813) <= '0';
    layer1_outputs(1814) <= not((layer0_outputs(1833)) or (layer0_outputs(2923)));
    layer1_outputs(1815) <= layer0_outputs(3682);
    layer1_outputs(1816) <= not((layer0_outputs(114)) or (layer0_outputs(4132)));
    layer1_outputs(1817) <= '0';
    layer1_outputs(1818) <= (layer0_outputs(1161)) and (layer0_outputs(3581));
    layer1_outputs(1819) <= (layer0_outputs(2812)) and (layer0_outputs(1411));
    layer1_outputs(1820) <= not(layer0_outputs(4364)) or (layer0_outputs(1067));
    layer1_outputs(1821) <= not(layer0_outputs(114)) or (layer0_outputs(4068));
    layer1_outputs(1822) <= (layer0_outputs(2591)) and (layer0_outputs(981));
    layer1_outputs(1823) <= (layer0_outputs(1508)) and not (layer0_outputs(3201));
    layer1_outputs(1824) <= not((layer0_outputs(1839)) and (layer0_outputs(3361)));
    layer1_outputs(1825) <= not(layer0_outputs(3956));
    layer1_outputs(1826) <= not(layer0_outputs(4105)) or (layer0_outputs(2778));
    layer1_outputs(1827) <= (layer0_outputs(138)) and not (layer0_outputs(2464));
    layer1_outputs(1828) <= layer0_outputs(3570);
    layer1_outputs(1829) <= not((layer0_outputs(616)) and (layer0_outputs(2665)));
    layer1_outputs(1830) <= (layer0_outputs(2563)) and (layer0_outputs(3266));
    layer1_outputs(1831) <= not((layer0_outputs(4796)) or (layer0_outputs(3717)));
    layer1_outputs(1832) <= not(layer0_outputs(3852)) or (layer0_outputs(355));
    layer1_outputs(1833) <= '0';
    layer1_outputs(1834) <= '0';
    layer1_outputs(1835) <= '1';
    layer1_outputs(1836) <= (layer0_outputs(2217)) or (layer0_outputs(2032));
    layer1_outputs(1837) <= (layer0_outputs(4882)) and not (layer0_outputs(1816));
    layer1_outputs(1838) <= (layer0_outputs(548)) or (layer0_outputs(829));
    layer1_outputs(1839) <= not((layer0_outputs(374)) and (layer0_outputs(1257)));
    layer1_outputs(1840) <= '0';
    layer1_outputs(1841) <= '0';
    layer1_outputs(1842) <= (layer0_outputs(4718)) or (layer0_outputs(4950));
    layer1_outputs(1843) <= not(layer0_outputs(637)) or (layer0_outputs(1175));
    layer1_outputs(1844) <= (layer0_outputs(3698)) and not (layer0_outputs(333));
    layer1_outputs(1845) <= '0';
    layer1_outputs(1846) <= not(layer0_outputs(3821));
    layer1_outputs(1847) <= (layer0_outputs(4041)) or (layer0_outputs(3384));
    layer1_outputs(1848) <= layer0_outputs(3667);
    layer1_outputs(1849) <= not((layer0_outputs(350)) and (layer0_outputs(3536)));
    layer1_outputs(1850) <= not(layer0_outputs(1584));
    layer1_outputs(1851) <= not((layer0_outputs(1590)) and (layer0_outputs(2284)));
    layer1_outputs(1852) <= not(layer0_outputs(1842)) or (layer0_outputs(1686));
    layer1_outputs(1853) <= (layer0_outputs(921)) and not (layer0_outputs(898));
    layer1_outputs(1854) <= (layer0_outputs(399)) and not (layer0_outputs(4212));
    layer1_outputs(1855) <= (layer0_outputs(127)) or (layer0_outputs(2146));
    layer1_outputs(1856) <= layer0_outputs(3572);
    layer1_outputs(1857) <= (layer0_outputs(1859)) and not (layer0_outputs(1310));
    layer1_outputs(1858) <= not(layer0_outputs(4698)) or (layer0_outputs(446));
    layer1_outputs(1859) <= layer0_outputs(4921);
    layer1_outputs(1860) <= not(layer0_outputs(3664)) or (layer0_outputs(2417));
    layer1_outputs(1861) <= layer0_outputs(4124);
    layer1_outputs(1862) <= layer0_outputs(4538);
    layer1_outputs(1863) <= '1';
    layer1_outputs(1864) <= '0';
    layer1_outputs(1865) <= '0';
    layer1_outputs(1866) <= '0';
    layer1_outputs(1867) <= not(layer0_outputs(3642));
    layer1_outputs(1868) <= not(layer0_outputs(4198)) or (layer0_outputs(4681));
    layer1_outputs(1869) <= (layer0_outputs(3465)) and not (layer0_outputs(2282));
    layer1_outputs(1870) <= '1';
    layer1_outputs(1871) <= (layer0_outputs(5119)) and not (layer0_outputs(535));
    layer1_outputs(1872) <= (layer0_outputs(3869)) and not (layer0_outputs(3891));
    layer1_outputs(1873) <= not((layer0_outputs(3065)) or (layer0_outputs(4109)));
    layer1_outputs(1874) <= not(layer0_outputs(2546));
    layer1_outputs(1875) <= (layer0_outputs(4828)) or (layer0_outputs(753));
    layer1_outputs(1876) <= not((layer0_outputs(5006)) or (layer0_outputs(2698)));
    layer1_outputs(1877) <= not(layer0_outputs(2454));
    layer1_outputs(1878) <= not((layer0_outputs(2454)) or (layer0_outputs(3679)));
    layer1_outputs(1879) <= '1';
    layer1_outputs(1880) <= '1';
    layer1_outputs(1881) <= '1';
    layer1_outputs(1882) <= layer0_outputs(161);
    layer1_outputs(1883) <= (layer0_outputs(2603)) and not (layer0_outputs(4249));
    layer1_outputs(1884) <= not((layer0_outputs(4871)) and (layer0_outputs(3885)));
    layer1_outputs(1885) <= not(layer0_outputs(2498));
    layer1_outputs(1886) <= layer0_outputs(3579);
    layer1_outputs(1887) <= (layer0_outputs(3114)) or (layer0_outputs(2652));
    layer1_outputs(1888) <= '1';
    layer1_outputs(1889) <= not((layer0_outputs(4707)) or (layer0_outputs(4454)));
    layer1_outputs(1890) <= not((layer0_outputs(934)) and (layer0_outputs(1768)));
    layer1_outputs(1891) <= '0';
    layer1_outputs(1892) <= (layer0_outputs(2551)) and not (layer0_outputs(2641));
    layer1_outputs(1893) <= '1';
    layer1_outputs(1894) <= (layer0_outputs(2806)) and not (layer0_outputs(999));
    layer1_outputs(1895) <= not(layer0_outputs(2)) or (layer0_outputs(1134));
    layer1_outputs(1896) <= '0';
    layer1_outputs(1897) <= not((layer0_outputs(417)) or (layer0_outputs(2580)));
    layer1_outputs(1898) <= '0';
    layer1_outputs(1899) <= not(layer0_outputs(3681)) or (layer0_outputs(834));
    layer1_outputs(1900) <= (layer0_outputs(2007)) and not (layer0_outputs(2210));
    layer1_outputs(1901) <= layer0_outputs(4325);
    layer1_outputs(1902) <= not((layer0_outputs(4121)) and (layer0_outputs(1307)));
    layer1_outputs(1903) <= not((layer0_outputs(2391)) or (layer0_outputs(4155)));
    layer1_outputs(1904) <= '1';
    layer1_outputs(1905) <= '1';
    layer1_outputs(1906) <= not(layer0_outputs(281)) or (layer0_outputs(721));
    layer1_outputs(1907) <= (layer0_outputs(4351)) and not (layer0_outputs(36));
    layer1_outputs(1908) <= (layer0_outputs(16)) and not (layer0_outputs(720));
    layer1_outputs(1909) <= layer0_outputs(204);
    layer1_outputs(1910) <= not(layer0_outputs(2272));
    layer1_outputs(1911) <= not((layer0_outputs(786)) and (layer0_outputs(4037)));
    layer1_outputs(1912) <= (layer0_outputs(4036)) and not (layer0_outputs(4059));
    layer1_outputs(1913) <= not(layer0_outputs(202)) or (layer0_outputs(670));
    layer1_outputs(1914) <= (layer0_outputs(282)) or (layer0_outputs(1654));
    layer1_outputs(1915) <= '0';
    layer1_outputs(1916) <= not(layer0_outputs(3013)) or (layer0_outputs(3412));
    layer1_outputs(1917) <= (layer0_outputs(1232)) and not (layer0_outputs(1651));
    layer1_outputs(1918) <= not((layer0_outputs(2509)) and (layer0_outputs(221)));
    layer1_outputs(1919) <= '0';
    layer1_outputs(1920) <= layer0_outputs(919);
    layer1_outputs(1921) <= layer0_outputs(2136);
    layer1_outputs(1922) <= not((layer0_outputs(4478)) and (layer0_outputs(2437)));
    layer1_outputs(1923) <= '0';
    layer1_outputs(1924) <= not((layer0_outputs(4994)) or (layer0_outputs(4486)));
    layer1_outputs(1925) <= not(layer0_outputs(3872));
    layer1_outputs(1926) <= '0';
    layer1_outputs(1927) <= not((layer0_outputs(4865)) or (layer0_outputs(1190)));
    layer1_outputs(1928) <= not((layer0_outputs(827)) or (layer0_outputs(5107)));
    layer1_outputs(1929) <= not(layer0_outputs(1532)) or (layer0_outputs(1485));
    layer1_outputs(1930) <= '0';
    layer1_outputs(1931) <= not(layer0_outputs(3384));
    layer1_outputs(1932) <= not(layer0_outputs(1187));
    layer1_outputs(1933) <= '1';
    layer1_outputs(1934) <= '0';
    layer1_outputs(1935) <= (layer0_outputs(1906)) and (layer0_outputs(1401));
    layer1_outputs(1936) <= '1';
    layer1_outputs(1937) <= (layer0_outputs(3008)) and not (layer0_outputs(1467));
    layer1_outputs(1938) <= not((layer0_outputs(3537)) or (layer0_outputs(3434)));
    layer1_outputs(1939) <= (layer0_outputs(4388)) xor (layer0_outputs(3482));
    layer1_outputs(1940) <= layer0_outputs(4424);
    layer1_outputs(1941) <= '0';
    layer1_outputs(1942) <= '1';
    layer1_outputs(1943) <= '1';
    layer1_outputs(1944) <= layer0_outputs(3701);
    layer1_outputs(1945) <= (layer0_outputs(2582)) and not (layer0_outputs(4840));
    layer1_outputs(1946) <= not(layer0_outputs(3781)) or (layer0_outputs(2440));
    layer1_outputs(1947) <= not(layer0_outputs(3973));
    layer1_outputs(1948) <= not(layer0_outputs(1663)) or (layer0_outputs(2813));
    layer1_outputs(1949) <= not(layer0_outputs(4154)) or (layer0_outputs(1268));
    layer1_outputs(1950) <= not((layer0_outputs(1320)) or (layer0_outputs(2279)));
    layer1_outputs(1951) <= (layer0_outputs(4417)) and not (layer0_outputs(1890));
    layer1_outputs(1952) <= layer0_outputs(2800);
    layer1_outputs(1953) <= layer0_outputs(3031);
    layer1_outputs(1954) <= not(layer0_outputs(1168)) or (layer0_outputs(3343));
    layer1_outputs(1955) <= '0';
    layer1_outputs(1956) <= not((layer0_outputs(3642)) or (layer0_outputs(1934)));
    layer1_outputs(1957) <= '0';
    layer1_outputs(1958) <= layer0_outputs(3586);
    layer1_outputs(1959) <= '0';
    layer1_outputs(1960) <= layer0_outputs(1740);
    layer1_outputs(1961) <= (layer0_outputs(744)) and (layer0_outputs(1239));
    layer1_outputs(1962) <= (layer0_outputs(4834)) and not (layer0_outputs(1720));
    layer1_outputs(1963) <= layer0_outputs(1124);
    layer1_outputs(1964) <= (layer0_outputs(4402)) and not (layer0_outputs(401));
    layer1_outputs(1965) <= (layer0_outputs(3138)) and (layer0_outputs(1050));
    layer1_outputs(1966) <= not(layer0_outputs(3392)) or (layer0_outputs(522));
    layer1_outputs(1967) <= (layer0_outputs(4703)) or (layer0_outputs(1930));
    layer1_outputs(1968) <= not((layer0_outputs(3256)) and (layer0_outputs(3996)));
    layer1_outputs(1969) <= layer0_outputs(29);
    layer1_outputs(1970) <= '0';
    layer1_outputs(1971) <= layer0_outputs(1588);
    layer1_outputs(1972) <= '1';
    layer1_outputs(1973) <= not(layer0_outputs(3805));
    layer1_outputs(1974) <= (layer0_outputs(206)) and not (layer0_outputs(2744));
    layer1_outputs(1975) <= not((layer0_outputs(2277)) and (layer0_outputs(3711)));
    layer1_outputs(1976) <= layer0_outputs(1514);
    layer1_outputs(1977) <= layer0_outputs(2876);
    layer1_outputs(1978) <= '0';
    layer1_outputs(1979) <= '0';
    layer1_outputs(1980) <= layer0_outputs(40);
    layer1_outputs(1981) <= (layer0_outputs(1668)) or (layer0_outputs(265));
    layer1_outputs(1982) <= '0';
    layer1_outputs(1983) <= (layer0_outputs(531)) and not (layer0_outputs(606));
    layer1_outputs(1984) <= '0';
    layer1_outputs(1985) <= (layer0_outputs(1410)) xor (layer0_outputs(1950));
    layer1_outputs(1986) <= (layer0_outputs(211)) or (layer0_outputs(2400));
    layer1_outputs(1987) <= (layer0_outputs(3546)) or (layer0_outputs(3401));
    layer1_outputs(1988) <= (layer0_outputs(4438)) or (layer0_outputs(953));
    layer1_outputs(1989) <= '1';
    layer1_outputs(1990) <= not(layer0_outputs(4236)) or (layer0_outputs(1110));
    layer1_outputs(1991) <= (layer0_outputs(887)) and not (layer0_outputs(4858));
    layer1_outputs(1992) <= not(layer0_outputs(58)) or (layer0_outputs(4250));
    layer1_outputs(1993) <= not(layer0_outputs(482)) or (layer0_outputs(4428));
    layer1_outputs(1994) <= not((layer0_outputs(432)) and (layer0_outputs(2400)));
    layer1_outputs(1995) <= layer0_outputs(3346);
    layer1_outputs(1996) <= not(layer0_outputs(4306)) or (layer0_outputs(550));
    layer1_outputs(1997) <= layer0_outputs(3596);
    layer1_outputs(1998) <= '1';
    layer1_outputs(1999) <= '1';
    layer1_outputs(2000) <= layer0_outputs(825);
    layer1_outputs(2001) <= not(layer0_outputs(3860)) or (layer0_outputs(2712));
    layer1_outputs(2002) <= (layer0_outputs(2264)) xor (layer0_outputs(985));
    layer1_outputs(2003) <= '0';
    layer1_outputs(2004) <= (layer0_outputs(4216)) and (layer0_outputs(4394));
    layer1_outputs(2005) <= layer0_outputs(917);
    layer1_outputs(2006) <= not(layer0_outputs(2823)) or (layer0_outputs(119));
    layer1_outputs(2007) <= not((layer0_outputs(1557)) and (layer0_outputs(5012)));
    layer1_outputs(2008) <= (layer0_outputs(3174)) and (layer0_outputs(2115));
    layer1_outputs(2009) <= not((layer0_outputs(1128)) and (layer0_outputs(1735)));
    layer1_outputs(2010) <= not((layer0_outputs(4931)) and (layer0_outputs(5026)));
    layer1_outputs(2011) <= not(layer0_outputs(742)) or (layer0_outputs(2154));
    layer1_outputs(2012) <= '0';
    layer1_outputs(2013) <= '0';
    layer1_outputs(2014) <= not((layer0_outputs(2443)) and (layer0_outputs(4440)));
    layer1_outputs(2015) <= '0';
    layer1_outputs(2016) <= (layer0_outputs(2929)) and not (layer0_outputs(5066));
    layer1_outputs(2017) <= (layer0_outputs(2795)) and not (layer0_outputs(2555));
    layer1_outputs(2018) <= (layer0_outputs(4127)) or (layer0_outputs(2336));
    layer1_outputs(2019) <= '0';
    layer1_outputs(2020) <= '0';
    layer1_outputs(2021) <= (layer0_outputs(4715)) and not (layer0_outputs(1412));
    layer1_outputs(2022) <= not(layer0_outputs(3410));
    layer1_outputs(2023) <= '0';
    layer1_outputs(2024) <= '1';
    layer1_outputs(2025) <= (layer0_outputs(4548)) and (layer0_outputs(2456));
    layer1_outputs(2026) <= (layer0_outputs(1265)) and (layer0_outputs(3696));
    layer1_outputs(2027) <= not(layer0_outputs(515));
    layer1_outputs(2028) <= not(layer0_outputs(2325)) or (layer0_outputs(1102));
    layer1_outputs(2029) <= '0';
    layer1_outputs(2030) <= '0';
    layer1_outputs(2031) <= (layer0_outputs(4173)) and not (layer0_outputs(295));
    layer1_outputs(2032) <= '0';
    layer1_outputs(2033) <= (layer0_outputs(4688)) and not (layer0_outputs(1023));
    layer1_outputs(2034) <= not((layer0_outputs(1863)) and (layer0_outputs(2831)));
    layer1_outputs(2035) <= layer0_outputs(4040);
    layer1_outputs(2036) <= not(layer0_outputs(2883)) or (layer0_outputs(5108));
    layer1_outputs(2037) <= not(layer0_outputs(854));
    layer1_outputs(2038) <= '0';
    layer1_outputs(2039) <= not(layer0_outputs(1770));
    layer1_outputs(2040) <= not(layer0_outputs(1932));
    layer1_outputs(2041) <= not((layer0_outputs(3988)) or (layer0_outputs(4411)));
    layer1_outputs(2042) <= not((layer0_outputs(2521)) and (layer0_outputs(1085)));
    layer1_outputs(2043) <= (layer0_outputs(2520)) and (layer0_outputs(4067));
    layer1_outputs(2044) <= not(layer0_outputs(4525));
    layer1_outputs(2045) <= '1';
    layer1_outputs(2046) <= '0';
    layer1_outputs(2047) <= '0';
    layer1_outputs(2048) <= '1';
    layer1_outputs(2049) <= not((layer0_outputs(1954)) or (layer0_outputs(319)));
    layer1_outputs(2050) <= not(layer0_outputs(1536));
    layer1_outputs(2051) <= (layer0_outputs(2898)) xor (layer0_outputs(1418));
    layer1_outputs(2052) <= '0';
    layer1_outputs(2053) <= layer0_outputs(4008);
    layer1_outputs(2054) <= not(layer0_outputs(3936)) or (layer0_outputs(1702));
    layer1_outputs(2055) <= not(layer0_outputs(3140));
    layer1_outputs(2056) <= not(layer0_outputs(2353)) or (layer0_outputs(2331));
    layer1_outputs(2057) <= not(layer0_outputs(88));
    layer1_outputs(2058) <= layer0_outputs(3014);
    layer1_outputs(2059) <= (layer0_outputs(1713)) and not (layer0_outputs(1248));
    layer1_outputs(2060) <= not(layer0_outputs(4732));
    layer1_outputs(2061) <= not((layer0_outputs(646)) and (layer0_outputs(2702)));
    layer1_outputs(2062) <= not(layer0_outputs(4046)) or (layer0_outputs(2011));
    layer1_outputs(2063) <= '0';
    layer1_outputs(2064) <= not(layer0_outputs(255)) or (layer0_outputs(4987));
    layer1_outputs(2065) <= not(layer0_outputs(2777));
    layer1_outputs(2066) <= (layer0_outputs(3016)) and not (layer0_outputs(1388));
    layer1_outputs(2067) <= not((layer0_outputs(2042)) or (layer0_outputs(1850)));
    layer1_outputs(2068) <= layer0_outputs(755);
    layer1_outputs(2069) <= (layer0_outputs(3624)) and (layer0_outputs(1322));
    layer1_outputs(2070) <= (layer0_outputs(4541)) or (layer0_outputs(448));
    layer1_outputs(2071) <= '0';
    layer1_outputs(2072) <= not((layer0_outputs(2571)) and (layer0_outputs(4058)));
    layer1_outputs(2073) <= not(layer0_outputs(3383)) or (layer0_outputs(707));
    layer1_outputs(2074) <= (layer0_outputs(4845)) and not (layer0_outputs(3893));
    layer1_outputs(2075) <= not(layer0_outputs(4935)) or (layer0_outputs(767));
    layer1_outputs(2076) <= '0';
    layer1_outputs(2077) <= not(layer0_outputs(1163)) or (layer0_outputs(3370));
    layer1_outputs(2078) <= '1';
    layer1_outputs(2079) <= (layer0_outputs(3490)) and not (layer0_outputs(3139));
    layer1_outputs(2080) <= layer0_outputs(1049);
    layer1_outputs(2081) <= '0';
    layer1_outputs(2082) <= not(layer0_outputs(2599));
    layer1_outputs(2083) <= layer0_outputs(984);
    layer1_outputs(2084) <= not((layer0_outputs(4188)) xor (layer0_outputs(2118)));
    layer1_outputs(2085) <= not(layer0_outputs(4386));
    layer1_outputs(2086) <= not((layer0_outputs(3425)) and (layer0_outputs(386)));
    layer1_outputs(2087) <= not((layer0_outputs(4948)) or (layer0_outputs(5023)));
    layer1_outputs(2088) <= '1';
    layer1_outputs(2089) <= '0';
    layer1_outputs(2090) <= layer0_outputs(5074);
    layer1_outputs(2091) <= '0';
    layer1_outputs(2092) <= layer0_outputs(1682);
    layer1_outputs(2093) <= (layer0_outputs(423)) and not (layer0_outputs(5065));
    layer1_outputs(2094) <= '0';
    layer1_outputs(2095) <= (layer0_outputs(3247)) and not (layer0_outputs(123));
    layer1_outputs(2096) <= (layer0_outputs(3760)) or (layer0_outputs(522));
    layer1_outputs(2097) <= '1';
    layer1_outputs(2098) <= not(layer0_outputs(2416)) or (layer0_outputs(3173));
    layer1_outputs(2099) <= (layer0_outputs(3120)) and not (layer0_outputs(2390));
    layer1_outputs(2100) <= not(layer0_outputs(2308)) or (layer0_outputs(2726));
    layer1_outputs(2101) <= (layer0_outputs(1922)) and (layer0_outputs(3444));
    layer1_outputs(2102) <= not((layer0_outputs(1851)) and (layer0_outputs(4668)));
    layer1_outputs(2103) <= not(layer0_outputs(4938)) or (layer0_outputs(1202));
    layer1_outputs(2104) <= (layer0_outputs(1630)) or (layer0_outputs(4599));
    layer1_outputs(2105) <= not(layer0_outputs(2525)) or (layer0_outputs(3635));
    layer1_outputs(2106) <= layer0_outputs(2767);
    layer1_outputs(2107) <= not(layer0_outputs(4920)) or (layer0_outputs(3728));
    layer1_outputs(2108) <= '0';
    layer1_outputs(2109) <= (layer0_outputs(3873)) xor (layer0_outputs(106));
    layer1_outputs(2110) <= not(layer0_outputs(3973));
    layer1_outputs(2111) <= not(layer0_outputs(3199)) or (layer0_outputs(4119));
    layer1_outputs(2112) <= (layer0_outputs(2648)) and (layer0_outputs(1759));
    layer1_outputs(2113) <= not(layer0_outputs(1580));
    layer1_outputs(2114) <= not((layer0_outputs(4865)) and (layer0_outputs(3835)));
    layer1_outputs(2115) <= not(layer0_outputs(468)) or (layer0_outputs(2418));
    layer1_outputs(2116) <= layer0_outputs(4577);
    layer1_outputs(2117) <= '0';
    layer1_outputs(2118) <= not((layer0_outputs(625)) and (layer0_outputs(4244)));
    layer1_outputs(2119) <= '0';
    layer1_outputs(2120) <= (layer0_outputs(103)) and (layer0_outputs(3552));
    layer1_outputs(2121) <= '0';
    layer1_outputs(2122) <= not(layer0_outputs(3668)) or (layer0_outputs(3074));
    layer1_outputs(2123) <= not(layer0_outputs(540)) or (layer0_outputs(257));
    layer1_outputs(2124) <= layer0_outputs(3451);
    layer1_outputs(2125) <= not((layer0_outputs(4643)) and (layer0_outputs(992)));
    layer1_outputs(2126) <= layer0_outputs(404);
    layer1_outputs(2127) <= (layer0_outputs(1050)) and not (layer0_outputs(4691));
    layer1_outputs(2128) <= (layer0_outputs(1999)) and not (layer0_outputs(2598));
    layer1_outputs(2129) <= not(layer0_outputs(3198)) or (layer0_outputs(3879));
    layer1_outputs(2130) <= not(layer0_outputs(4890));
    layer1_outputs(2131) <= (layer0_outputs(2853)) and not (layer0_outputs(111));
    layer1_outputs(2132) <= '0';
    layer1_outputs(2133) <= (layer0_outputs(1689)) and not (layer0_outputs(798));
    layer1_outputs(2134) <= not(layer0_outputs(878));
    layer1_outputs(2135) <= not(layer0_outputs(2567));
    layer1_outputs(2136) <= not(layer0_outputs(1033));
    layer1_outputs(2137) <= '0';
    layer1_outputs(2138) <= (layer0_outputs(3261)) or (layer0_outputs(4329));
    layer1_outputs(2139) <= layer0_outputs(3460);
    layer1_outputs(2140) <= not((layer0_outputs(1047)) or (layer0_outputs(2119)));
    layer1_outputs(2141) <= not((layer0_outputs(3439)) and (layer0_outputs(3502)));
    layer1_outputs(2142) <= '0';
    layer1_outputs(2143) <= layer0_outputs(2489);
    layer1_outputs(2144) <= not(layer0_outputs(4939)) or (layer0_outputs(3147));
    layer1_outputs(2145) <= layer0_outputs(363);
    layer1_outputs(2146) <= (layer0_outputs(5105)) and (layer0_outputs(2318));
    layer1_outputs(2147) <= '1';
    layer1_outputs(2148) <= not((layer0_outputs(803)) and (layer0_outputs(5016)));
    layer1_outputs(2149) <= layer0_outputs(4213);
    layer1_outputs(2150) <= '0';
    layer1_outputs(2151) <= (layer0_outputs(330)) and (layer0_outputs(1843));
    layer1_outputs(2152) <= not((layer0_outputs(2886)) or (layer0_outputs(4437)));
    layer1_outputs(2153) <= '0';
    layer1_outputs(2154) <= '0';
    layer1_outputs(2155) <= (layer0_outputs(654)) and not (layer0_outputs(3418));
    layer1_outputs(2156) <= (layer0_outputs(4176)) and (layer0_outputs(4078));
    layer1_outputs(2157) <= not((layer0_outputs(5043)) xor (layer0_outputs(4259)));
    layer1_outputs(2158) <= (layer0_outputs(1729)) or (layer0_outputs(479));
    layer1_outputs(2159) <= not((layer0_outputs(1972)) and (layer0_outputs(1327)));
    layer1_outputs(2160) <= (layer0_outputs(3363)) and (layer0_outputs(3229));
    layer1_outputs(2161) <= not((layer0_outputs(2743)) and (layer0_outputs(1709)));
    layer1_outputs(2162) <= layer0_outputs(7);
    layer1_outputs(2163) <= '0';
    layer1_outputs(2164) <= (layer0_outputs(3029)) and (layer0_outputs(3202));
    layer1_outputs(2165) <= not(layer0_outputs(3480)) or (layer0_outputs(21));
    layer1_outputs(2166) <= '0';
    layer1_outputs(2167) <= '0';
    layer1_outputs(2168) <= not(layer0_outputs(270));
    layer1_outputs(2169) <= '0';
    layer1_outputs(2170) <= not(layer0_outputs(4093)) or (layer0_outputs(1599));
    layer1_outputs(2171) <= (layer0_outputs(2292)) and not (layer0_outputs(151));
    layer1_outputs(2172) <= not(layer0_outputs(1997));
    layer1_outputs(2173) <= '0';
    layer1_outputs(2174) <= layer0_outputs(105);
    layer1_outputs(2175) <= '0';
    layer1_outputs(2176) <= (layer0_outputs(2433)) xor (layer0_outputs(4785));
    layer1_outputs(2177) <= '0';
    layer1_outputs(2178) <= '1';
    layer1_outputs(2179) <= not(layer0_outputs(4147));
    layer1_outputs(2180) <= '1';
    layer1_outputs(2181) <= (layer0_outputs(63)) and not (layer0_outputs(893));
    layer1_outputs(2182) <= (layer0_outputs(1968)) and (layer0_outputs(651));
    layer1_outputs(2183) <= (layer0_outputs(4819)) and (layer0_outputs(3339));
    layer1_outputs(2184) <= '0';
    layer1_outputs(2185) <= '1';
    layer1_outputs(2186) <= (layer0_outputs(469)) and not (layer0_outputs(2466));
    layer1_outputs(2187) <= layer0_outputs(3184);
    layer1_outputs(2188) <= (layer0_outputs(4728)) and (layer0_outputs(911));
    layer1_outputs(2189) <= '1';
    layer1_outputs(2190) <= layer0_outputs(4584);
    layer1_outputs(2191) <= '0';
    layer1_outputs(2192) <= layer0_outputs(861);
    layer1_outputs(2193) <= not((layer0_outputs(4590)) and (layer0_outputs(4384)));
    layer1_outputs(2194) <= (layer0_outputs(1263)) and (layer0_outputs(1362));
    layer1_outputs(2195) <= (layer0_outputs(4778)) and (layer0_outputs(1637));
    layer1_outputs(2196) <= not((layer0_outputs(362)) and (layer0_outputs(1340)));
    layer1_outputs(2197) <= not(layer0_outputs(3803));
    layer1_outputs(2198) <= '0';
    layer1_outputs(2199) <= '0';
    layer1_outputs(2200) <= not((layer0_outputs(4941)) and (layer0_outputs(1189)));
    layer1_outputs(2201) <= not(layer0_outputs(2151)) or (layer0_outputs(3160));
    layer1_outputs(2202) <= not(layer0_outputs(1038));
    layer1_outputs(2203) <= (layer0_outputs(3799)) and (layer0_outputs(3263));
    layer1_outputs(2204) <= (layer0_outputs(4614)) and (layer0_outputs(1999));
    layer1_outputs(2205) <= layer0_outputs(3831);
    layer1_outputs(2206) <= '0';
    layer1_outputs(2207) <= not((layer0_outputs(3287)) and (layer0_outputs(3345)));
    layer1_outputs(2208) <= '0';
    layer1_outputs(2209) <= '0';
    layer1_outputs(2210) <= not(layer0_outputs(95));
    layer1_outputs(2211) <= layer0_outputs(3566);
    layer1_outputs(2212) <= not(layer0_outputs(2501)) or (layer0_outputs(3926));
    layer1_outputs(2213) <= not((layer0_outputs(4286)) and (layer0_outputs(4602)));
    layer1_outputs(2214) <= '1';
    layer1_outputs(2215) <= '0';
    layer1_outputs(2216) <= '1';
    layer1_outputs(2217) <= '1';
    layer1_outputs(2218) <= layer0_outputs(3501);
    layer1_outputs(2219) <= not(layer0_outputs(2774));
    layer1_outputs(2220) <= (layer0_outputs(1302)) and not (layer0_outputs(4393));
    layer1_outputs(2221) <= not((layer0_outputs(4618)) and (layer0_outputs(1347)));
    layer1_outputs(2222) <= not((layer0_outputs(4345)) or (layer0_outputs(2047)));
    layer1_outputs(2223) <= not((layer0_outputs(201)) and (layer0_outputs(1114)));
    layer1_outputs(2224) <= (layer0_outputs(3793)) and (layer0_outputs(664));
    layer1_outputs(2225) <= not(layer0_outputs(4336)) or (layer0_outputs(3450));
    layer1_outputs(2226) <= not((layer0_outputs(2380)) xor (layer0_outputs(3108)));
    layer1_outputs(2227) <= '1';
    layer1_outputs(2228) <= (layer0_outputs(4583)) and (layer0_outputs(663));
    layer1_outputs(2229) <= (layer0_outputs(1519)) or (layer0_outputs(193));
    layer1_outputs(2230) <= (layer0_outputs(1374)) or (layer0_outputs(4236));
    layer1_outputs(2231) <= not(layer0_outputs(2715));
    layer1_outputs(2232) <= not((layer0_outputs(2836)) and (layer0_outputs(2123)));
    layer1_outputs(2233) <= layer0_outputs(764);
    layer1_outputs(2234) <= not((layer0_outputs(1801)) or (layer0_outputs(4801)));
    layer1_outputs(2235) <= (layer0_outputs(2399)) and not (layer0_outputs(3672));
    layer1_outputs(2236) <= not((layer0_outputs(1293)) and (layer0_outputs(229)));
    layer1_outputs(2237) <= not((layer0_outputs(3531)) or (layer0_outputs(1453)));
    layer1_outputs(2238) <= '1';
    layer1_outputs(2239) <= not((layer0_outputs(837)) or (layer0_outputs(4265)));
    layer1_outputs(2240) <= not((layer0_outputs(2473)) or (layer0_outputs(4011)));
    layer1_outputs(2241) <= not(layer0_outputs(3206)) or (layer0_outputs(3638));
    layer1_outputs(2242) <= not(layer0_outputs(3963));
    layer1_outputs(2243) <= (layer0_outputs(1825)) and not (layer0_outputs(1985));
    layer1_outputs(2244) <= '1';
    layer1_outputs(2245) <= not((layer0_outputs(5025)) or (layer0_outputs(4450)));
    layer1_outputs(2246) <= (layer0_outputs(1770)) and (layer0_outputs(1021));
    layer1_outputs(2247) <= '1';
    layer1_outputs(2248) <= '0';
    layer1_outputs(2249) <= (layer0_outputs(2035)) or (layer0_outputs(654));
    layer1_outputs(2250) <= '0';
    layer1_outputs(2251) <= not((layer0_outputs(3247)) and (layer0_outputs(970)));
    layer1_outputs(2252) <= '1';
    layer1_outputs(2253) <= '1';
    layer1_outputs(2254) <= '1';
    layer1_outputs(2255) <= layer0_outputs(2649);
    layer1_outputs(2256) <= not((layer0_outputs(4156)) or (layer0_outputs(3849)));
    layer1_outputs(2257) <= layer0_outputs(1515);
    layer1_outputs(2258) <= (layer0_outputs(4475)) or (layer0_outputs(1353));
    layer1_outputs(2259) <= not(layer0_outputs(3026));
    layer1_outputs(2260) <= not(layer0_outputs(4688)) or (layer0_outputs(2178));
    layer1_outputs(2261) <= (layer0_outputs(3898)) and (layer0_outputs(1104));
    layer1_outputs(2262) <= '1';
    layer1_outputs(2263) <= '0';
    layer1_outputs(2264) <= (layer0_outputs(1948)) or (layer0_outputs(122));
    layer1_outputs(2265) <= not(layer0_outputs(3721)) or (layer0_outputs(5000));
    layer1_outputs(2266) <= '1';
    layer1_outputs(2267) <= not(layer0_outputs(4364));
    layer1_outputs(2268) <= '0';
    layer1_outputs(2269) <= '1';
    layer1_outputs(2270) <= not((layer0_outputs(3565)) or (layer0_outputs(3217)));
    layer1_outputs(2271) <= not((layer0_outputs(4781)) and (layer0_outputs(2024)));
    layer1_outputs(2272) <= not(layer0_outputs(539));
    layer1_outputs(2273) <= not(layer0_outputs(3603));
    layer1_outputs(2274) <= layer0_outputs(4074);
    layer1_outputs(2275) <= (layer0_outputs(3071)) and not (layer0_outputs(496));
    layer1_outputs(2276) <= layer0_outputs(78);
    layer1_outputs(2277) <= (layer0_outputs(929)) and not (layer0_outputs(4038));
    layer1_outputs(2278) <= (layer0_outputs(2906)) and not (layer0_outputs(2787));
    layer1_outputs(2279) <= '0';
    layer1_outputs(2280) <= not((layer0_outputs(2959)) and (layer0_outputs(2430)));
    layer1_outputs(2281) <= not(layer0_outputs(3820)) or (layer0_outputs(2280));
    layer1_outputs(2282) <= not((layer0_outputs(4825)) and (layer0_outputs(222)));
    layer1_outputs(2283) <= (layer0_outputs(4765)) or (layer0_outputs(3457));
    layer1_outputs(2284) <= layer0_outputs(692);
    layer1_outputs(2285) <= '1';
    layer1_outputs(2286) <= (layer0_outputs(347)) and not (layer0_outputs(4197));
    layer1_outputs(2287) <= layer0_outputs(2517);
    layer1_outputs(2288) <= not((layer0_outputs(3437)) and (layer0_outputs(2601)));
    layer1_outputs(2289) <= '1';
    layer1_outputs(2290) <= layer0_outputs(4630);
    layer1_outputs(2291) <= (layer0_outputs(1152)) and (layer0_outputs(2142));
    layer1_outputs(2292) <= layer0_outputs(4015);
    layer1_outputs(2293) <= '0';
    layer1_outputs(2294) <= '1';
    layer1_outputs(2295) <= '0';
    layer1_outputs(2296) <= (layer0_outputs(3420)) and not (layer0_outputs(400));
    layer1_outputs(2297) <= not(layer0_outputs(2381)) or (layer0_outputs(464));
    layer1_outputs(2298) <= not(layer0_outputs(4608));
    layer1_outputs(2299) <= (layer0_outputs(4815)) or (layer0_outputs(2139));
    layer1_outputs(2300) <= '1';
    layer1_outputs(2301) <= (layer0_outputs(3183)) and (layer0_outputs(4898));
    layer1_outputs(2302) <= (layer0_outputs(555)) and not (layer0_outputs(4949));
    layer1_outputs(2303) <= '1';
    layer1_outputs(2304) <= '0';
    layer1_outputs(2305) <= not(layer0_outputs(575)) or (layer0_outputs(1053));
    layer1_outputs(2306) <= not((layer0_outputs(3705)) and (layer0_outputs(1629)));
    layer1_outputs(2307) <= not(layer0_outputs(2752)) or (layer0_outputs(1697));
    layer1_outputs(2308) <= layer0_outputs(4547);
    layer1_outputs(2309) <= '0';
    layer1_outputs(2310) <= layer0_outputs(3888);
    layer1_outputs(2311) <= (layer0_outputs(4791)) and not (layer0_outputs(3762));
    layer1_outputs(2312) <= not(layer0_outputs(1397));
    layer1_outputs(2313) <= not((layer0_outputs(407)) and (layer0_outputs(605)));
    layer1_outputs(2314) <= not(layer0_outputs(2875));
    layer1_outputs(2315) <= not(layer0_outputs(4933));
    layer1_outputs(2316) <= not(layer0_outputs(923)) or (layer0_outputs(2489));
    layer1_outputs(2317) <= '0';
    layer1_outputs(2318) <= not((layer0_outputs(4997)) or (layer0_outputs(431)));
    layer1_outputs(2319) <= layer0_outputs(1414);
    layer1_outputs(2320) <= '1';
    layer1_outputs(2321) <= not(layer0_outputs(2441)) or (layer0_outputs(2312));
    layer1_outputs(2322) <= '0';
    layer1_outputs(2323) <= (layer0_outputs(3593)) and not (layer0_outputs(183));
    layer1_outputs(2324) <= (layer0_outputs(1248)) or (layer0_outputs(3529));
    layer1_outputs(2325) <= '0';
    layer1_outputs(2326) <= (layer0_outputs(1583)) or (layer0_outputs(4455));
    layer1_outputs(2327) <= not(layer0_outputs(4497)) or (layer0_outputs(4793));
    layer1_outputs(2328) <= '0';
    layer1_outputs(2329) <= '0';
    layer1_outputs(2330) <= '1';
    layer1_outputs(2331) <= layer0_outputs(2065);
    layer1_outputs(2332) <= layer0_outputs(2719);
    layer1_outputs(2333) <= not(layer0_outputs(1565)) or (layer0_outputs(2133));
    layer1_outputs(2334) <= not(layer0_outputs(5044));
    layer1_outputs(2335) <= layer0_outputs(632);
    layer1_outputs(2336) <= not((layer0_outputs(3049)) or (layer0_outputs(4362)));
    layer1_outputs(2337) <= not(layer0_outputs(3585)) or (layer0_outputs(1379));
    layer1_outputs(2338) <= (layer0_outputs(1713)) and (layer0_outputs(918));
    layer1_outputs(2339) <= '1';
    layer1_outputs(2340) <= (layer0_outputs(939)) and (layer0_outputs(1120));
    layer1_outputs(2341) <= layer0_outputs(612);
    layer1_outputs(2342) <= '1';
    layer1_outputs(2343) <= '1';
    layer1_outputs(2344) <= layer0_outputs(959);
    layer1_outputs(2345) <= layer0_outputs(3865);
    layer1_outputs(2346) <= '1';
    layer1_outputs(2347) <= (layer0_outputs(97)) and not (layer0_outputs(798));
    layer1_outputs(2348) <= (layer0_outputs(3965)) and not (layer0_outputs(3267));
    layer1_outputs(2349) <= '0';
    layer1_outputs(2350) <= not(layer0_outputs(4243));
    layer1_outputs(2351) <= (layer0_outputs(782)) and not (layer0_outputs(663));
    layer1_outputs(2352) <= not(layer0_outputs(471));
    layer1_outputs(2353) <= '1';
    layer1_outputs(2354) <= (layer0_outputs(438)) and not (layer0_outputs(1041));
    layer1_outputs(2355) <= not(layer0_outputs(3719));
    layer1_outputs(2356) <= not(layer0_outputs(714));
    layer1_outputs(2357) <= (layer0_outputs(2349)) and (layer0_outputs(38));
    layer1_outputs(2358) <= layer0_outputs(989);
    layer1_outputs(2359) <= (layer0_outputs(794)) and not (layer0_outputs(579));
    layer1_outputs(2360) <= (layer0_outputs(2890)) and not (layer0_outputs(2979));
    layer1_outputs(2361) <= (layer0_outputs(2745)) xor (layer0_outputs(168));
    layer1_outputs(2362) <= '0';
    layer1_outputs(2363) <= (layer0_outputs(3598)) and (layer0_outputs(2478));
    layer1_outputs(2364) <= not(layer0_outputs(221));
    layer1_outputs(2365) <= (layer0_outputs(3527)) and not (layer0_outputs(3293));
    layer1_outputs(2366) <= (layer0_outputs(4771)) or (layer0_outputs(4928));
    layer1_outputs(2367) <= '1';
    layer1_outputs(2368) <= (layer0_outputs(1902)) and (layer0_outputs(2305));
    layer1_outputs(2369) <= (layer0_outputs(3409)) and not (layer0_outputs(119));
    layer1_outputs(2370) <= (layer0_outputs(4126)) and not (layer0_outputs(224));
    layer1_outputs(2371) <= not(layer0_outputs(3155)) or (layer0_outputs(2876));
    layer1_outputs(2372) <= '0';
    layer1_outputs(2373) <= (layer0_outputs(3684)) and (layer0_outputs(1060));
    layer1_outputs(2374) <= not((layer0_outputs(2004)) or (layer0_outputs(4655)));
    layer1_outputs(2375) <= (layer0_outputs(4243)) and not (layer0_outputs(1321));
    layer1_outputs(2376) <= (layer0_outputs(3509)) or (layer0_outputs(3430));
    layer1_outputs(2377) <= (layer0_outputs(2516)) or (layer0_outputs(2759));
    layer1_outputs(2378) <= not(layer0_outputs(2737)) or (layer0_outputs(594));
    layer1_outputs(2379) <= (layer0_outputs(3827)) and (layer0_outputs(2250));
    layer1_outputs(2380) <= '1';
    layer1_outputs(2381) <= '1';
    layer1_outputs(2382) <= layer0_outputs(1864);
    layer1_outputs(2383) <= (layer0_outputs(1020)) or (layer0_outputs(4775));
    layer1_outputs(2384) <= not((layer0_outputs(1945)) or (layer0_outputs(4826)));
    layer1_outputs(2385) <= not(layer0_outputs(2267));
    layer1_outputs(2386) <= (layer0_outputs(71)) or (layer0_outputs(4496));
    layer1_outputs(2387) <= (layer0_outputs(1836)) and (layer0_outputs(1164));
    layer1_outputs(2388) <= '1';
    layer1_outputs(2389) <= not(layer0_outputs(2881));
    layer1_outputs(2390) <= (layer0_outputs(4653)) and (layer0_outputs(1216));
    layer1_outputs(2391) <= not(layer0_outputs(3886));
    layer1_outputs(2392) <= '1';
    layer1_outputs(2393) <= layer0_outputs(4810);
    layer1_outputs(2394) <= (layer0_outputs(3649)) xor (layer0_outputs(2151));
    layer1_outputs(2395) <= layer0_outputs(2986);
    layer1_outputs(2396) <= '0';
    layer1_outputs(2397) <= '1';
    layer1_outputs(2398) <= not(layer0_outputs(346));
    layer1_outputs(2399) <= (layer0_outputs(4420)) or (layer0_outputs(446));
    layer1_outputs(2400) <= (layer0_outputs(671)) or (layer0_outputs(952));
    layer1_outputs(2401) <= '0';
    layer1_outputs(2402) <= layer0_outputs(97);
    layer1_outputs(2403) <= (layer0_outputs(5094)) and not (layer0_outputs(3590));
    layer1_outputs(2404) <= not(layer0_outputs(2186));
    layer1_outputs(2405) <= '0';
    layer1_outputs(2406) <= not(layer0_outputs(527));
    layer1_outputs(2407) <= (layer0_outputs(2410)) and not (layer0_outputs(3360));
    layer1_outputs(2408) <= not(layer0_outputs(4584)) or (layer0_outputs(1896));
    layer1_outputs(2409) <= not((layer0_outputs(1794)) or (layer0_outputs(2904)));
    layer1_outputs(2410) <= not((layer0_outputs(4552)) or (layer0_outputs(2175)));
    layer1_outputs(2411) <= not((layer0_outputs(618)) or (layer0_outputs(4500)));
    layer1_outputs(2412) <= (layer0_outputs(3807)) and not (layer0_outputs(2846));
    layer1_outputs(2413) <= not(layer0_outputs(1645));
    layer1_outputs(2414) <= not(layer0_outputs(3432)) or (layer0_outputs(4637));
    layer1_outputs(2415) <= not((layer0_outputs(2817)) xor (layer0_outputs(73)));
    layer1_outputs(2416) <= (layer0_outputs(5060)) and not (layer0_outputs(2374));
    layer1_outputs(2417) <= (layer0_outputs(2064)) and not (layer0_outputs(610));
    layer1_outputs(2418) <= layer0_outputs(1097);
    layer1_outputs(2419) <= not((layer0_outputs(1313)) or (layer0_outputs(3766)));
    layer1_outputs(2420) <= not(layer0_outputs(1730)) or (layer0_outputs(3195));
    layer1_outputs(2421) <= not(layer0_outputs(4611));
    layer1_outputs(2422) <= not(layer0_outputs(1344));
    layer1_outputs(2423) <= not((layer0_outputs(4545)) and (layer0_outputs(493)));
    layer1_outputs(2424) <= layer0_outputs(4899);
    layer1_outputs(2425) <= (layer0_outputs(2104)) or (layer0_outputs(2615));
    layer1_outputs(2426) <= '1';
    layer1_outputs(2427) <= not((layer0_outputs(393)) or (layer0_outputs(3685)));
    layer1_outputs(2428) <= '1';
    layer1_outputs(2429) <= not((layer0_outputs(4903)) and (layer0_outputs(3464)));
    layer1_outputs(2430) <= (layer0_outputs(1823)) or (layer0_outputs(3895));
    layer1_outputs(2431) <= (layer0_outputs(3177)) or (layer0_outputs(425));
    layer1_outputs(2432) <= not((layer0_outputs(4005)) or (layer0_outputs(2920)));
    layer1_outputs(2433) <= '1';
    layer1_outputs(2434) <= '0';
    layer1_outputs(2435) <= layer0_outputs(1242);
    layer1_outputs(2436) <= not(layer0_outputs(512));
    layer1_outputs(2437) <= layer0_outputs(2567);
    layer1_outputs(2438) <= '0';
    layer1_outputs(2439) <= not(layer0_outputs(2094));
    layer1_outputs(2440) <= '0';
    layer1_outputs(2441) <= (layer0_outputs(3575)) or (layer0_outputs(4946));
    layer1_outputs(2442) <= (layer0_outputs(2735)) or (layer0_outputs(1884));
    layer1_outputs(2443) <= not(layer0_outputs(997)) or (layer0_outputs(2367));
    layer1_outputs(2444) <= '1';
    layer1_outputs(2445) <= not(layer0_outputs(1623));
    layer1_outputs(2446) <= (layer0_outputs(3150)) and not (layer0_outputs(2182));
    layer1_outputs(2447) <= layer0_outputs(1011);
    layer1_outputs(2448) <= not((layer0_outputs(3255)) and (layer0_outputs(3715)));
    layer1_outputs(2449) <= not(layer0_outputs(3044));
    layer1_outputs(2450) <= '1';
    layer1_outputs(2451) <= layer0_outputs(628);
    layer1_outputs(2452) <= '0';
    layer1_outputs(2453) <= (layer0_outputs(2408)) and not (layer0_outputs(2397));
    layer1_outputs(2454) <= '1';
    layer1_outputs(2455) <= layer0_outputs(1635);
    layer1_outputs(2456) <= '1';
    layer1_outputs(2457) <= (layer0_outputs(3702)) and (layer0_outputs(2540));
    layer1_outputs(2458) <= (layer0_outputs(4188)) and (layer0_outputs(3308));
    layer1_outputs(2459) <= not(layer0_outputs(1955));
    layer1_outputs(2460) <= (layer0_outputs(2138)) and (layer0_outputs(1608));
    layer1_outputs(2461) <= '1';
    layer1_outputs(2462) <= (layer0_outputs(4262)) or (layer0_outputs(1619));
    layer1_outputs(2463) <= not((layer0_outputs(4061)) or (layer0_outputs(2200)));
    layer1_outputs(2464) <= not(layer0_outputs(3261));
    layer1_outputs(2465) <= not(layer0_outputs(2026)) or (layer0_outputs(1855));
    layer1_outputs(2466) <= not(layer0_outputs(2984)) or (layer0_outputs(863));
    layer1_outputs(2467) <= (layer0_outputs(4655)) and (layer0_outputs(4638));
    layer1_outputs(2468) <= not(layer0_outputs(1129));
    layer1_outputs(2469) <= not((layer0_outputs(3192)) or (layer0_outputs(4045)));
    layer1_outputs(2470) <= (layer0_outputs(2226)) and (layer0_outputs(4492));
    layer1_outputs(2471) <= '0';
    layer1_outputs(2472) <= '0';
    layer1_outputs(2473) <= '1';
    layer1_outputs(2474) <= layer0_outputs(3459);
    layer1_outputs(2475) <= layer0_outputs(1246);
    layer1_outputs(2476) <= (layer0_outputs(2486)) and (layer0_outputs(4368));
    layer1_outputs(2477) <= '1';
    layer1_outputs(2478) <= not(layer0_outputs(3695));
    layer1_outputs(2479) <= '1';
    layer1_outputs(2480) <= '0';
    layer1_outputs(2481) <= not(layer0_outputs(1837)) or (layer0_outputs(4098));
    layer1_outputs(2482) <= not(layer0_outputs(2851)) or (layer0_outputs(2385));
    layer1_outputs(2483) <= not(layer0_outputs(45)) or (layer0_outputs(2819));
    layer1_outputs(2484) <= (layer0_outputs(3242)) and not (layer0_outputs(2087));
    layer1_outputs(2485) <= '0';
    layer1_outputs(2486) <= layer0_outputs(666);
    layer1_outputs(2487) <= not(layer0_outputs(2794)) or (layer0_outputs(4189));
    layer1_outputs(2488) <= (layer0_outputs(268)) and (layer0_outputs(4288));
    layer1_outputs(2489) <= layer0_outputs(4569);
    layer1_outputs(2490) <= not(layer0_outputs(4759));
    layer1_outputs(2491) <= (layer0_outputs(2794)) and (layer0_outputs(1881));
    layer1_outputs(2492) <= '1';
    layer1_outputs(2493) <= not((layer0_outputs(4585)) or (layer0_outputs(3594)));
    layer1_outputs(2494) <= '0';
    layer1_outputs(2495) <= not(layer0_outputs(1707)) or (layer0_outputs(631));
    layer1_outputs(2496) <= (layer0_outputs(2561)) and not (layer0_outputs(4185));
    layer1_outputs(2497) <= (layer0_outputs(5088)) or (layer0_outputs(1224));
    layer1_outputs(2498) <= (layer0_outputs(2798)) or (layer0_outputs(260));
    layer1_outputs(2499) <= not((layer0_outputs(4805)) xor (layer0_outputs(51)));
    layer1_outputs(2500) <= (layer0_outputs(1252)) and (layer0_outputs(1407));
    layer1_outputs(2501) <= (layer0_outputs(4484)) xor (layer0_outputs(336));
    layer1_outputs(2502) <= '1';
    layer1_outputs(2503) <= '0';
    layer1_outputs(2504) <= not(layer0_outputs(348)) or (layer0_outputs(2791));
    layer1_outputs(2505) <= not(layer0_outputs(3222)) or (layer0_outputs(1597));
    layer1_outputs(2506) <= '1';
    layer1_outputs(2507) <= (layer0_outputs(4284)) and not (layer0_outputs(831));
    layer1_outputs(2508) <= '0';
    layer1_outputs(2509) <= layer0_outputs(3098);
    layer1_outputs(2510) <= not(layer0_outputs(1746)) or (layer0_outputs(3022));
    layer1_outputs(2511) <= not(layer0_outputs(3360));
    layer1_outputs(2512) <= '0';
    layer1_outputs(2513) <= not((layer0_outputs(3870)) or (layer0_outputs(3605)));
    layer1_outputs(2514) <= (layer0_outputs(4183)) and not (layer0_outputs(4645));
    layer1_outputs(2515) <= not(layer0_outputs(1022));
    layer1_outputs(2516) <= layer0_outputs(4709);
    layer1_outputs(2517) <= not(layer0_outputs(2242)) or (layer0_outputs(4910));
    layer1_outputs(2518) <= (layer0_outputs(1469)) and not (layer0_outputs(3645));
    layer1_outputs(2519) <= '0';
    layer1_outputs(2520) <= not((layer0_outputs(2175)) and (layer0_outputs(4585)));
    layer1_outputs(2521) <= '0';
    layer1_outputs(2522) <= layer0_outputs(4660);
    layer1_outputs(2523) <= (layer0_outputs(1217)) and not (layer0_outputs(3009));
    layer1_outputs(2524) <= (layer0_outputs(2678)) xor (layer0_outputs(1433));
    layer1_outputs(2525) <= not(layer0_outputs(4574));
    layer1_outputs(2526) <= '0';
    layer1_outputs(2527) <= (layer0_outputs(2854)) and (layer0_outputs(3028));
    layer1_outputs(2528) <= (layer0_outputs(3627)) or (layer0_outputs(950));
    layer1_outputs(2529) <= '1';
    layer1_outputs(2530) <= not(layer0_outputs(238)) or (layer0_outputs(4257));
    layer1_outputs(2531) <= not(layer0_outputs(212)) or (layer0_outputs(2597));
    layer1_outputs(2532) <= layer0_outputs(638);
    layer1_outputs(2533) <= not(layer0_outputs(1331)) or (layer0_outputs(1130));
    layer1_outputs(2534) <= (layer0_outputs(566)) and not (layer0_outputs(1828));
    layer1_outputs(2535) <= not(layer0_outputs(1478));
    layer1_outputs(2536) <= not(layer0_outputs(3445)) or (layer0_outputs(1021));
    layer1_outputs(2537) <= '0';
    layer1_outputs(2538) <= '0';
    layer1_outputs(2539) <= (layer0_outputs(5072)) or (layer0_outputs(3600));
    layer1_outputs(2540) <= (layer0_outputs(3889)) or (layer0_outputs(1861));
    layer1_outputs(2541) <= not((layer0_outputs(950)) or (layer0_outputs(2790)));
    layer1_outputs(2542) <= not(layer0_outputs(3796));
    layer1_outputs(2543) <= '0';
    layer1_outputs(2544) <= not(layer0_outputs(463));
    layer1_outputs(2545) <= '1';
    layer1_outputs(2546) <= not((layer0_outputs(1141)) and (layer0_outputs(2852)));
    layer1_outputs(2547) <= not(layer0_outputs(3672));
    layer1_outputs(2548) <= '1';
    layer1_outputs(2549) <= (layer0_outputs(212)) and not (layer0_outputs(2556));
    layer1_outputs(2550) <= layer0_outputs(4866);
    layer1_outputs(2551) <= '0';
    layer1_outputs(2552) <= not(layer0_outputs(2369));
    layer1_outputs(2553) <= (layer0_outputs(2539)) or (layer0_outputs(2153));
    layer1_outputs(2554) <= (layer0_outputs(964)) and (layer0_outputs(4206));
    layer1_outputs(2555) <= not(layer0_outputs(2285)) or (layer0_outputs(238));
    layer1_outputs(2556) <= (layer0_outputs(1821)) and (layer0_outputs(4316));
    layer1_outputs(2557) <= (layer0_outputs(4984)) and (layer0_outputs(4208));
    layer1_outputs(2558) <= not(layer0_outputs(3640));
    layer1_outputs(2559) <= not((layer0_outputs(2753)) and (layer0_outputs(1961)));
    layer1_outputs(2560) <= '0';
    layer1_outputs(2561) <= '1';
    layer1_outputs(2562) <= '1';
    layer1_outputs(2563) <= '1';
    layer1_outputs(2564) <= '1';
    layer1_outputs(2565) <= not((layer0_outputs(3149)) or (layer0_outputs(138)));
    layer1_outputs(2566) <= not((layer0_outputs(4774)) xor (layer0_outputs(2727)));
    layer1_outputs(2567) <= not(layer0_outputs(621));
    layer1_outputs(2568) <= not(layer0_outputs(827)) or (layer0_outputs(1226));
    layer1_outputs(2569) <= layer0_outputs(3585);
    layer1_outputs(2570) <= (layer0_outputs(2671)) xor (layer0_outputs(1039));
    layer1_outputs(2571) <= not(layer0_outputs(2340)) or (layer0_outputs(56));
    layer1_outputs(2572) <= (layer0_outputs(3896)) and not (layer0_outputs(379));
    layer1_outputs(2573) <= (layer0_outputs(4535)) and (layer0_outputs(1479));
    layer1_outputs(2574) <= (layer0_outputs(1053)) or (layer0_outputs(54));
    layer1_outputs(2575) <= (layer0_outputs(4010)) and not (layer0_outputs(3942));
    layer1_outputs(2576) <= '0';
    layer1_outputs(2577) <= '1';
    layer1_outputs(2578) <= layer0_outputs(679);
    layer1_outputs(2579) <= not(layer0_outputs(3235));
    layer1_outputs(2580) <= '0';
    layer1_outputs(2581) <= '0';
    layer1_outputs(2582) <= (layer0_outputs(1398)) and not (layer0_outputs(3908));
    layer1_outputs(2583) <= layer0_outputs(4432);
    layer1_outputs(2584) <= '1';
    layer1_outputs(2585) <= (layer0_outputs(747)) xor (layer0_outputs(4331));
    layer1_outputs(2586) <= (layer0_outputs(862)) and (layer0_outputs(1478));
    layer1_outputs(2587) <= (layer0_outputs(3248)) or (layer0_outputs(1548));
    layer1_outputs(2588) <= (layer0_outputs(3549)) and not (layer0_outputs(4276));
    layer1_outputs(2589) <= not((layer0_outputs(5117)) and (layer0_outputs(3181)));
    layer1_outputs(2590) <= not(layer0_outputs(4004)) or (layer0_outputs(879));
    layer1_outputs(2591) <= (layer0_outputs(949)) and (layer0_outputs(4956));
    layer1_outputs(2592) <= layer0_outputs(2557);
    layer1_outputs(2593) <= (layer0_outputs(170)) and not (layer0_outputs(1733));
    layer1_outputs(2594) <= not(layer0_outputs(806)) or (layer0_outputs(2399));
    layer1_outputs(2595) <= '0';
    layer1_outputs(2596) <= (layer0_outputs(645)) and (layer0_outputs(3001));
    layer1_outputs(2597) <= (layer0_outputs(4342)) and not (layer0_outputs(3110));
    layer1_outputs(2598) <= '0';
    layer1_outputs(2599) <= not(layer0_outputs(662));
    layer1_outputs(2600) <= not(layer0_outputs(3800));
    layer1_outputs(2601) <= (layer0_outputs(523)) and not (layer0_outputs(4666));
    layer1_outputs(2602) <= not(layer0_outputs(5093)) or (layer0_outputs(990));
    layer1_outputs(2603) <= not(layer0_outputs(4016));
    layer1_outputs(2604) <= (layer0_outputs(4007)) or (layer0_outputs(4914));
    layer1_outputs(2605) <= not((layer0_outputs(2675)) and (layer0_outputs(4486)));
    layer1_outputs(2606) <= '1';
    layer1_outputs(2607) <= not(layer0_outputs(1476));
    layer1_outputs(2608) <= '1';
    layer1_outputs(2609) <= not(layer0_outputs(4044));
    layer1_outputs(2610) <= (layer0_outputs(1678)) and not (layer0_outputs(913));
    layer1_outputs(2611) <= '1';
    layer1_outputs(2612) <= not(layer0_outputs(4577)) or (layer0_outputs(198));
    layer1_outputs(2613) <= (layer0_outputs(1148)) or (layer0_outputs(257));
    layer1_outputs(2614) <= '0';
    layer1_outputs(2615) <= '0';
    layer1_outputs(2616) <= not(layer0_outputs(181)) or (layer0_outputs(3437));
    layer1_outputs(2617) <= not(layer0_outputs(1150));
    layer1_outputs(2618) <= not((layer0_outputs(1366)) or (layer0_outputs(2463)));
    layer1_outputs(2619) <= not((layer0_outputs(1255)) xor (layer0_outputs(262)));
    layer1_outputs(2620) <= (layer0_outputs(3691)) and (layer0_outputs(505));
    layer1_outputs(2621) <= layer0_outputs(3423);
    layer1_outputs(2622) <= '1';
    layer1_outputs(2623) <= (layer0_outputs(3364)) and not (layer0_outputs(2217));
    layer1_outputs(2624) <= not((layer0_outputs(2662)) or (layer0_outputs(1427)));
    layer1_outputs(2625) <= '1';
    layer1_outputs(2626) <= '1';
    layer1_outputs(2627) <= '1';
    layer1_outputs(2628) <= '0';
    layer1_outputs(2629) <= (layer0_outputs(3876)) or (layer0_outputs(3966));
    layer1_outputs(2630) <= '1';
    layer1_outputs(2631) <= (layer0_outputs(1514)) or (layer0_outputs(4955));
    layer1_outputs(2632) <= '1';
    layer1_outputs(2633) <= '1';
    layer1_outputs(2634) <= not((layer0_outputs(3802)) and (layer0_outputs(4776)));
    layer1_outputs(2635) <= not(layer0_outputs(3464)) or (layer0_outputs(297));
    layer1_outputs(2636) <= (layer0_outputs(536)) and not (layer0_outputs(2270));
    layer1_outputs(2637) <= layer0_outputs(4787);
    layer1_outputs(2638) <= '1';
    layer1_outputs(2639) <= '0';
    layer1_outputs(2640) <= (layer0_outputs(1974)) or (layer0_outputs(2168));
    layer1_outputs(2641) <= '0';
    layer1_outputs(2642) <= not((layer0_outputs(1579)) and (layer0_outputs(1348)));
    layer1_outputs(2643) <= layer0_outputs(897);
    layer1_outputs(2644) <= not(layer0_outputs(1154));
    layer1_outputs(2645) <= not((layer0_outputs(1918)) and (layer0_outputs(1538)));
    layer1_outputs(2646) <= not(layer0_outputs(2171)) or (layer0_outputs(1971));
    layer1_outputs(2647) <= '1';
    layer1_outputs(2648) <= layer0_outputs(3365);
    layer1_outputs(2649) <= (layer0_outputs(118)) and not (layer0_outputs(5105));
    layer1_outputs(2650) <= (layer0_outputs(5080)) and not (layer0_outputs(4883));
    layer1_outputs(2651) <= '0';
    layer1_outputs(2652) <= '1';
    layer1_outputs(2653) <= layer0_outputs(1924);
    layer1_outputs(2654) <= not(layer0_outputs(2995)) or (layer0_outputs(4472));
    layer1_outputs(2655) <= not(layer0_outputs(3961)) or (layer0_outputs(186));
    layer1_outputs(2656) <= not(layer0_outputs(4297));
    layer1_outputs(2657) <= layer0_outputs(2602);
    layer1_outputs(2658) <= not(layer0_outputs(4866));
    layer1_outputs(2659) <= '1';
    layer1_outputs(2660) <= '1';
    layer1_outputs(2661) <= not((layer0_outputs(2664)) and (layer0_outputs(23)));
    layer1_outputs(2662) <= (layer0_outputs(1019)) and not (layer0_outputs(1462));
    layer1_outputs(2663) <= (layer0_outputs(3037)) and (layer0_outputs(973));
    layer1_outputs(2664) <= not(layer0_outputs(370)) or (layer0_outputs(551));
    layer1_outputs(2665) <= not((layer0_outputs(2884)) or (layer0_outputs(3741)));
    layer1_outputs(2666) <= layer0_outputs(308);
    layer1_outputs(2667) <= (layer0_outputs(3051)) and not (layer0_outputs(1593));
    layer1_outputs(2668) <= (layer0_outputs(2978)) and not (layer0_outputs(3073));
    layer1_outputs(2669) <= not(layer0_outputs(5030)) or (layer0_outputs(214));
    layer1_outputs(2670) <= '1';
    layer1_outputs(2671) <= '1';
    layer1_outputs(2672) <= layer0_outputs(3782);
    layer1_outputs(2673) <= '0';
    layer1_outputs(2674) <= not((layer0_outputs(109)) xor (layer0_outputs(3883)));
    layer1_outputs(2675) <= not(layer0_outputs(2626)) or (layer0_outputs(927));
    layer1_outputs(2676) <= not(layer0_outputs(4385)) or (layer0_outputs(3501));
    layer1_outputs(2677) <= '1';
    layer1_outputs(2678) <= '1';
    layer1_outputs(2679) <= not((layer0_outputs(2031)) or (layer0_outputs(4823)));
    layer1_outputs(2680) <= '1';
    layer1_outputs(2681) <= (layer0_outputs(3365)) and not (layer0_outputs(4650));
    layer1_outputs(2682) <= layer0_outputs(223);
    layer1_outputs(2683) <= (layer0_outputs(2657)) and not (layer0_outputs(294));
    layer1_outputs(2684) <= '0';
    layer1_outputs(2685) <= (layer0_outputs(3494)) and not (layer0_outputs(1828));
    layer1_outputs(2686) <= '1';
    layer1_outputs(2687) <= '0';
    layer1_outputs(2688) <= (layer0_outputs(4414)) or (layer0_outputs(167));
    layer1_outputs(2689) <= layer0_outputs(4302);
    layer1_outputs(2690) <= not(layer0_outputs(2950));
    layer1_outputs(2691) <= not((layer0_outputs(276)) and (layer0_outputs(3881)));
    layer1_outputs(2692) <= not(layer0_outputs(2702)) or (layer0_outputs(4934));
    layer1_outputs(2693) <= '1';
    layer1_outputs(2694) <= not(layer0_outputs(3432)) or (layer0_outputs(3235));
    layer1_outputs(2695) <= layer0_outputs(58);
    layer1_outputs(2696) <= '0';
    layer1_outputs(2697) <= '1';
    layer1_outputs(2698) <= not(layer0_outputs(1621));
    layer1_outputs(2699) <= not(layer0_outputs(874)) or (layer0_outputs(1119));
    layer1_outputs(2700) <= not(layer0_outputs(1642));
    layer1_outputs(2701) <= not((layer0_outputs(4808)) and (layer0_outputs(3203)));
    layer1_outputs(2702) <= not(layer0_outputs(1456)) or (layer0_outputs(2934));
    layer1_outputs(2703) <= not(layer0_outputs(3103)) or (layer0_outputs(3142));
    layer1_outputs(2704) <= '1';
    layer1_outputs(2705) <= not(layer0_outputs(1912));
    layer1_outputs(2706) <= not((layer0_outputs(3396)) and (layer0_outputs(763)));
    layer1_outputs(2707) <= '1';
    layer1_outputs(2708) <= (layer0_outputs(2781)) and (layer0_outputs(1454));
    layer1_outputs(2709) <= not(layer0_outputs(2659));
    layer1_outputs(2710) <= (layer0_outputs(1588)) and not (layer0_outputs(4851));
    layer1_outputs(2711) <= '0';
    layer1_outputs(2712) <= not(layer0_outputs(1757)) or (layer0_outputs(2782));
    layer1_outputs(2713) <= '1';
    layer1_outputs(2714) <= '1';
    layer1_outputs(2715) <= not(layer0_outputs(4277));
    layer1_outputs(2716) <= (layer0_outputs(1440)) xor (layer0_outputs(4857));
    layer1_outputs(2717) <= layer0_outputs(3647);
    layer1_outputs(2718) <= not(layer0_outputs(704));
    layer1_outputs(2719) <= not(layer0_outputs(998));
    layer1_outputs(2720) <= (layer0_outputs(4589)) and not (layer0_outputs(977));
    layer1_outputs(2721) <= layer0_outputs(3362);
    layer1_outputs(2722) <= not(layer0_outputs(758));
    layer1_outputs(2723) <= (layer0_outputs(3606)) and (layer0_outputs(3000));
    layer1_outputs(2724) <= not((layer0_outputs(299)) and (layer0_outputs(251)));
    layer1_outputs(2725) <= '0';
    layer1_outputs(2726) <= layer0_outputs(1967);
    layer1_outputs(2727) <= not((layer0_outputs(1612)) and (layer0_outputs(3828)));
    layer1_outputs(2728) <= '0';
    layer1_outputs(2729) <= '0';
    layer1_outputs(2730) <= (layer0_outputs(3684)) and not (layer0_outputs(2509));
    layer1_outputs(2731) <= (layer0_outputs(3602)) and not (layer0_outputs(1040));
    layer1_outputs(2732) <= '1';
    layer1_outputs(2733) <= layer0_outputs(4795);
    layer1_outputs(2734) <= not((layer0_outputs(3097)) and (layer0_outputs(3438)));
    layer1_outputs(2735) <= not(layer0_outputs(4463)) or (layer0_outputs(4184));
    layer1_outputs(2736) <= '1';
    layer1_outputs(2737) <= '0';
    layer1_outputs(2738) <= (layer0_outputs(3519)) or (layer0_outputs(3699));
    layer1_outputs(2739) <= layer0_outputs(1046);
    layer1_outputs(2740) <= not(layer0_outputs(2695));
    layer1_outputs(2741) <= not(layer0_outputs(1914)) or (layer0_outputs(2663));
    layer1_outputs(2742) <= '0';
    layer1_outputs(2743) <= not(layer0_outputs(1126));
    layer1_outputs(2744) <= layer0_outputs(1492);
    layer1_outputs(2745) <= not(layer0_outputs(2369)) or (layer0_outputs(2996));
    layer1_outputs(2746) <= (layer0_outputs(1975)) and (layer0_outputs(876));
    layer1_outputs(2747) <= (layer0_outputs(1430)) or (layer0_outputs(3088));
    layer1_outputs(2748) <= '1';
    layer1_outputs(2749) <= '1';
    layer1_outputs(2750) <= '1';
    layer1_outputs(2751) <= (layer0_outputs(1285)) and not (layer0_outputs(1147));
    layer1_outputs(2752) <= not(layer0_outputs(1712));
    layer1_outputs(2753) <= not((layer0_outputs(4270)) or (layer0_outputs(1406)));
    layer1_outputs(2754) <= (layer0_outputs(421)) or (layer0_outputs(3121));
    layer1_outputs(2755) <= '0';
    layer1_outputs(2756) <= (layer0_outputs(1278)) and (layer0_outputs(4358));
    layer1_outputs(2757) <= not(layer0_outputs(4027));
    layer1_outputs(2758) <= not((layer0_outputs(4689)) or (layer0_outputs(3417)));
    layer1_outputs(2759) <= (layer0_outputs(1080)) and (layer0_outputs(715));
    layer1_outputs(2760) <= not((layer0_outputs(1378)) and (layer0_outputs(4489)));
    layer1_outputs(2761) <= not((layer0_outputs(376)) and (layer0_outputs(4413)));
    layer1_outputs(2762) <= (layer0_outputs(1064)) and (layer0_outputs(3782));
    layer1_outputs(2763) <= not(layer0_outputs(3901));
    layer1_outputs(2764) <= '1';
    layer1_outputs(2765) <= not((layer0_outputs(40)) and (layer0_outputs(1581)));
    layer1_outputs(2766) <= '0';
    layer1_outputs(2767) <= (layer0_outputs(275)) and (layer0_outputs(678));
    layer1_outputs(2768) <= '0';
    layer1_outputs(2769) <= '1';
    layer1_outputs(2770) <= not(layer0_outputs(5084));
    layer1_outputs(2771) <= layer0_outputs(2232);
    layer1_outputs(2772) <= '1';
    layer1_outputs(2773) <= layer0_outputs(4974);
    layer1_outputs(2774) <= not((layer0_outputs(811)) and (layer0_outputs(2438)));
    layer1_outputs(2775) <= '0';
    layer1_outputs(2776) <= (layer0_outputs(3557)) and not (layer0_outputs(154));
    layer1_outputs(2777) <= (layer0_outputs(1504)) and not (layer0_outputs(4035));
    layer1_outputs(2778) <= layer0_outputs(3080);
    layer1_outputs(2779) <= '0';
    layer1_outputs(2780) <= layer0_outputs(1602);
    layer1_outputs(2781) <= not(layer0_outputs(4363)) or (layer0_outputs(102));
    layer1_outputs(2782) <= (layer0_outputs(487)) and (layer0_outputs(3083));
    layer1_outputs(2783) <= '0';
    layer1_outputs(2784) <= not((layer0_outputs(3079)) or (layer0_outputs(3937)));
    layer1_outputs(2785) <= (layer0_outputs(4877)) or (layer0_outputs(1929));
    layer1_outputs(2786) <= layer0_outputs(2073);
    layer1_outputs(2787) <= not(layer0_outputs(3325)) or (layer0_outputs(3547));
    layer1_outputs(2788) <= not(layer0_outputs(1382));
    layer1_outputs(2789) <= '0';
    layer1_outputs(2790) <= (layer0_outputs(4560)) and not (layer0_outputs(2701));
    layer1_outputs(2791) <= (layer0_outputs(3925)) and (layer0_outputs(4925));
    layer1_outputs(2792) <= (layer0_outputs(1736)) or (layer0_outputs(633));
    layer1_outputs(2793) <= not(layer0_outputs(1799)) or (layer0_outputs(2975));
    layer1_outputs(2794) <= (layer0_outputs(4929)) or (layer0_outputs(1060));
    layer1_outputs(2795) <= layer0_outputs(4955);
    layer1_outputs(2796) <= (layer0_outputs(2180)) and not (layer0_outputs(4674));
    layer1_outputs(2797) <= '0';
    layer1_outputs(2798) <= '1';
    layer1_outputs(2799) <= (layer0_outputs(3906)) or (layer0_outputs(1633));
    layer1_outputs(2800) <= (layer0_outputs(1752)) or (layer0_outputs(2480));
    layer1_outputs(2801) <= layer0_outputs(3571);
    layer1_outputs(2802) <= (layer0_outputs(3231)) and (layer0_outputs(468));
    layer1_outputs(2803) <= layer0_outputs(3580);
    layer1_outputs(2804) <= not((layer0_outputs(1279)) and (layer0_outputs(3210)));
    layer1_outputs(2805) <= not(layer0_outputs(1496));
    layer1_outputs(2806) <= '1';
    layer1_outputs(2807) <= not((layer0_outputs(4017)) and (layer0_outputs(549)));
    layer1_outputs(2808) <= (layer0_outputs(184)) xor (layer0_outputs(2632));
    layer1_outputs(2809) <= '1';
    layer1_outputs(2810) <= '1';
    layer1_outputs(2811) <= not(layer0_outputs(574)) or (layer0_outputs(4369));
    layer1_outputs(2812) <= not((layer0_outputs(3767)) xor (layer0_outputs(2615)));
    layer1_outputs(2813) <= (layer0_outputs(4064)) or (layer0_outputs(4598));
    layer1_outputs(2814) <= '1';
    layer1_outputs(2815) <= not(layer0_outputs(4981));
    layer1_outputs(2816) <= not(layer0_outputs(3096)) or (layer0_outputs(2460));
    layer1_outputs(2817) <= '0';
    layer1_outputs(2818) <= (layer0_outputs(676)) xor (layer0_outputs(4415));
    layer1_outputs(2819) <= not((layer0_outputs(2357)) or (layer0_outputs(2540)));
    layer1_outputs(2820) <= (layer0_outputs(1298)) and not (layer0_outputs(4003));
    layer1_outputs(2821) <= not(layer0_outputs(4426));
    layer1_outputs(2822) <= not(layer0_outputs(585));
    layer1_outputs(2823) <= layer0_outputs(4351);
    layer1_outputs(2824) <= layer0_outputs(4235);
    layer1_outputs(2825) <= (layer0_outputs(2546)) or (layer0_outputs(3480));
    layer1_outputs(2826) <= not((layer0_outputs(943)) or (layer0_outputs(691)));
    layer1_outputs(2827) <= not(layer0_outputs(2225));
    layer1_outputs(2828) <= (layer0_outputs(3076)) and not (layer0_outputs(5057));
    layer1_outputs(2829) <= not((layer0_outputs(4848)) or (layer0_outputs(4753)));
    layer1_outputs(2830) <= not((layer0_outputs(277)) or (layer0_outputs(4670)));
    layer1_outputs(2831) <= layer0_outputs(1779);
    layer1_outputs(2832) <= '1';
    layer1_outputs(2833) <= (layer0_outputs(3461)) and (layer0_outputs(2086));
    layer1_outputs(2834) <= layer0_outputs(4675);
    layer1_outputs(2835) <= '0';
    layer1_outputs(2836) <= layer0_outputs(4877);
    layer1_outputs(2837) <= '0';
    layer1_outputs(2838) <= '0';
    layer1_outputs(2839) <= not(layer0_outputs(2459));
    layer1_outputs(2840) <= '1';
    layer1_outputs(2841) <= '1';
    layer1_outputs(2842) <= not(layer0_outputs(2598)) or (layer0_outputs(3023));
    layer1_outputs(2843) <= not(layer0_outputs(1375));
    layer1_outputs(2844) <= '1';
    layer1_outputs(2845) <= (layer0_outputs(1223)) and (layer0_outputs(1054));
    layer1_outputs(2846) <= layer0_outputs(748);
    layer1_outputs(2847) <= '0';
    layer1_outputs(2848) <= layer0_outputs(3382);
    layer1_outputs(2849) <= '1';
    layer1_outputs(2850) <= not(layer0_outputs(1553));
    layer1_outputs(2851) <= layer0_outputs(2137);
    layer1_outputs(2852) <= not(layer0_outputs(5111));
    layer1_outputs(2853) <= layer0_outputs(1316);
    layer1_outputs(2854) <= '1';
    layer1_outputs(2855) <= (layer0_outputs(72)) and not (layer0_outputs(3843));
    layer1_outputs(2856) <= not(layer0_outputs(5));
    layer1_outputs(2857) <= (layer0_outputs(1644)) and not (layer0_outputs(4383));
    layer1_outputs(2858) <= not((layer0_outputs(1419)) and (layer0_outputs(4242)));
    layer1_outputs(2859) <= layer0_outputs(2586);
    layer1_outputs(2860) <= '1';
    layer1_outputs(2861) <= not((layer0_outputs(2203)) or (layer0_outputs(1852)));
    layer1_outputs(2862) <= (layer0_outputs(83)) and not (layer0_outputs(1461));
    layer1_outputs(2863) <= '0';
    layer1_outputs(2864) <= not((layer0_outputs(2348)) or (layer0_outputs(91)));
    layer1_outputs(2865) <= not((layer0_outputs(1517)) and (layer0_outputs(3713)));
    layer1_outputs(2866) <= (layer0_outputs(4313)) and not (layer0_outputs(213));
    layer1_outputs(2867) <= (layer0_outputs(2494)) or (layer0_outputs(3924));
    layer1_outputs(2868) <= layer0_outputs(413);
    layer1_outputs(2869) <= not(layer0_outputs(2769)) or (layer0_outputs(2174));
    layer1_outputs(2870) <= layer0_outputs(4377);
    layer1_outputs(2871) <= not((layer0_outputs(3306)) and (layer0_outputs(4209)));
    layer1_outputs(2872) <= '0';
    layer1_outputs(2873) <= (layer0_outputs(1793)) and not (layer0_outputs(4005));
    layer1_outputs(2874) <= layer0_outputs(4930);
    layer1_outputs(2875) <= '1';
    layer1_outputs(2876) <= (layer0_outputs(1164)) and not (layer0_outputs(2064));
    layer1_outputs(2877) <= not((layer0_outputs(2958)) and (layer0_outputs(4929)));
    layer1_outputs(2878) <= not((layer0_outputs(1684)) and (layer0_outputs(2453)));
    layer1_outputs(2879) <= not(layer0_outputs(2313)) or (layer0_outputs(235));
    layer1_outputs(2880) <= '1';
    layer1_outputs(2881) <= layer0_outputs(4600);
    layer1_outputs(2882) <= (layer0_outputs(510)) and (layer0_outputs(1264));
    layer1_outputs(2883) <= (layer0_outputs(3666)) and not (layer0_outputs(951));
    layer1_outputs(2884) <= not(layer0_outputs(3504)) or (layer0_outputs(3288));
    layer1_outputs(2885) <= not(layer0_outputs(2711)) or (layer0_outputs(4139));
    layer1_outputs(2886) <= '1';
    layer1_outputs(2887) <= not(layer0_outputs(3090)) or (layer0_outputs(4702));
    layer1_outputs(2888) <= '1';
    layer1_outputs(2889) <= not((layer0_outputs(3076)) or (layer0_outputs(2675)));
    layer1_outputs(2890) <= (layer0_outputs(1807)) and not (layer0_outputs(484));
    layer1_outputs(2891) <= '1';
    layer1_outputs(2892) <= not((layer0_outputs(132)) or (layer0_outputs(195)));
    layer1_outputs(2893) <= '1';
    layer1_outputs(2894) <= '0';
    layer1_outputs(2895) <= layer0_outputs(2811);
    layer1_outputs(2896) <= not(layer0_outputs(4123));
    layer1_outputs(2897) <= (layer0_outputs(2583)) and not (layer0_outputs(5042));
    layer1_outputs(2898) <= not(layer0_outputs(5063)) or (layer0_outputs(3563));
    layer1_outputs(2899) <= (layer0_outputs(967)) or (layer0_outputs(4467));
    layer1_outputs(2900) <= layer0_outputs(4042);
    layer1_outputs(2901) <= not((layer0_outputs(3329)) and (layer0_outputs(4105)));
    layer1_outputs(2902) <= '1';
    layer1_outputs(2903) <= '1';
    layer1_outputs(2904) <= not(layer0_outputs(4380)) or (layer0_outputs(3420));
    layer1_outputs(2905) <= (layer0_outputs(2389)) or (layer0_outputs(4762));
    layer1_outputs(2906) <= layer0_outputs(3458);
    layer1_outputs(2907) <= not(layer0_outputs(4595));
    layer1_outputs(2908) <= not(layer0_outputs(955)) or (layer0_outputs(4412));
    layer1_outputs(2909) <= layer0_outputs(3544);
    layer1_outputs(2910) <= (layer0_outputs(994)) and not (layer0_outputs(3609));
    layer1_outputs(2911) <= not(layer0_outputs(2413));
    layer1_outputs(2912) <= not(layer0_outputs(2362));
    layer1_outputs(2913) <= not((layer0_outputs(1037)) and (layer0_outputs(807)));
    layer1_outputs(2914) <= not(layer0_outputs(2713));
    layer1_outputs(2915) <= '1';
    layer1_outputs(2916) <= not((layer0_outputs(4664)) or (layer0_outputs(3433)));
    layer1_outputs(2917) <= layer0_outputs(1120);
    layer1_outputs(2918) <= (layer0_outputs(1434)) and (layer0_outputs(582));
    layer1_outputs(2919) <= not((layer0_outputs(3871)) or (layer0_outputs(4725)));
    layer1_outputs(2920) <= (layer0_outputs(1188)) and (layer0_outputs(2482));
    layer1_outputs(2921) <= not((layer0_outputs(4878)) and (layer0_outputs(4604)));
    layer1_outputs(2922) <= (layer0_outputs(3923)) and not (layer0_outputs(1404));
    layer1_outputs(2923) <= '1';
    layer1_outputs(2924) <= not((layer0_outputs(2548)) or (layer0_outputs(193)));
    layer1_outputs(2925) <= '1';
    layer1_outputs(2926) <= '0';
    layer1_outputs(2927) <= (layer0_outputs(2093)) and (layer0_outputs(1523));
    layer1_outputs(2928) <= not(layer0_outputs(1933));
    layer1_outputs(2929) <= '1';
    layer1_outputs(2930) <= not(layer0_outputs(3483)) or (layer0_outputs(2905));
    layer1_outputs(2931) <= not(layer0_outputs(1197)) or (layer0_outputs(2442));
    layer1_outputs(2932) <= (layer0_outputs(2030)) and (layer0_outputs(1354));
    layer1_outputs(2933) <= '1';
    layer1_outputs(2934) <= not((layer0_outputs(3146)) and (layer0_outputs(65)));
    layer1_outputs(2935) <= not((layer0_outputs(4069)) and (layer0_outputs(3643)));
    layer1_outputs(2936) <= (layer0_outputs(4549)) and not (layer0_outputs(2518));
    layer1_outputs(2937) <= (layer0_outputs(4604)) and (layer0_outputs(2265));
    layer1_outputs(2938) <= not(layer0_outputs(4803)) or (layer0_outputs(3776));
    layer1_outputs(2939) <= not((layer0_outputs(5055)) or (layer0_outputs(1622)));
    layer1_outputs(2940) <= (layer0_outputs(4275)) xor (layer0_outputs(4208));
    layer1_outputs(2941) <= '1';
    layer1_outputs(2942) <= not(layer0_outputs(2298)) or (layer0_outputs(1169));
    layer1_outputs(2943) <= not(layer0_outputs(4398)) or (layer0_outputs(2774));
    layer1_outputs(2944) <= (layer0_outputs(3555)) and (layer0_outputs(1798));
    layer1_outputs(2945) <= '0';
    layer1_outputs(2946) <= '1';
    layer1_outputs(2947) <= not(layer0_outputs(2716));
    layer1_outputs(2948) <= (layer0_outputs(3425)) or (layer0_outputs(4976));
    layer1_outputs(2949) <= layer0_outputs(2190);
    layer1_outputs(2950) <= not(layer0_outputs(735)) or (layer0_outputs(4546));
    layer1_outputs(2951) <= layer0_outputs(888);
    layer1_outputs(2952) <= (layer0_outputs(5027)) and (layer0_outputs(375));
    layer1_outputs(2953) <= layer0_outputs(5056);
    layer1_outputs(2954) <= not(layer0_outputs(1667));
    layer1_outputs(2955) <= not(layer0_outputs(3675)) or (layer0_outputs(4843));
    layer1_outputs(2956) <= '1';
    layer1_outputs(2957) <= '1';
    layer1_outputs(2958) <= (layer0_outputs(180)) and not (layer0_outputs(1564));
    layer1_outputs(2959) <= '1';
    layer1_outputs(2960) <= not(layer0_outputs(1109)) or (layer0_outputs(4435));
    layer1_outputs(2961) <= not(layer0_outputs(3024)) or (layer0_outputs(2630));
    layer1_outputs(2962) <= '1';
    layer1_outputs(2963) <= not(layer0_outputs(3810)) or (layer0_outputs(1634));
    layer1_outputs(2964) <= layer0_outputs(1518);
    layer1_outputs(2965) <= not((layer0_outputs(3987)) or (layer0_outputs(3923)));
    layer1_outputs(2966) <= not(layer0_outputs(2092));
    layer1_outputs(2967) <= (layer0_outputs(4029)) and (layer0_outputs(4485));
    layer1_outputs(2968) <= not(layer0_outputs(4222));
    layer1_outputs(2969) <= layer0_outputs(811);
    layer1_outputs(2970) <= not((layer0_outputs(2245)) and (layer0_outputs(2107)));
    layer1_outputs(2971) <= not((layer0_outputs(4630)) xor (layer0_outputs(4063)));
    layer1_outputs(2972) <= (layer0_outputs(2761)) and not (layer0_outputs(2294));
    layer1_outputs(2973) <= not(layer0_outputs(2122)) or (layer0_outputs(4840));
    layer1_outputs(2974) <= '1';
    layer1_outputs(2975) <= layer0_outputs(4549);
    layer1_outputs(2976) <= '0';
    layer1_outputs(2977) <= (layer0_outputs(2437)) and (layer0_outputs(4909));
    layer1_outputs(2978) <= layer0_outputs(4026);
    layer1_outputs(2979) <= (layer0_outputs(3744)) and not (layer0_outputs(5110));
    layer1_outputs(2980) <= not((layer0_outputs(1527)) and (layer0_outputs(3932)));
    layer1_outputs(2981) <= '0';
    layer1_outputs(2982) <= (layer0_outputs(1300)) or (layer0_outputs(3715));
    layer1_outputs(2983) <= not((layer0_outputs(1204)) xor (layer0_outputs(4896)));
    layer1_outputs(2984) <= (layer0_outputs(906)) and (layer0_outputs(1938));
    layer1_outputs(2985) <= not((layer0_outputs(2840)) and (layer0_outputs(4870)));
    layer1_outputs(2986) <= not(layer0_outputs(4967));
    layer1_outputs(2987) <= (layer0_outputs(4804)) xor (layer0_outputs(1913));
    layer1_outputs(2988) <= '0';
    layer1_outputs(2989) <= not((layer0_outputs(4879)) and (layer0_outputs(4846)));
    layer1_outputs(2990) <= layer0_outputs(3046);
    layer1_outputs(2991) <= not((layer0_outputs(444)) and (layer0_outputs(177)));
    layer1_outputs(2992) <= '1';
    layer1_outputs(2993) <= '1';
    layer1_outputs(2994) <= layer0_outputs(3944);
    layer1_outputs(2995) <= not((layer0_outputs(1937)) and (layer0_outputs(1137)));
    layer1_outputs(2996) <= '1';
    layer1_outputs(2997) <= not((layer0_outputs(2920)) or (layer0_outputs(1878)));
    layer1_outputs(2998) <= not(layer0_outputs(5012));
    layer1_outputs(2999) <= (layer0_outputs(4226)) and not (layer0_outputs(226));
    layer1_outputs(3000) <= '0';
    layer1_outputs(3001) <= '1';
    layer1_outputs(3002) <= not(layer0_outputs(2191)) or (layer0_outputs(524));
    layer1_outputs(3003) <= '1';
    layer1_outputs(3004) <= not((layer0_outputs(497)) and (layer0_outputs(2755)));
    layer1_outputs(3005) <= not(layer0_outputs(3670)) or (layer0_outputs(4238));
    layer1_outputs(3006) <= '0';
    layer1_outputs(3007) <= (layer0_outputs(4716)) and not (layer0_outputs(1522));
    layer1_outputs(3008) <= '0';
    layer1_outputs(3009) <= (layer0_outputs(5047)) or (layer0_outputs(2333));
    layer1_outputs(3010) <= not((layer0_outputs(780)) and (layer0_outputs(4081)));
    layer1_outputs(3011) <= (layer0_outputs(4884)) and not (layer0_outputs(1233));
    layer1_outputs(3012) <= not(layer0_outputs(675)) or (layer0_outputs(2908));
    layer1_outputs(3013) <= (layer0_outputs(1013)) and (layer0_outputs(70));
    layer1_outputs(3014) <= not((layer0_outputs(4344)) or (layer0_outputs(0)));
    layer1_outputs(3015) <= (layer0_outputs(485)) and (layer0_outputs(2352));
    layer1_outputs(3016) <= '0';
    layer1_outputs(3017) <= (layer0_outputs(739)) and (layer0_outputs(3467));
    layer1_outputs(3018) <= (layer0_outputs(4738)) and not (layer0_outputs(4133));
    layer1_outputs(3019) <= '1';
    layer1_outputs(3020) <= not((layer0_outputs(4668)) and (layer0_outputs(359)));
    layer1_outputs(3021) <= '0';
    layer1_outputs(3022) <= not(layer0_outputs(5046));
    layer1_outputs(3023) <= (layer0_outputs(3617)) and not (layer0_outputs(2155));
    layer1_outputs(3024) <= not(layer0_outputs(50)) or (layer0_outputs(2426));
    layer1_outputs(3025) <= layer0_outputs(3865);
    layer1_outputs(3026) <= '0';
    layer1_outputs(3027) <= layer0_outputs(2952);
    layer1_outputs(3028) <= '0';
    layer1_outputs(3029) <= layer0_outputs(1371);
    layer1_outputs(3030) <= layer0_outputs(722);
    layer1_outputs(3031) <= (layer0_outputs(1642)) or (layer0_outputs(4026));
    layer1_outputs(3032) <= not(layer0_outputs(3517));
    layer1_outputs(3033) <= (layer0_outputs(3149)) and not (layer0_outputs(1501));
    layer1_outputs(3034) <= not(layer0_outputs(2778)) or (layer0_outputs(310));
    layer1_outputs(3035) <= (layer0_outputs(1398)) or (layer0_outputs(4824));
    layer1_outputs(3036) <= not(layer0_outputs(3726)) or (layer0_outputs(1956));
    layer1_outputs(3037) <= '1';
    layer1_outputs(3038) <= not((layer0_outputs(349)) and (layer0_outputs(5064)));
    layer1_outputs(3039) <= '1';
    layer1_outputs(3040) <= not(layer0_outputs(4171)) or (layer0_outputs(3915));
    layer1_outputs(3041) <= not((layer0_outputs(1179)) or (layer0_outputs(3749)));
    layer1_outputs(3042) <= (layer0_outputs(4187)) or (layer0_outputs(5043));
    layer1_outputs(3043) <= not((layer0_outputs(756)) and (layer0_outputs(788)));
    layer1_outputs(3044) <= not((layer0_outputs(165)) or (layer0_outputs(4968)));
    layer1_outputs(3045) <= (layer0_outputs(5103)) and not (layer0_outputs(3626));
    layer1_outputs(3046) <= '1';
    layer1_outputs(3047) <= (layer0_outputs(2228)) and not (layer0_outputs(2897));
    layer1_outputs(3048) <= not(layer0_outputs(1199));
    layer1_outputs(3049) <= (layer0_outputs(1684)) and not (layer0_outputs(366));
    layer1_outputs(3050) <= '0';
    layer1_outputs(3051) <= not((layer0_outputs(3322)) and (layer0_outputs(2974)));
    layer1_outputs(3052) <= '0';
    layer1_outputs(3053) <= layer0_outputs(2275);
    layer1_outputs(3054) <= not(layer0_outputs(1192));
    layer1_outputs(3055) <= not((layer0_outputs(3522)) or (layer0_outputs(93)));
    layer1_outputs(3056) <= (layer0_outputs(3419)) and not (layer0_outputs(4694));
    layer1_outputs(3057) <= '0';
    layer1_outputs(3058) <= not((layer0_outputs(4165)) and (layer0_outputs(3054)));
    layer1_outputs(3059) <= not(layer0_outputs(4378));
    layer1_outputs(3060) <= '0';
    layer1_outputs(3061) <= not(layer0_outputs(2781));
    layer1_outputs(3062) <= layer0_outputs(4616);
    layer1_outputs(3063) <= layer0_outputs(2651);
    layer1_outputs(3064) <= (layer0_outputs(3588)) and (layer0_outputs(4964));
    layer1_outputs(3065) <= layer0_outputs(2285);
    layer1_outputs(3066) <= (layer0_outputs(3473)) or (layer0_outputs(4434));
    layer1_outputs(3067) <= not(layer0_outputs(3461)) or (layer0_outputs(1066));
    layer1_outputs(3068) <= '1';
    layer1_outputs(3069) <= not(layer0_outputs(156));
    layer1_outputs(3070) <= layer0_outputs(2456);
    layer1_outputs(3071) <= layer0_outputs(3411);
    layer1_outputs(3072) <= '0';
    layer1_outputs(3073) <= not(layer0_outputs(718)) or (layer0_outputs(1196));
    layer1_outputs(3074) <= not((layer0_outputs(1964)) or (layer0_outputs(1565)));
    layer1_outputs(3075) <= not(layer0_outputs(1057)) or (layer0_outputs(2889));
    layer1_outputs(3076) <= '0';
    layer1_outputs(3077) <= (layer0_outputs(3548)) or (layer0_outputs(3984));
    layer1_outputs(3078) <= not(layer0_outputs(1927));
    layer1_outputs(3079) <= '0';
    layer1_outputs(3080) <= layer0_outputs(3269);
    layer1_outputs(3081) <= '0';
    layer1_outputs(3082) <= '0';
    layer1_outputs(3083) <= (layer0_outputs(5078)) or (layer0_outputs(867));
    layer1_outputs(3084) <= '0';
    layer1_outputs(3085) <= not(layer0_outputs(4893));
    layer1_outputs(3086) <= layer0_outputs(1129);
    layer1_outputs(3087) <= (layer0_outputs(2475)) and not (layer0_outputs(2406));
    layer1_outputs(3088) <= (layer0_outputs(998)) and (layer0_outputs(1547));
    layer1_outputs(3089) <= '1';
    layer1_outputs(3090) <= '1';
    layer1_outputs(3091) <= not((layer0_outputs(1326)) and (layer0_outputs(3761)));
    layer1_outputs(3092) <= (layer0_outputs(1325)) and not (layer0_outputs(2815));
    layer1_outputs(3093) <= layer0_outputs(4807);
    layer1_outputs(3094) <= layer0_outputs(878);
    layer1_outputs(3095) <= not(layer0_outputs(4374));
    layer1_outputs(3096) <= (layer0_outputs(2865)) and not (layer0_outputs(4089));
    layer1_outputs(3097) <= (layer0_outputs(1399)) and not (layer0_outputs(3129));
    layer1_outputs(3098) <= not((layer0_outputs(3710)) and (layer0_outputs(1493)));
    layer1_outputs(3099) <= (layer0_outputs(3268)) and not (layer0_outputs(2695));
    layer1_outputs(3100) <= not((layer0_outputs(4550)) and (layer0_outputs(2543)));
    layer1_outputs(3101) <= '0';
    layer1_outputs(3102) <= (layer0_outputs(1525)) or (layer0_outputs(2202));
    layer1_outputs(3103) <= not(layer0_outputs(3881));
    layer1_outputs(3104) <= not(layer0_outputs(3851));
    layer1_outputs(3105) <= not((layer0_outputs(394)) or (layer0_outputs(2683)));
    layer1_outputs(3106) <= '0';
    layer1_outputs(3107) <= layer0_outputs(3764);
    layer1_outputs(3108) <= (layer0_outputs(4977)) and not (layer0_outputs(1835));
    layer1_outputs(3109) <= '0';
    layer1_outputs(3110) <= '1';
    layer1_outputs(3111) <= not(layer0_outputs(538)) or (layer0_outputs(3877));
    layer1_outputs(3112) <= '1';
    layer1_outputs(3113) <= '1';
    layer1_outputs(3114) <= '0';
    layer1_outputs(3115) <= not((layer0_outputs(5013)) xor (layer0_outputs(334)));
    layer1_outputs(3116) <= not(layer0_outputs(3696));
    layer1_outputs(3117) <= '0';
    layer1_outputs(3118) <= (layer0_outputs(4641)) and not (layer0_outputs(2170));
    layer1_outputs(3119) <= '1';
    layer1_outputs(3120) <= '0';
    layer1_outputs(3121) <= '0';
    layer1_outputs(3122) <= not(layer0_outputs(1865)) or (layer0_outputs(1665));
    layer1_outputs(3123) <= (layer0_outputs(2731)) or (layer0_outputs(46));
    layer1_outputs(3124) <= (layer0_outputs(3293)) or (layer0_outputs(4299));
    layer1_outputs(3125) <= (layer0_outputs(4961)) and not (layer0_outputs(1385));
    layer1_outputs(3126) <= (layer0_outputs(383)) and not (layer0_outputs(4886));
    layer1_outputs(3127) <= not(layer0_outputs(3758)) or (layer0_outputs(974));
    layer1_outputs(3128) <= layer0_outputs(4211);
    layer1_outputs(3129) <= '0';
    layer1_outputs(3130) <= '1';
    layer1_outputs(3131) <= '1';
    layer1_outputs(3132) <= not(layer0_outputs(2436)) or (layer0_outputs(1706));
    layer1_outputs(3133) <= not((layer0_outputs(790)) and (layer0_outputs(4480)));
    layer1_outputs(3134) <= not(layer0_outputs(3038));
    layer1_outputs(3135) <= not(layer0_outputs(4639));
    layer1_outputs(3136) <= layer0_outputs(4965);
    layer1_outputs(3137) <= (layer0_outputs(541)) and not (layer0_outputs(3096));
    layer1_outputs(3138) <= layer0_outputs(4270);
    layer1_outputs(3139) <= '0';
    layer1_outputs(3140) <= '0';
    layer1_outputs(3141) <= not(layer0_outputs(4158));
    layer1_outputs(3142) <= not((layer0_outputs(4244)) and (layer0_outputs(4524)));
    layer1_outputs(3143) <= '1';
    layer1_outputs(3144) <= not(layer0_outputs(4930));
    layer1_outputs(3145) <= '1';
    layer1_outputs(3146) <= (layer0_outputs(2763)) or (layer0_outputs(3654));
    layer1_outputs(3147) <= not((layer0_outputs(1655)) or (layer0_outputs(4081)));
    layer1_outputs(3148) <= not(layer0_outputs(2497));
    layer1_outputs(3149) <= not(layer0_outputs(5038));
    layer1_outputs(3150) <= not((layer0_outputs(2921)) and (layer0_outputs(4566)));
    layer1_outputs(3151) <= '1';
    layer1_outputs(3152) <= not((layer0_outputs(830)) or (layer0_outputs(4536)));
    layer1_outputs(3153) <= '0';
    layer1_outputs(3154) <= (layer0_outputs(4881)) and not (layer0_outputs(797));
    layer1_outputs(3155) <= (layer0_outputs(1115)) and not (layer0_outputs(4340));
    layer1_outputs(3156) <= '0';
    layer1_outputs(3157) <= not((layer0_outputs(1133)) xor (layer0_outputs(3426)));
    layer1_outputs(3158) <= not(layer0_outputs(4328)) or (layer0_outputs(4651));
    layer1_outputs(3159) <= '0';
    layer1_outputs(3160) <= (layer0_outputs(234)) and not (layer0_outputs(5109));
    layer1_outputs(3161) <= (layer0_outputs(4367)) xor (layer0_outputs(5015));
    layer1_outputs(3162) <= '0';
    layer1_outputs(3163) <= not((layer0_outputs(2727)) or (layer0_outputs(2395)));
    layer1_outputs(3164) <= layer0_outputs(2492);
    layer1_outputs(3165) <= '1';
    layer1_outputs(3166) <= layer0_outputs(2271);
    layer1_outputs(3167) <= (layer0_outputs(3334)) and not (layer0_outputs(4894));
    layer1_outputs(3168) <= layer0_outputs(4600);
    layer1_outputs(3169) <= layer0_outputs(3565);
    layer1_outputs(3170) <= not((layer0_outputs(1910)) and (layer0_outputs(1342)));
    layer1_outputs(3171) <= not((layer0_outputs(4661)) and (layer0_outputs(3724)));
    layer1_outputs(3172) <= '1';
    layer1_outputs(3173) <= '0';
    layer1_outputs(3174) <= (layer0_outputs(1144)) or (layer0_outputs(1421));
    layer1_outputs(3175) <= not(layer0_outputs(1372));
    layer1_outputs(3176) <= (layer0_outputs(110)) and not (layer0_outputs(2002));
    layer1_outputs(3177) <= (layer0_outputs(489)) and (layer0_outputs(3659));
    layer1_outputs(3178) <= layer0_outputs(3824);
    layer1_outputs(3179) <= '0';
    layer1_outputs(3180) <= (layer0_outputs(3207)) and not (layer0_outputs(1028));
    layer1_outputs(3181) <= '0';
    layer1_outputs(3182) <= '1';
    layer1_outputs(3183) <= (layer0_outputs(2502)) and not (layer0_outputs(2640));
    layer1_outputs(3184) <= not(layer0_outputs(2162));
    layer1_outputs(3185) <= '0';
    layer1_outputs(3186) <= (layer0_outputs(3408)) and not (layer0_outputs(4513));
    layer1_outputs(3187) <= '0';
    layer1_outputs(3188) <= not(layer0_outputs(4636)) or (layer0_outputs(1944));
    layer1_outputs(3189) <= not(layer0_outputs(3017));
    layer1_outputs(3190) <= '0';
    layer1_outputs(3191) <= (layer0_outputs(5032)) and not (layer0_outputs(3369));
    layer1_outputs(3192) <= (layer0_outputs(4151)) or (layer0_outputs(2051));
    layer1_outputs(3193) <= (layer0_outputs(3472)) and not (layer0_outputs(427));
    layer1_outputs(3194) <= layer0_outputs(4693);
    layer1_outputs(3195) <= not(layer0_outputs(2061)) or (layer0_outputs(586));
    layer1_outputs(3196) <= '0';
    layer1_outputs(3197) <= '0';
    layer1_outputs(3198) <= '0';
    layer1_outputs(3199) <= not(layer0_outputs(1389)) or (layer0_outputs(4911));
    layer1_outputs(3200) <= (layer0_outputs(911)) or (layer0_outputs(2152));
    layer1_outputs(3201) <= not((layer0_outputs(3535)) and (layer0_outputs(4842)));
    layer1_outputs(3202) <= (layer0_outputs(1784)) or (layer0_outputs(3550));
    layer1_outputs(3203) <= (layer0_outputs(1735)) and not (layer0_outputs(3304));
    layer1_outputs(3204) <= '0';
    layer1_outputs(3205) <= (layer0_outputs(2414)) and not (layer0_outputs(3184));
    layer1_outputs(3206) <= not(layer0_outputs(3719)) or (layer0_outputs(2993));
    layer1_outputs(3207) <= '0';
    layer1_outputs(3208) <= not(layer0_outputs(3344)) or (layer0_outputs(2287));
    layer1_outputs(3209) <= (layer0_outputs(1409)) and not (layer0_outputs(265));
    layer1_outputs(3210) <= (layer0_outputs(944)) or (layer0_outputs(1205));
    layer1_outputs(3211) <= '1';
    layer1_outputs(3212) <= '0';
    layer1_outputs(3213) <= not((layer0_outputs(2224)) and (layer0_outputs(345)));
    layer1_outputs(3214) <= not((layer0_outputs(4018)) or (layer0_outputs(4219)));
    layer1_outputs(3215) <= '1';
    layer1_outputs(3216) <= (layer0_outputs(3332)) or (layer0_outputs(4239));
    layer1_outputs(3217) <= not((layer0_outputs(3722)) and (layer0_outputs(1582)));
    layer1_outputs(3218) <= (layer0_outputs(4963)) and (layer0_outputs(1925));
    layer1_outputs(3219) <= (layer0_outputs(2988)) and not (layer0_outputs(360));
    layer1_outputs(3220) <= (layer0_outputs(3750)) and not (layer0_outputs(4765));
    layer1_outputs(3221) <= not(layer0_outputs(1499)) or (layer0_outputs(1396));
    layer1_outputs(3222) <= '0';
    layer1_outputs(3223) <= not((layer0_outputs(4891)) or (layer0_outputs(866)));
    layer1_outputs(3224) <= (layer0_outputs(4453)) or (layer0_outputs(747));
    layer1_outputs(3225) <= (layer0_outputs(4659)) and not (layer0_outputs(3952));
    layer1_outputs(3226) <= not(layer0_outputs(3834));
    layer1_outputs(3227) <= layer0_outputs(1743);
    layer1_outputs(3228) <= not(layer0_outputs(1775));
    layer1_outputs(3229) <= not((layer0_outputs(1718)) or (layer0_outputs(86)));
    layer1_outputs(3230) <= layer0_outputs(3644);
    layer1_outputs(3231) <= layer0_outputs(96);
    layer1_outputs(3232) <= not(layer0_outputs(5023)) or (layer0_outputs(4928));
    layer1_outputs(3233) <= not((layer0_outputs(1677)) and (layer0_outputs(1315)));
    layer1_outputs(3234) <= '1';
    layer1_outputs(3235) <= not(layer0_outputs(4563)) or (layer0_outputs(287));
    layer1_outputs(3236) <= (layer0_outputs(3104)) xor (layer0_outputs(1731));
    layer1_outputs(3237) <= '0';
    layer1_outputs(3238) <= layer0_outputs(3411);
    layer1_outputs(3239) <= not((layer0_outputs(3330)) or (layer0_outputs(2341)));
    layer1_outputs(3240) <= (layer0_outputs(4576)) xor (layer0_outputs(517));
    layer1_outputs(3241) <= not(layer0_outputs(227));
    layer1_outputs(3242) <= not(layer0_outputs(3740));
    layer1_outputs(3243) <= '1';
    layer1_outputs(3244) <= '1';
    layer1_outputs(3245) <= not(layer0_outputs(3986)) or (layer0_outputs(128));
    layer1_outputs(3246) <= layer0_outputs(2835);
    layer1_outputs(3247) <= (layer0_outputs(3826)) and not (layer0_outputs(2746));
    layer1_outputs(3248) <= not(layer0_outputs(4294));
    layer1_outputs(3249) <= '1';
    layer1_outputs(3250) <= layer0_outputs(2283);
    layer1_outputs(3251) <= '0';
    layer1_outputs(3252) <= not((layer0_outputs(3166)) and (layer0_outputs(200)));
    layer1_outputs(3253) <= not(layer0_outputs(3578));
    layer1_outputs(3254) <= not(layer0_outputs(2149));
    layer1_outputs(3255) <= not(layer0_outputs(3906)) or (layer0_outputs(3200));
    layer1_outputs(3256) <= '0';
    layer1_outputs(3257) <= layer0_outputs(337);
    layer1_outputs(3258) <= not(layer0_outputs(2463));
    layer1_outputs(3259) <= '0';
    layer1_outputs(3260) <= not(layer0_outputs(4562)) or (layer0_outputs(2819));
    layer1_outputs(3261) <= layer0_outputs(2390);
    layer1_outputs(3262) <= (layer0_outputs(1932)) and (layer0_outputs(1820));
    layer1_outputs(3263) <= not(layer0_outputs(4381)) or (layer0_outputs(1907));
    layer1_outputs(3264) <= not(layer0_outputs(1516)) or (layer0_outputs(4953));
    layer1_outputs(3265) <= not(layer0_outputs(1688)) or (layer0_outputs(1886));
    layer1_outputs(3266) <= not((layer0_outputs(1571)) and (layer0_outputs(4723)));
    layer1_outputs(3267) <= '1';
    layer1_outputs(3268) <= (layer0_outputs(1727)) and not (layer0_outputs(674));
    layer1_outputs(3269) <= '1';
    layer1_outputs(3270) <= '1';
    layer1_outputs(3271) <= (layer0_outputs(4476)) and not (layer0_outputs(4733));
    layer1_outputs(3272) <= not(layer0_outputs(4032));
    layer1_outputs(3273) <= (layer0_outputs(1558)) and (layer0_outputs(1178));
    layer1_outputs(3274) <= not((layer0_outputs(173)) or (layer0_outputs(2329)));
    layer1_outputs(3275) <= layer0_outputs(1827);
    layer1_outputs(3276) <= (layer0_outputs(1574)) or (layer0_outputs(3407));
    layer1_outputs(3277) <= not(layer0_outputs(4038));
    layer1_outputs(3278) <= not(layer0_outputs(3527)) or (layer0_outputs(2530));
    layer1_outputs(3279) <= not((layer0_outputs(1641)) or (layer0_outputs(3225)));
    layer1_outputs(3280) <= layer0_outputs(1749);
    layer1_outputs(3281) <= not(layer0_outputs(4936));
    layer1_outputs(3282) <= '0';
    layer1_outputs(3283) <= '1';
    layer1_outputs(3284) <= (layer0_outputs(3629)) and not (layer0_outputs(1128));
    layer1_outputs(3285) <= '1';
    layer1_outputs(3286) <= not(layer0_outputs(954)) or (layer0_outputs(1394));
    layer1_outputs(3287) <= layer0_outputs(4713);
    layer1_outputs(3288) <= layer0_outputs(2967);
    layer1_outputs(3289) <= not(layer0_outputs(3929));
    layer1_outputs(3290) <= layer0_outputs(3750);
    layer1_outputs(3291) <= (layer0_outputs(355)) and not (layer0_outputs(2729));
    layer1_outputs(3292) <= not((layer0_outputs(2717)) or (layer0_outputs(273)));
    layer1_outputs(3293) <= not(layer0_outputs(4607));
    layer1_outputs(3294) <= '0';
    layer1_outputs(3295) <= not(layer0_outputs(4676));
    layer1_outputs(3296) <= '0';
    layer1_outputs(3297) <= '0';
    layer1_outputs(3298) <= layer0_outputs(2972);
    layer1_outputs(3299) <= '1';
    layer1_outputs(3300) <= (layer0_outputs(3490)) and (layer0_outputs(4282));
    layer1_outputs(3301) <= not(layer0_outputs(4800)) or (layer0_outputs(1644));
    layer1_outputs(3302) <= (layer0_outputs(4658)) and not (layer0_outputs(210));
    layer1_outputs(3303) <= (layer0_outputs(2760)) or (layer0_outputs(1131));
    layer1_outputs(3304) <= not((layer0_outputs(1290)) xor (layer0_outputs(3336)));
    layer1_outputs(3305) <= not((layer0_outputs(1679)) or (layer0_outputs(1032)));
    layer1_outputs(3306) <= (layer0_outputs(748)) and not (layer0_outputs(4875));
    layer1_outputs(3307) <= (layer0_outputs(957)) and (layer0_outputs(190));
    layer1_outputs(3308) <= layer0_outputs(3204);
    layer1_outputs(3309) <= layer0_outputs(3320);
    layer1_outputs(3310) <= (layer0_outputs(521)) and not (layer0_outputs(1159));
    layer1_outputs(3311) <= '1';
    layer1_outputs(3312) <= layer0_outputs(3727);
    layer1_outputs(3313) <= not(layer0_outputs(4672)) or (layer0_outputs(1211));
    layer1_outputs(3314) <= not((layer0_outputs(2840)) or (layer0_outputs(645)));
    layer1_outputs(3315) <= not((layer0_outputs(4371)) and (layer0_outputs(142)));
    layer1_outputs(3316) <= (layer0_outputs(2562)) and not (layer0_outputs(4293));
    layer1_outputs(3317) <= not(layer0_outputs(1811));
    layer1_outputs(3318) <= '1';
    layer1_outputs(3319) <= not(layer0_outputs(3274)) or (layer0_outputs(4002));
    layer1_outputs(3320) <= (layer0_outputs(358)) or (layer0_outputs(374));
    layer1_outputs(3321) <= (layer0_outputs(3374)) and not (layer0_outputs(2386));
    layer1_outputs(3322) <= not((layer0_outputs(999)) xor (layer0_outputs(4430)));
    layer1_outputs(3323) <= '0';
    layer1_outputs(3324) <= not(layer0_outputs(4601));
    layer1_outputs(3325) <= '0';
    layer1_outputs(3326) <= (layer0_outputs(3257)) and not (layer0_outputs(5050));
    layer1_outputs(3327) <= '1';
    layer1_outputs(3328) <= not(layer0_outputs(3970)) or (layer0_outputs(2903));
    layer1_outputs(3329) <= (layer0_outputs(772)) and (layer0_outputs(4356));
    layer1_outputs(3330) <= not(layer0_outputs(2616)) or (layer0_outputs(1420));
    layer1_outputs(3331) <= layer0_outputs(1886);
    layer1_outputs(3332) <= not((layer0_outputs(1658)) and (layer0_outputs(82)));
    layer1_outputs(3333) <= not((layer0_outputs(3999)) and (layer0_outputs(3185)));
    layer1_outputs(3334) <= not(layer0_outputs(251));
    layer1_outputs(3335) <= layer0_outputs(346);
    layer1_outputs(3336) <= '0';
    layer1_outputs(3337) <= not(layer0_outputs(3801)) or (layer0_outputs(1595));
    layer1_outputs(3338) <= (layer0_outputs(2754)) and not (layer0_outputs(2549));
    layer1_outputs(3339) <= '1';
    layer1_outputs(3340) <= layer0_outputs(2154);
    layer1_outputs(3341) <= layer0_outputs(261);
    layer1_outputs(3342) <= not(layer0_outputs(5082)) or (layer0_outputs(4482));
    layer1_outputs(3343) <= '1';
    layer1_outputs(3344) <= '0';
    layer1_outputs(3345) <= '1';
    layer1_outputs(3346) <= layer0_outputs(1674);
    layer1_outputs(3347) <= '1';
    layer1_outputs(3348) <= layer0_outputs(2045);
    layer1_outputs(3349) <= not(layer0_outputs(3276)) or (layer0_outputs(4533));
    layer1_outputs(3350) <= (layer0_outputs(1200)) xor (layer0_outputs(2575));
    layer1_outputs(3351) <= not(layer0_outputs(4365)) or (layer0_outputs(4958));
    layer1_outputs(3352) <= not((layer0_outputs(146)) and (layer0_outputs(2340)));
    layer1_outputs(3353) <= not(layer0_outputs(4505));
    layer1_outputs(3354) <= not(layer0_outputs(2850)) or (layer0_outputs(2336));
    layer1_outputs(3355) <= '0';
    layer1_outputs(3356) <= (layer0_outputs(1020)) and not (layer0_outputs(117));
    layer1_outputs(3357) <= (layer0_outputs(1452)) or (layer0_outputs(3688));
    layer1_outputs(3358) <= '0';
    layer1_outputs(3359) <= not(layer0_outputs(3692)) or (layer0_outputs(1859));
    layer1_outputs(3360) <= (layer0_outputs(3524)) and (layer0_outputs(4553));
    layer1_outputs(3361) <= '1';
    layer1_outputs(3362) <= (layer0_outputs(4115)) or (layer0_outputs(1894));
    layer1_outputs(3363) <= '0';
    layer1_outputs(3364) <= not(layer0_outputs(3695));
    layer1_outputs(3365) <= layer0_outputs(2164);
    layer1_outputs(3366) <= '1';
    layer1_outputs(3367) <= not(layer0_outputs(4905)) or (layer0_outputs(1318));
    layer1_outputs(3368) <= (layer0_outputs(4620)) and (layer0_outputs(3078));
    layer1_outputs(3369) <= (layer0_outputs(883)) or (layer0_outputs(32));
    layer1_outputs(3370) <= (layer0_outputs(666)) and not (layer0_outputs(232));
    layer1_outputs(3371) <= '0';
    layer1_outputs(3372) <= not(layer0_outputs(2729));
    layer1_outputs(3373) <= not(layer0_outputs(1764)) or (layer0_outputs(3863));
    layer1_outputs(3374) <= (layer0_outputs(3690)) and (layer0_outputs(3619));
    layer1_outputs(3375) <= '1';
    layer1_outputs(3376) <= '1';
    layer1_outputs(3377) <= (layer0_outputs(3944)) or (layer0_outputs(4571));
    layer1_outputs(3378) <= not((layer0_outputs(791)) xor (layer0_outputs(971)));
    layer1_outputs(3379) <= not(layer0_outputs(465)) or (layer0_outputs(2886));
    layer1_outputs(3380) <= not(layer0_outputs(4227));
    layer1_outputs(3381) <= layer0_outputs(896);
    layer1_outputs(3382) <= layer0_outputs(4327);
    layer1_outputs(3383) <= '1';
    layer1_outputs(3384) <= not((layer0_outputs(1333)) or (layer0_outputs(3752)));
    layer1_outputs(3385) <= not(layer0_outputs(4163)) or (layer0_outputs(799));
    layer1_outputs(3386) <= not(layer0_outputs(4730));
    layer1_outputs(3387) <= layer0_outputs(4052);
    layer1_outputs(3388) <= not((layer0_outputs(3717)) or (layer0_outputs(4442)));
    layer1_outputs(3389) <= '0';
    layer1_outputs(3390) <= (layer0_outputs(1554)) and not (layer0_outputs(983));
    layer1_outputs(3391) <= '1';
    layer1_outputs(3392) <= not((layer0_outputs(253)) or (layer0_outputs(4893)));
    layer1_outputs(3393) <= layer0_outputs(4000);
    layer1_outputs(3394) <= layer0_outputs(2103);
    layer1_outputs(3395) <= layer0_outputs(2955);
    layer1_outputs(3396) <= not((layer0_outputs(1581)) and (layer0_outputs(1627)));
    layer1_outputs(3397) <= '0';
    layer1_outputs(3398) <= '0';
    layer1_outputs(3399) <= not(layer0_outputs(706)) or (layer0_outputs(2975));
    layer1_outputs(3400) <= not(layer0_outputs(1824)) or (layer0_outputs(591));
    layer1_outputs(3401) <= '1';
    layer1_outputs(3402) <= (layer0_outputs(4285)) and not (layer0_outputs(3310));
    layer1_outputs(3403) <= not(layer0_outputs(3753)) or (layer0_outputs(209));
    layer1_outputs(3404) <= layer0_outputs(353);
    layer1_outputs(3405) <= '0';
    layer1_outputs(3406) <= layer0_outputs(768);
    layer1_outputs(3407) <= '1';
    layer1_outputs(3408) <= '1';
    layer1_outputs(3409) <= (layer0_outputs(4582)) and (layer0_outputs(1838));
    layer1_outputs(3410) <= not(layer0_outputs(861));
    layer1_outputs(3411) <= '0';
    layer1_outputs(3412) <= '0';
    layer1_outputs(3413) <= not((layer0_outputs(3389)) and (layer0_outputs(3125)));
    layer1_outputs(3414) <= '1';
    layer1_outputs(3415) <= '1';
    layer1_outputs(3416) <= '1';
    layer1_outputs(3417) <= '1';
    layer1_outputs(3418) <= '0';
    layer1_outputs(3419) <= '0';
    layer1_outputs(3420) <= '1';
    layer1_outputs(3421) <= '0';
    layer1_outputs(3422) <= not(layer0_outputs(3393));
    layer1_outputs(3423) <= '1';
    layer1_outputs(3424) <= not(layer0_outputs(4832));
    layer1_outputs(3425) <= (layer0_outputs(3785)) and (layer0_outputs(4661));
    layer1_outputs(3426) <= (layer0_outputs(2027)) or (layer0_outputs(232));
    layer1_outputs(3427) <= '0';
    layer1_outputs(3428) <= (layer0_outputs(3739)) and not (layer0_outputs(1210));
    layer1_outputs(3429) <= not(layer0_outputs(4022));
    layer1_outputs(3430) <= '1';
    layer1_outputs(3431) <= not(layer0_outputs(78)) or (layer0_outputs(245));
    layer1_outputs(3432) <= '1';
    layer1_outputs(3433) <= not(layer0_outputs(5030));
    layer1_outputs(3434) <= not(layer0_outputs(1636));
    layer1_outputs(3435) <= (layer0_outputs(3007)) and not (layer0_outputs(1318));
    layer1_outputs(3436) <= '1';
    layer1_outputs(3437) <= layer0_outputs(11);
    layer1_outputs(3438) <= not((layer0_outputs(4195)) and (layer0_outputs(2560)));
    layer1_outputs(3439) <= (layer0_outputs(4551)) and not (layer0_outputs(4323));
    layer1_outputs(3440) <= layer0_outputs(4756);
    layer1_outputs(3441) <= '0';
    layer1_outputs(3442) <= (layer0_outputs(1919)) and not (layer0_outputs(4622));
    layer1_outputs(3443) <= not((layer0_outputs(4682)) and (layer0_outputs(4532)));
    layer1_outputs(3444) <= layer0_outputs(2627);
    layer1_outputs(3445) <= not(layer0_outputs(225)) or (layer0_outputs(2605));
    layer1_outputs(3446) <= '0';
    layer1_outputs(3447) <= '1';
    layer1_outputs(3448) <= not((layer0_outputs(4914)) and (layer0_outputs(3371)));
    layer1_outputs(3449) <= layer0_outputs(2609);
    layer1_outputs(3450) <= not((layer0_outputs(4084)) or (layer0_outputs(3151)));
    layer1_outputs(3451) <= '0';
    layer1_outputs(3452) <= '0';
    layer1_outputs(3453) <= layer0_outputs(424);
    layer1_outputs(3454) <= (layer0_outputs(393)) and (layer0_outputs(2647));
    layer1_outputs(3455) <= layer0_outputs(2863);
    layer1_outputs(3456) <= layer0_outputs(4487);
    layer1_outputs(3457) <= not(layer0_outputs(1339));
    layer1_outputs(3458) <= not(layer0_outputs(2738)) or (layer0_outputs(567));
    layer1_outputs(3459) <= layer0_outputs(4095);
    layer1_outputs(3460) <= not((layer0_outputs(2496)) or (layer0_outputs(2515)));
    layer1_outputs(3461) <= (layer0_outputs(903)) or (layer0_outputs(258));
    layer1_outputs(3462) <= (layer0_outputs(409)) or (layer0_outputs(428));
    layer1_outputs(3463) <= '0';
    layer1_outputs(3464) <= not(layer0_outputs(442)) or (layer0_outputs(3561));
    layer1_outputs(3465) <= not(layer0_outputs(4594));
    layer1_outputs(3466) <= not((layer0_outputs(3912)) or (layer0_outputs(2842)));
    layer1_outputs(3467) <= (layer0_outputs(4735)) and (layer0_outputs(1708));
    layer1_outputs(3468) <= '0';
    layer1_outputs(3469) <= '1';
    layer1_outputs(3470) <= not(layer0_outputs(292));
    layer1_outputs(3471) <= not(layer0_outputs(2019)) or (layer0_outputs(4567));
    layer1_outputs(3472) <= not(layer0_outputs(1063));
    layer1_outputs(3473) <= layer0_outputs(4511);
    layer1_outputs(3474) <= (layer0_outputs(4153)) and (layer0_outputs(4093));
    layer1_outputs(3475) <= '1';
    layer1_outputs(3476) <= (layer0_outputs(4710)) and (layer0_outputs(525));
    layer1_outputs(3477) <= not(layer0_outputs(1998)) or (layer0_outputs(3354));
    layer1_outputs(3478) <= not(layer0_outputs(2676));
    layer1_outputs(3479) <= not(layer0_outputs(3340)) or (layer0_outputs(938));
    layer1_outputs(3480) <= (layer0_outputs(4882)) and (layer0_outputs(3407));
    layer1_outputs(3481) <= '1';
    layer1_outputs(3482) <= not((layer0_outputs(2335)) and (layer0_outputs(2863)));
    layer1_outputs(3483) <= '0';
    layer1_outputs(3484) <= not(layer0_outputs(1897));
    layer1_outputs(3485) <= '1';
    layer1_outputs(3486) <= not((layer0_outputs(2111)) or (layer0_outputs(4773)));
    layer1_outputs(3487) <= not((layer0_outputs(3668)) and (layer0_outputs(840)));
    layer1_outputs(3488) <= not(layer0_outputs(252)) or (layer0_outputs(480));
    layer1_outputs(3489) <= not((layer0_outputs(2173)) or (layer0_outputs(377)));
    layer1_outputs(3490) <= not(layer0_outputs(1803));
    layer1_outputs(3491) <= not((layer0_outputs(2780)) or (layer0_outputs(3406)));
    layer1_outputs(3492) <= (layer0_outputs(1863)) and not (layer0_outputs(2864));
    layer1_outputs(3493) <= layer0_outputs(2098);
    layer1_outputs(3494) <= not((layer0_outputs(1570)) or (layer0_outputs(4521)));
    layer1_outputs(3495) <= not(layer0_outputs(3748)) or (layer0_outputs(3379));
    layer1_outputs(3496) <= '0';
    layer1_outputs(3497) <= not(layer0_outputs(1928));
    layer1_outputs(3498) <= '1';
    layer1_outputs(3499) <= not((layer0_outputs(2558)) and (layer0_outputs(4169)));
    layer1_outputs(3500) <= not((layer0_outputs(2786)) or (layer0_outputs(1091)));
    layer1_outputs(3501) <= '0';
    layer1_outputs(3502) <= (layer0_outputs(3808)) and not (layer0_outputs(3711));
    layer1_outputs(3503) <= '1';
    layer1_outputs(3504) <= '0';
    layer1_outputs(3505) <= '1';
    layer1_outputs(3506) <= not(layer0_outputs(3868));
    layer1_outputs(3507) <= not(layer0_outputs(3002)) or (layer0_outputs(2436));
    layer1_outputs(3508) <= '0';
    layer1_outputs(3509) <= not((layer0_outputs(1586)) and (layer0_outputs(808)));
    layer1_outputs(3510) <= (layer0_outputs(1796)) and not (layer0_outputs(2592));
    layer1_outputs(3511) <= not((layer0_outputs(1553)) or (layer0_outputs(2785)));
    layer1_outputs(3512) <= not(layer0_outputs(2282));
    layer1_outputs(3513) <= not(layer0_outputs(752)) or (layer0_outputs(4035));
    layer1_outputs(3514) <= '1';
    layer1_outputs(3515) <= not(layer0_outputs(4333));
    layer1_outputs(3516) <= '1';
    layer1_outputs(3517) <= '0';
    layer1_outputs(3518) <= (layer0_outputs(4626)) and not (layer0_outputs(4435));
    layer1_outputs(3519) <= (layer0_outputs(1405)) and (layer0_outputs(2686));
    layer1_outputs(3520) <= not((layer0_outputs(4880)) or (layer0_outputs(4397)));
    layer1_outputs(3521) <= not(layer0_outputs(3219));
    layer1_outputs(3522) <= (layer0_outputs(1952)) or (layer0_outputs(3683));
    layer1_outputs(3523) <= '1';
    layer1_outputs(3524) <= (layer0_outputs(3664)) and not (layer0_outputs(2012));
    layer1_outputs(3525) <= not(layer0_outputs(847)) or (layer0_outputs(3606));
    layer1_outputs(3526) <= not(layer0_outputs(2468));
    layer1_outputs(3527) <= '0';
    layer1_outputs(3528) <= layer0_outputs(2963);
    layer1_outputs(3529) <= (layer0_outputs(4849)) and (layer0_outputs(1288));
    layer1_outputs(3530) <= (layer0_outputs(3731)) and (layer0_outputs(1424));
    layer1_outputs(3531) <= not(layer0_outputs(2041)) or (layer0_outputs(971));
    layer1_outputs(3532) <= '0';
    layer1_outputs(3533) <= not(layer0_outputs(3188)) or (layer0_outputs(4373));
    layer1_outputs(3534) <= '1';
    layer1_outputs(3535) <= '1';
    layer1_outputs(3536) <= not((layer0_outputs(744)) or (layer0_outputs(3243)));
    layer1_outputs(3537) <= not(layer0_outputs(5040)) or (layer0_outputs(4815));
    layer1_outputs(3538) <= (layer0_outputs(1266)) or (layer0_outputs(3085));
    layer1_outputs(3539) <= (layer0_outputs(634)) xor (layer0_outputs(4621));
    layer1_outputs(3540) <= layer0_outputs(3978);
    layer1_outputs(3541) <= (layer0_outputs(5110)) or (layer0_outputs(2135));
    layer1_outputs(3542) <= not(layer0_outputs(2161)) or (layer0_outputs(2917));
    layer1_outputs(3543) <= not(layer0_outputs(4654));
    layer1_outputs(3544) <= '1';
    layer1_outputs(3545) <= '0';
    layer1_outputs(3546) <= '1';
    layer1_outputs(3547) <= '1';
    layer1_outputs(3548) <= not(layer0_outputs(3992));
    layer1_outputs(3549) <= (layer0_outputs(4724)) and not (layer0_outputs(2434));
    layer1_outputs(3550) <= '0';
    layer1_outputs(3551) <= (layer0_outputs(1048)) xor (layer0_outputs(600));
    layer1_outputs(3552) <= layer0_outputs(1996);
    layer1_outputs(3553) <= not((layer0_outputs(108)) or (layer0_outputs(2651)));
    layer1_outputs(3554) <= '0';
    layer1_outputs(3555) <= not((layer0_outputs(4102)) or (layer0_outputs(4264)));
    layer1_outputs(3556) <= (layer0_outputs(3921)) or (layer0_outputs(3777));
    layer1_outputs(3557) <= (layer0_outputs(3894)) and not (layer0_outputs(916));
    layer1_outputs(3558) <= not((layer0_outputs(2490)) xor (layer0_outputs(94)));
    layer1_outputs(3559) <= '0';
    layer1_outputs(3560) <= '1';
    layer1_outputs(3561) <= not(layer0_outputs(2447)) or (layer0_outputs(3788));
    layer1_outputs(3562) <= (layer0_outputs(4872)) and not (layer0_outputs(2762));
    layer1_outputs(3563) <= (layer0_outputs(803)) and not (layer0_outputs(167));
    layer1_outputs(3564) <= (layer0_outputs(5021)) and not (layer0_outputs(1722));
    layer1_outputs(3565) <= not(layer0_outputs(2144)) or (layer0_outputs(2018));
    layer1_outputs(3566) <= (layer0_outputs(1416)) and not (layer0_outputs(2212));
    layer1_outputs(3567) <= '0';
    layer1_outputs(3568) <= (layer0_outputs(696)) or (layer0_outputs(1380));
    layer1_outputs(3569) <= '0';
    layer1_outputs(3570) <= '1';
    layer1_outputs(3571) <= layer0_outputs(436);
    layer1_outputs(3572) <= not(layer0_outputs(2902)) or (layer0_outputs(979));
    layer1_outputs(3573) <= (layer0_outputs(4417)) and (layer0_outputs(4252));
    layer1_outputs(3574) <= '0';
    layer1_outputs(3575) <= not(layer0_outputs(1448));
    layer1_outputs(3576) <= not(layer0_outputs(3481));
    layer1_outputs(3577) <= not(layer0_outputs(43)) or (layer0_outputs(2351));
    layer1_outputs(3578) <= not((layer0_outputs(4644)) or (layer0_outputs(745)));
    layer1_outputs(3579) <= (layer0_outputs(3264)) or (layer0_outputs(2512));
    layer1_outputs(3580) <= '0';
    layer1_outputs(3581) <= '1';
    layer1_outputs(3582) <= '1';
    layer1_outputs(3583) <= layer0_outputs(498);
    layer1_outputs(3584) <= (layer0_outputs(16)) or (layer0_outputs(1343));
    layer1_outputs(3585) <= not((layer0_outputs(2252)) and (layer0_outputs(2240)));
    layer1_outputs(3586) <= (layer0_outputs(4986)) and not (layer0_outputs(1809));
    layer1_outputs(3587) <= not((layer0_outputs(3256)) or (layer0_outputs(130)));
    layer1_outputs(3588) <= (layer0_outputs(2561)) or (layer0_outputs(270));
    layer1_outputs(3589) <= layer0_outputs(1882);
    layer1_outputs(3590) <= not(layer0_outputs(1810)) or (layer0_outputs(1858));
    layer1_outputs(3591) <= not(layer0_outputs(1488));
    layer1_outputs(3592) <= not((layer0_outputs(2635)) and (layer0_outputs(2735)));
    layer1_outputs(3593) <= layer0_outputs(3435);
    layer1_outputs(3594) <= '1';
    layer1_outputs(3595) <= '1';
    layer1_outputs(3596) <= '1';
    layer1_outputs(3597) <= not(layer0_outputs(2777));
    layer1_outputs(3598) <= layer0_outputs(2922);
    layer1_outputs(3599) <= '1';
    layer1_outputs(3600) <= '1';
    layer1_outputs(3601) <= not(layer0_outputs(702));
    layer1_outputs(3602) <= (layer0_outputs(706)) and not (layer0_outputs(2337));
    layer1_outputs(3603) <= not(layer0_outputs(2559)) or (layer0_outputs(4360));
    layer1_outputs(3604) <= (layer0_outputs(3752)) and not (layer0_outputs(3980));
    layer1_outputs(3605) <= layer0_outputs(146);
    layer1_outputs(3606) <= (layer0_outputs(4352)) and not (layer0_outputs(4));
    layer1_outputs(3607) <= (layer0_outputs(1033)) and (layer0_outputs(619));
    layer1_outputs(3608) <= layer0_outputs(650);
    layer1_outputs(3609) <= not((layer0_outputs(2972)) or (layer0_outputs(2783)));
    layer1_outputs(3610) <= '0';
    layer1_outputs(3611) <= not((layer0_outputs(1870)) or (layer0_outputs(4547)));
    layer1_outputs(3612) <= (layer0_outputs(4747)) and (layer0_outputs(929));
    layer1_outputs(3613) <= '0';
    layer1_outputs(3614) <= not((layer0_outputs(1264)) and (layer0_outputs(2927)));
    layer1_outputs(3615) <= not((layer0_outputs(3367)) and (layer0_outputs(5108)));
    layer1_outputs(3616) <= not((layer0_outputs(2096)) and (layer0_outputs(325)));
    layer1_outputs(3617) <= not(layer0_outputs(1444)) or (layer0_outputs(3357));
    layer1_outputs(3618) <= '1';
    layer1_outputs(3619) <= layer0_outputs(14);
    layer1_outputs(3620) <= not((layer0_outputs(417)) or (layer0_outputs(2743)));
    layer1_outputs(3621) <= not(layer0_outputs(4522)) or (layer0_outputs(1363));
    layer1_outputs(3622) <= (layer0_outputs(403)) and not (layer0_outputs(730));
    layer1_outputs(3623) <= not((layer0_outputs(1917)) and (layer0_outputs(2747)));
    layer1_outputs(3624) <= (layer0_outputs(2793)) or (layer0_outputs(2719));
    layer1_outputs(3625) <= layer0_outputs(3105);
    layer1_outputs(3626) <= not(layer0_outputs(4111));
    layer1_outputs(3627) <= (layer0_outputs(366)) and (layer0_outputs(2060));
    layer1_outputs(3628) <= not((layer0_outputs(2132)) and (layer0_outputs(2057)));
    layer1_outputs(3629) <= '0';
    layer1_outputs(3630) <= '0';
    layer1_outputs(3631) <= '1';
    layer1_outputs(3632) <= (layer0_outputs(3298)) and not (layer0_outputs(3523));
    layer1_outputs(3633) <= layer0_outputs(1802);
    layer1_outputs(3634) <= '1';
    layer1_outputs(3635) <= not(layer0_outputs(2159));
    layer1_outputs(3636) <= layer0_outputs(494);
    layer1_outputs(3637) <= '1';
    layer1_outputs(3638) <= (layer0_outputs(1470)) and (layer0_outputs(3686));
    layer1_outputs(3639) <= '1';
    layer1_outputs(3640) <= not(layer0_outputs(1121));
    layer1_outputs(3641) <= not((layer0_outputs(2109)) and (layer0_outputs(4264)));
    layer1_outputs(3642) <= (layer0_outputs(3260)) and not (layer0_outputs(542));
    layer1_outputs(3643) <= '1';
    layer1_outputs(3644) <= '1';
    layer1_outputs(3645) <= not(layer0_outputs(2495)) or (layer0_outputs(1943));
    layer1_outputs(3646) <= (layer0_outputs(2682)) xor (layer0_outputs(3534));
    layer1_outputs(3647) <= not(layer0_outputs(2948));
    layer1_outputs(3648) <= '0';
    layer1_outputs(3649) <= layer0_outputs(4792);
    layer1_outputs(3650) <= not(layer0_outputs(4474)) or (layer0_outputs(802));
    layer1_outputs(3651) <= (layer0_outputs(3317)) and not (layer0_outputs(1765));
    layer1_outputs(3652) <= not((layer0_outputs(306)) xor (layer0_outputs(1968)));
    layer1_outputs(3653) <= '1';
    layer1_outputs(3654) <= (layer0_outputs(3467)) and not (layer0_outputs(282));
    layer1_outputs(3655) <= not((layer0_outputs(2365)) xor (layer0_outputs(3630)));
    layer1_outputs(3656) <= layer0_outputs(4425);
    layer1_outputs(3657) <= layer0_outputs(963);
    layer1_outputs(3658) <= not((layer0_outputs(749)) or (layer0_outputs(2931)));
    layer1_outputs(3659) <= not((layer0_outputs(4141)) or (layer0_outputs(2069)));
    layer1_outputs(3660) <= (layer0_outputs(4336)) or (layer0_outputs(4082));
    layer1_outputs(3661) <= layer0_outputs(2029);
    layer1_outputs(3662) <= (layer0_outputs(3107)) and not (layer0_outputs(2707));
    layer1_outputs(3663) <= (layer0_outputs(190)) and not (layer0_outputs(3326));
    layer1_outputs(3664) <= layer0_outputs(4375);
    layer1_outputs(3665) <= (layer0_outputs(239)) xor (layer0_outputs(3614));
    layer1_outputs(3666) <= (layer0_outputs(322)) and not (layer0_outputs(2612));
    layer1_outputs(3667) <= (layer0_outputs(3823)) and (layer0_outputs(4491));
    layer1_outputs(3668) <= not(layer0_outputs(4099)) or (layer0_outputs(2241));
    layer1_outputs(3669) <= layer0_outputs(3414);
    layer1_outputs(3670) <= '0';
    layer1_outputs(3671) <= '0';
    layer1_outputs(3672) <= (layer0_outputs(157)) and not (layer0_outputs(3872));
    layer1_outputs(3673) <= not(layer0_outputs(4240));
    layer1_outputs(3674) <= not((layer0_outputs(637)) and (layer0_outputs(3869)));
    layer1_outputs(3675) <= not((layer0_outputs(229)) and (layer0_outputs(2665)));
    layer1_outputs(3676) <= not(layer0_outputs(4072)) or (layer0_outputs(2353));
    layer1_outputs(3677) <= not(layer0_outputs(701)) or (layer0_outputs(3189));
    layer1_outputs(3678) <= not(layer0_outputs(1975));
    layer1_outputs(3679) <= layer0_outputs(2801);
    layer1_outputs(3680) <= '0';
    layer1_outputs(3681) <= (layer0_outputs(969)) and (layer0_outputs(2240));
    layer1_outputs(3682) <= layer0_outputs(1202);
    layer1_outputs(3683) <= '1';
    layer1_outputs(3684) <= (layer0_outputs(3839)) and not (layer0_outputs(1382));
    layer1_outputs(3685) <= '0';
    layer1_outputs(3686) <= not(layer0_outputs(1733)) or (layer0_outputs(4043));
    layer1_outputs(3687) <= (layer0_outputs(2447)) and (layer0_outputs(3066));
    layer1_outputs(3688) <= not((layer0_outputs(669)) and (layer0_outputs(1105)));
    layer1_outputs(3689) <= not((layer0_outputs(2734)) and (layer0_outputs(3094)));
    layer1_outputs(3690) <= not((layer0_outputs(105)) or (layer0_outputs(382)));
    layer1_outputs(3691) <= '1';
    layer1_outputs(3692) <= layer0_outputs(4017);
    layer1_outputs(3693) <= not(layer0_outputs(4346));
    layer1_outputs(3694) <= '1';
    layer1_outputs(3695) <= layer0_outputs(4925);
    layer1_outputs(3696) <= (layer0_outputs(3583)) or (layer0_outputs(4237));
    layer1_outputs(3697) <= not((layer0_outputs(1381)) or (layer0_outputs(2363)));
    layer1_outputs(3698) <= not(layer0_outputs(4065)) or (layer0_outputs(2235));
    layer1_outputs(3699) <= '0';
    layer1_outputs(3700) <= '0';
    layer1_outputs(3701) <= (layer0_outputs(3116)) and not (layer0_outputs(864));
    layer1_outputs(3702) <= (layer0_outputs(1177)) or (layer0_outputs(1424));
    layer1_outputs(3703) <= (layer0_outputs(635)) and not (layer0_outputs(1156));
    layer1_outputs(3704) <= layer0_outputs(2067);
    layer1_outputs(3705) <= '1';
    layer1_outputs(3706) <= not((layer0_outputs(3521)) and (layer0_outputs(2046)));
    layer1_outputs(3707) <= not(layer0_outputs(449)) or (layer0_outputs(871));
    layer1_outputs(3708) <= '0';
    layer1_outputs(3709) <= '0';
    layer1_outputs(3710) <= (layer0_outputs(493)) or (layer0_outputs(1271));
    layer1_outputs(3711) <= (layer0_outputs(2620)) and not (layer0_outputs(1893));
    layer1_outputs(3712) <= not((layer0_outputs(2083)) and (layer0_outputs(159)));
    layer1_outputs(3713) <= (layer0_outputs(3939)) and (layer0_outputs(2007));
    layer1_outputs(3714) <= not((layer0_outputs(1887)) and (layer0_outputs(388)));
    layer1_outputs(3715) <= (layer0_outputs(2994)) and (layer0_outputs(275));
    layer1_outputs(3716) <= '1';
    layer1_outputs(3717) <= '0';
    layer1_outputs(3718) <= (layer0_outputs(1002)) or (layer0_outputs(1475));
    layer1_outputs(3719) <= (layer0_outputs(3983)) and not (layer0_outputs(2181));
    layer1_outputs(3720) <= not(layer0_outputs(4361));
    layer1_outputs(3721) <= layer0_outputs(4594);
    layer1_outputs(3722) <= '0';
    layer1_outputs(3723) <= not(layer0_outputs(1186));
    layer1_outputs(3724) <= not((layer0_outputs(1078)) or (layer0_outputs(3845)));
    layer1_outputs(3725) <= (layer0_outputs(2953)) and not (layer0_outputs(2143));
    layer1_outputs(3726) <= (layer0_outputs(2867)) or (layer0_outputs(1614));
    layer1_outputs(3727) <= (layer0_outputs(1490)) and not (layer0_outputs(4083));
    layer1_outputs(3728) <= '1';
    layer1_outputs(3729) <= not(layer0_outputs(4215)) or (layer0_outputs(2940));
    layer1_outputs(3730) <= not((layer0_outputs(2565)) or (layer0_outputs(4099)));
    layer1_outputs(3731) <= not(layer0_outputs(912));
    layer1_outputs(3732) <= not(layer0_outputs(1703)) or (layer0_outputs(4224));
    layer1_outputs(3733) <= layer0_outputs(1029);
    layer1_outputs(3734) <= '0';
    layer1_outputs(3735) <= (layer0_outputs(741)) and (layer0_outputs(511));
    layer1_outputs(3736) <= not(layer0_outputs(2085));
    layer1_outputs(3737) <= '1';
    layer1_outputs(3738) <= '1';
    layer1_outputs(3739) <= (layer0_outputs(4505)) and not (layer0_outputs(2458));
    layer1_outputs(3740) <= '0';
    layer1_outputs(3741) <= '1';
    layer1_outputs(3742) <= '1';
    layer1_outputs(3743) <= not((layer0_outputs(2507)) or (layer0_outputs(940)));
    layer1_outputs(3744) <= '0';
    layer1_outputs(3745) <= (layer0_outputs(2856)) and not (layer0_outputs(668));
    layer1_outputs(3746) <= layer0_outputs(2258);
    layer1_outputs(3747) <= (layer0_outputs(3341)) and not (layer0_outputs(1432));
    layer1_outputs(3748) <= not(layer0_outputs(699));
    layer1_outputs(3749) <= not(layer0_outputs(5048)) or (layer0_outputs(1086));
    layer1_outputs(3750) <= '0';
    layer1_outputs(3751) <= not(layer0_outputs(3525)) or (layer0_outputs(2470));
    layer1_outputs(3752) <= layer0_outputs(1959);
    layer1_outputs(3753) <= not(layer0_outputs(1093)) or (layer0_outputs(148));
    layer1_outputs(3754) <= not(layer0_outputs(4947)) or (layer0_outputs(1444));
    layer1_outputs(3755) <= not(layer0_outputs(3946));
    layer1_outputs(3756) <= '0';
    layer1_outputs(3757) <= layer0_outputs(1769);
    layer1_outputs(3758) <= '1';
    layer1_outputs(3759) <= '0';
    layer1_outputs(3760) <= not(layer0_outputs(1121)) or (layer0_outputs(4118));
    layer1_outputs(3761) <= '0';
    layer1_outputs(3762) <= (layer0_outputs(1321)) and (layer0_outputs(61));
    layer1_outputs(3763) <= layer0_outputs(3748);
    layer1_outputs(3764) <= (layer0_outputs(2827)) and not (layer0_outputs(205));
    layer1_outputs(3765) <= layer0_outputs(4451);
    layer1_outputs(3766) <= not(layer0_outputs(4885));
    layer1_outputs(3767) <= '0';
    layer1_outputs(3768) <= '1';
    layer1_outputs(3769) <= not((layer0_outputs(4985)) and (layer0_outputs(3547)));
    layer1_outputs(3770) <= not(layer0_outputs(3751)) or (layer0_outputs(3381));
    layer1_outputs(3771) <= '0';
    layer1_outputs(3772) <= layer0_outputs(2221);
    layer1_outputs(3773) <= '0';
    layer1_outputs(3774) <= '0';
    layer1_outputs(3775) <= not(layer0_outputs(1372));
    layer1_outputs(3776) <= (layer0_outputs(2114)) xor (layer0_outputs(1671));
    layer1_outputs(3777) <= layer0_outputs(491);
    layer1_outputs(3778) <= layer0_outputs(5006);
    layer1_outputs(3779) <= (layer0_outputs(782)) and not (layer0_outputs(2779));
    layer1_outputs(3780) <= not(layer0_outputs(1816));
    layer1_outputs(3781) <= not((layer0_outputs(2033)) and (layer0_outputs(4964)));
    layer1_outputs(3782) <= not(layer0_outputs(4009));
    layer1_outputs(3783) <= not(layer0_outputs(1841));
    layer1_outputs(3784) <= not(layer0_outputs(4729)) or (layer0_outputs(4696));
    layer1_outputs(3785) <= not(layer0_outputs(380));
    layer1_outputs(3786) <= not(layer0_outputs(4754));
    layer1_outputs(3787) <= not(layer0_outputs(4874));
    layer1_outputs(3788) <= not(layer0_outputs(2345)) or (layer0_outputs(3861));
    layer1_outputs(3789) <= not(layer0_outputs(3643)) or (layer0_outputs(3015));
    layer1_outputs(3790) <= '0';
    layer1_outputs(3791) <= '1';
    layer1_outputs(3792) <= not(layer0_outputs(3068));
    layer1_outputs(3793) <= (layer0_outputs(838)) and not (layer0_outputs(1222));
    layer1_outputs(3794) <= not(layer0_outputs(2070)) or (layer0_outputs(1090));
    layer1_outputs(3795) <= layer0_outputs(2716);
    layer1_outputs(3796) <= '1';
    layer1_outputs(3797) <= '1';
    layer1_outputs(3798) <= not((layer0_outputs(4192)) or (layer0_outputs(196)));
    layer1_outputs(3799) <= not((layer0_outputs(4466)) and (layer0_outputs(1214)));
    layer1_outputs(3800) <= (layer0_outputs(4050)) and not (layer0_outputs(3882));
    layer1_outputs(3801) <= '0';
    layer1_outputs(3802) <= (layer0_outputs(2263)) and not (layer0_outputs(1370));
    layer1_outputs(3803) <= not((layer0_outputs(1291)) or (layer0_outputs(1803)));
    layer1_outputs(3804) <= not((layer0_outputs(3866)) and (layer0_outputs(3151)));
    layer1_outputs(3805) <= (layer0_outputs(4605)) and (layer0_outputs(461));
    layer1_outputs(3806) <= not(layer0_outputs(2162)) or (layer0_outputs(3284));
    layer1_outputs(3807) <= '0';
    layer1_outputs(3808) <= layer0_outputs(2645);
    layer1_outputs(3809) <= '1';
    layer1_outputs(3810) <= (layer0_outputs(178)) and (layer0_outputs(2822));
    layer1_outputs(3811) <= '1';
    layer1_outputs(3812) <= '0';
    layer1_outputs(3813) <= layer0_outputs(1208);
    layer1_outputs(3814) <= (layer0_outputs(2075)) and not (layer0_outputs(2544));
    layer1_outputs(3815) <= not(layer0_outputs(1741)) or (layer0_outputs(4907));
    layer1_outputs(3816) <= not(layer0_outputs(2223)) or (layer0_outputs(4538));
    layer1_outputs(3817) <= layer0_outputs(961);
    layer1_outputs(3818) <= not(layer0_outputs(980)) or (layer0_outputs(568));
    layer1_outputs(3819) <= not(layer0_outputs(1559));
    layer1_outputs(3820) <= not((layer0_outputs(2412)) and (layer0_outputs(534)));
    layer1_outputs(3821) <= (layer0_outputs(818)) xor (layer0_outputs(1151));
    layer1_outputs(3822) <= (layer0_outputs(314)) and not (layer0_outputs(3113));
    layer1_outputs(3823) <= '1';
    layer1_outputs(3824) <= '0';
    layer1_outputs(3825) <= '1';
    layer1_outputs(3826) <= '1';
    layer1_outputs(3827) <= not(layer0_outputs(4460)) or (layer0_outputs(2526));
    layer1_outputs(3828) <= (layer0_outputs(1537)) or (layer0_outputs(2453));
    layer1_outputs(3829) <= not(layer0_outputs(2783));
    layer1_outputs(3830) <= '0';
    layer1_outputs(3831) <= layer0_outputs(2089);
    layer1_outputs(3832) <= not((layer0_outputs(3400)) and (layer0_outputs(1648)));
    layer1_outputs(3833) <= '1';
    layer1_outputs(3834) <= (layer0_outputs(472)) and (layer0_outputs(1350));
    layer1_outputs(3835) <= not(layer0_outputs(433)) or (layer0_outputs(4508));
    layer1_outputs(3836) <= '1';
    layer1_outputs(3837) <= (layer0_outputs(1941)) and not (layer0_outputs(1889));
    layer1_outputs(3838) <= '1';
    layer1_outputs(3839) <= layer0_outputs(1734);
    layer1_outputs(3840) <= not(layer0_outputs(1510));
    layer1_outputs(3841) <= (layer0_outputs(4053)) and not (layer0_outputs(3394));
    layer1_outputs(3842) <= (layer0_outputs(4851)) and not (layer0_outputs(3229));
    layer1_outputs(3843) <= not(layer0_outputs(3596)) or (layer0_outputs(1551));
    layer1_outputs(3844) <= not((layer0_outputs(3712)) or (layer0_outputs(3575)));
    layer1_outputs(3845) <= '1';
    layer1_outputs(3846) <= (layer0_outputs(4239)) or (layer0_outputs(947));
    layer1_outputs(3847) <= not(layer0_outputs(1364)) or (layer0_outputs(4907));
    layer1_outputs(3848) <= (layer0_outputs(4071)) and not (layer0_outputs(3495));
    layer1_outputs(3849) <= not(layer0_outputs(3128));
    layer1_outputs(3850) <= '1';
    layer1_outputs(3851) <= not(layer0_outputs(5096)) or (layer0_outputs(4436));
    layer1_outputs(3852) <= not((layer0_outputs(1643)) xor (layer0_outputs(3098)));
    layer1_outputs(3853) <= not(layer0_outputs(5057));
    layer1_outputs(3854) <= (layer0_outputs(3530)) or (layer0_outputs(1911));
    layer1_outputs(3855) <= (layer0_outputs(1526)) or (layer0_outputs(640));
    layer1_outputs(3856) <= '1';
    layer1_outputs(3857) <= '1';
    layer1_outputs(3858) <= layer0_outputs(3874);
    layer1_outputs(3859) <= '1';
    layer1_outputs(3860) <= not(layer0_outputs(4470));
    layer1_outputs(3861) <= (layer0_outputs(4961)) and (layer0_outputs(3379));
    layer1_outputs(3862) <= not(layer0_outputs(1861));
    layer1_outputs(3863) <= layer0_outputs(796);
    layer1_outputs(3864) <= (layer0_outputs(129)) and not (layer0_outputs(3515));
    layer1_outputs(3865) <= '0';
    layer1_outputs(3866) <= not((layer0_outputs(3819)) or (layer0_outputs(4529)));
    layer1_outputs(3867) <= '1';
    layer1_outputs(3868) <= '1';
    layer1_outputs(3869) <= not(layer0_outputs(4014)) or (layer0_outputs(3179));
    layer1_outputs(3870) <= (layer0_outputs(4872)) and (layer0_outputs(4347));
    layer1_outputs(3871) <= layer0_outputs(1875);
    layer1_outputs(3872) <= layer0_outputs(886);
    layer1_outputs(3873) <= (layer0_outputs(20)) and not (layer0_outputs(1790));
    layer1_outputs(3874) <= '1';
    layer1_outputs(3875) <= not((layer0_outputs(609)) and (layer0_outputs(4153)));
    layer1_outputs(3876) <= not(layer0_outputs(4057));
    layer1_outputs(3877) <= not((layer0_outputs(3150)) or (layer0_outputs(2962)));
    layer1_outputs(3878) <= '1';
    layer1_outputs(3879) <= (layer0_outputs(1633)) and (layer0_outputs(2739));
    layer1_outputs(3880) <= layer0_outputs(2259);
    layer1_outputs(3881) <= (layer0_outputs(2848)) and not (layer0_outputs(4501));
    layer1_outputs(3882) <= (layer0_outputs(1926)) and not (layer0_outputs(414));
    layer1_outputs(3883) <= layer0_outputs(5040);
    layer1_outputs(3884) <= (layer0_outputs(2417)) xor (layer0_outputs(593));
    layer1_outputs(3885) <= '1';
    layer1_outputs(3886) <= '0';
    layer1_outputs(3887) <= not((layer0_outputs(287)) or (layer0_outputs(4095)));
    layer1_outputs(3888) <= layer0_outputs(249);
    layer1_outputs(3889) <= '0';
    layer1_outputs(3890) <= (layer0_outputs(4918)) and (layer0_outputs(1920));
    layer1_outputs(3891) <= '0';
    layer1_outputs(3892) <= '1';
    layer1_outputs(3893) <= layer0_outputs(4432);
    layer1_outputs(3894) <= not(layer0_outputs(1670)) or (layer0_outputs(858));
    layer1_outputs(3895) <= not((layer0_outputs(3834)) or (layer0_outputs(4002)));
    layer1_outputs(3896) <= (layer0_outputs(528)) and (layer0_outputs(4624));
    layer1_outputs(3897) <= not(layer0_outputs(29)) or (layer0_outputs(4339));
    layer1_outputs(3898) <= '1';
    layer1_outputs(3899) <= layer0_outputs(1653);
    layer1_outputs(3900) <= not((layer0_outputs(627)) xor (layer0_outputs(3577)));
    layer1_outputs(3901) <= '0';
    layer1_outputs(3902) <= not((layer0_outputs(4579)) and (layer0_outputs(2995)));
    layer1_outputs(3903) <= not(layer0_outputs(4646));
    layer1_outputs(3904) <= not(layer0_outputs(2205)) or (layer0_outputs(1329));
    layer1_outputs(3905) <= (layer0_outputs(268)) and not (layer0_outputs(3470));
    layer1_outputs(3906) <= not((layer0_outputs(4004)) or (layer0_outputs(2117)));
    layer1_outputs(3907) <= (layer0_outputs(79)) and (layer0_outputs(1194));
    layer1_outputs(3908) <= '0';
    layer1_outputs(3909) <= (layer0_outputs(2359)) and not (layer0_outputs(2352));
    layer1_outputs(3910) <= (layer0_outputs(2639)) and (layer0_outputs(371));
    layer1_outputs(3911) <= not(layer0_outputs(124));
    layer1_outputs(3912) <= '1';
    layer1_outputs(3913) <= not(layer0_outputs(3816)) or (layer0_outputs(4537));
    layer1_outputs(3914) <= layer0_outputs(821);
    layer1_outputs(3915) <= (layer0_outputs(4037)) and not (layer0_outputs(719));
    layer1_outputs(3916) <= '1';
    layer1_outputs(3917) <= not((layer0_outputs(1116)) or (layer0_outputs(2569)));
    layer1_outputs(3918) <= '1';
    layer1_outputs(3919) <= not(layer0_outputs(405));
    layer1_outputs(3920) <= not(layer0_outputs(1865)) or (layer0_outputs(3175));
    layer1_outputs(3921) <= (layer0_outputs(4587)) and (layer0_outputs(4352));
    layer1_outputs(3922) <= layer0_outputs(2813);
    layer1_outputs(3923) <= not((layer0_outputs(4800)) and (layer0_outputs(2880)));
    layer1_outputs(3924) <= not((layer0_outputs(301)) or (layer0_outputs(291)));
    layer1_outputs(3925) <= '0';
    layer1_outputs(3926) <= not(layer0_outputs(1385));
    layer1_outputs(3927) <= (layer0_outputs(766)) and not (layer0_outputs(3102));
    layer1_outputs(3928) <= (layer0_outputs(674)) and not (layer0_outputs(3152));
    layer1_outputs(3929) <= (layer0_outputs(90)) and (layer0_outputs(3975));
    layer1_outputs(3930) <= not(layer0_outputs(1562)) or (layer0_outputs(3551));
    layer1_outputs(3931) <= layer0_outputs(5);
    layer1_outputs(3932) <= not(layer0_outputs(2432));
    layer1_outputs(3933) <= '0';
    layer1_outputs(3934) <= '0';
    layer1_outputs(3935) <= (layer0_outputs(2231)) and not (layer0_outputs(813));
    layer1_outputs(3936) <= not(layer0_outputs(2832));
    layer1_outputs(3937) <= not((layer0_outputs(2537)) xor (layer0_outputs(855)));
    layer1_outputs(3938) <= (layer0_outputs(283)) or (layer0_outputs(2409));
    layer1_outputs(3939) <= '1';
    layer1_outputs(3940) <= layer0_outputs(3907);
    layer1_outputs(3941) <= '0';
    layer1_outputs(3942) <= not(layer0_outputs(649)) or (layer0_outputs(384));
    layer1_outputs(3943) <= (layer0_outputs(4527)) and not (layer0_outputs(1428));
    layer1_outputs(3944) <= layer0_outputs(2378);
    layer1_outputs(3945) <= (layer0_outputs(1354)) or (layer0_outputs(3174));
    layer1_outputs(3946) <= not(layer0_outputs(783));
    layer1_outputs(3947) <= '0';
    layer1_outputs(3948) <= (layer0_outputs(4051)) or (layer0_outputs(1431));
    layer1_outputs(3949) <= not(layer0_outputs(3173));
    layer1_outputs(3950) <= not(layer0_outputs(2821)) or (layer0_outputs(1090));
    layer1_outputs(3951) <= not(layer0_outputs(2837)) or (layer0_outputs(4534));
    layer1_outputs(3952) <= layer0_outputs(1168);
    layer1_outputs(3953) <= '0';
    layer1_outputs(3954) <= (layer0_outputs(4674)) and not (layer0_outputs(860));
    layer1_outputs(3955) <= (layer0_outputs(3019)) and not (layer0_outputs(4128));
    layer1_outputs(3956) <= not(layer0_outputs(5087));
    layer1_outputs(3957) <= not((layer0_outputs(928)) and (layer0_outputs(1390)));
    layer1_outputs(3958) <= (layer0_outputs(19)) and not (layer0_outputs(2605));
    layer1_outputs(3959) <= not(layer0_outputs(4254));
    layer1_outputs(3960) <= (layer0_outputs(4814)) and (layer0_outputs(4764));
    layer1_outputs(3961) <= not((layer0_outputs(938)) or (layer0_outputs(1314)));
    layer1_outputs(3962) <= (layer0_outputs(4936)) and (layer0_outputs(2160));
    layer1_outputs(3963) <= (layer0_outputs(4562)) and not (layer0_outputs(2974));
    layer1_outputs(3964) <= '0';
    layer1_outputs(3965) <= not(layer0_outputs(1801)) or (layer0_outputs(4758));
    layer1_outputs(3966) <= not((layer0_outputs(2491)) or (layer0_outputs(2457)));
    layer1_outputs(3967) <= (layer0_outputs(4945)) or (layer0_outputs(2935));
    layer1_outputs(3968) <= '1';
    layer1_outputs(3969) <= '1';
    layer1_outputs(3970) <= '0';
    layer1_outputs(3971) <= (layer0_outputs(3569)) and not (layer0_outputs(323));
    layer1_outputs(3972) <= not(layer0_outputs(824)) or (layer0_outputs(3925));
    layer1_outputs(3973) <= not(layer0_outputs(531)) or (layer0_outputs(686));
    layer1_outputs(3974) <= not((layer0_outputs(4856)) xor (layer0_outputs(230)));
    layer1_outputs(3975) <= '0';
    layer1_outputs(3976) <= '0';
    layer1_outputs(3977) <= not(layer0_outputs(2789)) or (layer0_outputs(2141));
    layer1_outputs(3978) <= not((layer0_outputs(4648)) or (layer0_outputs(5118)));
    layer1_outputs(3979) <= '1';
    layer1_outputs(3980) <= (layer0_outputs(5094)) or (layer0_outputs(2081));
    layer1_outputs(3981) <= '1';
    layer1_outputs(3982) <= (layer0_outputs(1377)) and not (layer0_outputs(2999));
    layer1_outputs(3983) <= layer0_outputs(1105);
    layer1_outputs(3984) <= not(layer0_outputs(2083)) or (layer0_outputs(1625));
    layer1_outputs(3985) <= layer0_outputs(1667);
    layer1_outputs(3986) <= '0';
    layer1_outputs(3987) <= layer0_outputs(4709);
    layer1_outputs(3988) <= (layer0_outputs(2796)) and not (layer0_outputs(4286));
    layer1_outputs(3989) <= '1';
    layer1_outputs(3990) <= '0';
    layer1_outputs(3991) <= not((layer0_outputs(4260)) and (layer0_outputs(4309)));
    layer1_outputs(3992) <= (layer0_outputs(4385)) and not (layer0_outputs(1755));
    layer1_outputs(3993) <= not(layer0_outputs(2621));
    layer1_outputs(3994) <= '1';
    layer1_outputs(3995) <= (layer0_outputs(2677)) and not (layer0_outputs(1543));
    layer1_outputs(3996) <= not(layer0_outputs(692)) or (layer0_outputs(1827));
    layer1_outputs(3997) <= (layer0_outputs(5037)) or (layer0_outputs(4634));
    layer1_outputs(3998) <= not((layer0_outputs(2894)) and (layer0_outputs(805)));
    layer1_outputs(3999) <= not(layer0_outputs(3000)) or (layer0_outputs(1466));
    layer1_outputs(4000) <= layer0_outputs(4128);
    layer1_outputs(4001) <= (layer0_outputs(603)) and (layer0_outputs(10));
    layer1_outputs(4002) <= '1';
    layer1_outputs(4003) <= (layer0_outputs(3781)) and (layer0_outputs(2360));
    layer1_outputs(4004) <= '1';
    layer1_outputs(4005) <= not(layer0_outputs(732)) or (layer0_outputs(2147));
    layer1_outputs(4006) <= not(layer0_outputs(341)) or (layer0_outputs(1610));
    layer1_outputs(4007) <= (layer0_outputs(3787)) or (layer0_outputs(859));
    layer1_outputs(4008) <= not(layer0_outputs(5021));
    layer1_outputs(4009) <= not(layer0_outputs(303)) or (layer0_outputs(3562));
    layer1_outputs(4010) <= (layer0_outputs(4485)) and (layer0_outputs(3302));
    layer1_outputs(4011) <= not((layer0_outputs(3847)) and (layer0_outputs(4605)));
    layer1_outputs(4012) <= (layer0_outputs(1902)) or (layer0_outputs(1331));
    layer1_outputs(4013) <= layer0_outputs(576);
    layer1_outputs(4014) <= not(layer0_outputs(533));
    layer1_outputs(4015) <= not(layer0_outputs(4625));
    layer1_outputs(4016) <= not(layer0_outputs(617)) or (layer0_outputs(3559));
    layer1_outputs(4017) <= not(layer0_outputs(4233));
    layer1_outputs(4018) <= not((layer0_outputs(1269)) or (layer0_outputs(3131)));
    layer1_outputs(4019) <= '1';
    layer1_outputs(4020) <= '0';
    layer1_outputs(4021) <= (layer0_outputs(4581)) and not (layer0_outputs(3404));
    layer1_outputs(4022) <= layer0_outputs(760);
    layer1_outputs(4023) <= not(layer0_outputs(413)) or (layer0_outputs(1469));
    layer1_outputs(4024) <= (layer0_outputs(2854)) or (layer0_outputs(3441));
    layer1_outputs(4025) <= '1';
    layer1_outputs(4026) <= '0';
    layer1_outputs(4027) <= '1';
    layer1_outputs(4028) <= not((layer0_outputs(4214)) or (layer0_outputs(3665)));
    layer1_outputs(4029) <= (layer0_outputs(913)) and not (layer0_outputs(4094));
    layer1_outputs(4030) <= layer0_outputs(3567);
    layer1_outputs(4031) <= '1';
    layer1_outputs(4032) <= '0';
    layer1_outputs(4033) <= (layer0_outputs(746)) and not (layer0_outputs(4642));
    layer1_outputs(4034) <= layer0_outputs(1402);
    layer1_outputs(4035) <= not((layer0_outputs(1036)) and (layer0_outputs(3656)));
    layer1_outputs(4036) <= not(layer0_outputs(4996));
    layer1_outputs(4037) <= (layer0_outputs(889)) and not (layer0_outputs(1270));
    layer1_outputs(4038) <= '1';
    layer1_outputs(4039) <= not((layer0_outputs(4954)) or (layer0_outputs(2314)));
    layer1_outputs(4040) <= not((layer0_outputs(4421)) or (layer0_outputs(5117)));
    layer1_outputs(4041) <= '1';
    layer1_outputs(4042) <= layer0_outputs(690);
    layer1_outputs(4043) <= not(layer0_outputs(1732)) or (layer0_outputs(2739));
    layer1_outputs(4044) <= (layer0_outputs(1776)) or (layer0_outputs(135));
    layer1_outputs(4045) <= layer0_outputs(736);
    layer1_outputs(4046) <= '0';
    layer1_outputs(4047) <= not(layer0_outputs(2902)) or (layer0_outputs(62));
    layer1_outputs(4048) <= (layer0_outputs(4284)) and not (layer0_outputs(2113));
    layer1_outputs(4049) <= layer0_outputs(1117);
    layer1_outputs(4050) <= '1';
    layer1_outputs(4051) <= not(layer0_outputs(3455));
    layer1_outputs(4052) <= layer0_outputs(4323);
    layer1_outputs(4053) <= (layer0_outputs(2467)) and not (layer0_outputs(392));
    layer1_outputs(4054) <= not((layer0_outputs(1974)) or (layer0_outputs(2246)));
    layer1_outputs(4055) <= layer0_outputs(1140);
    layer1_outputs(4056) <= '0';
    layer1_outputs(4057) <= layer0_outputs(312);
    layer1_outputs(4058) <= '0';
    layer1_outputs(4059) <= '1';
    layer1_outputs(4060) <= not(layer0_outputs(4923));
    layer1_outputs(4061) <= not((layer0_outputs(230)) and (layer0_outputs(1787)));
    layer1_outputs(4062) <= layer0_outputs(2218);
    layer1_outputs(4063) <= not(layer0_outputs(4143));
    layer1_outputs(4064) <= not(layer0_outputs(2552)) or (layer0_outputs(3471));
    layer1_outputs(4065) <= not((layer0_outputs(4363)) and (layer0_outputs(2176)));
    layer1_outputs(4066) <= (layer0_outputs(542)) and not (layer0_outputs(1690));
    layer1_outputs(4067) <= '0';
    layer1_outputs(4068) <= '1';
    layer1_outputs(4069) <= '0';
    layer1_outputs(4070) <= (layer0_outputs(2403)) and not (layer0_outputs(112));
    layer1_outputs(4071) <= '1';
    layer1_outputs(4072) <= (layer0_outputs(4246)) and not (layer0_outputs(1340));
    layer1_outputs(4073) <= '1';
    layer1_outputs(4074) <= not(layer0_outputs(436));
    layer1_outputs(4075) <= layer0_outputs(856);
    layer1_outputs(4076) <= not(layer0_outputs(2445)) or (layer0_outputs(655));
    layer1_outputs(4077) <= not((layer0_outputs(2724)) or (layer0_outputs(1728)));
    layer1_outputs(4078) <= '1';
    layer1_outputs(4079) <= (layer0_outputs(104)) and not (layer0_outputs(1672));
    layer1_outputs(4080) <= not(layer0_outputs(4372));
    layer1_outputs(4081) <= '1';
    layer1_outputs(4082) <= '1';
    layer1_outputs(4083) <= not(layer0_outputs(2613)) or (layer0_outputs(1775));
    layer1_outputs(4084) <= not((layer0_outputs(3830)) or (layer0_outputs(2685)));
    layer1_outputs(4085) <= not(layer0_outputs(1949)) or (layer0_outputs(1961));
    layer1_outputs(4086) <= not((layer0_outputs(87)) and (layer0_outputs(3313)));
    layer1_outputs(4087) <= '1';
    layer1_outputs(4088) <= not(layer0_outputs(3634));
    layer1_outputs(4089) <= not((layer0_outputs(822)) and (layer0_outputs(3735)));
    layer1_outputs(4090) <= '0';
    layer1_outputs(4091) <= layer0_outputs(3328);
    layer1_outputs(4092) <= '0';
    layer1_outputs(4093) <= layer0_outputs(398);
    layer1_outputs(4094) <= not(layer0_outputs(801)) or (layer0_outputs(3362));
    layer1_outputs(4095) <= layer0_outputs(1127);
    layer1_outputs(4096) <= not((layer0_outputs(814)) or (layer0_outputs(1520)));
    layer1_outputs(4097) <= not(layer0_outputs(4642)) or (layer0_outputs(4528));
    layer1_outputs(4098) <= '0';
    layer1_outputs(4099) <= (layer0_outputs(3522)) xor (layer0_outputs(1515));
    layer1_outputs(4100) <= (layer0_outputs(3928)) and not (layer0_outputs(1556));
    layer1_outputs(4101) <= layer0_outputs(4335);
    layer1_outputs(4102) <= not(layer0_outputs(116));
    layer1_outputs(4103) <= not((layer0_outputs(4673)) or (layer0_outputs(5100)));
    layer1_outputs(4104) <= '1';
    layer1_outputs(4105) <= not(layer0_outputs(3050)) or (layer0_outputs(3294));
    layer1_outputs(4106) <= not((layer0_outputs(2301)) or (layer0_outputs(1427)));
    layer1_outputs(4107) <= not((layer0_outputs(860)) xor (layer0_outputs(4822)));
    layer1_outputs(4108) <= '1';
    layer1_outputs(4109) <= not(layer0_outputs(2899));
    layer1_outputs(4110) <= (layer0_outputs(2046)) and not (layer0_outputs(80));
    layer1_outputs(4111) <= not((layer0_outputs(2025)) and (layer0_outputs(4995)));
    layer1_outputs(4112) <= not(layer0_outputs(587)) or (layer0_outputs(177));
    layer1_outputs(4113) <= not(layer0_outputs(2095)) or (layer0_outputs(2176));
    layer1_outputs(4114) <= layer0_outputs(839);
    layer1_outputs(4115) <= (layer0_outputs(1175)) or (layer0_outputs(4864));
    layer1_outputs(4116) <= '1';
    layer1_outputs(4117) <= not(layer0_outputs(2343));
    layer1_outputs(4118) <= '0';
    layer1_outputs(4119) <= '0';
    layer1_outputs(4120) <= not((layer0_outputs(165)) and (layer0_outputs(3479)));
    layer1_outputs(4121) <= '0';
    layer1_outputs(4122) <= (layer0_outputs(4431)) or (layer0_outputs(4234));
    layer1_outputs(4123) <= layer0_outputs(3157);
    layer1_outputs(4124) <= '1';
    layer1_outputs(4125) <= not((layer0_outputs(2021)) and (layer0_outputs(771)));
    layer1_outputs(4126) <= '1';
    layer1_outputs(4127) <= (layer0_outputs(925)) and (layer0_outputs(1884));
    layer1_outputs(4128) <= not(layer0_outputs(1749));
    layer1_outputs(4129) <= (layer0_outputs(113)) or (layer0_outputs(804));
    layer1_outputs(4130) <= not(layer0_outputs(1592)) or (layer0_outputs(1227));
    layer1_outputs(4131) <= not((layer0_outputs(4551)) or (layer0_outputs(3742)));
    layer1_outputs(4132) <= (layer0_outputs(47)) and not (layer0_outputs(589));
    layer1_outputs(4133) <= '1';
    layer1_outputs(4134) <= not(layer0_outputs(2413)) or (layer0_outputs(1935));
    layer1_outputs(4135) <= not((layer0_outputs(1495)) or (layer0_outputs(4580)));
    layer1_outputs(4136) <= (layer0_outputs(481)) and not (layer0_outputs(2393));
    layer1_outputs(4137) <= layer0_outputs(3375);
    layer1_outputs(4138) <= '1';
    layer1_outputs(4139) <= not(layer0_outputs(2725)) or (layer0_outputs(2094));
    layer1_outputs(4140) <= not((layer0_outputs(3725)) and (layer0_outputs(241)));
    layer1_outputs(4141) <= not(layer0_outputs(2372));
    layer1_outputs(4142) <= layer0_outputs(4632);
    layer1_outputs(4143) <= '1';
    layer1_outputs(4144) <= not((layer0_outputs(1030)) and (layer0_outputs(708)));
    layer1_outputs(4145) <= '1';
    layer1_outputs(4146) <= layer0_outputs(4892);
    layer1_outputs(4147) <= '0';
    layer1_outputs(4148) <= '0';
    layer1_outputs(4149) <= not((layer0_outputs(3542)) and (layer0_outputs(3277)));
    layer1_outputs(4150) <= not(layer0_outputs(2660));
    layer1_outputs(4151) <= layer0_outputs(2324);
    layer1_outputs(4152) <= '1';
    layer1_outputs(4153) <= (layer0_outputs(4565)) or (layer0_outputs(1306));
    layer1_outputs(4154) <= not((layer0_outputs(4707)) or (layer0_outputs(2008)));
    layer1_outputs(4155) <= not(layer0_outputs(1198)) or (layer0_outputs(842));
    layer1_outputs(4156) <= '0';
    layer1_outputs(4157) <= (layer0_outputs(2507)) and (layer0_outputs(4669));
    layer1_outputs(4158) <= not((layer0_outputs(4228)) or (layer0_outputs(2751)));
    layer1_outputs(4159) <= layer0_outputs(1557);
    layer1_outputs(4160) <= not(layer0_outputs(4061)) or (layer0_outputs(351));
    layer1_outputs(4161) <= '0';
    layer1_outputs(4162) <= not((layer0_outputs(2214)) or (layer0_outputs(437)));
    layer1_outputs(4163) <= (layer0_outputs(4687)) and (layer0_outputs(2660));
    layer1_outputs(4164) <= layer0_outputs(5017);
    layer1_outputs(4165) <= (layer0_outputs(1218)) and (layer0_outputs(1274));
    layer1_outputs(4166) <= layer0_outputs(4342);
    layer1_outputs(4167) <= not(layer0_outputs(778)) or (layer0_outputs(258));
    layer1_outputs(4168) <= (layer0_outputs(4757)) and not (layer0_outputs(4332));
    layer1_outputs(4169) <= layer0_outputs(2832);
    layer1_outputs(4170) <= not(layer0_outputs(1064));
    layer1_outputs(4171) <= (layer0_outputs(1707)) and (layer0_outputs(340));
    layer1_outputs(4172) <= '1';
    layer1_outputs(4173) <= '0';
    layer1_outputs(4174) <= not(layer0_outputs(3792)) or (layer0_outputs(4304));
    layer1_outputs(4175) <= not(layer0_outputs(1338));
    layer1_outputs(4176) <= (layer0_outputs(1457)) and not (layer0_outputs(3931));
    layer1_outputs(4177) <= (layer0_outputs(4301)) and (layer0_outputs(1613));
    layer1_outputs(4178) <= not((layer0_outputs(1439)) and (layer0_outputs(3521)));
    layer1_outputs(4179) <= not(layer0_outputs(3802));
    layer1_outputs(4180) <= not((layer0_outputs(2844)) and (layer0_outputs(4561)));
    layer1_outputs(4181) <= layer0_outputs(1353);
    layer1_outputs(4182) <= '1';
    layer1_outputs(4183) <= not(layer0_outputs(3022)) or (layer0_outputs(599));
    layer1_outputs(4184) <= '1';
    layer1_outputs(4185) <= layer0_outputs(4704);
    layer1_outputs(4186) <= not(layer0_outputs(1589));
    layer1_outputs(4187) <= '0';
    layer1_outputs(4188) <= not((layer0_outputs(4306)) and (layer0_outputs(2458)));
    layer1_outputs(4189) <= '0';
    layer1_outputs(4190) <= layer0_outputs(2421);
    layer1_outputs(4191) <= '0';
    layer1_outputs(4192) <= not((layer0_outputs(4392)) or (layer0_outputs(737)));
    layer1_outputs(4193) <= not(layer0_outputs(1866));
    layer1_outputs(4194) <= not(layer0_outputs(1545)) or (layer0_outputs(872));
    layer1_outputs(4195) <= (layer0_outputs(3816)) and not (layer0_outputs(1555));
    layer1_outputs(4196) <= not(layer0_outputs(3700));
    layer1_outputs(4197) <= not(layer0_outputs(3185)) or (layer0_outputs(3808));
    layer1_outputs(4198) <= (layer0_outputs(1261)) and not (layer0_outputs(4530));
    layer1_outputs(4199) <= '0';
    layer1_outputs(4200) <= '1';
    layer1_outputs(4201) <= '0';
    layer1_outputs(4202) <= (layer0_outputs(4074)) and (layer0_outputs(4356));
    layer1_outputs(4203) <= layer0_outputs(2607);
    layer1_outputs(4204) <= not(layer0_outputs(3602)) or (layer0_outputs(4911));
    layer1_outputs(4205) <= (layer0_outputs(4917)) or (layer0_outputs(4749));
    layer1_outputs(4206) <= not((layer0_outputs(3600)) and (layer0_outputs(1366)));
    layer1_outputs(4207) <= not((layer0_outputs(3176)) and (layer0_outputs(3769)));
    layer1_outputs(4208) <= (layer0_outputs(1239)) and not (layer0_outputs(752));
    layer1_outputs(4209) <= '0';
    layer1_outputs(4210) <= not(layer0_outputs(4853)) or (layer0_outputs(1008));
    layer1_outputs(4211) <= '0';
    layer1_outputs(4212) <= not((layer0_outputs(1166)) and (layer0_outputs(1122)));
    layer1_outputs(4213) <= '1';
    layer1_outputs(4214) <= not(layer0_outputs(904));
    layer1_outputs(4215) <= '0';
    layer1_outputs(4216) <= layer0_outputs(2020);
    layer1_outputs(4217) <= not((layer0_outputs(1106)) or (layer0_outputs(4025)));
    layer1_outputs(4218) <= '0';
    layer1_outputs(4219) <= '0';
    layer1_outputs(4220) <= not((layer0_outputs(1071)) xor (layer0_outputs(884)));
    layer1_outputs(4221) <= '0';
    layer1_outputs(4222) <= '0';
    layer1_outputs(4223) <= not(layer0_outputs(1395));
    layer1_outputs(4224) <= not(layer0_outputs(131));
    layer1_outputs(4225) <= not(layer0_outputs(4876)) or (layer0_outputs(927));
    layer1_outputs(4226) <= '1';
    layer1_outputs(4227) <= (layer0_outputs(1487)) and not (layer0_outputs(1893));
    layer1_outputs(4228) <= not((layer0_outputs(3974)) and (layer0_outputs(185)));
    layer1_outputs(4229) <= '1';
    layer1_outputs(4230) <= not(layer0_outputs(2406)) or (layer0_outputs(2499));
    layer1_outputs(4231) <= not(layer0_outputs(4123));
    layer1_outputs(4232) <= not(layer0_outputs(1800)) or (layer0_outputs(3979));
    layer1_outputs(4233) <= '0';
    layer1_outputs(4234) <= not(layer0_outputs(1142));
    layer1_outputs(4235) <= not((layer0_outputs(4459)) and (layer0_outputs(194)));
    layer1_outputs(4236) <= not(layer0_outputs(3875)) or (layer0_outputs(2034));
    layer1_outputs(4237) <= (layer0_outputs(3537)) or (layer0_outputs(1142));
    layer1_outputs(4238) <= (layer0_outputs(689)) and (layer0_outputs(387));
    layer1_outputs(4239) <= not(layer0_outputs(896));
    layer1_outputs(4240) <= (layer0_outputs(1760)) or (layer0_outputs(902));
    layer1_outputs(4241) <= '0';
    layer1_outputs(4242) <= not(layer0_outputs(4805)) or (layer0_outputs(3615));
    layer1_outputs(4243) <= not(layer0_outputs(4794)) or (layer0_outputs(1986));
    layer1_outputs(4244) <= not(layer0_outputs(791));
    layer1_outputs(4245) <= not(layer0_outputs(1253)) or (layer0_outputs(300));
    layer1_outputs(4246) <= not((layer0_outputs(3968)) and (layer0_outputs(1572)));
    layer1_outputs(4247) <= (layer0_outputs(1087)) or (layer0_outputs(3353));
    layer1_outputs(4248) <= layer0_outputs(650);
    layer1_outputs(4249) <= not(layer0_outputs(45));
    layer1_outputs(4250) <= '0';
    layer1_outputs(4251) <= layer0_outputs(2294);
    layer1_outputs(4252) <= '0';
    layer1_outputs(4253) <= '1';
    layer1_outputs(4254) <= not(layer0_outputs(1882));
    layer1_outputs(4255) <= not(layer0_outputs(1781)) or (layer0_outputs(179));
    layer1_outputs(4256) <= not((layer0_outputs(2982)) and (layer0_outputs(2043)));
    layer1_outputs(4257) <= layer0_outputs(1345);
    layer1_outputs(4258) <= (layer0_outputs(4826)) and not (layer0_outputs(2866));
    layer1_outputs(4259) <= not(layer0_outputs(2669));
    layer1_outputs(4260) <= not(layer0_outputs(1073)) or (layer0_outputs(2385));
    layer1_outputs(4261) <= not(layer0_outputs(1911)) or (layer0_outputs(71));
    layer1_outputs(4262) <= (layer0_outputs(4229)) and not (layer0_outputs(2028));
    layer1_outputs(4263) <= not(layer0_outputs(3231)) or (layer0_outputs(1753));
    layer1_outputs(4264) <= not((layer0_outputs(1740)) and (layer0_outputs(4789)));
    layer1_outputs(4265) <= layer0_outputs(3241);
    layer1_outputs(4266) <= not(layer0_outputs(438)) or (layer0_outputs(3145));
    layer1_outputs(4267) <= not(layer0_outputs(4256)) or (layer0_outputs(917));
    layer1_outputs(4268) <= (layer0_outputs(775)) or (layer0_outputs(910));
    layer1_outputs(4269) <= (layer0_outputs(330)) and not (layer0_outputs(326));
    layer1_outputs(4270) <= '0';
    layer1_outputs(4271) <= (layer0_outputs(1343)) and (layer0_outputs(3622));
    layer1_outputs(4272) <= (layer0_outputs(396)) and not (layer0_outputs(3795));
    layer1_outputs(4273) <= layer0_outputs(1419);
    layer1_outputs(4274) <= (layer0_outputs(4943)) or (layer0_outputs(2628));
    layer1_outputs(4275) <= '1';
    layer1_outputs(4276) <= '0';
    layer1_outputs(4277) <= not(layer0_outputs(933));
    layer1_outputs(4278) <= not(layer0_outputs(4020)) or (layer0_outputs(3703));
    layer1_outputs(4279) <= layer0_outputs(1003);
    layer1_outputs(4280) <= '0';
    layer1_outputs(4281) <= not(layer0_outputs(4516));
    layer1_outputs(4282) <= not((layer0_outputs(2885)) and (layer0_outputs(808)));
    layer1_outputs(4283) <= layer0_outputs(4088);
    layer1_outputs(4284) <= (layer0_outputs(1560)) and (layer0_outputs(1980));
    layer1_outputs(4285) <= '1';
    layer1_outputs(4286) <= '1';
    layer1_outputs(4287) <= (layer0_outputs(3532)) and not (layer0_outputs(4512));
    layer1_outputs(4288) <= not((layer0_outputs(4957)) and (layer0_outputs(1941)));
    layer1_outputs(4289) <= (layer0_outputs(4345)) or (layer0_outputs(2900));
    layer1_outputs(4290) <= '1';
    layer1_outputs(4291) <= (layer0_outputs(1901)) xor (layer0_outputs(3786));
    layer1_outputs(4292) <= not(layer0_outputs(3841));
    layer1_outputs(4293) <= layer0_outputs(2429);
    layer1_outputs(4294) <= not(layer0_outputs(1596));
    layer1_outputs(4295) <= (layer0_outputs(3388)) or (layer0_outputs(2445));
    layer1_outputs(4296) <= not(layer0_outputs(3670));
    layer1_outputs(4297) <= layer0_outputs(4319);
    layer1_outputs(4298) <= layer0_outputs(3932);
    layer1_outputs(4299) <= not((layer0_outputs(486)) xor (layer0_outputs(3989)));
    layer1_outputs(4300) <= not(layer0_outputs(2708)) or (layer0_outputs(389));
    layer1_outputs(4301) <= not((layer0_outputs(2062)) or (layer0_outputs(3372)));
    layer1_outputs(4302) <= '0';
    layer1_outputs(4303) <= (layer0_outputs(2243)) and not (layer0_outputs(928));
    layer1_outputs(4304) <= layer0_outputs(3335);
    layer1_outputs(4305) <= not(layer0_outputs(1966)) or (layer0_outputs(2951));
    layer1_outputs(4306) <= '0';
    layer1_outputs(4307) <= not(layer0_outputs(130));
    layer1_outputs(4308) <= (layer0_outputs(2545)) or (layer0_outputs(1017));
    layer1_outputs(4309) <= (layer0_outputs(3191)) and (layer0_outputs(3331));
    layer1_outputs(4310) <= not(layer0_outputs(4788));
    layer1_outputs(4311) <= not(layer0_outputs(1572)) or (layer0_outputs(3964));
    layer1_outputs(4312) <= '1';
    layer1_outputs(4313) <= (layer0_outputs(4772)) or (layer0_outputs(3891));
    layer1_outputs(4314) <= (layer0_outputs(1606)) and (layer0_outputs(3511));
    layer1_outputs(4315) <= not(layer0_outputs(1115));
    layer1_outputs(4316) <= not((layer0_outputs(4810)) xor (layer0_outputs(3842)));
    layer1_outputs(4317) <= layer0_outputs(3397);
    layer1_outputs(4318) <= not(layer0_outputs(4712)) or (layer0_outputs(3291));
    layer1_outputs(4319) <= not(layer0_outputs(3496));
    layer1_outputs(4320) <= (layer0_outputs(3999)) and not (layer0_outputs(4288));
    layer1_outputs(4321) <= (layer0_outputs(3091)) or (layer0_outputs(2187));
    layer1_outputs(4322) <= layer0_outputs(2344);
    layer1_outputs(4323) <= (layer0_outputs(4986)) and (layer0_outputs(694));
    layer1_outputs(4324) <= not(layer0_outputs(297)) or (layer0_outputs(2058));
    layer1_outputs(4325) <= '1';
    layer1_outputs(4326) <= not(layer0_outputs(3601));
    layer1_outputs(4327) <= '0';
    layer1_outputs(4328) <= '1';
    layer1_outputs(4329) <= '1';
    layer1_outputs(4330) <= not((layer0_outputs(700)) and (layer0_outputs(2947)));
    layer1_outputs(4331) <= (layer0_outputs(3524)) and (layer0_outputs(4704));
    layer1_outputs(4332) <= not(layer0_outputs(4588));
    layer1_outputs(4333) <= '1';
    layer1_outputs(4334) <= not((layer0_outputs(820)) and (layer0_outputs(4321)));
    layer1_outputs(4335) <= (layer0_outputs(3349)) and (layer0_outputs(2309));
    layer1_outputs(4336) <= (layer0_outputs(1392)) or (layer0_outputs(80));
    layer1_outputs(4337) <= (layer0_outputs(410)) and not (layer0_outputs(4933));
    layer1_outputs(4338) <= (layer0_outputs(186)) or (layer0_outputs(3214));
    layer1_outputs(4339) <= (layer0_outputs(2476)) and not (layer0_outputs(2087));
    layer1_outputs(4340) <= not((layer0_outputs(1848)) or (layer0_outputs(3177)));
    layer1_outputs(4341) <= (layer0_outputs(3218)) and not (layer0_outputs(4201));
    layer1_outputs(4342) <= (layer0_outputs(2396)) or (layer0_outputs(288));
    layer1_outputs(4343) <= '0';
    layer1_outputs(4344) <= (layer0_outputs(3298)) and not (layer0_outputs(2159));
    layer1_outputs(4345) <= not(layer0_outputs(3220)) or (layer0_outputs(1207));
    layer1_outputs(4346) <= not(layer0_outputs(2126)) or (layer0_outputs(2060));
    layer1_outputs(4347) <= not(layer0_outputs(4291)) or (layer0_outputs(2044));
    layer1_outputs(4348) <= (layer0_outputs(1287)) and (layer0_outputs(532));
    layer1_outputs(4349) <= (layer0_outputs(2914)) or (layer0_outputs(850));
    layer1_outputs(4350) <= not((layer0_outputs(52)) or (layer0_outputs(4996)));
    layer1_outputs(4351) <= not(layer0_outputs(1831)) or (layer0_outputs(810));
    layer1_outputs(4352) <= not((layer0_outputs(4836)) and (layer0_outputs(241)));
    layer1_outputs(4353) <= '1';
    layer1_outputs(4354) <= layer0_outputs(3657);
    layer1_outputs(4355) <= '1';
    layer1_outputs(4356) <= not(layer0_outputs(2780)) or (layer0_outputs(3046));
    layer1_outputs(4357) <= not(layer0_outputs(4217)) or (layer0_outputs(123));
    layer1_outputs(4358) <= not((layer0_outputs(1361)) or (layer0_outputs(3530)));
    layer1_outputs(4359) <= '1';
    layer1_outputs(4360) <= not(layer0_outputs(3822)) or (layer0_outputs(2446));
    layer1_outputs(4361) <= (layer0_outputs(2230)) or (layer0_outputs(2192));
    layer1_outputs(4362) <= not(layer0_outputs(843)) or (layer0_outputs(1181));
    layer1_outputs(4363) <= layer0_outputs(4433);
    layer1_outputs(4364) <= (layer0_outputs(1871)) and not (layer0_outputs(1852));
    layer1_outputs(4365) <= not(layer0_outputs(1089));
    layer1_outputs(4366) <= (layer0_outputs(3791)) and not (layer0_outputs(831));
    layer1_outputs(4367) <= (layer0_outputs(4752)) and not (layer0_outputs(2824));
    layer1_outputs(4368) <= (layer0_outputs(2024)) and (layer0_outputs(4677));
    layer1_outputs(4369) <= '1';
    layer1_outputs(4370) <= (layer0_outputs(1448)) and (layer0_outputs(2971));
    layer1_outputs(4371) <= not((layer0_outputs(3826)) xor (layer0_outputs(3358)));
    layer1_outputs(4372) <= layer0_outputs(1465);
    layer1_outputs(4373) <= (layer0_outputs(2105)) or (layer0_outputs(855));
    layer1_outputs(4374) <= not(layer0_outputs(1963)) or (layer0_outputs(4572));
    layer1_outputs(4375) <= (layer0_outputs(4075)) and (layer0_outputs(4761));
    layer1_outputs(4376) <= '0';
    layer1_outputs(4377) <= not(layer0_outputs(1948)) or (layer0_outputs(2427));
    layer1_outputs(4378) <= '1';
    layer1_outputs(4379) <= '1';
    layer1_outputs(4380) <= (layer0_outputs(1832)) and not (layer0_outputs(3466));
    layer1_outputs(4381) <= '1';
    layer1_outputs(4382) <= (layer0_outputs(3489)) and not (layer0_outputs(1434));
    layer1_outputs(4383) <= (layer0_outputs(2487)) and not (layer0_outputs(3484));
    layer1_outputs(4384) <= not((layer0_outputs(1315)) and (layer0_outputs(3133)));
    layer1_outputs(4385) <= not(layer0_outputs(3453)) or (layer0_outputs(33));
    layer1_outputs(4386) <= '0';
    layer1_outputs(4387) <= '0';
    layer1_outputs(4388) <= (layer0_outputs(3236)) and (layer0_outputs(1554));
    layer1_outputs(4389) <= not((layer0_outputs(4550)) and (layer0_outputs(3172)));
    layer1_outputs(4390) <= not(layer0_outputs(3574)) or (layer0_outputs(974));
    layer1_outputs(4391) <= not(layer0_outputs(4062)) or (layer0_outputs(1609));
    layer1_outputs(4392) <= not(layer0_outputs(3978)) or (layer0_outputs(2670));
    layer1_outputs(4393) <= '0';
    layer1_outputs(4394) <= (layer0_outputs(2544)) or (layer0_outputs(4822));
    layer1_outputs(4395) <= not(layer0_outputs(4924)) or (layer0_outputs(4497));
    layer1_outputs(4396) <= (layer0_outputs(434)) or (layer0_outputs(3827));
    layer1_outputs(4397) <= (layer0_outputs(4863)) and not (layer0_outputs(2522));
    layer1_outputs(4398) <= not((layer0_outputs(2649)) or (layer0_outputs(1330)));
    layer1_outputs(4399) <= (layer0_outputs(2121)) and not (layer0_outputs(643));
    layer1_outputs(4400) <= layer0_outputs(3397);
    layer1_outputs(4401) <= layer0_outputs(4034);
    layer1_outputs(4402) <= '0';
    layer1_outputs(4403) <= not(layer0_outputs(3204));
    layer1_outputs(4404) <= not((layer0_outputs(794)) or (layer0_outputs(2163)));
    layer1_outputs(4405) <= not(layer0_outputs(2346));
    layer1_outputs(4406) <= not(layer0_outputs(734)) or (layer0_outputs(1888));
    layer1_outputs(4407) <= (layer0_outputs(930)) or (layer0_outputs(2405));
    layer1_outputs(4408) <= '1';
    layer1_outputs(4409) <= '1';
    layer1_outputs(4410) <= not((layer0_outputs(4401)) and (layer0_outputs(2638)));
    layer1_outputs(4411) <= '0';
    layer1_outputs(4412) <= '1';
    layer1_outputs(4413) <= '0';
    layer1_outputs(4414) <= (layer0_outputs(1409)) and not (layer0_outputs(4685));
    layer1_outputs(4415) <= not(layer0_outputs(1486));
    layer1_outputs(4416) <= (layer0_outputs(4427)) and not (layer0_outputs(2260));
    layer1_outputs(4417) <= (layer0_outputs(3101)) xor (layer0_outputs(5058));
    layer1_outputs(4418) <= (layer0_outputs(1546)) and not (layer0_outputs(3910));
    layer1_outputs(4419) <= not(layer0_outputs(1660)) or (layer0_outputs(1994));
    layer1_outputs(4420) <= (layer0_outputs(2933)) and not (layer0_outputs(2870));
    layer1_outputs(4421) <= '1';
    layer1_outputs(4422) <= not(layer0_outputs(2839));
    layer1_outputs(4423) <= not(layer0_outputs(10)) or (layer0_outputs(1193));
    layer1_outputs(4424) <= '1';
    layer1_outputs(4425) <= not(layer0_outputs(1191));
    layer1_outputs(4426) <= '0';
    layer1_outputs(4427) <= '0';
    layer1_outputs(4428) <= layer0_outputs(3094);
    layer1_outputs(4429) <= not(layer0_outputs(2077));
    layer1_outputs(4430) <= (layer0_outputs(390)) and (layer0_outputs(3951));
    layer1_outputs(4431) <= not((layer0_outputs(4839)) and (layer0_outputs(1076)));
    layer1_outputs(4432) <= layer0_outputs(3493);
    layer1_outputs(4433) <= '0';
    layer1_outputs(4434) <= '1';
    layer1_outputs(4435) <= (layer0_outputs(968)) or (layer0_outputs(4512));
    layer1_outputs(4436) <= not(layer0_outputs(1944)) or (layer0_outputs(2508));
    layer1_outputs(4437) <= not(layer0_outputs(4024)) or (layer0_outputs(2356));
    layer1_outputs(4438) <= not(layer0_outputs(140)) or (layer0_outputs(3465));
    layer1_outputs(4439) <= '1';
    layer1_outputs(4440) <= '1';
    layer1_outputs(4441) <= '0';
    layer1_outputs(4442) <= '1';
    layer1_outputs(4443) <= not(layer0_outputs(1867));
    layer1_outputs(4444) <= '0';
    layer1_outputs(4445) <= not(layer0_outputs(120));
    layer1_outputs(4446) <= layer0_outputs(2714);
    layer1_outputs(4447) <= not(layer0_outputs(2191));
    layer1_outputs(4448) <= (layer0_outputs(3315)) and not (layer0_outputs(1834));
    layer1_outputs(4449) <= not(layer0_outputs(875));
    layer1_outputs(4450) <= layer0_outputs(1209);
    layer1_outputs(4451) <= not(layer0_outputs(4968)) or (layer0_outputs(4204));
    layer1_outputs(4452) <= '0';
    layer1_outputs(4453) <= '1';
    layer1_outputs(4454) <= '0';
    layer1_outputs(4455) <= '0';
    layer1_outputs(4456) <= layer0_outputs(696);
    layer1_outputs(4457) <= not(layer0_outputs(3053)) or (layer0_outputs(1062));
    layer1_outputs(4458) <= not((layer0_outputs(2860)) or (layer0_outputs(3626)));
    layer1_outputs(4459) <= (layer0_outputs(4888)) and not (layer0_outputs(1271));
    layer1_outputs(4460) <= not((layer0_outputs(2814)) and (layer0_outputs(3706)));
    layer1_outputs(4461) <= not(layer0_outputs(35));
    layer1_outputs(4462) <= '0';
    layer1_outputs(4463) <= '1';
    layer1_outputs(4464) <= not((layer0_outputs(3297)) and (layer0_outputs(600)));
    layer1_outputs(4465) <= layer0_outputs(2909);
    layer1_outputs(4466) <= (layer0_outputs(1211)) and not (layer0_outputs(1333));
    layer1_outputs(4467) <= '0';
    layer1_outputs(4468) <= (layer0_outputs(4383)) or (layer0_outputs(174));
    layer1_outputs(4469) <= not((layer0_outputs(4645)) or (layer0_outputs(2896)));
    layer1_outputs(4470) <= '0';
    layer1_outputs(4471) <= (layer0_outputs(3512)) and not (layer0_outputs(846));
    layer1_outputs(4472) <= not(layer0_outputs(7)) or (layer0_outputs(1732));
    layer1_outputs(4473) <= not(layer0_outputs(3006));
    layer1_outputs(4474) <= '0';
    layer1_outputs(4475) <= not((layer0_outputs(419)) and (layer0_outputs(3895)));
    layer1_outputs(4476) <= layer0_outputs(2900);
    layer1_outputs(4477) <= '0';
    layer1_outputs(4478) <= not((layer0_outputs(4055)) or (layer0_outputs(1042)));
    layer1_outputs(4479) <= not((layer0_outputs(1079)) or (layer0_outputs(2602)));
    layer1_outputs(4480) <= (layer0_outputs(2956)) and not (layer0_outputs(423));
    layer1_outputs(4481) <= not(layer0_outputs(2455)) or (layer0_outputs(823));
    layer1_outputs(4482) <= (layer0_outputs(972)) and (layer0_outputs(1743));
    layer1_outputs(4483) <= '1';
    layer1_outputs(4484) <= not((layer0_outputs(1384)) and (layer0_outputs(4729)));
    layer1_outputs(4485) <= '0';
    layer1_outputs(4486) <= not(layer0_outputs(3426)) or (layer0_outputs(3992));
    layer1_outputs(4487) <= layer0_outputs(4271);
    layer1_outputs(4488) <= not((layer0_outputs(3382)) or (layer0_outputs(1795)));
    layer1_outputs(4489) <= (layer0_outputs(3628)) and (layer0_outputs(2312));
    layer1_outputs(4490) <= not((layer0_outputs(3305)) or (layer0_outputs(285)));
    layer1_outputs(4491) <= '1';
    layer1_outputs(4492) <= not(layer0_outputs(281)) or (layer0_outputs(4780));
    layer1_outputs(4493) <= '1';
    layer1_outputs(4494) <= not(layer0_outputs(4087));
    layer1_outputs(4495) <= '1';
    layer1_outputs(4496) <= (layer0_outputs(3324)) or (layer0_outputs(1192));
    layer1_outputs(4497) <= (layer0_outputs(2648)) and not (layer0_outputs(1807));
    layer1_outputs(4498) <= not(layer0_outputs(1026)) or (layer0_outputs(5068));
    layer1_outputs(4499) <= not(layer0_outputs(4181)) or (layer0_outputs(1953));
    layer1_outputs(4500) <= '0';
    layer1_outputs(4501) <= not(layer0_outputs(3884)) or (layer0_outputs(4318));
    layer1_outputs(4502) <= not(layer0_outputs(2831)) or (layer0_outputs(4576));
    layer1_outputs(4503) <= (layer0_outputs(3246)) or (layer0_outputs(4359));
    layer1_outputs(4504) <= layer0_outputs(86);
    layer1_outputs(4505) <= (layer0_outputs(144)) and not (layer0_outputs(225));
    layer1_outputs(4506) <= '0';
    layer1_outputs(4507) <= layer0_outputs(4265);
    layer1_outputs(4508) <= not(layer0_outputs(2427)) or (layer0_outputs(1552));
    layer1_outputs(4509) <= (layer0_outputs(3265)) or (layer0_outputs(411));
    layer1_outputs(4510) <= not((layer0_outputs(90)) or (layer0_outputs(3314)));
    layer1_outputs(4511) <= layer0_outputs(4041);
    layer1_outputs(4512) <= '0';
    layer1_outputs(4513) <= not((layer0_outputs(2630)) or (layer0_outputs(2566)));
    layer1_outputs(4514) <= not(layer0_outputs(2261));
    layer1_outputs(4515) <= layer0_outputs(1927);
    layer1_outputs(4516) <= '1';
    layer1_outputs(4517) <= (layer0_outputs(4619)) and not (layer0_outputs(99));
    layer1_outputs(4518) <= not(layer0_outputs(1048)) or (layer0_outputs(1246));
    layer1_outputs(4519) <= not(layer0_outputs(1710)) or (layer0_outputs(4101));
    layer1_outputs(4520) <= layer0_outputs(602);
    layer1_outputs(4521) <= not(layer0_outputs(3036)) or (layer0_outputs(2490));
    layer1_outputs(4522) <= '0';
    layer1_outputs(4523) <= not((layer0_outputs(4649)) or (layer0_outputs(3514)));
    layer1_outputs(4524) <= (layer0_outputs(4464)) or (layer0_outputs(4087));
    layer1_outputs(4525) <= '0';
    layer1_outputs(4526) <= layer0_outputs(4660);
    layer1_outputs(4527) <= '1';
    layer1_outputs(4528) <= layer0_outputs(169);
    layer1_outputs(4529) <= not(layer0_outputs(3624)) or (layer0_outputs(5112));
    layer1_outputs(4530) <= (layer0_outputs(2653)) xor (layer0_outputs(1345));
    layer1_outputs(4531) <= '1';
    layer1_outputs(4532) <= not(layer0_outputs(3340)) or (layer0_outputs(2667));
    layer1_outputs(4533) <= not(layer0_outputs(3929)) or (layer0_outputs(1104));
    layer1_outputs(4534) <= '1';
    layer1_outputs(4535) <= (layer0_outputs(84)) and not (layer0_outputs(2076));
    layer1_outputs(4536) <= (layer0_outputs(25)) and not (layer0_outputs(3639));
    layer1_outputs(4537) <= (layer0_outputs(584)) and not (layer0_outputs(3914));
    layer1_outputs(4538) <= '1';
    layer1_outputs(4539) <= (layer0_outputs(2988)) and not (layer0_outputs(675));
    layer1_outputs(4540) <= not((layer0_outputs(3674)) or (layer0_outputs(1913)));
    layer1_outputs(4541) <= (layer0_outputs(4940)) and not (layer0_outputs(5066));
    layer1_outputs(4542) <= '0';
    layer1_outputs(4543) <= '0';
    layer1_outputs(4544) <= not(layer0_outputs(2398)) or (layer0_outputs(869));
    layer1_outputs(4545) <= not(layer0_outputs(1174)) or (layer0_outputs(4937));
    layer1_outputs(4546) <= (layer0_outputs(1155)) and not (layer0_outputs(2823));
    layer1_outputs(4547) <= '0';
    layer1_outputs(4548) <= not(layer0_outputs(4523));
    layer1_outputs(4549) <= '1';
    layer1_outputs(4550) <= '0';
    layer1_outputs(4551) <= layer0_outputs(2620);
    layer1_outputs(4552) <= not((layer0_outputs(914)) and (layer0_outputs(1725)));
    layer1_outputs(4553) <= (layer0_outputs(4113)) and not (layer0_outputs(1158));
    layer1_outputs(4554) <= layer0_outputs(1131);
    layer1_outputs(4555) <= '0';
    layer1_outputs(4556) <= (layer0_outputs(781)) and not (layer0_outputs(4380));
    layer1_outputs(4557) <= '1';
    layer1_outputs(4558) <= not((layer0_outputs(547)) or (layer0_outputs(4253)));
    layer1_outputs(4559) <= not(layer0_outputs(3732)) or (layer0_outputs(2903));
    layer1_outputs(4560) <= not(layer0_outputs(2296));
    layer1_outputs(4561) <= layer0_outputs(1783);
    layer1_outputs(4562) <= '1';
    layer1_outputs(4563) <= (layer0_outputs(4422)) and not (layer0_outputs(1839));
    layer1_outputs(4564) <= layer0_outputs(4794);
    layer1_outputs(4565) <= (layer0_outputs(5020)) or (layer0_outputs(1438));
    layer1_outputs(4566) <= not(layer0_outputs(4156)) or (layer0_outputs(660));
    layer1_outputs(4567) <= not(layer0_outputs(755));
    layer1_outputs(4568) <= (layer0_outputs(3246)) or (layer0_outputs(1403));
    layer1_outputs(4569) <= not(layer0_outputs(2145)) or (layer0_outputs(2379));
    layer1_outputs(4570) <= (layer0_outputs(1307)) or (layer0_outputs(4515));
    layer1_outputs(4571) <= '1';
    layer1_outputs(4572) <= not(layer0_outputs(806)) or (layer0_outputs(2122));
    layer1_outputs(4573) <= layer0_outputs(3662);
    layer1_outputs(4574) <= '1';
    layer1_outputs(4575) <= not((layer0_outputs(2582)) or (layer0_outputs(1958)));
    layer1_outputs(4576) <= not(layer0_outputs(3366)) or (layer0_outputs(4434));
    layer1_outputs(4577) <= '1';
    layer1_outputs(4578) <= not(layer0_outputs(1051)) or (layer0_outputs(1659));
    layer1_outputs(4579) <= not((layer0_outputs(3652)) or (layer0_outputs(2247)));
    layer1_outputs(4580) <= not((layer0_outputs(4687)) and (layer0_outputs(1546)));
    layer1_outputs(4581) <= layer0_outputs(2883);
    layer1_outputs(4582) <= layer0_outputs(376);
    layer1_outputs(4583) <= layer0_outputs(31);
    layer1_outputs(4584) <= '0';
    layer1_outputs(4585) <= (layer0_outputs(104)) and (layer0_outputs(2216));
    layer1_outputs(4586) <= layer0_outputs(4889);
    layer1_outputs(4587) <= (layer0_outputs(3451)) and not (layer0_outputs(4506));
    layer1_outputs(4588) <= (layer0_outputs(2879)) and not (layer0_outputs(3314));
    layer1_outputs(4589) <= layer0_outputs(3850);
    layer1_outputs(4590) <= '0';
    layer1_outputs(4591) <= not(layer0_outputs(2674)) or (layer0_outputs(705));
    layer1_outputs(4592) <= '1';
    layer1_outputs(4593) <= '0';
    layer1_outputs(4594) <= not(layer0_outputs(1597)) or (layer0_outputs(4814));
    layer1_outputs(4595) <= '1';
    layer1_outputs(4596) <= not(layer0_outputs(4592)) or (layer0_outputs(2945));
    layer1_outputs(4597) <= (layer0_outputs(216)) and (layer0_outputs(470));
    layer1_outputs(4598) <= (layer0_outputs(4859)) or (layer0_outputs(1283));
    layer1_outputs(4599) <= (layer0_outputs(3898)) and (layer0_outputs(1152));
    layer1_outputs(4600) <= not(layer0_outputs(3969));
    layer1_outputs(4601) <= not((layer0_outputs(2965)) and (layer0_outputs(2479)));
    layer1_outputs(4602) <= '1';
    layer1_outputs(4603) <= (layer0_outputs(1098)) and not (layer0_outputs(2522));
    layer1_outputs(4604) <= layer0_outputs(290);
    layer1_outputs(4605) <= '1';
    layer1_outputs(4606) <= not(layer0_outputs(4405));
    layer1_outputs(4607) <= '1';
    layer1_outputs(4608) <= layer0_outputs(3809);
    layer1_outputs(4609) <= not((layer0_outputs(4112)) or (layer0_outputs(509)));
    layer1_outputs(4610) <= (layer0_outputs(1139)) and not (layer0_outputs(137));
    layer1_outputs(4611) <= layer0_outputs(1503);
    layer1_outputs(4612) <= (layer0_outputs(3959)) xor (layer0_outputs(5106));
    layer1_outputs(4613) <= not((layer0_outputs(561)) and (layer0_outputs(1981)));
    layer1_outputs(4614) <= layer0_outputs(1088);
    layer1_outputs(4615) <= (layer0_outputs(5092)) and (layer0_outputs(964));
    layer1_outputs(4616) <= '0';
    layer1_outputs(4617) <= not(layer0_outputs(3323));
    layer1_outputs(4618) <= (layer0_outputs(1634)) or (layer0_outputs(1474));
    layer1_outputs(4619) <= not(layer0_outputs(4727)) or (layer0_outputs(133));
    layer1_outputs(4620) <= '0';
    layer1_outputs(4621) <= (layer0_outputs(357)) and (layer0_outputs(3095));
    layer1_outputs(4622) <= not(layer0_outputs(1853)) or (layer0_outputs(2326));
    layer1_outputs(4623) <= '0';
    layer1_outputs(4624) <= (layer0_outputs(2276)) and (layer0_outputs(4232));
    layer1_outputs(4625) <= layer0_outputs(3114);
    layer1_outputs(4626) <= '0';
    layer1_outputs(4627) <= layer0_outputs(4402);
    layer1_outputs(4628) <= layer0_outputs(247);
    layer1_outputs(4629) <= (layer0_outputs(4436)) and not (layer0_outputs(2344));
    layer1_outputs(4630) <= not((layer0_outputs(945)) and (layer0_outputs(658)));
    layer1_outputs(4631) <= not(layer0_outputs(3087));
    layer1_outputs(4632) <= not((layer0_outputs(2754)) or (layer0_outputs(1576)));
    layer1_outputs(4633) <= '1';
    layer1_outputs(4634) <= '1';
    layer1_outputs(4635) <= (layer0_outputs(3571)) and (layer0_outputs(1270));
    layer1_outputs(4636) <= '1';
    layer1_outputs(4637) <= '0';
    layer1_outputs(4638) <= not((layer0_outputs(1260)) or (layer0_outputs(2954)));
    layer1_outputs(4639) <= not(layer0_outputs(2048));
    layer1_outputs(4640) <= (layer0_outputs(3893)) and not (layer0_outputs(4431));
    layer1_outputs(4641) <= layer0_outputs(5102);
    layer1_outputs(4642) <= not((layer0_outputs(2371)) or (layer0_outputs(2703)));
    layer1_outputs(4643) <= not(layer0_outputs(502));
    layer1_outputs(4644) <= layer0_outputs(4066);
    layer1_outputs(4645) <= not(layer0_outputs(147)) or (layer0_outputs(2373));
    layer1_outputs(4646) <= not((layer0_outputs(931)) and (layer0_outputs(2219)));
    layer1_outputs(4647) <= (layer0_outputs(3863)) and not (layer0_outputs(2220));
    layer1_outputs(4648) <= (layer0_outputs(4304)) and not (layer0_outputs(2531));
    layer1_outputs(4649) <= not(layer0_outputs(785));
    layer1_outputs(4650) <= (layer0_outputs(1058)) xor (layer0_outputs(777));
    layer1_outputs(4651) <= not((layer0_outputs(925)) xor (layer0_outputs(4353)));
    layer1_outputs(4652) <= (layer0_outputs(2634)) or (layer0_outputs(2208));
    layer1_outputs(4653) <= '0';
    layer1_outputs(4654) <= not(layer0_outputs(2733)) or (layer0_outputs(3172));
    layer1_outputs(4655) <= not((layer0_outputs(4708)) or (layer0_outputs(2868)));
    layer1_outputs(4656) <= not((layer0_outputs(1933)) or (layer0_outputs(1569)));
    layer1_outputs(4657) <= '0';
    layer1_outputs(4658) <= not((layer0_outputs(900)) and (layer0_outputs(616)));
    layer1_outputs(4659) <= not((layer0_outputs(1329)) and (layer0_outputs(749)));
    layer1_outputs(4660) <= layer0_outputs(347);
    layer1_outputs(4661) <= '0';
    layer1_outputs(4662) <= '0';
    layer1_outputs(4663) <= not(layer0_outputs(1014)) or (layer0_outputs(2124));
    layer1_outputs(4664) <= not(layer0_outputs(3965));
    layer1_outputs(4665) <= not((layer0_outputs(948)) and (layer0_outputs(3474)));
    layer1_outputs(4666) <= not((layer0_outputs(5091)) or (layer0_outputs(1680)));
    layer1_outputs(4667) <= (layer0_outputs(2928)) and not (layer0_outputs(20));
    layer1_outputs(4668) <= not(layer0_outputs(3055)) or (layer0_outputs(2619));
    layer1_outputs(4669) <= layer0_outputs(1235);
    layer1_outputs(4670) <= '1';
    layer1_outputs(4671) <= not(layer0_outputs(2554)) or (layer0_outputs(2537));
    layer1_outputs(4672) <= '1';
    layer1_outputs(4673) <= not(layer0_outputs(4096)) or (layer0_outputs(1785));
    layer1_outputs(4674) <= (layer0_outputs(1391)) and not (layer0_outputs(5034));
    layer1_outputs(4675) <= (layer0_outputs(3226)) and not (layer0_outputs(3882));
    layer1_outputs(4676) <= not(layer0_outputs(2721)) or (layer0_outputs(3221));
    layer1_outputs(4677) <= not((layer0_outputs(1436)) and (layer0_outputs(351)));
    layer1_outputs(4678) <= layer0_outputs(3694);
    layer1_outputs(4679) <= not(layer0_outputs(3832));
    layer1_outputs(4680) <= '1';
    layer1_outputs(4681) <= not((layer0_outputs(3628)) or (layer0_outputs(60)));
    layer1_outputs(4682) <= '1';
    layer1_outputs(4683) <= not(layer0_outputs(2420)) or (layer0_outputs(2424));
    layer1_outputs(4684) <= not(layer0_outputs(2696)) or (layer0_outputs(508));
    layer1_outputs(4685) <= '0';
    layer1_outputs(4686) <= '0';
    layer1_outputs(4687) <= not(layer0_outputs(3205)) or (layer0_outputs(5053));
    layer1_outputs(4688) <= '1';
    layer1_outputs(4689) <= (layer0_outputs(648)) and not (layer0_outputs(2321));
    layer1_outputs(4690) <= (layer0_outputs(2134)) or (layer0_outputs(1990));
    layer1_outputs(4691) <= (layer0_outputs(930)) and not (layer0_outputs(1437));
    layer1_outputs(4692) <= '0';
    layer1_outputs(4693) <= (layer0_outputs(1086)) or (layer0_outputs(3633));
    layer1_outputs(4694) <= not(layer0_outputs(3697)) or (layer0_outputs(1056));
    layer1_outputs(4695) <= not(layer0_outputs(1896)) or (layer0_outputs(1796));
    layer1_outputs(4696) <= not(layer0_outputs(1408)) or (layer0_outputs(3158));
    layer1_outputs(4697) <= not(layer0_outputs(98)) or (layer0_outputs(5079));
    layer1_outputs(4698) <= not((layer0_outputs(2269)) or (layer0_outputs(3564)));
    layer1_outputs(4699) <= '0';
    layer1_outputs(4700) <= not(layer0_outputs(581));
    layer1_outputs(4701) <= (layer0_outputs(2642)) and not (layer0_outputs(2503));
    layer1_outputs(4702) <= not((layer0_outputs(3560)) xor (layer0_outputs(93)));
    layer1_outputs(4703) <= (layer0_outputs(924)) and not (layer0_outputs(3561));
    layer1_outputs(4704) <= not(layer0_outputs(4334)) or (layer0_outputs(2560));
    layer1_outputs(4705) <= '1';
    layer1_outputs(4706) <= (layer0_outputs(4831)) and (layer0_outputs(1593));
    layer1_outputs(4707) <= not(layer0_outputs(2348)) or (layer0_outputs(4088));
    layer1_outputs(4708) <= not(layer0_outputs(4525));
    layer1_outputs(4709) <= '1';
    layer1_outputs(4710) <= '1';
    layer1_outputs(4711) <= not(layer0_outputs(2893));
    layer1_outputs(4712) <= '0';
    layer1_outputs(4713) <= '0';
    layer1_outputs(4714) <= '1';
    layer1_outputs(4715) <= '1';
    layer1_outputs(4716) <= '1';
    layer1_outputs(4717) <= '0';
    layer1_outputs(4718) <= layer0_outputs(647);
    layer1_outputs(4719) <= (layer0_outputs(440)) and not (layer0_outputs(1610));
    layer1_outputs(4720) <= '0';
    layer1_outputs(4721) <= not(layer0_outputs(2807));
    layer1_outputs(4722) <= (layer0_outputs(4596)) and not (layer0_outputs(2746));
    layer1_outputs(4723) <= not(layer0_outputs(4050));
    layer1_outputs(4724) <= (layer0_outputs(2563)) and not (layer0_outputs(1629));
    layer1_outputs(4725) <= not((layer0_outputs(3938)) or (layer0_outputs(4769)));
    layer1_outputs(4726) <= not(layer0_outputs(2377)) or (layer0_outputs(3305));
    layer1_outputs(4727) <= '1';
    layer1_outputs(4728) <= '0';
    layer1_outputs(4729) <= not(layer0_outputs(2265)) or (layer0_outputs(2332));
    layer1_outputs(4730) <= not((layer0_outputs(697)) and (layer0_outputs(555)));
    layer1_outputs(4731) <= layer0_outputs(341);
    layer1_outputs(4732) <= '0';
    layer1_outputs(4733) <= (layer0_outputs(2131)) and not (layer0_outputs(4589));
    layer1_outputs(4734) <= layer0_outputs(1134);
    layer1_outputs(4735) <= '1';
    layer1_outputs(4736) <= not(layer0_outputs(1826)) or (layer0_outputs(4450));
    layer1_outputs(4737) <= (layer0_outputs(2302)) and not (layer0_outputs(1876));
    layer1_outputs(4738) <= not(layer0_outputs(2251)) or (layer0_outputs(2610));
    layer1_outputs(4739) <= not((layer0_outputs(720)) or (layer0_outputs(1363)));
    layer1_outputs(4740) <= (layer0_outputs(2668)) and not (layer0_outputs(2112));
    layer1_outputs(4741) <= '1';
    layer1_outputs(4742) <= '0';
    layer1_outputs(4743) <= (layer0_outputs(3440)) or (layer0_outputs(2916));
    layer1_outputs(4744) <= not(layer0_outputs(1229)) or (layer0_outputs(2190));
    layer1_outputs(4745) <= not(layer0_outputs(1625));
    layer1_outputs(4746) <= not(layer0_outputs(2322));
    layer1_outputs(4747) <= not(layer0_outputs(589));
    layer1_outputs(4748) <= not((layer0_outputs(2658)) and (layer0_outputs(1544)));
    layer1_outputs(4749) <= '0';
    layer1_outputs(4750) <= not(layer0_outputs(64)) or (layer0_outputs(1687));
    layer1_outputs(4751) <= (layer0_outputs(2752)) or (layer0_outputs(3836));
    layer1_outputs(4752) <= (layer0_outputs(4597)) or (layer0_outputs(4530));
    layer1_outputs(4753) <= '0';
    layer1_outputs(4754) <= '0';
    layer1_outputs(4755) <= '0';
    layer1_outputs(4756) <= (layer0_outputs(3817)) and not (layer0_outputs(4543));
    layer1_outputs(4757) <= (layer0_outputs(1231)) and (layer0_outputs(2394));
    layer1_outputs(4758) <= not(layer0_outputs(3756)) or (layer0_outputs(4606));
    layer1_outputs(4759) <= not(layer0_outputs(1637));
    layer1_outputs(4760) <= not(layer0_outputs(2728));
    layer1_outputs(4761) <= not(layer0_outputs(3048)) or (layer0_outputs(1376));
    layer1_outputs(4762) <= (layer0_outputs(4439)) and (layer0_outputs(4305));
    layer1_outputs(4763) <= (layer0_outputs(545)) and not (layer0_outputs(2109));
    layer1_outputs(4764) <= not(layer0_outputs(2382)) or (layer0_outputs(3930));
    layer1_outputs(4765) <= not(layer0_outputs(4182)) or (layer0_outputs(3854));
    layer1_outputs(4766) <= (layer0_outputs(1400)) and not (layer0_outputs(868));
    layer1_outputs(4767) <= not((layer0_outputs(3721)) and (layer0_outputs(2594)));
    layer1_outputs(4768) <= '1';
    layer1_outputs(4769) <= not(layer0_outputs(3278)) or (layer0_outputs(5056));
    layer1_outputs(4770) <= (layer0_outputs(3232)) and not (layer0_outputs(826));
    layer1_outputs(4771) <= (layer0_outputs(3640)) and not (layer0_outputs(939));
    layer1_outputs(4772) <= '1';
    layer1_outputs(4773) <= (layer0_outputs(1209)) and not (layer0_outputs(3408));
    layer1_outputs(4774) <= layer0_outputs(3774);
    layer1_outputs(4775) <= not((layer0_outputs(3070)) and (layer0_outputs(316)));
    layer1_outputs(4776) <= (layer0_outputs(3295)) and (layer0_outputs(1221));
    layer1_outputs(4777) <= (layer0_outputs(3164)) and not (layer0_outputs(857));
    layer1_outputs(4778) <= (layer0_outputs(4440)) or (layer0_outputs(2448));
    layer1_outputs(4779) <= not((layer0_outputs(201)) xor (layer0_outputs(3442)));
    layer1_outputs(4780) <= (layer0_outputs(2177)) and not (layer0_outputs(1982));
    layer1_outputs(4781) <= layer0_outputs(284);
    layer1_outputs(4782) <= not((layer0_outputs(921)) and (layer0_outputs(3977)));
    layer1_outputs(4783) <= (layer0_outputs(908)) and not (layer0_outputs(2934));
    layer1_outputs(4784) <= '0';
    layer1_outputs(4785) <= '1';
    layer1_outputs(4786) <= (layer0_outputs(4016)) and (layer0_outputs(1558));
    layer1_outputs(4787) <= not(layer0_outputs(4237)) or (layer0_outputs(4603));
    layer1_outputs(4788) <= '0';
    layer1_outputs(4789) <= not(layer0_outputs(1240));
    layer1_outputs(4790) <= (layer0_outputs(3337)) and not (layer0_outputs(1604));
    layer1_outputs(4791) <= not(layer0_outputs(2784)) or (layer0_outputs(1737));
    layer1_outputs(4792) <= (layer0_outputs(2820)) xor (layer0_outputs(3169));
    layer1_outputs(4793) <= not((layer0_outputs(4393)) or (layer0_outputs(1885)));
    layer1_outputs(4794) <= '0';
    layer1_outputs(4795) <= not((layer0_outputs(4310)) or (layer0_outputs(2953)));
    layer1_outputs(4796) <= '0';
    layer1_outputs(4797) <= (layer0_outputs(164)) and not (layer0_outputs(5093));
    layer1_outputs(4798) <= '1';
    layer1_outputs(4799) <= '0';
    layer1_outputs(4800) <= '0';
    layer1_outputs(4801) <= not((layer0_outputs(2334)) and (layer0_outputs(1904)));
    layer1_outputs(4802) <= layer0_outputs(3733);
    layer1_outputs(4803) <= '0';
    layer1_outputs(4804) <= '0';
    layer1_outputs(4805) <= not(layer0_outputs(1556)) or (layer0_outputs(2156));
    layer1_outputs(4806) <= '0';
    layer1_outputs(4807) <= (layer0_outputs(210)) or (layer0_outputs(3542));
    layer1_outputs(4808) <= (layer0_outputs(836)) and not (layer0_outputs(3180));
    layer1_outputs(4809) <= (layer0_outputs(4308)) and (layer0_outputs(1498));
    layer1_outputs(4810) <= (layer0_outputs(609)) or (layer0_outputs(944));
    layer1_outputs(4811) <= layer0_outputs(4140);
    layer1_outputs(4812) <= '0';
    layer1_outputs(4813) <= '1';
    layer1_outputs(4814) <= layer0_outputs(2869);
    layer1_outputs(4815) <= layer0_outputs(4129);
    layer1_outputs(4816) <= not((layer0_outputs(1393)) or (layer0_outputs(4528)));
    layer1_outputs(4817) <= '0';
    layer1_outputs(4818) <= (layer0_outputs(2513)) and not (layer0_outputs(1603));
    layer1_outputs(4819) <= '0';
    layer1_outputs(4820) <= (layer0_outputs(4152)) and (layer0_outputs(406));
    layer1_outputs(4821) <= (layer0_outputs(2614)) and not (layer0_outputs(244));
    layer1_outputs(4822) <= (layer0_outputs(354)) or (layer0_outputs(3862));
    layer1_outputs(4823) <= '0';
    layer1_outputs(4824) <= '0';
    layer1_outputs(4825) <= '1';
    layer1_outputs(4826) <= not((layer0_outputs(1240)) and (layer0_outputs(565)));
    layer1_outputs(4827) <= not(layer0_outputs(818)) or (layer0_outputs(4255));
    layer1_outputs(4828) <= '1';
    layer1_outputs(4829) <= (layer0_outputs(1150)) and not (layer0_outputs(227));
    layer1_outputs(4830) <= not((layer0_outputs(2139)) or (layer0_outputs(1598)));
    layer1_outputs(4831) <= (layer0_outputs(4172)) and (layer0_outputs(2371));
    layer1_outputs(4832) <= not((layer0_outputs(1669)) or (layer0_outputs(797)));
    layer1_outputs(4833) <= '0';
    layer1_outputs(4834) <= (layer0_outputs(1112)) and not (layer0_outputs(1009));
    layer1_outputs(4835) <= not((layer0_outputs(311)) and (layer0_outputs(3462)));
    layer1_outputs(4836) <= '0';
    layer1_outputs(4837) <= not(layer0_outputs(1992)) or (layer0_outputs(766));
    layer1_outputs(4838) <= '1';
    layer1_outputs(4839) <= not((layer0_outputs(3538)) or (layer0_outputs(4962)));
    layer1_outputs(4840) <= (layer0_outputs(1031)) or (layer0_outputs(5010));
    layer1_outputs(4841) <= not(layer0_outputs(4257)) or (layer0_outputs(4290));
    layer1_outputs(4842) <= not(layer0_outputs(1662));
    layer1_outputs(4843) <= '0';
    layer1_outputs(4844) <= (layer0_outputs(1550)) and not (layer0_outputs(571));
    layer1_outputs(4845) <= (layer0_outputs(2655)) and not (layer0_outputs(2127));
    layer1_outputs(4846) <= (layer0_outputs(5112)) or (layer0_outputs(3354));
    layer1_outputs(4847) <= (layer0_outputs(3141)) and not (layer0_outputs(4799));
    layer1_outputs(4848) <= not((layer0_outputs(3226)) and (layer0_outputs(3985)));
    layer1_outputs(4849) <= not(layer0_outputs(4802));
    layer1_outputs(4850) <= not((layer0_outputs(3295)) or (layer0_outputs(4743)));
    layer1_outputs(4851) <= not(layer0_outputs(1751));
    layer1_outputs(4852) <= (layer0_outputs(4259)) and not (layer0_outputs(701));
    layer1_outputs(4853) <= (layer0_outputs(4554)) or (layer0_outputs(1267));
    layer1_outputs(4854) <= '0';
    layer1_outputs(4855) <= '0';
    layer1_outputs(4856) <= '0';
    layer1_outputs(4857) <= layer0_outputs(3378);
    layer1_outputs(4858) <= '0';
    layer1_outputs(4859) <= '0';
    layer1_outputs(4860) <= not(layer0_outputs(459)) or (layer0_outputs(897));
    layer1_outputs(4861) <= not((layer0_outputs(3618)) or (layer0_outputs(667)));
    layer1_outputs(4862) <= (layer0_outputs(3792)) and (layer0_outputs(2241));
    layer1_outputs(4863) <= (layer0_outputs(4031)) or (layer0_outputs(4279));
    layer1_outputs(4864) <= not(layer0_outputs(2398)) or (layer0_outputs(1416));
    layer1_outputs(4865) <= not(layer0_outputs(5073)) or (layer0_outputs(832));
    layer1_outputs(4866) <= layer0_outputs(5059);
    layer1_outputs(4867) <= (layer0_outputs(3142)) and not (layer0_outputs(2958));
    layer1_outputs(4868) <= not(layer0_outputs(5107));
    layer1_outputs(4869) <= not(layer0_outputs(2165)) or (layer0_outputs(426));
    layer1_outputs(4870) <= layer0_outputs(563);
    layer1_outputs(4871) <= layer0_outputs(288);
    layer1_outputs(4872) <= (layer0_outputs(465)) and (layer0_outputs(4146));
    layer1_outputs(4873) <= (layer0_outputs(1822)) and not (layer0_outputs(2968));
    layer1_outputs(4874) <= (layer0_outputs(598)) and (layer0_outputs(557));
    layer1_outputs(4875) <= (layer0_outputs(552)) and not (layer0_outputs(817));
    layer1_outputs(4876) <= '0';
    layer1_outputs(4877) <= (layer0_outputs(1491)) and not (layer0_outputs(2347));
    layer1_outputs(4878) <= (layer0_outputs(2491)) and not (layer0_outputs(250));
    layer1_outputs(4879) <= (layer0_outputs(1415)) and not (layer0_outputs(2756));
    layer1_outputs(4880) <= '1';
    layer1_outputs(4881) <= not(layer0_outputs(722)) or (layer0_outputs(3545));
    layer1_outputs(4882) <= (layer0_outputs(4340)) and (layer0_outputs(3794));
    layer1_outputs(4883) <= '1';
    layer1_outputs(4884) <= '1';
    layer1_outputs(4885) <= not((layer0_outputs(1218)) and (layer0_outputs(5115)));
    layer1_outputs(4886) <= (layer0_outputs(655)) and (layer0_outputs(4272));
    layer1_outputs(4887) <= not((layer0_outputs(3217)) and (layer0_outputs(2986)));
    layer1_outputs(4888) <= not((layer0_outputs(1631)) or (layer0_outputs(4777)));
    layer1_outputs(4889) <= '0';
    layer1_outputs(4890) <= '1';
    layer1_outputs(4891) <= not(layer0_outputs(4330)) or (layer0_outputs(3259));
    layer1_outputs(4892) <= not((layer0_outputs(4029)) and (layer0_outputs(62)));
    layer1_outputs(4893) <= not(layer0_outputs(2121)) or (layer0_outputs(379));
    layer1_outputs(4894) <= (layer0_outputs(895)) and (layer0_outputs(1965));
    layer1_outputs(4895) <= not((layer0_outputs(488)) or (layer0_outputs(1103)));
    layer1_outputs(4896) <= (layer0_outputs(2310)) and not (layer0_outputs(1447));
    layer1_outputs(4897) <= not(layer0_outputs(2937));
    layer1_outputs(4898) <= '0';
    layer1_outputs(4899) <= (layer0_outputs(5092)) and not (layer0_outputs(4028));
    layer1_outputs(4900) <= not((layer0_outputs(4058)) or (layer0_outputs(1636)));
    layer1_outputs(4901) <= (layer0_outputs(2805)) or (layer0_outputs(4461));
    layer1_outputs(4902) <= (layer0_outputs(1650)) and (layer0_outputs(1489));
    layer1_outputs(4903) <= '1';
    layer1_outputs(4904) <= '0';
    layer1_outputs(4905) <= layer0_outputs(2468);
    layer1_outputs(4906) <= layer0_outputs(2496);
    layer1_outputs(4907) <= '1';
    layer1_outputs(4908) <= not(layer0_outputs(3438)) or (layer0_outputs(714));
    layer1_outputs(4909) <= (layer0_outputs(3948)) and (layer0_outputs(2107));
    layer1_outputs(4910) <= not((layer0_outputs(1612)) and (layer0_outputs(1951)));
    layer1_outputs(4911) <= (layer0_outputs(2022)) and (layer0_outputs(2080));
    layer1_outputs(4912) <= not((layer0_outputs(3042)) or (layer0_outputs(3786)));
    layer1_outputs(4913) <= (layer0_outputs(4774)) or (layer0_outputs(4734));
    layer1_outputs(4914) <= (layer0_outputs(3558)) and not (layer0_outputs(2206));
    layer1_outputs(4915) <= (layer0_outputs(2759)) and not (layer0_outputs(1562));
    layer1_outputs(4916) <= '1';
    layer1_outputs(4917) <= not((layer0_outputs(4746)) and (layer0_outputs(4253)));
    layer1_outputs(4918) <= (layer0_outputs(1096)) or (layer0_outputs(2644));
    layer1_outputs(4919) <= (layer0_outputs(259)) and not (layer0_outputs(1973));
    layer1_outputs(4920) <= (layer0_outputs(1286)) or (layer0_outputs(3147));
    layer1_outputs(4921) <= not((layer0_outputs(2551)) or (layer0_outputs(4027)));
    layer1_outputs(4922) <= layer0_outputs(3332);
    layer1_outputs(4923) <= not(layer0_outputs(3083)) or (layer0_outputs(1808));
    layer1_outputs(4924) <= (layer0_outputs(3422)) and not (layer0_outputs(543));
    layer1_outputs(4925) <= not(layer0_outputs(2000));
    layer1_outputs(4926) <= not((layer0_outputs(3785)) or (layer0_outputs(4252)));
    layer1_outputs(4927) <= '0';
    layer1_outputs(4928) <= not((layer0_outputs(2825)) and (layer0_outputs(2654)));
    layer1_outputs(4929) <= not((layer0_outputs(2657)) and (layer0_outputs(4714)));
    layer1_outputs(4930) <= not(layer0_outputs(2859)) or (layer0_outputs(3592));
    layer1_outputs(4931) <= '1';
    layer1_outputs(4932) <= (layer0_outputs(1311)) or (layer0_outputs(2741));
    layer1_outputs(4933) <= not((layer0_outputs(982)) and (layer0_outputs(1703)));
    layer1_outputs(4934) <= '0';
    layer1_outputs(4935) <= '1';
    layer1_outputs(4936) <= '0';
    layer1_outputs(4937) <= (layer0_outputs(4856)) and not (layer0_outputs(2091));
    layer1_outputs(4938) <= (layer0_outputs(1365)) and not (layer0_outputs(4507));
    layer1_outputs(4939) <= layer0_outputs(4073);
    layer1_outputs(4940) <= '0';
    layer1_outputs(4941) <= layer0_outputs(1016);
    layer1_outputs(4942) <= (layer0_outputs(2839)) and not (layer0_outputs(21));
    layer1_outputs(4943) <= '0';
    layer1_outputs(4944) <= (layer0_outputs(2207)) and not (layer0_outputs(4537));
    layer1_outputs(4945) <= (layer0_outputs(1178)) and (layer0_outputs(740));
    layer1_outputs(4946) <= not(layer0_outputs(1976)) or (layer0_outputs(3385));
    layer1_outputs(4947) <= not(layer0_outputs(1847)) or (layer0_outputs(571));
    layer1_outputs(4948) <= (layer0_outputs(4797)) or (layer0_outputs(5017));
    layer1_outputs(4949) <= not(layer0_outputs(4663));
    layer1_outputs(4950) <= not(layer0_outputs(1367));
    layer1_outputs(4951) <= '1';
    layer1_outputs(4952) <= layer0_outputs(4913);
    layer1_outputs(4953) <= not((layer0_outputs(5005)) and (layer0_outputs(630)));
    layer1_outputs(4954) <= not(layer0_outputs(1969)) or (layer0_outputs(1369));
    layer1_outputs(4955) <= not(layer0_outputs(2078)) or (layer0_outputs(2768));
    layer1_outputs(4956) <= not(layer0_outputs(3307));
    layer1_outputs(4957) <= '0';
    layer1_outputs(4958) <= (layer0_outputs(3069)) and (layer0_outputs(4703));
    layer1_outputs(4959) <= '0';
    layer1_outputs(4960) <= not(layer0_outputs(1977));
    layer1_outputs(4961) <= not((layer0_outputs(1606)) and (layer0_outputs(3765)));
    layer1_outputs(4962) <= not(layer0_outputs(4263));
    layer1_outputs(4963) <= '0';
    layer1_outputs(4964) <= (layer0_outputs(4705)) and not (layer0_outputs(4908));
    layer1_outputs(4965) <= '0';
    layer1_outputs(4966) <= layer0_outputs(2227);
    layer1_outputs(4967) <= layer0_outputs(3497);
    layer1_outputs(4968) <= '0';
    layer1_outputs(4969) <= layer0_outputs(1663);
    layer1_outputs(4970) <= not(layer0_outputs(2431)) or (layer0_outputs(4458));
    layer1_outputs(4971) <= not(layer0_outputs(5100));
    layer1_outputs(4972) <= layer0_outputs(4100);
    layer1_outputs(4973) <= '0';
    layer1_outputs(4974) <= '0';
    layer1_outputs(4975) <= (layer0_outputs(1762)) and (layer0_outputs(1567));
    layer1_outputs(4976) <= (layer0_outputs(2574)) and not (layer0_outputs(3804));
    layer1_outputs(4977) <= (layer0_outputs(1746)) and not (layer0_outputs(3252));
    layer1_outputs(4978) <= (layer0_outputs(2085)) and not (layer0_outputs(1792));
    layer1_outputs(4979) <= not((layer0_outputs(4582)) and (layer0_outputs(763)));
    layer1_outputs(4980) <= not((layer0_outputs(222)) and (layer0_outputs(4812)));
    layer1_outputs(4981) <= not((layer0_outputs(495)) and (layer0_outputs(2372)));
    layer1_outputs(4982) <= (layer0_outputs(3693)) and not (layer0_outputs(2829));
    layer1_outputs(4983) <= not(layer0_outputs(1059));
    layer1_outputs(4984) <= layer0_outputs(4204);
    layer1_outputs(4985) <= (layer0_outputs(1341)) and not (layer0_outputs(1692));
    layer1_outputs(4986) <= '0';
    layer1_outputs(4987) <= layer0_outputs(1727);
    layer1_outputs(4988) <= (layer0_outputs(4115)) and not (layer0_outputs(914));
    layer1_outputs(4989) <= (layer0_outputs(2203)) and not (layer0_outputs(3789));
    layer1_outputs(4990) <= (layer0_outputs(4997)) or (layer0_outputs(933));
    layer1_outputs(4991) <= (layer0_outputs(1826)) and (layer0_outputs(2004));
    layer1_outputs(4992) <= '1';
    layer1_outputs(4993) <= not(layer0_outputs(1918));
    layer1_outputs(4994) <= not((layer0_outputs(700)) or (layer0_outputs(3036)));
    layer1_outputs(4995) <= (layer0_outputs(946)) or (layer0_outputs(1425));
    layer1_outputs(4996) <= not((layer0_outputs(912)) or (layer0_outputs(1916)));
    layer1_outputs(4997) <= not((layer0_outputs(4201)) or (layer0_outputs(501)));
    layer1_outputs(4998) <= (layer0_outputs(1983)) and not (layer0_outputs(783));
    layer1_outputs(4999) <= '0';
    layer1_outputs(5000) <= '1';
    layer1_outputs(5001) <= (layer0_outputs(4523)) or (layer0_outputs(1183));
    layer1_outputs(5002) <= (layer0_outputs(234)) or (layer0_outputs(4078));
    layer1_outputs(5003) <= not(layer0_outputs(246));
    layer1_outputs(5004) <= (layer0_outputs(4850)) or (layer0_outputs(3040));
    layer1_outputs(5005) <= not((layer0_outputs(298)) and (layer0_outputs(3689)));
    layer1_outputs(5006) <= not(layer0_outputs(3595)) or (layer0_outputs(1029));
    layer1_outputs(5007) <= not((layer0_outputs(4760)) or (layer0_outputs(164)));
    layer1_outputs(5008) <= not(layer0_outputs(3263));
    layer1_outputs(5009) <= not(layer0_outputs(4260));
    layer1_outputs(5010) <= layer0_outputs(4307);
    layer1_outputs(5011) <= (layer0_outputs(3682)) and not (layer0_outputs(3356));
    layer1_outputs(5012) <= (layer0_outputs(1359)) xor (layer0_outputs(4588));
    layer1_outputs(5013) <= not(layer0_outputs(948));
    layer1_outputs(5014) <= not(layer0_outputs(4922));
    layer1_outputs(5015) <= (layer0_outputs(1456)) and (layer0_outputs(4080));
    layer1_outputs(5016) <= '1';
    layer1_outputs(5017) <= not(layer0_outputs(2662)) or (layer0_outputs(3539));
    layer1_outputs(5018) <= '0';
    layer1_outputs(5019) <= (layer0_outputs(4086)) and not (layer0_outputs(799));
    layer1_outputs(5020) <= layer0_outputs(3578);
    layer1_outputs(5021) <= layer0_outputs(1408);
    layer1_outputs(5022) <= (layer0_outputs(4411)) and not (layer0_outputs(242));
    layer1_outputs(5023) <= (layer0_outputs(4165)) and (layer0_outputs(4960));
    layer1_outputs(5024) <= '1';
    layer1_outputs(5025) <= not((layer0_outputs(4394)) or (layer0_outputs(4442)));
    layer1_outputs(5026) <= not(layer0_outputs(3590)) or (layer0_outputs(2938));
    layer1_outputs(5027) <= (layer0_outputs(2097)) and (layer0_outputs(4735));
    layer1_outputs(5028) <= '0';
    layer1_outputs(5029) <= '0';
    layer1_outputs(5030) <= '1';
    layer1_outputs(5031) <= layer0_outputs(2055);
    layer1_outputs(5032) <= '1';
    layer1_outputs(5033) <= layer0_outputs(2423);
    layer1_outputs(5034) <= '1';
    layer1_outputs(5035) <= (layer0_outputs(4536)) and not (layer0_outputs(3003));
    layer1_outputs(5036) <= not(layer0_outputs(3734)) or (layer0_outputs(101));
    layer1_outputs(5037) <= layer0_outputs(2050);
    layer1_outputs(5038) <= '1';
    layer1_outputs(5039) <= not(layer0_outputs(2666)) or (layer0_outputs(875));
    layer1_outputs(5040) <= (layer0_outputs(324)) and (layer0_outputs(3068));
    layer1_outputs(5041) <= not(layer0_outputs(4132)) or (layer0_outputs(3589));
    layer1_outputs(5042) <= not((layer0_outputs(4743)) or (layer0_outputs(2861)));
    layer1_outputs(5043) <= layer0_outputs(1018);
    layer1_outputs(5044) <= not((layer0_outputs(2099)) and (layer0_outputs(3364)));
    layer1_outputs(5045) <= not((layer0_outputs(902)) or (layer0_outputs(4289)));
    layer1_outputs(5046) <= not(layer0_outputs(2912)) or (layer0_outputs(908));
    layer1_outputs(5047) <= '0';
    layer1_outputs(5048) <= layer0_outputs(3938);
    layer1_outputs(5049) <= '0';
    layer1_outputs(5050) <= not(layer0_outputs(758));
    layer1_outputs(5051) <= not(layer0_outputs(1337));
    layer1_outputs(5052) <= layer0_outputs(2205);
    layer1_outputs(5053) <= (layer0_outputs(1862)) or (layer0_outputs(750));
    layer1_outputs(5054) <= layer0_outputs(3555);
    layer1_outputs(5055) <= not((layer0_outputs(4648)) or (layer0_outputs(2361)));
    layer1_outputs(5056) <= '1';
    layer1_outputs(5057) <= layer0_outputs(4514);
    layer1_outputs(5058) <= not((layer0_outputs(3947)) and (layer0_outputs(2978)));
    layer1_outputs(5059) <= '1';
    layer1_outputs(5060) <= not(layer0_outputs(5119));
    layer1_outputs(5061) <= layer0_outputs(3650);
    layer1_outputs(5062) <= (layer0_outputs(1310)) or (layer0_outputs(5059));
    layer1_outputs(5063) <= '1';
    layer1_outputs(5064) <= not((layer0_outputs(3052)) or (layer0_outputs(2315)));
    layer1_outputs(5065) <= not(layer0_outputs(319)) or (layer0_outputs(2867));
    layer1_outputs(5066) <= (layer0_outputs(3303)) or (layer0_outputs(3683));
    layer1_outputs(5067) <= not(layer0_outputs(862)) or (layer0_outputs(1854));
    layer1_outputs(5068) <= (layer0_outputs(2071)) or (layer0_outputs(4008));
    layer1_outputs(5069) <= not((layer0_outputs(3587)) and (layer0_outputs(5018)));
    layer1_outputs(5070) <= (layer0_outputs(4811)) and not (layer0_outputs(4157));
    layer1_outputs(5071) <= (layer0_outputs(2480)) or (layer0_outputs(1638));
    layer1_outputs(5072) <= not(layer0_outputs(1990)) or (layer0_outputs(1446));
    layer1_outputs(5073) <= not(layer0_outputs(887));
    layer1_outputs(5074) <= '1';
    layer1_outputs(5075) <= not((layer0_outputs(3762)) or (layer0_outputs(3291)));
    layer1_outputs(5076) <= (layer0_outputs(4439)) and not (layer0_outputs(3111));
    layer1_outputs(5077) <= '1';
    layer1_outputs(5078) <= '0';
    layer1_outputs(5079) <= not((layer0_outputs(2673)) or (layer0_outputs(1183)));
    layer1_outputs(5080) <= not((layer0_outputs(2339)) or (layer0_outputs(3780)));
    layer1_outputs(5081) <= not(layer0_outputs(3769)) or (layer0_outputs(4347));
    layer1_outputs(5082) <= '1';
    layer1_outputs(5083) <= layer0_outputs(2347);
    layer1_outputs(5084) <= '1';
    layer1_outputs(5085) <= not((layer0_outputs(4779)) or (layer0_outputs(280)));
    layer1_outputs(5086) <= not(layer0_outputs(3081)) or (layer0_outputs(1083));
    layer1_outputs(5087) <= (layer0_outputs(2116)) and (layer0_outputs(272));
    layer1_outputs(5088) <= (layer0_outputs(4221)) or (layer0_outputs(3859));
    layer1_outputs(5089) <= (layer0_outputs(3662)) and not (layer0_outputs(5007));
    layer1_outputs(5090) <= '1';
    layer1_outputs(5091) <= not((layer0_outputs(3058)) or (layer0_outputs(2541)));
    layer1_outputs(5092) <= (layer0_outputs(4613)) or (layer0_outputs(4186));
    layer1_outputs(5093) <= not((layer0_outputs(1959)) or (layer0_outputs(3593)));
    layer1_outputs(5094) <= '1';
    layer1_outputs(5095) <= layer0_outputs(2304);
    layer1_outputs(5096) <= '0';
    layer1_outputs(5097) <= (layer0_outputs(1350)) and not (layer0_outputs(3543));
    layer1_outputs(5098) <= layer0_outputs(2401);
    layer1_outputs(5099) <= (layer0_outputs(709)) and not (layer0_outputs(256));
    layer1_outputs(5100) <= '1';
    layer1_outputs(5101) <= '0';
    layer1_outputs(5102) <= layer0_outputs(1627);
    layer1_outputs(5103) <= '0';
    layer1_outputs(5104) <= '1';
    layer1_outputs(5105) <= '0';
    layer1_outputs(5106) <= not(layer0_outputs(1422)) or (layer0_outputs(2980));
    layer1_outputs(5107) <= layer0_outputs(2178);
    layer1_outputs(5108) <= '0';
    layer1_outputs(5109) <= (layer0_outputs(95)) and not (layer0_outputs(2766));
    layer1_outputs(5110) <= not(layer0_outputs(3311)) or (layer0_outputs(2956));
    layer1_outputs(5111) <= not((layer0_outputs(3053)) and (layer0_outputs(239)));
    layer1_outputs(5112) <= '1';
    layer1_outputs(5113) <= layer0_outputs(2907);
    layer1_outputs(5114) <= not(layer0_outputs(1224));
    layer1_outputs(5115) <= not(layer0_outputs(1817));
    layer1_outputs(5116) <= '1';
    layer1_outputs(5117) <= not(layer0_outputs(1731)) or (layer0_outputs(3779));
    layer1_outputs(5118) <= layer0_outputs(3864);
    layer1_outputs(5119) <= not(layer0_outputs(1641));
    layer2_outputs(0) <= (layer1_outputs(4628)) and not (layer1_outputs(3490));
    layer2_outputs(1) <= not(layer1_outputs(2296)) or (layer1_outputs(4041));
    layer2_outputs(2) <= not(layer1_outputs(4292));
    layer2_outputs(3) <= layer1_outputs(196);
    layer2_outputs(4) <= (layer1_outputs(497)) or (layer1_outputs(3521));
    layer2_outputs(5) <= '0';
    layer2_outputs(6) <= not(layer1_outputs(2073));
    layer2_outputs(7) <= layer1_outputs(1190);
    layer2_outputs(8) <= (layer1_outputs(2921)) and not (layer1_outputs(771));
    layer2_outputs(9) <= '1';
    layer2_outputs(10) <= not((layer1_outputs(2062)) or (layer1_outputs(3600)));
    layer2_outputs(11) <= (layer1_outputs(529)) xor (layer1_outputs(131));
    layer2_outputs(12) <= not(layer1_outputs(1994)) or (layer1_outputs(486));
    layer2_outputs(13) <= layer1_outputs(374);
    layer2_outputs(14) <= '1';
    layer2_outputs(15) <= not(layer1_outputs(3451)) or (layer1_outputs(4961));
    layer2_outputs(16) <= (layer1_outputs(397)) or (layer1_outputs(4516));
    layer2_outputs(17) <= layer1_outputs(3008);
    layer2_outputs(18) <= '0';
    layer2_outputs(19) <= not(layer1_outputs(371)) or (layer1_outputs(2788));
    layer2_outputs(20) <= '0';
    layer2_outputs(21) <= not(layer1_outputs(2286));
    layer2_outputs(22) <= not((layer1_outputs(336)) xor (layer1_outputs(3875)));
    layer2_outputs(23) <= not((layer1_outputs(2068)) and (layer1_outputs(685)));
    layer2_outputs(24) <= not((layer1_outputs(3589)) and (layer1_outputs(1198)));
    layer2_outputs(25) <= '1';
    layer2_outputs(26) <= not(layer1_outputs(887)) or (layer1_outputs(1585));
    layer2_outputs(27) <= '0';
    layer2_outputs(28) <= not(layer1_outputs(1163)) or (layer1_outputs(1456));
    layer2_outputs(29) <= not((layer1_outputs(4056)) or (layer1_outputs(581)));
    layer2_outputs(30) <= not((layer1_outputs(4015)) and (layer1_outputs(776)));
    layer2_outputs(31) <= (layer1_outputs(1754)) and (layer1_outputs(4034));
    layer2_outputs(32) <= (layer1_outputs(1934)) and (layer1_outputs(2614));
    layer2_outputs(33) <= not(layer1_outputs(3987));
    layer2_outputs(34) <= not(layer1_outputs(2709));
    layer2_outputs(35) <= '0';
    layer2_outputs(36) <= not(layer1_outputs(261)) or (layer1_outputs(4318));
    layer2_outputs(37) <= (layer1_outputs(1467)) or (layer1_outputs(4548));
    layer2_outputs(38) <= layer1_outputs(94);
    layer2_outputs(39) <= (layer1_outputs(1737)) and not (layer1_outputs(2671));
    layer2_outputs(40) <= '1';
    layer2_outputs(41) <= layer1_outputs(920);
    layer2_outputs(42) <= (layer1_outputs(5099)) and not (layer1_outputs(4411));
    layer2_outputs(43) <= not(layer1_outputs(205));
    layer2_outputs(44) <= not(layer1_outputs(4882)) or (layer1_outputs(661));
    layer2_outputs(45) <= '1';
    layer2_outputs(46) <= not(layer1_outputs(3977)) or (layer1_outputs(2630));
    layer2_outputs(47) <= (layer1_outputs(3532)) and (layer1_outputs(3733));
    layer2_outputs(48) <= layer1_outputs(1091);
    layer2_outputs(49) <= (layer1_outputs(3469)) and not (layer1_outputs(4671));
    layer2_outputs(50) <= (layer1_outputs(3390)) and not (layer1_outputs(4756));
    layer2_outputs(51) <= '0';
    layer2_outputs(52) <= (layer1_outputs(2614)) and not (layer1_outputs(1547));
    layer2_outputs(53) <= not(layer1_outputs(4148)) or (layer1_outputs(4447));
    layer2_outputs(54) <= (layer1_outputs(4749)) and not (layer1_outputs(1332));
    layer2_outputs(55) <= not(layer1_outputs(2155));
    layer2_outputs(56) <= (layer1_outputs(4131)) and not (layer1_outputs(771));
    layer2_outputs(57) <= not(layer1_outputs(4123)) or (layer1_outputs(3611));
    layer2_outputs(58) <= '1';
    layer2_outputs(59) <= not((layer1_outputs(3177)) and (layer1_outputs(2279)));
    layer2_outputs(60) <= not(layer1_outputs(3116));
    layer2_outputs(61) <= not((layer1_outputs(3990)) and (layer1_outputs(901)));
    layer2_outputs(62) <= not((layer1_outputs(1826)) or (layer1_outputs(129)));
    layer2_outputs(63) <= (layer1_outputs(2740)) and not (layer1_outputs(3328));
    layer2_outputs(64) <= not((layer1_outputs(168)) xor (layer1_outputs(1491)));
    layer2_outputs(65) <= layer1_outputs(3675);
    layer2_outputs(66) <= '0';
    layer2_outputs(67) <= (layer1_outputs(2991)) or (layer1_outputs(1739));
    layer2_outputs(68) <= not(layer1_outputs(3536)) or (layer1_outputs(4235));
    layer2_outputs(69) <= not(layer1_outputs(2227)) or (layer1_outputs(1459));
    layer2_outputs(70) <= (layer1_outputs(3533)) xor (layer1_outputs(1153));
    layer2_outputs(71) <= '1';
    layer2_outputs(72) <= layer1_outputs(210);
    layer2_outputs(73) <= (layer1_outputs(2611)) and not (layer1_outputs(397));
    layer2_outputs(74) <= not(layer1_outputs(1249)) or (layer1_outputs(2311));
    layer2_outputs(75) <= (layer1_outputs(4133)) or (layer1_outputs(1114));
    layer2_outputs(76) <= '0';
    layer2_outputs(77) <= '1';
    layer2_outputs(78) <= not(layer1_outputs(2741));
    layer2_outputs(79) <= '1';
    layer2_outputs(80) <= layer1_outputs(4851);
    layer2_outputs(81) <= not(layer1_outputs(4367)) or (layer1_outputs(4297));
    layer2_outputs(82) <= not((layer1_outputs(153)) or (layer1_outputs(3341)));
    layer2_outputs(83) <= not((layer1_outputs(598)) xor (layer1_outputs(4519)));
    layer2_outputs(84) <= not(layer1_outputs(2816)) or (layer1_outputs(2082));
    layer2_outputs(85) <= '1';
    layer2_outputs(86) <= not((layer1_outputs(1863)) or (layer1_outputs(2704)));
    layer2_outputs(87) <= '1';
    layer2_outputs(88) <= not((layer1_outputs(3816)) xor (layer1_outputs(4693)));
    layer2_outputs(89) <= not(layer1_outputs(2005));
    layer2_outputs(90) <= (layer1_outputs(3445)) or (layer1_outputs(3572));
    layer2_outputs(91) <= '0';
    layer2_outputs(92) <= not((layer1_outputs(4891)) and (layer1_outputs(3079)));
    layer2_outputs(93) <= (layer1_outputs(4363)) and (layer1_outputs(927));
    layer2_outputs(94) <= not(layer1_outputs(1893)) or (layer1_outputs(394));
    layer2_outputs(95) <= (layer1_outputs(778)) or (layer1_outputs(3869));
    layer2_outputs(96) <= '1';
    layer2_outputs(97) <= (layer1_outputs(4808)) and (layer1_outputs(3061));
    layer2_outputs(98) <= (layer1_outputs(844)) xor (layer1_outputs(1806));
    layer2_outputs(99) <= (layer1_outputs(4217)) and not (layer1_outputs(2884));
    layer2_outputs(100) <= (layer1_outputs(1897)) and not (layer1_outputs(1935));
    layer2_outputs(101) <= (layer1_outputs(3177)) and (layer1_outputs(210));
    layer2_outputs(102) <= '0';
    layer2_outputs(103) <= layer1_outputs(856);
    layer2_outputs(104) <= layer1_outputs(4397);
    layer2_outputs(105) <= (layer1_outputs(1169)) and (layer1_outputs(812));
    layer2_outputs(106) <= '0';
    layer2_outputs(107) <= (layer1_outputs(2095)) and not (layer1_outputs(1820));
    layer2_outputs(108) <= not((layer1_outputs(4841)) or (layer1_outputs(1653)));
    layer2_outputs(109) <= not(layer1_outputs(3041)) or (layer1_outputs(476));
    layer2_outputs(110) <= layer1_outputs(3254);
    layer2_outputs(111) <= not((layer1_outputs(1397)) or (layer1_outputs(1395)));
    layer2_outputs(112) <= '0';
    layer2_outputs(113) <= '1';
    layer2_outputs(114) <= (layer1_outputs(4743)) or (layer1_outputs(5036));
    layer2_outputs(115) <= not(layer1_outputs(4135)) or (layer1_outputs(2754));
    layer2_outputs(116) <= layer1_outputs(1302);
    layer2_outputs(117) <= '1';
    layer2_outputs(118) <= not(layer1_outputs(1327)) or (layer1_outputs(5044));
    layer2_outputs(119) <= '0';
    layer2_outputs(120) <= (layer1_outputs(4017)) and not (layer1_outputs(1229));
    layer2_outputs(121) <= not((layer1_outputs(1486)) and (layer1_outputs(456)));
    layer2_outputs(122) <= layer1_outputs(4293);
    layer2_outputs(123) <= (layer1_outputs(2863)) and not (layer1_outputs(452));
    layer2_outputs(124) <= not(layer1_outputs(2195)) or (layer1_outputs(3257));
    layer2_outputs(125) <= not(layer1_outputs(3478));
    layer2_outputs(126) <= layer1_outputs(2274);
    layer2_outputs(127) <= not(layer1_outputs(737)) or (layer1_outputs(1252));
    layer2_outputs(128) <= '0';
    layer2_outputs(129) <= not(layer1_outputs(3459));
    layer2_outputs(130) <= '0';
    layer2_outputs(131) <= not(layer1_outputs(2359));
    layer2_outputs(132) <= (layer1_outputs(3887)) and not (layer1_outputs(2893));
    layer2_outputs(133) <= layer1_outputs(1011);
    layer2_outputs(134) <= not(layer1_outputs(2350)) or (layer1_outputs(3738));
    layer2_outputs(135) <= (layer1_outputs(2363)) and not (layer1_outputs(2320));
    layer2_outputs(136) <= (layer1_outputs(2515)) and (layer1_outputs(353));
    layer2_outputs(137) <= not(layer1_outputs(2447));
    layer2_outputs(138) <= not(layer1_outputs(4836));
    layer2_outputs(139) <= not((layer1_outputs(1138)) or (layer1_outputs(1454)));
    layer2_outputs(140) <= '0';
    layer2_outputs(141) <= not(layer1_outputs(418)) or (layer1_outputs(2227));
    layer2_outputs(142) <= (layer1_outputs(1357)) or (layer1_outputs(1063));
    layer2_outputs(143) <= not(layer1_outputs(1388));
    layer2_outputs(144) <= not(layer1_outputs(675));
    layer2_outputs(145) <= not(layer1_outputs(2441));
    layer2_outputs(146) <= '1';
    layer2_outputs(147) <= '1';
    layer2_outputs(148) <= (layer1_outputs(480)) and (layer1_outputs(2733));
    layer2_outputs(149) <= '0';
    layer2_outputs(150) <= '1';
    layer2_outputs(151) <= '0';
    layer2_outputs(152) <= '0';
    layer2_outputs(153) <= (layer1_outputs(2468)) and (layer1_outputs(4029));
    layer2_outputs(154) <= '0';
    layer2_outputs(155) <= not(layer1_outputs(3573));
    layer2_outputs(156) <= not(layer1_outputs(4213));
    layer2_outputs(157) <= (layer1_outputs(2675)) and (layer1_outputs(3318));
    layer2_outputs(158) <= '1';
    layer2_outputs(159) <= layer1_outputs(2315);
    layer2_outputs(160) <= (layer1_outputs(1270)) and (layer1_outputs(2648));
    layer2_outputs(161) <= (layer1_outputs(4342)) and not (layer1_outputs(2875));
    layer2_outputs(162) <= (layer1_outputs(3404)) and not (layer1_outputs(4930));
    layer2_outputs(163) <= (layer1_outputs(3016)) and not (layer1_outputs(1214));
    layer2_outputs(164) <= '0';
    layer2_outputs(165) <= (layer1_outputs(3231)) and (layer1_outputs(4923));
    layer2_outputs(166) <= '0';
    layer2_outputs(167) <= not(layer1_outputs(1976));
    layer2_outputs(168) <= not(layer1_outputs(4533));
    layer2_outputs(169) <= not((layer1_outputs(513)) or (layer1_outputs(3679)));
    layer2_outputs(170) <= not(layer1_outputs(81)) or (layer1_outputs(1939));
    layer2_outputs(171) <= (layer1_outputs(4984)) or (layer1_outputs(1370));
    layer2_outputs(172) <= layer1_outputs(1278);
    layer2_outputs(173) <= not((layer1_outputs(628)) or (layer1_outputs(4504)));
    layer2_outputs(174) <= '0';
    layer2_outputs(175) <= (layer1_outputs(3464)) and not (layer1_outputs(1909));
    layer2_outputs(176) <= not(layer1_outputs(404));
    layer2_outputs(177) <= not(layer1_outputs(331)) or (layer1_outputs(14));
    layer2_outputs(178) <= not((layer1_outputs(2027)) or (layer1_outputs(285)));
    layer2_outputs(179) <= layer1_outputs(4384);
    layer2_outputs(180) <= not(layer1_outputs(3078)) or (layer1_outputs(469));
    layer2_outputs(181) <= layer1_outputs(3637);
    layer2_outputs(182) <= not(layer1_outputs(906));
    layer2_outputs(183) <= not(layer1_outputs(813)) or (layer1_outputs(793));
    layer2_outputs(184) <= layer1_outputs(2293);
    layer2_outputs(185) <= '1';
    layer2_outputs(186) <= not(layer1_outputs(3843));
    layer2_outputs(187) <= layer1_outputs(1343);
    layer2_outputs(188) <= layer1_outputs(734);
    layer2_outputs(189) <= '1';
    layer2_outputs(190) <= not(layer1_outputs(3573)) or (layer1_outputs(2764));
    layer2_outputs(191) <= '1';
    layer2_outputs(192) <= not(layer1_outputs(3718)) or (layer1_outputs(4347));
    layer2_outputs(193) <= '1';
    layer2_outputs(194) <= (layer1_outputs(4190)) and not (layer1_outputs(3000));
    layer2_outputs(195) <= not(layer1_outputs(887)) or (layer1_outputs(1587));
    layer2_outputs(196) <= '1';
    layer2_outputs(197) <= '0';
    layer2_outputs(198) <= not((layer1_outputs(1431)) or (layer1_outputs(3027)));
    layer2_outputs(199) <= not(layer1_outputs(2119));
    layer2_outputs(200) <= '0';
    layer2_outputs(201) <= layer1_outputs(291);
    layer2_outputs(202) <= not((layer1_outputs(2701)) or (layer1_outputs(4893)));
    layer2_outputs(203) <= '0';
    layer2_outputs(204) <= not(layer1_outputs(302)) or (layer1_outputs(4830));
    layer2_outputs(205) <= '0';
    layer2_outputs(206) <= not(layer1_outputs(858)) or (layer1_outputs(3828));
    layer2_outputs(207) <= (layer1_outputs(4978)) and not (layer1_outputs(2886));
    layer2_outputs(208) <= (layer1_outputs(2233)) and (layer1_outputs(881));
    layer2_outputs(209) <= (layer1_outputs(2259)) and (layer1_outputs(4950));
    layer2_outputs(210) <= not(layer1_outputs(932)) or (layer1_outputs(4955));
    layer2_outputs(211) <= '0';
    layer2_outputs(212) <= layer1_outputs(2900);
    layer2_outputs(213) <= not(layer1_outputs(2035)) or (layer1_outputs(3727));
    layer2_outputs(214) <= not(layer1_outputs(3441)) or (layer1_outputs(1990));
    layer2_outputs(215) <= not((layer1_outputs(3332)) and (layer1_outputs(43)));
    layer2_outputs(216) <= (layer1_outputs(4702)) or (layer1_outputs(2640));
    layer2_outputs(217) <= '1';
    layer2_outputs(218) <= (layer1_outputs(1053)) or (layer1_outputs(4992));
    layer2_outputs(219) <= not(layer1_outputs(2004)) or (layer1_outputs(593));
    layer2_outputs(220) <= (layer1_outputs(4449)) or (layer1_outputs(1140));
    layer2_outputs(221) <= '1';
    layer2_outputs(222) <= not(layer1_outputs(3045)) or (layer1_outputs(3928));
    layer2_outputs(223) <= '0';
    layer2_outputs(224) <= '1';
    layer2_outputs(225) <= layer1_outputs(1633);
    layer2_outputs(226) <= not(layer1_outputs(4985)) or (layer1_outputs(238));
    layer2_outputs(227) <= not(layer1_outputs(3895));
    layer2_outputs(228) <= not(layer1_outputs(4146)) or (layer1_outputs(3944));
    layer2_outputs(229) <= not(layer1_outputs(3269)) or (layer1_outputs(2178));
    layer2_outputs(230) <= '0';
    layer2_outputs(231) <= '0';
    layer2_outputs(232) <= (layer1_outputs(3031)) or (layer1_outputs(3379));
    layer2_outputs(233) <= '0';
    layer2_outputs(234) <= '0';
    layer2_outputs(235) <= (layer1_outputs(4674)) and (layer1_outputs(4069));
    layer2_outputs(236) <= layer1_outputs(1719);
    layer2_outputs(237) <= not((layer1_outputs(791)) and (layer1_outputs(2843)));
    layer2_outputs(238) <= (layer1_outputs(4296)) or (layer1_outputs(4099));
    layer2_outputs(239) <= '0';
    layer2_outputs(240) <= (layer1_outputs(3731)) and (layer1_outputs(933));
    layer2_outputs(241) <= '1';
    layer2_outputs(242) <= not(layer1_outputs(4479)) or (layer1_outputs(1454));
    layer2_outputs(243) <= not((layer1_outputs(3656)) or (layer1_outputs(4216)));
    layer2_outputs(244) <= not(layer1_outputs(5057));
    layer2_outputs(245) <= '1';
    layer2_outputs(246) <= '0';
    layer2_outputs(247) <= layer1_outputs(1527);
    layer2_outputs(248) <= not(layer1_outputs(3715)) or (layer1_outputs(4846));
    layer2_outputs(249) <= not(layer1_outputs(1360));
    layer2_outputs(250) <= '0';
    layer2_outputs(251) <= layer1_outputs(3437);
    layer2_outputs(252) <= not(layer1_outputs(4591));
    layer2_outputs(253) <= '1';
    layer2_outputs(254) <= '0';
    layer2_outputs(255) <= not(layer1_outputs(3593));
    layer2_outputs(256) <= (layer1_outputs(2183)) and not (layer1_outputs(4805));
    layer2_outputs(257) <= not(layer1_outputs(1548));
    layer2_outputs(258) <= not(layer1_outputs(4762)) or (layer1_outputs(823));
    layer2_outputs(259) <= '0';
    layer2_outputs(260) <= (layer1_outputs(4070)) and (layer1_outputs(4090));
    layer2_outputs(261) <= not(layer1_outputs(1375)) or (layer1_outputs(1913));
    layer2_outputs(262) <= not(layer1_outputs(2757));
    layer2_outputs(263) <= not(layer1_outputs(4357));
    layer2_outputs(264) <= layer1_outputs(5075);
    layer2_outputs(265) <= '0';
    layer2_outputs(266) <= layer1_outputs(656);
    layer2_outputs(267) <= '0';
    layer2_outputs(268) <= layer1_outputs(3330);
    layer2_outputs(269) <= layer1_outputs(5003);
    layer2_outputs(270) <= '1';
    layer2_outputs(271) <= layer1_outputs(317);
    layer2_outputs(272) <= not(layer1_outputs(1560));
    layer2_outputs(273) <= not((layer1_outputs(1024)) and (layer1_outputs(196)));
    layer2_outputs(274) <= (layer1_outputs(461)) and (layer1_outputs(2407));
    layer2_outputs(275) <= (layer1_outputs(142)) or (layer1_outputs(897));
    layer2_outputs(276) <= '1';
    layer2_outputs(277) <= '1';
    layer2_outputs(278) <= not(layer1_outputs(1635));
    layer2_outputs(279) <= not((layer1_outputs(581)) or (layer1_outputs(4557)));
    layer2_outputs(280) <= not(layer1_outputs(4243));
    layer2_outputs(281) <= (layer1_outputs(3539)) and not (layer1_outputs(1964));
    layer2_outputs(282) <= layer1_outputs(1416);
    layer2_outputs(283) <= not(layer1_outputs(3054));
    layer2_outputs(284) <= not((layer1_outputs(641)) and (layer1_outputs(2665)));
    layer2_outputs(285) <= not((layer1_outputs(431)) or (layer1_outputs(4228)));
    layer2_outputs(286) <= (layer1_outputs(1569)) or (layer1_outputs(329));
    layer2_outputs(287) <= not(layer1_outputs(4279)) or (layer1_outputs(998));
    layer2_outputs(288) <= layer1_outputs(3513);
    layer2_outputs(289) <= not((layer1_outputs(727)) or (layer1_outputs(1129)));
    layer2_outputs(290) <= not(layer1_outputs(3810));
    layer2_outputs(291) <= not(layer1_outputs(1943));
    layer2_outputs(292) <= not(layer1_outputs(2080)) or (layer1_outputs(483));
    layer2_outputs(293) <= layer1_outputs(944);
    layer2_outputs(294) <= not(layer1_outputs(5053));
    layer2_outputs(295) <= (layer1_outputs(703)) and not (layer1_outputs(4286));
    layer2_outputs(296) <= (layer1_outputs(4773)) or (layer1_outputs(2805));
    layer2_outputs(297) <= '1';
    layer2_outputs(298) <= not((layer1_outputs(4844)) or (layer1_outputs(4532)));
    layer2_outputs(299) <= (layer1_outputs(3717)) and not (layer1_outputs(4634));
    layer2_outputs(300) <= (layer1_outputs(4038)) xor (layer1_outputs(3788));
    layer2_outputs(301) <= '1';
    layer2_outputs(302) <= (layer1_outputs(2039)) and (layer1_outputs(1885));
    layer2_outputs(303) <= not(layer1_outputs(5116));
    layer2_outputs(304) <= not(layer1_outputs(1199)) or (layer1_outputs(2851));
    layer2_outputs(305) <= not(layer1_outputs(4510)) or (layer1_outputs(3120));
    layer2_outputs(306) <= not(layer1_outputs(403));
    layer2_outputs(307) <= (layer1_outputs(3162)) and not (layer1_outputs(1459));
    layer2_outputs(308) <= not(layer1_outputs(233));
    layer2_outputs(309) <= not(layer1_outputs(1526));
    layer2_outputs(310) <= (layer1_outputs(2037)) and (layer1_outputs(2125));
    layer2_outputs(311) <= not((layer1_outputs(86)) or (layer1_outputs(1540)));
    layer2_outputs(312) <= (layer1_outputs(5085)) and (layer1_outputs(2149));
    layer2_outputs(313) <= (layer1_outputs(484)) and (layer1_outputs(1594));
    layer2_outputs(314) <= (layer1_outputs(761)) xor (layer1_outputs(3032));
    layer2_outputs(315) <= not((layer1_outputs(2270)) or (layer1_outputs(3594)));
    layer2_outputs(316) <= (layer1_outputs(4700)) and (layer1_outputs(4873));
    layer2_outputs(317) <= '1';
    layer2_outputs(318) <= (layer1_outputs(374)) or (layer1_outputs(2461));
    layer2_outputs(319) <= layer1_outputs(3893);
    layer2_outputs(320) <= not(layer1_outputs(1965)) or (layer1_outputs(2019));
    layer2_outputs(321) <= not((layer1_outputs(4229)) or (layer1_outputs(1017)));
    layer2_outputs(322) <= (layer1_outputs(2169)) and not (layer1_outputs(90));
    layer2_outputs(323) <= (layer1_outputs(2414)) and (layer1_outputs(3853));
    layer2_outputs(324) <= (layer1_outputs(4734)) or (layer1_outputs(1060));
    layer2_outputs(325) <= not((layer1_outputs(2057)) and (layer1_outputs(3139)));
    layer2_outputs(326) <= not(layer1_outputs(2620));
    layer2_outputs(327) <= (layer1_outputs(4959)) and not (layer1_outputs(2361));
    layer2_outputs(328) <= layer1_outputs(4947);
    layer2_outputs(329) <= not(layer1_outputs(969)) or (layer1_outputs(2755));
    layer2_outputs(330) <= '1';
    layer2_outputs(331) <= (layer1_outputs(2206)) and not (layer1_outputs(701));
    layer2_outputs(332) <= (layer1_outputs(1349)) and not (layer1_outputs(3258));
    layer2_outputs(333) <= layer1_outputs(4205);
    layer2_outputs(334) <= layer1_outputs(173);
    layer2_outputs(335) <= '1';
    layer2_outputs(336) <= not(layer1_outputs(270));
    layer2_outputs(337) <= '1';
    layer2_outputs(338) <= '0';
    layer2_outputs(339) <= layer1_outputs(3304);
    layer2_outputs(340) <= layer1_outputs(222);
    layer2_outputs(341) <= not((layer1_outputs(4684)) or (layer1_outputs(1340)));
    layer2_outputs(342) <= '0';
    layer2_outputs(343) <= not(layer1_outputs(5068));
    layer2_outputs(344) <= layer1_outputs(2643);
    layer2_outputs(345) <= layer1_outputs(3669);
    layer2_outputs(346) <= layer1_outputs(1305);
    layer2_outputs(347) <= not((layer1_outputs(229)) and (layer1_outputs(4514)));
    layer2_outputs(348) <= (layer1_outputs(3105)) and not (layer1_outputs(4013));
    layer2_outputs(349) <= layer1_outputs(1714);
    layer2_outputs(350) <= '1';
    layer2_outputs(351) <= not((layer1_outputs(3313)) or (layer1_outputs(3710)));
    layer2_outputs(352) <= '1';
    layer2_outputs(353) <= not(layer1_outputs(1230));
    layer2_outputs(354) <= not(layer1_outputs(133)) or (layer1_outputs(67));
    layer2_outputs(355) <= (layer1_outputs(1712)) and not (layer1_outputs(2908));
    layer2_outputs(356) <= not(layer1_outputs(4461)) or (layer1_outputs(2427));
    layer2_outputs(357) <= '1';
    layer2_outputs(358) <= layer1_outputs(641);
    layer2_outputs(359) <= (layer1_outputs(1210)) and (layer1_outputs(716));
    layer2_outputs(360) <= not(layer1_outputs(3159)) or (layer1_outputs(4436));
    layer2_outputs(361) <= not((layer1_outputs(747)) or (layer1_outputs(1947)));
    layer2_outputs(362) <= layer1_outputs(1736);
    layer2_outputs(363) <= '1';
    layer2_outputs(364) <= (layer1_outputs(4301)) and not (layer1_outputs(2241));
    layer2_outputs(365) <= not((layer1_outputs(3943)) or (layer1_outputs(450)));
    layer2_outputs(366) <= (layer1_outputs(4220)) and not (layer1_outputs(2927));
    layer2_outputs(367) <= layer1_outputs(118);
    layer2_outputs(368) <= '1';
    layer2_outputs(369) <= layer1_outputs(563);
    layer2_outputs(370) <= layer1_outputs(1118);
    layer2_outputs(371) <= not((layer1_outputs(2120)) and (layer1_outputs(1553)));
    layer2_outputs(372) <= (layer1_outputs(2260)) and not (layer1_outputs(2767));
    layer2_outputs(373) <= not(layer1_outputs(4410));
    layer2_outputs(374) <= (layer1_outputs(2620)) and not (layer1_outputs(905));
    layer2_outputs(375) <= not((layer1_outputs(733)) and (layer1_outputs(4497)));
    layer2_outputs(376) <= '0';
    layer2_outputs(377) <= (layer1_outputs(1529)) and not (layer1_outputs(1785));
    layer2_outputs(378) <= (layer1_outputs(271)) and not (layer1_outputs(186));
    layer2_outputs(379) <= '0';
    layer2_outputs(380) <= (layer1_outputs(2992)) or (layer1_outputs(2841));
    layer2_outputs(381) <= '0';
    layer2_outputs(382) <= not(layer1_outputs(3235));
    layer2_outputs(383) <= not(layer1_outputs(4857));
    layer2_outputs(384) <= layer1_outputs(4348);
    layer2_outputs(385) <= '1';
    layer2_outputs(386) <= not(layer1_outputs(3746));
    layer2_outputs(387) <= (layer1_outputs(1538)) and (layer1_outputs(3053));
    layer2_outputs(388) <= not((layer1_outputs(218)) or (layer1_outputs(2432)));
    layer2_outputs(389) <= '1';
    layer2_outputs(390) <= (layer1_outputs(3296)) and (layer1_outputs(4965));
    layer2_outputs(391) <= not((layer1_outputs(1629)) and (layer1_outputs(518)));
    layer2_outputs(392) <= not(layer1_outputs(2327)) or (layer1_outputs(470));
    layer2_outputs(393) <= (layer1_outputs(189)) and (layer1_outputs(3795));
    layer2_outputs(394) <= not(layer1_outputs(2217));
    layer2_outputs(395) <= not((layer1_outputs(539)) or (layer1_outputs(2670)));
    layer2_outputs(396) <= not((layer1_outputs(3212)) and (layer1_outputs(554)));
    layer2_outputs(397) <= '0';
    layer2_outputs(398) <= '0';
    layer2_outputs(399) <= (layer1_outputs(2122)) and not (layer1_outputs(3178));
    layer2_outputs(400) <= not(layer1_outputs(2667)) or (layer1_outputs(1643));
    layer2_outputs(401) <= not(layer1_outputs(4139));
    layer2_outputs(402) <= '0';
    layer2_outputs(403) <= layer1_outputs(1890);
    layer2_outputs(404) <= not(layer1_outputs(2954));
    layer2_outputs(405) <= not((layer1_outputs(540)) and (layer1_outputs(82)));
    layer2_outputs(406) <= (layer1_outputs(4223)) and (layer1_outputs(4189));
    layer2_outputs(407) <= (layer1_outputs(1578)) or (layer1_outputs(4408));
    layer2_outputs(408) <= (layer1_outputs(3641)) and (layer1_outputs(3808));
    layer2_outputs(409) <= not(layer1_outputs(2864)) or (layer1_outputs(5016));
    layer2_outputs(410) <= not((layer1_outputs(3462)) or (layer1_outputs(1988)));
    layer2_outputs(411) <= not(layer1_outputs(2469));
    layer2_outputs(412) <= layer1_outputs(1892);
    layer2_outputs(413) <= not(layer1_outputs(3779)) or (layer1_outputs(2762));
    layer2_outputs(414) <= layer1_outputs(888);
    layer2_outputs(415) <= not(layer1_outputs(1616)) or (layer1_outputs(596));
    layer2_outputs(416) <= not((layer1_outputs(125)) and (layer1_outputs(4631)));
    layer2_outputs(417) <= (layer1_outputs(941)) and (layer1_outputs(1713));
    layer2_outputs(418) <= (layer1_outputs(2662)) and not (layer1_outputs(4707));
    layer2_outputs(419) <= '0';
    layer2_outputs(420) <= not((layer1_outputs(4484)) and (layer1_outputs(2245)));
    layer2_outputs(421) <= (layer1_outputs(3554)) and not (layer1_outputs(1743));
    layer2_outputs(422) <= '1';
    layer2_outputs(423) <= (layer1_outputs(4455)) and (layer1_outputs(3767));
    layer2_outputs(424) <= not((layer1_outputs(5003)) and (layer1_outputs(1656)));
    layer2_outputs(425) <= not((layer1_outputs(413)) or (layer1_outputs(2627)));
    layer2_outputs(426) <= not(layer1_outputs(854));
    layer2_outputs(427) <= (layer1_outputs(3862)) or (layer1_outputs(3556));
    layer2_outputs(428) <= not(layer1_outputs(59)) or (layer1_outputs(2196));
    layer2_outputs(429) <= (layer1_outputs(2131)) and not (layer1_outputs(4717));
    layer2_outputs(430) <= (layer1_outputs(4008)) or (layer1_outputs(444));
    layer2_outputs(431) <= (layer1_outputs(3181)) and not (layer1_outputs(2269));
    layer2_outputs(432) <= (layer1_outputs(142)) or (layer1_outputs(708));
    layer2_outputs(433) <= not(layer1_outputs(4989)) or (layer1_outputs(3868));
    layer2_outputs(434) <= (layer1_outputs(3734)) and not (layer1_outputs(1487));
    layer2_outputs(435) <= not((layer1_outputs(855)) or (layer1_outputs(3950)));
    layer2_outputs(436) <= (layer1_outputs(4030)) and not (layer1_outputs(760));
    layer2_outputs(437) <= '1';
    layer2_outputs(438) <= '0';
    layer2_outputs(439) <= layer1_outputs(2686);
    layer2_outputs(440) <= '1';
    layer2_outputs(441) <= not(layer1_outputs(4505));
    layer2_outputs(442) <= (layer1_outputs(707)) and (layer1_outputs(3748));
    layer2_outputs(443) <= (layer1_outputs(3277)) and not (layer1_outputs(20));
    layer2_outputs(444) <= not(layer1_outputs(3257));
    layer2_outputs(445) <= (layer1_outputs(4795)) and not (layer1_outputs(2769));
    layer2_outputs(446) <= not(layer1_outputs(3686)) or (layer1_outputs(4519));
    layer2_outputs(447) <= not((layer1_outputs(3513)) or (layer1_outputs(811)));
    layer2_outputs(448) <= not((layer1_outputs(3098)) or (layer1_outputs(1809)));
    layer2_outputs(449) <= (layer1_outputs(2327)) and (layer1_outputs(1462));
    layer2_outputs(450) <= (layer1_outputs(950)) or (layer1_outputs(5061));
    layer2_outputs(451) <= not(layer1_outputs(2081)) or (layer1_outputs(1109));
    layer2_outputs(452) <= '0';
    layer2_outputs(453) <= not(layer1_outputs(1683));
    layer2_outputs(454) <= (layer1_outputs(3881)) and not (layer1_outputs(3768));
    layer2_outputs(455) <= not((layer1_outputs(4827)) xor (layer1_outputs(4526)));
    layer2_outputs(456) <= not(layer1_outputs(493)) or (layer1_outputs(1606));
    layer2_outputs(457) <= not((layer1_outputs(2743)) or (layer1_outputs(1995)));
    layer2_outputs(458) <= layer1_outputs(1558);
    layer2_outputs(459) <= not(layer1_outputs(1268)) or (layer1_outputs(2694));
    layer2_outputs(460) <= (layer1_outputs(1634)) or (layer1_outputs(3141));
    layer2_outputs(461) <= (layer1_outputs(4430)) and not (layer1_outputs(3779));
    layer2_outputs(462) <= not((layer1_outputs(861)) or (layer1_outputs(2481)));
    layer2_outputs(463) <= not(layer1_outputs(4358)) or (layer1_outputs(137));
    layer2_outputs(464) <= '1';
    layer2_outputs(465) <= layer1_outputs(4431);
    layer2_outputs(466) <= (layer1_outputs(4643)) and not (layer1_outputs(2159));
    layer2_outputs(467) <= (layer1_outputs(2077)) or (layer1_outputs(3371));
    layer2_outputs(468) <= '1';
    layer2_outputs(469) <= (layer1_outputs(4452)) and (layer1_outputs(447));
    layer2_outputs(470) <= (layer1_outputs(1428)) and not (layer1_outputs(1797));
    layer2_outputs(471) <= (layer1_outputs(2861)) and not (layer1_outputs(21));
    layer2_outputs(472) <= (layer1_outputs(500)) and (layer1_outputs(2573));
    layer2_outputs(473) <= '0';
    layer2_outputs(474) <= (layer1_outputs(2233)) or (layer1_outputs(619));
    layer2_outputs(475) <= '1';
    layer2_outputs(476) <= '1';
    layer2_outputs(477) <= not((layer1_outputs(2299)) xor (layer1_outputs(3510)));
    layer2_outputs(478) <= layer1_outputs(1262);
    layer2_outputs(479) <= not(layer1_outputs(4543)) or (layer1_outputs(28));
    layer2_outputs(480) <= not((layer1_outputs(3255)) and (layer1_outputs(2669)));
    layer2_outputs(481) <= '0';
    layer2_outputs(482) <= '1';
    layer2_outputs(483) <= not((layer1_outputs(350)) and (layer1_outputs(3371)));
    layer2_outputs(484) <= not(layer1_outputs(1331));
    layer2_outputs(485) <= '0';
    layer2_outputs(486) <= not((layer1_outputs(3498)) or (layer1_outputs(3003)));
    layer2_outputs(487) <= (layer1_outputs(1632)) and (layer1_outputs(180));
    layer2_outputs(488) <= (layer1_outputs(3983)) or (layer1_outputs(4342));
    layer2_outputs(489) <= '1';
    layer2_outputs(490) <= '0';
    layer2_outputs(491) <= '0';
    layer2_outputs(492) <= (layer1_outputs(1224)) and (layer1_outputs(1223));
    layer2_outputs(493) <= not(layer1_outputs(1128)) or (layer1_outputs(3380));
    layer2_outputs(494) <= (layer1_outputs(2075)) or (layer1_outputs(4710));
    layer2_outputs(495) <= '1';
    layer2_outputs(496) <= not((layer1_outputs(3790)) and (layer1_outputs(2151)));
    layer2_outputs(497) <= layer1_outputs(2054);
    layer2_outputs(498) <= not(layer1_outputs(4016));
    layer2_outputs(499) <= (layer1_outputs(4858)) and not (layer1_outputs(3473));
    layer2_outputs(500) <= not((layer1_outputs(621)) and (layer1_outputs(974)));
    layer2_outputs(501) <= not(layer1_outputs(4603)) or (layer1_outputs(1675));
    layer2_outputs(502) <= (layer1_outputs(1805)) and (layer1_outputs(1180));
    layer2_outputs(503) <= '1';
    layer2_outputs(504) <= '0';
    layer2_outputs(505) <= '1';
    layer2_outputs(506) <= layer1_outputs(3025);
    layer2_outputs(507) <= layer1_outputs(1997);
    layer2_outputs(508) <= not(layer1_outputs(919));
    layer2_outputs(509) <= not(layer1_outputs(4660)) or (layer1_outputs(676));
    layer2_outputs(510) <= (layer1_outputs(1755)) or (layer1_outputs(2135));
    layer2_outputs(511) <= not((layer1_outputs(864)) or (layer1_outputs(4103)));
    layer2_outputs(512) <= not((layer1_outputs(2852)) and (layer1_outputs(2066)));
    layer2_outputs(513) <= (layer1_outputs(2790)) and not (layer1_outputs(4897));
    layer2_outputs(514) <= not((layer1_outputs(1237)) and (layer1_outputs(3879)));
    layer2_outputs(515) <= not((layer1_outputs(1886)) and (layer1_outputs(2014)));
    layer2_outputs(516) <= not((layer1_outputs(639)) or (layer1_outputs(4107)));
    layer2_outputs(517) <= (layer1_outputs(1221)) and not (layer1_outputs(1957));
    layer2_outputs(518) <= not(layer1_outputs(5028)) or (layer1_outputs(3403));
    layer2_outputs(519) <= not((layer1_outputs(1351)) and (layer1_outputs(1768)));
    layer2_outputs(520) <= (layer1_outputs(1621)) or (layer1_outputs(599));
    layer2_outputs(521) <= layer1_outputs(3784);
    layer2_outputs(522) <= not(layer1_outputs(2969)) or (layer1_outputs(5008));
    layer2_outputs(523) <= not((layer1_outputs(2483)) or (layer1_outputs(3838)));
    layer2_outputs(524) <= (layer1_outputs(739)) and not (layer1_outputs(4831));
    layer2_outputs(525) <= not(layer1_outputs(1061)) or (layer1_outputs(4813));
    layer2_outputs(526) <= (layer1_outputs(1423)) and not (layer1_outputs(1695));
    layer2_outputs(527) <= not((layer1_outputs(3553)) xor (layer1_outputs(375)));
    layer2_outputs(528) <= (layer1_outputs(4219)) or (layer1_outputs(4419));
    layer2_outputs(529) <= not(layer1_outputs(1487));
    layer2_outputs(530) <= (layer1_outputs(528)) and not (layer1_outputs(37));
    layer2_outputs(531) <= '1';
    layer2_outputs(532) <= '1';
    layer2_outputs(533) <= not(layer1_outputs(1965)) or (layer1_outputs(1811));
    layer2_outputs(534) <= not(layer1_outputs(4449)) or (layer1_outputs(4678));
    layer2_outputs(535) <= (layer1_outputs(4022)) and (layer1_outputs(4306));
    layer2_outputs(536) <= '0';
    layer2_outputs(537) <= (layer1_outputs(321)) and not (layer1_outputs(4682));
    layer2_outputs(538) <= (layer1_outputs(1312)) and (layer1_outputs(3603));
    layer2_outputs(539) <= '1';
    layer2_outputs(540) <= not((layer1_outputs(3746)) and (layer1_outputs(2831)));
    layer2_outputs(541) <= (layer1_outputs(3569)) and not (layer1_outputs(3576));
    layer2_outputs(542) <= not((layer1_outputs(973)) or (layer1_outputs(4892)));
    layer2_outputs(543) <= not((layer1_outputs(2544)) and (layer1_outputs(2953)));
    layer2_outputs(544) <= not(layer1_outputs(3145));
    layer2_outputs(545) <= (layer1_outputs(3363)) and not (layer1_outputs(2192));
    layer2_outputs(546) <= not(layer1_outputs(348)) or (layer1_outputs(2422));
    layer2_outputs(547) <= (layer1_outputs(3916)) or (layer1_outputs(2333));
    layer2_outputs(548) <= not(layer1_outputs(2718)) or (layer1_outputs(905));
    layer2_outputs(549) <= (layer1_outputs(4503)) or (layer1_outputs(4247));
    layer2_outputs(550) <= not(layer1_outputs(3425)) or (layer1_outputs(3357));
    layer2_outputs(551) <= (layer1_outputs(3668)) and (layer1_outputs(1955));
    layer2_outputs(552) <= (layer1_outputs(73)) and not (layer1_outputs(1036));
    layer2_outputs(553) <= not(layer1_outputs(736)) or (layer1_outputs(3739));
    layer2_outputs(554) <= not(layer1_outputs(3358)) or (layer1_outputs(440));
    layer2_outputs(555) <= not((layer1_outputs(3765)) or (layer1_outputs(4348)));
    layer2_outputs(556) <= '1';
    layer2_outputs(557) <= '0';
    layer2_outputs(558) <= layer1_outputs(1257);
    layer2_outputs(559) <= not(layer1_outputs(4559));
    layer2_outputs(560) <= (layer1_outputs(1871)) and not (layer1_outputs(3745));
    layer2_outputs(561) <= (layer1_outputs(3812)) and not (layer1_outputs(4061));
    layer2_outputs(562) <= (layer1_outputs(3988)) and not (layer1_outputs(896));
    layer2_outputs(563) <= (layer1_outputs(2020)) and (layer1_outputs(4855));
    layer2_outputs(564) <= (layer1_outputs(2955)) and not (layer1_outputs(2525));
    layer2_outputs(565) <= '1';
    layer2_outputs(566) <= '1';
    layer2_outputs(567) <= layer1_outputs(880);
    layer2_outputs(568) <= layer1_outputs(2753);
    layer2_outputs(569) <= (layer1_outputs(3484)) and (layer1_outputs(2540));
    layer2_outputs(570) <= '0';
    layer2_outputs(571) <= (layer1_outputs(4723)) and not (layer1_outputs(2748));
    layer2_outputs(572) <= not((layer1_outputs(2554)) xor (layer1_outputs(43)));
    layer2_outputs(573) <= (layer1_outputs(1828)) and not (layer1_outputs(316));
    layer2_outputs(574) <= not(layer1_outputs(386)) or (layer1_outputs(4830));
    layer2_outputs(575) <= '0';
    layer2_outputs(576) <= '0';
    layer2_outputs(577) <= '1';
    layer2_outputs(578) <= not((layer1_outputs(2547)) or (layer1_outputs(1356)));
    layer2_outputs(579) <= (layer1_outputs(3979)) xor (layer1_outputs(4818));
    layer2_outputs(580) <= '1';
    layer2_outputs(581) <= not((layer1_outputs(5084)) xor (layer1_outputs(1642)));
    layer2_outputs(582) <= not((layer1_outputs(1409)) or (layer1_outputs(2116)));
    layer2_outputs(583) <= not((layer1_outputs(5001)) and (layer1_outputs(4757)));
    layer2_outputs(584) <= (layer1_outputs(2452)) and not (layer1_outputs(273));
    layer2_outputs(585) <= not((layer1_outputs(816)) or (layer1_outputs(1373)));
    layer2_outputs(586) <= not((layer1_outputs(2320)) and (layer1_outputs(224)));
    layer2_outputs(587) <= '1';
    layer2_outputs(588) <= (layer1_outputs(584)) and (layer1_outputs(4168));
    layer2_outputs(589) <= (layer1_outputs(1405)) and not (layer1_outputs(3321));
    layer2_outputs(590) <= '0';
    layer2_outputs(591) <= layer1_outputs(1590);
    layer2_outputs(592) <= '1';
    layer2_outputs(593) <= (layer1_outputs(3238)) and not (layer1_outputs(2334));
    layer2_outputs(594) <= not((layer1_outputs(21)) or (layer1_outputs(4154)));
    layer2_outputs(595) <= (layer1_outputs(586)) and not (layer1_outputs(349));
    layer2_outputs(596) <= (layer1_outputs(171)) or (layer1_outputs(548));
    layer2_outputs(597) <= not(layer1_outputs(572)) or (layer1_outputs(2056));
    layer2_outputs(598) <= (layer1_outputs(3263)) or (layer1_outputs(1765));
    layer2_outputs(599) <= (layer1_outputs(2572)) and (layer1_outputs(567));
    layer2_outputs(600) <= (layer1_outputs(2526)) and not (layer1_outputs(2824));
    layer2_outputs(601) <= not(layer1_outputs(3648));
    layer2_outputs(602) <= (layer1_outputs(2899)) or (layer1_outputs(2973));
    layer2_outputs(603) <= not((layer1_outputs(2840)) or (layer1_outputs(267)));
    layer2_outputs(604) <= '0';
    layer2_outputs(605) <= (layer1_outputs(921)) or (layer1_outputs(3742));
    layer2_outputs(606) <= '0';
    layer2_outputs(607) <= (layer1_outputs(313)) and (layer1_outputs(1944));
    layer2_outputs(608) <= '1';
    layer2_outputs(609) <= not(layer1_outputs(1654)) or (layer1_outputs(87));
    layer2_outputs(610) <= not(layer1_outputs(3678));
    layer2_outputs(611) <= '0';
    layer2_outputs(612) <= (layer1_outputs(2200)) or (layer1_outputs(3665));
    layer2_outputs(613) <= not(layer1_outputs(1412));
    layer2_outputs(614) <= '1';
    layer2_outputs(615) <= layer1_outputs(4958);
    layer2_outputs(616) <= (layer1_outputs(860)) and (layer1_outputs(3352));
    layer2_outputs(617) <= (layer1_outputs(2167)) and not (layer1_outputs(1373));
    layer2_outputs(618) <= (layer1_outputs(2052)) and not (layer1_outputs(1704));
    layer2_outputs(619) <= not(layer1_outputs(2775)) or (layer1_outputs(1636));
    layer2_outputs(620) <= (layer1_outputs(2947)) or (layer1_outputs(2169));
    layer2_outputs(621) <= (layer1_outputs(4562)) and (layer1_outputs(4991));
    layer2_outputs(622) <= not(layer1_outputs(4480));
    layer2_outputs(623) <= '0';
    layer2_outputs(624) <= not((layer1_outputs(2111)) xor (layer1_outputs(2710)));
    layer2_outputs(625) <= layer1_outputs(314);
    layer2_outputs(626) <= not(layer1_outputs(3098));
    layer2_outputs(627) <= not((layer1_outputs(3908)) and (layer1_outputs(15)));
    layer2_outputs(628) <= (layer1_outputs(3477)) and not (layer1_outputs(2240));
    layer2_outputs(629) <= not((layer1_outputs(1710)) or (layer1_outputs(3150)));
    layer2_outputs(630) <= (layer1_outputs(1251)) or (layer1_outputs(717));
    layer2_outputs(631) <= (layer1_outputs(790)) and not (layer1_outputs(38));
    layer2_outputs(632) <= not(layer1_outputs(2534)) or (layer1_outputs(2660));
    layer2_outputs(633) <= not((layer1_outputs(2950)) or (layer1_outputs(4987)));
    layer2_outputs(634) <= (layer1_outputs(4904)) and (layer1_outputs(77));
    layer2_outputs(635) <= (layer1_outputs(3007)) and not (layer1_outputs(158));
    layer2_outputs(636) <= not(layer1_outputs(1948));
    layer2_outputs(637) <= not(layer1_outputs(5097)) or (layer1_outputs(1832));
    layer2_outputs(638) <= '1';
    layer2_outputs(639) <= (layer1_outputs(1422)) and not (layer1_outputs(1936));
    layer2_outputs(640) <= (layer1_outputs(2424)) and not (layer1_outputs(4313));
    layer2_outputs(641) <= (layer1_outputs(2396)) and not (layer1_outputs(2878));
    layer2_outputs(642) <= layer1_outputs(2337);
    layer2_outputs(643) <= (layer1_outputs(3793)) or (layer1_outputs(2310));
    layer2_outputs(644) <= (layer1_outputs(592)) and not (layer1_outputs(2978));
    layer2_outputs(645) <= (layer1_outputs(2147)) or (layer1_outputs(3968));
    layer2_outputs(646) <= not((layer1_outputs(2507)) xor (layer1_outputs(1537)));
    layer2_outputs(647) <= layer1_outputs(2175);
    layer2_outputs(648) <= (layer1_outputs(2242)) and (layer1_outputs(3382));
    layer2_outputs(649) <= not(layer1_outputs(1881));
    layer2_outputs(650) <= not(layer1_outputs(4815)) or (layer1_outputs(4880));
    layer2_outputs(651) <= not((layer1_outputs(1460)) xor (layer1_outputs(2870)));
    layer2_outputs(652) <= (layer1_outputs(4569)) or (layer1_outputs(2655));
    layer2_outputs(653) <= not(layer1_outputs(3821)) or (layer1_outputs(1290));
    layer2_outputs(654) <= (layer1_outputs(3121)) or (layer1_outputs(1344));
    layer2_outputs(655) <= not(layer1_outputs(3858)) or (layer1_outputs(2732));
    layer2_outputs(656) <= '0';
    layer2_outputs(657) <= '1';
    layer2_outputs(658) <= not(layer1_outputs(1790));
    layer2_outputs(659) <= (layer1_outputs(2997)) or (layer1_outputs(4179));
    layer2_outputs(660) <= layer1_outputs(4937);
    layer2_outputs(661) <= '0';
    layer2_outputs(662) <= layer1_outputs(3855);
    layer2_outputs(663) <= not(layer1_outputs(3818));
    layer2_outputs(664) <= (layer1_outputs(2475)) or (layer1_outputs(2970));
    layer2_outputs(665) <= (layer1_outputs(4646)) and not (layer1_outputs(3310));
    layer2_outputs(666) <= layer1_outputs(1330);
    layer2_outputs(667) <= layer1_outputs(1277);
    layer2_outputs(668) <= not((layer1_outputs(4887)) or (layer1_outputs(3286)));
    layer2_outputs(669) <= not(layer1_outputs(4093)) or (layer1_outputs(4551));
    layer2_outputs(670) <= not((layer1_outputs(1458)) and (layer1_outputs(1038)));
    layer2_outputs(671) <= '1';
    layer2_outputs(672) <= '1';
    layer2_outputs(673) <= not(layer1_outputs(2566));
    layer2_outputs(674) <= '0';
    layer2_outputs(675) <= (layer1_outputs(1346)) or (layer1_outputs(3500));
    layer2_outputs(676) <= not(layer1_outputs(3127));
    layer2_outputs(677) <= (layer1_outputs(4555)) and (layer1_outputs(831));
    layer2_outputs(678) <= '1';
    layer2_outputs(679) <= not(layer1_outputs(4320)) or (layer1_outputs(692));
    layer2_outputs(680) <= not((layer1_outputs(684)) or (layer1_outputs(222)));
    layer2_outputs(681) <= (layer1_outputs(2786)) and (layer1_outputs(1379));
    layer2_outputs(682) <= (layer1_outputs(4625)) and not (layer1_outputs(2593));
    layer2_outputs(683) <= not((layer1_outputs(3355)) xor (layer1_outputs(2905)));
    layer2_outputs(684) <= '1';
    layer2_outputs(685) <= not(layer1_outputs(1791)) or (layer1_outputs(2353));
    layer2_outputs(686) <= not(layer1_outputs(1153)) or (layer1_outputs(4178));
    layer2_outputs(687) <= not((layer1_outputs(4470)) and (layer1_outputs(3633)));
    layer2_outputs(688) <= (layer1_outputs(3418)) and not (layer1_outputs(262));
    layer2_outputs(689) <= '0';
    layer2_outputs(690) <= '1';
    layer2_outputs(691) <= '1';
    layer2_outputs(692) <= not((layer1_outputs(3226)) and (layer1_outputs(3840)));
    layer2_outputs(693) <= (layer1_outputs(1185)) and (layer1_outputs(3721));
    layer2_outputs(694) <= (layer1_outputs(904)) or (layer1_outputs(1090));
    layer2_outputs(695) <= (layer1_outputs(1133)) and not (layer1_outputs(3992));
    layer2_outputs(696) <= '0';
    layer2_outputs(697) <= (layer1_outputs(918)) and not (layer1_outputs(3947));
    layer2_outputs(698) <= not(layer1_outputs(1101));
    layer2_outputs(699) <= not(layer1_outputs(1684)) or (layer1_outputs(1188));
    layer2_outputs(700) <= '1';
    layer2_outputs(701) <= '0';
    layer2_outputs(702) <= not((layer1_outputs(4267)) or (layer1_outputs(706)));
    layer2_outputs(703) <= (layer1_outputs(317)) and not (layer1_outputs(3876));
    layer2_outputs(704) <= not(layer1_outputs(3426));
    layer2_outputs(705) <= not(layer1_outputs(3806));
    layer2_outputs(706) <= not(layer1_outputs(1063));
    layer2_outputs(707) <= not((layer1_outputs(2538)) and (layer1_outputs(1047)));
    layer2_outputs(708) <= layer1_outputs(4294);
    layer2_outputs(709) <= (layer1_outputs(4854)) and (layer1_outputs(871));
    layer2_outputs(710) <= '1';
    layer2_outputs(711) <= (layer1_outputs(1616)) xor (layer1_outputs(3934));
    layer2_outputs(712) <= (layer1_outputs(2323)) or (layer1_outputs(1068));
    layer2_outputs(713) <= not((layer1_outputs(532)) or (layer1_outputs(4151)));
    layer2_outputs(714) <= '1';
    layer2_outputs(715) <= not((layer1_outputs(851)) xor (layer1_outputs(882)));
    layer2_outputs(716) <= '0';
    layer2_outputs(717) <= not(layer1_outputs(648));
    layer2_outputs(718) <= (layer1_outputs(1068)) and not (layer1_outputs(3364));
    layer2_outputs(719) <= not(layer1_outputs(4132)) or (layer1_outputs(2881));
    layer2_outputs(720) <= not(layer1_outputs(4674)) or (layer1_outputs(541));
    layer2_outputs(721) <= not((layer1_outputs(2250)) or (layer1_outputs(1398)));
    layer2_outputs(722) <= not(layer1_outputs(3647));
    layer2_outputs(723) <= (layer1_outputs(4207)) and not (layer1_outputs(702));
    layer2_outputs(724) <= (layer1_outputs(2913)) or (layer1_outputs(2721));
    layer2_outputs(725) <= not(layer1_outputs(2708));
    layer2_outputs(726) <= layer1_outputs(3334);
    layer2_outputs(727) <= not(layer1_outputs(2519));
    layer2_outputs(728) <= not((layer1_outputs(278)) and (layer1_outputs(4629)));
    layer2_outputs(729) <= not((layer1_outputs(2767)) or (layer1_outputs(158)));
    layer2_outputs(730) <= not((layer1_outputs(3972)) or (layer1_outputs(4325)));
    layer2_outputs(731) <= not((layer1_outputs(989)) or (layer1_outputs(3740)));
    layer2_outputs(732) <= '0';
    layer2_outputs(733) <= layer1_outputs(2257);
    layer2_outputs(734) <= (layer1_outputs(3550)) and not (layer1_outputs(3462));
    layer2_outputs(735) <= (layer1_outputs(32)) and not (layer1_outputs(385));
    layer2_outputs(736) <= (layer1_outputs(2723)) or (layer1_outputs(2294));
    layer2_outputs(737) <= layer1_outputs(3243);
    layer2_outputs(738) <= not((layer1_outputs(4768)) or (layer1_outputs(2670)));
    layer2_outputs(739) <= (layer1_outputs(1147)) or (layer1_outputs(5109));
    layer2_outputs(740) <= layer1_outputs(2050);
    layer2_outputs(741) <= not(layer1_outputs(600));
    layer2_outputs(742) <= layer1_outputs(1328);
    layer2_outputs(743) <= not((layer1_outputs(3174)) and (layer1_outputs(3103)));
    layer2_outputs(744) <= not((layer1_outputs(4115)) or (layer1_outputs(3717)));
    layer2_outputs(745) <= layer1_outputs(858);
    layer2_outputs(746) <= (layer1_outputs(4399)) xor (layer1_outputs(1822));
    layer2_outputs(747) <= not(layer1_outputs(490));
    layer2_outputs(748) <= (layer1_outputs(4608)) or (layer1_outputs(1687));
    layer2_outputs(749) <= (layer1_outputs(3190)) and not (layer1_outputs(1577));
    layer2_outputs(750) <= not(layer1_outputs(2390)) or (layer1_outputs(5071));
    layer2_outputs(751) <= not(layer1_outputs(1691)) or (layer1_outputs(5072));
    layer2_outputs(752) <= (layer1_outputs(1324)) or (layer1_outputs(5));
    layer2_outputs(753) <= (layer1_outputs(3644)) or (layer1_outputs(3035));
    layer2_outputs(754) <= (layer1_outputs(2576)) and (layer1_outputs(2285));
    layer2_outputs(755) <= (layer1_outputs(3000)) and not (layer1_outputs(916));
    layer2_outputs(756) <= '1';
    layer2_outputs(757) <= not(layer1_outputs(3398)) or (layer1_outputs(2107));
    layer2_outputs(758) <= (layer1_outputs(382)) or (layer1_outputs(3728));
    layer2_outputs(759) <= not((layer1_outputs(1635)) or (layer1_outputs(1533)));
    layer2_outputs(760) <= not(layer1_outputs(4307));
    layer2_outputs(761) <= layer1_outputs(2938);
    layer2_outputs(762) <= '1';
    layer2_outputs(763) <= '1';
    layer2_outputs(764) <= not(layer1_outputs(41)) or (layer1_outputs(3132));
    layer2_outputs(765) <= (layer1_outputs(219)) or (layer1_outputs(3592));
    layer2_outputs(766) <= (layer1_outputs(2646)) or (layer1_outputs(4697));
    layer2_outputs(767) <= not((layer1_outputs(4128)) or (layer1_outputs(2597)));
    layer2_outputs(768) <= not((layer1_outputs(2078)) and (layer1_outputs(1565)));
    layer2_outputs(769) <= '0';
    layer2_outputs(770) <= (layer1_outputs(1164)) and not (layer1_outputs(4843));
    layer2_outputs(771) <= '1';
    layer2_outputs(772) <= '0';
    layer2_outputs(773) <= not(layer1_outputs(3405)) or (layer1_outputs(180));
    layer2_outputs(774) <= '1';
    layer2_outputs(775) <= '1';
    layer2_outputs(776) <= '1';
    layer2_outputs(777) <= not(layer1_outputs(3395)) or (layer1_outputs(1936));
    layer2_outputs(778) <= (layer1_outputs(2560)) and (layer1_outputs(4320));
    layer2_outputs(779) <= '1';
    layer2_outputs(780) <= layer1_outputs(4045);
    layer2_outputs(781) <= '0';
    layer2_outputs(782) <= not(layer1_outputs(4922));
    layer2_outputs(783) <= '0';
    layer2_outputs(784) <= (layer1_outputs(693)) and (layer1_outputs(4663));
    layer2_outputs(785) <= '1';
    layer2_outputs(786) <= not((layer1_outputs(1060)) and (layer1_outputs(4633)));
    layer2_outputs(787) <= not((layer1_outputs(3210)) or (layer1_outputs(3391)));
    layer2_outputs(788) <= not(layer1_outputs(4499)) or (layer1_outputs(1029));
    layer2_outputs(789) <= (layer1_outputs(524)) and not (layer1_outputs(4600));
    layer2_outputs(790) <= not((layer1_outputs(61)) or (layer1_outputs(4581)));
    layer2_outputs(791) <= (layer1_outputs(774)) and (layer1_outputs(4599));
    layer2_outputs(792) <= not(layer1_outputs(3830));
    layer2_outputs(793) <= not((layer1_outputs(4640)) and (layer1_outputs(3626)));
    layer2_outputs(794) <= not(layer1_outputs(2112));
    layer2_outputs(795) <= layer1_outputs(1243);
    layer2_outputs(796) <= not(layer1_outputs(3480)) or (layer1_outputs(1848));
    layer2_outputs(797) <= (layer1_outputs(4636)) and not (layer1_outputs(1862));
    layer2_outputs(798) <= not((layer1_outputs(2965)) or (layer1_outputs(4337)));
    layer2_outputs(799) <= not(layer1_outputs(930)) or (layer1_outputs(942));
    layer2_outputs(800) <= (layer1_outputs(4896)) and (layer1_outputs(139));
    layer2_outputs(801) <= '1';
    layer2_outputs(802) <= (layer1_outputs(4790)) and (layer1_outputs(3125));
    layer2_outputs(803) <= not(layer1_outputs(4732)) or (layer1_outputs(557));
    layer2_outputs(804) <= (layer1_outputs(281)) and not (layer1_outputs(3543));
    layer2_outputs(805) <= (layer1_outputs(1411)) and not (layer1_outputs(3965));
    layer2_outputs(806) <= not(layer1_outputs(3537));
    layer2_outputs(807) <= not((layer1_outputs(2917)) or (layer1_outputs(517)));
    layer2_outputs(808) <= not(layer1_outputs(4144));
    layer2_outputs(809) <= (layer1_outputs(2278)) and not (layer1_outputs(1692));
    layer2_outputs(810) <= not(layer1_outputs(3465)) or (layer1_outputs(4333));
    layer2_outputs(811) <= '1';
    layer2_outputs(812) <= not((layer1_outputs(12)) or (layer1_outputs(4833)));
    layer2_outputs(813) <= (layer1_outputs(3505)) and not (layer1_outputs(3056));
    layer2_outputs(814) <= not(layer1_outputs(3624));
    layer2_outputs(815) <= layer1_outputs(2022);
    layer2_outputs(816) <= (layer1_outputs(3803)) or (layer1_outputs(1319));
    layer2_outputs(817) <= not((layer1_outputs(2993)) and (layer1_outputs(3118)));
    layer2_outputs(818) <= '0';
    layer2_outputs(819) <= (layer1_outputs(2741)) or (layer1_outputs(4838));
    layer2_outputs(820) <= (layer1_outputs(4508)) and not (layer1_outputs(3260));
    layer2_outputs(821) <= (layer1_outputs(2249)) or (layer1_outputs(242));
    layer2_outputs(822) <= (layer1_outputs(1120)) and (layer1_outputs(2730));
    layer2_outputs(823) <= '1';
    layer2_outputs(824) <= (layer1_outputs(1929)) and (layer1_outputs(4876));
    layer2_outputs(825) <= (layer1_outputs(1316)) and not (layer1_outputs(1479));
    layer2_outputs(826) <= (layer1_outputs(4762)) and not (layer1_outputs(3388));
    layer2_outputs(827) <= (layer1_outputs(356)) and not (layer1_outputs(1135));
    layer2_outputs(828) <= not((layer1_outputs(2796)) and (layer1_outputs(4686)));
    layer2_outputs(829) <= not(layer1_outputs(4979)) or (layer1_outputs(231));
    layer2_outputs(830) <= not((layer1_outputs(3203)) and (layer1_outputs(2668)));
    layer2_outputs(831) <= (layer1_outputs(4452)) and (layer1_outputs(935));
    layer2_outputs(832) <= not((layer1_outputs(4624)) or (layer1_outputs(2305)));
    layer2_outputs(833) <= not(layer1_outputs(4197)) or (layer1_outputs(781));
    layer2_outputs(834) <= (layer1_outputs(4125)) and (layer1_outputs(1577));
    layer2_outputs(835) <= '1';
    layer2_outputs(836) <= not((layer1_outputs(4890)) and (layer1_outputs(2672)));
    layer2_outputs(837) <= not(layer1_outputs(3497));
    layer2_outputs(838) <= not((layer1_outputs(1662)) or (layer1_outputs(2742)));
    layer2_outputs(839) <= not(layer1_outputs(3438)) or (layer1_outputs(3055));
    layer2_outputs(840) <= not((layer1_outputs(1097)) and (layer1_outputs(1612)));
    layer2_outputs(841) <= '0';
    layer2_outputs(842) <= not(layer1_outputs(1709)) or (layer1_outputs(769));
    layer2_outputs(843) <= not((layer1_outputs(1314)) xor (layer1_outputs(787)));
    layer2_outputs(844) <= '0';
    layer2_outputs(845) <= (layer1_outputs(972)) or (layer1_outputs(605));
    layer2_outputs(846) <= '0';
    layer2_outputs(847) <= (layer1_outputs(1581)) and not (layer1_outputs(2852));
    layer2_outputs(848) <= '1';
    layer2_outputs(849) <= (layer1_outputs(1955)) and not (layer1_outputs(4014));
    layer2_outputs(850) <= '1';
    layer2_outputs(851) <= '0';
    layer2_outputs(852) <= not((layer1_outputs(1593)) xor (layer1_outputs(874)));
    layer2_outputs(853) <= '0';
    layer2_outputs(854) <= '1';
    layer2_outputs(855) <= not(layer1_outputs(2488)) or (layer1_outputs(4571));
    layer2_outputs(856) <= not((layer1_outputs(5080)) and (layer1_outputs(4614)));
    layer2_outputs(857) <= not(layer1_outputs(1723));
    layer2_outputs(858) <= (layer1_outputs(2830)) xor (layer1_outputs(1518));
    layer2_outputs(859) <= '1';
    layer2_outputs(860) <= layer1_outputs(873);
    layer2_outputs(861) <= (layer1_outputs(4062)) and not (layer1_outputs(871));
    layer2_outputs(862) <= layer1_outputs(2095);
    layer2_outputs(863) <= not((layer1_outputs(5100)) or (layer1_outputs(2993)));
    layer2_outputs(864) <= '1';
    layer2_outputs(865) <= '1';
    layer2_outputs(866) <= '1';
    layer2_outputs(867) <= '0';
    layer2_outputs(868) <= layer1_outputs(883);
    layer2_outputs(869) <= layer1_outputs(3762);
    layer2_outputs(870) <= layer1_outputs(1984);
    layer2_outputs(871) <= '1';
    layer2_outputs(872) <= not((layer1_outputs(46)) or (layer1_outputs(1849)));
    layer2_outputs(873) <= '0';
    layer2_outputs(874) <= '1';
    layer2_outputs(875) <= layer1_outputs(426);
    layer2_outputs(876) <= (layer1_outputs(1108)) and not (layer1_outputs(4798));
    layer2_outputs(877) <= not(layer1_outputs(3160)) or (layer1_outputs(1634));
    layer2_outputs(878) <= layer1_outputs(239);
    layer2_outputs(879) <= not(layer1_outputs(3247)) or (layer1_outputs(2391));
    layer2_outputs(880) <= not((layer1_outputs(5017)) or (layer1_outputs(399)));
    layer2_outputs(881) <= (layer1_outputs(3116)) and (layer1_outputs(1850));
    layer2_outputs(882) <= (layer1_outputs(4130)) and not (layer1_outputs(2245));
    layer2_outputs(883) <= layer1_outputs(4869);
    layer2_outputs(884) <= layer1_outputs(4408);
    layer2_outputs(885) <= (layer1_outputs(2906)) and not (layer1_outputs(3564));
    layer2_outputs(886) <= not(layer1_outputs(1723)) or (layer1_outputs(4268));
    layer2_outputs(887) <= not((layer1_outputs(402)) and (layer1_outputs(4635)));
    layer2_outputs(888) <= '1';
    layer2_outputs(889) <= (layer1_outputs(1045)) or (layer1_outputs(1494));
    layer2_outputs(890) <= '0';
    layer2_outputs(891) <= not((layer1_outputs(2814)) or (layer1_outputs(2811)));
    layer2_outputs(892) <= (layer1_outputs(205)) xor (layer1_outputs(4700));
    layer2_outputs(893) <= '1';
    layer2_outputs(894) <= not(layer1_outputs(2680)) or (layer1_outputs(4763));
    layer2_outputs(895) <= not(layer1_outputs(2568));
    layer2_outputs(896) <= not(layer1_outputs(1312)) or (layer1_outputs(18));
    layer2_outputs(897) <= not((layer1_outputs(1458)) or (layer1_outputs(675)));
    layer2_outputs(898) <= (layer1_outputs(1930)) and not (layer1_outputs(3288));
    layer2_outputs(899) <= layer1_outputs(4994);
    layer2_outputs(900) <= '0';
    layer2_outputs(901) <= '0';
    layer2_outputs(902) <= '1';
    layer2_outputs(903) <= '1';
    layer2_outputs(904) <= not((layer1_outputs(5095)) or (layer1_outputs(23)));
    layer2_outputs(905) <= (layer1_outputs(3490)) and (layer1_outputs(249));
    layer2_outputs(906) <= layer1_outputs(410);
    layer2_outputs(907) <= (layer1_outputs(1255)) and not (layer1_outputs(4841));
    layer2_outputs(908) <= not((layer1_outputs(4273)) xor (layer1_outputs(2505)));
    layer2_outputs(909) <= not(layer1_outputs(1558)) or (layer1_outputs(4197));
    layer2_outputs(910) <= not(layer1_outputs(1738)) or (layer1_outputs(1533));
    layer2_outputs(911) <= layer1_outputs(5009);
    layer2_outputs(912) <= layer1_outputs(4187);
    layer2_outputs(913) <= not(layer1_outputs(1421)) or (layer1_outputs(5050));
    layer2_outputs(914) <= not(layer1_outputs(4929));
    layer2_outputs(915) <= (layer1_outputs(4811)) xor (layer1_outputs(4412));
    layer2_outputs(916) <= (layer1_outputs(71)) and (layer1_outputs(2869));
    layer2_outputs(917) <= not((layer1_outputs(3284)) and (layer1_outputs(3108)));
    layer2_outputs(918) <= (layer1_outputs(2897)) and not (layer1_outputs(484));
    layer2_outputs(919) <= (layer1_outputs(117)) and (layer1_outputs(1694));
    layer2_outputs(920) <= '1';
    layer2_outputs(921) <= '1';
    layer2_outputs(922) <= (layer1_outputs(1907)) and not (layer1_outputs(4518));
    layer2_outputs(923) <= not(layer1_outputs(4316)) or (layer1_outputs(2975));
    layer2_outputs(924) <= '0';
    layer2_outputs(925) <= not(layer1_outputs(2367)) or (layer1_outputs(4782));
    layer2_outputs(926) <= layer1_outputs(1432);
    layer2_outputs(927) <= not(layer1_outputs(801)) or (layer1_outputs(411));
    layer2_outputs(928) <= not(layer1_outputs(3250)) or (layer1_outputs(4048));
    layer2_outputs(929) <= '0';
    layer2_outputs(930) <= (layer1_outputs(240)) and not (layer1_outputs(4772));
    layer2_outputs(931) <= '0';
    layer2_outputs(932) <= '1';
    layer2_outputs(933) <= not(layer1_outputs(890));
    layer2_outputs(934) <= '1';
    layer2_outputs(935) <= layer1_outputs(1121);
    layer2_outputs(936) <= (layer1_outputs(4244)) or (layer1_outputs(1966));
    layer2_outputs(937) <= not((layer1_outputs(4760)) or (layer1_outputs(878)));
    layer2_outputs(938) <= not(layer1_outputs(4038)) or (layer1_outputs(2587));
    layer2_outputs(939) <= layer1_outputs(3075);
    layer2_outputs(940) <= (layer1_outputs(758)) or (layer1_outputs(2603));
    layer2_outputs(941) <= not(layer1_outputs(994)) or (layer1_outputs(3459));
    layer2_outputs(942) <= not((layer1_outputs(4072)) and (layer1_outputs(3237)));
    layer2_outputs(943) <= (layer1_outputs(2451)) or (layer1_outputs(2394));
    layer2_outputs(944) <= '0';
    layer2_outputs(945) <= (layer1_outputs(2318)) and not (layer1_outputs(1908));
    layer2_outputs(946) <= (layer1_outputs(2898)) or (layer1_outputs(1958));
    layer2_outputs(947) <= (layer1_outputs(786)) or (layer1_outputs(704));
    layer2_outputs(948) <= (layer1_outputs(3844)) and (layer1_outputs(457));
    layer2_outputs(949) <= not(layer1_outputs(3150));
    layer2_outputs(950) <= not((layer1_outputs(1659)) or (layer1_outputs(5102)));
    layer2_outputs(951) <= '0';
    layer2_outputs(952) <= not(layer1_outputs(3664));
    layer2_outputs(953) <= layer1_outputs(2489);
    layer2_outputs(954) <= '1';
    layer2_outputs(955) <= not(layer1_outputs(799)) or (layer1_outputs(2849));
    layer2_outputs(956) <= '0';
    layer2_outputs(957) <= not(layer1_outputs(798));
    layer2_outputs(958) <= not((layer1_outputs(2940)) and (layer1_outputs(4969)));
    layer2_outputs(959) <= '1';
    layer2_outputs(960) <= layer1_outputs(1740);
    layer2_outputs(961) <= not((layer1_outputs(490)) or (layer1_outputs(2836)));
    layer2_outputs(962) <= layer1_outputs(2571);
    layer2_outputs(963) <= layer1_outputs(1974);
    layer2_outputs(964) <= not(layer1_outputs(2413));
    layer2_outputs(965) <= (layer1_outputs(1831)) or (layer1_outputs(4362));
    layer2_outputs(966) <= not((layer1_outputs(1676)) xor (layer1_outputs(1629)));
    layer2_outputs(967) <= layer1_outputs(4912);
    layer2_outputs(968) <= (layer1_outputs(2603)) and not (layer1_outputs(1338));
    layer2_outputs(969) <= not((layer1_outputs(4120)) and (layer1_outputs(658)));
    layer2_outputs(970) <= not(layer1_outputs(1906));
    layer2_outputs(971) <= (layer1_outputs(3495)) and (layer1_outputs(4837));
    layer2_outputs(972) <= '1';
    layer2_outputs(973) <= layer1_outputs(1022);
    layer2_outputs(974) <= not((layer1_outputs(2755)) and (layer1_outputs(3690)));
    layer2_outputs(975) <= not((layer1_outputs(301)) or (layer1_outputs(2888)));
    layer2_outputs(976) <= '1';
    layer2_outputs(977) <= (layer1_outputs(4443)) and not (layer1_outputs(1583));
    layer2_outputs(978) <= '0';
    layer2_outputs(979) <= '1';
    layer2_outputs(980) <= (layer1_outputs(1074)) and (layer1_outputs(4227));
    layer2_outputs(981) <= not(layer1_outputs(61)) or (layer1_outputs(2181));
    layer2_outputs(982) <= not((layer1_outputs(2180)) or (layer1_outputs(4932)));
    layer2_outputs(983) <= (layer1_outputs(1825)) and not (layer1_outputs(4607));
    layer2_outputs(984) <= not(layer1_outputs(427));
    layer2_outputs(985) <= (layer1_outputs(5053)) and (layer1_outputs(1339));
    layer2_outputs(986) <= not(layer1_outputs(912)) or (layer1_outputs(4371));
    layer2_outputs(987) <= layer1_outputs(3915);
    layer2_outputs(988) <= (layer1_outputs(2588)) and (layer1_outputs(42));
    layer2_outputs(989) <= (layer1_outputs(3346)) and not (layer1_outputs(552));
    layer2_outputs(990) <= not((layer1_outputs(4663)) or (layer1_outputs(3783)));
    layer2_outputs(991) <= (layer1_outputs(3500)) and not (layer1_outputs(3223));
    layer2_outputs(992) <= (layer1_outputs(3670)) and not (layer1_outputs(2442));
    layer2_outputs(993) <= (layer1_outputs(2706)) and not (layer1_outputs(1191));
    layer2_outputs(994) <= (layer1_outputs(4052)) or (layer1_outputs(4863));
    layer2_outputs(995) <= not((layer1_outputs(3360)) or (layer1_outputs(1480)));
    layer2_outputs(996) <= (layer1_outputs(1762)) and (layer1_outputs(616));
    layer2_outputs(997) <= not(layer1_outputs(1512));
    layer2_outputs(998) <= '1';
    layer2_outputs(999) <= (layer1_outputs(4842)) or (layer1_outputs(13));
    layer2_outputs(1000) <= not((layer1_outputs(953)) and (layer1_outputs(597)));
    layer2_outputs(1001) <= (layer1_outputs(1983)) and not (layer1_outputs(4459));
    layer2_outputs(1002) <= not(layer1_outputs(97)) or (layer1_outputs(1085));
    layer2_outputs(1003) <= '1';
    layer2_outputs(1004) <= not(layer1_outputs(4992)) or (layer1_outputs(4933));
    layer2_outputs(1005) <= layer1_outputs(2785);
    layer2_outputs(1006) <= '0';
    layer2_outputs(1007) <= (layer1_outputs(995)) and (layer1_outputs(1749));
    layer2_outputs(1008) <= (layer1_outputs(837)) and (layer1_outputs(4218));
    layer2_outputs(1009) <= not(layer1_outputs(1323));
    layer2_outputs(1010) <= (layer1_outputs(1871)) and not (layer1_outputs(1821));
    layer2_outputs(1011) <= '0';
    layer2_outputs(1012) <= (layer1_outputs(3044)) and (layer1_outputs(4648));
    layer2_outputs(1013) <= '1';
    layer2_outputs(1014) <= not((layer1_outputs(4870)) and (layer1_outputs(4651)));
    layer2_outputs(1015) <= (layer1_outputs(2857)) and not (layer1_outputs(2793));
    layer2_outputs(1016) <= (layer1_outputs(3947)) and (layer1_outputs(3105));
    layer2_outputs(1017) <= '0';
    layer2_outputs(1018) <= not(layer1_outputs(4399));
    layer2_outputs(1019) <= not(layer1_outputs(4232)) or (layer1_outputs(1969));
    layer2_outputs(1020) <= '1';
    layer2_outputs(1021) <= '1';
    layer2_outputs(1022) <= '1';
    layer2_outputs(1023) <= '0';
    layer2_outputs(1024) <= not(layer1_outputs(900)) or (layer1_outputs(432));
    layer2_outputs(1025) <= '1';
    layer2_outputs(1026) <= not(layer1_outputs(4138));
    layer2_outputs(1027) <= '1';
    layer2_outputs(1028) <= not(layer1_outputs(2348));
    layer2_outputs(1029) <= not(layer1_outputs(3662)) or (layer1_outputs(3613));
    layer2_outputs(1030) <= (layer1_outputs(3465)) and (layer1_outputs(3542));
    layer2_outputs(1031) <= '1';
    layer2_outputs(1032) <= not(layer1_outputs(3826)) or (layer1_outputs(957));
    layer2_outputs(1033) <= layer1_outputs(286);
    layer2_outputs(1034) <= (layer1_outputs(4170)) and not (layer1_outputs(354));
    layer2_outputs(1035) <= (layer1_outputs(1991)) or (layer1_outputs(884));
    layer2_outputs(1036) <= not((layer1_outputs(4835)) or (layer1_outputs(5115)));
    layer2_outputs(1037) <= '0';
    layer2_outputs(1038) <= (layer1_outputs(3885)) and not (layer1_outputs(2062));
    layer2_outputs(1039) <= not(layer1_outputs(3714));
    layer2_outputs(1040) <= not(layer1_outputs(365)) or (layer1_outputs(215));
    layer2_outputs(1041) <= layer1_outputs(4615);
    layer2_outputs(1042) <= '1';
    layer2_outputs(1043) <= not((layer1_outputs(2864)) and (layer1_outputs(1394)));
    layer2_outputs(1044) <= (layer1_outputs(137)) or (layer1_outputs(4410));
    layer2_outputs(1045) <= '1';
    layer2_outputs(1046) <= '0';
    layer2_outputs(1047) <= not(layer1_outputs(4424));
    layer2_outputs(1048) <= (layer1_outputs(4068)) or (layer1_outputs(3275));
    layer2_outputs(1049) <= (layer1_outputs(1199)) and not (layer1_outputs(1557));
    layer2_outputs(1050) <= not((layer1_outputs(3350)) or (layer1_outputs(836)));
    layer2_outputs(1051) <= (layer1_outputs(1597)) and not (layer1_outputs(561));
    layer2_outputs(1052) <= not(layer1_outputs(2694));
    layer2_outputs(1053) <= (layer1_outputs(2423)) and (layer1_outputs(2255));
    layer2_outputs(1054) <= not(layer1_outputs(3576)) or (layer1_outputs(4160));
    layer2_outputs(1055) <= layer1_outputs(4346);
    layer2_outputs(1056) <= '1';
    layer2_outputs(1057) <= layer1_outputs(881);
    layer2_outputs(1058) <= layer1_outputs(1344);
    layer2_outputs(1059) <= (layer1_outputs(461)) and not (layer1_outputs(2702));
    layer2_outputs(1060) <= (layer1_outputs(2586)) and not (layer1_outputs(863));
    layer2_outputs(1061) <= layer1_outputs(842);
    layer2_outputs(1062) <= (layer1_outputs(2766)) and not (layer1_outputs(3179));
    layer2_outputs(1063) <= (layer1_outputs(2872)) and (layer1_outputs(2922));
    layer2_outputs(1064) <= not((layer1_outputs(2443)) and (layer1_outputs(2372)));
    layer2_outputs(1065) <= not(layer1_outputs(975)) or (layer1_outputs(40));
    layer2_outputs(1066) <= layer1_outputs(166);
    layer2_outputs(1067) <= not(layer1_outputs(3482));
    layer2_outputs(1068) <= layer1_outputs(1474);
    layer2_outputs(1069) <= layer1_outputs(4162);
    layer2_outputs(1070) <= '1';
    layer2_outputs(1071) <= '1';
    layer2_outputs(1072) <= layer1_outputs(2778);
    layer2_outputs(1073) <= not((layer1_outputs(322)) or (layer1_outputs(1293)));
    layer2_outputs(1074) <= layer1_outputs(2389);
    layer2_outputs(1075) <= not(layer1_outputs(3641)) or (layer1_outputs(1755));
    layer2_outputs(1076) <= (layer1_outputs(1834)) and not (layer1_outputs(2077));
    layer2_outputs(1077) <= '0';
    layer2_outputs(1078) <= layer1_outputs(3092);
    layer2_outputs(1079) <= not((layer1_outputs(956)) and (layer1_outputs(2314)));
    layer2_outputs(1080) <= layer1_outputs(2400);
    layer2_outputs(1081) <= (layer1_outputs(2419)) and not (layer1_outputs(3541));
    layer2_outputs(1082) <= layer1_outputs(598);
    layer2_outputs(1083) <= (layer1_outputs(1489)) and not (layer1_outputs(2064));
    layer2_outputs(1084) <= layer1_outputs(4935);
    layer2_outputs(1085) <= not((layer1_outputs(2812)) and (layer1_outputs(4456)));
    layer2_outputs(1086) <= '0';
    layer2_outputs(1087) <= (layer1_outputs(2650)) and (layer1_outputs(2219));
    layer2_outputs(1088) <= layer1_outputs(3241);
    layer2_outputs(1089) <= '0';
    layer2_outputs(1090) <= (layer1_outputs(4305)) and not (layer1_outputs(3453));
    layer2_outputs(1091) <= not(layer1_outputs(3209));
    layer2_outputs(1092) <= (layer1_outputs(1455)) or (layer1_outputs(4332));
    layer2_outputs(1093) <= not((layer1_outputs(2987)) and (layer1_outputs(643)));
    layer2_outputs(1094) <= not((layer1_outputs(1385)) and (layer1_outputs(120)));
    layer2_outputs(1095) <= '1';
    layer2_outputs(1096) <= not(layer1_outputs(3959)) or (layer1_outputs(4301));
    layer2_outputs(1097) <= '0';
    layer2_outputs(1098) <= not((layer1_outputs(4483)) and (layer1_outputs(665)));
    layer2_outputs(1099) <= (layer1_outputs(275)) and not (layer1_outputs(406));
    layer2_outputs(1100) <= (layer1_outputs(1555)) or (layer1_outputs(3082));
    layer2_outputs(1101) <= '1';
    layer2_outputs(1102) <= not((layer1_outputs(2704)) and (layer1_outputs(4259)));
    layer2_outputs(1103) <= not(layer1_outputs(2806));
    layer2_outputs(1104) <= '1';
    layer2_outputs(1105) <= layer1_outputs(4248);
    layer2_outputs(1106) <= not(layer1_outputs(4060)) or (layer1_outputs(4639));
    layer2_outputs(1107) <= (layer1_outputs(356)) or (layer1_outputs(4567));
    layer2_outputs(1108) <= not(layer1_outputs(2684)) or (layer1_outputs(333));
    layer2_outputs(1109) <= '1';
    layer2_outputs(1110) <= not((layer1_outputs(3547)) or (layer1_outputs(3143)));
    layer2_outputs(1111) <= '0';
    layer2_outputs(1112) <= (layer1_outputs(1433)) or (layer1_outputs(4019));
    layer2_outputs(1113) <= not((layer1_outputs(3671)) and (layer1_outputs(2033)));
    layer2_outputs(1114) <= not(layer1_outputs(4163));
    layer2_outputs(1115) <= (layer1_outputs(3657)) and not (layer1_outputs(4719));
    layer2_outputs(1116) <= not((layer1_outputs(1207)) and (layer1_outputs(2999)));
    layer2_outputs(1117) <= '0';
    layer2_outputs(1118) <= (layer1_outputs(4816)) and not (layer1_outputs(2090));
    layer2_outputs(1119) <= '1';
    layer2_outputs(1120) <= '0';
    layer2_outputs(1121) <= (layer1_outputs(2401)) and (layer1_outputs(105));
    layer2_outputs(1122) <= not(layer1_outputs(1465)) or (layer1_outputs(1403));
    layer2_outputs(1123) <= (layer1_outputs(1325)) and (layer1_outputs(1392));
    layer2_outputs(1124) <= not(layer1_outputs(907)) or (layer1_outputs(5014));
    layer2_outputs(1125) <= not(layer1_outputs(2130)) or (layer1_outputs(1707));
    layer2_outputs(1126) <= '1';
    layer2_outputs(1127) <= not(layer1_outputs(817)) or (layer1_outputs(1823));
    layer2_outputs(1128) <= not((layer1_outputs(3757)) and (layer1_outputs(2582)));
    layer2_outputs(1129) <= '1';
    layer2_outputs(1130) <= layer1_outputs(3416);
    layer2_outputs(1131) <= not(layer1_outputs(729));
    layer2_outputs(1132) <= '0';
    layer2_outputs(1133) <= '1';
    layer2_outputs(1134) <= not(layer1_outputs(656)) or (layer1_outputs(160));
    layer2_outputs(1135) <= not(layer1_outputs(4645));
    layer2_outputs(1136) <= not(layer1_outputs(293)) or (layer1_outputs(685));
    layer2_outputs(1137) <= (layer1_outputs(3516)) and not (layer1_outputs(1596));
    layer2_outputs(1138) <= not(layer1_outputs(3135));
    layer2_outputs(1139) <= '1';
    layer2_outputs(1140) <= not(layer1_outputs(310)) or (layer1_outputs(1598));
    layer2_outputs(1141) <= (layer1_outputs(176)) and not (layer1_outputs(405));
    layer2_outputs(1142) <= (layer1_outputs(4704)) and not (layer1_outputs(4656));
    layer2_outputs(1143) <= not(layer1_outputs(2664));
    layer2_outputs(1144) <= '1';
    layer2_outputs(1145) <= not(layer1_outputs(2638)) or (layer1_outputs(955));
    layer2_outputs(1146) <= not((layer1_outputs(2569)) and (layer1_outputs(216)));
    layer2_outputs(1147) <= '1';
    layer2_outputs(1148) <= (layer1_outputs(512)) and not (layer1_outputs(1680));
    layer2_outputs(1149) <= '0';
    layer2_outputs(1150) <= not(layer1_outputs(4183)) or (layer1_outputs(3038));
    layer2_outputs(1151) <= (layer1_outputs(3427)) and not (layer1_outputs(2441));
    layer2_outputs(1152) <= '1';
    layer2_outputs(1153) <= not((layer1_outputs(2079)) and (layer1_outputs(4049)));
    layer2_outputs(1154) <= '1';
    layer2_outputs(1155) <= not(layer1_outputs(1377)) or (layer1_outputs(662));
    layer2_outputs(1156) <= not(layer1_outputs(2791)) or (layer1_outputs(3295));
    layer2_outputs(1157) <= not(layer1_outputs(3615));
    layer2_outputs(1158) <= '0';
    layer2_outputs(1159) <= '1';
    layer2_outputs(1160) <= '1';
    layer2_outputs(1161) <= not(layer1_outputs(3521));
    layer2_outputs(1162) <= '0';
    layer2_outputs(1163) <= not(layer1_outputs(4728));
    layer2_outputs(1164) <= (layer1_outputs(2200)) or (layer1_outputs(2750));
    layer2_outputs(1165) <= layer1_outputs(4239);
    layer2_outputs(1166) <= (layer1_outputs(4507)) and not (layer1_outputs(4754));
    layer2_outputs(1167) <= '1';
    layer2_outputs(1168) <= '0';
    layer2_outputs(1169) <= layer1_outputs(2368);
    layer2_outputs(1170) <= (layer1_outputs(1651)) or (layer1_outputs(1824));
    layer2_outputs(1171) <= '0';
    layer2_outputs(1172) <= layer1_outputs(3154);
    layer2_outputs(1173) <= (layer1_outputs(2609)) and not (layer1_outputs(4993));
    layer2_outputs(1174) <= not((layer1_outputs(4383)) and (layer1_outputs(4571)));
    layer2_outputs(1175) <= not((layer1_outputs(3365)) and (layer1_outputs(864)));
    layer2_outputs(1176) <= '1';
    layer2_outputs(1177) <= '0';
    layer2_outputs(1178) <= '0';
    layer2_outputs(1179) <= layer1_outputs(1449);
    layer2_outputs(1180) <= not((layer1_outputs(3525)) or (layer1_outputs(879)));
    layer2_outputs(1181) <= not(layer1_outputs(32)) or (layer1_outputs(4721));
    layer2_outputs(1182) <= not((layer1_outputs(4593)) or (layer1_outputs(3672)));
    layer2_outputs(1183) <= not(layer1_outputs(3518)) or (layer1_outputs(3594));
    layer2_outputs(1184) <= not(layer1_outputs(511));
    layer2_outputs(1185) <= layer1_outputs(3198);
    layer2_outputs(1186) <= (layer1_outputs(4708)) and not (layer1_outputs(400));
    layer2_outputs(1187) <= not(layer1_outputs(3302));
    layer2_outputs(1188) <= not(layer1_outputs(1310));
    layer2_outputs(1189) <= not(layer1_outputs(1461));
    layer2_outputs(1190) <= not((layer1_outputs(4177)) and (layer1_outputs(1578)));
    layer2_outputs(1191) <= not(layer1_outputs(3527)) or (layer1_outputs(2568));
    layer2_outputs(1192) <= not(layer1_outputs(1410)) or (layer1_outputs(2093));
    layer2_outputs(1193) <= layer1_outputs(5037);
    layer2_outputs(1194) <= '1';
    layer2_outputs(1195) <= '1';
    layer2_outputs(1196) <= (layer1_outputs(3499)) and not (layer1_outputs(3916));
    layer2_outputs(1197) <= not((layer1_outputs(2190)) and (layer1_outputs(2047)));
    layer2_outputs(1198) <= '0';
    layer2_outputs(1199) <= (layer1_outputs(4845)) and (layer1_outputs(939));
    layer2_outputs(1200) <= (layer1_outputs(2716)) and (layer1_outputs(1212));
    layer2_outputs(1201) <= not(layer1_outputs(1815));
    layer2_outputs(1202) <= not((layer1_outputs(4160)) and (layer1_outputs(3095)));
    layer2_outputs(1203) <= '0';
    layer2_outputs(1204) <= not(layer1_outputs(954));
    layer2_outputs(1205) <= '0';
    layer2_outputs(1206) <= not(layer1_outputs(3276)) or (layer1_outputs(4605));
    layer2_outputs(1207) <= not(layer1_outputs(1451)) or (layer1_outputs(2241));
    layer2_outputs(1208) <= not((layer1_outputs(2640)) xor (layer1_outputs(816)));
    layer2_outputs(1209) <= not((layer1_outputs(1341)) and (layer1_outputs(838)));
    layer2_outputs(1210) <= layer1_outputs(1594);
    layer2_outputs(1211) <= not(layer1_outputs(244));
    layer2_outputs(1212) <= (layer1_outputs(362)) and not (layer1_outputs(2924));
    layer2_outputs(1213) <= (layer1_outputs(3338)) and (layer1_outputs(2781));
    layer2_outputs(1214) <= not((layer1_outputs(365)) or (layer1_outputs(3354)));
    layer2_outputs(1215) <= not(layer1_outputs(795)) or (layer1_outputs(3108));
    layer2_outputs(1216) <= '1';
    layer2_outputs(1217) <= not(layer1_outputs(4167)) or (layer1_outputs(1353));
    layer2_outputs(1218) <= '0';
    layer2_outputs(1219) <= not(layer1_outputs(578)) or (layer1_outputs(3284));
    layer2_outputs(1220) <= layer1_outputs(2410);
    layer2_outputs(1221) <= not(layer1_outputs(5111)) or (layer1_outputs(1179));
    layer2_outputs(1222) <= not(layer1_outputs(1081)) or (layer1_outputs(1087));
    layer2_outputs(1223) <= not(layer1_outputs(1974));
    layer2_outputs(1224) <= layer1_outputs(4824);
    layer2_outputs(1225) <= not((layer1_outputs(2344)) and (layer1_outputs(4164)));
    layer2_outputs(1226) <= not(layer1_outputs(2157)) or (layer1_outputs(3719));
    layer2_outputs(1227) <= layer1_outputs(916);
    layer2_outputs(1228) <= (layer1_outputs(1882)) and not (layer1_outputs(4945));
    layer2_outputs(1229) <= not((layer1_outputs(2362)) and (layer1_outputs(2819)));
    layer2_outputs(1230) <= (layer1_outputs(1496)) and not (layer1_outputs(3651));
    layer2_outputs(1231) <= not(layer1_outputs(3136));
    layer2_outputs(1232) <= not(layer1_outputs(69));
    layer2_outputs(1233) <= '1';
    layer2_outputs(1234) <= not(layer1_outputs(4937)) or (layer1_outputs(2956));
    layer2_outputs(1235) <= not(layer1_outputs(3957));
    layer2_outputs(1236) <= not(layer1_outputs(1938)) or (layer1_outputs(1208));
    layer2_outputs(1237) <= not((layer1_outputs(2210)) or (layer1_outputs(4369)));
    layer2_outputs(1238) <= not((layer1_outputs(3560)) and (layer1_outputs(1509)));
    layer2_outputs(1239) <= not((layer1_outputs(2063)) and (layer1_outputs(1045)));
    layer2_outputs(1240) <= not((layer1_outputs(3965)) and (layer1_outputs(4696)));
    layer2_outputs(1241) <= not((layer1_outputs(3611)) and (layer1_outputs(4624)));
    layer2_outputs(1242) <= not(layer1_outputs(2108));
    layer2_outputs(1243) <= '0';
    layer2_outputs(1244) <= (layer1_outputs(2663)) and not (layer1_outputs(550));
    layer2_outputs(1245) <= (layer1_outputs(4465)) or (layer1_outputs(1481));
    layer2_outputs(1246) <= layer1_outputs(1205);
    layer2_outputs(1247) <= not(layer1_outputs(3572));
    layer2_outputs(1248) <= layer1_outputs(2518);
    layer2_outputs(1249) <= not(layer1_outputs(3808));
    layer2_outputs(1250) <= '0';
    layer2_outputs(1251) <= layer1_outputs(3732);
    layer2_outputs(1252) <= not(layer1_outputs(1604));
    layer2_outputs(1253) <= '0';
    layer2_outputs(1254) <= not(layer1_outputs(183));
    layer2_outputs(1255) <= layer1_outputs(2108);
    layer2_outputs(1256) <= not(layer1_outputs(4802)) or (layer1_outputs(4644));
    layer2_outputs(1257) <= '1';
    layer2_outputs(1258) <= not(layer1_outputs(1132));
    layer2_outputs(1259) <= (layer1_outputs(2046)) and not (layer1_outputs(4006));
    layer2_outputs(1260) <= (layer1_outputs(2983)) and (layer1_outputs(2730));
    layer2_outputs(1261) <= '0';
    layer2_outputs(1262) <= not(layer1_outputs(4535)) or (layer1_outputs(1741));
    layer2_outputs(1263) <= (layer1_outputs(4067)) and (layer1_outputs(3843));
    layer2_outputs(1264) <= '0';
    layer2_outputs(1265) <= layer1_outputs(4834);
    layer2_outputs(1266) <= (layer1_outputs(84)) and (layer1_outputs(4991));
    layer2_outputs(1267) <= not((layer1_outputs(2188)) or (layer1_outputs(295)));
    layer2_outputs(1268) <= not(layer1_outputs(4428)) or (layer1_outputs(846));
    layer2_outputs(1269) <= not(layer1_outputs(4169)) or (layer1_outputs(4309));
    layer2_outputs(1270) <= '1';
    layer2_outputs(1271) <= '0';
    layer2_outputs(1272) <= not(layer1_outputs(1271));
    layer2_outputs(1273) <= '0';
    layer2_outputs(1274) <= not(layer1_outputs(3274)) or (layer1_outputs(1251));
    layer2_outputs(1275) <= '0';
    layer2_outputs(1276) <= not((layer1_outputs(4944)) and (layer1_outputs(1954)));
    layer2_outputs(1277) <= (layer1_outputs(2680)) or (layer1_outputs(3301));
    layer2_outputs(1278) <= (layer1_outputs(1900)) and not (layer1_outputs(2466));
    layer2_outputs(1279) <= not(layer1_outputs(2164));
    layer2_outputs(1280) <= not(layer1_outputs(4858));
    layer2_outputs(1281) <= '1';
    layer2_outputs(1282) <= layer1_outputs(2881);
    layer2_outputs(1283) <= not(layer1_outputs(3096)) or (layer1_outputs(3473));
    layer2_outputs(1284) <= layer1_outputs(4447);
    layer2_outputs(1285) <= not(layer1_outputs(3310)) or (layer1_outputs(974));
    layer2_outputs(1286) <= (layer1_outputs(1855)) and (layer1_outputs(3023));
    layer2_outputs(1287) <= layer1_outputs(965);
    layer2_outputs(1288) <= '1';
    layer2_outputs(1289) <= '0';
    layer2_outputs(1290) <= '1';
    layer2_outputs(1291) <= (layer1_outputs(169)) or (layer1_outputs(4396));
    layer2_outputs(1292) <= (layer1_outputs(4287)) or (layer1_outputs(1056));
    layer2_outputs(1293) <= not((layer1_outputs(1358)) or (layer1_outputs(126)));
    layer2_outputs(1294) <= not((layer1_outputs(277)) and (layer1_outputs(2522)));
    layer2_outputs(1295) <= (layer1_outputs(1524)) and not (layer1_outputs(1326));
    layer2_outputs(1296) <= not((layer1_outputs(280)) or (layer1_outputs(4308)));
    layer2_outputs(1297) <= '1';
    layer2_outputs(1298) <= layer1_outputs(971);
    layer2_outputs(1299) <= not(layer1_outputs(54)) or (layer1_outputs(1102));
    layer2_outputs(1300) <= (layer1_outputs(2263)) and not (layer1_outputs(1387));
    layer2_outputs(1301) <= layer1_outputs(4154);
    layer2_outputs(1302) <= (layer1_outputs(209)) or (layer1_outputs(4021));
    layer2_outputs(1303) <= not((layer1_outputs(3245)) or (layer1_outputs(4885)));
    layer2_outputs(1304) <= not(layer1_outputs(1674));
    layer2_outputs(1305) <= layer1_outputs(3482);
    layer2_outputs(1306) <= (layer1_outputs(3834)) and not (layer1_outputs(3058));
    layer2_outputs(1307) <= layer1_outputs(256);
    layer2_outputs(1308) <= (layer1_outputs(1915)) and (layer1_outputs(4339));
    layer2_outputs(1309) <= not(layer1_outputs(652)) or (layer1_outputs(3561));
    layer2_outputs(1310) <= '1';
    layer2_outputs(1311) <= (layer1_outputs(4046)) and not (layer1_outputs(4027));
    layer2_outputs(1312) <= not(layer1_outputs(4990));
    layer2_outputs(1313) <= (layer1_outputs(4303)) and not (layer1_outputs(714));
    layer2_outputs(1314) <= '0';
    layer2_outputs(1315) <= (layer1_outputs(4973)) and not (layer1_outputs(5034));
    layer2_outputs(1316) <= not(layer1_outputs(4014));
    layer2_outputs(1317) <= layer1_outputs(161);
    layer2_outputs(1318) <= '0';
    layer2_outputs(1319) <= not(layer1_outputs(2516));
    layer2_outputs(1320) <= (layer1_outputs(1089)) and (layer1_outputs(4385));
    layer2_outputs(1321) <= (layer1_outputs(2042)) and (layer1_outputs(2464));
    layer2_outputs(1322) <= '1';
    layer2_outputs(1323) <= not(layer1_outputs(3738)) or (layer1_outputs(4229));
    layer2_outputs(1324) <= '0';
    layer2_outputs(1325) <= not(layer1_outputs(3769));
    layer2_outputs(1326) <= (layer1_outputs(3695)) and not (layer1_outputs(635));
    layer2_outputs(1327) <= not(layer1_outputs(2043));
    layer2_outputs(1328) <= (layer1_outputs(5039)) or (layer1_outputs(3494));
    layer2_outputs(1329) <= (layer1_outputs(488)) or (layer1_outputs(3289));
    layer2_outputs(1330) <= (layer1_outputs(2081)) and (layer1_outputs(4047));
    layer2_outputs(1331) <= layer1_outputs(2391);
    layer2_outputs(1332) <= not(layer1_outputs(3873)) or (layer1_outputs(476));
    layer2_outputs(1333) <= '0';
    layer2_outputs(1334) <= not(layer1_outputs(312)) or (layer1_outputs(167));
    layer2_outputs(1335) <= '0';
    layer2_outputs(1336) <= (layer1_outputs(3570)) or (layer1_outputs(3590));
    layer2_outputs(1337) <= not(layer1_outputs(1661)) or (layer1_outputs(938));
    layer2_outputs(1338) <= not(layer1_outputs(744));
    layer2_outputs(1339) <= '0';
    layer2_outputs(1340) <= layer1_outputs(423);
    layer2_outputs(1341) <= '1';
    layer2_outputs(1342) <= '1';
    layer2_outputs(1343) <= not(layer1_outputs(2218));
    layer2_outputs(1344) <= not((layer1_outputs(2523)) and (layer1_outputs(2735)));
    layer2_outputs(1345) <= not((layer1_outputs(1711)) and (layer1_outputs(3415)));
    layer2_outputs(1346) <= (layer1_outputs(4550)) and (layer1_outputs(1752));
    layer2_outputs(1347) <= (layer1_outputs(2312)) and not (layer1_outputs(2289));
    layer2_outputs(1348) <= (layer1_outputs(4876)) and not (layer1_outputs(2300));
    layer2_outputs(1349) <= not(layer1_outputs(4972)) or (layer1_outputs(4652));
    layer2_outputs(1350) <= (layer1_outputs(680)) and not (layer1_outputs(3874));
    layer2_outputs(1351) <= '0';
    layer2_outputs(1352) <= (layer1_outputs(2982)) and (layer1_outputs(3386));
    layer2_outputs(1353) <= '1';
    layer2_outputs(1354) <= (layer1_outputs(3156)) and not (layer1_outputs(4025));
    layer2_outputs(1355) <= '0';
    layer2_outputs(1356) <= (layer1_outputs(110)) and not (layer1_outputs(2114));
    layer2_outputs(1357) <= not(layer1_outputs(283));
    layer2_outputs(1358) <= not(layer1_outputs(719));
    layer2_outputs(1359) <= layer1_outputs(4204);
    layer2_outputs(1360) <= not(layer1_outputs(4034)) or (layer1_outputs(3489));
    layer2_outputs(1361) <= not(layer1_outputs(2815));
    layer2_outputs(1362) <= not(layer1_outputs(1704)) or (layer1_outputs(1745));
    layer2_outputs(1363) <= '1';
    layer2_outputs(1364) <= '1';
    layer2_outputs(1365) <= layer1_outputs(2368);
    layer2_outputs(1366) <= (layer1_outputs(2060)) xor (layer1_outputs(2991));
    layer2_outputs(1367) <= '1';
    layer2_outputs(1368) <= not(layer1_outputs(5064)) or (layer1_outputs(2707));
    layer2_outputs(1369) <= not((layer1_outputs(2376)) or (layer1_outputs(555)));
    layer2_outputs(1370) <= not(layer1_outputs(4526)) or (layer1_outputs(2671));
    layer2_outputs(1371) <= not(layer1_outputs(1603)) or (layer1_outputs(3477));
    layer2_outputs(1372) <= '0';
    layer2_outputs(1373) <= (layer1_outputs(5082)) and not (layer1_outputs(1430));
    layer2_outputs(1374) <= layer1_outputs(2500);
    layer2_outputs(1375) <= (layer1_outputs(4551)) and not (layer1_outputs(1742));
    layer2_outputs(1376) <= (layer1_outputs(1605)) and not (layer1_outputs(3509));
    layer2_outputs(1377) <= (layer1_outputs(986)) or (layer1_outputs(3627));
    layer2_outputs(1378) <= not(layer1_outputs(2758));
    layer2_outputs(1379) <= (layer1_outputs(2141)) or (layer1_outputs(1731));
    layer2_outputs(1380) <= '1';
    layer2_outputs(1381) <= (layer1_outputs(958)) and not (layer1_outputs(4583));
    layer2_outputs(1382) <= not(layer1_outputs(4057));
    layer2_outputs(1383) <= not(layer1_outputs(520)) or (layer1_outputs(4212));
    layer2_outputs(1384) <= (layer1_outputs(4692)) and (layer1_outputs(1447));
    layer2_outputs(1385) <= not((layer1_outputs(3434)) or (layer1_outputs(788)));
    layer2_outputs(1386) <= layer1_outputs(4506);
    layer2_outputs(1387) <= not((layer1_outputs(19)) and (layer1_outputs(262)));
    layer2_outputs(1388) <= not(layer1_outputs(1083));
    layer2_outputs(1389) <= layer1_outputs(508);
    layer2_outputs(1390) <= layer1_outputs(3914);
    layer2_outputs(1391) <= not(layer1_outputs(1283)) or (layer1_outputs(1489));
    layer2_outputs(1392) <= (layer1_outputs(988)) and not (layer1_outputs(4062));
    layer2_outputs(1393) <= '0';
    layer2_outputs(1394) <= (layer1_outputs(2074)) and not (layer1_outputs(2506));
    layer2_outputs(1395) <= not((layer1_outputs(4705)) or (layer1_outputs(72)));
    layer2_outputs(1396) <= (layer1_outputs(1983)) and (layer1_outputs(335));
    layer2_outputs(1397) <= (layer1_outputs(4532)) and not (layer1_outputs(2734));
    layer2_outputs(1398) <= '0';
    layer2_outputs(1399) <= layer1_outputs(885);
    layer2_outputs(1400) <= '1';
    layer2_outputs(1401) <= not((layer1_outputs(4698)) and (layer1_outputs(3384)));
    layer2_outputs(1402) <= not((layer1_outputs(4174)) or (layer1_outputs(4353)));
    layer2_outputs(1403) <= (layer1_outputs(3013)) and not (layer1_outputs(2181));
    layer2_outputs(1404) <= (layer1_outputs(3264)) or (layer1_outputs(1879));
    layer2_outputs(1405) <= (layer1_outputs(4913)) or (layer1_outputs(2450));
    layer2_outputs(1406) <= not(layer1_outputs(697));
    layer2_outputs(1407) <= not(layer1_outputs(1113));
    layer2_outputs(1408) <= not(layer1_outputs(3337)) or (layer1_outputs(766));
    layer2_outputs(1409) <= not((layer1_outputs(2265)) or (layer1_outputs(3066)));
    layer2_outputs(1410) <= (layer1_outputs(2065)) or (layer1_outputs(413));
    layer2_outputs(1411) <= (layer1_outputs(3765)) and not (layer1_outputs(2470));
    layer2_outputs(1412) <= not(layer1_outputs(2920)) or (layer1_outputs(4108));
    layer2_outputs(1413) <= '1';
    layer2_outputs(1414) <= layer1_outputs(4750);
    layer2_outputs(1415) <= (layer1_outputs(334)) and not (layer1_outputs(4114));
    layer2_outputs(1416) <= (layer1_outputs(504)) and not (layer1_outputs(4852));
    layer2_outputs(1417) <= '0';
    layer2_outputs(1418) <= not((layer1_outputs(797)) and (layer1_outputs(1767)));
    layer2_outputs(1419) <= not(layer1_outputs(2688));
    layer2_outputs(1420) <= layer1_outputs(917);
    layer2_outputs(1421) <= layer1_outputs(3847);
    layer2_outputs(1422) <= not((layer1_outputs(2321)) or (layer1_outputs(928)));
    layer2_outputs(1423) <= (layer1_outputs(2805)) and (layer1_outputs(2592));
    layer2_outputs(1424) <= '1';
    layer2_outputs(1425) <= not(layer1_outputs(4064)) or (layer1_outputs(4242));
    layer2_outputs(1426) <= not(layer1_outputs(3034)) or (layer1_outputs(3600));
    layer2_outputs(1427) <= layer1_outputs(3737);
    layer2_outputs(1428) <= (layer1_outputs(1190)) and (layer1_outputs(79));
    layer2_outputs(1429) <= (layer1_outputs(3906)) and (layer1_outputs(772));
    layer2_outputs(1430) <= not(layer1_outputs(1809)) or (layer1_outputs(4486));
    layer2_outputs(1431) <= layer1_outputs(2357);
    layer2_outputs(1432) <= '1';
    layer2_outputs(1433) <= not((layer1_outputs(4780)) and (layer1_outputs(852)));
    layer2_outputs(1434) <= (layer1_outputs(369)) or (layer1_outputs(2453));
    layer2_outputs(1435) <= (layer1_outputs(1051)) and (layer1_outputs(4315));
    layer2_outputs(1436) <= not(layer1_outputs(3621)) or (layer1_outputs(2051));
    layer2_outputs(1437) <= (layer1_outputs(1423)) and not (layer1_outputs(3751));
    layer2_outputs(1438) <= not((layer1_outputs(427)) and (layer1_outputs(3630)));
    layer2_outputs(1439) <= '0';
    layer2_outputs(1440) <= (layer1_outputs(1099)) and (layer1_outputs(285));
    layer2_outputs(1441) <= not(layer1_outputs(1396));
    layer2_outputs(1442) <= not(layer1_outputs(1254)) or (layer1_outputs(3158));
    layer2_outputs(1443) <= (layer1_outputs(4462)) and not (layer1_outputs(3203));
    layer2_outputs(1444) <= (layer1_outputs(3959)) or (layer1_outputs(4112));
    layer2_outputs(1445) <= not(layer1_outputs(2554)) or (layer1_outputs(3570));
    layer2_outputs(1446) <= not((layer1_outputs(3593)) xor (layer1_outputs(4524)));
    layer2_outputs(1447) <= (layer1_outputs(1962)) and not (layer1_outputs(451));
    layer2_outputs(1448) <= '1';
    layer2_outputs(1449) <= not(layer1_outputs(2541)) or (layer1_outputs(4665));
    layer2_outputs(1450) <= '1';
    layer2_outputs(1451) <= (layer1_outputs(2789)) and not (layer1_outputs(1082));
    layer2_outputs(1452) <= not((layer1_outputs(820)) and (layer1_outputs(91)));
    layer2_outputs(1453) <= (layer1_outputs(2478)) and not (layer1_outputs(3677));
    layer2_outputs(1454) <= not(layer1_outputs(832));
    layer2_outputs(1455) <= layer1_outputs(342);
    layer2_outputs(1456) <= (layer1_outputs(1064)) or (layer1_outputs(4567));
    layer2_outputs(1457) <= (layer1_outputs(4227)) and not (layer1_outputs(924));
    layer2_outputs(1458) <= not(layer1_outputs(3251)) or (layer1_outputs(2714));
    layer2_outputs(1459) <= (layer1_outputs(2029)) and not (layer1_outputs(2589));
    layer2_outputs(1460) <= not(layer1_outputs(1279)) or (layer1_outputs(3682));
    layer2_outputs(1461) <= not(layer1_outputs(1443));
    layer2_outputs(1462) <= not((layer1_outputs(3879)) and (layer1_outputs(4047)));
    layer2_outputs(1463) <= (layer1_outputs(2695)) and (layer1_outputs(1080));
    layer2_outputs(1464) <= not(layer1_outputs(4075));
    layer2_outputs(1465) <= (layer1_outputs(3378)) and not (layer1_outputs(1469));
    layer2_outputs(1466) <= not(layer1_outputs(4237));
    layer2_outputs(1467) <= not(layer1_outputs(4921));
    layer2_outputs(1468) <= not(layer1_outputs(3932));
    layer2_outputs(1469) <= layer1_outputs(1103);
    layer2_outputs(1470) <= not(layer1_outputs(1794)) or (layer1_outputs(4980));
    layer2_outputs(1471) <= not(layer1_outputs(4157)) or (layer1_outputs(1428));
    layer2_outputs(1472) <= not((layer1_outputs(3412)) or (layer1_outputs(3364)));
    layer2_outputs(1473) <= not((layer1_outputs(1488)) and (layer1_outputs(13)));
    layer2_outputs(1474) <= '1';
    layer2_outputs(1475) <= not(layer1_outputs(3529));
    layer2_outputs(1476) <= not(layer1_outputs(4640)) or (layer1_outputs(3110));
    layer2_outputs(1477) <= (layer1_outputs(2469)) and not (layer1_outputs(5071));
    layer2_outputs(1478) <= '1';
    layer2_outputs(1479) <= '1';
    layer2_outputs(1480) <= not(layer1_outputs(4965)) or (layer1_outputs(2013));
    layer2_outputs(1481) <= not(layer1_outputs(238));
    layer2_outputs(1482) <= (layer1_outputs(800)) and not (layer1_outputs(4949));
    layer2_outputs(1483) <= (layer1_outputs(2279)) and not (layer1_outputs(3143));
    layer2_outputs(1484) <= (layer1_outputs(601)) and not (layer1_outputs(2381));
    layer2_outputs(1485) <= (layer1_outputs(3844)) and not (layer1_outputs(458));
    layer2_outputs(1486) <= '0';
    layer2_outputs(1487) <= (layer1_outputs(510)) and not (layer1_outputs(3539));
    layer2_outputs(1488) <= not(layer1_outputs(1309)) or (layer1_outputs(3736));
    layer2_outputs(1489) <= not((layer1_outputs(4164)) and (layer1_outputs(4839)));
    layer2_outputs(1490) <= not(layer1_outputs(3402)) or (layer1_outputs(1399));
    layer2_outputs(1491) <= '1';
    layer2_outputs(1492) <= (layer1_outputs(3026)) and (layer1_outputs(1827));
    layer2_outputs(1493) <= not(layer1_outputs(2599));
    layer2_outputs(1494) <= layer1_outputs(3481);
    layer2_outputs(1495) <= (layer1_outputs(4618)) xor (layer1_outputs(2859));
    layer2_outputs(1496) <= not(layer1_outputs(933)) or (layer1_outputs(2887));
    layer2_outputs(1497) <= '0';
    layer2_outputs(1498) <= (layer1_outputs(1992)) and not (layer1_outputs(726));
    layer2_outputs(1499) <= not((layer1_outputs(99)) xor (layer1_outputs(4183)));
    layer2_outputs(1500) <= not(layer1_outputs(3339));
    layer2_outputs(1501) <= '1';
    layer2_outputs(1502) <= (layer1_outputs(4070)) and not (layer1_outputs(88));
    layer2_outputs(1503) <= (layer1_outputs(3901)) and not (layer1_outputs(650));
    layer2_outputs(1504) <= '0';
    layer2_outputs(1505) <= not((layer1_outputs(1313)) and (layer1_outputs(4710)));
    layer2_outputs(1506) <= not(layer1_outputs(1945)) or (layer1_outputs(289));
    layer2_outputs(1507) <= not(layer1_outputs(1984)) or (layer1_outputs(1065));
    layer2_outputs(1508) <= (layer1_outputs(1498)) or (layer1_outputs(243));
    layer2_outputs(1509) <= (layer1_outputs(4777)) and (layer1_outputs(2607));
    layer2_outputs(1510) <= not(layer1_outputs(3713)) or (layer1_outputs(232));
    layer2_outputs(1511) <= layer1_outputs(2612);
    layer2_outputs(1512) <= '0';
    layer2_outputs(1513) <= not(layer1_outputs(2264));
    layer2_outputs(1514) <= not(layer1_outputs(1124));
    layer2_outputs(1515) <= '0';
    layer2_outputs(1516) <= layer1_outputs(2190);
    layer2_outputs(1517) <= (layer1_outputs(1297)) and (layer1_outputs(1520));
    layer2_outputs(1518) <= not(layer1_outputs(3726)) or (layer1_outputs(815));
    layer2_outputs(1519) <= (layer1_outputs(4591)) or (layer1_outputs(496));
    layer2_outputs(1520) <= '0';
    layer2_outputs(1521) <= '0';
    layer2_outputs(1522) <= not(layer1_outputs(2416)) or (layer1_outputs(2813));
    layer2_outputs(1523) <= '0';
    layer2_outputs(1524) <= (layer1_outputs(2635)) or (layer1_outputs(4828));
    layer2_outputs(1525) <= (layer1_outputs(3146)) or (layer1_outputs(1768));
    layer2_outputs(1526) <= '0';
    layer2_outputs(1527) <= not(layer1_outputs(1127)) or (layer1_outputs(4487));
    layer2_outputs(1528) <= not(layer1_outputs(2511));
    layer2_outputs(1529) <= not(layer1_outputs(3167));
    layer2_outputs(1530) <= (layer1_outputs(3496)) and (layer1_outputs(4612));
    layer2_outputs(1531) <= (layer1_outputs(834)) and not (layer1_outputs(1835));
    layer2_outputs(1532) <= (layer1_outputs(145)) or (layer1_outputs(2764));
    layer2_outputs(1533) <= layer1_outputs(2006);
    layer2_outputs(1534) <= layer1_outputs(2822);
    layer2_outputs(1535) <= layer1_outputs(3628);
    layer2_outputs(1536) <= (layer1_outputs(2626)) or (layer1_outputs(4324));
    layer2_outputs(1537) <= (layer1_outputs(2448)) and not (layer1_outputs(3778));
    layer2_outputs(1538) <= (layer1_outputs(90)) or (layer1_outputs(1715));
    layer2_outputs(1539) <= not(layer1_outputs(1567)) or (layer1_outputs(2389));
    layer2_outputs(1540) <= not((layer1_outputs(2358)) and (layer1_outputs(3228)));
    layer2_outputs(1541) <= not(layer1_outputs(1874));
    layer2_outputs(1542) <= not(layer1_outputs(2217));
    layer2_outputs(1543) <= not(layer1_outputs(3036)) or (layer1_outputs(1215));
    layer2_outputs(1544) <= not(layer1_outputs(4739)) or (layer1_outputs(785));
    layer2_outputs(1545) <= (layer1_outputs(190)) and (layer1_outputs(3007));
    layer2_outputs(1546) <= not((layer1_outputs(2254)) or (layer1_outputs(3438)));
    layer2_outputs(1547) <= not((layer1_outputs(2337)) or (layer1_outputs(2253)));
    layer2_outputs(1548) <= not(layer1_outputs(2303)) or (layer1_outputs(3239));
    layer2_outputs(1549) <= not(layer1_outputs(634)) or (layer1_outputs(2842));
    layer2_outputs(1550) <= (layer1_outputs(3894)) and not (layer1_outputs(3460));
    layer2_outputs(1551) <= not((layer1_outputs(2746)) and (layer1_outputs(2682)));
    layer2_outputs(1552) <= '1';
    layer2_outputs(1553) <= '0';
    layer2_outputs(1554) <= not((layer1_outputs(4176)) or (layer1_outputs(4495)));
    layer2_outputs(1555) <= not(layer1_outputs(4715));
    layer2_outputs(1556) <= not((layer1_outputs(1697)) and (layer1_outputs(126)));
    layer2_outputs(1557) <= layer1_outputs(3526);
    layer2_outputs(1558) <= not(layer1_outputs(1134));
    layer2_outputs(1559) <= '1';
    layer2_outputs(1560) <= layer1_outputs(998);
    layer2_outputs(1561) <= (layer1_outputs(2900)) or (layer1_outputs(1696));
    layer2_outputs(1562) <= (layer1_outputs(340)) and not (layer1_outputs(4917));
    layer2_outputs(1563) <= not(layer1_outputs(3743)) or (layer1_outputs(2961));
    layer2_outputs(1564) <= not((layer1_outputs(3213)) xor (layer1_outputs(3151)));
    layer2_outputs(1565) <= not((layer1_outputs(525)) xor (layer1_outputs(4626)));
    layer2_outputs(1566) <= not(layer1_outputs(765)) or (layer1_outputs(2247));
    layer2_outputs(1567) <= layer1_outputs(2861);
    layer2_outputs(1568) <= layer1_outputs(1071);
    layer2_outputs(1569) <= not((layer1_outputs(4615)) and (layer1_outputs(2151)));
    layer2_outputs(1570) <= layer1_outputs(4575);
    layer2_outputs(1571) <= (layer1_outputs(1622)) and (layer1_outputs(417));
    layer2_outputs(1572) <= not(layer1_outputs(2877)) or (layer1_outputs(3070));
    layer2_outputs(1573) <= not(layer1_outputs(4675)) or (layer1_outputs(115));
    layer2_outputs(1574) <= layer1_outputs(2497);
    layer2_outputs(1575) <= not(layer1_outputs(3886));
    layer2_outputs(1576) <= not((layer1_outputs(3951)) and (layer1_outputs(190)));
    layer2_outputs(1577) <= not(layer1_outputs(559)) or (layer1_outputs(2280));
    layer2_outputs(1578) <= (layer1_outputs(530)) and not (layer1_outputs(3387));
    layer2_outputs(1579) <= not(layer1_outputs(3872));
    layer2_outputs(1580) <= not(layer1_outputs(1842));
    layer2_outputs(1581) <= (layer1_outputs(1549)) or (layer1_outputs(1887));
    layer2_outputs(1582) <= '0';
    layer2_outputs(1583) <= not(layer1_outputs(4420));
    layer2_outputs(1584) <= '1';
    layer2_outputs(1585) <= '0';
    layer2_outputs(1586) <= (layer1_outputs(897)) and not (layer1_outputs(398));
    layer2_outputs(1587) <= not(layer1_outputs(2895));
    layer2_outputs(1588) <= not(layer1_outputs(2792));
    layer2_outputs(1589) <= '0';
    layer2_outputs(1590) <= (layer1_outputs(3053)) or (layer1_outputs(1987));
    layer2_outputs(1591) <= (layer1_outputs(1521)) or (layer1_outputs(1586));
    layer2_outputs(1592) <= not((layer1_outputs(3851)) and (layer1_outputs(4565)));
    layer2_outputs(1593) <= '0';
    layer2_outputs(1594) <= (layer1_outputs(3976)) and not (layer1_outputs(2713));
    layer2_outputs(1595) <= not(layer1_outputs(2473)) or (layer1_outputs(1056));
    layer2_outputs(1596) <= not((layer1_outputs(3069)) or (layer1_outputs(127)));
    layer2_outputs(1597) <= '1';
    layer2_outputs(1598) <= '0';
    layer2_outputs(1599) <= (layer1_outputs(653)) and not (layer1_outputs(2033));
    layer2_outputs(1600) <= layer1_outputs(3211);
    layer2_outputs(1601) <= layer1_outputs(22);
    layer2_outputs(1602) <= '0';
    layer2_outputs(1603) <= (layer1_outputs(3550)) and not (layer1_outputs(375));
    layer2_outputs(1604) <= not((layer1_outputs(4093)) and (layer1_outputs(4817)));
    layer2_outputs(1605) <= not((layer1_outputs(1671)) and (layer1_outputs(741)));
    layer2_outputs(1606) <= not(layer1_outputs(420)) or (layer1_outputs(2789));
    layer2_outputs(1607) <= (layer1_outputs(984)) and not (layer1_outputs(1671));
    layer2_outputs(1608) <= not(layer1_outputs(4337)) or (layer1_outputs(4901));
    layer2_outputs(1609) <= '1';
    layer2_outputs(1610) <= (layer1_outputs(3376)) and not (layer1_outputs(3582));
    layer2_outputs(1611) <= '0';
    layer2_outputs(1612) <= (layer1_outputs(560)) and not (layer1_outputs(3938));
    layer2_outputs(1613) <= '0';
    layer2_outputs(1614) <= not(layer1_outputs(2137)) or (layer1_outputs(4727));
    layer2_outputs(1615) <= not(layer1_outputs(2874));
    layer2_outputs(1616) <= '0';
    layer2_outputs(1617) <= '1';
    layer2_outputs(1618) <= '1';
    layer2_outputs(1619) <= (layer1_outputs(3800)) and not (layer1_outputs(3048));
    layer2_outputs(1620) <= '1';
    layer2_outputs(1621) <= not((layer1_outputs(4149)) and (layer1_outputs(2705)));
    layer2_outputs(1622) <= (layer1_outputs(3152)) and not (layer1_outputs(2435));
    layer2_outputs(1623) <= (layer1_outputs(2976)) and (layer1_outputs(3824));
    layer2_outputs(1624) <= '0';
    layer2_outputs(1625) <= not((layer1_outputs(2559)) and (layer1_outputs(640)));
    layer2_outputs(1626) <= (layer1_outputs(1687)) and not (layer1_outputs(2213));
    layer2_outputs(1627) <= (layer1_outputs(3193)) and (layer1_outputs(2623));
    layer2_outputs(1628) <= not(layer1_outputs(2338));
    layer2_outputs(1629) <= '0';
    layer2_outputs(1630) <= (layer1_outputs(2335)) and not (layer1_outputs(2101));
    layer2_outputs(1631) <= (layer1_outputs(5032)) and (layer1_outputs(2609));
    layer2_outputs(1632) <= not((layer1_outputs(2006)) or (layer1_outputs(1627)));
    layer2_outputs(1633) <= layer1_outputs(2110);
    layer2_outputs(1634) <= (layer1_outputs(257)) xor (layer1_outputs(27));
    layer2_outputs(1635) <= '0';
    layer2_outputs(1636) <= (layer1_outputs(481)) and not (layer1_outputs(103));
    layer2_outputs(1637) <= '0';
    layer2_outputs(1638) <= not((layer1_outputs(831)) and (layer1_outputs(71)));
    layer2_outputs(1639) <= not((layer1_outputs(3296)) and (layer1_outputs(2229)));
    layer2_outputs(1640) <= (layer1_outputs(2328)) and (layer1_outputs(1511));
    layer2_outputs(1641) <= not((layer1_outputs(645)) and (layer1_outputs(4582)));
    layer2_outputs(1642) <= (layer1_outputs(159)) and not (layer1_outputs(3819));
    layer2_outputs(1643) <= (layer1_outputs(450)) or (layer1_outputs(2851));
    layer2_outputs(1644) <= not((layer1_outputs(2598)) and (layer1_outputs(575)));
    layer2_outputs(1645) <= layer1_outputs(367);
    layer2_outputs(1646) <= not((layer1_outputs(2055)) and (layer1_outputs(1872)));
    layer2_outputs(1647) <= (layer1_outputs(3386)) and (layer1_outputs(2815));
    layer2_outputs(1648) <= (layer1_outputs(321)) or (layer1_outputs(489));
    layer2_outputs(1649) <= '1';
    layer2_outputs(1650) <= not(layer1_outputs(1607)) or (layer1_outputs(4879));
    layer2_outputs(1651) <= not(layer1_outputs(3911)) or (layer1_outputs(551));
    layer2_outputs(1652) <= '1';
    layer2_outputs(1653) <= layer1_outputs(4149);
    layer2_outputs(1654) <= '1';
    layer2_outputs(1655) <= (layer1_outputs(3887)) and (layer1_outputs(4198));
    layer2_outputs(1656) <= layer1_outputs(4460);
    layer2_outputs(1657) <= (layer1_outputs(3741)) or (layer1_outputs(677));
    layer2_outputs(1658) <= layer1_outputs(1221);
    layer2_outputs(1659) <= not((layer1_outputs(3391)) and (layer1_outputs(325)));
    layer2_outputs(1660) <= not((layer1_outputs(2005)) or (layer1_outputs(2123)));
    layer2_outputs(1661) <= not(layer1_outputs(4546));
    layer2_outputs(1662) <= not(layer1_outputs(2844));
    layer2_outputs(1663) <= (layer1_outputs(1790)) and not (layer1_outputs(3316));
    layer2_outputs(1664) <= '0';
    layer2_outputs(1665) <= (layer1_outputs(3277)) and (layer1_outputs(65));
    layer2_outputs(1666) <= '1';
    layer2_outputs(1667) <= (layer1_outputs(3949)) and not (layer1_outputs(3216));
    layer2_outputs(1668) <= (layer1_outputs(2860)) or (layer1_outputs(1059));
    layer2_outputs(1669) <= layer1_outputs(3192);
    layer2_outputs(1670) <= '1';
    layer2_outputs(1671) <= not(layer1_outputs(2988)) or (layer1_outputs(2613));
    layer2_outputs(1672) <= not(layer1_outputs(2856));
    layer2_outputs(1673) <= not((layer1_outputs(3854)) or (layer1_outputs(258)));
    layer2_outputs(1674) <= not((layer1_outputs(455)) or (layer1_outputs(4716)));
    layer2_outputs(1675) <= (layer1_outputs(5092)) and not (layer1_outputs(2347));
    layer2_outputs(1676) <= not(layer1_outputs(1941));
    layer2_outputs(1677) <= not((layer1_outputs(1632)) and (layer1_outputs(616)));
    layer2_outputs(1678) <= layer1_outputs(2909);
    layer2_outputs(1679) <= (layer1_outputs(4942)) and not (layer1_outputs(1939));
    layer2_outputs(1680) <= '1';
    layer2_outputs(1681) <= not(layer1_outputs(3710));
    layer2_outputs(1682) <= '0';
    layer2_outputs(1683) <= (layer1_outputs(3952)) and not (layer1_outputs(1159));
    layer2_outputs(1684) <= (layer1_outputs(1617)) or (layer1_outputs(4409));
    layer2_outputs(1685) <= '0';
    layer2_outputs(1686) <= not((layer1_outputs(1935)) or (layer1_outputs(2482)));
    layer2_outputs(1687) <= '1';
    layer2_outputs(1688) <= '1';
    layer2_outputs(1689) <= not(layer1_outputs(1529));
    layer2_outputs(1690) <= not((layer1_outputs(3029)) or (layer1_outputs(4934)));
    layer2_outputs(1691) <= not((layer1_outputs(5063)) and (layer1_outputs(131)));
    layer2_outputs(1692) <= (layer1_outputs(4819)) and not (layer1_outputs(909));
    layer2_outputs(1693) <= (layer1_outputs(5108)) or (layer1_outputs(4196));
    layer2_outputs(1694) <= not(layer1_outputs(1273)) or (layer1_outputs(2104));
    layer2_outputs(1695) <= not(layer1_outputs(2726));
    layer2_outputs(1696) <= '1';
    layer2_outputs(1697) <= layer1_outputs(2706);
    layer2_outputs(1698) <= not((layer1_outputs(612)) or (layer1_outputs(4478)));
    layer2_outputs(1699) <= '1';
    layer2_outputs(1700) <= layer1_outputs(1020);
    layer2_outputs(1701) <= not(layer1_outputs(2853)) or (layer1_outputs(2732));
    layer2_outputs(1702) <= not(layer1_outputs(755)) or (layer1_outputs(3187));
    layer2_outputs(1703) <= (layer1_outputs(2888)) or (layer1_outputs(5031));
    layer2_outputs(1704) <= not(layer1_outputs(2723));
    layer2_outputs(1705) <= not(layer1_outputs(2739));
    layer2_outputs(1706) <= '1';
    layer2_outputs(1707) <= (layer1_outputs(3978)) and (layer1_outputs(980));
    layer2_outputs(1708) <= not(layer1_outputs(2276)) or (layer1_outputs(1420));
    layer2_outputs(1709) <= layer1_outputs(5119);
    layer2_outputs(1710) <= (layer1_outputs(825)) or (layer1_outputs(3666));
    layer2_outputs(1711) <= '0';
    layer2_outputs(1712) <= (layer1_outputs(1443)) and not (layer1_outputs(2826));
    layer2_outputs(1713) <= layer1_outputs(2210);
    layer2_outputs(1714) <= not(layer1_outputs(2023));
    layer2_outputs(1715) <= not((layer1_outputs(3767)) or (layer1_outputs(2284)));
    layer2_outputs(1716) <= (layer1_outputs(2100)) and not (layer1_outputs(1294));
    layer2_outputs(1717) <= not(layer1_outputs(2363)) or (layer1_outputs(4684));
    layer2_outputs(1718) <= '1';
    layer2_outputs(1719) <= '0';
    layer2_outputs(1720) <= not(layer1_outputs(3291));
    layer2_outputs(1721) <= not(layer1_outputs(3014));
    layer2_outputs(1722) <= (layer1_outputs(1162)) and not (layer1_outputs(1367));
    layer2_outputs(1723) <= not(layer1_outputs(3285));
    layer2_outputs(1724) <= not(layer1_outputs(914)) or (layer1_outputs(46));
    layer2_outputs(1725) <= not(layer1_outputs(3410)) or (layer1_outputs(694));
    layer2_outputs(1726) <= layer1_outputs(2357);
    layer2_outputs(1727) <= '0';
    layer2_outputs(1728) <= (layer1_outputs(4310)) or (layer1_outputs(1532));
    layer2_outputs(1729) <= layer1_outputs(3566);
    layer2_outputs(1730) <= not(layer1_outputs(3259));
    layer2_outputs(1731) <= layer1_outputs(5112);
    layer2_outputs(1732) <= (layer1_outputs(2923)) or (layer1_outputs(1167));
    layer2_outputs(1733) <= not(layer1_outputs(2040)) or (layer1_outputs(1166));
    layer2_outputs(1734) <= layer1_outputs(3145);
    layer2_outputs(1735) <= not((layer1_outputs(2985)) or (layer1_outputs(4064)));
    layer2_outputs(1736) <= (layer1_outputs(161)) and not (layer1_outputs(1589));
    layer2_outputs(1737) <= '1';
    layer2_outputs(1738) <= not(layer1_outputs(3569)) or (layer1_outputs(4194));
    layer2_outputs(1739) <= layer1_outputs(4664);
    layer2_outputs(1740) <= (layer1_outputs(2349)) and not (layer1_outputs(3383));
    layer2_outputs(1741) <= '1';
    layer2_outputs(1742) <= '0';
    layer2_outputs(1743) <= (layer1_outputs(671)) xor (layer1_outputs(3424));
    layer2_outputs(1744) <= (layer1_outputs(653)) or (layer1_outputs(2139));
    layer2_outputs(1745) <= '1';
    layer2_outputs(1746) <= not(layer1_outputs(1301)) or (layer1_outputs(4787));
    layer2_outputs(1747) <= not((layer1_outputs(2574)) and (layer1_outputs(3215)));
    layer2_outputs(1748) <= '0';
    layer2_outputs(1749) <= layer1_outputs(2409);
    layer2_outputs(1750) <= (layer1_outputs(63)) and (layer1_outputs(2302));
    layer2_outputs(1751) <= '1';
    layer2_outputs(1752) <= (layer1_outputs(1125)) or (layer1_outputs(4078));
    layer2_outputs(1753) <= not(layer1_outputs(4392));
    layer2_outputs(1754) <= (layer1_outputs(3776)) and not (layer1_outputs(3653));
    layer2_outputs(1755) <= (layer1_outputs(3104)) and not (layer1_outputs(2212));
    layer2_outputs(1756) <= not(layer1_outputs(911));
    layer2_outputs(1757) <= (layer1_outputs(487)) or (layer1_outputs(3414));
    layer2_outputs(1758) <= '0';
    layer2_outputs(1759) <= (layer1_outputs(3050)) and (layer1_outputs(2163));
    layer2_outputs(1760) <= (layer1_outputs(2360)) and not (layer1_outputs(3447));
    layer2_outputs(1761) <= '0';
    layer2_outputs(1762) <= not(layer1_outputs(166)) or (layer1_outputs(1264));
    layer2_outputs(1763) <= '0';
    layer2_outputs(1764) <= not((layer1_outputs(3200)) and (layer1_outputs(3764)));
    layer2_outputs(1765) <= (layer1_outputs(3934)) and not (layer1_outputs(2772));
    layer2_outputs(1766) <= layer1_outputs(4266);
    layer2_outputs(1767) <= '0';
    layer2_outputs(1768) <= not(layer1_outputs(2011));
    layer2_outputs(1769) <= (layer1_outputs(4253)) or (layer1_outputs(4072));
    layer2_outputs(1770) <= layer1_outputs(4059);
    layer2_outputs(1771) <= (layer1_outputs(1799)) or (layer1_outputs(710));
    layer2_outputs(1772) <= not(layer1_outputs(4241)) or (layer1_outputs(2369));
    layer2_outputs(1773) <= not((layer1_outputs(236)) and (layer1_outputs(4983)));
    layer2_outputs(1774) <= (layer1_outputs(4272)) and not (layer1_outputs(78));
    layer2_outputs(1775) <= not(layer1_outputs(3028)) or (layer1_outputs(1247));
    layer2_outputs(1776) <= not(layer1_outputs(2786)) or (layer1_outputs(3270));
    layer2_outputs(1777) <= not((layer1_outputs(1256)) or (layer1_outputs(151)));
    layer2_outputs(1778) <= not(layer1_outputs(524));
    layer2_outputs(1779) <= (layer1_outputs(3963)) and not (layer1_outputs(3031));
    layer2_outputs(1780) <= not((layer1_outputs(2101)) and (layer1_outputs(3439)));
    layer2_outputs(1781) <= (layer1_outputs(2779)) or (layer1_outputs(3929));
    layer2_outputs(1782) <= (layer1_outputs(2208)) and not (layer1_outputs(1048));
    layer2_outputs(1783) <= layer1_outputs(2809);
    layer2_outputs(1784) <= layer1_outputs(2655);
    layer2_outputs(1785) <= not(layer1_outputs(502)) or (layer1_outputs(3124));
    layer2_outputs(1786) <= not(layer1_outputs(4904));
    layer2_outputs(1787) <= not(layer1_outputs(1079));
    layer2_outputs(1788) <= not(layer1_outputs(3645));
    layer2_outputs(1789) <= (layer1_outputs(1875)) and not (layer1_outputs(4823));
    layer2_outputs(1790) <= (layer1_outputs(3350)) and not (layer1_outputs(2127));
    layer2_outputs(1791) <= '1';
    layer2_outputs(1792) <= not((layer1_outputs(2298)) and (layer1_outputs(3685)));
    layer2_outputs(1793) <= (layer1_outputs(2021)) and not (layer1_outputs(4405));
    layer2_outputs(1794) <= '1';
    layer2_outputs(1795) <= not((layer1_outputs(885)) or (layer1_outputs(2583)));
    layer2_outputs(1796) <= '1';
    layer2_outputs(1797) <= not(layer1_outputs(3548));
    layer2_outputs(1798) <= layer1_outputs(1932);
    layer2_outputs(1799) <= not(layer1_outputs(2862));
    layer2_outputs(1800) <= '0';
    layer2_outputs(1801) <= '1';
    layer2_outputs(1802) <= (layer1_outputs(4578)) and (layer1_outputs(3776));
    layer2_outputs(1803) <= not(layer1_outputs(373)) or (layer1_outputs(3599));
    layer2_outputs(1804) <= (layer1_outputs(3107)) and not (layer1_outputs(1682));
    layer2_outputs(1805) <= (layer1_outputs(1148)) and not (layer1_outputs(1160));
    layer2_outputs(1806) <= layer1_outputs(4969);
    layer2_outputs(1807) <= '0';
    layer2_outputs(1808) <= not((layer1_outputs(1654)) and (layer1_outputs(1554)));
    layer2_outputs(1809) <= (layer1_outputs(741)) xor (layer1_outputs(4632));
    layer2_outputs(1810) <= '0';
    layer2_outputs(1811) <= (layer1_outputs(3002)) or (layer1_outputs(1342));
    layer2_outputs(1812) <= (layer1_outputs(1123)) and not (layer1_outputs(3417));
    layer2_outputs(1813) <= (layer1_outputs(2990)) and (layer1_outputs(1370));
    layer2_outputs(1814) <= '1';
    layer2_outputs(1815) <= not(layer1_outputs(2189)) or (layer1_outputs(4463));
    layer2_outputs(1816) <= (layer1_outputs(1567)) or (layer1_outputs(2378));
    layer2_outputs(1817) <= (layer1_outputs(4371)) or (layer1_outputs(2980));
    layer2_outputs(1818) <= not(layer1_outputs(777));
    layer2_outputs(1819) <= not((layer1_outputs(1631)) or (layer1_outputs(369)));
    layer2_outputs(1820) <= (layer1_outputs(2555)) and not (layer1_outputs(338));
    layer2_outputs(1821) <= not(layer1_outputs(791)) or (layer1_outputs(952));
    layer2_outputs(1822) <= layer1_outputs(3122);
    layer2_outputs(1823) <= (layer1_outputs(2085)) or (layer1_outputs(3219));
    layer2_outputs(1824) <= (layer1_outputs(1001)) xor (layer1_outputs(3441));
    layer2_outputs(1825) <= '0';
    layer2_outputs(1826) <= not(layer1_outputs(3920)) or (layer1_outputs(1070));
    layer2_outputs(1827) <= '1';
    layer2_outputs(1828) <= not(layer1_outputs(2932));
    layer2_outputs(1829) <= not(layer1_outputs(1543)) or (layer1_outputs(4721));
    layer2_outputs(1830) <= (layer1_outputs(1524)) or (layer1_outputs(4479));
    layer2_outputs(1831) <= '0';
    layer2_outputs(1832) <= not(layer1_outputs(176));
    layer2_outputs(1833) <= not(layer1_outputs(4403));
    layer2_outputs(1834) <= not(layer1_outputs(1544));
    layer2_outputs(1835) <= (layer1_outputs(892)) and not (layer1_outputs(4694));
    layer2_outputs(1836) <= (layer1_outputs(4941)) and not (layer1_outputs(1878));
    layer2_outputs(1837) <= '0';
    layer2_outputs(1838) <= not(layer1_outputs(2663));
    layer2_outputs(1839) <= layer1_outputs(1878);
    layer2_outputs(1840) <= (layer1_outputs(915)) or (layer1_outputs(4576));
    layer2_outputs(1841) <= (layer1_outputs(1224)) and (layer1_outputs(4909));
    layer2_outputs(1842) <= (layer1_outputs(4957)) xor (layer1_outputs(3006));
    layer2_outputs(1843) <= (layer1_outputs(4809)) and (layer1_outputs(1544));
    layer2_outputs(1844) <= (layer1_outputs(3663)) and not (layer1_outputs(2929));
    layer2_outputs(1845) <= not((layer1_outputs(4724)) and (layer1_outputs(4032)));
    layer2_outputs(1846) <= not((layer1_outputs(333)) or (layer1_outputs(4448)));
    layer2_outputs(1847) <= not(layer1_outputs(4224));
    layer2_outputs(1848) <= (layer1_outputs(2493)) and not (layer1_outputs(255));
    layer2_outputs(1849) <= '0';
    layer2_outputs(1850) <= '1';
    layer2_outputs(1851) <= (layer1_outputs(1116)) xor (layer1_outputs(3701));
    layer2_outputs(1852) <= not(layer1_outputs(2935)) or (layer1_outputs(3194));
    layer2_outputs(1853) <= '0';
    layer2_outputs(1854) <= not(layer1_outputs(1330)) or (layer1_outputs(346));
    layer2_outputs(1855) <= (layer1_outputs(2910)) and not (layer1_outputs(2203));
    layer2_outputs(1856) <= (layer1_outputs(1369)) and not (layer1_outputs(459));
    layer2_outputs(1857) <= not(layer1_outputs(3305)) or (layer1_outputs(4634));
    layer2_outputs(1858) <= (layer1_outputs(1135)) and not (layer1_outputs(1301));
    layer2_outputs(1859) <= (layer1_outputs(2574)) or (layer1_outputs(3889));
    layer2_outputs(1860) <= not((layer1_outputs(850)) xor (layer1_outputs(1966)));
    layer2_outputs(1861) <= '1';
    layer2_outputs(1862) <= not((layer1_outputs(329)) or (layer1_outputs(3945)));
    layer2_outputs(1863) <= layer1_outputs(1895);
    layer2_outputs(1864) <= not(layer1_outputs(1209));
    layer2_outputs(1865) <= (layer1_outputs(3348)) and (layer1_outputs(2716));
    layer2_outputs(1866) <= not((layer1_outputs(3538)) xor (layer1_outputs(1845)));
    layer2_outputs(1867) <= (layer1_outputs(3860)) and (layer1_outputs(1884));
    layer2_outputs(1868) <= not(layer1_outputs(875)) or (layer1_outputs(2408));
    layer2_outputs(1869) <= '1';
    layer2_outputs(1870) <= not(layer1_outputs(2416)) or (layer1_outputs(2757));
    layer2_outputs(1871) <= (layer1_outputs(763)) and not (layer1_outputs(4977));
    layer2_outputs(1872) <= (layer1_outputs(76)) or (layer1_outputs(4931));
    layer2_outputs(1873) <= not((layer1_outputs(220)) and (layer1_outputs(6)));
    layer2_outputs(1874) <= '0';
    layer2_outputs(1875) <= (layer1_outputs(4152)) or (layer1_outputs(194));
    layer2_outputs(1876) <= (layer1_outputs(4712)) and not (layer1_outputs(1676));
    layer2_outputs(1877) <= layer1_outputs(4024);
    layer2_outputs(1878) <= '0';
    layer2_outputs(1879) <= '0';
    layer2_outputs(1880) <= not(layer1_outputs(2542)) or (layer1_outputs(3653));
    layer2_outputs(1881) <= (layer1_outputs(1244)) or (layer1_outputs(3946));
    layer2_outputs(1882) <= not((layer1_outputs(618)) or (layer1_outputs(337)));
    layer2_outputs(1883) <= not((layer1_outputs(2173)) and (layer1_outputs(1307)));
    layer2_outputs(1884) <= not(layer1_outputs(3681));
    layer2_outputs(1885) <= '1';
    layer2_outputs(1886) <= '0';
    layer2_outputs(1887) <= layer1_outputs(1222);
    layer2_outputs(1888) <= not((layer1_outputs(4794)) and (layer1_outputs(237)));
    layer2_outputs(1889) <= layer1_outputs(3383);
    layer2_outputs(1890) <= (layer1_outputs(861)) and (layer1_outputs(4276));
    layer2_outputs(1891) <= layer1_outputs(1783);
    layer2_outputs(1892) <= (layer1_outputs(2582)) and not (layer1_outputs(3754));
    layer2_outputs(1893) <= layer1_outputs(865);
    layer2_outputs(1894) <= (layer1_outputs(2254)) or (layer1_outputs(2657));
    layer2_outputs(1895) <= not(layer1_outputs(202)) or (layer1_outputs(3281));
    layer2_outputs(1896) <= not((layer1_outputs(464)) and (layer1_outputs(1713)));
    layer2_outputs(1897) <= '0';
    layer2_outputs(1898) <= '1';
    layer2_outputs(1899) <= '0';
    layer2_outputs(1900) <= layer1_outputs(4334);
    layer2_outputs(1901) <= (layer1_outputs(1315)) and not (layer1_outputs(60));
    layer2_outputs(1902) <= not((layer1_outputs(2470)) and (layer1_outputs(1774)));
    layer2_outputs(1903) <= '0';
    layer2_outputs(1904) <= not(layer1_outputs(876)) or (layer1_outputs(4836));
    layer2_outputs(1905) <= '1';
    layer2_outputs(1906) <= not((layer1_outputs(3646)) and (layer1_outputs(3207)));
    layer2_outputs(1907) <= not(layer1_outputs(2324)) or (layer1_outputs(4380));
    layer2_outputs(1908) <= '0';
    layer2_outputs(1909) <= (layer1_outputs(1207)) and (layer1_outputs(4430));
    layer2_outputs(1910) <= '1';
    layer2_outputs(1911) <= (layer1_outputs(531)) and (layer1_outputs(800));
    layer2_outputs(1912) <= not(layer1_outputs(1379)) or (layer1_outputs(5024));
    layer2_outputs(1913) <= not(layer1_outputs(1172));
    layer2_outputs(1914) <= not((layer1_outputs(2184)) and (layer1_outputs(5076)));
    layer2_outputs(1915) <= (layer1_outputs(769)) and not (layer1_outputs(4528));
    layer2_outputs(1916) <= not(layer1_outputs(29));
    layer2_outputs(1917) <= (layer1_outputs(3417)) or (layer1_outputs(1324));
    layer2_outputs(1918) <= (layer1_outputs(2071)) and not (layer1_outputs(4483));
    layer2_outputs(1919) <= '0';
    layer2_outputs(1920) <= not((layer1_outputs(2042)) xor (layer1_outputs(3983)));
    layer2_outputs(1921) <= (layer1_outputs(4558)) and not (layer1_outputs(3595));
    layer2_outputs(1922) <= (layer1_outputs(2222)) and not (layer1_outputs(3950));
    layer2_outputs(1923) <= not((layer1_outputs(1702)) or (layer1_outputs(1353)));
    layer2_outputs(1924) <= (layer1_outputs(2839)) and (layer1_outputs(3280));
    layer2_outputs(1925) <= not((layer1_outputs(710)) or (layer1_outputs(3554)));
    layer2_outputs(1926) <= (layer1_outputs(2756)) and (layer1_outputs(2367));
    layer2_outputs(1927) <= not(layer1_outputs(3483));
    layer2_outputs(1928) <= not(layer1_outputs(1709)) or (layer1_outputs(1618));
    layer2_outputs(1929) <= '1';
    layer2_outputs(1930) <= (layer1_outputs(2794)) and not (layer1_outputs(3089));
    layer2_outputs(1931) <= '1';
    layer2_outputs(1932) <= (layer1_outputs(1492)) or (layer1_outputs(2034));
    layer2_outputs(1933) <= layer1_outputs(3340);
    layer2_outputs(1934) <= not(layer1_outputs(4003)) or (layer1_outputs(1602));
    layer2_outputs(1935) <= not(layer1_outputs(4781)) or (layer1_outputs(4542));
    layer2_outputs(1936) <= '0';
    layer2_outputs(1937) <= not(layer1_outputs(4776)) or (layer1_outputs(3489));
    layer2_outputs(1938) <= '1';
    layer2_outputs(1939) <= not(layer1_outputs(3837));
    layer2_outputs(1940) <= not(layer1_outputs(1750));
    layer2_outputs(1941) <= not(layer1_outputs(594)) or (layer1_outputs(2803));
    layer2_outputs(1942) <= not(layer1_outputs(902)) or (layer1_outputs(4848));
    layer2_outputs(1943) <= '0';
    layer2_outputs(1944) <= layer1_outputs(3142);
    layer2_outputs(1945) <= not(layer1_outputs(1770));
    layer2_outputs(1946) <= '1';
    layer2_outputs(1947) <= not(layer1_outputs(1822)) or (layer1_outputs(1483));
    layer2_outputs(1948) <= not((layer1_outputs(3891)) and (layer1_outputs(310)));
    layer2_outputs(1949) <= '0';
    layer2_outputs(1950) <= layer1_outputs(4113);
    layer2_outputs(1951) <= layer1_outputs(3167);
    layer2_outputs(1952) <= not(layer1_outputs(3307));
    layer2_outputs(1953) <= not(layer1_outputs(5055)) or (layer1_outputs(899));
    layer2_outputs(1954) <= '0';
    layer2_outputs(1955) <= not(layer1_outputs(4803)) or (layer1_outputs(3639));
    layer2_outputs(1956) <= not((layer1_outputs(2044)) or (layer1_outputs(1543)));
    layer2_outputs(1957) <= not(layer1_outputs(844)) or (layer1_outputs(590));
    layer2_outputs(1958) <= not(layer1_outputs(3226)) or (layer1_outputs(4560));
    layer2_outputs(1959) <= layer1_outputs(4147);
    layer2_outputs(1960) <= layer1_outputs(4050);
    layer2_outputs(1961) <= not((layer1_outputs(4374)) or (layer1_outputs(4570)));
    layer2_outputs(1962) <= '1';
    layer2_outputs(1963) <= not((layer1_outputs(3279)) or (layer1_outputs(620)));
    layer2_outputs(1964) <= '1';
    layer2_outputs(1965) <= '0';
    layer2_outputs(1966) <= '0';
    layer2_outputs(1967) <= layer1_outputs(2855);
    layer2_outputs(1968) <= not(layer1_outputs(230)) or (layer1_outputs(3265));
    layer2_outputs(1969) <= not(layer1_outputs(705)) or (layer1_outputs(187));
    layer2_outputs(1970) <= not((layer1_outputs(4868)) and (layer1_outputs(2776)));
    layer2_outputs(1971) <= '1';
    layer2_outputs(1972) <= '0';
    layer2_outputs(1973) <= '1';
    layer2_outputs(1974) <= '0';
    layer2_outputs(1975) <= '0';
    layer2_outputs(1976) <= '1';
    layer2_outputs(1977) <= not((layer1_outputs(758)) and (layer1_outputs(910)));
    layer2_outputs(1978) <= not((layer1_outputs(541)) or (layer1_outputs(718)));
    layer2_outputs(1979) <= (layer1_outputs(4351)) and (layer1_outputs(4482));
    layer2_outputs(1980) <= layer1_outputs(4330);
    layer2_outputs(1981) <= '1';
    layer2_outputs(1982) <= (layer1_outputs(996)) and not (layer1_outputs(1023));
    layer2_outputs(1983) <= (layer1_outputs(1794)) and not (layer1_outputs(2964));
    layer2_outputs(1984) <= (layer1_outputs(3318)) or (layer1_outputs(599));
    layer2_outputs(1985) <= not(layer1_outputs(2622));
    layer2_outputs(1986) <= not(layer1_outputs(3506));
    layer2_outputs(1987) <= (layer1_outputs(1386)) and not (layer1_outputs(4478));
    layer2_outputs(1988) <= not(layer1_outputs(1996));
    layer2_outputs(1989) <= layer1_outputs(4692);
    layer2_outputs(1990) <= '0';
    layer2_outputs(1991) <= (layer1_outputs(2417)) and not (layer1_outputs(3523));
    layer2_outputs(1992) <= not((layer1_outputs(3429)) and (layer1_outputs(4360)));
    layer2_outputs(1993) <= (layer1_outputs(4127)) and not (layer1_outputs(1702));
    layer2_outputs(1994) <= not((layer1_outputs(3353)) and (layer1_outputs(3677)));
    layer2_outputs(1995) <= '1';
    layer2_outputs(1996) <= (layer1_outputs(3753)) and (layer1_outputs(3409));
    layer2_outputs(1997) <= not(layer1_outputs(4139));
    layer2_outputs(1998) <= not(layer1_outputs(738)) or (layer1_outputs(5095));
    layer2_outputs(1999) <= not(layer1_outputs(1410));
    layer2_outputs(2000) <= '1';
    layer2_outputs(2001) <= (layer1_outputs(5079)) and not (layer1_outputs(3139));
    layer2_outputs(2002) <= (layer1_outputs(2843)) and not (layer1_outputs(3408));
    layer2_outputs(2003) <= (layer1_outputs(4470)) and (layer1_outputs(2434));
    layer2_outputs(2004) <= not(layer1_outputs(2010));
    layer2_outputs(2005) <= not(layer1_outputs(2636)) or (layer1_outputs(178));
    layer2_outputs(2006) <= '1';
    layer2_outputs(2007) <= not(layer1_outputs(2556)) or (layer1_outputs(485));
    layer2_outputs(2008) <= (layer1_outputs(3157)) xor (layer1_outputs(4840));
    layer2_outputs(2009) <= not((layer1_outputs(1484)) or (layer1_outputs(736)));
    layer2_outputs(2010) <= layer1_outputs(2800);
    layer2_outputs(2011) <= not(layer1_outputs(1178)) or (layer1_outputs(3004));
    layer2_outputs(2012) <= layer1_outputs(3553);
    layer2_outputs(2013) <= '1';
    layer2_outputs(2014) <= '0';
    layer2_outputs(2015) <= not(layer1_outputs(3557)) or (layer1_outputs(3688));
    layer2_outputs(2016) <= '0';
    layer2_outputs(2017) <= not((layer1_outputs(4068)) xor (layer1_outputs(2091)));
    layer2_outputs(2018) <= (layer1_outputs(1209)) or (layer1_outputs(3400));
    layer2_outputs(2019) <= (layer1_outputs(4552)) or (layer1_outputs(3369));
    layer2_outputs(2020) <= (layer1_outputs(1441)) and not (layer1_outputs(4518));
    layer2_outputs(2021) <= not((layer1_outputs(2725)) xor (layer1_outputs(4085)));
    layer2_outputs(2022) <= not(layer1_outputs(1087)) or (layer1_outputs(2140));
    layer2_outputs(2023) <= not((layer1_outputs(1472)) or (layer1_outputs(182)));
    layer2_outputs(2024) <= (layer1_outputs(4272)) and (layer1_outputs(3721));
    layer2_outputs(2025) <= (layer1_outputs(2366)) or (layer1_outputs(850));
    layer2_outputs(2026) <= not(layer1_outputs(3591)) or (layer1_outputs(2866));
    layer2_outputs(2027) <= '1';
    layer2_outputs(2028) <= (layer1_outputs(3040)) or (layer1_outputs(552));
    layer2_outputs(2029) <= '1';
    layer2_outputs(2030) <= '0';
    layer2_outputs(2031) <= not(layer1_outputs(4084)) or (layer1_outputs(1288));
    layer2_outputs(2032) <= (layer1_outputs(5055)) and (layer1_outputs(2460));
    layer2_outputs(2033) <= layer1_outputs(1804);
    layer2_outputs(2034) <= not(layer1_outputs(2016));
    layer2_outputs(2035) <= not((layer1_outputs(3479)) or (layer1_outputs(3090)));
    layer2_outputs(2036) <= not((layer1_outputs(2600)) and (layer1_outputs(3442)));
    layer2_outputs(2037) <= not((layer1_outputs(1402)) and (layer1_outputs(4997)));
    layer2_outputs(2038) <= not(layer1_outputs(4826));
    layer2_outputs(2039) <= not((layer1_outputs(3998)) or (layer1_outputs(4416)));
    layer2_outputs(2040) <= '0';
    layer2_outputs(2041) <= '1';
    layer2_outputs(2042) <= '0';
    layer2_outputs(2043) <= '1';
    layer2_outputs(2044) <= layer1_outputs(1576);
    layer2_outputs(2045) <= (layer1_outputs(3096)) and not (layer1_outputs(1600));
    layer2_outputs(2046) <= not(layer1_outputs(1335));
    layer2_outputs(2047) <= layer1_outputs(549);
    layer2_outputs(2048) <= layer1_outputs(2418);
    layer2_outputs(2049) <= not((layer1_outputs(3448)) and (layer1_outputs(3977)));
    layer2_outputs(2050) <= not((layer1_outputs(1646)) or (layer1_outputs(3221)));
    layer2_outputs(2051) <= '0';
    layer2_outputs(2052) <= not((layer1_outputs(2926)) and (layer1_outputs(4844)));
    layer2_outputs(2053) <= '1';
    layer2_outputs(2054) <= not((layer1_outputs(380)) and (layer1_outputs(482)));
    layer2_outputs(2055) <= (layer1_outputs(3342)) or (layer1_outputs(4724));
    layer2_outputs(2056) <= '0';
    layer2_outputs(2057) <= '0';
    layer2_outputs(2058) <= '0';
    layer2_outputs(2059) <= '0';
    layer2_outputs(2060) <= (layer1_outputs(5093)) and not (layer1_outputs(1053));
    layer2_outputs(2061) <= (layer1_outputs(2916)) and not (layer1_outputs(3568));
    layer2_outputs(2062) <= not((layer1_outputs(2674)) and (layer1_outputs(4809)));
    layer2_outputs(2063) <= (layer1_outputs(98)) and not (layer1_outputs(559));
    layer2_outputs(2064) <= not((layer1_outputs(2004)) or (layer1_outputs(2584)));
    layer2_outputs(2065) <= layer1_outputs(45);
    layer2_outputs(2066) <= (layer1_outputs(1904)) and (layer1_outputs(2939));
    layer2_outputs(2067) <= layer1_outputs(1530);
    layer2_outputs(2068) <= '0';
    layer2_outputs(2069) <= not((layer1_outputs(3639)) or (layer1_outputs(4588)));
    layer2_outputs(2070) <= not((layer1_outputs(1735)) or (layer1_outputs(5056)));
    layer2_outputs(2071) <= not(layer1_outputs(2787));
    layer2_outputs(2072) <= not(layer1_outputs(1689));
    layer2_outputs(2073) <= not((layer1_outputs(3993)) or (layer1_outputs(3649)));
    layer2_outputs(2074) <= not(layer1_outputs(1058));
    layer2_outputs(2075) <= not((layer1_outputs(1308)) or (layer1_outputs(4004)));
    layer2_outputs(2076) <= (layer1_outputs(4402)) and not (layer1_outputs(2661));
    layer2_outputs(2077) <= (layer1_outputs(2579)) and (layer1_outputs(3591));
    layer2_outputs(2078) <= (layer1_outputs(1142)) and not (layer1_outputs(3924));
    layer2_outputs(2079) <= (layer1_outputs(1793)) and not (layer1_outputs(2343));
    layer2_outputs(2080) <= (layer1_outputs(1615)) or (layer1_outputs(3171));
    layer2_outputs(2081) <= not((layer1_outputs(3839)) and (layer1_outputs(3453)));
    layer2_outputs(2082) <= (layer1_outputs(3212)) and (layer1_outputs(1510));
    layer2_outputs(2083) <= (layer1_outputs(4675)) and not (layer1_outputs(4069));
    layer2_outputs(2084) <= not(layer1_outputs(1242)) or (layer1_outputs(553));
    layer2_outputs(2085) <= layer1_outputs(3691);
    layer2_outputs(2086) <= '0';
    layer2_outputs(2087) <= '0';
    layer2_outputs(2088) <= not(layer1_outputs(3214));
    layer2_outputs(2089) <= layer1_outputs(3829);
    layer2_outputs(2090) <= not(layer1_outputs(1340));
    layer2_outputs(2091) <= '0';
    layer2_outputs(2092) <= not(layer1_outputs(354));
    layer2_outputs(2093) <= not((layer1_outputs(986)) or (layer1_outputs(2236)));
    layer2_outputs(2094) <= (layer1_outputs(5100)) and not (layer1_outputs(3835));
    layer2_outputs(2095) <= not(layer1_outputs(1678));
    layer2_outputs(2096) <= (layer1_outputs(2522)) and (layer1_outputs(170));
    layer2_outputs(2097) <= not(layer1_outputs(4331));
    layer2_outputs(2098) <= '1';
    layer2_outputs(2099) <= not(layer1_outputs(2853));
    layer2_outputs(2100) <= '1';
    layer2_outputs(2101) <= '0';
    layer2_outputs(2102) <= not(layer1_outputs(132));
    layer2_outputs(2103) <= '1';
    layer2_outputs(2104) <= layer1_outputs(3086);
    layer2_outputs(2105) <= '0';
    layer2_outputs(2106) <= '0';
    layer2_outputs(2107) <= (layer1_outputs(505)) or (layer1_outputs(3919));
    layer2_outputs(2108) <= layer1_outputs(3819);
    layer2_outputs(2109) <= not((layer1_outputs(1652)) or (layer1_outputs(4032)));
    layer2_outputs(2110) <= '1';
    layer2_outputs(2111) <= not(layer1_outputs(4420)) or (layer1_outputs(4594));
    layer2_outputs(2112) <= (layer1_outputs(3080)) or (layer1_outputs(3220));
    layer2_outputs(2113) <= (layer1_outputs(4011)) or (layer1_outputs(4428));
    layer2_outputs(2114) <= not((layer1_outputs(4789)) and (layer1_outputs(49)));
    layer2_outputs(2115) <= '1';
    layer2_outputs(2116) <= not(layer1_outputs(1765));
    layer2_outputs(2117) <= not(layer1_outputs(2126));
    layer2_outputs(2118) <= (layer1_outputs(269)) and (layer1_outputs(2336));
    layer2_outputs(2119) <= (layer1_outputs(4325)) and not (layer1_outputs(4063));
    layer2_outputs(2120) <= layer1_outputs(627);
    layer2_outputs(2121) <= (layer1_outputs(2825)) and (layer1_outputs(3861));
    layer2_outputs(2122) <= not((layer1_outputs(1140)) and (layer1_outputs(3929)));
    layer2_outputs(2123) <= '1';
    layer2_outputs(2124) <= '1';
    layer2_outputs(2125) <= (layer1_outputs(3971)) or (layer1_outputs(3777));
    layer2_outputs(2126) <= (layer1_outputs(975)) and (layer1_outputs(1389));
    layer2_outputs(2127) <= '0';
    layer2_outputs(2128) <= (layer1_outputs(5087)) and (layer1_outputs(1151));
    layer2_outputs(2129) <= (layer1_outputs(3896)) xor (layer1_outputs(3312));
    layer2_outputs(2130) <= layer1_outputs(4775);
    layer2_outputs(2131) <= not(layer1_outputs(4146)) or (layer1_outputs(2840));
    layer2_outputs(2132) <= (layer1_outputs(1518)) and (layer1_outputs(2995));
    layer2_outputs(2133) <= not((layer1_outputs(3673)) and (layer1_outputs(638)));
    layer2_outputs(2134) <= not(layer1_outputs(101)) or (layer1_outputs(2400));
    layer2_outputs(2135) <= not((layer1_outputs(4039)) and (layer1_outputs(1864)));
    layer2_outputs(2136) <= not(layer1_outputs(3049)) or (layer1_outputs(3846));
    layer2_outputs(2137) <= not(layer1_outputs(296)) or (layer1_outputs(1686));
    layer2_outputs(2138) <= '1';
    layer2_outputs(2139) <= not(layer1_outputs(1408)) or (layer1_outputs(1287));
    layer2_outputs(2140) <= layer1_outputs(384);
    layer2_outputs(2141) <= not(layer1_outputs(4638));
    layer2_outputs(2142) <= layer1_outputs(4036);
    layer2_outputs(2143) <= '0';
    layer2_outputs(2144) <= (layer1_outputs(1119)) and not (layer1_outputs(3067));
    layer2_outputs(2145) <= layer1_outputs(4117);
    layer2_outputs(2146) <= not(layer1_outputs(2146));
    layer2_outputs(2147) <= '1';
    layer2_outputs(2148) <= (layer1_outputs(1144)) and (layer1_outputs(1572));
    layer2_outputs(2149) <= (layer1_outputs(1847)) or (layer1_outputs(4487));
    layer2_outputs(2150) <= '1';
    layer2_outputs(2151) <= (layer1_outputs(3936)) or (layer1_outputs(3154));
    layer2_outputs(2152) <= not((layer1_outputs(1405)) or (layer1_outputs(2748)));
    layer2_outputs(2153) <= (layer1_outputs(4984)) and not (layer1_outputs(1308));
    layer2_outputs(2154) <= not((layer1_outputs(326)) and (layer1_outputs(300)));
    layer2_outputs(2155) <= (layer1_outputs(206)) and not (layer1_outputs(5048));
    layer2_outputs(2156) <= (layer1_outputs(4310)) and not (layer1_outputs(4587));
    layer2_outputs(2157) <= layer1_outputs(754);
    layer2_outputs(2158) <= '0';
    layer2_outputs(2159) <= (layer1_outputs(418)) and (layer1_outputs(3106));
    layer2_outputs(2160) <= (layer1_outputs(538)) xor (layer1_outputs(4839));
    layer2_outputs(2161) <= not((layer1_outputs(4136)) xor (layer1_outputs(2812)));
    layer2_outputs(2162) <= '1';
    layer2_outputs(2163) <= not(layer1_outputs(1016));
    layer2_outputs(2164) <= layer1_outputs(3395);
    layer2_outputs(2165) <= not(layer1_outputs(2182)) or (layer1_outputs(4772));
    layer2_outputs(2166) <= not(layer1_outputs(4344));
    layer2_outputs(2167) <= (layer1_outputs(3458)) or (layer1_outputs(4501));
    layer2_outputs(2168) <= not(layer1_outputs(4225));
    layer2_outputs(2169) <= (layer1_outputs(3690)) and (layer1_outputs(712));
    layer2_outputs(2170) <= '1';
    layer2_outputs(2171) <= (layer1_outputs(3014)) xor (layer1_outputs(108));
    layer2_outputs(2172) <= (layer1_outputs(4094)) or (layer1_outputs(330));
    layer2_outputs(2173) <= layer1_outputs(3917);
    layer2_outputs(2174) <= (layer1_outputs(3863)) and not (layer1_outputs(4208));
    layer2_outputs(2175) <= not((layer1_outputs(4668)) or (layer1_outputs(1971)));
    layer2_outputs(2176) <= not((layer1_outputs(4947)) or (layer1_outputs(4406)));
    layer2_outputs(2177) <= not(layer1_outputs(5047));
    layer2_outputs(2178) <= not((layer1_outputs(2049)) xor (layer1_outputs(2045)));
    layer2_outputs(2179) <= '1';
    layer2_outputs(2180) <= '0';
    layer2_outputs(2181) <= '0';
    layer2_outputs(2182) <= not(layer1_outputs(514));
    layer2_outputs(2183) <= not((layer1_outputs(1424)) or (layer1_outputs(1401)));
    layer2_outputs(2184) <= (layer1_outputs(1651)) and not (layer1_outputs(4143));
    layer2_outputs(2185) <= '1';
    layer2_outputs(2186) <= '1';
    layer2_outputs(2187) <= not(layer1_outputs(3074)) or (layer1_outputs(4877));
    layer2_outputs(2188) <= (layer1_outputs(1276)) and not (layer1_outputs(4928));
    layer2_outputs(2189) <= '1';
    layer2_outputs(2190) <= (layer1_outputs(3230)) and (layer1_outputs(1570));
    layer2_outputs(2191) <= not((layer1_outputs(2232)) or (layer1_outputs(88)));
    layer2_outputs(2192) <= (layer1_outputs(2977)) and (layer1_outputs(4363));
    layer2_outputs(2193) <= (layer1_outputs(4933)) or (layer1_outputs(1564));
    layer2_outputs(2194) <= (layer1_outputs(2904)) and (layer1_outputs(5106));
    layer2_outputs(2195) <= (layer1_outputs(2329)) or (layer1_outputs(1217));
    layer2_outputs(2196) <= (layer1_outputs(2142)) and not (layer1_outputs(2160));
    layer2_outputs(2197) <= not((layer1_outputs(3722)) and (layer1_outputs(958)));
    layer2_outputs(2198) <= '1';
    layer2_outputs(2199) <= '1';
    layer2_outputs(2200) <= layer1_outputs(2666);
    layer2_outputs(2201) <= not(layer1_outputs(4790)) or (layer1_outputs(1429));
    layer2_outputs(2202) <= layer1_outputs(4915);
    layer2_outputs(2203) <= layer1_outputs(594);
    layer2_outputs(2204) <= not(layer1_outputs(3715)) or (layer1_outputs(2287));
    layer2_outputs(2205) <= '1';
    layer2_outputs(2206) <= not(layer1_outputs(1841)) or (layer1_outputs(4345));
    layer2_outputs(2207) <= layer1_outputs(2573);
    layer2_outputs(2208) <= not(layer1_outputs(4099)) or (layer1_outputs(3614));
    layer2_outputs(2209) <= not(layer1_outputs(4767));
    layer2_outputs(2210) <= (layer1_outputs(5010)) and (layer1_outputs(806));
    layer2_outputs(2211) <= not((layer1_outputs(3381)) or (layer1_outputs(1200)));
    layer2_outputs(2212) <= '0';
    layer2_outputs(2213) <= (layer1_outputs(1775)) and (layer1_outputs(3214));
    layer2_outputs(2214) <= (layer1_outputs(2834)) and not (layer1_outputs(1098));
    layer2_outputs(2215) <= '1';
    layer2_outputs(2216) <= not(layer1_outputs(1475)) or (layer1_outputs(506));
    layer2_outputs(2217) <= (layer1_outputs(2936)) and not (layer1_outputs(3736));
    layer2_outputs(2218) <= '0';
    layer2_outputs(2219) <= not(layer1_outputs(129));
    layer2_outputs(2220) <= (layer1_outputs(3388)) and (layer1_outputs(4800));
    layer2_outputs(2221) <= (layer1_outputs(4474)) and (layer1_outputs(2021));
    layer2_outputs(2222) <= not(layer1_outputs(2886));
    layer2_outputs(2223) <= '1';
    layer2_outputs(2224) <= not(layer1_outputs(3609)) or (layer1_outputs(2040));
    layer2_outputs(2225) <= (layer1_outputs(4076)) or (layer1_outputs(3111));
    layer2_outputs(2226) <= not((layer1_outputs(4390)) or (layer1_outputs(344)));
    layer2_outputs(2227) <= '0';
    layer2_outputs(2228) <= (layer1_outputs(1744)) and not (layer1_outputs(3067));
    layer2_outputs(2229) <= (layer1_outputs(1223)) and not (layer1_outputs(2508));
    layer2_outputs(2230) <= '0';
    layer2_outputs(2231) <= '0';
    layer2_outputs(2232) <= (layer1_outputs(2698)) and (layer1_outputs(4103));
    layer2_outputs(2233) <= (layer1_outputs(1112)) and not (layer1_outputs(1022));
    layer2_outputs(2234) <= '0';
    layer2_outputs(2235) <= not(layer1_outputs(2159));
    layer2_outputs(2236) <= (layer1_outputs(4401)) and not (layer1_outputs(324));
    layer2_outputs(2237) <= layer1_outputs(4629);
    layer2_outputs(2238) <= not(layer1_outputs(3377));
    layer2_outputs(2239) <= layer1_outputs(2717);
    layer2_outputs(2240) <= not((layer1_outputs(2476)) and (layer1_outputs(922)));
    layer2_outputs(2241) <= (layer1_outputs(4960)) and not (layer1_outputs(364));
    layer2_outputs(2242) <= (layer1_outputs(2089)) or (layer1_outputs(5117));
    layer2_outputs(2243) <= (layer1_outputs(3073)) and not (layer1_outputs(1488));
    layer2_outputs(2244) <= not(layer1_outputs(4121)) or (layer1_outputs(395));
    layer2_outputs(2245) <= (layer1_outputs(3015)) and not (layer1_outputs(2642));
    layer2_outputs(2246) <= '0';
    layer2_outputs(2247) <= (layer1_outputs(4847)) and (layer1_outputs(199));
    layer2_outputs(2248) <= layer1_outputs(672);
    layer2_outputs(2249) <= not((layer1_outputs(4511)) or (layer1_outputs(1606)));
    layer2_outputs(2250) <= '1';
    layer2_outputs(2251) <= '1';
    layer2_outputs(2252) <= (layer1_outputs(2848)) and not (layer1_outputs(3945));
    layer2_outputs(2253) <= (layer1_outputs(629)) xor (layer1_outputs(419));
    layer2_outputs(2254) <= not((layer1_outputs(248)) and (layer1_outputs(1034)));
    layer2_outputs(2255) <= '0';
    layer2_outputs(2256) <= layer1_outputs(820);
    layer2_outputs(2257) <= (layer1_outputs(2237)) and (layer1_outputs(968));
    layer2_outputs(2258) <= not((layer1_outputs(4733)) and (layer1_outputs(3047)));
    layer2_outputs(2259) <= not((layer1_outputs(4664)) or (layer1_outputs(3062)));
    layer2_outputs(2260) <= '0';
    layer2_outputs(2261) <= '1';
    layer2_outputs(2262) <= '1';
    layer2_outputs(2263) <= (layer1_outputs(3540)) and not (layer1_outputs(4580));
    layer2_outputs(2264) <= not(layer1_outputs(1158));
    layer2_outputs(2265) <= not(layer1_outputs(1708)) or (layer1_outputs(274));
    layer2_outputs(2266) <= (layer1_outputs(3730)) and not (layer1_outputs(441));
    layer2_outputs(2267) <= layer1_outputs(2160);
    layer2_outputs(2268) <= not(layer1_outputs(3948)) or (layer1_outputs(930));
    layer2_outputs(2269) <= layer1_outputs(5072);
    layer2_outputs(2270) <= (layer1_outputs(1613)) and not (layer1_outputs(3475));
    layer2_outputs(2271) <= (layer1_outputs(1092)) or (layer1_outputs(1273));
    layer2_outputs(2272) <= (layer1_outputs(1821)) or (layer1_outputs(4456));
    layer2_outputs(2273) <= layer1_outputs(152);
    layer2_outputs(2274) <= (layer1_outputs(2055)) and (layer1_outputs(1770));
    layer2_outputs(2275) <= (layer1_outputs(2116)) and not (layer1_outputs(2530));
    layer2_outputs(2276) <= not(layer1_outputs(377)) or (layer1_outputs(4936));
    layer2_outputs(2277) <= not(layer1_outputs(964)) or (layer1_outputs(1956));
    layer2_outputs(2278) <= '0';
    layer2_outputs(2279) <= not(layer1_outputs(2262));
    layer2_outputs(2280) <= not(layer1_outputs(2471));
    layer2_outputs(2281) <= '0';
    layer2_outputs(2282) <= '1';
    layer2_outputs(2283) <= not((layer1_outputs(767)) and (layer1_outputs(1442)));
    layer2_outputs(2284) <= '1';
    layer2_outputs(2285) <= not((layer1_outputs(2082)) or (layer1_outputs(1701)));
    layer2_outputs(2286) <= (layer1_outputs(3598)) and (layer1_outputs(4820));
    layer2_outputs(2287) <= not(layer1_outputs(2701));
    layer2_outputs(2288) <= '0';
    layer2_outputs(2289) <= not((layer1_outputs(4280)) or (layer1_outputs(4853)));
    layer2_outputs(2290) <= '1';
    layer2_outputs(2291) <= '0';
    layer2_outputs(2292) <= (layer1_outputs(2476)) or (layer1_outputs(4013));
    layer2_outputs(2293) <= layer1_outputs(4046);
    layer2_outputs(2294) <= not(layer1_outputs(2268)) or (layer1_outputs(4469));
    layer2_outputs(2295) <= layer1_outputs(1464);
    layer2_outputs(2296) <= (layer1_outputs(16)) and not (layer1_outputs(3592));
    layer2_outputs(2297) <= (layer1_outputs(1482)) and (layer1_outputs(3107));
    layer2_outputs(2298) <= (layer1_outputs(19)) and (layer1_outputs(2446));
    layer2_outputs(2299) <= not(layer1_outputs(3176));
    layer2_outputs(2300) <= (layer1_outputs(4527)) and (layer1_outputs(1561));
    layer2_outputs(2301) <= not(layer1_outputs(4914)) or (layer1_outputs(3531));
    layer2_outputs(2302) <= not(layer1_outputs(3712));
    layer2_outputs(2303) <= (layer1_outputs(762)) and not (layer1_outputs(3112));
    layer2_outputs(2304) <= '1';
    layer2_outputs(2305) <= not((layer1_outputs(1079)) xor (layer1_outputs(157)));
    layer2_outputs(2306) <= (layer1_outputs(1815)) and (layer1_outputs(3805));
    layer2_outputs(2307) <= not((layer1_outputs(2393)) or (layer1_outputs(3723)));
    layer2_outputs(2308) <= layer1_outputs(175);
    layer2_outputs(2309) <= not(layer1_outputs(1115));
    layer2_outputs(2310) <= '0';
    layer2_outputs(2311) <= (layer1_outputs(1504)) or (layer1_outputs(1665));
    layer2_outputs(2312) <= layer1_outputs(435);
    layer2_outputs(2313) <= not((layer1_outputs(3418)) or (layer1_outputs(2553)));
    layer2_outputs(2314) <= not((layer1_outputs(1683)) or (layer1_outputs(1200)));
    layer2_outputs(2315) <= '1';
    layer2_outputs(2316) <= layer1_outputs(4471);
    layer2_outputs(2317) <= not((layer1_outputs(2364)) and (layer1_outputs(4365)));
    layer2_outputs(2318) <= not((layer1_outputs(342)) or (layer1_outputs(551)));
    layer2_outputs(2319) <= (layer1_outputs(434)) and (layer1_outputs(3658));
    layer2_outputs(2320) <= '0';
    layer2_outputs(2321) <= not((layer1_outputs(2989)) and (layer1_outputs(1800)));
    layer2_outputs(2322) <= (layer1_outputs(3831)) and not (layer1_outputs(315));
    layer2_outputs(2323) <= (layer1_outputs(869)) or (layer1_outputs(2539));
    layer2_outputs(2324) <= '1';
    layer2_outputs(2325) <= (layer1_outputs(2258)) and not (layer1_outputs(2288));
    layer2_outputs(2326) <= (layer1_outputs(5038)) or (layer1_outputs(1519));
    layer2_outputs(2327) <= not((layer1_outputs(2963)) or (layer1_outputs(1912)));
    layer2_outputs(2328) <= not(layer1_outputs(3180)) or (layer1_outputs(884));
    layer2_outputs(2329) <= not(layer1_outputs(4810));
    layer2_outputs(2330) <= not((layer1_outputs(1354)) or (layer1_outputs(1438)));
    layer2_outputs(2331) <= not(layer1_outputs(3985)) or (layer1_outputs(3048));
    layer2_outputs(2332) <= layer1_outputs(4475);
    layer2_outputs(2333) <= layer1_outputs(4466);
    layer2_outputs(2334) <= (layer1_outputs(1398)) and not (layer1_outputs(5002));
    layer2_outputs(2335) <= '1';
    layer2_outputs(2336) <= not(layer1_outputs(1362)) or (layer1_outputs(550));
    layer2_outputs(2337) <= not((layer1_outputs(2150)) and (layer1_outputs(4198)));
    layer2_outputs(2338) <= '1';
    layer2_outputs(2339) <= not(layer1_outputs(1502)) or (layer1_outputs(4438));
    layer2_outputs(2340) <= '0';
    layer2_outputs(2341) <= '0';
    layer2_outputs(2342) <= '0';
    layer2_outputs(2343) <= not(layer1_outputs(3305)) or (layer1_outputs(3769));
    layer2_outputs(2344) <= not(layer1_outputs(2567));
    layer2_outputs(2345) <= layer1_outputs(1998);
    layer2_outputs(2346) <= not(layer1_outputs(1041)) or (layer1_outputs(1636));
    layer2_outputs(2347) <= '0';
    layer2_outputs(2348) <= (layer1_outputs(3691)) or (layer1_outputs(3271));
    layer2_outputs(2349) <= (layer1_outputs(3240)) and (layer1_outputs(1106));
    layer2_outputs(2350) <= not(layer1_outputs(4617));
    layer2_outputs(2351) <= (layer1_outputs(1412)) and not (layer1_outputs(4911));
    layer2_outputs(2352) <= (layer1_outputs(4611)) and (layer1_outputs(4158));
    layer2_outputs(2353) <= '0';
    layer2_outputs(2354) <= '1';
    layer2_outputs(2355) <= (layer1_outputs(173)) and (layer1_outputs(3695));
    layer2_outputs(2356) <= not((layer1_outputs(4202)) and (layer1_outputs(2687)));
    layer2_outputs(2357) <= not(layer1_outputs(1332));
    layer2_outputs(2358) <= not(layer1_outputs(1625)) or (layer1_outputs(4333));
    layer2_outputs(2359) <= layer1_outputs(4476);
    layer2_outputs(2360) <= not(layer1_outputs(4446)) or (layer1_outputs(3869));
    layer2_outputs(2361) <= (layer1_outputs(2468)) and not (layer1_outputs(3584));
    layer2_outputs(2362) <= (layer1_outputs(879)) and (layer1_outputs(1166));
    layer2_outputs(2363) <= (layer1_outputs(3735)) and (layer1_outputs(192));
    layer2_outputs(2364) <= '0';
    layer2_outputs(2365) <= not(layer1_outputs(1679)) or (layer1_outputs(102));
    layer2_outputs(2366) <= layer1_outputs(3676);
    layer2_outputs(2367) <= (layer1_outputs(128)) and not (layer1_outputs(2100));
    layer2_outputs(2368) <= (layer1_outputs(3168)) and not (layer1_outputs(1668));
    layer2_outputs(2369) <= (layer1_outputs(2059)) and not (layer1_outputs(4002));
    layer2_outputs(2370) <= '1';
    layer2_outputs(2371) <= (layer1_outputs(1006)) and not (layer1_outputs(1914));
    layer2_outputs(2372) <= (layer1_outputs(2740)) and (layer1_outputs(1010));
    layer2_outputs(2373) <= not(layer1_outputs(109)) or (layer1_outputs(528));
    layer2_outputs(2374) <= (layer1_outputs(1778)) and not (layer1_outputs(1210));
    layer2_outputs(2375) <= not(layer1_outputs(4940));
    layer2_outputs(2376) <= layer1_outputs(4144);
    layer2_outputs(2377) <= layer1_outputs(3367);
    layer2_outputs(2378) <= layer1_outputs(360);
    layer2_outputs(2379) <= not((layer1_outputs(2564)) or (layer1_outputs(2677)));
    layer2_outputs(2380) <= '1';
    layer2_outputs(2381) <= '1';
    layer2_outputs(2382) <= not((layer1_outputs(2251)) and (layer1_outputs(2312)));
    layer2_outputs(2383) <= '0';
    layer2_outputs(2384) <= (layer1_outputs(3805)) and not (layer1_outputs(2388));
    layer2_outputs(2385) <= not((layer1_outputs(4302)) and (layer1_outputs(4426)));
    layer2_outputs(2386) <= (layer1_outputs(4172)) and not (layer1_outputs(1777));
    layer2_outputs(2387) <= (layer1_outputs(3696)) and not (layer1_outputs(821));
    layer2_outputs(2388) <= not(layer1_outputs(493)) or (layer1_outputs(2813));
    layer2_outputs(2389) <= not((layer1_outputs(4397)) or (layer1_outputs(1471)));
    layer2_outputs(2390) <= not(layer1_outputs(683)) or (layer1_outputs(1128));
    layer2_outputs(2391) <= (layer1_outputs(4262)) and not (layer1_outputs(868));
    layer2_outputs(2392) <= '0';
    layer2_outputs(2393) <= not(layer1_outputs(4993));
    layer2_outputs(2394) <= (layer1_outputs(1023)) and (layer1_outputs(22));
    layer2_outputs(2395) <= not(layer1_outputs(2307)) or (layer1_outputs(2489));
    layer2_outputs(2396) <= not((layer1_outputs(521)) and (layer1_outputs(3774)));
    layer2_outputs(2397) <= '1';
    layer2_outputs(2398) <= '0';
    layer2_outputs(2399) <= layer1_outputs(3921);
    layer2_outputs(2400) <= not((layer1_outputs(4693)) or (layer1_outputs(4472)));
    layer2_outputs(2401) <= (layer1_outputs(3956)) and (layer1_outputs(1674));
    layer2_outputs(2402) <= '1';
    layer2_outputs(2403) <= (layer1_outputs(163)) and not (layer1_outputs(4925));
    layer2_outputs(2404) <= layer1_outputs(4498);
    layer2_outputs(2405) <= not(layer1_outputs(319)) or (layer1_outputs(1948));
    layer2_outputs(2406) <= layer1_outputs(2711);
    layer2_outputs(2407) <= (layer1_outputs(4805)) or (layer1_outputs(5059));
    layer2_outputs(2408) <= (layer1_outputs(1630)) and (layer1_outputs(4078));
    layer2_outputs(2409) <= layer1_outputs(4952);
    layer2_outputs(2410) <= layer1_outputs(276);
    layer2_outputs(2411) <= (layer1_outputs(1782)) and (layer1_outputs(1803));
    layer2_outputs(2412) <= (layer1_outputs(1271)) and (layer1_outputs(4821));
    layer2_outputs(2413) <= (layer1_outputs(2208)) and (layer1_outputs(4067));
    layer2_outputs(2414) <= not((layer1_outputs(3813)) or (layer1_outputs(842)));
    layer2_outputs(2415) <= layer1_outputs(4037);
    layer2_outputs(2416) <= (layer1_outputs(4587)) and (layer1_outputs(1372));
    layer2_outputs(2417) <= not(layer1_outputs(351));
    layer2_outputs(2418) <= not((layer1_outputs(1258)) and (layer1_outputs(4271)));
    layer2_outputs(2419) <= not(layer1_outputs(3005)) or (layer1_outputs(610));
    layer2_outputs(2420) <= '0';
    layer2_outputs(2421) <= (layer1_outputs(899)) or (layer1_outputs(1725));
    layer2_outputs(2422) <= not(layer1_outputs(1376));
    layer2_outputs(2423) <= not(layer1_outputs(3187));
    layer2_outputs(2424) <= not(layer1_outputs(4017));
    layer2_outputs(2425) <= (layer1_outputs(4814)) and not (layer1_outputs(436));
    layer2_outputs(2426) <= layer1_outputs(1600);
    layer2_outputs(2427) <= (layer1_outputs(3921)) or (layer1_outputs(299));
    layer2_outputs(2428) <= (layer1_outputs(2121)) and not (layer1_outputs(2583));
    layer2_outputs(2429) <= not((layer1_outputs(3087)) and (layer1_outputs(1604)));
    layer2_outputs(2430) <= not((layer1_outputs(3046)) and (layer1_outputs(730)));
    layer2_outputs(2431) <= '0';
    layer2_outputs(2432) <= (layer1_outputs(5066)) and not (layer1_outputs(2735));
    layer2_outputs(2433) <= not((layer1_outputs(225)) or (layer1_outputs(664)));
    layer2_outputs(2434) <= '1';
    layer2_outputs(2435) <= not((layer1_outputs(3487)) or (layer1_outputs(1842)));
    layer2_outputs(2436) <= (layer1_outputs(96)) and not (layer1_outputs(2690));
    layer2_outputs(2437) <= (layer1_outputs(614)) and not (layer1_outputs(4995));
    layer2_outputs(2438) <= '0';
    layer2_outputs(2439) <= (layer1_outputs(4657)) and (layer1_outputs(4195));
    layer2_outputs(2440) <= not(layer1_outputs(3156)) or (layer1_outputs(2898));
    layer2_outputs(2441) <= (layer1_outputs(2738)) or (layer1_outputs(1497));
    layer2_outputs(2442) <= (layer1_outputs(4819)) and not (layer1_outputs(3514));
    layer2_outputs(2443) <= not(layer1_outputs(937));
    layer2_outputs(2444) <= '0';
    layer2_outputs(2445) <= not(layer1_outputs(52)) or (layer1_outputs(4065));
    layer2_outputs(2446) <= not(layer1_outputs(1194)) or (layer1_outputs(4429));
    layer2_outputs(2447) <= not((layer1_outputs(571)) and (layer1_outputs(2901)));
    layer2_outputs(2448) <= '1';
    layer2_outputs(2449) <= '1';
    layer2_outputs(2450) <= not((layer1_outputs(1779)) and (layer1_outputs(1551)));
    layer2_outputs(2451) <= (layer1_outputs(188)) or (layer1_outputs(4670));
    layer2_outputs(2452) <= not((layer1_outputs(1559)) and (layer1_outputs(3478)));
    layer2_outputs(2453) <= '0';
    layer2_outputs(2454) <= not((layer1_outputs(4701)) and (layer1_outputs(2845)));
    layer2_outputs(2455) <= not(layer1_outputs(3605));
    layer2_outputs(2456) <= not((layer1_outputs(1307)) or (layer1_outputs(85)));
    layer2_outputs(2457) <= layer1_outputs(3926);
    layer2_outputs(2458) <= not(layer1_outputs(3953)) or (layer1_outputs(2612));
    layer2_outputs(2459) <= not((layer1_outputs(2558)) and (layer1_outputs(4186)));
    layer2_outputs(2460) <= not(layer1_outputs(4860));
    layer2_outputs(2461) <= (layer1_outputs(3894)) and (layer1_outputs(3189));
    layer2_outputs(2462) <= '0';
    layer2_outputs(2463) <= layer1_outputs(4177);
    layer2_outputs(2464) <= not((layer1_outputs(1378)) or (layer1_outputs(2931)));
    layer2_outputs(2465) <= not((layer1_outputs(1359)) xor (layer1_outputs(3315)));
    layer2_outputs(2466) <= '1';
    layer2_outputs(2467) <= not((layer1_outputs(4231)) and (layer1_outputs(803)));
    layer2_outputs(2468) <= not(layer1_outputs(4192)) or (layer1_outputs(3361));
    layer2_outputs(2469) <= not(layer1_outputs(2133));
    layer2_outputs(2470) <= '1';
    layer2_outputs(2471) <= not((layer1_outputs(4994)) and (layer1_outputs(1514)));
    layer2_outputs(2472) <= '1';
    layer2_outputs(2473) <= '0';
    layer2_outputs(2474) <= not((layer1_outputs(4833)) or (layer1_outputs(4857)));
    layer2_outputs(2475) <= not((layer1_outputs(1241)) or (layer1_outputs(3994)));
    layer2_outputs(2476) <= '0';
    layer2_outputs(2477) <= (layer1_outputs(1780)) and (layer1_outputs(3192));
    layer2_outputs(2478) <= not(layer1_outputs(4803));
    layer2_outputs(2479) <= '0';
    layer2_outputs(2480) <= not(layer1_outputs(284)) or (layer1_outputs(4971));
    layer2_outputs(2481) <= not(layer1_outputs(1051)) or (layer1_outputs(1052));
    layer2_outputs(2482) <= layer1_outputs(2461);
    layer2_outputs(2483) <= not((layer1_outputs(3966)) and (layer1_outputs(3483)));
    layer2_outputs(2484) <= (layer1_outputs(1035)) and not (layer1_outputs(323));
    layer2_outputs(2485) <= not(layer1_outputs(1268));
    layer2_outputs(2486) <= not(layer1_outputs(4927)) or (layer1_outputs(2739));
    layer2_outputs(2487) <= '0';
    layer2_outputs(2488) <= not(layer1_outputs(474)) or (layer1_outputs(2231));
    layer2_outputs(2489) <= (layer1_outputs(63)) and not (layer1_outputs(1380));
    layer2_outputs(2490) <= (layer1_outputs(3670)) and not (layer1_outputs(2625));
    layer2_outputs(2491) <= not(layer1_outputs(2511));
    layer2_outputs(2492) <= not((layer1_outputs(4995)) or (layer1_outputs(1868)));
    layer2_outputs(2493) <= not((layer1_outputs(485)) or (layer1_outputs(4683)));
    layer2_outputs(2494) <= not(layer1_outputs(2287)) or (layer1_outputs(2310));
    layer2_outputs(2495) <= '0';
    layer2_outputs(2496) <= not(layer1_outputs(1088)) or (layer1_outputs(5091));
    layer2_outputs(2497) <= not((layer1_outputs(5054)) and (layer1_outputs(4035)));
    layer2_outputs(2498) <= not((layer1_outputs(775)) and (layer1_outputs(2372)));
    layer2_outputs(2499) <= not(layer1_outputs(4494)) or (layer1_outputs(3501));
    layer2_outputs(2500) <= (layer1_outputs(739)) and (layer1_outputs(2342));
    layer2_outputs(2501) <= (layer1_outputs(2958)) and not (layer1_outputs(1669));
    layer2_outputs(2502) <= (layer1_outputs(682)) and (layer1_outputs(221));
    layer2_outputs(2503) <= '0';
    layer2_outputs(2504) <= (layer1_outputs(358)) xor (layer1_outputs(2691));
    layer2_outputs(2505) <= not((layer1_outputs(3184)) and (layer1_outputs(1311)));
    layer2_outputs(2506) <= '1';
    layer2_outputs(2507) <= not(layer1_outputs(408)) or (layer1_outputs(3432));
    layer2_outputs(2508) <= (layer1_outputs(1257)) and not (layer1_outputs(4016));
    layer2_outputs(2509) <= not(layer1_outputs(2648)) or (layer1_outputs(4278));
    layer2_outputs(2510) <= '1';
    layer2_outputs(2511) <= not((layer1_outputs(2253)) and (layer1_outputs(2387)));
    layer2_outputs(2512) <= not((layer1_outputs(1073)) and (layer1_outputs(744)));
    layer2_outputs(2513) <= '0';
    layer2_outputs(2514) <= layer1_outputs(3597);
    layer2_outputs(2515) <= (layer1_outputs(3457)) and (layer1_outputs(1937));
    layer2_outputs(2516) <= layer1_outputs(568);
    layer2_outputs(2517) <= not(layer1_outputs(1502));
    layer2_outputs(2518) <= not(layer1_outputs(1112)) or (layer1_outputs(189));
    layer2_outputs(2519) <= '1';
    layer2_outputs(2520) <= '0';
    layer2_outputs(2521) <= layer1_outputs(1571);
    layer2_outputs(2522) <= (layer1_outputs(2154)) and (layer1_outputs(3368));
    layer2_outputs(2523) <= not((layer1_outputs(4897)) or (layer1_outputs(4419)));
    layer2_outputs(2524) <= (layer1_outputs(2588)) and not (layer1_outputs(4906));
    layer2_outputs(2525) <= not(layer1_outputs(3099));
    layer2_outputs(2526) <= not((layer1_outputs(2196)) or (layer1_outputs(4568)));
    layer2_outputs(2527) <= not((layer1_outputs(3077)) or (layer1_outputs(4502)));
    layer2_outputs(2528) <= (layer1_outputs(1777)) or (layer1_outputs(1514));
    layer2_outputs(2529) <= not(layer1_outputs(4635)) or (layer1_outputs(4934));
    layer2_outputs(2530) <= not((layer1_outputs(2048)) or (layer1_outputs(2858)));
    layer2_outputs(2531) <= (layer1_outputs(1040)) or (layer1_outputs(4596));
    layer2_outputs(2532) <= (layer1_outputs(2188)) and not (layer1_outputs(3011));
    layer2_outputs(2533) <= (layer1_outputs(2768)) and (layer1_outputs(4413));
    layer2_outputs(2534) <= (layer1_outputs(1814)) and not (layer1_outputs(3012));
    layer2_outputs(2535) <= '0';
    layer2_outputs(2536) <= (layer1_outputs(1841)) and not (layer1_outputs(2467));
    layer2_outputs(2537) <= '0';
    layer2_outputs(2538) <= not((layer1_outputs(1352)) and (layer1_outputs(4709)));
    layer2_outputs(2539) <= (layer1_outputs(2517)) and not (layer1_outputs(1846));
    layer2_outputs(2540) <= not((layer1_outputs(4445)) or (layer1_outputs(3056)));
    layer2_outputs(2541) <= not(layer1_outputs(1261));
    layer2_outputs(2542) <= layer1_outputs(1381);
    layer2_outputs(2543) <= not((layer1_outputs(898)) and (layer1_outputs(2291)));
    layer2_outputs(2544) <= layer1_outputs(4496);
    layer2_outputs(2545) <= layer1_outputs(97);
    layer2_outputs(2546) <= not(layer1_outputs(4473));
    layer2_outputs(2547) <= (layer1_outputs(200)) and not (layer1_outputs(2230));
    layer2_outputs(2548) <= not((layer1_outputs(3023)) and (layer1_outputs(5007)));
    layer2_outputs(2549) <= layer1_outputs(4151);
    layer2_outputs(2550) <= layer1_outputs(4827);
    layer2_outputs(2551) <= '1';
    layer2_outputs(2552) <= not(layer1_outputs(2503)) or (layer1_outputs(18));
    layer2_outputs(2553) <= not(layer1_outputs(284)) or (layer1_outputs(4979));
    layer2_outputs(2554) <= '1';
    layer2_outputs(2555) <= (layer1_outputs(5078)) and (layer1_outputs(982));
    layer2_outputs(2556) <= '0';
    layer2_outputs(2557) <= not((layer1_outputs(856)) or (layer1_outputs(1149)));
    layer2_outputs(2558) <= (layer1_outputs(1254)) and not (layer1_outputs(4359));
    layer2_outputs(2559) <= (layer1_outputs(2651)) and not (layer1_outputs(2642));
    layer2_outputs(2560) <= layer1_outputs(5022);
    layer2_outputs(2561) <= (layer1_outputs(1432)) or (layer1_outputs(2407));
    layer2_outputs(2562) <= not(layer1_outputs(1392)) or (layer1_outputs(5067));
    layer2_outputs(2563) <= not(layer1_outputs(164));
    layer2_outputs(2564) <= layer1_outputs(1355);
    layer2_outputs(2565) <= not(layer1_outputs(4983));
    layer2_outputs(2566) <= (layer1_outputs(3394)) and not (layer1_outputs(4369));
    layer2_outputs(2567) <= '1';
    layer2_outputs(2568) <= '1';
    layer2_outputs(2569) <= (layer1_outputs(1967)) and (layer1_outputs(4206));
    layer2_outputs(2570) <= (layer1_outputs(2425)) or (layer1_outputs(1500));
    layer2_outputs(2571) <= not((layer1_outputs(740)) or (layer1_outputs(1289)));
    layer2_outputs(2572) <= not((layer1_outputs(3803)) and (layer1_outputs(3692)));
    layer2_outputs(2573) <= layer1_outputs(230);
    layer2_outputs(2574) <= '1';
    layer2_outputs(2575) <= (layer1_outputs(4637)) and (layer1_outputs(4717));
    layer2_outputs(2576) <= (layer1_outputs(3814)) and not (layer1_outputs(1062));
    layer2_outputs(2577) <= '0';
    layer2_outputs(2578) <= (layer1_outputs(4797)) and not (layer1_outputs(2705));
    layer2_outputs(2579) <= not((layer1_outputs(742)) and (layer1_outputs(3205)));
    layer2_outputs(2580) <= not(layer1_outputs(3131));
    layer2_outputs(2581) <= not(layer1_outputs(1284)) or (layer1_outputs(1175));
    layer2_outputs(2582) <= '0';
    layer2_outputs(2583) <= (layer1_outputs(4388)) and (layer1_outputs(2868));
    layer2_outputs(2584) <= (layer1_outputs(5083)) or (layer1_outputs(121));
    layer2_outputs(2585) <= not(layer1_outputs(4747)) or (layer1_outputs(2940));
    layer2_outputs(2586) <= '1';
    layer2_outputs(2587) <= '0';
    layer2_outputs(2588) <= '0';
    layer2_outputs(2589) <= not((layer1_outputs(2753)) or (layer1_outputs(223)));
    layer2_outputs(2590) <= (layer1_outputs(3880)) xor (layer1_outputs(634));
    layer2_outputs(2591) <= layer1_outputs(3580);
    layer2_outputs(2592) <= '1';
    layer2_outputs(2593) <= '0';
    layer2_outputs(2594) <= not((layer1_outputs(3346)) xor (layer1_outputs(4732)));
    layer2_outputs(2595) <= (layer1_outputs(1253)) and not (layer1_outputs(3227));
    layer2_outputs(2596) <= '1';
    layer2_outputs(2597) <= not(layer1_outputs(1377)) or (layer1_outputs(4282));
    layer2_outputs(2598) <= '1';
    layer2_outputs(2599) <= (layer1_outputs(3069)) xor (layer1_outputs(1470));
    layer2_outputs(2600) <= layer1_outputs(4669);
    layer2_outputs(2601) <= (layer1_outputs(5089)) and (layer1_outputs(1213));
    layer2_outputs(2602) <= layer1_outputs(1507);
    layer2_outputs(2603) <= '0';
    layer2_outputs(2604) <= not((layer1_outputs(477)) or (layer1_outputs(468)));
    layer2_outputs(2605) <= not(layer1_outputs(2980));
    layer2_outputs(2606) <= (layer1_outputs(4137)) xor (layer1_outputs(3914));
    layer2_outputs(2607) <= not(layer1_outputs(4946)) or (layer1_outputs(4554));
    layer2_outputs(2608) <= not(layer1_outputs(1499)) or (layer1_outputs(566));
    layer2_outputs(2609) <= layer1_outputs(1402);
    layer2_outputs(2610) <= '1';
    layer2_outputs(2611) <= not(layer1_outputs(3306)) or (layer1_outputs(5081));
    layer2_outputs(2612) <= not((layer1_outputs(2028)) or (layer1_outputs(579)));
    layer2_outputs(2613) <= not((layer1_outputs(3787)) xor (layer1_outputs(2643)));
    layer2_outputs(2614) <= not(layer1_outputs(5009));
    layer2_outputs(2615) <= '1';
    layer2_outputs(2616) <= '1';
    layer2_outputs(2617) <= not(layer1_outputs(1840)) or (layer1_outputs(1646));
    layer2_outputs(2618) <= '0';
    layer2_outputs(2619) <= not(layer1_outputs(439));
    layer2_outputs(2620) <= not(layer1_outputs(3693));
    layer2_outputs(2621) <= layer1_outputs(3960);
    layer2_outputs(2622) <= (layer1_outputs(2187)) and not (layer1_outputs(3906));
    layer2_outputs(2623) <= not(layer1_outputs(847)) or (layer1_outputs(3571));
    layer2_outputs(2624) <= '1';
    layer2_outputs(2625) <= (layer1_outputs(2543)) and not (layer1_outputs(4153));
    layer2_outputs(2626) <= '0';
    layer2_outputs(2627) <= '1';
    layer2_outputs(2628) <= not((layer1_outputs(1304)) or (layer1_outputs(3293)));
    layer2_outputs(2629) <= '1';
    layer2_outputs(2630) <= (layer1_outputs(1163)) and not (layer1_outputs(1921));
    layer2_outputs(2631) <= not(layer1_outputs(2967)) or (layer1_outputs(1812));
    layer2_outputs(2632) <= (layer1_outputs(1889)) and not (layer1_outputs(1259));
    layer2_outputs(2633) <= not(layer1_outputs(4143));
    layer2_outputs(2634) <= layer1_outputs(2390);
    layer2_outputs(2635) <= not((layer1_outputs(610)) xor (layer1_outputs(1044)));
    layer2_outputs(2636) <= (layer1_outputs(1064)) and (layer1_outputs(3958));
    layer2_outputs(2637) <= layer1_outputs(3969);
    layer2_outputs(2638) <= '1';
    layer2_outputs(2639) <= not(layer1_outputs(4757));
    layer2_outputs(2640) <= not(layer1_outputs(1098)) or (layer1_outputs(1117));
    layer2_outputs(2641) <= not(layer1_outputs(3811));
    layer2_outputs(2642) <= (layer1_outputs(459)) or (layer1_outputs(2689));
    layer2_outputs(2643) <= not(layer1_outputs(3720)) or (layer1_outputs(4370));
    layer2_outputs(2644) <= '0';
    layer2_outputs(2645) <= not((layer1_outputs(3392)) and (layer1_outputs(3173)));
    layer2_outputs(2646) <= not((layer1_outputs(5027)) and (layer1_outputs(4098)));
    layer2_outputs(2647) <= not(layer1_outputs(1197)) or (layer1_outputs(651));
    layer2_outputs(2648) <= layer1_outputs(1413);
    layer2_outputs(2649) <= not((layer1_outputs(601)) and (layer1_outputs(123)));
    layer2_outputs(2650) <= layer1_outputs(2086);
    layer2_outputs(2651) <= (layer1_outputs(1833)) or (layer1_outputs(3899));
    layer2_outputs(2652) <= '0';
    layer2_outputs(2653) <= not(layer1_outputs(626));
    layer2_outputs(2654) <= (layer1_outputs(3604)) and (layer1_outputs(3574));
    layer2_outputs(2655) <= not(layer1_outputs(193)) or (layer1_outputs(2891));
    layer2_outputs(2656) <= not(layer1_outputs(3510));
    layer2_outputs(2657) <= layer1_outputs(3512);
    layer2_outputs(2658) <= '0';
    layer2_outputs(2659) <= (layer1_outputs(617)) and (layer1_outputs(5040));
    layer2_outputs(2660) <= '1';
    layer2_outputs(2661) <= '0';
    layer2_outputs(2662) <= not(layer1_outputs(1368)) or (layer1_outputs(2428));
    layer2_outputs(2663) <= not(layer1_outputs(766)) or (layer1_outputs(2798));
    layer2_outputs(2664) <= (layer1_outputs(363)) and (layer1_outputs(3437));
    layer2_outputs(2665) <= (layer1_outputs(2027)) or (layer1_outputs(2418));
    layer2_outputs(2666) <= (layer1_outputs(2632)) or (layer1_outputs(2548));
    layer2_outputs(2667) <= (layer1_outputs(945)) and (layer1_outputs(426));
    layer2_outputs(2668) <= not(layer1_outputs(3935));
    layer2_outputs(2669) <= '0';
    layer2_outputs(2670) <= not(layer1_outputs(4203));
    layer2_outputs(2671) <= (layer1_outputs(3529)) and (layer1_outputs(1910));
    layer2_outputs(2672) <= not((layer1_outputs(604)) or (layer1_outputs(5098)));
    layer2_outputs(2673) <= '1';
    layer2_outputs(2674) <= '1';
    layer2_outputs(2675) <= (layer1_outputs(1919)) and not (layer1_outputs(4436));
    layer2_outputs(2676) <= not(layer1_outputs(4127)) or (layer1_outputs(1804));
    layer2_outputs(2677) <= not(layer1_outputs(108));
    layer2_outputs(2678) <= (layer1_outputs(3241)) and (layer1_outputs(2500));
    layer2_outputs(2679) <= layer1_outputs(3431);
    layer2_outputs(2680) <= (layer1_outputs(1553)) and not (layer1_outputs(3051));
    layer2_outputs(2681) <= not(layer1_outputs(478)) or (layer1_outputs(714));
    layer2_outputs(2682) <= layer1_outputs(4500);
    layer2_outputs(2683) <= not(layer1_outputs(4100));
    layer2_outputs(2684) <= '1';
    layer2_outputs(2685) <= (layer1_outputs(3621)) and not (layer1_outputs(3312));
    layer2_outputs(2686) <= (layer1_outputs(3222)) or (layer1_outputs(2722));
    layer2_outputs(2687) <= (layer1_outputs(1219)) and not (layer1_outputs(306));
    layer2_outputs(2688) <= not((layer1_outputs(4731)) xor (layer1_outputs(3251)));
    layer2_outputs(2689) <= (layer1_outputs(900)) and not (layer1_outputs(982));
    layer2_outputs(2690) <= not(layer1_outputs(1095)) or (layer1_outputs(42));
    layer2_outputs(2691) <= (layer1_outputs(3518)) and (layer1_outputs(3384));
    layer2_outputs(2692) <= (layer1_outputs(4968)) and not (layer1_outputs(3964));
    layer2_outputs(2693) <= '0';
    layer2_outputs(2694) <= not((layer1_outputs(3309)) or (layer1_outputs(4565)));
    layer2_outputs(2695) <= not(layer1_outputs(3860)) or (layer1_outputs(4493));
    layer2_outputs(2696) <= (layer1_outputs(3129)) and (layer1_outputs(2351));
    layer2_outputs(2697) <= (layer1_outputs(1999)) or (layer1_outputs(361));
    layer2_outputs(2698) <= not(layer1_outputs(288)) or (layer1_outputs(4878));
    layer2_outputs(2699) <= not(layer1_outputs(4258)) or (layer1_outputs(3973));
    layer2_outputs(2700) <= layer1_outputs(428);
    layer2_outputs(2701) <= not(layer1_outputs(1450)) or (layer1_outputs(1331));
    layer2_outputs(2702) <= (layer1_outputs(1155)) and (layer1_outputs(4750));
    layer2_outputs(2703) <= (layer1_outputs(2164)) and not (layer1_outputs(4778));
    layer2_outputs(2704) <= (layer1_outputs(4784)) and not (layer1_outputs(1071));
    layer2_outputs(2705) <= (layer1_outputs(4095)) and not (layer1_outputs(637));
    layer2_outputs(2706) <= (layer1_outputs(4472)) or (layer1_outputs(1418));
    layer2_outputs(2707) <= not(layer1_outputs(2104)) or (layer1_outputs(3974));
    layer2_outputs(2708) <= not(layer1_outputs(2370));
    layer2_outputs(2709) <= not(layer1_outputs(1468)) or (layer1_outputs(3798));
    layer2_outputs(2710) <= not(layer1_outputs(2801));
    layer2_outputs(2711) <= (layer1_outputs(1953)) and not (layer1_outputs(2981));
    layer2_outputs(2712) <= '0';
    layer2_outputs(2713) <= (layer1_outputs(437)) and not (layer1_outputs(2807));
    layer2_outputs(2714) <= not((layer1_outputs(3344)) and (layer1_outputs(2246)));
    layer2_outputs(2715) <= (layer1_outputs(4434)) or (layer1_outputs(542));
    layer2_outputs(2716) <= (layer1_outputs(1124)) and (layer1_outputs(4978));
    layer2_outputs(2717) <= layer1_outputs(3085);
    layer2_outputs(2718) <= layer1_outputs(917);
    layer2_outputs(2719) <= '0';
    layer2_outputs(2720) <= '0';
    layer2_outputs(2721) <= '0';
    layer2_outputs(2722) <= (layer1_outputs(1817)) and (layer1_outputs(133));
    layer2_outputs(2723) <= not(layer1_outputs(4295)) or (layer1_outputs(1838));
    layer2_outputs(2724) <= not(layer1_outputs(1046)) or (layer1_outputs(2268));
    layer2_outputs(2725) <= '1';
    layer2_outputs(2726) <= '1';
    layer2_outputs(2727) <= not((layer1_outputs(3357)) and (layer1_outputs(4898)));
    layer2_outputs(2728) <= not(layer1_outputs(1823)) or (layer1_outputs(1472));
    layer2_outputs(2729) <= '0';
    layer2_outputs(2730) <= (layer1_outputs(256)) or (layer1_outputs(4057));
    layer2_outputs(2731) <= (layer1_outputs(2880)) or (layer1_outputs(2297));
    layer2_outputs(2732) <= (layer1_outputs(3941)) and not (layer1_outputs(4792));
    layer2_outputs(2733) <= (layer1_outputs(3597)) and not (layer1_outputs(4789));
    layer2_outputs(2734) <= not(layer1_outputs(953));
    layer2_outputs(2735) <= '1';
    layer2_outputs(2736) <= not((layer1_outputs(3022)) and (layer1_outputs(4585)));
    layer2_outputs(2737) <= (layer1_outputs(2802)) and not (layer1_outputs(4012));
    layer2_outputs(2738) <= (layer1_outputs(2017)) xor (layer1_outputs(1304));
    layer2_outputs(2739) <= (layer1_outputs(4415)) and not (layer1_outputs(4500));
    layer2_outputs(2740) <= not((layer1_outputs(253)) and (layer1_outputs(3021)));
    layer2_outputs(2741) <= '1';
    layer2_outputs(2742) <= not(layer1_outputs(2039));
    layer2_outputs(2743) <= (layer1_outputs(3488)) and not (layer1_outputs(3579));
    layer2_outputs(2744) <= (layer1_outputs(3642)) and (layer1_outputs(4274));
    layer2_outputs(2745) <= '0';
    layer2_outputs(2746) <= not(layer1_outputs(3837));
    layer2_outputs(2747) <= layer1_outputs(898);
    layer2_outputs(2748) <= layer1_outputs(1021);
    layer2_outputs(2749) <= '0';
    layer2_outputs(2750) <= '1';
    layer2_outputs(2751) <= not(layer1_outputs(4734)) or (layer1_outputs(3293));
    layer2_outputs(2752) <= '1';
    layer2_outputs(2753) <= (layer1_outputs(4162)) and not (layer1_outputs(135));
    layer2_outputs(2754) <= not((layer1_outputs(2984)) xor (layer1_outputs(2216)));
    layer2_outputs(2755) <= '0';
    layer2_outputs(2756) <= layer1_outputs(3449);
    layer2_outputs(2757) <= not(layer1_outputs(4257));
    layer2_outputs(2758) <= (layer1_outputs(2659)) or (layer1_outputs(4260));
    layer2_outputs(2759) <= layer1_outputs(3999);
    layer2_outputs(2760) <= '0';
    layer2_outputs(2761) <= '1';
    layer2_outputs(2762) <= '0';
    layer2_outputs(2763) <= (layer1_outputs(2765)) or (layer1_outputs(4848));
    layer2_outputs(2764) <= not(layer1_outputs(2437));
    layer2_outputs(2765) <= (layer1_outputs(4595)) or (layer1_outputs(2024));
    layer2_outputs(2766) <= (layer1_outputs(4364)) and not (layer1_outputs(883));
    layer2_outputs(2767) <= (layer1_outputs(259)) and not (layer1_outputs(1193));
    layer2_outputs(2768) <= (layer1_outputs(3933)) and not (layer1_outputs(4783));
    layer2_outputs(2769) <= (layer1_outputs(2471)) and not (layer1_outputs(2654));
    layer2_outputs(2770) <= not((layer1_outputs(4824)) xor (layer1_outputs(2047)));
    layer2_outputs(2771) <= '0';
    layer2_outputs(2772) <= '1';
    layer2_outputs(2773) <= (layer1_outputs(2681)) and not (layer1_outputs(2561));
    layer2_outputs(2774) <= (layer1_outputs(4350)) and not (layer1_outputs(4913));
    layer2_outputs(2775) <= (layer1_outputs(2276)) and not (layer1_outputs(1753));
    layer2_outputs(2776) <= layer1_outputs(4880);
    layer2_outputs(2777) <= not(layer1_outputs(3183));
    layer2_outputs(2778) <= (layer1_outputs(3234)) or (layer1_outputs(4578));
    layer2_outputs(2779) <= (layer1_outputs(4020)) and not (layer1_outputs(877));
    layer2_outputs(2780) <= (layer1_outputs(156)) or (layer1_outputs(888));
    layer2_outputs(2781) <= (layer1_outputs(3694)) or (layer1_outputs(2849));
    layer2_outputs(2782) <= '0';
    layer2_outputs(2783) <= layer1_outputs(155);
    layer2_outputs(2784) <= not(layer1_outputs(3468)) or (layer1_outputs(1929));
    layer2_outputs(2785) <= not((layer1_outputs(2644)) and (layer1_outputs(1807)));
    layer2_outputs(2786) <= '1';
    layer2_outputs(2787) <= (layer1_outputs(3555)) and (layer1_outputs(3463));
    layer2_outputs(2788) <= (layer1_outputs(74)) xor (layer1_outputs(4804));
    layer2_outputs(2789) <= (layer1_outputs(1493)) and not (layer1_outputs(4000));
    layer2_outputs(2790) <= (layer1_outputs(3426)) or (layer1_outputs(2109));
    layer2_outputs(2791) <= '0';
    layer2_outputs(2792) <= '0';
    layer2_outputs(2793) <= '0';
    layer2_outputs(2794) <= not((layer1_outputs(1136)) xor (layer1_outputs(2482)));
    layer2_outputs(2795) <= '0';
    layer2_outputs(2796) <= layer1_outputs(5083);
    layer2_outputs(2797) <= not(layer1_outputs(4187)) or (layer1_outputs(674));
    layer2_outputs(2798) <= not(layer1_outputs(761));
    layer2_outputs(2799) <= not(layer1_outputs(3704));
    layer2_outputs(2800) <= '1';
    layer2_outputs(2801) <= '0';
    layer2_outputs(2802) <= '1';
    layer2_outputs(2803) <= not((layer1_outputs(2862)) and (layer1_outputs(4725)));
    layer2_outputs(2804) <= layer1_outputs(2187);
    layer2_outputs(2805) <= (layer1_outputs(3294)) and not (layer1_outputs(3811));
    layer2_outputs(2806) <= (layer1_outputs(2308)) and (layer1_outputs(534));
    layer2_outputs(2807) <= not((layer1_outputs(4462)) and (layer1_outputs(134)));
    layer2_outputs(2808) <= '0';
    layer2_outputs(2809) <= '1';
    layer2_outputs(2810) <= (layer1_outputs(4280)) and not (layer1_outputs(2885));
    layer2_outputs(2811) <= not((layer1_outputs(1019)) or (layer1_outputs(4907)));
    layer2_outputs(2812) <= (layer1_outputs(3961)) and not (layer1_outputs(2850));
    layer2_outputs(2813) <= not(layer1_outputs(5000)) or (layer1_outputs(3987));
    layer2_outputs(2814) <= not(layer1_outputs(1830));
    layer2_outputs(2815) <= layer1_outputs(2744);
    layer2_outputs(2816) <= (layer1_outputs(1033)) or (layer1_outputs(320));
    layer2_outputs(2817) <= (layer1_outputs(1160)) and not (layer1_outputs(929));
    layer2_outputs(2818) <= (layer1_outputs(1655)) and not (layer1_outputs(2378));
    layer2_outputs(2819) <= '1';
    layer2_outputs(2820) <= '1';
    layer2_outputs(2821) <= not(layer1_outputs(4080));
    layer2_outputs(2822) <= (layer1_outputs(1706)) and not (layer1_outputs(3799));
    layer2_outputs(2823) <= not((layer1_outputs(2446)) and (layer1_outputs(2194)));
    layer2_outputs(2824) <= layer1_outputs(1265);
    layer2_outputs(2825) <= (layer1_outputs(2313)) and not (layer1_outputs(549));
    layer2_outputs(2826) <= (layer1_outputs(1991)) and not (layer1_outputs(4948));
    layer2_outputs(2827) <= '1';
    layer2_outputs(2828) <= layer1_outputs(4730);
    layer2_outputs(2829) <= not(layer1_outputs(1031));
    layer2_outputs(2830) <= not(layer1_outputs(570));
    layer2_outputs(2831) <= '1';
    layer2_outputs(2832) <= not((layer1_outputs(2552)) or (layer1_outputs(3414)));
    layer2_outputs(2833) <= (layer1_outputs(4443)) and not (layer1_outputs(588));
    layer2_outputs(2834) <= layer1_outputs(2907);
    layer2_outputs(2835) <= '1';
    layer2_outputs(2836) <= not((layer1_outputs(2171)) and (layer1_outputs(1817)));
    layer2_outputs(2837) <= (layer1_outputs(571)) and (layer1_outputs(2079));
    layer2_outputs(2838) <= not((layer1_outputs(1250)) and (layer1_outputs(2728)));
    layer2_outputs(2839) <= not(layer1_outputs(513)) or (layer1_outputs(3699));
    layer2_outputs(2840) <= not(layer1_outputs(162)) or (layer1_outputs(4759));
    layer2_outputs(2841) <= '0';
    layer2_outputs(2842) <= '0';
    layer2_outputs(2843) <= (layer1_outputs(1927)) and not (layer1_outputs(4373));
    layer2_outputs(2844) <= (layer1_outputs(677)) and (layer1_outputs(1408));
    layer2_outputs(2845) <= not(layer1_outputs(87)) or (layer1_outputs(1437));
    layer2_outputs(2846) <= '1';
    layer2_outputs(2847) <= '0';
    layer2_outputs(2848) <= not(layer1_outputs(3750)) or (layer1_outputs(9));
    layer2_outputs(2849) <= not((layer1_outputs(3163)) and (layer1_outputs(4946)));
    layer2_outputs(2850) <= (layer1_outputs(2580)) and not (layer1_outputs(4547));
    layer2_outputs(2851) <= not(layer1_outputs(307)) or (layer1_outputs(2919));
    layer2_outputs(2852) <= not(layer1_outputs(216)) or (layer1_outputs(1248));
    layer2_outputs(2853) <= '1';
    layer2_outputs(2854) <= '1';
    layer2_outputs(2855) <= not(layer1_outputs(2098)) or (layer1_outputs(1829));
    layer2_outputs(2856) <= layer1_outputs(4641);
    layer2_outputs(2857) <= not((layer1_outputs(445)) or (layer1_outputs(1513)));
    layer2_outputs(2858) <= not(layer1_outputs(3378));
    layer2_outputs(2859) <= not((layer1_outputs(2742)) and (layer1_outputs(5101)));
    layer2_outputs(2860) <= not(layer1_outputs(253)) or (layer1_outputs(539));
    layer2_outputs(2861) <= (layer1_outputs(2142)) or (layer1_outputs(3684));
    layer2_outputs(2862) <= '0';
    layer2_outputs(2863) <= '0';
    layer2_outputs(2864) <= '0';
    layer2_outputs(2865) <= not((layer1_outputs(1982)) and (layer1_outputs(4821)));
    layer2_outputs(2866) <= not((layer1_outputs(3399)) and (layer1_outputs(402)));
    layer2_outputs(2867) <= '0';
    layer2_outputs(2868) <= not(layer1_outputs(3649)) or (layer1_outputs(3520));
    layer2_outputs(2869) <= '0';
    layer2_outputs(2870) <= (layer1_outputs(764)) and not (layer1_outputs(2973));
    layer2_outputs(2871) <= '0';
    layer2_outputs(2872) <= (layer1_outputs(2972)) and not (layer1_outputs(2873));
    layer2_outputs(2873) <= (layer1_outputs(3698)) and not (layer1_outputs(241));
    layer2_outputs(2874) <= not(layer1_outputs(3725));
    layer2_outputs(2875) <= (layer1_outputs(3045)) and not (layer1_outputs(4900));
    layer2_outputs(2876) <= (layer1_outputs(1441)) and not (layer1_outputs(3216));
    layer2_outputs(2877) <= '1';
    layer2_outputs(2878) <= not((layer1_outputs(502)) and (layer1_outputs(4444)));
    layer2_outputs(2879) <= not(layer1_outputs(1964));
    layer2_outputs(2880) <= '0';
    layer2_outputs(2881) <= not((layer1_outputs(1401)) and (layer1_outputs(4795)));
    layer2_outputs(2882) <= not(layer1_outputs(4215));
    layer2_outputs(2883) <= not(layer1_outputs(1898)) or (layer1_outputs(3643));
    layer2_outputs(2884) <= not(layer1_outputs(4110)) or (layer1_outputs(2333));
    layer2_outputs(2885) <= '0';
    layer2_outputs(2886) <= '1';
    layer2_outputs(2887) <= not((layer1_outputs(30)) and (layer1_outputs(3802)));
    layer2_outputs(2888) <= (layer1_outputs(3224)) or (layer1_outputs(606));
    layer2_outputs(2889) <= layer1_outputs(1912);
    layer2_outputs(2890) <= not(layer1_outputs(2437));
    layer2_outputs(2891) <= (layer1_outputs(4545)) and not (layer1_outputs(2392));
    layer2_outputs(2892) <= not((layer1_outputs(4714)) or (layer1_outputs(3369)));
    layer2_outputs(2893) <= '1';
    layer2_outputs(2894) <= (layer1_outputs(4266)) and not (layer1_outputs(415));
    layer2_outputs(2895) <= (layer1_outputs(124)) or (layer1_outputs(4577));
    layer2_outputs(2896) <= not((layer1_outputs(3680)) and (layer1_outputs(3585)));
    layer2_outputs(2897) <= not((layer1_outputs(2474)) or (layer1_outputs(206)));
    layer2_outputs(2898) <= not(layer1_outputs(976));
    layer2_outputs(2899) <= (layer1_outputs(1062)) or (layer1_outputs(4081));
    layer2_outputs(2900) <= '0';
    layer2_outputs(2901) <= '1';
    layer2_outputs(2902) <= layer1_outputs(826);
    layer2_outputs(2903) <= (layer1_outputs(3199)) and not (layer1_outputs(1944));
    layer2_outputs(2904) <= not((layer1_outputs(3132)) and (layer1_outputs(3064)));
    layer2_outputs(2905) <= not((layer1_outputs(2966)) or (layer1_outputs(3942)));
    layer2_outputs(2906) <= '0';
    layer2_outputs(2907) <= not((layer1_outputs(4885)) or (layer1_outputs(4545)));
    layer2_outputs(2908) <= not((layer1_outputs(3832)) or (layer1_outputs(809)));
    layer2_outputs(2909) <= not(layer1_outputs(2246));
    layer2_outputs(2910) <= '1';
    layer2_outputs(2911) <= layer1_outputs(1201);
    layer2_outputs(2912) <= '0';
    layer2_outputs(2913) <= (layer1_outputs(4485)) or (layer1_outputs(584));
    layer2_outputs(2914) <= not((layer1_outputs(3202)) and (layer1_outputs(5035)));
    layer2_outputs(2915) <= layer1_outputs(3498);
    layer2_outputs(2916) <= (layer1_outputs(3036)) and (layer1_outputs(4389));
    layer2_outputs(2917) <= '1';
    layer2_outputs(2918) <= not(layer1_outputs(4437)) or (layer1_outputs(2145));
    layer2_outputs(2919) <= '1';
    layer2_outputs(2920) <= '1';
    layer2_outputs(2921) <= not(layer1_outputs(1203)) or (layer1_outputs(2765));
    layer2_outputs(2922) <= not(layer1_outputs(1960));
    layer2_outputs(2923) <= layer1_outputs(702);
    layer2_outputs(2924) <= '0';
    layer2_outputs(2925) <= not(layer1_outputs(4314)) or (layer1_outputs(4004));
    layer2_outputs(2926) <= (layer1_outputs(3476)) and not (layer1_outputs(708));
    layer2_outputs(2927) <= (layer1_outputs(1137)) or (layer1_outputs(2915));
    layer2_outputs(2928) <= '1';
    layer2_outputs(2929) <= not(layer1_outputs(3619));
    layer2_outputs(2930) <= layer1_outputs(4711);
    layer2_outputs(2931) <= (layer1_outputs(4677)) and not (layer1_outputs(3969));
    layer2_outputs(2932) <= '0';
    layer2_outputs(2933) <= '1';
    layer2_outputs(2934) <= layer1_outputs(3729);
    layer2_outputs(2935) <= (layer1_outputs(34)) and not (layer1_outputs(2383));
    layer2_outputs(2936) <= not(layer1_outputs(2457));
    layer2_outputs(2937) <= '1';
    layer2_outputs(2938) <= '1';
    layer2_outputs(2939) <= '0';
    layer2_outputs(2940) <= '1';
    layer2_outputs(2941) <= '0';
    layer2_outputs(2942) <= not(layer1_outputs(2248));
    layer2_outputs(2943) <= not(layer1_outputs(4878));
    layer2_outputs(2944) <= (layer1_outputs(4018)) xor (layer1_outputs(623));
    layer2_outputs(2945) <= (layer1_outputs(3559)) or (layer1_outputs(1391));
    layer2_outputs(2946) <= not(layer1_outputs(5094));
    layer2_outputs(2947) <= not((layer1_outputs(1961)) xor (layer1_outputs(1931)));
    layer2_outputs(2948) <= not((layer1_outputs(1185)) and (layer1_outputs(686)));
    layer2_outputs(2949) <= layer1_outputs(611);
    layer2_outputs(2950) <= not(layer1_outputs(4899)) or (layer1_outputs(3400));
    layer2_outputs(2951) <= not((layer1_outputs(2504)) and (layer1_outputs(3925)));
    layer2_outputs(2952) <= layer1_outputs(117);
    layer2_outputs(2953) <= not(layer1_outputs(1442)) or (layer1_outputs(2103));
    layer2_outputs(2954) <= not(layer1_outputs(1916));
    layer2_outputs(2955) <= not(layer1_outputs(5061)) or (layer1_outputs(2947));
    layer2_outputs(2956) <= '1';
    layer2_outputs(2957) <= not((layer1_outputs(2383)) or (layer1_outputs(242)));
    layer2_outputs(2958) <= not((layer1_outputs(2673)) or (layer1_outputs(1041)));
    layer2_outputs(2959) <= not((layer1_outputs(4547)) and (layer1_outputs(3162)));
    layer2_outputs(2960) <= layer1_outputs(3149);
    layer2_outputs(2961) <= '0';
    layer2_outputs(2962) <= (layer1_outputs(1973)) or (layer1_outputs(2784));
    layer2_outputs(2963) <= '0';
    layer2_outputs(2964) <= '0';
    layer2_outputs(2965) <= '1';
    layer2_outputs(2966) <= layer1_outputs(4866);
    layer2_outputs(2967) <= '0';
    layer2_outputs(2968) <= '1';
    layer2_outputs(2969) <= not(layer1_outputs(2682)) or (layer1_outputs(4403));
    layer2_outputs(2970) <= (layer1_outputs(1184)) and not (layer1_outputs(1164));
    layer2_outputs(2971) <= not(layer1_outputs(393));
    layer2_outputs(2972) <= not(layer1_outputs(207)) or (layer1_outputs(1238));
    layer2_outputs(2973) <= not(layer1_outputs(4131)) or (layer1_outputs(4832));
    layer2_outputs(2974) <= (layer1_outputs(4136)) and (layer1_outputs(4963));
    layer2_outputs(2975) <= not(layer1_outputs(127)) or (layer1_outputs(966));
    layer2_outputs(2976) <= (layer1_outputs(967)) and not (layer1_outputs(3997));
    layer2_outputs(2977) <= (layer1_outputs(604)) and not (layer1_outputs(2141));
    layer2_outputs(2978) <= not((layer1_outputs(4095)) or (layer1_outputs(66)));
    layer2_outputs(2979) <= not(layer1_outputs(4655));
    layer2_outputs(2980) <= not(layer1_outputs(537)) or (layer1_outputs(1136));
    layer2_outputs(2981) <= layer1_outputs(689);
    layer2_outputs(2982) <= '0';
    layer2_outputs(2983) <= (layer1_outputs(4871)) and (layer1_outputs(3229));
    layer2_outputs(2984) <= not(layer1_outputs(3102));
    layer2_outputs(2985) <= (layer1_outputs(1788)) and not (layer1_outputs(4073));
    layer2_outputs(2986) <= not(layer1_outputs(478)) or (layer1_outputs(3797));
    layer2_outputs(2987) <= (layer1_outputs(4453)) and not (layer1_outputs(1751));
    layer2_outputs(2988) <= (layer1_outputs(4847)) and (layer1_outputs(3870));
    layer2_outputs(2989) <= not(layer1_outputs(4666));
    layer2_outputs(2990) <= (layer1_outputs(4873)) and (layer1_outputs(410));
    layer2_outputs(2991) <= not((layer1_outputs(297)) or (layer1_outputs(1333)));
    layer2_outputs(2992) <= '0';
    layer2_outputs(2993) <= (layer1_outputs(257)) and not (layer1_outputs(937));
    layer2_outputs(2994) <= layer1_outputs(4330);
    layer2_outputs(2995) <= not(layer1_outputs(1625)) or (layer1_outputs(793));
    layer2_outputs(2996) <= not(layer1_outputs(4747)) or (layer1_outputs(2565));
    layer2_outputs(2997) <= (layer1_outputs(1184)) and (layer1_outputs(1556));
    layer2_outputs(2998) <= (layer1_outputs(690)) and (layer1_outputs(3324));
    layer2_outputs(2999) <= '1';
    layer2_outputs(3000) <= (layer1_outputs(2010)) xor (layer1_outputs(2955));
    layer2_outputs(3001) <= '0';
    layer2_outputs(3002) <= (layer1_outputs(507)) and not (layer1_outputs(442));
    layer2_outputs(3003) <= '0';
    layer2_outputs(3004) <= (layer1_outputs(1482)) and (layer1_outputs(1791));
    layer2_outputs(3005) <= (layer1_outputs(4216)) and not (layer1_outputs(130));
    layer2_outputs(3006) <= layer1_outputs(1531);
    layer2_outputs(3007) <= not(layer1_outputs(3392)) or (layer1_outputs(3680));
    layer2_outputs(3008) <= layer1_outputs(3275);
    layer2_outputs(3009) <= (layer1_outputs(2484)) and not (layer1_outputs(1234));
    layer2_outputs(3010) <= not(layer1_outputs(2883)) or (layer1_outputs(208));
    layer2_outputs(3011) <= not(layer1_outputs(3025)) or (layer1_outputs(214));
    layer2_outputs(3012) <= layer1_outputs(4533);
    layer2_outputs(3013) <= not((layer1_outputs(2639)) or (layer1_outputs(1065)));
    layer2_outputs(3014) <= '1';
    layer2_outputs(3015) <= not(layer1_outputs(4340));
    layer2_outputs(3016) <= not(layer1_outputs(2379));
    layer2_outputs(3017) <= '1';
    layer2_outputs(3018) <= not(layer1_outputs(110));
    layer2_outputs(3019) <= (layer1_outputs(4539)) and not (layer1_outputs(3503));
    layer2_outputs(3020) <= layer1_outputs(2949);
    layer2_outputs(3021) <= not(layer1_outputs(3499));
    layer2_outputs(3022) <= (layer1_outputs(3222)) and not (layer1_outputs(2305));
    layer2_outputs(3023) <= '0';
    layer2_outputs(3024) <= '0';
    layer2_outputs(3025) <= not(layer1_outputs(4166)) or (layer1_outputs(3917));
    layer2_outputs(3026) <= '1';
    layer2_outputs(3027) <= not(layer1_outputs(1994)) or (layer1_outputs(3070));
    layer2_outputs(3028) <= (layer1_outputs(1542)) and not (layer1_outputs(2366));
    layer2_outputs(3029) <= '1';
    layer2_outputs(3030) <= not(layer1_outputs(3689)) or (layer1_outputs(456));
    layer2_outputs(3031) <= not(layer1_outputs(1647));
    layer2_outputs(3032) <= not(layer1_outputs(3901));
    layer2_outputs(3033) <= not(layer1_outputs(3379)) or (layer1_outputs(4024));
    layer2_outputs(3034) <= not((layer1_outputs(182)) or (layer1_outputs(3443)));
    layer2_outputs(3035) <= (layer1_outputs(424)) and not (layer1_outputs(721));
    layer2_outputs(3036) <= not((layer1_outputs(4531)) xor (layer1_outputs(2521)));
    layer2_outputs(3037) <= (layer1_outputs(4398)) and not (layer1_outputs(1303));
    layer2_outputs(3038) <= layer1_outputs(1226);
    layer2_outputs(3039) <= '1';
    layer2_outputs(3040) <= not(layer1_outputs(2517)) or (layer1_outputs(3880));
    layer2_outputs(3041) <= (layer1_outputs(1696)) and (layer1_outputs(1265));
    layer2_outputs(3042) <= '1';
    layer2_outputs(3043) <= (layer1_outputs(4328)) or (layer1_outputs(4243));
    layer2_outputs(3044) <= not((layer1_outputs(3416)) or (layer1_outputs(3040)));
    layer2_outputs(3045) <= (layer1_outputs(860)) and (layer1_outputs(1414));
    layer2_outputs(3046) <= '1';
    layer2_outputs(3047) <= layer1_outputs(4222);
    layer2_outputs(3048) <= not(layer1_outputs(4962)) or (layer1_outputs(751));
    layer2_outputs(3049) <= (layer1_outputs(585)) or (layer1_outputs(2762));
    layer2_outputs(3050) <= not((layer1_outputs(3041)) and (layer1_outputs(582)));
    layer2_outputs(3051) <= '1';
    layer2_outputs(3052) <= '1';
    layer2_outputs(3053) <= not((layer1_outputs(4829)) and (layer1_outputs(4223)));
    layer2_outputs(3054) <= not(layer1_outputs(2041)) or (layer1_outputs(4887));
    layer2_outputs(3055) <= not(layer1_outputs(4169));
    layer2_outputs(3056) <= layer1_outputs(2514);
    layer2_outputs(3057) <= not(layer1_outputs(2224)) or (layer1_outputs(1957));
    layer2_outputs(3058) <= not(layer1_outputs(2132)) or (layer1_outputs(2892));
    layer2_outputs(3059) <= '0';
    layer2_outputs(3060) <= '0';
    layer2_outputs(3061) <= layer1_outputs(1424);
    layer2_outputs(3062) <= not((layer1_outputs(11)) and (layer1_outputs(1562)));
    layer2_outputs(3063) <= not((layer1_outputs(1528)) or (layer1_outputs(2225)));
    layer2_outputs(3064) <= (layer1_outputs(3886)) or (layer1_outputs(4786));
    layer2_outputs(3065) <= not((layer1_outputs(379)) and (layer1_outputs(1435)));
    layer2_outputs(3066) <= not(layer1_outputs(3913));
    layer2_outputs(3067) <= '1';
    layer2_outputs(3068) <= not((layer1_outputs(361)) or (layer1_outputs(4417)));
    layer2_outputs(3069) <= (layer1_outputs(2729)) and not (layer1_outputs(2749));
    layer2_outputs(3070) <= (layer1_outputs(207)) and not (layer1_outputs(3951));
    layer2_outputs(3071) <= not(layer1_outputs(4569));
    layer2_outputs(3072) <= (layer1_outputs(1346)) and not (layer1_outputs(3248));
    layer2_outputs(3073) <= '1';
    layer2_outputs(3074) <= layer1_outputs(4865);
    layer2_outputs(3075) <= not((layer1_outputs(3232)) and (layer1_outputs(2325)));
    layer2_outputs(3076) <= not((layer1_outputs(989)) and (layer1_outputs(291)));
    layer2_outputs(3077) <= '0';
    layer2_outputs(3078) <= '0';
    layer2_outputs(3079) <= not(layer1_outputs(3854));
    layer2_outputs(3080) <= '0';
    layer2_outputs(3081) <= (layer1_outputs(730)) xor (layer1_outputs(1455));
    layer2_outputs(3082) <= not((layer1_outputs(3238)) and (layer1_outputs(5113)));
    layer2_outputs(3083) <= '0';
    layer2_outputs(3084) <= not(layer1_outputs(4870)) or (layer1_outputs(687));
    layer2_outputs(3085) <= '0';
    layer2_outputs(3086) <= (layer1_outputs(229)) or (layer1_outputs(1357));
    layer2_outputs(3087) <= layer1_outputs(2467);
    layer2_outputs(3088) <= layer1_outputs(2681);
    layer2_outputs(3089) <= '1';
    layer2_outputs(3090) <= not((layer1_outputs(1773)) and (layer1_outputs(3982)));
    layer2_outputs(3091) <= '0';
    layer2_outputs(3092) <= (layer1_outputs(469)) and not (layer1_outputs(4577));
    layer2_outputs(3093) <= (layer1_outputs(2219)) or (layer1_outputs(3380));
    layer2_outputs(3094) <= not((layer1_outputs(4089)) and (layer1_outputs(462)));
    layer2_outputs(3095) <= layer1_outputs(240);
    layer2_outputs(3096) <= '0';
    layer2_outputs(3097) <= '0';
    layer2_outputs(3098) <= not(layer1_outputs(2092)) or (layer1_outputs(3706));
    layer2_outputs(3099) <= not(layer1_outputs(3457));
    layer2_outputs(3100) <= not(layer1_outputs(611)) or (layer1_outputs(4610));
    layer2_outputs(3101) <= not(layer1_outputs(306));
    layer2_outputs(3102) <= not(layer1_outputs(44));
    layer2_outputs(3103) <= '0';
    layer2_outputs(3104) <= not((layer1_outputs(3100)) or (layer1_outputs(794)));
    layer2_outputs(3105) <= not((layer1_outputs(3033)) or (layer1_outputs(3792)));
    layer2_outputs(3106) <= '1';
    layer2_outputs(3107) <= not(layer1_outputs(1121));
    layer2_outputs(3108) <= '0';
    layer2_outputs(3109) <= not(layer1_outputs(343)) or (layer1_outputs(720));
    layer2_outputs(3110) <= not((layer1_outputs(0)) or (layer1_outputs(3179)));
    layer2_outputs(3111) <= not(layer1_outputs(997)) or (layer1_outputs(4783));
    layer2_outputs(3112) <= '1';
    layer2_outputs(3113) <= '0';
    layer2_outputs(3114) <= (layer1_outputs(1515)) and not (layer1_outputs(4432));
    layer2_outputs(3115) <= (layer1_outputs(3674)) xor (layer1_outputs(392));
    layer2_outputs(3116) <= not((layer1_outputs(3171)) and (layer1_outputs(3922)));
    layer2_outputs(3117) <= '1';
    layer2_outputs(3118) <= layer1_outputs(1321);
    layer2_outputs(3119) <= layer1_outputs(4217);
    layer2_outputs(3120) <= '1';
    layer2_outputs(3121) <= '0';
    layer2_outputs(3122) <= not((layer1_outputs(818)) or (layer1_outputs(1211)));
    layer2_outputs(3123) <= not(layer1_outputs(4593)) or (layer1_outputs(1317));
    layer2_outputs(3124) <= layer1_outputs(2914);
    layer2_outputs(3125) <= '1';
    layer2_outputs(3126) <= (layer1_outputs(2297)) or (layer1_outputs(3991));
    layer2_outputs(3127) <= (layer1_outputs(2683)) and (layer1_outputs(569));
    layer2_outputs(3128) <= (layer1_outputs(1364)) and not (layer1_outputs(2624));
    layer2_outputs(3129) <= not(layer1_outputs(4238)) or (layer1_outputs(1456));
    layer2_outputs(3130) <= not((layer1_outputs(3558)) or (layer1_outputs(3980)));
    layer2_outputs(3131) <= not(layer1_outputs(1858));
    layer2_outputs(3132) <= (layer1_outputs(2752)) and not (layer1_outputs(2435));
    layer2_outputs(3133) <= not(layer1_outputs(983)) or (layer1_outputs(2068));
    layer2_outputs(3134) <= not(layer1_outputs(519));
    layer2_outputs(3135) <= not(layer1_outputs(4972));
    layer2_outputs(3136) <= (layer1_outputs(116)) and (layer1_outputs(3770));
    layer2_outputs(3137) <= (layer1_outputs(2131)) and (layer1_outputs(1623));
    layer2_outputs(3138) <= not((layer1_outputs(4295)) and (layer1_outputs(287)));
    layer2_outputs(3139) <= '1';
    layer2_outputs(3140) <= '0';
    layer2_outputs(3141) <= not((layer1_outputs(2370)) or (layer1_outputs(2402)));
    layer2_outputs(3142) <= '1';
    layer2_outputs(3143) <= (layer1_outputs(2795)) and not (layer1_outputs(4807));
    layer2_outputs(3144) <= layer1_outputs(4464);
    layer2_outputs(3145) <= layer1_outputs(1195);
    layer2_outputs(3146) <= (layer1_outputs(4306)) xor (layer1_outputs(1285));
    layer2_outputs(3147) <= layer1_outputs(2289);
    layer2_outputs(3148) <= not((layer1_outputs(2773)) and (layer1_outputs(3563)));
    layer2_outputs(3149) <= not((layer1_outputs(2577)) or (layer1_outputs(1018)));
    layer2_outputs(3150) <= not((layer1_outputs(2341)) or (layer1_outputs(3326)));
    layer2_outputs(3151) <= not((layer1_outputs(1690)) or (layer1_outputs(1239)));
    layer2_outputs(3152) <= (layer1_outputs(1315)) and not (layer1_outputs(3403));
    layer2_outputs(3153) <= not(layer1_outputs(2149));
    layer2_outputs(3154) <= not(layer1_outputs(3225));
    layer2_outputs(3155) <= '0';
    layer2_outputs(3156) <= not(layer1_outputs(72));
    layer2_outputs(3157) <= (layer1_outputs(283)) or (layer1_outputs(2865));
    layer2_outputs(3158) <= not(layer1_outputs(3909)) or (layer1_outputs(3543));
    layer2_outputs(3159) <= not(layer1_outputs(1703));
    layer2_outputs(3160) <= '0';
    layer2_outputs(3161) <= not(layer1_outputs(2553)) or (layer1_outputs(843));
    layer2_outputs(3162) <= '1';
    layer2_outputs(3163) <= '1';
    layer2_outputs(3164) <= not((layer1_outputs(1206)) or (layer1_outputs(4063)));
    layer2_outputs(3165) <= '1';
    layer2_outputs(3166) <= (layer1_outputs(204)) and (layer1_outputs(4808));
    layer2_outputs(3167) <= layer1_outputs(2099);
    layer2_outputs(3168) <= layer1_outputs(4176);
    layer2_outputs(3169) <= layer1_outputs(2869);
    layer2_outputs(3170) <= (layer1_outputs(2096)) and not (layer1_outputs(1801));
    layer2_outputs(3171) <= layer1_outputs(4894);
    layer2_outputs(3172) <= (layer1_outputs(2882)) and not (layer1_outputs(2102));
    layer2_outputs(3173) <= '1';
    layer2_outputs(3174) <= not((layer1_outputs(195)) or (layer1_outputs(3763)));
    layer2_outputs(3175) <= '0';
    layer2_outputs(3176) <= not(layer1_outputs(3958)) or (layer1_outputs(4589));
    layer2_outputs(3177) <= not((layer1_outputs(80)) or (layer1_outputs(2129)));
    layer2_outputs(3178) <= not((layer1_outputs(3328)) or (layer1_outputs(3009)));
    layer2_outputs(3179) <= '1';
    layer2_outputs(3180) <= (layer1_outputs(1092)) and not (layer1_outputs(2494));
    layer2_outputs(3181) <= (layer1_outputs(1187)) or (layer1_outputs(4617));
    layer2_outputs(3182) <= '1';
    layer2_outputs(3183) <= not(layer1_outputs(501));
    layer2_outputs(3184) <= layer1_outputs(4407);
    layer2_outputs(3185) <= not(layer1_outputs(2053));
    layer2_outputs(3186) <= '1';
    layer2_outputs(3187) <= '0';
    layer2_outputs(3188) <= (layer1_outputs(3827)) and not (layer1_outputs(4393));
    layer2_outputs(3189) <= (layer1_outputs(1917)) and not (layer1_outputs(3157));
    layer2_outputs(3190) <= (layer1_outputs(2890)) and not (layer1_outputs(2179));
    layer2_outputs(3191) <= (layer1_outputs(1942)) or (layer1_outputs(562));
    layer2_outputs(3192) <= (layer1_outputs(3016)) and not (layer1_outputs(1362));
    layer2_outputs(3193) <= not(layer1_outputs(1837)) or (layer1_outputs(2401));
    layer2_outputs(3194) <= '1';
    layer2_outputs(3195) <= layer1_outputs(4030);
    layer2_outputs(3196) <= (layer1_outputs(1322)) and not (layer1_outputs(4822));
    layer2_outputs(3197) <= not((layer1_outputs(2412)) and (layer1_outputs(1355)));
    layer2_outputs(3198) <= (layer1_outputs(807)) and not (layer1_outputs(405));
    layer2_outputs(3199) <= (layer1_outputs(1078)) and not (layer1_outputs(1662));
    layer2_outputs(3200) <= not(layer1_outputs(1486)) or (layer1_outputs(3825));
    layer2_outputs(3201) <= (layer1_outputs(2823)) and not (layer1_outputs(1546));
    layer2_outputs(3202) <= (layer1_outputs(138)) or (layer1_outputs(3297));
    layer2_outputs(3203) <= not(layer1_outputs(266)) or (layer1_outputs(4600));
    layer2_outputs(3204) <= '0';
    layer2_outputs(3205) <= '0';
    layer2_outputs(3206) <= not((layer1_outputs(1431)) and (layer1_outputs(1771)));
    layer2_outputs(3207) <= not(layer1_outputs(3303)) or (layer1_outputs(849));
    layer2_outputs(3208) <= '1';
    layer2_outputs(3209) <= '1';
    layer2_outputs(3210) <= '0';
    layer2_outputs(3211) <= (layer1_outputs(467)) and (layer1_outputs(4806));
    layer2_outputs(3212) <= not(layer1_outputs(4250)) or (layer1_outputs(2352));
    layer2_outputs(3213) <= '0';
    layer2_outputs(3214) <= layer1_outputs(345);
    layer2_outputs(3215) <= (layer1_outputs(2202)) and (layer1_outputs(2369));
    layer2_outputs(3216) <= (layer1_outputs(893)) and not (layer1_outputs(312));
    layer2_outputs(3217) <= (layer1_outputs(467)) and not (layer1_outputs(1568));
    layer2_outputs(3218) <= '0';
    layer2_outputs(3219) <= (layer1_outputs(1857)) and not (layer1_outputs(3568));
    layer2_outputs(3220) <= not(layer1_outputs(1154)) or (layer1_outputs(607));
    layer2_outputs(3221) <= (layer1_outputs(1105)) and not (layer1_outputs(2462));
    layer2_outputs(3222) <= (layer1_outputs(828)) and not (layer1_outputs(2845));
    layer2_outputs(3223) <= not(layer1_outputs(4153));
    layer2_outputs(3224) <= not(layer1_outputs(1147));
    layer2_outputs(3225) <= not(layer1_outputs(4040)) or (layer1_outputs(3979));
    layer2_outputs(3226) <= '1';
    layer2_outputs(3227) <= not(layer1_outputs(2538)) or (layer1_outputs(1859));
    layer2_outputs(3228) <= (layer1_outputs(2546)) and (layer1_outputs(1980));
    layer2_outputs(3229) <= '0';
    layer2_outputs(3230) <= (layer1_outputs(3515)) and not (layer1_outputs(2479));
    layer2_outputs(3231) <= '0';
    layer2_outputs(3232) <= not(layer1_outputs(4806)) or (layer1_outputs(3330));
    layer2_outputs(3233) <= (layer1_outputs(3517)) and not (layer1_outputs(3158));
    layer2_outputs(3234) <= (layer1_outputs(2496)) or (layer1_outputs(1299));
    layer2_outputs(3235) <= '0';
    layer2_outputs(3236) <= not((layer1_outputs(3758)) and (layer1_outputs(3549)));
    layer2_outputs(3237) <= (layer1_outputs(833)) and not (layer1_outputs(4621));
    layer2_outputs(3238) <= not((layer1_outputs(823)) and (layer1_outputs(372)));
    layer2_outputs(3239) <= (layer1_outputs(2952)) and (layer1_outputs(4465));
    layer2_outputs(3240) <= (layer1_outputs(1539)) or (layer1_outputs(368));
    layer2_outputs(3241) <= not((layer1_outputs(4322)) xor (layer1_outputs(2228)));
    layer2_outputs(3242) <= not((layer1_outputs(1503)) and (layer1_outputs(1655)));
    layer2_outputs(3243) <= (layer1_outputs(3361)) xor (layer1_outputs(2968));
    layer2_outputs(3244) <= not(layer1_outputs(4058)) or (layer1_outputs(2204));
    layer2_outputs(3245) <= '0';
    layer2_outputs(3246) <= '0';
    layer2_outputs(3247) <= not((layer1_outputs(148)) or (layer1_outputs(983)));
    layer2_outputs(3248) <= '1';
    layer2_outputs(3249) <= not(layer1_outputs(1390)) or (layer1_outputs(1082));
    layer2_outputs(3250) <= layer1_outputs(3815);
    layer2_outputs(3251) <= not((layer1_outputs(509)) and (layer1_outputs(3903)));
    layer2_outputs(3252) <= (layer1_outputs(4528)) or (layer1_outputs(3367));
    layer2_outputs(3253) <= (layer1_outputs(2773)) or (layer1_outputs(1789));
    layer2_outputs(3254) <= not(layer1_outputs(3227));
    layer2_outputs(3255) <= (layer1_outputs(3407)) xor (layer1_outputs(2262));
    layer2_outputs(3256) <= (layer1_outputs(1205)) and (layer1_outputs(1162));
    layer2_outputs(3257) <= (layer1_outputs(4976)) and not (layer1_outputs(1243));
    layer2_outputs(3258) <= '0';
    layer2_outputs(3259) <= (layer1_outputs(4981)) or (layer1_outputs(2533));
    layer2_outputs(3260) <= (layer1_outputs(1597)) and not (layer1_outputs(4679));
    layer2_outputs(3261) <= not(layer1_outputs(2239));
    layer2_outputs(3262) <= not((layer1_outputs(2641)) and (layer1_outputs(4081)));
    layer2_outputs(3263) <= (layer1_outputs(3582)) or (layer1_outputs(1300));
    layer2_outputs(3264) <= not((layer1_outputs(2036)) or (layer1_outputs(2756)));
    layer2_outputs(3265) <= '1';
    layer2_outputs(3266) <= not(layer1_outputs(2518)) or (layer1_outputs(4744));
    layer2_outputs(3267) <= '0';
    layer2_outputs(3268) <= not(layer1_outputs(2790)) or (layer1_outputs(553));
    layer2_outputs(3269) <= '1';
    layer2_outputs(3270) <= '1';
    layer2_outputs(3271) <= '0';
    layer2_outputs(3272) <= not((layer1_outputs(2537)) or (layer1_outputs(1167)));
    layer2_outputs(3273) <= not(layer1_outputs(124));
    layer2_outputs(3274) <= '1';
    layer2_outputs(3275) <= (layer1_outputs(2959)) and not (layer1_outputs(2381));
    layer2_outputs(3276) <= (layer1_outputs(4175)) xor (layer1_outputs(258));
    layer2_outputs(3277) <= layer1_outputs(5031);
    layer2_outputs(3278) <= not(layer1_outputs(3433));
    layer2_outputs(3279) <= layer1_outputs(4902);
    layer2_outputs(3280) <= not(layer1_outputs(103));
    layer2_outputs(3281) <= (layer1_outputs(4264)) and not (layer1_outputs(3782));
    layer2_outputs(3282) <= not(layer1_outputs(1029)) or (layer1_outputs(483));
    layer2_outputs(3283) <= not((layer1_outputs(3784)) or (layer1_outputs(2201)));
    layer2_outputs(3284) <= layer1_outputs(2933);
    layer2_outputs(3285) <= '0';
    layer2_outputs(3286) <= '1';
    layer2_outputs(3287) <= not((layer1_outputs(1354)) and (layer1_outputs(926)));
    layer2_outputs(3288) <= '1';
    layer2_outputs(3289) <= not(layer1_outputs(1851)) or (layer1_outputs(2621));
    layer2_outputs(3290) <= '0';
    layer2_outputs(3291) <= '0';
    layer2_outputs(3292) <= (layer1_outputs(2589)) and (layer1_outputs(5048));
    layer2_outputs(3293) <= not(layer1_outputs(1813));
    layer2_outputs(3294) <= '1';
    layer2_outputs(3295) <= (layer1_outputs(3515)) and (layer1_outputs(4166));
    layer2_outputs(3296) <= (layer1_outputs(4077)) and not (layer1_outputs(261));
    layer2_outputs(3297) <= not(layer1_outputs(201)) or (layer1_outputs(1857));
    layer2_outputs(3298) <= not(layer1_outputs(1043)) or (layer1_outputs(4673));
    layer2_outputs(3299) <= layer1_outputs(743);
    layer2_outputs(3300) <= '1';
    layer2_outputs(3301) <= not(layer1_outputs(1840)) or (layer1_outputs(1013));
    layer2_outputs(3302) <= (layer1_outputs(2384)) and (layer1_outputs(2665));
    layer2_outputs(3303) <= not((layer1_outputs(4394)) and (layer1_outputs(1306)));
    layer2_outputs(3304) <= (layer1_outputs(1368)) and not (layer1_outputs(1579));
    layer2_outputs(3305) <= (layer1_outputs(4645)) or (layer1_outputs(979));
    layer2_outputs(3306) <= '1';
    layer2_outputs(3307) <= not((layer1_outputs(4564)) or (layer1_outputs(4312)));
    layer2_outputs(3308) <= '1';
    layer2_outputs(3309) <= '1';
    layer2_outputs(3310) <= '1';
    layer2_outputs(3311) <= '0';
    layer2_outputs(3312) <= (layer1_outputs(2318)) xor (layer1_outputs(1298));
    layer2_outputs(3313) <= layer1_outputs(1483);
    layer2_outputs(3314) <= not(layer1_outputs(1619));
    layer2_outputs(3315) <= '1';
    layer2_outputs(3316) <= (layer1_outputs(2857)) and (layer1_outputs(1869));
    layer2_outputs(3317) <= (layer1_outputs(241)) and (layer1_outputs(2879));
    layer2_outputs(3318) <= layer1_outputs(4204);
    layer2_outputs(3319) <= layer1_outputs(2525);
    layer2_outputs(3320) <= not(layer1_outputs(2231)) or (layer1_outputs(1493));
    layer2_outputs(3321) <= not((layer1_outputs(1176)) and (layer1_outputs(939)));
    layer2_outputs(3322) <= layer1_outputs(2787);
    layer2_outputs(3323) <= layer1_outputs(2685);
    layer2_outputs(3324) <= not(layer1_outputs(1786)) or (layer1_outputs(3428));
    layer2_outputs(3325) <= not(layer1_outputs(3882)) or (layer1_outputs(940));
    layer2_outputs(3326) <= '0';
    layer2_outputs(3327) <= layer1_outputs(1677);
    layer2_outputs(3328) <= (layer1_outputs(4163)) and not (layer1_outputs(1076));
    layer2_outputs(3329) <= (layer1_outputs(2307)) and not (layer1_outputs(789));
    layer2_outputs(3330) <= '0';
    layer2_outputs(3331) <= not((layer1_outputs(3624)) or (layer1_outputs(4055)));
    layer2_outputs(3332) <= (layer1_outputs(4522)) and not (layer1_outputs(728));
    layer2_outputs(3333) <= not((layer1_outputs(4269)) and (layer1_outputs(3723)));
    layer2_outputs(3334) <= (layer1_outputs(4639)) xor (layer1_outputs(4101));
    layer2_outputs(3335) <= '1';
    layer2_outputs(3336) <= '1';
    layer2_outputs(3337) <= (layer1_outputs(3632)) and not (layer1_outputs(2720));
    layer2_outputs(3338) <= (layer1_outputs(2275)) and not (layer1_outputs(2118));
    layer2_outputs(3339) <= (layer1_outputs(3491)) and not (layer1_outputs(4613));
    layer2_outputs(3340) <= not((layer1_outputs(3735)) and (layer1_outputs(1907)));
    layer2_outputs(3341) <= (layer1_outputs(3059)) and not (layer1_outputs(2002));
    layer2_outputs(3342) <= (layer1_outputs(5105)) and not (layer1_outputs(2449));
    layer2_outputs(3343) <= '1';
    layer2_outputs(3344) <= not(layer1_outputs(4412));
    layer2_outputs(3345) <= layer1_outputs(2423);
    layer2_outputs(3346) <= layer1_outputs(633);
    layer2_outputs(3347) <= not((layer1_outputs(3032)) xor (layer1_outputs(449)));
    layer2_outputs(3348) <= not(layer1_outputs(2610)) or (layer1_outputs(4725));
    layer2_outputs(3349) <= not(layer1_outputs(2084)) or (layer1_outputs(5113));
    layer2_outputs(3350) <= (layer1_outputs(4801)) and not (layer1_outputs(4382));
    layer2_outputs(3351) <= not(layer1_outputs(1406));
    layer2_outputs(3352) <= not(layer1_outputs(1476));
    layer2_outputs(3353) <= not(layer1_outputs(2910)) or (layer1_outputs(3514));
    layer2_outputs(3354) <= (layer1_outputs(3008)) and (layer1_outputs(1698));
    layer2_outputs(3355) <= not(layer1_outputs(1415)) or (layer1_outputs(4289));
    layer2_outputs(3356) <= '1';
    layer2_outputs(3357) <= '1';
    layer2_outputs(3358) <= (layer1_outputs(1883)) and not (layer1_outputs(2281));
    layer2_outputs(3359) <= layer1_outputs(4315);
    layer2_outputs(3360) <= (layer1_outputs(866)) or (layer1_outputs(1386));
    layer2_outputs(3361) <= '1';
    layer2_outputs(3362) <= not((layer1_outputs(2534)) xor (layer1_outputs(3783)));
    layer2_outputs(3363) <= layer1_outputs(4211);
    layer2_outputs(3364) <= (layer1_outputs(314)) and not (layer1_outputs(4276));
    layer2_outputs(3365) <= not(layer1_outputs(1371));
    layer2_outputs(3366) <= '1';
    layer2_outputs(3367) <= '1';
    layer2_outputs(3368) <= (layer1_outputs(1348)) or (layer1_outputs(3024));
    layer2_outputs(3369) <= '1';
    layer2_outputs(3370) <= '0';
    layer2_outputs(3371) <= layer1_outputs(5039);
    layer2_outputs(3372) <= '0';
    layer2_outputs(3373) <= layer1_outputs(4463);
    layer2_outputs(3374) <= '0';
    layer2_outputs(3375) <= not(layer1_outputs(357));
    layer2_outputs(3376) <= not(layer1_outputs(2751));
    layer2_outputs(3377) <= not((layer1_outputs(3186)) or (layer1_outputs(100)));
    layer2_outputs(3378) <= (layer1_outputs(38)) and not (layer1_outputs(4735));
    layer2_outputs(3379) <= (layer1_outputs(4597)) and not (layer1_outputs(4263));
    layer2_outputs(3380) <= (layer1_outputs(525)) and not (layer1_outputs(2836));
    layer2_outputs(3381) <= '1';
    layer2_outputs(3382) <= layer1_outputs(750);
    layer2_outputs(3383) <= not((layer1_outputs(3957)) and (layer1_outputs(2135)));
    layer2_outputs(3384) <= not(layer1_outputs(4627)) or (layer1_outputs(334));
    layer2_outputs(3385) <= '1';
    layer2_outputs(3386) <= (layer1_outputs(2385)) and not (layer1_outputs(116));
    layer2_outputs(3387) <= not((layer1_outputs(1899)) or (layer1_outputs(3307)));
    layer2_outputs(3388) <= not(layer1_outputs(3636)) or (layer1_outputs(3228));
    layer2_outputs(3389) <= (layer1_outputs(4088)) xor (layer1_outputs(2319));
    layer2_outputs(3390) <= '0';
    layer2_outputs(3391) <= not(layer1_outputs(4341)) or (layer1_outputs(4230));
    layer2_outputs(3392) <= (layer1_outputs(4588)) and (layer1_outputs(1282));
    layer2_outputs(3393) <= not(layer1_outputs(4454)) or (layer1_outputs(3842));
    layer2_outputs(3394) <= not(layer1_outputs(654)) or (layer1_outputs(3973));
    layer2_outputs(3395) <= not((layer1_outputs(436)) and (layer1_outputs(2585)));
    layer2_outputs(3396) <= '0';
    layer2_outputs(3397) <= (layer1_outputs(1669)) and not (layer1_outputs(802));
    layer2_outputs(3398) <= '0';
    layer2_outputs(3399) <= '0';
    layer2_outputs(3400) <= not(layer1_outputs(3424)) or (layer1_outputs(2601));
    layer2_outputs(3401) <= '0';
    layer2_outputs(3402) <= not(layer1_outputs(3299)) or (layer1_outputs(4455));
    layer2_outputs(3403) <= (layer1_outputs(3265)) or (layer1_outputs(3351));
    layer2_outputs(3404) <= (layer1_outputs(4298)) and not (layer1_outputs(1463));
    layer2_outputs(3405) <= (layer1_outputs(4335)) xor (layer1_outputs(1446));
    layer2_outputs(3406) <= not((layer1_outputs(1552)) or (layer1_outputs(2510)));
    layer2_outputs(3407) <= (layer1_outputs(2025)) and not (layer1_outputs(4184));
    layer2_outputs(3408) <= not(layer1_outputs(1122)) or (layer1_outputs(2299));
    layer2_outputs(3409) <= '0';
    layer2_outputs(3410) <= '1';
    layer2_outputs(3411) <= '0';
    layer2_outputs(3412) <= (layer1_outputs(4899)) and not (layer1_outputs(3101));
    layer2_outputs(3413) <= '0';
    layer2_outputs(3414) <= not(layer1_outputs(3524));
    layer2_outputs(3415) <= (layer1_outputs(1820)) or (layer1_outputs(2931));
    layer2_outputs(3416) <= (layer1_outputs(451)) or (layer1_outputs(1427));
    layer2_outputs(3417) <= '1';
    layer2_outputs(3418) <= '1';
    layer2_outputs(3419) <= not(layer1_outputs(4859));
    layer2_outputs(3420) <= not(layer1_outputs(2154)) or (layer1_outputs(2346));
    layer2_outputs(3421) <= '1';
    layer2_outputs(3422) <= not(layer1_outputs(4090)) or (layer1_outputs(1843));
    layer2_outputs(3423) <= not((layer1_outputs(3317)) or (layer1_outputs(673)));
    layer2_outputs(3424) <= '1';
    layer2_outputs(3425) <= (layer1_outputs(721)) and not (layer1_outputs(2683));
    layer2_outputs(3426) <= (layer1_outputs(4279)) and not (layer1_outputs(2440));
    layer2_outputs(3427) <= not(layer1_outputs(784)) or (layer1_outputs(1191));
    layer2_outputs(3428) <= not((layer1_outputs(3137)) or (layer1_outputs(3587)));
    layer2_outputs(3429) <= (layer1_outputs(5045)) or (layer1_outputs(1641));
    layer2_outputs(3430) <= not(layer1_outputs(3399));
    layer2_outputs(3431) <= '0';
    layer2_outputs(3432) <= layer1_outputs(3974);
    layer2_outputs(3433) <= not((layer1_outputs(2067)) and (layer1_outputs(3756)));
    layer2_outputs(3434) <= (layer1_outputs(3042)) and not (layer1_outputs(2458));
    layer2_outputs(3435) <= '0';
    layer2_outputs(3436) <= not((layer1_outputs(1132)) or (layer1_outputs(1781)));
    layer2_outputs(3437) <= (layer1_outputs(3261)) and (layer1_outputs(1801));
    layer2_outputs(3438) <= not(layer1_outputs(4215)) or (layer1_outputs(732));
    layer2_outputs(3439) <= (layer1_outputs(3714)) and not (layer1_outputs(1580));
    layer2_outputs(3440) <= not(layer1_outputs(4956));
    layer2_outputs(3441) <= layer1_outputs(1072);
    layer2_outputs(3442) <= '0';
    layer2_outputs(3443) <= '1';
    layer2_outputs(3444) <= '1';
    layer2_outputs(3445) <= not(layer1_outputs(3744)) or (layer1_outputs(3182));
    layer2_outputs(3446) <= (layer1_outputs(2177)) and (layer1_outputs(3336));
    layer2_outputs(3447) <= not(layer1_outputs(3419)) or (layer1_outputs(55));
    layer2_outputs(3448) <= '1';
    layer2_outputs(3449) <= (layer1_outputs(425)) and not (layer1_outputs(667));
    layer2_outputs(3450) <= (layer1_outputs(2121)) and not (layer1_outputs(3415));
    layer2_outputs(3451) <= not((layer1_outputs(2311)) and (layer1_outputs(4948)));
    layer2_outputs(3452) <= (layer1_outputs(4598)) or (layer1_outputs(3940));
    layer2_outputs(3453) <= (layer1_outputs(1699)) or (layer1_outputs(4618));
    layer2_outputs(3454) <= not((layer1_outputs(655)) and (layer1_outputs(2924)));
    layer2_outputs(3455) <= layer1_outputs(752);
    layer2_outputs(3456) <= (layer1_outputs(2524)) and not (layer1_outputs(1813));
    layer2_outputs(3457) <= not(layer1_outputs(1536));
    layer2_outputs(3458) <= not((layer1_outputs(4874)) or (layer1_outputs(5112)));
    layer2_outputs(3459) <= (layer1_outputs(4)) xor (layer1_outputs(4594));
    layer2_outputs(3460) <= (layer1_outputs(3809)) xor (layer1_outputs(4304));
    layer2_outputs(3461) <= not(layer1_outputs(64));
    layer2_outputs(3462) <= not(layer1_outputs(4581));
    layer2_outputs(3463) <= '0';
    layer2_outputs(3464) <= not((layer1_outputs(1461)) or (layer1_outputs(2858)));
    layer2_outputs(3465) <= not(layer1_outputs(346)) or (layer1_outputs(1406));
    layer2_outputs(3466) <= layer1_outputs(729);
    layer2_outputs(3467) <= not((layer1_outputs(4711)) xor (layer1_outputs(5023)));
    layer2_outputs(3468) <= not(layer1_outputs(70)) or (layer1_outputs(1061));
    layer2_outputs(3469) <= not((layer1_outputs(1115)) and (layer1_outputs(3274)));
    layer2_outputs(3470) <= (layer1_outputs(2535)) or (layer1_outputs(2157));
    layer2_outputs(3471) <= layer1_outputs(147);
    layer2_outputs(3472) <= not((layer1_outputs(387)) or (layer1_outputs(2657)));
    layer2_outputs(3473) <= not(layer1_outputs(4386)) or (layer1_outputs(305));
    layer2_outputs(3474) <= (layer1_outputs(1069)) or (layer1_outputs(3208));
    layer2_outputs(3475) <= not(layer1_outputs(1118));
    layer2_outputs(3476) <= '0';
    layer2_outputs(3477) <= (layer1_outputs(4453)) or (layer1_outputs(58));
    layer2_outputs(3478) <= not((layer1_outputs(4893)) or (layer1_outputs(1772)));
    layer2_outputs(3479) <= (layer1_outputs(1850)) and not (layer1_outputs(4727));
    layer2_outputs(3480) <= not(layer1_outputs(2713)) or (layer1_outputs(589));
    layer2_outputs(3481) <= '1';
    layer2_outputs(3482) <= '1';
    layer2_outputs(3483) <= not((layer1_outputs(4699)) and (layer1_outputs(3256)));
    layer2_outputs(3484) <= not((layer1_outputs(3663)) and (layer1_outputs(870)));
    layer2_outputs(3485) <= not(layer1_outputs(2465));
    layer2_outputs(3486) <= (layer1_outputs(2197)) and (layer1_outputs(419));
    layer2_outputs(3487) <= layer1_outputs(1901);
    layer2_outputs(3488) <= not(layer1_outputs(3948)) or (layer1_outputs(2703));
    layer2_outputs(3489) <= (layer1_outputs(1466)) and not (layer1_outputs(3821));
    layer2_outputs(3490) <= not(layer1_outputs(2235)) or (layer1_outputs(2769));
    layer2_outputs(3491) <= not(layer1_outputs(1779));
    layer2_outputs(3492) <= (layer1_outputs(625)) xor (layer1_outputs(466));
    layer2_outputs(3493) <= (layer1_outputs(2508)) and not (layer1_outputs(3474));
    layer2_outputs(3494) <= (layer1_outputs(3244)) and not (layer1_outputs(268));
    layer2_outputs(3495) <= not(layer1_outputs(2797)) or (layer1_outputs(3577));
    layer2_outputs(3496) <= (layer1_outputs(3320)) or (layer1_outputs(3125));
    layer2_outputs(3497) <= not(layer1_outputs(2134)) or (layer1_outputs(1059));
    layer2_outputs(3498) <= (layer1_outputs(3809)) or (layer1_outputs(977));
    layer2_outputs(3499) <= '0';
    layer2_outputs(3500) <= not(layer1_outputs(2251));
    layer2_outputs(3501) <= not(layer1_outputs(3562)) or (layer1_outputs(2115));
    layer2_outputs(3502) <= not((layer1_outputs(282)) or (layer1_outputs(4835)));
    layer2_outputs(3503) <= not((layer1_outputs(1660)) and (layer1_outputs(1296)));
    layer2_outputs(3504) <= '1';
    layer2_outputs(3505) <= (layer1_outputs(4049)) and not (layer1_outputs(1320));
    layer2_outputs(3506) <= not(layer1_outputs(389)) or (layer1_outputs(3253));
    layer2_outputs(3507) <= (layer1_outputs(2822)) or (layer1_outputs(2520));
    layer2_outputs(3508) <= (layer1_outputs(1070)) or (layer1_outputs(2622));
    layer2_outputs(3509) <= (layer1_outputs(2330)) or (layer1_outputs(1641));
    layer2_outputs(3510) <= not(layer1_outputs(857));
    layer2_outputs(3511) <= not(layer1_outputs(1743));
    layer2_outputs(3512) <= '1';
    layer2_outputs(3513) <= '1';
    layer2_outputs(3514) <= not(layer1_outputs(4071)) or (layer1_outputs(1793));
    layer2_outputs(3515) <= '0';
    layer2_outputs(3516) <= '0';
    layer2_outputs(3517) <= not(layer1_outputs(3602)) or (layer1_outputs(3533));
    layer2_outputs(3518) <= not((layer1_outputs(1457)) or (layer1_outputs(2605)));
    layer2_outputs(3519) <= (layer1_outputs(669)) or (layer1_outputs(1019));
    layer2_outputs(3520) <= not(layer1_outputs(1173));
    layer2_outputs(3521) <= (layer1_outputs(3702)) and (layer1_outputs(275));
    layer2_outputs(3522) <= not((layer1_outputs(309)) and (layer1_outputs(4895)));
    layer2_outputs(3523) <= '0';
    layer2_outputs(3524) <= not((layer1_outputs(4924)) or (layer1_outputs(4673)));
    layer2_outputs(3525) <= (layer1_outputs(2847)) and not (layer1_outputs(4355));
    layer2_outputs(3526) <= '0';
    layer2_outputs(3527) <= '1';
    layer2_outputs(3528) <= (layer1_outputs(2270)) and not (layer1_outputs(644));
    layer2_outputs(3529) <= not((layer1_outputs(2374)) and (layer1_outputs(951)));
    layer2_outputs(3530) <= not(layer1_outputs(2186));
    layer2_outputs(3531) <= '0';
    layer2_outputs(3532) <= layer1_outputs(733);
    layer2_outputs(3533) <= (layer1_outputs(668)) and (layer1_outputs(3708));
    layer2_outputs(3534) <= layer1_outputs(2921);
    layer2_outputs(3535) <= not((layer1_outputs(665)) and (layer1_outputs(1970)));
    layer2_outputs(3536) <= '1';
    layer2_outputs(3537) <= not((layer1_outputs(949)) and (layer1_outputs(195)));
    layer2_outputs(3538) <= (layer1_outputs(48)) and not (layer1_outputs(659));
    layer2_outputs(3539) <= (layer1_outputs(1919)) and (layer1_outputs(633));
    layer2_outputs(3540) <= (layer1_outputs(2829)) or (layer1_outputs(873));
    layer2_outputs(3541) <= '1';
    layer2_outputs(3542) <= not(layer1_outputs(2143)) or (layer1_outputs(3393));
    layer2_outputs(3543) <= not(layer1_outputs(2532)) or (layer1_outputs(1694));
    layer2_outputs(3544) <= not(layer1_outputs(2395));
    layer2_outputs(3545) <= not((layer1_outputs(4224)) or (layer1_outputs(3406)));
    layer2_outputs(3546) <= not(layer1_outputs(1426)) or (layer1_outputs(1476));
    layer2_outputs(3547) <= not((layer1_outputs(327)) and (layer1_outputs(4246)));
    layer2_outputs(3548) <= (layer1_outputs(886)) and (layer1_outputs(4704));
    layer2_outputs(3549) <= not(layer1_outputs(707));
    layer2_outputs(3550) <= '0';
    layer2_outputs(3551) <= (layer1_outputs(3622)) xor (layer1_outputs(1924));
    layer2_outputs(3552) <= (layer1_outputs(786)) xor (layer1_outputs(2194));
    layer2_outputs(3553) <= not(layer1_outputs(867)) or (layer1_outputs(3133));
    layer2_outputs(3554) <= (layer1_outputs(2969)) or (layer1_outputs(859));
    layer2_outputs(3555) <= (layer1_outputs(3633)) and (layer1_outputs(2422));
    layer2_outputs(3556) <= not((layer1_outputs(4566)) or (layer1_outputs(82)));
    layer2_outputs(3557) <= '0';
    layer2_outputs(3558) <= '0';
    layer2_outputs(3559) <= '1';
    layer2_outputs(3560) <= layer1_outputs(1854);
    layer2_outputs(3561) <= not(layer1_outputs(3372)) or (layer1_outputs(1008));
    layer2_outputs(3562) <= '1';
    layer2_outputs(3563) <= not(layer1_outputs(360)) or (layer1_outputs(4468));
    layer2_outputs(3564) <= not(layer1_outputs(1192)) or (layer1_outputs(636));
    layer2_outputs(3565) <= (layer1_outputs(1439)) or (layer1_outputs(4220));
    layer2_outputs(3566) <= '0';
    layer2_outputs(3567) <= not(layer1_outputs(652));
    layer2_outputs(3568) <= not(layer1_outputs(12));
    layer2_outputs(3569) <= '1';
    layer2_outputs(3570) <= (layer1_outputs(3272)) and not (layer1_outputs(1663));
    layer2_outputs(3571) <= not(layer1_outputs(4570));
    layer2_outputs(3572) <= (layer1_outputs(2800)) xor (layer1_outputs(2259));
    layer2_outputs(3573) <= not((layer1_outputs(1796)) and (layer1_outputs(3311)));
    layer2_outputs(3574) <= '1';
    layer2_outputs(3575) <= (layer1_outputs(219)) and not (layer1_outputs(1274));
    layer2_outputs(3576) <= (layer1_outputs(2842)) and (layer1_outputs(1169));
    layer2_outputs(3577) <= not(layer1_outputs(1985));
    layer2_outputs(3578) <= not(layer1_outputs(3516)) or (layer1_outputs(4574));
    layer2_outputs(3579) <= not((layer1_outputs(3182)) or (layer1_outputs(1652)));
    layer2_outputs(3580) <= not(layer1_outputs(2331));
    layer2_outputs(3581) <= not((layer1_outputs(4497)) and (layer1_outputs(2956)));
    layer2_outputs(3582) <= not(layer1_outputs(215)) or (layer1_outputs(5002));
    layer2_outputs(3583) <= layer1_outputs(1708);
    layer2_outputs(3584) <= layer1_outputs(1120);
    layer2_outputs(3585) <= (layer1_outputs(2948)) and not (layer1_outputs(3818));
    layer2_outputs(3586) <= '1';
    layer2_outputs(3587) <= (layer1_outputs(660)) and (layer1_outputs(2491));
    layer2_outputs(3588) <= '0';
    layer2_outputs(3589) <= not((layer1_outputs(2738)) or (layer1_outputs(2894)));
    layer2_outputs(3590) <= (layer1_outputs(438)) and not (layer1_outputs(1664));
    layer2_outputs(3591) <= '1';
    layer2_outputs(3592) <= '1';
    layer2_outputs(3593) <= not((layer1_outputs(399)) and (layer1_outputs(249)));
    layer2_outputs(3594) <= not(layer1_outputs(3927)) or (layer1_outputs(4633));
    layer2_outputs(3595) <= (layer1_outputs(3722)) and (layer1_outputs(1145));
    layer2_outputs(3596) <= layer1_outputs(4763);
    layer2_outputs(3597) <= layer1_outputs(4641);
    layer2_outputs(3598) <= '1';
    layer2_outputs(3599) <= '0';
    layer2_outputs(3600) <= '1';
    layer2_outputs(3601) <= layer1_outputs(2752);
    layer2_outputs(3602) <= not(layer1_outputs(4582));
    layer2_outputs(3603) <= not(layer1_outputs(4691)) or (layer1_outputs(4743));
    layer2_outputs(3604) <= layer1_outputs(4905);
    layer2_outputs(3605) <= (layer1_outputs(209)) and not (layer1_outputs(2594));
    layer2_outputs(3606) <= not(layer1_outputs(4368));
    layer2_outputs(3607) <= (layer1_outputs(1854)) and not (layer1_outputs(4608));
    layer2_outputs(3608) <= not(layer1_outputs(2874)) or (layer1_outputs(2966));
    layer2_outputs(3609) <= not(layer1_outputs(3170));
    layer2_outputs(3610) <= not(layer1_outputs(3524)) or (layer1_outputs(3694));
    layer2_outputs(3611) <= layer1_outputs(278);
    layer2_outputs(3612) <= not(layer1_outputs(977));
    layer2_outputs(3613) <= '1';
    layer2_outputs(3614) <= '1';
    layer2_outputs(3615) <= not(layer1_outputs(3752));
    layer2_outputs(3616) <= (layer1_outputs(1796)) and not (layer1_outputs(5030));
    layer2_outputs(3617) <= layer1_outputs(4680);
    layer2_outputs(3618) <= '1';
    layer2_outputs(3619) <= '1';
    layer2_outputs(3620) <= (layer1_outputs(4959)) and not (layer1_outputs(731));
    layer2_outputs(3621) <= not((layer1_outputs(4168)) and (layer1_outputs(4940)));
    layer2_outputs(3622) <= (layer1_outputs(1260)) and (layer1_outputs(1626));
    layer2_outputs(3623) <= '1';
    layer2_outputs(3624) <= (layer1_outputs(383)) and not (layer1_outputs(3758));
    layer2_outputs(3625) <= layer1_outputs(4060);
    layer2_outputs(3626) <= (layer1_outputs(2810)) and (layer1_outputs(1573));
    layer2_outputs(3627) <= '0';
    layer2_outputs(3628) <= layer1_outputs(3083);
    layer2_outputs(3629) <= not(layer1_outputs(2198)) or (layer1_outputs(4355));
    layer2_outputs(3630) <= layer1_outputs(4886);
    layer2_outputs(3631) <= not(layer1_outputs(4794)) or (layer1_outputs(54));
    layer2_outputs(3632) <= not(layer1_outputs(3874));
    layer2_outputs(3633) <= not((layer1_outputs(609)) or (layer1_outputs(2860)));
    layer2_outputs(3634) <= not(layer1_outputs(2406));
    layer2_outputs(3635) <= not((layer1_outputs(2551)) and (layer1_outputs(4731)));
    layer2_outputs(3636) <= layer1_outputs(2808);
    layer2_outputs(3637) <= layer1_outputs(5033);
    layer2_outputs(3638) <= '1';
    layer2_outputs(3639) <= (layer1_outputs(2201)) or (layer1_outputs(3812));
    layer2_outputs(3640) <= (layer1_outputs(1171)) and not (layer1_outputs(2941));
    layer2_outputs(3641) <= (layer1_outputs(2487)) or (layer1_outputs(818));
    layer2_outputs(3642) <= (layer1_outputs(1762)) and not (layer1_outputs(5087));
    layer2_outputs(3643) <= not(layer1_outputs(1637));
    layer2_outputs(3644) <= not(layer1_outputs(608)) or (layer1_outputs(3760));
    layer2_outputs(3645) <= not((layer1_outputs(4360)) or (layer1_outputs(3857)));
    layer2_outputs(3646) <= '1';
    layer2_outputs(3647) <= '1';
    layer2_outputs(3648) <= (layer1_outputs(700)) and not (layer1_outputs(2361));
    layer2_outputs(3649) <= '1';
    layer2_outputs(3650) <= not((layer1_outputs(3519)) and (layer1_outputs(4490)));
    layer2_outputs(3651) <= not((layer1_outputs(990)) and (layer1_outputs(1044)));
    layer2_outputs(3652) <= not((layer1_outputs(814)) or (layer1_outputs(4391)));
    layer2_outputs(3653) <= not((layer1_outputs(3548)) and (layer1_outputs(2610)));
    layer2_outputs(3654) <= not((layer1_outputs(695)) or (layer1_outputs(4541)));
    layer2_outputs(3655) <= layer1_outputs(2495);
    layer2_outputs(3656) <= not(layer1_outputs(4987));
    layer2_outputs(3657) <= not(layer1_outputs(3817)) or (layer1_outputs(4372));
    layer2_outputs(3658) <= not((layer1_outputs(4729)) or (layer1_outputs(154)));
    layer2_outputs(3659) <= '1';
    layer2_outputs(3660) <= (layer1_outputs(3673)) or (layer1_outputs(2692));
    layer2_outputs(3661) <= (layer1_outputs(4179)) and (layer1_outputs(3287));
    layer2_outputs(3662) <= not(layer1_outputs(2722)) or (layer1_outputs(1986));
    layer2_outputs(3663) <= '0';
    layer2_outputs(3664) <= '1';
    layer2_outputs(3665) <= not((layer1_outputs(500)) xor (layer1_outputs(1110)));
    layer2_outputs(3666) <= not((layer1_outputs(4541)) and (layer1_outputs(2737)));
    layer2_outputs(3667) <= not(layer1_outputs(1638)) or (layer1_outputs(2932));
    layer2_outputs(3668) <= not((layer1_outputs(1526)) or (layer1_outputs(2714)));
    layer2_outputs(3669) <= not((layer1_outputs(1981)) and (layer1_outputs(2041)));
    layer2_outputs(3670) <= (layer1_outputs(3733)) or (layer1_outputs(1996));
    layer2_outputs(3671) <= layer1_outputs(1575);
    layer2_outputs(3672) <= not(layer1_outputs(4865));
    layer2_outputs(3673) <= (layer1_outputs(728)) and not (layer1_outputs(1525));
    layer2_outputs(3674) <= '1';
    layer2_outputs(3675) <= '1';
    layer2_outputs(3676) <= (layer1_outputs(1511)) xor (layer1_outputs(1139));
    layer2_outputs(3677) <= '0';
    layer2_outputs(3678) <= not((layer1_outputs(2634)) or (layer1_outputs(2303)));
    layer2_outputs(3679) <= not(layer1_outputs(566));
    layer2_outputs(3680) <= (layer1_outputs(2833)) or (layer1_outputs(2092));
    layer2_outputs(3681) <= not(layer1_outputs(2763));
    layer2_outputs(3682) <= not(layer1_outputs(273));
    layer2_outputs(3683) <= (layer1_outputs(2105)) and not (layer1_outputs(4361));
    layer2_outputs(3684) <= layer1_outputs(3724);
    layer2_outputs(3685) <= layer1_outputs(4534);
    layer2_outputs(3686) <= layer1_outputs(3263);
    layer2_outputs(3687) <= (layer1_outputs(1151)) and not (layer1_outputs(1722));
    layer2_outputs(3688) <= not(layer1_outputs(3559)) or (layer1_outputs(4237));
    layer2_outputs(3689) <= layer1_outputs(2008);
    layer2_outputs(3690) <= not(layer1_outputs(1310)) or (layer1_outputs(3522));
    layer2_outputs(3691) <= '1';
    layer2_outputs(3692) <= (layer1_outputs(2799)) and not (layer1_outputs(4307));
    layer2_outputs(3693) <= not((layer1_outputs(3825)) and (layer1_outputs(4985)));
    layer2_outputs(3694) <= '0';
    layer2_outputs(3695) <= (layer1_outputs(50)) or (layer1_outputs(3063));
    layer2_outputs(3696) <= '0';
    layer2_outputs(3697) <= (layer1_outputs(1042)) and not (layer1_outputs(3607));
    layer2_outputs(3698) <= layer1_outputs(366);
    layer2_outputs(3699) <= not(layer1_outputs(114)) or (layer1_outputs(1904));
    layer2_outputs(3700) <= '1';
    layer2_outputs(3701) <= not(layer1_outputs(3720)) or (layer1_outputs(4774));
    layer2_outputs(3702) <= layer1_outputs(1216);
    layer2_outputs(3703) <= '1';
    layer2_outputs(3704) <= (layer1_outputs(1926)) and (layer1_outputs(3629));
    layer2_outputs(3705) <= not(layer1_outputs(1009)) or (layer1_outputs(1495));
    layer2_outputs(3706) <= '0';
    layer2_outputs(3707) <= not(layer1_outputs(4760));
    layer2_outputs(3708) <= '1';
    layer2_outputs(3709) <= layer1_outputs(1759);
    layer2_outputs(3710) <= (layer1_outputs(1334)) or (layer1_outputs(5020));
    layer2_outputs(3711) <= '1';
    layer2_outputs(3712) <= '0';
    layer2_outputs(3713) <= '0';
    layer2_outputs(3714) <= (layer1_outputs(1598)) and not (layer1_outputs(2617));
    layer2_outputs(3715) <= (layer1_outputs(684)) and (layer1_outputs(4595));
    layer2_outputs(3716) <= not(layer1_outputs(3763)) or (layer1_outputs(3726));
    layer2_outputs(3717) <= not((layer1_outputs(2438)) or (layer1_outputs(3583)));
    layer2_outputs(3718) <= not(layer1_outputs(632)) or (layer1_outputs(2232));
    layer2_outputs(3719) <= layer1_outputs(1091);
    layer2_outputs(3720) <= not(layer1_outputs(4862));
    layer2_outputs(3721) <= layer1_outputs(3625);
    layer2_outputs(3722) <= '1';
    layer2_outputs(3723) <= not(layer1_outputs(3393)) or (layer1_outputs(4395));
    layer2_outputs(3724) <= '1';
    layer2_outputs(3725) <= not(layer1_outputs(4460)) or (layer1_outputs(2098));
    layer2_outputs(3726) <= (layer1_outputs(5024)) or (layer1_outputs(4491));
    layer2_outputs(3727) <= layer1_outputs(587);
    layer2_outputs(3728) <= (layer1_outputs(89)) and not (layer1_outputs(1866));
    layer2_outputs(3729) <= not(layer1_outputs(4620));
    layer2_outputs(3730) <= (layer1_outputs(4042)) and not (layer1_outputs(2474));
    layer2_outputs(3731) <= not((layer1_outputs(2036)) or (layer1_outputs(4695)));
    layer2_outputs(3732) <= '0';
    layer2_outputs(3733) <= layer1_outputs(4861);
    layer2_outputs(3734) <= '1';
    layer2_outputs(3735) <= not(layer1_outputs(4697));
    layer2_outputs(3736) <= '1';
    layer2_outputs(3737) <= not(layer1_outputs(57));
    layer2_outputs(3738) <= not(layer1_outputs(1947));
    layer2_outputs(3739) <= '0';
    layer2_outputs(3740) <= (layer1_outputs(4359)) xor (layer1_outputs(1695));
    layer2_outputs(3741) <= '0';
    layer2_outputs(3742) <= '1';
    layer2_outputs(3743) <= not(layer1_outputs(403));
    layer2_outputs(3744) <= '1';
    layer2_outputs(3745) <= not((layer1_outputs(639)) or (layer1_outputs(3628)));
    layer2_outputs(3746) <= '0';
    layer2_outputs(3747) <= not((layer1_outputs(495)) or (layer1_outputs(3078)));
    layer2_outputs(3748) <= not((layer1_outputs(1180)) or (layer1_outputs(4277)));
    layer2_outputs(3749) <= (layer1_outputs(1582)) and (layer1_outputs(1421));
    layer2_outputs(3750) <= '1';
    layer2_outputs(3751) <= layer1_outputs(694);
    layer2_outputs(3752) <= not(layer1_outputs(1748));
    layer2_outputs(3753) <= not(layer1_outputs(4874));
    layer2_outputs(3754) <= not(layer1_outputs(429));
    layer2_outputs(3755) <= layer1_outputs(3747);
    layer2_outputs(3756) <= '0';
    layer2_outputs(3757) <= (layer1_outputs(3578)) and (layer1_outputs(4649));
    layer2_outputs(3758) <= '0';
    layer2_outputs(3759) <= layer1_outputs(803);
    layer2_outputs(3760) <= not(layer1_outputs(4109));
    layer2_outputs(3761) <= not((layer1_outputs(3315)) or (layer1_outputs(3581)));
    layer2_outputs(3762) <= not((layer1_outputs(4475)) or (layer1_outputs(773)));
    layer2_outputs(3763) <= (layer1_outputs(37)) and (layer1_outputs(2432));
    layer2_outputs(3764) <= (layer1_outputs(4602)) or (layer1_outputs(4576));
    layer2_outputs(3765) <= not(layer1_outputs(3283)) or (layer1_outputs(1374));
    layer2_outputs(3766) <= not(layer1_outputs(2990)) or (layer1_outputs(2780));
    layer2_outputs(3767) <= layer1_outputs(3022);
    layer2_outputs(3768) <= (layer1_outputs(4323)) and not (layer1_outputs(68));
    layer2_outputs(3769) <= (layer1_outputs(3057)) and not (layer1_outputs(4415));
    layer2_outputs(3770) <= '0';
    layer2_outputs(3771) <= layer1_outputs(2828);
    layer2_outputs(3772) <= (layer1_outputs(2016)) and not (layer1_outputs(3785));
    layer2_outputs(3773) <= (layer1_outputs(632)) or (layer1_outputs(2928));
    layer2_outputs(3774) <= layer1_outputs(2120);
    layer2_outputs(3775) <= '1';
    layer2_outputs(3776) <= (layer1_outputs(1278)) and not (layer1_outputs(1719));
    layer2_outputs(3777) <= (layer1_outputs(3862)) xor (layer1_outputs(4150));
    layer2_outputs(3778) <= not(layer1_outputs(3276)) or (layer1_outputs(1325));
    layer2_outputs(3779) <= (layer1_outputs(4289)) or (layer1_outputs(4043));
    layer2_outputs(3780) <= (layer1_outputs(749)) and (layer1_outputs(2015));
    layer2_outputs(3781) <= (layer1_outputs(2599)) and (layer1_outputs(3254));
    layer2_outputs(3782) <= (layer1_outputs(4031)) or (layer1_outputs(5073));
    layer2_outputs(3783) <= '0';
    layer2_outputs(3784) <= layer1_outputs(2488);
    layer2_outputs(3785) <= not((layer1_outputs(2480)) and (layer1_outputs(5064)));
    layer2_outputs(3786) <= not(layer1_outputs(2832));
    layer2_outputs(3787) <= not(layer1_outputs(4302)) or (layer1_outputs(3039));
    layer2_outputs(3788) <= (layer1_outputs(961)) and not (layer1_outputs(609));
    layer2_outputs(3789) <= (layer1_outputs(2649)) and not (layer1_outputs(128));
    layer2_outputs(3790) <= not((layer1_outputs(1844)) or (layer1_outputs(1490)));
    layer2_outputs(3791) <= not(layer1_outputs(31));
    layer2_outputs(3792) <= layer1_outputs(1928);
    layer2_outputs(3793) <= (layer1_outputs(3665)) or (layer1_outputs(1747));
    layer2_outputs(3794) <= '1';
    layer2_outputs(3795) <= not(layer1_outputs(307)) or (layer1_outputs(2645));
    layer2_outputs(3796) <= '0';
    layer2_outputs(3797) <= '0';
    layer2_outputs(3798) <= '1';
    layer2_outputs(3799) <= '1';
    layer2_outputs(3800) <= (layer1_outputs(4284)) and (layer1_outputs(2994));
    layer2_outputs(3801) <= (layer1_outputs(1961)) and not (layer1_outputs(4623));
    layer2_outputs(3802) <= not(layer1_outputs(927)) or (layer1_outputs(3421));
    layer2_outputs(3803) <= not(layer1_outputs(2153)) or (layer1_outputs(3020));
    layer2_outputs(3804) <= not(layer1_outputs(423));
    layer2_outputs(3805) <= (layer1_outputs(1864)) and not (layer1_outputs(1633));
    layer2_outputs(3806) <= (layer1_outputs(934)) and not (layer1_outputs(151));
    layer2_outputs(3807) <= layer1_outputs(3828);
    layer2_outputs(3808) <= (layer1_outputs(3858)) and not (layer1_outputs(5069));
    layer2_outputs(3809) <= not((layer1_outputs(4097)) or (layer1_outputs(1020)));
    layer2_outputs(3810) <= (layer1_outputs(920)) or (layer1_outputs(936));
    layer2_outputs(3811) <= '0';
    layer2_outputs(3812) <= not(layer1_outputs(4241));
    layer2_outputs(3813) <= (layer1_outputs(1839)) and not (layer1_outputs(1845));
    layer2_outputs(3814) <= not(layer1_outputs(2414));
    layer2_outputs(3815) <= not((layer1_outputs(2058)) and (layer1_outputs(1189)));
    layer2_outputs(3816) <= '0';
    layer2_outputs(3817) <= not((layer1_outputs(303)) and (layer1_outputs(3517)));
    layer2_outputs(3818) <= not(layer1_outputs(965));
    layer2_outputs(3819) <= (layer1_outputs(3262)) and (layer1_outputs(28));
    layer2_outputs(3820) <= '0';
    layer2_outputs(3821) <= not(layer1_outputs(1366)) or (layer1_outputs(3271));
    layer2_outputs(3822) <= '1';
    layer2_outputs(3823) <= not(layer1_outputs(1363));
    layer2_outputs(3824) <= (layer1_outputs(3181)) and not (layer1_outputs(499));
    layer2_outputs(3825) <= not(layer1_outputs(556)) or (layer1_outputs(260));
    layer2_outputs(3826) <= '1';
    layer2_outputs(3827) <= not(layer1_outputs(4817)) or (layer1_outputs(1693));
    layer2_outputs(3828) <= not(layer1_outputs(5001));
    layer2_outputs(3829) <= not(layer1_outputs(4111)) or (layer1_outputs(5118));
    layer2_outputs(3830) <= '0';
    layer2_outputs(3831) <= not(layer1_outputs(2430));
    layer2_outputs(3832) <= not(layer1_outputs(2427));
    layer2_outputs(3833) <= not((layer1_outputs(2193)) or (layer1_outputs(4932)));
    layer2_outputs(3834) <= not(layer1_outputs(2551));
    layer2_outputs(3835) <= (layer1_outputs(4181)) and not (layer1_outputs(4356));
    layer2_outputs(3836) <= not(layer1_outputs(3363)) or (layer1_outputs(2777));
    layer2_outputs(3837) <= '1';
    layer2_outputs(3838) <= (layer1_outputs(3248)) or (layer1_outputs(3278));
    layer2_outputs(3839) <= not(layer1_outputs(3759)) or (layer1_outputs(2281));
    layer2_outputs(3840) <= (layer1_outputs(422)) and not (layer1_outputs(756));
    layer2_outputs(3841) <= (layer1_outputs(3751)) or (layer1_outputs(3552));
    layer2_outputs(3842) <= layer1_outputs(3822);
    layer2_outputs(3843) <= layer1_outputs(554);
    layer2_outputs(3844) <= not(layer1_outputs(4597)) or (layer1_outputs(4764));
    layer2_outputs(3845) <= not(layer1_outputs(947));
    layer2_outputs(3846) <= not(layer1_outputs(2600)) or (layer1_outputs(867));
    layer2_outputs(3847) <= not(layer1_outputs(1517)) or (layer1_outputs(2445));
    layer2_outputs(3848) <= '1';
    layer2_outputs(3849) <= not(layer1_outputs(212)) or (layer1_outputs(1430));
    layer2_outputs(3850) <= (layer1_outputs(3412)) or (layer1_outputs(4660));
    layer2_outputs(3851) <= layer1_outputs(3193);
    layer2_outputs(3852) <= not(layer1_outputs(4542)) or (layer1_outputs(1420));
    layer2_outputs(3853) <= not(layer1_outputs(4417));
    layer2_outputs(3854) <= (layer1_outputs(4796)) and not (layer1_outputs(4520));
    layer2_outputs(3855) <= (layer1_outputs(4211)) and (layer1_outputs(2605));
    layer2_outputs(3856) <= '1';
    layer2_outputs(3857) <= (layer1_outputs(2344)) and (layer1_outputs(4579));
    layer2_outputs(3858) <= '0';
    layer2_outputs(3859) <= (layer1_outputs(3295)) and (layer1_outputs(1649));
    layer2_outputs(3860) <= not((layer1_outputs(2963)) and (layer1_outputs(2644)));
    layer2_outputs(3861) <= (layer1_outputs(570)) and (layer1_outputs(1083));
    layer2_outputs(3862) <= not(layer1_outputs(2725)) or (layer1_outputs(2859));
    layer2_outputs(3863) <= '1';
    layer2_outputs(3864) <= '0';
    layer2_outputs(3865) <= (layer1_outputs(2175)) and not (layer1_outputs(2109));
    layer2_outputs(3866) <= (layer1_outputs(4689)) and not (layer1_outputs(2867));
    layer2_outputs(3867) <= (layer1_outputs(3169)) and not (layer1_outputs(3282));
    layer2_outputs(3868) <= '1';
    layer2_outputs(3869) <= not(layer1_outputs(1506)) or (layer1_outputs(111));
    layer2_outputs(3870) <= not((layer1_outputs(183)) or (layer1_outputs(589)));
    layer2_outputs(3871) <= not(layer1_outputs(4040)) or (layer1_outputs(1240));
    layer2_outputs(3872) <= (layer1_outputs(2111)) and not (layer1_outputs(2960));
    layer2_outputs(3873) <= not(layer1_outputs(3080));
    layer2_outputs(3874) <= not((layer1_outputs(904)) and (layer1_outputs(4956)));
    layer2_outputs(3875) <= (layer1_outputs(3138)) and (layer1_outputs(3161));
    layer2_outputs(3876) <= '0';
    layer2_outputs(3877) <= '0';
    layer2_outputs(3878) <= not(layer1_outputs(1172));
    layer2_outputs(3879) <= (layer1_outputs(3749)) and not (layer1_outputs(2439));
    layer2_outputs(3880) <= not(layer1_outputs(755));
    layer2_outputs(3881) <= layer1_outputs(1977);
    layer2_outputs(3882) <= '1';
    layer2_outputs(3883) <= not(layer1_outputs(2152));
    layer2_outputs(3884) <= not((layer1_outputs(1415)) or (layer1_outputs(8)));
    layer2_outputs(3885) <= (layer1_outputs(3912)) and (layer1_outputs(2780));
    layer2_outputs(3886) <= '0';
    layer2_outputs(3887) <= '0';
    layer2_outputs(3888) <= not((layer1_outputs(267)) and (layer1_outputs(3115)));
    layer2_outputs(3889) <= not(layer1_outputs(3631)) or (layer1_outputs(231));
    layer2_outputs(3890) <= (layer1_outputs(3625)) and (layer1_outputs(3993));
    layer2_outputs(3891) <= '0';
    layer2_outputs(3892) <= (layer1_outputs(1534)) and not (layer1_outputs(3907));
    layer2_outputs(3893) <= not(layer1_outputs(3451)) or (layer1_outputs(3224));
    layer2_outputs(3894) <= (layer1_outputs(4012)) and (layer1_outputs(5073));
    layer2_outputs(3895) <= '0';
    layer2_outputs(3896) <= '0';
    layer2_outputs(3897) <= not((layer1_outputs(704)) or (layer1_outputs(4966)));
    layer2_outputs(3898) <= (layer1_outputs(889)) or (layer1_outputs(3904));
    layer2_outputs(3899) <= not(layer1_outputs(2375));
    layer2_outputs(3900) <= not(layer1_outputs(308)) or (layer1_outputs(2429));
    layer2_outputs(3901) <= '1';
    layer2_outputs(3902) <= not(layer1_outputs(2280));
    layer2_outputs(3903) <= (layer1_outputs(491)) and not (layer1_outputs(785));
    layer2_outputs(3904) <= '0';
    layer2_outputs(3905) <= '1';
    layer2_outputs(3906) <= (layer1_outputs(4745)) and (layer1_outputs(4778));
    layer2_outputs(3907) <= not((layer1_outputs(1867)) or (layer1_outputs(4404)));
    layer2_outputs(3908) <= (layer1_outputs(1040)) and (layer1_outputs(4258));
    layer2_outputs(3909) <= not((layer1_outputs(3997)) or (layer1_outputs(1400)));
    layer2_outputs(3910) <= '0';
    layer2_outputs(3911) <= (layer1_outputs(3601)) and not (layer1_outputs(635));
    layer2_outputs(3912) <= '1';
    layer2_outputs(3913) <= '0';
    layer2_outputs(3914) <= '1';
    layer2_outputs(3915) <= (layer1_outputs(3279)) and not (layer1_outputs(2908));
    layer2_outputs(3916) <= '0';
    layer2_outputs(3917) <= not((layer1_outputs(4523)) and (layer1_outputs(4603)));
    layer2_outputs(3918) <= not(layer1_outputs(213)) or (layer1_outputs(2570));
    layer2_outputs(3919) <= (layer1_outputs(2243)) and not (layer1_outputs(4079));
    layer2_outputs(3920) <= not((layer1_outputs(960)) or (layer1_outputs(2115)));
    layer2_outputs(3921) <= not((layer1_outputs(1193)) xor (layer1_outputs(3586)));
    layer2_outputs(3922) <= not((layer1_outputs(1738)) xor (layer1_outputs(5086)));
    layer2_outputs(3923) <= layer1_outputs(1626);
    layer2_outputs(3924) <= (layer1_outputs(1220)) and (layer1_outputs(2171));
    layer2_outputs(3925) <= not((layer1_outputs(4722)) and (layer1_outputs(562)));
    layer2_outputs(3926) <= not((layer1_outputs(3445)) and (layer1_outputs(2277)));
    layer2_outputs(3927) <= layer1_outputs(4159);
    layer2_outputs(3928) <= layer1_outputs(1758);
    layer2_outputs(3929) <= '1';
    layer2_outputs(3930) <= layer1_outputs(2465);
    layer2_outputs(3931) <= '1';
    layer2_outputs(3932) <= layer1_outputs(2700);
    layer2_outputs(3933) <= not(layer1_outputs(854)) or (layer1_outputs(2319));
    layer2_outputs(3934) <= not(layer1_outputs(2798));
    layer2_outputs(3935) <= '1';
    layer2_outputs(3936) <= (layer1_outputs(4924)) and not (layer1_outputs(535));
    layer2_outputs(3937) <= not((layer1_outputs(2260)) or (layer1_outputs(4891)));
    layer2_outputs(3938) <= (layer1_outputs(3082)) and not (layer1_outputs(3244));
    layer2_outputs(3939) <= not(layer1_outputs(4822)) or (layer1_outputs(3004));
    layer2_outputs(3940) <= (layer1_outputs(2425)) and (layer1_outputs(3065));
    layer2_outputs(3941) <= '1';
    layer2_outputs(3942) <= not((layer1_outputs(1196)) or (layer1_outputs(4234)));
    layer2_outputs(3943) <= layer1_outputs(2211);
    layer2_outputs(3944) <= not(layer1_outputs(4926)) or (layer1_outputs(3354));
    layer2_outputs(3945) <= layer1_outputs(748);
    layer2_outputs(3946) <= not((layer1_outputs(2726)) and (layer1_outputs(1756)));
    layer2_outputs(3947) <= '0';
    layer2_outputs(3948) <= (layer1_outputs(2215)) and (layer1_outputs(5103));
    layer2_outputs(3949) <= not((layer1_outputs(1812)) or (layer1_outputs(3137)));
    layer2_outputs(3950) <= not((layer1_outputs(4888)) and (layer1_outputs(4165)));
    layer2_outputs(3951) <= not(layer1_outputs(1900)) or (layer1_outputs(2096));
    layer2_outputs(3952) <= '0';
    layer2_outputs(3953) <= '0';
    layer2_outputs(3954) <= not(layer1_outputs(4477)) or (layer1_outputs(2814));
    layer2_outputs(3955) <= not(layer1_outputs(798)) or (layer1_outputs(527));
    layer2_outputs(3956) <= '0';
    layer2_outputs(3957) <= layer1_outputs(3606);
    layer2_outputs(3958) <= '1';
    layer2_outputs(3959) <= (layer1_outputs(3256)) and not (layer1_outputs(1142));
    layer2_outputs(3960) <= (layer1_outputs(432)) and not (layer1_outputs(3128));
    layer2_outputs(3961) <= '1';
    layer2_outputs(3962) <= not((layer1_outputs(4025)) or (layer1_outputs(3376)));
    layer2_outputs(3963) <= (layer1_outputs(395)) and not (layer1_outputs(4564));
    layer2_outputs(3964) <= '0';
    layer2_outputs(3965) <= not(layer1_outputs(2146));
    layer2_outputs(3966) <= '0';
    layer2_outputs(3967) <= not(layer1_outputs(4896));
    layer2_outputs(3968) <= '0';
    layer2_outputs(3969) <= '0';
    layer2_outputs(3970) <= not(layer1_outputs(3836));
    layer2_outputs(3971) <= not(layer1_outputs(4467)) or (layer1_outputs(1916));
    layer2_outputs(3972) <= not(layer1_outputs(3961)) or (layer1_outputs(364));
    layer2_outputs(3973) <= layer1_outputs(4638);
    layer2_outputs(3974) <= not((layer1_outputs(1288)) or (layer1_outputs(5021)));
    layer2_outputs(3975) <= '0';
    layer2_outputs(3976) <= not(layer1_outputs(1818));
    layer2_outputs(3977) <= not((layer1_outputs(3466)) and (layer1_outputs(2340)));
    layer2_outputs(3978) <= not((layer1_outputs(3718)) or (layer1_outputs(4695)));
    layer2_outputs(3979) <= (layer1_outputs(2957)) or (layer1_outputs(3707));
    layer2_outputs(3980) <= (layer1_outputs(3435)) and not (layer1_outputs(4501));
    layer2_outputs(3981) <= (layer1_outputs(1293)) or (layer1_outputs(2283));
    layer2_outputs(3982) <= layer1_outputs(471);
    layer2_outputs(3983) <= (layer1_outputs(3370)) and not (layer1_outputs(62));
    layer2_outputs(3984) <= not((layer1_outputs(2637)) and (layer1_outputs(970)));
    layer2_outputs(3985) <= (layer1_outputs(2003)) and (layer1_outputs(2703));
    layer2_outputs(3986) <= not((layer1_outputs(3924)) and (layer1_outputs(2334)));
    layer2_outputs(3987) <= layer1_outputs(2974);
    layer2_outputs(3988) <= '1';
    layer2_outputs(3989) <= layer1_outputs(2905);
    layer2_outputs(3990) <= (layer1_outputs(2679)) or (layer1_outputs(4358));
    layer2_outputs(3991) <= not(layer1_outputs(2563));
    layer2_outputs(3992) <= '0';
    layer2_outputs(3993) <= layer1_outputs(4077);
    layer2_outputs(3994) <= '0';
    layer2_outputs(3995) <= '0';
    layer2_outputs(3996) <= (layer1_outputs(2265)) and not (layer1_outputs(3493));
    layer2_outputs(3997) <= '1';
    layer2_outputs(3998) <= (layer1_outputs(3700)) and not (layer1_outputs(4329));
    layer2_outputs(3999) <= (layer1_outputs(355)) or (layer1_outputs(515));
    layer2_outputs(4000) <= layer1_outputs(4572);
    layer2_outputs(4001) <= not(layer1_outputs(3581));
    layer2_outputs(4002) <= not(layer1_outputs(2292)) or (layer1_outputs(286));
    layer2_outputs(4003) <= not((layer1_outputs(4489)) or (layer1_outputs(3985)));
    layer2_outputs(4004) <= not(layer1_outputs(668)) or (layer1_outputs(4766));
    layer2_outputs(4005) <= not((layer1_outputs(498)) xor (layer1_outputs(101)));
    layer2_outputs(4006) <= '1';
    layer2_outputs(4007) <= (layer1_outputs(4860)) xor (layer1_outputs(892));
    layer2_outputs(4008) <= '0';
    layer2_outputs(4009) <= '1';
    layer2_outputs(4010) <= not((layer1_outputs(4150)) and (layer1_outputs(3085)));
    layer2_outputs(4011) <= '0';
    layer2_outputs(4012) <= not((layer1_outputs(681)) and (layer1_outputs(3097)));
    layer2_outputs(4013) <= (layer1_outputs(1033)) or (layer1_outputs(2009));
    layer2_outputs(4014) <= not(layer1_outputs(2575)) or (layer1_outputs(3781));
    layer2_outputs(4015) <= (layer1_outputs(1888)) and not (layer1_outputs(445));
    layer2_outputs(4016) <= not(layer1_outputs(1561)) or (layer1_outputs(2486));
    layer2_outputs(4017) <= '0';
    layer2_outputs(4018) <= layer1_outputs(5014);
    layer2_outputs(4019) <= not((layer1_outputs(1034)) or (layer1_outputs(2887)));
    layer2_outputs(4020) <= not((layer1_outputs(4619)) or (layer1_outputs(1825)));
    layer2_outputs(4021) <= (layer1_outputs(1846)) and (layer1_outputs(3642));
    layer2_outputs(4022) <= '1';
    layer2_outputs(4023) <= '0';
    layer2_outputs(4024) <= layer1_outputs(2282);
    layer2_outputs(4025) <= not((layer1_outputs(2953)) or (layer1_outputs(4384)));
    layer2_outputs(4026) <= (layer1_outputs(3956)) and not (layer1_outputs(1450));
    layer2_outputs(4027) <= (layer1_outputs(3)) or (layer1_outputs(4336));
    layer2_outputs(4028) <= (layer1_outputs(3126)) and (layer1_outputs(4974));
    layer2_outputs(4029) <= '1';
    layer2_outputs(4030) <= not(layer1_outputs(3630)) or (layer1_outputs(1720));
    layer2_outputs(4031) <= (layer1_outputs(5004)) and (layer1_outputs(376));
    layer2_outputs(4032) <= '1';
    layer2_outputs(4033) <= (layer1_outputs(3164)) or (layer1_outputs(327));
    layer2_outputs(4034) <= not(layer1_outputs(4877)) or (layer1_outputs(3206));
    layer2_outputs(4035) <= (layer1_outputs(3552)) or (layer1_outputs(1532));
    layer2_outputs(4036) <= '0';
    layer2_outputs(4037) <= (layer1_outputs(193)) xor (layer1_outputs(926));
    layer2_outputs(4038) <= '0';
    layer2_outputs(4039) <= layer1_outputs(4354);
    layer2_outputs(4040) <= layer1_outputs(394);
    layer2_outputs(4041) <= '1';
    layer2_outputs(4042) <= '1';
    layer2_outputs(4043) <= '0';
    layer2_outputs(4044) <= '0';
    layer2_outputs(4045) <= layer1_outputs(1666);
    layer2_outputs(4046) <= (layer1_outputs(1803)) and not (layer1_outputs(3616));
    layer2_outputs(4047) <= '1';
    layer2_outputs(4048) <= not(layer1_outputs(2927));
    layer2_outputs(4049) <= '0';
    layer2_outputs(4050) <= not(layer1_outputs(3204)) or (layer1_outputs(3456));
    layer2_outputs(4051) <= not((layer1_outputs(143)) or (layer1_outputs(3590)));
    layer2_outputs(4052) <= (layer1_outputs(2371)) and not (layer1_outputs(1292));
    layer2_outputs(4053) <= not(layer1_outputs(3566)) or (layer1_outputs(3034));
    layer2_outputs(4054) <= not(layer1_outputs(713));
    layer2_outputs(4055) <= '1';
    layer2_outputs(4056) <= '0';
    layer2_outputs(4057) <= (layer1_outputs(4902)) and (layer1_outputs(2067));
    layer2_outputs(4058) <= (layer1_outputs(1730)) and (layer1_outputs(2166));
    layer2_outputs(4059) <= (layer1_outputs(4044)) or (layer1_outputs(4134));
    layer2_outputs(4060) <= (layer1_outputs(4718)) or (layer1_outputs(3015));
    layer2_outputs(4061) <= '0';
    layer2_outputs(4062) <= '0';
    layer2_outputs(4063) <= not((layer1_outputs(2602)) and (layer1_outputs(981)));
    layer2_outputs(4064) <= '0';
    layer2_outputs(4065) <= (layer1_outputs(4446)) and not (layer1_outputs(2306));
    layer2_outputs(4066) <= not((layer1_outputs(155)) and (layer1_outputs(4405)));
    layer2_outputs(4067) <= (layer1_outputs(3308)) and not (layer1_outputs(711));
    layer2_outputs(4068) <= not((layer1_outputs(1645)) xor (layer1_outputs(2321)));
    layer2_outputs(4069) <= (layer1_outputs(4332)) xor (layer1_outputs(2099));
    layer2_outputs(4070) <= not((layer1_outputs(1171)) and (layer1_outputs(622)));
    layer2_outputs(4071) <= (layer1_outputs(4875)) and not (layer1_outputs(1275));
    layer2_outputs(4072) <= (layer1_outputs(1782)) or (layer1_outputs(4748));
    layer2_outputs(4073) <= not(layer1_outputs(3930));
    layer2_outputs(4074) <= not((layer1_outputs(113)) or (layer1_outputs(4970)));
    layer2_outputs(4075) <= not((layer1_outputs(959)) and (layer1_outputs(4621)));
    layer2_outputs(4076) <= (layer1_outputs(787)) and not (layer1_outputs(3148));
    layer2_outputs(4077) <= not(layer1_outputs(4357));
    layer2_outputs(4078) <= (layer1_outputs(2356)) or (layer1_outputs(1453));
    layer2_outputs(4079) <= not(layer1_outputs(3298));
    layer2_outputs(4080) <= (layer1_outputs(4346)) and not (layer1_outputs(3528));
    layer2_outputs(4081) <= '1';
    layer2_outputs(4082) <= not(layer1_outputs(1099));
    layer2_outputs(4083) <= (layer1_outputs(3189)) and not (layer1_outputs(3994));
    layer2_outputs(4084) <= layer1_outputs(1130);
    layer2_outputs(4085) <= (layer1_outputs(576)) or (layer1_outputs(687));
    layer2_outputs(4086) <= not(layer1_outputs(931));
    layer2_outputs(4087) <= layer1_outputs(3575);
    layer2_outputs(4088) <= not(layer1_outputs(2406));
    layer2_outputs(4089) <= not(layer1_outputs(1550));
    layer2_outputs(4090) <= '1';
    layer2_outputs(4091) <= '0';
    layer2_outputs(4092) <= layer1_outputs(2266);
    layer2_outputs(4093) <= not(layer1_outputs(1371));
    layer2_outputs(4094) <= '1';
    layer2_outputs(4095) <= (layer1_outputs(1299)) and (layer1_outputs(3235));
    layer2_outputs(4096) <= not((layer1_outputs(5089)) or (layer1_outputs(903)));
    layer2_outputs(4097) <= layer1_outputs(3246);
    layer2_outputs(4098) <= (layer1_outputs(3623)) or (layer1_outputs(2380));
    layer2_outputs(4099) <= (layer1_outputs(5096)) and (layer1_outputs(3397));
    layer2_outputs(4100) <= not((layer1_outputs(4182)) and (layer1_outputs(4657)));
    layer2_outputs(4101) <= not((layer1_outputs(3989)) or (layer1_outputs(3579)));
    layer2_outputs(4102) <= not(layer1_outputs(646)) or (layer1_outputs(750));
    layer2_outputs(4103) <= (layer1_outputs(2937)) or (layer1_outputs(4511));
    layer2_outputs(4104) <= not((layer1_outputs(73)) and (layer1_outputs(1688)));
    layer2_outputs(4105) <= not(layer1_outputs(339)) or (layer1_outputs(556));
    layer2_outputs(4106) <= not((layer1_outputs(4510)) and (layer1_outputs(2803)));
    layer2_outputs(4107) <= '1';
    layer2_outputs(4108) <= (layer1_outputs(4687)) and (layer1_outputs(2846));
    layer2_outputs(4109) <= (layer1_outputs(2358)) and not (layer1_outputs(1954));
    layer2_outputs(4110) <= '1';
    layer2_outputs(4111) <= '0';
    layer2_outputs(4112) <= '1';
    layer2_outputs(4113) <= (layer1_outputs(353)) or (layer1_outputs(3535));
    layer2_outputs(4114) <= (layer1_outputs(3841)) and not (layer1_outputs(5109));
    layer2_outputs(4115) <= '1';
    layer2_outputs(4116) <= '1';
    layer2_outputs(4117) <= '0';
    layer2_outputs(4118) <= (layer1_outputs(4888)) and not (layer1_outputs(1686));
    layer2_outputs(4119) <= not(layer1_outputs(663));
    layer2_outputs(4120) <= (layer1_outputs(2658)) and not (layer1_outputs(891));
    layer2_outputs(4121) <= (layer1_outputs(1930)) and not (layer1_outputs(2837));
    layer2_outputs(4122) <= not(layer1_outputs(4974)) or (layer1_outputs(3172));
    layer2_outputs(4123) <= not(layer1_outputs(788));
    layer2_outputs(4124) <= not((layer1_outputs(232)) or (layer1_outputs(1802)));
    layer2_outputs(4125) <= '0';
    layer2_outputs(4126) <= '1';
    layer2_outputs(4127) <= '1';
    layer2_outputs(4128) <= not(layer1_outputs(2653)) or (layer1_outputs(2475));
    layer2_outputs(4129) <= '1';
    layer2_outputs(4130) <= not(layer1_outputs(1853)) or (layer1_outputs(2490));
    layer2_outputs(4131) <= (layer1_outputs(4022)) and not (layer1_outputs(2951));
    layer2_outputs(4132) <= not(layer1_outputs(5115)) or (layer1_outputs(3262));
    layer2_outputs(4133) <= (layer1_outputs(4540)) and (layer1_outputs(1004));
    layer2_outputs(4134) <= (layer1_outputs(833)) or (layer1_outputs(4583));
    layer2_outputs(4135) <= not(layer1_outputs(295)) or (layer1_outputs(5026));
    layer2_outputs(4136) <= not(layer1_outputs(946)) or (layer1_outputs(3165));
    layer2_outputs(4137) <= '1';
    layer2_outputs(4138) <= '1';
    layer2_outputs(4139) <= (layer1_outputs(2962)) xor (layer1_outputs(4414));
    layer2_outputs(4140) <= layer1_outputs(1901);
    layer2_outputs(4141) <= not(layer1_outputs(2550));
    layer2_outputs(4142) <= layer1_outputs(377);
    layer2_outputs(4143) <= not(layer1_outputs(4015));
    layer2_outputs(4144) <= '1';
    layer2_outputs(4145) <= (layer1_outputs(659)) and not (layer1_outputs(5058));
    layer2_outputs(4146) <= not(layer1_outputs(1727));
    layer2_outputs(4147) <= not(layer1_outputs(642)) or (layer1_outputs(2176));
    layer2_outputs(4148) <= (layer1_outputs(4740)) or (layer1_outputs(3848));
    layer2_outputs(4149) <= not(layer1_outputs(3749));
    layer2_outputs(4150) <= '1';
    layer2_outputs(4151) <= '1';
    layer2_outputs(4152) <= not((layer1_outputs(4156)) and (layer1_outputs(2410)));
    layer2_outputs(4153) <= (layer1_outputs(3839)) or (layer1_outputs(4699));
    layer2_outputs(4154) <= not(layer1_outputs(3712)) or (layer1_outputs(4744));
    layer2_outputs(4155) <= not((layer1_outputs(4053)) or (layer1_outputs(422)));
    layer2_outputs(4156) <= not((layer1_outputs(2630)) or (layer1_outputs(4011)));
    layer2_outputs(4157) <= '1';
    layer2_outputs(4158) <= '0';
    layer2_outputs(4159) <= '1';
    layer2_outputs(4160) <= '1';
    layer2_outputs(4161) <= not((layer1_outputs(4185)) or (layer1_outputs(3603)));
    layer2_outputs(4162) <= (layer1_outputs(1026)) or (layer1_outputs(1448));
    layer2_outputs(4163) <= (layer1_outputs(3703)) and not (layer1_outputs(4055));
    layer2_outputs(4164) <= '1';
    layer2_outputs(4165) <= not(layer1_outputs(4387)) or (layer1_outputs(4296));
    layer2_outputs(4166) <= not(layer1_outputs(2672));
    layer2_outputs(4167) <= not((layer1_outputs(5030)) and (layer1_outputs(3047)));
    layer2_outputs(4168) <= (layer1_outputs(1436)) and (layer1_outputs(2505));
    layer2_outputs(4169) <= not(layer1_outputs(2512)) or (layer1_outputs(272));
    layer2_outputs(4170) <= (layer1_outputs(2615)) and not (layer1_outputs(4138));
    layer2_outputs(4171) <= not((layer1_outputs(726)) and (layer1_outputs(4713)));
    layer2_outputs(4172) <= layer1_outputs(839);
    layer2_outputs(4173) <= (layer1_outputs(4515)) and not (layer1_outputs(2144));
    layer2_outputs(4174) <= not(layer1_outputs(1639));
    layer2_outputs(4175) <= not(layer1_outputs(3789)) or (layer1_outputs(4561));
    layer2_outputs(4176) <= layer1_outputs(4552);
    layer2_outputs(4177) <= (layer1_outputs(748)) and not (layer1_outputs(2150));
    layer2_outputs(4178) <= (layer1_outputs(1237)) and not (layer1_outputs(870));
    layer2_outputs(4179) <= '0';
    layer2_outputs(4180) <= '0';
    layer2_outputs(4181) <= (layer1_outputs(420)) and not (layer1_outputs(4378));
    layer2_outputs(4182) <= layer1_outputs(4);
    layer2_outputs(4183) <= (layer1_outputs(3760)) and not (layer1_outputs(2912));
    layer2_outputs(4184) <= layer1_outputs(203);
    layer2_outputs(4185) <= '1';
    layer2_outputs(4186) <= '1';
    layer2_outputs(4187) <= '1';
    layer2_outputs(4188) <= not(layer1_outputs(1717)) or (layer1_outputs(5032));
    layer2_outputs(4189) <= (layer1_outputs(4262)) and (layer1_outputs(4872));
    layer2_outputs(4190) <= '0';
    layer2_outputs(4191) <= not((layer1_outputs(1613)) or (layer1_outputs(200)));
    layer2_outputs(4192) <= '1';
    layer2_outputs(4193) <= (layer1_outputs(3372)) and (layer1_outputs(3313));
    layer2_outputs(4194) <= layer1_outputs(3333);
    layer2_outputs(4195) <= (layer1_outputs(3304)) xor (layer1_outputs(4840));
    layer2_outputs(4196) <= not(layer1_outputs(2920)) or (layer1_outputs(808));
    layer2_outputs(4197) <= not(layer1_outputs(2866)) or (layer1_outputs(753));
    layer2_outputs(4198) <= not(layer1_outputs(2889)) or (layer1_outputs(4563));
    layer2_outputs(4199) <= (layer1_outputs(4861)) and (layer1_outputs(3492));
    layer2_outputs(4200) <= layer1_outputs(3635);
    layer2_outputs(4201) <= (layer1_outputs(1108)) or (layer1_outputs(1968));
    layer2_outputs(4202) <= (layer1_outputs(734)) or (layer1_outputs(1583));
    layer2_outputs(4203) <= (layer1_outputs(4407)) or (layer1_outputs(1067));
    layer2_outputs(4204) <= not((layer1_outputs(2823)) and (layer1_outputs(2871)));
    layer2_outputs(4205) <= (layer1_outputs(119)) or (layer1_outputs(2102));
    layer2_outputs(4206) <= layer1_outputs(228);
    layer2_outputs(4207) <= (layer1_outputs(3826)) and (layer1_outputs(1228));
    layer2_outputs(4208) <= (layer1_outputs(1593)) and not (layer1_outputs(4123));
    layer2_outputs(4209) <= not((layer1_outputs(4917)) and (layer1_outputs(2946)));
    layer2_outputs(4210) <= not(layer1_outputs(106)) or (layer1_outputs(1239));
    layer2_outputs(4211) <= layer1_outputs(3650);
    layer2_outputs(4212) <= (layer1_outputs(1414)) and (layer1_outputs(1195));
    layer2_outputs(4213) <= (layer1_outputs(3955)) xor (layer1_outputs(3931));
    layer2_outputs(4214) <= not((layer1_outputs(4628)) and (layer1_outputs(1302)));
    layer2_outputs(4215) <= '0';
    layer2_outputs(4216) <= not(layer1_outputs(320)) or (layer1_outputs(4051));
    layer2_outputs(4217) <= not((layer1_outputs(2745)) or (layer1_outputs(3319)));
    layer2_outputs(4218) <= (layer1_outputs(597)) and not (layer1_outputs(2443));
    layer2_outputs(4219) <= '0';
    layer2_outputs(4220) <= (layer1_outputs(33)) or (layer1_outputs(2933));
    layer2_outputs(4221) <= (layer1_outputs(3807)) and not (layer1_outputs(725));
    layer2_outputs(4222) <= (layer1_outputs(4758)) and not (layer1_outputs(1234));
    layer2_outputs(4223) <= layer1_outputs(4094);
    layer2_outputs(4224) <= not(layer1_outputs(568));
    layer2_outputs(4225) <= not(layer1_outputs(282)) or (layer1_outputs(4506));
    layer2_outputs(4226) <= '1';
    layer2_outputs(4227) <= layer1_outputs(4976);
    layer2_outputs(4228) <= '0';
    layer2_outputs(4229) <= not((layer1_outputs(4818)) and (layer1_outputs(2838)));
    layer2_outputs(4230) <= not(layer1_outputs(862)) or (layer1_outputs(2273));
    layer2_outputs(4231) <= (layer1_outputs(2925)) or (layer1_outputs(4451));
    layer2_outputs(4232) <= '0';
    layer2_outputs(4233) <= '0';
    layer2_outputs(4234) <= (layer1_outputs(2636)) and not (layer1_outputs(4304));
    layer2_outputs(4235) <= '0';
    layer2_outputs(4236) <= '1';
    layer2_outputs(4237) <= layer1_outputs(2380);
    layer2_outputs(4238) <= '0';
    layer2_outputs(4239) <= not(layer1_outputs(4853));
    layer2_outputs(4240) <= not(layer1_outputs(1086)) or (layer1_outputs(2616));
    layer2_outputs(4241) <= not(layer1_outputs(2873)) or (layer1_outputs(1289));
    layer2_outputs(4242) <= (layer1_outputs(202)) and not (layer1_outputs(2001));
    layer2_outputs(4243) <= not(layer1_outputs(2528));
    layer2_outputs(4244) <= not(layer1_outputs(376));
    layer2_outputs(4245) <= not((layer1_outputs(357)) or (layer1_outputs(2230)));
    layer2_outputs(4246) <= not(layer1_outputs(804)) or (layer1_outputs(1805));
    layer2_outputs(4247) <= layer1_outputs(4044);
    layer2_outputs(4248) <= not(layer1_outputs(60));
    layer2_outputs(4249) <= layer1_outputs(1088);
    layer2_outputs(4250) <= '1';
    layer2_outputs(4251) <= (layer1_outputs(3298)) or (layer1_outputs(940));
    layer2_outputs(4252) <= layer1_outputs(2481);
    layer2_outputs(4253) <= (layer1_outputs(4161)) and not (layer1_outputs(1183));
    layer2_outputs(4254) <= (layer1_outputs(2724)) and not (layer1_outputs(2243));
    layer2_outputs(4255) <= layer1_outputs(36);
    layer2_outputs(4256) <= not(layer1_outputs(1658));
    layer2_outputs(4257) <= not((layer1_outputs(776)) and (layer1_outputs(522)));
    layer2_outputs(4258) <= (layer1_outputs(2529)) or (layer1_outputs(120));
    layer2_outputs(4259) <= (layer1_outputs(184)) and (layer1_outputs(4846));
    layer2_outputs(4260) <= not((layer1_outputs(1545)) xor (layer1_outputs(4375)));
    layer2_outputs(4261) <= not(layer1_outputs(4517));
    layer2_outputs(4262) <= (layer1_outputs(4879)) and not (layer1_outputs(4538));
    layer2_outputs(4263) <= not(layer1_outputs(913));
    layer2_outputs(4264) <= not((layer1_outputs(517)) or (layer1_outputs(955)));
    layer2_outputs(4265) <= not(layer1_outputs(4908)) or (layer1_outputs(2398));
    layer2_outputs(4266) <= '0';
    layer2_outputs(4267) <= not((layer1_outputs(1705)) or (layer1_outputs(1263)));
    layer2_outputs(4268) <= (layer1_outputs(2003)) and (layer1_outputs(2837));
    layer2_outputs(4269) <= '0';
    layer2_outputs(4270) <= (layer1_outputs(5076)) and not (layer1_outputs(3748));
    layer2_outputs(4271) <= layer1_outputs(802);
    layer2_outputs(4272) <= (layer1_outputs(4028)) xor (layer1_outputs(2592));
    layer2_outputs(4273) <= (layer1_outputs(3317)) xor (layer1_outputs(3981));
    layer2_outputs(4274) <= (layer1_outputs(3323)) and (layer1_outputs(3118));
    layer2_outputs(4275) <= '1';
    layer2_outputs(4276) <= layer1_outputs(1536);
    layer2_outputs(4277) <= '0';
    layer2_outputs(4278) <= (layer1_outputs(4186)) and (layer1_outputs(1187));
    layer2_outputs(4279) <= layer1_outputs(4884);
    layer2_outputs(4280) <= '1';
    layer2_outputs(4281) <= (layer1_outputs(2939)) and not (layer1_outputs(458));
    layer2_outputs(4282) <= not((layer1_outputs(2420)) and (layer1_outputs(666)));
    layer2_outputs(4283) <= not(layer1_outputs(613));
    layer2_outputs(4284) <= layer1_outputs(2911);
    layer2_outputs(4285) <= not(layer1_outputs(2743));
    layer2_outputs(4286) <= (layer1_outputs(3612)) and not (layer1_outputs(3406));
    layer2_outputs(4287) <= (layer1_outputs(1658)) and not (layer1_outputs(2449));
    layer2_outputs(4288) <= not((layer1_outputs(4083)) or (layer1_outputs(107)));
    layer2_outputs(4289) <= not(layer1_outputs(3166)) or (layer1_outputs(2161));
    layer2_outputs(4290) <= '0';
    layer2_outputs(4291) <= layer1_outputs(3211);
    layer2_outputs(4292) <= '1';
    layer2_outputs(4293) <= (layer1_outputs(1231)) and not (layer1_outputs(1874));
    layer2_outputs(4294) <= not(layer1_outputs(3288));
    layer2_outputs(4295) <= not((layer1_outputs(3895)) and (layer1_outputs(1097)));
    layer2_outputs(4296) <= (layer1_outputs(1521)) or (layer1_outputs(1832));
    layer2_outputs(4297) <= layer1_outputs(1094);
    layer2_outputs(4298) <= (layer1_outputs(3905)) and (layer1_outputs(1244));
    layer2_outputs(4299) <= (layer1_outputs(3925)) or (layer1_outputs(1653));
    layer2_outputs(4300) <= not(layer1_outputs(2184)) or (layer1_outputs(4752));
    layer2_outputs(4301) <= layer1_outputs(2114);
    layer2_outputs(4302) <= not((layer1_outputs(3077)) or (layer1_outputs(2761)));
    layer2_outputs(4303) <= '1';
    layer2_outputs(4304) <= not((layer1_outputs(1378)) or (layer1_outputs(4508)));
    layer2_outputs(4305) <= (layer1_outputs(3834)) and not (layer1_outputs(2097));
    layer2_outputs(4306) <= (layer1_outputs(1931)) and not (layer1_outputs(3981));
    layer2_outputs(4307) <= not((layer1_outputs(5052)) and (layer1_outputs(1342)));
    layer2_outputs(4308) <= '0';
    layer2_outputs(4309) <= (layer1_outputs(1291)) and (layer1_outputs(4530));
    layer2_outputs(4310) <= layer1_outputs(2883);
    layer2_outputs(4311) <= not(layer1_outputs(1690));
    layer2_outputs(4312) <= '1';
    layer2_outputs(4313) <= (layer1_outputs(722)) and not (layer1_outputs(5060));
    layer2_outputs(4314) <= not(layer1_outputs(2775)) or (layer1_outputs(2516));
    layer2_outputs(4315) <= (layer1_outputs(382)) or (layer1_outputs(4938));
    layer2_outputs(4316) <= '1';
    layer2_outputs(4317) <= (layer1_outputs(963)) and (layer1_outputs(3084));
    layer2_outputs(4318) <= not(layer1_outputs(3893)) or (layer1_outputs(3059));
    layer2_outputs(4319) <= '1';
    layer2_outputs(4320) <= '0';
    layer2_outputs(4321) <= not((layer1_outputs(2308)) or (layer1_outputs(4792)));
    layer2_outputs(4322) <= (layer1_outputs(1457)) and (layer1_outputs(3506));
    layer2_outputs(4323) <= '0';
    layer2_outputs(4324) <= '0';
    layer2_outputs(4325) <= not(layer1_outputs(4128));
    layer2_outputs(4326) <= not(layer1_outputs(3661)) or (layer1_outputs(4563));
    layer2_outputs(4327) <= (layer1_outputs(2404)) and not (layer1_outputs(804));
    layer2_outputs(4328) <= (layer1_outputs(2617)) and not (layer1_outputs(688));
    layer2_outputs(4329) <= not(layer1_outputs(3612));
    layer2_outputs(4330) <= not(layer1_outputs(1074));
    layer2_outputs(4331) <= (layer1_outputs(4423)) and not (layer1_outputs(596));
    layer2_outputs(4332) <= layer1_outputs(2676);
    layer2_outputs(4333) <= (layer1_outputs(4771)) and (layer1_outputs(373));
    layer2_outputs(4334) <= not(layer1_outputs(603));
    layer2_outputs(4335) <= not(layer1_outputs(23)) or (layer1_outputs(1111));
    layer2_outputs(4336) <= not((layer1_outputs(3618)) or (layer1_outputs(773)));
    layer2_outputs(4337) <= (layer1_outputs(2654)) xor (layer1_outputs(2744));
    layer2_outputs(4338) <= not((layer1_outputs(1852)) or (layer1_outputs(4008)));
    layer2_outputs(4339) <= (layer1_outputs(434)) and (layer1_outputs(177));
    layer2_outputs(4340) <= (layer1_outputs(4105)) or (layer1_outputs(263));
    layer2_outputs(4341) <= not(layer1_outputs(5000));
    layer2_outputs(4342) <= not(layer1_outputs(3377)) or (layer1_outputs(4457));
    layer2_outputs(4343) <= layer1_outputs(2972);
    layer2_outputs(4344) <= '0';
    layer2_outputs(4345) <= not((layer1_outputs(1673)) or (layer1_outputs(1830)));
    layer2_outputs(4346) <= (layer1_outputs(2404)) and not (layer1_outputs(4484));
    layer2_outputs(4347) <= (layer1_outputs(4738)) and (layer1_outputs(2125));
    layer2_outputs(4348) <= layer1_outputs(3816);
    layer2_outputs(4349) <= (layer1_outputs(1876)) and not (layer1_outputs(1757));
    layer2_outputs(4350) <= layer1_outputs(4740);
    layer2_outputs(4351) <= '0';
    layer2_outputs(4352) <= (layer1_outputs(2382)) or (layer1_outputs(2679));
    layer2_outputs(4353) <= (layer1_outputs(1920)) and not (layer1_outputs(147));
    layer2_outputs(4354) <= '0';
    layer2_outputs(4355) <= '1';
    layer2_outputs(4356) <= (layer1_outputs(3660)) and not (layer1_outputs(841));
    layer2_outputs(4357) <= not(layer1_outputs(2578));
    layer2_outputs(4358) <= (layer1_outputs(492)) and (layer1_outputs(768));
    layer2_outputs(4359) <= (layer1_outputs(3970)) and not (layer1_outputs(3512));
    layer2_outputs(4360) <= not(layer1_outputs(74)) or (layer1_outputs(3089));
    layer2_outputs(4361) <= (layer1_outputs(3188)) and not (layer1_outputs(908));
    layer2_outputs(4362) <= not((layer1_outputs(4781)) and (layer1_outputs(4026)));
    layer2_outputs(4363) <= not(layer1_outputs(4471)) or (layer1_outputs(2019));
    layer2_outputs(4364) <= layer1_outputs(2229);
    layer2_outputs(4365) <= (layer1_outputs(1280)) and not (layer1_outputs(4709));
    layer2_outputs(4366) <= not(layer1_outputs(3730)) or (layer1_outputs(1999));
    layer2_outputs(4367) <= '0';
    layer2_outputs(4368) <= not(layer1_outputs(2398)) or (layer1_outputs(2156));
    layer2_outputs(4369) <= not(layer1_outputs(1286)) or (layer1_outputs(2552));
    layer2_outputs(4370) <= (layer1_outputs(2084)) or (layer1_outputs(3564));
    layer2_outputs(4371) <= (layer1_outputs(1494)) and (layer1_outputs(716));
    layer2_outputs(4372) <= layer1_outputs(1993);
    layer2_outputs(4373) <= not(layer1_outputs(1657));
    layer2_outputs(4374) <= '1';
    layer2_outputs(4375) <= '0';
    layer2_outputs(4376) <= layer1_outputs(296);
    layer2_outputs(4377) <= layer1_outputs(1903);
    layer2_outputs(4378) <= layer1_outputs(4556);
    layer2_outputs(4379) <= '1';
    layer2_outputs(4380) <= not((layer1_outputs(3049)) and (layer1_outputs(3272)));
    layer2_outputs(4381) <= not((layer1_outputs(2064)) or (layer1_outputs(3596)));
    layer2_outputs(4382) <= not(layer1_outputs(1327)) or (layer1_outputs(876));
    layer2_outputs(4383) <= '1';
    layer2_outputs(4384) <= (layer1_outputs(409)) and not (layer1_outputs(809));
    layer2_outputs(4385) <= not(layer1_outputs(978));
    layer2_outputs(4386) <= not(layer1_outputs(2872)) or (layer1_outputs(4019));
    layer2_outputs(4387) <= '1';
    layer2_outputs(4388) <= '0';
    layer2_outputs(4389) <= '0';
    layer2_outputs(4390) <= '0';
    layer2_outputs(4391) <= (layer1_outputs(1143)) and not (layer1_outputs(1557));
    layer2_outputs(4392) <= layer1_outputs(1795);
    layer2_outputs(4393) <= '1';
    layer2_outputs(4394) <= '0';
    layer2_outputs(4395) <= '1';
    layer2_outputs(4396) <= (layer1_outputs(2456)) or (layer1_outputs(3472));
    layer2_outputs(4397) <= not(layer1_outputs(4856)) or (layer1_outputs(1444));
    layer2_outputs(4398) <= (layer1_outputs(4256)) or (layer1_outputs(782));
    layer2_outputs(4399) <= '0';
    layer2_outputs(4400) <= not((layer1_outputs(2960)) or (layer1_outputs(3928)));
    layer2_outputs(4401) <= '1';
    layer2_outputs(4402) <= '0';
    layer2_outputs(4403) <= (layer1_outputs(2613)) or (layer1_outputs(1222));
    layer2_outputs(4404) <= layer1_outputs(835);
    layer2_outputs(4405) <= not(layer1_outputs(2979)) or (layer1_outputs(486));
    layer2_outputs(4406) <= not(layer1_outputs(3168));
    layer2_outputs(4407) <= (layer1_outputs(2604)) or (layer1_outputs(4418));
    layer2_outputs(4408) <= not((layer1_outputs(1678)) or (layer1_outputs(2724)));
    layer2_outputs(4409) <= '1';
    layer2_outputs(4410) <= not((layer1_outputs(3194)) or (layer1_outputs(4494)));
    layer2_outputs(4411) <= (layer1_outputs(3087)) and not (layer1_outputs(2697));
    layer2_outputs(4412) <= layer1_outputs(4404);
    layer2_outputs(4413) <= (layer1_outputs(783)) and not (layer1_outputs(3689));
    layer2_outputs(4414) <= not((layer1_outputs(1732)) and (layer1_outputs(3410)));
    layer2_outputs(4415) <= '0';
    layer2_outputs(4416) <= (layer1_outputs(4135)) and not (layer1_outputs(1233));
    layer2_outputs(4417) <= '0';
    layer2_outputs(4418) <= layer1_outputs(1592);
    layer2_outputs(4419) <= (layer1_outputs(2166)) and (layer1_outputs(4658));
    layer2_outputs(4420) <= (layer1_outputs(2763)) and not (layer1_outputs(3918));
    layer2_outputs(4421) <= not(layer1_outputs(1952));
    layer2_outputs(4422) <= (layer1_outputs(3511)) and not (layer1_outputs(4549));
    layer2_outputs(4423) <= layer1_outputs(3658);
    layer2_outputs(4424) <= (layer1_outputs(1216)) xor (layer1_outputs(3030));
    layer2_outputs(4425) <= (layer1_outputs(3243)) and not (layer1_outputs(3018));
    layer2_outputs(4426) <= not(layer1_outputs(957)) or (layer1_outputs(3972));
    layer2_outputs(4427) <= not(layer1_outputs(2240));
    layer2_outputs(4428) <= not(layer1_outputs(1969)) or (layer1_outputs(3897));
    layer2_outputs(4429) <= layer1_outputs(3065);
    layer2_outputs(4430) <= layer1_outputs(2918);
    layer2_outputs(4431) <= (layer1_outputs(244)) and not (layer1_outputs(1685));
    layer2_outputs(4432) <= (layer1_outputs(969)) and not (layer1_outputs(2497));
    layer2_outputs(4433) <= layer1_outputs(3975);
    layer2_outputs(4434) <= not(layer1_outputs(3766));
    layer2_outputs(4435) <= not(layer1_outputs(946));
    layer2_outputs(4436) <= layer1_outputs(3026);
    layer2_outputs(4437) <= layer1_outputs(1995);
    layer2_outputs(4438) <= (layer1_outputs(165)) and not (layer1_outputs(2896));
    layer2_outputs(4439) <= (layer1_outputs(2496)) or (layer1_outputs(2711));
    layer2_outputs(4440) <= not(layer1_outputs(1873)) or (layer1_outputs(1807));
    layer2_outputs(4441) <= (layer1_outputs(211)) and (layer1_outputs(4102));
    layer2_outputs(4442) <= not(layer1_outputs(2439)) or (layer1_outputs(3935));
    layer2_outputs(4443) <= '0';
    layer2_outputs(4444) <= '0';
    layer2_outputs(4445) <= (layer1_outputs(772)) and not (layer1_outputs(587));
    layer2_outputs(4446) <= '0';
    layer2_outputs(4447) <= not((layer1_outputs(835)) xor (layer1_outputs(271)));
    layer2_outputs(4448) <= layer1_outputs(3586);
    layer2_outputs(4449) <= not(layer1_outputs(529)) or (layer1_outputs(3902));
    layer2_outputs(4450) <= '0';
    layer2_outputs(4451) <= not(layer1_outputs(2578)) or (layer1_outputs(3470));
    layer2_outputs(4452) <= (layer1_outputs(304)) and not (layer1_outputs(4918));
    layer2_outputs(4453) <= (layer1_outputs(1863)) and not (layer1_outputs(4864));
    layer2_outputs(4454) <= layer1_outputs(2090);
    layer2_outputs(4455) <= layer1_outputs(4925);
    layer2_outputs(4456) <= '1';
    layer2_outputs(4457) <= not(layer1_outputs(1810)) or (layer1_outputs(4646));
    layer2_outputs(4458) <= (layer1_outputs(3011)) and not (layer1_outputs(709));
    layer2_outputs(4459) <= '0';
    layer2_outputs(4460) <= not(layer1_outputs(3425)) or (layer1_outputs(2539));
    layer2_outputs(4461) <= '0';
    layer2_outputs(4462) <= '1';
    layer2_outputs(4463) <= (layer1_outputs(1520)) and (layer1_outputs(2238));
    layer2_outputs(4464) <= not(layer1_outputs(1011));
    layer2_outputs(4465) <= (layer1_outputs(4254)) and not (layer1_outputs(1599));
    layer2_outputs(4466) <= (layer1_outputs(2656)) or (layer1_outputs(923));
    layer2_outputs(4467) <= layer1_outputs(340);
    layer2_outputs(4468) <= '1';
    layer2_outputs(4469) <= not(layer1_outputs(3616)) or (layer1_outputs(4230));
    layer2_outputs(4470) <= layer1_outputs(1438);
    layer2_outputs(4471) <= layer1_outputs(4589);
    layer2_outputs(4472) <= '1';
    layer2_outputs(4473) <= '1';
    layer2_outputs(4474) <= not(layer1_outputs(2728)) or (layer1_outputs(874));
    layer2_outputs(4475) <= '0';
    layer2_outputs(4476) <= (layer1_outputs(390)) and not (layer1_outputs(5047));
    layer2_outputs(4477) <= (layer1_outputs(1979)) and not (layer1_outputs(2473));
    layer2_outputs(4478) <= (layer1_outputs(1305)) and (layer1_outputs(2070));
    layer2_outputs(4479) <= '0';
    layer2_outputs(4480) <= not(layer1_outputs(4614)) or (layer1_outputs(4395));
    layer2_outputs(4481) <= '1';
    layer2_outputs(4482) <= not((layer1_outputs(2124)) and (layer1_outputs(5108)));
    layer2_outputs(4483) <= (layer1_outputs(4091)) and (layer1_outputs(3442));
    layer2_outputs(4484) <= (layer1_outputs(2715)) and not (layer1_outputs(992));
    layer2_outputs(4485) <= (layer1_outputs(2408)) or (layer1_outputs(4349));
    layer2_outputs(4486) <= '1';
    layer2_outputs(4487) <= '1';
    layer2_outputs(4488) <= '0';
    layer2_outputs(4489) <= not(layer1_outputs(3996));
    layer2_outputs(4490) <= layer1_outputs(699);
    layer2_outputs(4491) <= layer1_outputs(4275);
    layer2_outputs(4492) <= '0';
    layer2_outputs(4493) <= (layer1_outputs(978)) and not (layer1_outputs(292));
    layer2_outputs(4494) <= (layer1_outputs(3303)) and (layer1_outputs(1566));
    layer2_outputs(4495) <= (layer1_outputs(463)) or (layer1_outputs(4903));
    layer2_outputs(4496) <= not((layer1_outputs(2395)) and (layer1_outputs(2249)));
    layer2_outputs(4497) <= not(layer1_outputs(252));
    layer2_outputs(4498) <= not(layer1_outputs(535));
    layer2_outputs(4499) <= '0';
    layer2_outputs(4500) <= (layer1_outputs(70)) or (layer1_outputs(2056));
    layer2_outputs(4501) <= '1';
    layer2_outputs(4502) <= not(layer1_outputs(34)) or (layer1_outputs(5016));
    layer2_outputs(4503) <= not(layer1_outputs(1203)) or (layer1_outputs(3484));
    layer2_outputs(4504) <= '1';
    layer2_outputs(4505) <= (layer1_outputs(1584)) and not (layer1_outputs(717));
    layer2_outputs(4506) <= not(layer1_outputs(2053));
    layer2_outputs(4507) <= (layer1_outputs(2203)) and not (layer1_outputs(25));
    layer2_outputs(4508) <= not((layer1_outputs(157)) and (layer1_outputs(2352)));
    layer2_outputs(4509) <= not(layer1_outputs(1677)) or (layer1_outputs(6));
    layer2_outputs(4510) <= layer1_outputs(3331);
    layer2_outputs(4511) <= (layer1_outputs(4082)) and (layer1_outputs(2514));
    layer2_outputs(4512) <= layer1_outputs(3546);
    layer2_outputs(4513) <= not((layer1_outputs(3856)) and (layer1_outputs(3571)));
    layer2_outputs(4514) <= (layer1_outputs(2997)) and not (layer1_outputs(2794));
    layer2_outputs(4515) <= layer1_outputs(1539);
    layer2_outputs(4516) <= '0';
    layer2_outputs(4517) <= (layer1_outputs(3583)) and not (layer1_outputs(1897));
    layer2_outputs(4518) <= '0';
    layer2_outputs(4519) <= not((layer1_outputs(1349)) or (layer1_outputs(911)));
    layer2_outputs(4520) <= '1';
    layer2_outputs(4521) <= not(layer1_outputs(4849));
    layer2_outputs(4522) <= layer1_outputs(480);
    layer2_outputs(4523) <= not(layer1_outputs(2460)) or (layer1_outputs(245));
    layer2_outputs(4524) <= not(layer1_outputs(3832)) or (layer1_outputs(1818));
    layer2_outputs(4525) <= '1';
    layer2_outputs(4526) <= not(layer1_outputs(2218)) or (layer1_outputs(3027));
    layer2_outputs(4527) <= '0';
    layer2_outputs(4528) <= '0';
    layer2_outputs(4529) <= '1';
    layer2_outputs(4530) <= (layer1_outputs(3349)) and not (layer1_outputs(4596));
    layer2_outputs(4531) <= '1';
    layer2_outputs(4532) <= not(layer1_outputs(789));
    layer2_outputs(4533) <= (layer1_outputs(4755)) xor (layer1_outputs(2144));
    layer2_outputs(4534) <= layer1_outputs(4240);
    layer2_outputs(4535) <= (layer1_outputs(139)) and not (layer1_outputs(3952));
    layer2_outputs(4536) <= not(layer1_outputs(4509));
    layer2_outputs(4537) <= '1';
    layer2_outputs(4538) <= not(layer1_outputs(1609)) or (layer1_outputs(1345));
    layer2_outputs(4539) <= not(layer1_outputs(4261));
    layer2_outputs(4540) <= not((layer1_outputs(4680)) xor (layer1_outputs(3678)));
    layer2_outputs(4541) <= layer1_outputs(4326);
    layer2_outputs(4542) <= '1';
    layer2_outputs(4543) <= not(layer1_outputs(1418)) or (layer1_outputs(5114));
    layer2_outputs(4544) <= (layer1_outputs(85)) and (layer1_outputs(4667));
    layer2_outputs(4545) <= (layer1_outputs(4097)) and not (layer1_outputs(1705));
    layer2_outputs(4546) <= not(layer1_outputs(2535));
    layer2_outputs(4547) <= not(layer1_outputs(5)) or (layer1_outputs(4285));
    layer2_outputs(4548) <= not((layer1_outputs(4190)) and (layer1_outputs(1501)));
    layer2_outputs(4549) <= '1';
    layer2_outputs(4550) <= not(layer1_outputs(3943));
    layer2_outputs(4551) <= '0';
    layer2_outputs(4552) <= not((layer1_outputs(4890)) or (layer1_outputs(3444)));
    layer2_outputs(4553) <= not((layer1_outputs(2426)) and (layer1_outputs(2662)));
    layer2_outputs(4554) <= not((layer1_outputs(4604)) and (layer1_outputs(3750)));
    layer2_outputs(4555) <= not(layer1_outputs(839)) or (layer1_outputs(669));
    layer2_outputs(4556) <= '0';
    layer2_outputs(4557) <= (layer1_outputs(1552)) or (layer1_outputs(2545));
    layer2_outputs(4558) <= not(layer1_outputs(4344)) or (layer1_outputs(1761));
    layer2_outputs(4559) <= (layer1_outputs(2155)) and not (layer1_outputs(2138));
    layer2_outputs(4560) <= not(layer1_outputs(5046)) or (layer1_outputs(1509));
    layer2_outputs(4561) <= not(layer1_outputs(2405)) or (layer1_outputs(2103));
    layer2_outputs(4562) <= '1';
    layer2_outputs(4563) <= (layer1_outputs(3830)) and not (layer1_outputs(1603));
    layer2_outputs(4564) <= not(layer1_outputs(370));
    layer2_outputs(4565) <= not(layer1_outputs(843)) or (layer1_outputs(519));
    layer2_outputs(4566) <= (layer1_outputs(3413)) or (layer1_outputs(1865));
    layer2_outputs(4567) <= not(layer1_outputs(4753)) or (layer1_outputs(1364));
    layer2_outputs(4568) <= '0';
    layer2_outputs(4569) <= not((layer1_outputs(2587)) or (layer1_outputs(5050)));
    layer2_outputs(4570) <= (layer1_outputs(1154)) and (layer1_outputs(1466));
    layer2_outputs(4571) <= (layer1_outputs(679)) and not (layer1_outputs(649));
    layer2_outputs(4572) <= layer1_outputs(3598);
    layer2_outputs(4573) <= layer1_outputs(1563);
    layer2_outputs(4574) <= (layer1_outputs(765)) and (layer1_outputs(2072));
    layer2_outputs(4575) <= not((layer1_outputs(55)) or (layer1_outputs(712)));
    layer2_outputs(4576) <= not((layer1_outputs(3801)) or (layer1_outputs(2498)));
    layer2_outputs(4577) <= not((layer1_outputs(1692)) or (layer1_outputs(1227)));
    layer2_outputs(4578) <= (layer1_outputs(2302)) and not (layer1_outputs(3430));
    layer2_outputs(4579) <= '1';
    layer2_outputs(4580) <= not(layer1_outputs(2746)) or (layer1_outputs(3683));
    layer2_outputs(4581) <= '0';
    layer2_outputs(4582) <= (layer1_outputs(2031)) and not (layer1_outputs(3615));
    layer2_outputs(4583) <= not((layer1_outputs(4167)) or (layer1_outputs(988)));
    layer2_outputs(4584) <= not(layer1_outputs(443)) or (layer1_outputs(3936));
    layer2_outputs(4585) <= (layer1_outputs(3117)) or (layer1_outputs(3876));
    layer2_outputs(4586) <= (layer1_outputs(2258)) or (layer1_outputs(3786));
    layer2_outputs(4587) <= layer1_outputs(3667);
    layer2_outputs(4588) <= (layer1_outputs(503)) and (layer1_outputs(2485));
    layer2_outputs(4589) <= not(layer1_outputs(2911)) or (layer1_outputs(3538));
    layer2_outputs(4590) <= (layer1_outputs(5051)) xor (layer1_outputs(178));
    layer2_outputs(4591) <= (layer1_outputs(1106)) and not (layer1_outputs(1732));
    layer2_outputs(4592) <= (layer1_outputs(1186)) or (layer1_outputs(3448));
    layer2_outputs(4593) <= not(layer1_outputs(4043));
    layer2_outputs(4594) <= '1';
    layer2_outputs(4595) <= (layer1_outputs(4906)) xor (layer1_outputs(4828));
    layer2_outputs(4596) <= (layer1_outputs(4390)) or (layer1_outputs(1615));
    layer2_outputs(4597) <= (layer1_outputs(840)) and (layer1_outputs(1066));
    layer2_outputs(4598) <= '1';
    layer2_outputs(4599) <= (layer1_outputs(3095)) or (layer1_outputs(3846));
    layer2_outputs(4600) <= '1';
    layer2_outputs(4601) <= (layer1_outputs(1523)) and not (layer1_outputs(715));
    layer2_outputs(4602) <= '0';
    layer2_outputs(4603) <= (layer1_outputs(4988)) and not (layer1_outputs(3184));
    layer2_outputs(4604) <= '1';
    layer2_outputs(4605) <= '1';
    layer2_outputs(4606) <= '0';
    layer2_outputs(4607) <= not((layer1_outputs(4742)) or (layer1_outputs(3488)));
    layer2_outputs(4608) <= layer1_outputs(3668);
    layer2_outputs(4609) <= not(layer1_outputs(1067));
    layer2_outputs(4610) <= (layer1_outputs(4010)) and not (layer1_outputs(3422));
    layer2_outputs(4611) <= '0';
    layer2_outputs(4612) <= layer1_outputs(3247);
    layer2_outputs(4613) <= not((layer1_outputs(2205)) and (layer1_outputs(1504)));
    layer2_outputs(4614) <= (layer1_outputs(4765)) and not (layer1_outputs(331));
    layer2_outputs(4615) <= '1';
    layer2_outputs(4616) <= '1';
    layer2_outputs(4617) <= not((layer1_outputs(1165)) or (layer1_outputs(1859)));
    layer2_outputs(4618) <= not((layer1_outputs(2057)) and (layer1_outputs(2501)));
    layer2_outputs(4619) <= not(layer1_outputs(759)) or (layer1_outputs(1760));
    layer2_outputs(4620) <= '1';
    layer2_outputs(4621) <= '1';
    layer2_outputs(4622) <= (layer1_outputs(1025)) and not (layer1_outputs(1761));
    layer2_outputs(4623) <= layer1_outputs(3223);
    layer2_outputs(4624) <= layer1_outputs(705);
    layer2_outputs(4625) <= not((layer1_outputs(1272)) or (layer1_outputs(105)));
    layer2_outputs(4626) <= not(layer1_outputs(438));
    layer2_outputs(4627) <= not((layer1_outputs(4193)) or (layer1_outputs(343)));
    layer2_outputs(4628) <= layer1_outputs(780);
    layer2_outputs(4629) <= layer1_outputs(2994);
    layer2_outputs(4630) <= (layer1_outputs(17)) and not (layer1_outputs(4923));
    layer2_outputs(4631) <= not(layer1_outputs(2464)) or (layer1_outputs(3534));
    layer2_outputs(4632) <= not(layer1_outputs(2524)) or (layer1_outputs(600));
    layer2_outputs(4633) <= not(layer1_outputs(4658));
    layer2_outputs(4634) <= not(layer1_outputs(834)) or (layer1_outputs(211));
    layer2_outputs(4635) <= '1';
    layer2_outputs(4636) <= not(layer1_outputs(4512)) or (layer1_outputs(1836));
    layer2_outputs(4637) <= not(layer1_outputs(889)) or (layer1_outputs(1266));
    layer2_outputs(4638) <= (layer1_outputs(1230)) or (layer1_outputs(3130));
    layer2_outputs(4639) <= not(layer1_outputs(2935));
    layer2_outputs(4640) <= (layer1_outputs(1384)) and not (layer1_outputs(3217));
    layer2_outputs(4641) <= not(layer1_outputs(1914));
    layer2_outputs(4642) <= not((layer1_outputs(4271)) and (layer1_outputs(2952)));
    layer2_outputs(4643) <= '1';
    layer2_outputs(4644) <= not(layer1_outputs(1941)) or (layer1_outputs(2207));
    layer2_outputs(4645) <= layer1_outputs(1006);
    layer2_outputs(4646) <= not((layer1_outputs(1425)) and (layer1_outputs(3349)));
    layer2_outputs(4647) <= not(layer1_outputs(585));
    layer2_outputs(4648) <= not((layer1_outputs(5022)) and (layer1_outputs(2093)));
    layer2_outputs(4649) <= not((layer1_outputs(4210)) and (layer1_outputs(4770)));
    layer2_outputs(4650) <= '1';
    layer2_outputs(4651) <= (layer1_outputs(4288)) or (layer1_outputs(4112));
    layer2_outputs(4652) <= not(layer1_outputs(26)) or (layer1_outputs(4255));
    layer2_outputs(4653) <= not(layer1_outputs(1786));
    layer2_outputs(4654) <= '1';
    layer2_outputs(4655) <= not(layer1_outputs(3711)) or (layer1_outputs(2239));
    layer2_outputs(4656) <= '0';
    layer2_outputs(4657) <= not(layer1_outputs(922)) or (layer1_outputs(477));
    layer2_outputs(4658) <= (layer1_outputs(893)) and (layer1_outputs(3374));
    layer2_outputs(4659) <= not(layer1_outputs(4389));
    layer2_outputs(4660) <= '0';
    layer2_outputs(4661) <= not((layer1_outputs(3990)) and (layer1_outputs(1516)));
    layer2_outputs(4662) <= layer1_outputs(1245);
    layer2_outputs(4663) <= (layer1_outputs(3946)) or (layer1_outputs(2193));
    layer2_outputs(4664) <= not(layer1_outputs(2651)) or (layer1_outputs(81));
    layer2_outputs(4665) <= '1';
    layer2_outputs(4666) <= not(layer1_outputs(481));
    layer2_outputs(4667) <= layer1_outputs(1902);
    layer2_outputs(4668) <= not(layer1_outputs(2202)) or (layer1_outputs(2699));
    layer2_outputs(4669) <= '1';
    layer2_outputs(4670) <= (layer1_outputs(4278)) or (layer1_outputs(1104));
    layer2_outputs(4671) <= not((layer1_outputs(3942)) or (layer1_outputs(3575)));
    layer2_outputs(4672) <= not(layer1_outputs(4231)) or (layer1_outputs(768));
    layer2_outputs(4673) <= (layer1_outputs(4661)) and not (layer1_outputs(602));
    layer2_outputs(4674) <= layer1_outputs(2896);
    layer2_outputs(4675) <= not((layer1_outputs(2885)) and (layer1_outputs(1640)));
    layer2_outputs(4676) <= not(layer1_outputs(2635)) or (layer1_outputs(2959));
    layer2_outputs(4677) <= not((layer1_outputs(125)) and (layer1_outputs(2627)));
    layer2_outputs(4678) <= '0';
    layer2_outputs(4679) <= '0';
    layer2_outputs(4680) <= (layer1_outputs(328)) and not (layer1_outputs(4935));
    layer2_outputs(4681) <= (layer1_outputs(4321)) or (layer1_outputs(3261));
    layer2_outputs(4682) <= '0';
    layer2_outputs(4683) <= not(layer1_outputs(1292)) or (layer1_outputs(4521));
    layer2_outputs(4684) <= (layer1_outputs(4920)) and (layer1_outputs(383));
    layer2_outputs(4685) <= '1';
    layer2_outputs(4686) <= (layer1_outputs(1116)) or (layer1_outputs(2781));
    layer2_outputs(4687) <= '1';
    layer2_outputs(4688) <= layer1_outputs(2971);
    layer2_outputs(4689) <= not(layer1_outputs(1728));
    layer2_outputs(4690) <= '1';
    layer2_outputs(4691) <= not((layer1_outputs(3698)) or (layer1_outputs(4492)));
    layer2_outputs(4692) <= '1';
    layer2_outputs(4693) <= not((layer1_outputs(3770)) or (layer1_outputs(1734)));
    layer2_outputs(4694) <= layer1_outputs(605);
    layer2_outputs(4695) <= layer1_outputs(2734);
    layer2_outputs(4696) <= '1';
    layer2_outputs(4697) <= layer1_outputs(1784);
    layer2_outputs(4698) <= layer1_outputs(1549);
    layer2_outputs(4699) <= '1';
    layer2_outputs(4700) <= (layer1_outputs(3753)) or (layer1_outputs(545));
    layer2_outputs(4701) <= not((layer1_outputs(3290)) and (layer1_outputs(2382)));
    layer2_outputs(4702) <= not(layer1_outputs(5043));
    layer2_outputs(4703) <= not((layer1_outputs(2396)) or (layer1_outputs(2575)));
    layer2_outputs(4704) <= not((layer1_outputs(4560)) and (layer1_outputs(941)));
    layer2_outputs(4705) <= '1';
    layer2_outputs(4706) <= layer1_outputs(2436);
    layer2_outputs(4707) <= (layer1_outputs(4764)) and (layer1_outputs(2076));
    layer2_outputs(4708) <= '1';
    layer2_outputs(4709) <= not((layer1_outputs(246)) or (layer1_outputs(1586)));
    layer2_outputs(4710) <= '1';
    layer2_outputs(4711) <= (layer1_outputs(4297)) or (layer1_outputs(1175));
    layer2_outputs(4712) <= not((layer1_outputs(1078)) or (layer1_outputs(4061)));
    layer2_outputs(4713) <= (layer1_outputs(4859)) and not (layer1_outputs(857));
    layer2_outputs(4714) <= not((layer1_outputs(425)) and (layer1_outputs(2526)));
    layer2_outputs(4715) <= '0';
    layer2_outputs(4716) <= layer1_outputs(1839);
    layer2_outputs(4717) <= layer1_outputs(4007);
    layer2_outputs(4718) <= '1';
    layer2_outputs(4719) <= (layer1_outputs(4837)) and not (layer1_outputs(3577));
    layer2_outputs(4720) <= '0';
    layer2_outputs(4721) <= not(layer1_outputs(415)) or (layer1_outputs(4955));
    layer2_outputs(4722) <= '0';
    layer2_outputs(4723) <= not((layer1_outputs(3716)) or (layer1_outputs(3558)));
    layer2_outputs(4724) <= not((layer1_outputs(1575)) or (layer1_outputs(1150)));
    layer2_outputs(4725) <= (layer1_outputs(2827)) and not (layer1_outputs(1284));
    layer2_outputs(4726) <= layer1_outputs(2607);
    layer2_outputs(4727) <= (layer1_outputs(3777)) and not (layer1_outputs(4970));
    layer2_outputs(4728) <= (layer1_outputs(670)) and not (layer1_outputs(4318));
    layer2_outputs(4729) <= '1';
    layer2_outputs(4730) <= not(layer1_outputs(1477));
    layer2_outputs(4731) <= layer1_outputs(2118);
    layer2_outputs(4732) <= not(layer1_outputs(1668)) or (layer1_outputs(69));
    layer2_outputs(4733) <= not(layer1_outputs(4171)) or (layer1_outputs(4178));
    layer2_outputs(4734) <= '0';
    layer2_outputs(4735) <= not((layer1_outputs(2770)) and (layer1_outputs(2417)));
    layer2_outputs(4736) <= '0';
    layer2_outputs(4737) <= '0';
    layer2_outputs(4738) <= not(layer1_outputs(2659)) or (layer1_outputs(1885));
    layer2_outputs(4739) <= '1';
    layer2_outputs(4740) <= not((layer1_outputs(251)) or (layer1_outputs(3206)));
    layer2_outputs(4741) <= not(layer1_outputs(2479));
    layer2_outputs(4742) <= (layer1_outputs(2484)) and not (layer1_outputs(2513));
    layer2_outputs(4743) <= (layer1_outputs(767)) and not (layer1_outputs(3667));
    layer2_outputs(4744) <= '1';
    layer2_outputs(4745) <= (layer1_outputs(2324)) or (layer1_outputs(250));
    layer2_outputs(4746) <= '0';
    layer2_outputs(4747) <= not((layer1_outputs(972)) and (layer1_outputs(1560)));
    layer2_outputs(4748) <= '0';
    layer2_outputs(4749) <= (layer1_outputs(4372)) and (layer1_outputs(1707));
    layer2_outputs(4750) <= (layer1_outputs(4586)) and not (layer1_outputs(1537));
    layer2_outputs(4751) <= not(layer1_outputs(4398));
    layer2_outputs(4752) <= not(layer1_outputs(3724));
    layer2_outputs(4753) <= not((layer1_outputs(591)) xor (layer1_outputs(516)));
    layer2_outputs(4754) <= (layer1_outputs(4386)) and not (layer1_outputs(92));
    layer2_outputs(4755) <= (layer1_outputs(378)) and not (layer1_outputs(2326));
    layer2_outputs(4756) <= not(layer1_outputs(1925)) or (layer1_outputs(472));
    layer2_outputs(4757) <= not(layer1_outputs(3268));
    layer2_outputs(4758) <= not(layer1_outputs(4247));
    layer2_outputs(4759) <= not(layer1_outputs(1225));
    layer2_outputs(4760) <= not(layer1_outputs(1703));
    layer2_outputs(4761) <= not((layer1_outputs(225)) or (layer1_outputs(4245)));
    layer2_outputs(4762) <= '0';
    layer2_outputs(4763) <= layer1_outputs(936);
    layer2_outputs(4764) <= layer1_outputs(4982);
    layer2_outputs(4765) <= not(layer1_outputs(855));
    layer2_outputs(4766) <= not(layer1_outputs(3097));
    layer2_outputs(4767) <= (layer1_outputs(2938)) and not (layer1_outputs(3329));
    layer2_outputs(4768) <= '0';
    layer2_outputs(4769) <= '0';
    layer2_outputs(4770) <= (layer1_outputs(2411)) and not (layer1_outputs(1157));
    layer2_outputs(4771) <= '0';
    layer2_outputs(4772) <= (layer1_outputs(3329)) and not (layer1_outputs(2676));
    layer2_outputs(4773) <= '1';
    layer2_outputs(4774) <= '1';
    layer2_outputs(4775) <= (layer1_outputs(1182)) or (layer1_outputs(921));
    layer2_outputs(4776) <= '1';
    layer2_outputs(4777) <= (layer1_outputs(1667)) or (layer1_outputs(4141));
    layer2_outputs(4778) <= '0';
    layer2_outputs(4779) <= (layer1_outputs(2022)) or (layer1_outputs(1499));
    layer2_outputs(4780) <= (layer1_outputs(163)) and not (layer1_outputs(24));
    layer2_outputs(4781) <= not(layer1_outputs(4051)) or (layer1_outputs(1535));
    layer2_outputs(4782) <= '0';
    layer2_outputs(4783) <= layer1_outputs(1318);
    layer2_outputs(4784) <= not(layer1_outputs(615)) or (layer1_outputs(68));
    layer2_outputs(4785) <= (layer1_outputs(2879)) or (layer1_outputs(1366));
    layer2_outputs(4786) <= (layer1_outputs(3060)) and not (layer1_outputs(2693));
    layer2_outputs(4787) <= not((layer1_outputs(1107)) or (layer1_outputs(1334)));
    layer2_outputs(4788) <= not(layer1_outputs(4234)) or (layer1_outputs(1375));
    layer2_outputs(4789) <= not((layer1_outputs(5019)) or (layer1_outputs(1730)));
    layer2_outputs(4790) <= '1';
    layer2_outputs(4791) <= not(layer1_outputs(4626));
    layer2_outputs(4792) <= layer1_outputs(4474);
    layer2_outputs(4793) <= '1';
    layer2_outputs(4794) <= not((layer1_outputs(1055)) and (layer1_outputs(475)));
    layer2_outputs(4795) <= layer1_outputs(3351);
    layer2_outputs(4796) <= (layer1_outputs(3195)) and not (layer1_outputs(5107));
    layer2_outputs(4797) <= not(layer1_outputs(4084));
    layer2_outputs(4798) <= not(layer1_outputs(3888));
    layer2_outputs(4799) <= '0';
    layer2_outputs(4800) <= (layer1_outputs(4631)) and not (layer1_outputs(2213));
    layer2_outputs(4801) <= '0';
    layer2_outputs(4802) <= not(layer1_outputs(3464)) or (layer1_outputs(595));
    layer2_outputs(4803) <= layer1_outputs(3270);
    layer2_outputs(4804) <= '1';
    layer2_outputs(4805) <= layer1_outputs(4102);
    layer2_outputs(4806) <= not((layer1_outputs(742)) or (layer1_outputs(1104)));
    layer2_outputs(4807) <= '0';
    layer2_outputs(4808) <= layer1_outputs(1894);
    layer2_outputs(4809) <= '0';
    layer2_outputs(4810) <= (layer1_outputs(2032)) and (layer1_outputs(4676));
    layer2_outputs(4811) <= (layer1_outputs(3549)) and not (layer1_outputs(4769));
    layer2_outputs(4812) <= '0';
    layer2_outputs(4813) <= '0';
    layer2_outputs(4814) <= not((layer1_outputs(2750)) or (layer1_outputs(3113)));
    layer2_outputs(4815) <= (layer1_outputs(2557)) and not (layer1_outputs(352));
    layer2_outputs(4816) <= not(layer1_outputs(2673));
    layer2_outputs(4817) <= not((layer1_outputs(4311)) or (layer1_outputs(505)));
    layer2_outputs(4818) <= not((layer1_outputs(2502)) or (layer1_outputs(696)));
    layer2_outputs(4819) <= '0';
    layer2_outputs(4820) <= not(layer1_outputs(4305)) or (layer1_outputs(2455));
    layer2_outputs(4821) <= '1';
    layer2_outputs(4822) <= (layer1_outputs(1397)) and not (layer1_outputs(3461));
    layer2_outputs(4823) <= not(layer1_outputs(4248)) or (layer1_outputs(4200));
    layer2_outputs(4824) <= not((layer1_outputs(2152)) and (layer1_outputs(2314)));
    layer2_outputs(4825) <= not((layer1_outputs(636)) or (layer1_outputs(4514)));
    layer2_outputs(4826) <= not(layer1_outputs(1932));
    layer2_outputs(4827) <= (layer1_outputs(2292)) and not (layer1_outputs(1419));
    layer2_outputs(4828) <= (layer1_outputs(3198)) and not (layer1_outputs(2608));
    layer2_outputs(4829) <= (layer1_outputs(1848)) and not (layer1_outputs(1849));
    layer2_outputs(4830) <= layer1_outputs(3795);
    layer2_outputs(4831) <= (layer1_outputs(89)) and (layer1_outputs(4548));
    layer2_outputs(4832) <= (layer1_outputs(372)) or (layer1_outputs(1714));
    layer2_outputs(4833) <= not(layer1_outputs(1938)) or (layer1_outputs(208));
    layer2_outputs(4834) <= layer1_outputs(691);
    layer2_outputs(4835) <= layer1_outputs(4402);
    layer2_outputs(4836) <= (layer1_outputs(141)) or (layer1_outputs(1300));
    layer2_outputs(4837) <= (layer1_outputs(4842)) and not (layer1_outputs(4290));
    layer2_outputs(4838) <= layer1_outputs(3253);
    layer2_outputs(4839) <= '1';
    layer2_outputs(4840) <= '1';
    layer2_outputs(4841) <= '0';
    layer2_outputs(4842) <= (layer1_outputs(4240)) and (layer1_outputs(2876));
    layer2_outputs(4843) <= (layer1_outputs(3455)) and (layer1_outputs(3823));
    layer2_outputs(4844) <= '0';
    layer2_outputs(4845) <= not(layer1_outputs(2431)) or (layer1_outputs(543));
    layer2_outputs(4846) <= '0';
    layer2_outputs(4847) <= not(layer1_outputs(1582));
    layer2_outputs(4848) <= not(layer1_outputs(2983));
    layer2_outputs(4849) <= (layer1_outputs(5038)) or (layer1_outputs(3149));
    layer2_outputs(4850) <= not(layer1_outputs(4601)) or (layer1_outputs(1232));
    layer2_outputs(4851) <= not((layer1_outputs(5111)) and (layer1_outputs(4048)));
    layer2_outputs(4852) <= (layer1_outputs(4988)) and (layer1_outputs(344));
    layer2_outputs(4853) <= '1';
    layer2_outputs(4854) <= not(layer1_outputs(992));
    layer2_outputs(4855) <= (layer1_outputs(792)) or (layer1_outputs(1718));
    layer2_outputs(4856) <= not(layer1_outputs(3068)) or (layer1_outputs(3075));
    layer2_outputs(4857) <= not(layer1_outputs(4647)) or (layer1_outputs(1877));
    layer2_outputs(4858) <= '0';
    layer2_outputs(4859) <= not((layer1_outputs(1855)) or (layer1_outputs(2074)));
    layer2_outputs(4860) <= (layer1_outputs(1639)) and not (layer1_outputs(5090));
    layer2_outputs(4861) <= not(layer1_outputs(4606));
    layer2_outputs(4862) <= (layer1_outputs(2269)) and not (layer1_outputs(2917));
    layer2_outputs(4863) <= not(layer1_outputs(670)) or (layer1_outputs(561));
    layer2_outputs(4864) <= (layer1_outputs(3890)) and (layer1_outputs(1352));
    layer2_outputs(4865) <= '1';
    layer2_outputs(4866) <= not(layer1_outputs(4368)) or (layer1_outputs(3930));
    layer2_outputs(4867) <= '1';
    layer2_outputs(4868) <= layer1_outputs(2198);
    layer2_outputs(4869) <= '1';
    layer2_outputs(4870) <= '1';
    layer2_outputs(4871) <= not(layer1_outputs(2745));
    layer2_outputs(4872) <= '1';
    layer2_outputs(4873) <= (layer1_outputs(2)) and (layer1_outputs(2543));
    layer2_outputs(4874) <= layer1_outputs(4683);
    layer2_outputs(4875) <= not((layer1_outputs(661)) or (layer1_outputs(5005)));
    layer2_outputs(4876) <= not((layer1_outputs(1962)) xor (layer1_outputs(33)));
    layer2_outputs(4877) <= (layer1_outputs(3995)) and not (layer1_outputs(3208));
    layer2_outputs(4878) <= '0';
    layer2_outputs(4879) <= '1';
    layer2_outputs(4880) <= (layer1_outputs(4756)) and (layer1_outputs(2984));
    layer2_outputs(4881) <= (layer1_outputs(3889)) and not (layer1_outputs(1437));
    layer2_outputs(4882) <= (layer1_outputs(48)) and not (layer1_outputs(3967));
    layer2_outputs(4883) <= layer1_outputs(3949);
    layer2_outputs(4884) <= not(layer1_outputs(4736));
    layer2_outputs(4885) <= '0';
    layer2_outputs(4886) <= not(layer1_outputs(3325)) or (layer1_outputs(2677));
    layer2_outputs(4887) <= (layer1_outputs(3545)) and (layer1_outputs(3747));
    layer2_outputs(4888) <= not(layer1_outputs(735)) or (layer1_outputs(318));
    layer2_outputs(4889) <= (layer1_outputs(2564)) or (layer1_outputs(4096));
    layer2_outputs(4890) <= layer1_outputs(4659);
    layer2_outputs(4891) <= layer1_outputs(3201);
    layer2_outputs(4892) <= not((layer1_outputs(5067)) xor (layer1_outputs(4185)));
    layer2_outputs(4893) <= layer1_outputs(3090);
    layer2_outputs(4894) <= (layer1_outputs(4677)) and not (layer1_outputs(1745));
    layer2_outputs(4895) <= not(layer1_outputs(1764));
    layer2_outputs(4896) <= '1';
    layer2_outputs(4897) <= not(layer1_outputs(1856)) or (layer1_outputs(2462));
    layer2_outputs(4898) <= '1';
    layer2_outputs(4899) <= '1';
    layer2_outputs(4900) <= '1';
    layer2_outputs(4901) <= (layer1_outputs(1550)) and not (layer1_outputs(1733));
    layer2_outputs(4902) <= (layer1_outputs(1000)) or (layer1_outputs(4920));
    layer2_outputs(4903) <= (layer1_outputs(2226)) and not (layer1_outputs(181));
    layer2_outputs(4904) <= not(layer1_outputs(2083));
    layer2_outputs(4905) <= (layer1_outputs(2944)) and not (layer1_outputs(1571));
    layer2_outputs(4906) <= '0';
    layer2_outputs(4907) <= (layer1_outputs(3360)) and (layer1_outputs(2277));
    layer2_outputs(4908) <= not(layer1_outputs(385));
    layer2_outputs(4909) <= '1';
    layer2_outputs(4910) <= (layer1_outputs(220)) and not (layer1_outputs(542));
    layer2_outputs(4911) <= '1';
    layer2_outputs(4912) <= (layer1_outputs(1416)) or (layer1_outputs(3373));
    layer2_outputs(4913) <= (layer1_outputs(4759)) and (layer1_outputs(4643));
    layer2_outputs(4914) <= (layer1_outputs(4377)) and not (layer1_outputs(3519));
    layer2_outputs(4915) <= not((layer1_outputs(3727)) or (layer1_outputs(3785)));
    layer2_outputs(4916) <= (layer1_outputs(300)) and not (layer1_outputs(428));
    layer2_outputs(4917) <= not((layer1_outputs(1679)) and (layer1_outputs(429)));
    layer2_outputs(4918) <= not(layer1_outputs(797));
    layer2_outputs(4919) <= (layer1_outputs(4184)) and (layer1_outputs(2855));
    layer2_outputs(4920) <= (layer1_outputs(191)) and not (layer1_outputs(3396));
    layer2_outputs(4921) <= '1';
    layer2_outputs(4922) <= (layer1_outputs(3647)) or (layer1_outputs(3654));
    layer2_outputs(4923) <= '1';
    layer2_outputs(4924) <= (layer1_outputs(4558)) and not (layer1_outputs(4075));
    layer2_outputs(4925) <= '1';
    layer2_outputs(4926) <= not((layer1_outputs(1741)) or (layer1_outputs(424)));
    layer2_outputs(4927) <= '0';
    layer2_outputs(4928) <= layer1_outputs(509);
    layer2_outputs(4929) <= layer1_outputs(181);
    layer2_outputs(4930) <= not(layer1_outputs(4206));
    layer2_outputs(4931) <= (layer1_outputs(4488)) and not (layer1_outputs(4779));
    layer2_outputs(4932) <= (layer1_outputs(3470)) or (layer1_outputs(3614));
    layer2_outputs(4933) <= not(layer1_outputs(918));
    layer2_outputs(4934) <= layer1_outputs(1724);
    layer2_outputs(4935) <= '0';
    layer2_outputs(4936) <= (layer1_outputs(5114)) and not (layer1_outputs(649));
    layer2_outputs(4937) <= '0';
    layer2_outputs(4938) <= '0';
    layer2_outputs(4939) <= '0';
    layer2_outputs(4940) <= layer1_outputs(289);
    layer2_outputs(4941) <= not(layer1_outputs(1279)) or (layer1_outputs(1181));
    layer2_outputs(4942) <= not((layer1_outputs(2029)) and (layer1_outputs(722)));
    layer2_outputs(4943) <= layer1_outputs(4317);
    layer2_outputs(4944) <= layer1_outputs(848);
    layer2_outputs(4945) <= not((layer1_outputs(2992)) or (layer1_outputs(3892)));
    layer2_outputs(4946) <= not((layer1_outputs(1131)) or (layer1_outputs(2106)));
    layer2_outputs(4947) <= (layer1_outputs(2261)) and not (layer1_outputs(4091));
    layer2_outputs(4948) <= layer1_outputs(1665);
    layer2_outputs(4949) <= (layer1_outputs(4998)) and not (layer1_outputs(2250));
    layer2_outputs(4950) <= '1';
    layer2_outputs(4951) <= layer1_outputs(3655);
    layer2_outputs(4952) <= (layer1_outputs(1280)) and not (layer1_outputs(4961));
    layer2_outputs(4953) <= (layer1_outputs(150)) and not (layer1_outputs(627));
    layer2_outputs(4954) <= not((layer1_outputs(2796)) or (layer1_outputs(100)));
    layer2_outputs(4955) <= (layer1_outputs(1858)) and not (layer1_outputs(3693));
    layer2_outputs(4956) <= layer1_outputs(3817);
    layer2_outputs(4957) <= layer1_outputs(3408);
    layer2_outputs(4958) <= (layer1_outputs(3810)) and not (layer1_outputs(3676));
    layer2_outputs(4959) <= (layer1_outputs(862)) and not (layer1_outputs(3875));
    layer2_outputs(4960) <= layer1_outputs(1174);
    layer2_outputs(4961) <= not((layer1_outputs(1989)) or (layer1_outputs(4381)));
    layer2_outputs(4962) <= (layer1_outputs(2566)) and not (layer1_outputs(3491));
    layer2_outputs(4963) <= '0';
    layer2_outputs(4964) <= not(layer1_outputs(3557));
    layer2_outputs(4965) <= not((layer1_outputs(2454)) or (layer1_outputs(1870)));
    layer2_outputs(4966) <= not((layer1_outputs(4881)) and (layer1_outputs(4513)));
    layer2_outputs(4967) <= not((layer1_outputs(2987)) or (layer1_outputs(3697)));
    layer2_outputs(4968) <= not(layer1_outputs(3687));
    layer2_outputs(4969) <= not(layer1_outputs(2444));
    layer2_outputs(4970) <= (layer1_outputs(1997)) xor (layer1_outputs(3820));
    layer2_outputs(4971) <= '1';
    layer2_outputs(4972) <= '1';
    layer2_outputs(4973) <= layer1_outputs(3130);
    layer2_outputs(4974) <= '0';
    layer2_outputs(4975) <= (layer1_outputs(3605)) or (layer1_outputs(4250));
    layer2_outputs(4976) <= (layer1_outputs(2700)) and not (layer1_outputs(3988));
    layer2_outputs(4977) <= (layer1_outputs(1896)) or (layer1_outputs(3541));
    layer2_outputs(4978) <= (layer1_outputs(3072)) and (layer1_outputs(2628));
    layer2_outputs(4979) <= not(layer1_outputs(3039));
    layer2_outputs(4980) <= not(layer1_outputs(4799)) or (layer1_outputs(2951));
    layer2_outputs(4981) <= layer1_outputs(1819);
    layer2_outputs(4982) <= not((layer1_outputs(10)) or (layer1_outputs(3429)));
    layer2_outputs(4983) <= not((layer1_outputs(967)) or (layer1_outputs(2531)));
    layer2_outputs(4984) <= (layer1_outputs(3941)) and not (layer1_outputs(2070));
    layer2_outputs(4985) <= layer1_outputs(308);
    layer2_outputs(4986) <= not((layer1_outputs(4787)) or (layer1_outputs(4107)));
    layer2_outputs(4987) <= (layer1_outputs(2087)) and (layer1_outputs(3128));
    layer2_outputs(4988) <= not((layer1_outputs(16)) and (layer1_outputs(680)));
    layer2_outputs(4989) <= '1';
    layer2_outputs(4990) <= not((layer1_outputs(4708)) or (layer1_outputs(2050)));
    layer2_outputs(4991) <= (layer1_outputs(379)) and not (layer1_outputs(4311));
    layer2_outputs(4992) <= '0';
    layer2_outputs(4993) <= (layer1_outputs(2590)) or (layer1_outputs(5075));
    layer2_outputs(4994) <= not(layer1_outputs(3486));
    layer2_outputs(4995) <= not((layer1_outputs(112)) and (layer1_outputs(4293)));
    layer2_outputs(4996) <= (layer1_outputs(3456)) or (layer1_outputs(1507));
    layer2_outputs(4997) <= not(layer1_outputs(3200));
    layer2_outputs(4998) <= not((layer1_outputs(824)) and (layer1_outputs(4919)));
    layer2_outputs(4999) <= not(layer1_outputs(1949)) or (layer1_outputs(3352));
    layer2_outputs(5000) <= '0';
    layer2_outputs(5001) <= (layer1_outputs(4098)) or (layer1_outputs(1758));
    layer2_outputs(5002) <= not((layer1_outputs(3230)) and (layer1_outputs(4473)));
    layer2_outputs(5003) <= (layer1_outputs(1734)) and not (layer1_outputs(1017));
    layer2_outputs(5004) <= '1';
    layer2_outputs(5005) <= not(layer1_outputs(1478)) or (layer1_outputs(4170));
    layer2_outputs(5006) <= (layer1_outputs(3711)) and not (layer1_outputs(3829));
    layer2_outputs(5007) <= (layer1_outputs(1159)) and (layer1_outputs(686));
    layer2_outputs(5008) <= not(layer1_outputs(1588)) or (layer1_outputs(4557));
    layer2_outputs(5009) <= not((layer1_outputs(326)) and (layer1_outputs(4620)));
    layer2_outputs(5010) <= not((layer1_outputs(4676)) xor (layer1_outputs(2895)));
    layer2_outputs(5011) <= (layer1_outputs(2774)) and not (layer1_outputs(593));
    layer2_outputs(5012) <= (layer1_outputs(3066)) or (layer1_outputs(5094));
    layer2_outputs(5013) <= not(layer1_outputs(5017)) or (layer1_outputs(3144));
    layer2_outputs(5014) <= not(layer1_outputs(603)) or (layer1_outputs(1282));
    layer2_outputs(5015) <= layer1_outputs(853);
    layer2_outputs(5016) <= (layer1_outputs(4650)) and (layer1_outputs(2360));
    layer2_outputs(5017) <= not(layer1_outputs(1811));
    layer2_outputs(5018) <= not((layer1_outputs(4986)) xor (layer1_outputs(3911)));
    layer2_outputs(5019) <= (layer1_outputs(4868)) and (layer1_outputs(531));
    layer2_outputs(5020) <= '1';
    layer2_outputs(5021) <= '1';
    layer2_outputs(5022) <= '1';
    layer2_outputs(5023) <= (layer1_outputs(0)) and (layer1_outputs(3799));
    layer2_outputs(5024) <= '0';
    layer2_outputs(5025) <= (layer1_outputs(1588)) or (layer1_outputs(454));
    layer2_outputs(5026) <= not((layer1_outputs(3756)) and (layer1_outputs(487)));
    layer2_outputs(5027) <= layer1_outputs(197);
    layer2_outputs(5028) <= not((layer1_outputs(932)) and (layer1_outputs(2948)));
    layer2_outputs(5029) <= (layer1_outputs(4252)) and (layer1_outputs(4118));
    layer2_outputs(5030) <= (layer1_outputs(4814)) and not (layer1_outputs(3502));
    layer2_outputs(5031) <= not(layer1_outputs(4572)) or (layer1_outputs(783));
    layer2_outputs(5032) <= layer1_outputs(3511);
    layer2_outputs(5033) <= not(layer1_outputs(4121)) or (layer1_outputs(213));
    layer2_outputs(5034) <= '1';
    layer2_outputs(5035) <= not(layer1_outputs(1027)) or (layer1_outputs(882));
    layer2_outputs(5036) <= not(layer1_outputs(1680)) or (layer1_outputs(3962));
    layer2_outputs(5037) <= '0';
    layer2_outputs(5038) <= '1';
    layer2_outputs(5039) <= not(layer1_outputs(2345));
    layer2_outputs(5040) <= not(layer1_outputs(3153)) or (layer1_outputs(2085));
    layer2_outputs(5041) <= layer1_outputs(2631);
    layer2_outputs(5042) <= not((layer1_outputs(462)) and (layer1_outputs(2206)));
    layer2_outputs(5043) <= '0';
    layer2_outputs(5044) <= not((layer1_outputs(2847)) and (layer1_outputs(1802)));
    layer2_outputs(5045) <= (layer1_outputs(4509)) and (layer1_outputs(57));
    layer2_outputs(5046) <= not(layer1_outputs(4281));
    layer2_outputs(5047) <= not(layer1_outputs(268)) or (layer1_outputs(1395));
    layer2_outputs(5048) <= layer1_outputs(1736);
    layer2_outputs(5049) <= '1';
    layer2_outputs(5050) <= not((layer1_outputs(4213)) or (layer1_outputs(1751)));
    layer2_outputs(5051) <= not((layer1_outputs(11)) or (layer1_outputs(3584)));
    layer2_outputs(5052) <= (layer1_outputs(1032)) and not (layer1_outputs(1246));
    layer2_outputs(5053) <= (layer1_outputs(4604)) and (layer1_outputs(468));
    layer2_outputs(5054) <= not((layer1_outputs(1393)) or (layer1_outputs(646)));
    layer2_outputs(5055) <= layer1_outputs(3703);
    layer2_outputs(5056) <= (layer1_outputs(608)) and (layer1_outputs(1095));
    layer2_outputs(5057) <= (layer1_outputs(3696)) and (layer1_outputs(2486));
    layer2_outputs(5058) <= '0';
    layer2_outputs(5059) <= not(layer1_outputs(1945));
    layer2_outputs(5060) <= not((layer1_outputs(1599)) and (layer1_outputs(698)));
    layer2_outputs(5061) <= '1';
    layer2_outputs(5062) <= not((layer1_outputs(3355)) and (layer1_outputs(1447)));
    layer2_outputs(5063) <= (layer1_outputs(1333)) and not (layer1_outputs(4374));
    layer2_outputs(5064) <= layer1_outputs(3233);
    layer2_outputs(5065) <= (layer1_outputs(3780)) and (layer1_outputs(1607));
    layer2_outputs(5066) <= layer1_outputs(2257);
    layer2_outputs(5067) <= layer1_outputs(3873);
    layer2_outputs(5068) <= not((layer1_outputs(2870)) or (layer1_outputs(4536)));
    layer2_outputs(5069) <= not(layer1_outputs(4450)) or (layer1_outputs(2355));
    layer2_outputs(5070) <= not(layer1_outputs(3664)) or (layer1_outputs(3252));
    layer2_outputs(5071) <= (layer1_outputs(4967)) or (layer1_outputs(1584));
    layer2_outputs(5072) <= not(layer1_outputs(2043)) or (layer1_outputs(1562));
    layer2_outputs(5073) <= not(layer1_outputs(1090)) or (layer1_outputs(1699));
    layer2_outputs(5074) <= (layer1_outputs(3560)) or (layer1_outputs(5040));
    layer2_outputs(5075) <= layer1_outputs(2512);
    layer2_outputs(5076) <= '1';
    layer2_outputs(5077) <= layer1_outputs(2112);
    layer2_outputs(5078) <= not((layer1_outputs(2298)) and (layer1_outputs(3012)));
    layer2_outputs(5079) <= '1';
    layer2_outputs(5080) <= (layer1_outputs(1908)) and not (layer1_outputs(3768));
    layer2_outputs(5081) <= (layer1_outputs(5080)) and (layer1_outputs(3389));
    layer2_outputs(5082) <= (layer1_outputs(718)) and not (layer1_outputs(2597));
    layer2_outputs(5083) <= '0';
    layer2_outputs(5084) <= not(layer1_outputs(2136));
    layer2_outputs(5085) <= '1';
    layer2_outputs(5086) <= (layer1_outputs(545)) and not (layer1_outputs(264));
    layer2_outputs(5087) <= (layer1_outputs(3074)) and not (layer1_outputs(543));
    layer2_outputs(5088) <= not(layer1_outputs(1570)) or (layer1_outputs(5117));
    layer2_outputs(5089) <= not((layer1_outputs(3385)) and (layer1_outputs(3883)));
    layer2_outputs(5090) <= not(layer1_outputs(960)) or (layer1_outputs(859));
    layer2_outputs(5091) <= not(layer1_outputs(26)) or (layer1_outputs(4881));
    layer2_outputs(5092) <= not((layer1_outputs(391)) or (layer1_outputs(3073)));
    layer2_outputs(5093) <= not((layer1_outputs(3503)) or (layer1_outputs(1498)));
    layer2_outputs(5094) <= (layer1_outputs(4939)) and (layer1_outputs(4632));
    layer2_outputs(5095) <= (layer1_outputs(1495)) xor (layer1_outputs(4096));
    layer2_outputs(5096) <= '1';
    layer2_outputs(5097) <= (layer1_outputs(2015)) and not (layer1_outputs(2180));
    layer2_outputs(5098) <= layer1_outputs(557);
    layer2_outputs(5099) <= (layer1_outputs(4689)) and not (layer1_outputs(3871));
    layer2_outputs(5100) <= '1';
    layer2_outputs(5101) <= '1';
    layer2_outputs(5102) <= layer1_outputs(4739);
    layer2_outputs(5103) <= (layer1_outputs(1877)) and not (layer1_outputs(1773));
    layer2_outputs(5104) <= (layer1_outputs(3353)) or (layer1_outputs(4424));
    layer2_outputs(5105) <= not(layer1_outputs(2348)) or (layer1_outputs(1645));
    layer2_outputs(5106) <= '1';
    layer2_outputs(5107) <= (layer1_outputs(3532)) and not (layer1_outputs(2294));
    layer2_outputs(5108) <= layer1_outputs(4825);
    layer2_outputs(5109) <= '0';
    layer2_outputs(5110) <= not((layer1_outputs(3337)) or (layer1_outputs(2759)));
    layer2_outputs(5111) <= not(layer1_outputs(1393));
    layer2_outputs(5112) <= not((layer1_outputs(3385)) or (layer1_outputs(3209)));
    layer2_outputs(5113) <= layer1_outputs(5042);
    layer2_outputs(5114) <= not(layer1_outputs(2783));
    layer2_outputs(5115) <= (layer1_outputs(3492)) and not (layer1_outputs(3509));
    layer2_outputs(5116) <= not(layer1_outputs(4366));
    layer2_outputs(5117) <= not((layer1_outputs(3683)) or (layer1_outputs(2174)));
    layer2_outputs(5118) <= not((layer1_outputs(2264)) and (layer1_outputs(3992)));
    layer2_outputs(5119) <= (layer1_outputs(4481)) or (layer1_outputs(2596));
    layer3_outputs(0) <= not(layer2_outputs(899)) or (layer2_outputs(3825));
    layer3_outputs(1) <= '0';
    layer3_outputs(2) <= not(layer2_outputs(3630));
    layer3_outputs(3) <= (layer2_outputs(168)) and (layer2_outputs(1848));
    layer3_outputs(4) <= not((layer2_outputs(3192)) and (layer2_outputs(3396)));
    layer3_outputs(5) <= '0';
    layer3_outputs(6) <= (layer2_outputs(1611)) or (layer2_outputs(2672));
    layer3_outputs(7) <= not((layer2_outputs(4136)) or (layer2_outputs(1688)));
    layer3_outputs(8) <= '0';
    layer3_outputs(9) <= layer2_outputs(2087);
    layer3_outputs(10) <= not((layer2_outputs(2109)) and (layer2_outputs(2017)));
    layer3_outputs(11) <= layer2_outputs(3806);
    layer3_outputs(12) <= (layer2_outputs(2629)) or (layer2_outputs(4428));
    layer3_outputs(13) <= '0';
    layer3_outputs(14) <= not((layer2_outputs(2877)) or (layer2_outputs(2280)));
    layer3_outputs(15) <= '0';
    layer3_outputs(16) <= (layer2_outputs(1218)) and not (layer2_outputs(1030));
    layer3_outputs(17) <= not(layer2_outputs(1874)) or (layer2_outputs(1399));
    layer3_outputs(18) <= layer2_outputs(3772);
    layer3_outputs(19) <= layer2_outputs(2532);
    layer3_outputs(20) <= (layer2_outputs(3713)) xor (layer2_outputs(1852));
    layer3_outputs(21) <= layer2_outputs(387);
    layer3_outputs(22) <= layer2_outputs(4335);
    layer3_outputs(23) <= not(layer2_outputs(2826));
    layer3_outputs(24) <= (layer2_outputs(445)) and not (layer2_outputs(684));
    layer3_outputs(25) <= (layer2_outputs(2999)) and not (layer2_outputs(572));
    layer3_outputs(26) <= '0';
    layer3_outputs(27) <= '0';
    layer3_outputs(28) <= not(layer2_outputs(3037));
    layer3_outputs(29) <= not((layer2_outputs(956)) and (layer2_outputs(3577)));
    layer3_outputs(30) <= layer2_outputs(3897);
    layer3_outputs(31) <= layer2_outputs(5002);
    layer3_outputs(32) <= '0';
    layer3_outputs(33) <= '1';
    layer3_outputs(34) <= not(layer2_outputs(172)) or (layer2_outputs(4462));
    layer3_outputs(35) <= '0';
    layer3_outputs(36) <= '1';
    layer3_outputs(37) <= layer2_outputs(309);
    layer3_outputs(38) <= (layer2_outputs(3786)) and not (layer2_outputs(1291));
    layer3_outputs(39) <= not(layer2_outputs(343));
    layer3_outputs(40) <= (layer2_outputs(4109)) and (layer2_outputs(2334));
    layer3_outputs(41) <= '0';
    layer3_outputs(42) <= not(layer2_outputs(3114));
    layer3_outputs(43) <= not(layer2_outputs(1096));
    layer3_outputs(44) <= '0';
    layer3_outputs(45) <= layer2_outputs(1907);
    layer3_outputs(46) <= (layer2_outputs(3335)) or (layer2_outputs(3799));
    layer3_outputs(47) <= '1';
    layer3_outputs(48) <= '1';
    layer3_outputs(49) <= (layer2_outputs(1439)) and (layer2_outputs(2703));
    layer3_outputs(50) <= (layer2_outputs(2877)) or (layer2_outputs(3191));
    layer3_outputs(51) <= '1';
    layer3_outputs(52) <= layer2_outputs(4016);
    layer3_outputs(53) <= layer2_outputs(2083);
    layer3_outputs(54) <= (layer2_outputs(1394)) and not (layer2_outputs(4967));
    layer3_outputs(55) <= not(layer2_outputs(2083)) or (layer2_outputs(141));
    layer3_outputs(56) <= not(layer2_outputs(3996)) or (layer2_outputs(647));
    layer3_outputs(57) <= (layer2_outputs(2763)) or (layer2_outputs(4821));
    layer3_outputs(58) <= not((layer2_outputs(2479)) and (layer2_outputs(3436)));
    layer3_outputs(59) <= layer2_outputs(557);
    layer3_outputs(60) <= not(layer2_outputs(2482)) or (layer2_outputs(1229));
    layer3_outputs(61) <= not((layer2_outputs(3726)) xor (layer2_outputs(4553)));
    layer3_outputs(62) <= '1';
    layer3_outputs(63) <= '0';
    layer3_outputs(64) <= '0';
    layer3_outputs(65) <= not(layer2_outputs(2920)) or (layer2_outputs(3366));
    layer3_outputs(66) <= layer2_outputs(550);
    layer3_outputs(67) <= (layer2_outputs(3943)) or (layer2_outputs(3427));
    layer3_outputs(68) <= (layer2_outputs(942)) or (layer2_outputs(1038));
    layer3_outputs(69) <= layer2_outputs(960);
    layer3_outputs(70) <= '1';
    layer3_outputs(71) <= (layer2_outputs(2745)) and (layer2_outputs(1261));
    layer3_outputs(72) <= '0';
    layer3_outputs(73) <= not((layer2_outputs(4924)) and (layer2_outputs(1500)));
    layer3_outputs(74) <= (layer2_outputs(486)) and not (layer2_outputs(2975));
    layer3_outputs(75) <= not(layer2_outputs(3530));
    layer3_outputs(76) <= layer2_outputs(3298);
    layer3_outputs(77) <= not(layer2_outputs(3218)) or (layer2_outputs(3416));
    layer3_outputs(78) <= layer2_outputs(3138);
    layer3_outputs(79) <= (layer2_outputs(888)) and not (layer2_outputs(2944));
    layer3_outputs(80) <= not(layer2_outputs(2628)) or (layer2_outputs(4816));
    layer3_outputs(81) <= not((layer2_outputs(2499)) and (layer2_outputs(3399)));
    layer3_outputs(82) <= (layer2_outputs(3508)) and not (layer2_outputs(1508));
    layer3_outputs(83) <= (layer2_outputs(1898)) and (layer2_outputs(1841));
    layer3_outputs(84) <= layer2_outputs(2670);
    layer3_outputs(85) <= not((layer2_outputs(4395)) or (layer2_outputs(2666)));
    layer3_outputs(86) <= not(layer2_outputs(668)) or (layer2_outputs(1837));
    layer3_outputs(87) <= (layer2_outputs(36)) and not (layer2_outputs(4838));
    layer3_outputs(88) <= '1';
    layer3_outputs(89) <= '1';
    layer3_outputs(90) <= '1';
    layer3_outputs(91) <= (layer2_outputs(4706)) and (layer2_outputs(3081));
    layer3_outputs(92) <= not(layer2_outputs(3487));
    layer3_outputs(93) <= '1';
    layer3_outputs(94) <= '1';
    layer3_outputs(95) <= not(layer2_outputs(345));
    layer3_outputs(96) <= layer2_outputs(4234);
    layer3_outputs(97) <= not((layer2_outputs(836)) and (layer2_outputs(2134)));
    layer3_outputs(98) <= not((layer2_outputs(2058)) and (layer2_outputs(623)));
    layer3_outputs(99) <= '0';
    layer3_outputs(100) <= (layer2_outputs(3339)) and not (layer2_outputs(2567));
    layer3_outputs(101) <= (layer2_outputs(1687)) or (layer2_outputs(4160));
    layer3_outputs(102) <= '1';
    layer3_outputs(103) <= (layer2_outputs(1275)) and not (layer2_outputs(637));
    layer3_outputs(104) <= not((layer2_outputs(2430)) or (layer2_outputs(1692)));
    layer3_outputs(105) <= '0';
    layer3_outputs(106) <= (layer2_outputs(1902)) and not (layer2_outputs(4467));
    layer3_outputs(107) <= (layer2_outputs(3541)) and not (layer2_outputs(3831));
    layer3_outputs(108) <= not((layer2_outputs(4255)) or (layer2_outputs(4354)));
    layer3_outputs(109) <= (layer2_outputs(486)) and not (layer2_outputs(75));
    layer3_outputs(110) <= layer2_outputs(1050);
    layer3_outputs(111) <= layer2_outputs(4254);
    layer3_outputs(112) <= (layer2_outputs(3254)) and (layer2_outputs(4214));
    layer3_outputs(113) <= (layer2_outputs(4311)) and not (layer2_outputs(4394));
    layer3_outputs(114) <= not((layer2_outputs(955)) or (layer2_outputs(921)));
    layer3_outputs(115) <= not(layer2_outputs(2805)) or (layer2_outputs(2441));
    layer3_outputs(116) <= not(layer2_outputs(973));
    layer3_outputs(117) <= (layer2_outputs(851)) and (layer2_outputs(1089));
    layer3_outputs(118) <= '1';
    layer3_outputs(119) <= not(layer2_outputs(1464)) or (layer2_outputs(348));
    layer3_outputs(120) <= '1';
    layer3_outputs(121) <= '0';
    layer3_outputs(122) <= (layer2_outputs(1508)) or (layer2_outputs(1879));
    layer3_outputs(123) <= layer2_outputs(3580);
    layer3_outputs(124) <= '0';
    layer3_outputs(125) <= not((layer2_outputs(3578)) or (layer2_outputs(1567)));
    layer3_outputs(126) <= '0';
    layer3_outputs(127) <= not((layer2_outputs(1580)) and (layer2_outputs(1871)));
    layer3_outputs(128) <= '0';
    layer3_outputs(129) <= layer2_outputs(1769);
    layer3_outputs(130) <= '0';
    layer3_outputs(131) <= not(layer2_outputs(3056)) or (layer2_outputs(287));
    layer3_outputs(132) <= '0';
    layer3_outputs(133) <= '1';
    layer3_outputs(134) <= not(layer2_outputs(3069)) or (layer2_outputs(2215));
    layer3_outputs(135) <= (layer2_outputs(3836)) and not (layer2_outputs(3474));
    layer3_outputs(136) <= '0';
    layer3_outputs(137) <= (layer2_outputs(3973)) and not (layer2_outputs(3930));
    layer3_outputs(138) <= (layer2_outputs(2832)) and (layer2_outputs(3756));
    layer3_outputs(139) <= (layer2_outputs(163)) and (layer2_outputs(563));
    layer3_outputs(140) <= not(layer2_outputs(4597));
    layer3_outputs(141) <= '1';
    layer3_outputs(142) <= not(layer2_outputs(2912));
    layer3_outputs(143) <= (layer2_outputs(3267)) and (layer2_outputs(207));
    layer3_outputs(144) <= not(layer2_outputs(4793));
    layer3_outputs(145) <= (layer2_outputs(4519)) or (layer2_outputs(2469));
    layer3_outputs(146) <= (layer2_outputs(3832)) and not (layer2_outputs(1813));
    layer3_outputs(147) <= '1';
    layer3_outputs(148) <= layer2_outputs(249);
    layer3_outputs(149) <= layer2_outputs(1132);
    layer3_outputs(150) <= not(layer2_outputs(1877));
    layer3_outputs(151) <= layer2_outputs(2517);
    layer3_outputs(152) <= '0';
    layer3_outputs(153) <= not((layer2_outputs(2181)) or (layer2_outputs(3452)));
    layer3_outputs(154) <= not((layer2_outputs(5064)) or (layer2_outputs(4899)));
    layer3_outputs(155) <= '0';
    layer3_outputs(156) <= not(layer2_outputs(1793));
    layer3_outputs(157) <= (layer2_outputs(2812)) and not (layer2_outputs(588));
    layer3_outputs(158) <= '1';
    layer3_outputs(159) <= (layer2_outputs(5018)) and (layer2_outputs(4590));
    layer3_outputs(160) <= layer2_outputs(2189);
    layer3_outputs(161) <= not(layer2_outputs(1492));
    layer3_outputs(162) <= (layer2_outputs(1231)) and not (layer2_outputs(3928));
    layer3_outputs(163) <= not(layer2_outputs(3753)) or (layer2_outputs(160));
    layer3_outputs(164) <= layer2_outputs(373);
    layer3_outputs(165) <= (layer2_outputs(4047)) or (layer2_outputs(3856));
    layer3_outputs(166) <= (layer2_outputs(4221)) and (layer2_outputs(603));
    layer3_outputs(167) <= not(layer2_outputs(4904));
    layer3_outputs(168) <= (layer2_outputs(91)) and (layer2_outputs(3406));
    layer3_outputs(169) <= (layer2_outputs(5)) or (layer2_outputs(2544));
    layer3_outputs(170) <= layer2_outputs(1661);
    layer3_outputs(171) <= '1';
    layer3_outputs(172) <= '1';
    layer3_outputs(173) <= not((layer2_outputs(4942)) and (layer2_outputs(4065)));
    layer3_outputs(174) <= (layer2_outputs(2843)) and not (layer2_outputs(707));
    layer3_outputs(175) <= layer2_outputs(3432);
    layer3_outputs(176) <= not(layer2_outputs(1671));
    layer3_outputs(177) <= not(layer2_outputs(4643)) or (layer2_outputs(2122));
    layer3_outputs(178) <= layer2_outputs(3627);
    layer3_outputs(179) <= '1';
    layer3_outputs(180) <= not((layer2_outputs(4866)) or (layer2_outputs(5009)));
    layer3_outputs(181) <= not((layer2_outputs(769)) or (layer2_outputs(2020)));
    layer3_outputs(182) <= '0';
    layer3_outputs(183) <= not(layer2_outputs(2988)) or (layer2_outputs(630));
    layer3_outputs(184) <= not((layer2_outputs(4912)) and (layer2_outputs(3564)));
    layer3_outputs(185) <= (layer2_outputs(1220)) and (layer2_outputs(3240));
    layer3_outputs(186) <= layer2_outputs(3253);
    layer3_outputs(187) <= not(layer2_outputs(1216));
    layer3_outputs(188) <= not(layer2_outputs(4766));
    layer3_outputs(189) <= layer2_outputs(3784);
    layer3_outputs(190) <= not(layer2_outputs(4780)) or (layer2_outputs(1215));
    layer3_outputs(191) <= (layer2_outputs(4974)) and (layer2_outputs(2850));
    layer3_outputs(192) <= '1';
    layer3_outputs(193) <= layer2_outputs(4731);
    layer3_outputs(194) <= not((layer2_outputs(4713)) and (layer2_outputs(2798)));
    layer3_outputs(195) <= (layer2_outputs(415)) and (layer2_outputs(1340));
    layer3_outputs(196) <= (layer2_outputs(105)) and not (layer2_outputs(4619));
    layer3_outputs(197) <= not(layer2_outputs(2007)) or (layer2_outputs(510));
    layer3_outputs(198) <= (layer2_outputs(1956)) and not (layer2_outputs(2587));
    layer3_outputs(199) <= '1';
    layer3_outputs(200) <= not(layer2_outputs(1050)) or (layer2_outputs(2350));
    layer3_outputs(201) <= layer2_outputs(3150);
    layer3_outputs(202) <= not(layer2_outputs(3132)) or (layer2_outputs(5021));
    layer3_outputs(203) <= '1';
    layer3_outputs(204) <= '0';
    layer3_outputs(205) <= not(layer2_outputs(743));
    layer3_outputs(206) <= '1';
    layer3_outputs(207) <= (layer2_outputs(4786)) and not (layer2_outputs(886));
    layer3_outputs(208) <= not((layer2_outputs(2937)) or (layer2_outputs(1913)));
    layer3_outputs(209) <= '1';
    layer3_outputs(210) <= '0';
    layer3_outputs(211) <= layer2_outputs(589);
    layer3_outputs(212) <= '0';
    layer3_outputs(213) <= layer2_outputs(120);
    layer3_outputs(214) <= (layer2_outputs(2243)) and not (layer2_outputs(3734));
    layer3_outputs(215) <= not((layer2_outputs(4681)) and (layer2_outputs(3733)));
    layer3_outputs(216) <= layer2_outputs(3016);
    layer3_outputs(217) <= '0';
    layer3_outputs(218) <= '1';
    layer3_outputs(219) <= '1';
    layer3_outputs(220) <= layer2_outputs(3215);
    layer3_outputs(221) <= not((layer2_outputs(1310)) or (layer2_outputs(878)));
    layer3_outputs(222) <= '1';
    layer3_outputs(223) <= not((layer2_outputs(4126)) or (layer2_outputs(1434)));
    layer3_outputs(224) <= not(layer2_outputs(3059));
    layer3_outputs(225) <= not(layer2_outputs(4351));
    layer3_outputs(226) <= '1';
    layer3_outputs(227) <= not(layer2_outputs(5050));
    layer3_outputs(228) <= layer2_outputs(2359);
    layer3_outputs(229) <= layer2_outputs(1169);
    layer3_outputs(230) <= not((layer2_outputs(4671)) or (layer2_outputs(828)));
    layer3_outputs(231) <= (layer2_outputs(455)) and not (layer2_outputs(718));
    layer3_outputs(232) <= '1';
    layer3_outputs(233) <= not(layer2_outputs(2093));
    layer3_outputs(234) <= layer2_outputs(3134);
    layer3_outputs(235) <= '0';
    layer3_outputs(236) <= (layer2_outputs(2891)) and (layer2_outputs(1966));
    layer3_outputs(237) <= not(layer2_outputs(4501)) or (layer2_outputs(1074));
    layer3_outputs(238) <= not((layer2_outputs(260)) and (layer2_outputs(3672)));
    layer3_outputs(239) <= not(layer2_outputs(658)) or (layer2_outputs(3291));
    layer3_outputs(240) <= not(layer2_outputs(835)) or (layer2_outputs(829));
    layer3_outputs(241) <= '1';
    layer3_outputs(242) <= '0';
    layer3_outputs(243) <= not(layer2_outputs(177)) or (layer2_outputs(4424));
    layer3_outputs(244) <= not(layer2_outputs(681)) or (layer2_outputs(1347));
    layer3_outputs(245) <= '0';
    layer3_outputs(246) <= '1';
    layer3_outputs(247) <= (layer2_outputs(1781)) and not (layer2_outputs(4072));
    layer3_outputs(248) <= (layer2_outputs(2824)) and (layer2_outputs(3092));
    layer3_outputs(249) <= (layer2_outputs(3816)) and not (layer2_outputs(3203));
    layer3_outputs(250) <= not((layer2_outputs(4454)) or (layer2_outputs(1072)));
    layer3_outputs(251) <= (layer2_outputs(1324)) and not (layer2_outputs(2029));
    layer3_outputs(252) <= (layer2_outputs(1622)) and not (layer2_outputs(4793));
    layer3_outputs(253) <= not(layer2_outputs(2355));
    layer3_outputs(254) <= not((layer2_outputs(4596)) or (layer2_outputs(3111)));
    layer3_outputs(255) <= '0';
    layer3_outputs(256) <= (layer2_outputs(3315)) or (layer2_outputs(2032));
    layer3_outputs(257) <= not((layer2_outputs(3277)) and (layer2_outputs(3272)));
    layer3_outputs(258) <= '0';
    layer3_outputs(259) <= (layer2_outputs(1419)) and not (layer2_outputs(3555));
    layer3_outputs(260) <= (layer2_outputs(2198)) and (layer2_outputs(2374));
    layer3_outputs(261) <= layer2_outputs(57);
    layer3_outputs(262) <= not(layer2_outputs(3217)) or (layer2_outputs(2199));
    layer3_outputs(263) <= '0';
    layer3_outputs(264) <= (layer2_outputs(2411)) xor (layer2_outputs(3612));
    layer3_outputs(265) <= '1';
    layer3_outputs(266) <= '1';
    layer3_outputs(267) <= (layer2_outputs(484)) and not (layer2_outputs(13));
    layer3_outputs(268) <= layer2_outputs(2893);
    layer3_outputs(269) <= (layer2_outputs(4691)) and not (layer2_outputs(2216));
    layer3_outputs(270) <= not(layer2_outputs(1700)) or (layer2_outputs(3765));
    layer3_outputs(271) <= layer2_outputs(2211);
    layer3_outputs(272) <= not(layer2_outputs(342)) or (layer2_outputs(1606));
    layer3_outputs(273) <= not((layer2_outputs(3608)) and (layer2_outputs(4293)));
    layer3_outputs(274) <= (layer2_outputs(5065)) and (layer2_outputs(2657));
    layer3_outputs(275) <= (layer2_outputs(2845)) and not (layer2_outputs(1914));
    layer3_outputs(276) <= not(layer2_outputs(2892)) or (layer2_outputs(352));
    layer3_outputs(277) <= '1';
    layer3_outputs(278) <= layer2_outputs(2059);
    layer3_outputs(279) <= not((layer2_outputs(1935)) xor (layer2_outputs(4944)));
    layer3_outputs(280) <= not(layer2_outputs(794));
    layer3_outputs(281) <= not((layer2_outputs(1490)) and (layer2_outputs(2958)));
    layer3_outputs(282) <= not(layer2_outputs(2286));
    layer3_outputs(283) <= '1';
    layer3_outputs(284) <= (layer2_outputs(1406)) and not (layer2_outputs(4094));
    layer3_outputs(285) <= not((layer2_outputs(1649)) or (layer2_outputs(1912)));
    layer3_outputs(286) <= not(layer2_outputs(4142)) or (layer2_outputs(885));
    layer3_outputs(287) <= not(layer2_outputs(655));
    layer3_outputs(288) <= (layer2_outputs(3873)) or (layer2_outputs(1740));
    layer3_outputs(289) <= '0';
    layer3_outputs(290) <= '0';
    layer3_outputs(291) <= not(layer2_outputs(2841)) or (layer2_outputs(203));
    layer3_outputs(292) <= not(layer2_outputs(4444)) or (layer2_outputs(4694));
    layer3_outputs(293) <= not((layer2_outputs(3523)) and (layer2_outputs(3870)));
    layer3_outputs(294) <= layer2_outputs(3121);
    layer3_outputs(295) <= not(layer2_outputs(186)) or (layer2_outputs(2650));
    layer3_outputs(296) <= not(layer2_outputs(4261));
    layer3_outputs(297) <= not(layer2_outputs(502)) or (layer2_outputs(4258));
    layer3_outputs(298) <= not((layer2_outputs(3239)) xor (layer2_outputs(4556)));
    layer3_outputs(299) <= not(layer2_outputs(1376)) or (layer2_outputs(1323));
    layer3_outputs(300) <= '1';
    layer3_outputs(301) <= not(layer2_outputs(1836)) or (layer2_outputs(2754));
    layer3_outputs(302) <= not((layer2_outputs(1491)) or (layer2_outputs(3091)));
    layer3_outputs(303) <= (layer2_outputs(1812)) or (layer2_outputs(1252));
    layer3_outputs(304) <= '1';
    layer3_outputs(305) <= not(layer2_outputs(570)) or (layer2_outputs(2519));
    layer3_outputs(306) <= not((layer2_outputs(3702)) and (layer2_outputs(250)));
    layer3_outputs(307) <= (layer2_outputs(2163)) and not (layer2_outputs(3459));
    layer3_outputs(308) <= (layer2_outputs(813)) and not (layer2_outputs(2805));
    layer3_outputs(309) <= not((layer2_outputs(4748)) and (layer2_outputs(2874)));
    layer3_outputs(310) <= (layer2_outputs(1492)) and not (layer2_outputs(811));
    layer3_outputs(311) <= '1';
    layer3_outputs(312) <= (layer2_outputs(588)) and not (layer2_outputs(1079));
    layer3_outputs(313) <= layer2_outputs(1337);
    layer3_outputs(314) <= (layer2_outputs(2016)) and not (layer2_outputs(3125));
    layer3_outputs(315) <= (layer2_outputs(1526)) and not (layer2_outputs(3255));
    layer3_outputs(316) <= (layer2_outputs(1069)) or (layer2_outputs(4405));
    layer3_outputs(317) <= not(layer2_outputs(2218)) or (layer2_outputs(2421));
    layer3_outputs(318) <= not(layer2_outputs(4587)) or (layer2_outputs(2940));
    layer3_outputs(319) <= not(layer2_outputs(3382));
    layer3_outputs(320) <= not(layer2_outputs(1415));
    layer3_outputs(321) <= '0';
    layer3_outputs(322) <= '0';
    layer3_outputs(323) <= (layer2_outputs(3539)) xor (layer2_outputs(1139));
    layer3_outputs(324) <= not(layer2_outputs(1159));
    layer3_outputs(325) <= not(layer2_outputs(4848));
    layer3_outputs(326) <= (layer2_outputs(2392)) and not (layer2_outputs(223));
    layer3_outputs(327) <= not((layer2_outputs(3539)) or (layer2_outputs(1201)));
    layer3_outputs(328) <= not(layer2_outputs(4747));
    layer3_outputs(329) <= (layer2_outputs(3939)) and not (layer2_outputs(2754));
    layer3_outputs(330) <= not((layer2_outputs(3468)) and (layer2_outputs(266)));
    layer3_outputs(331) <= '1';
    layer3_outputs(332) <= not(layer2_outputs(126)) or (layer2_outputs(476));
    layer3_outputs(333) <= '1';
    layer3_outputs(334) <= not((layer2_outputs(2750)) or (layer2_outputs(4992)));
    layer3_outputs(335) <= not(layer2_outputs(2169)) or (layer2_outputs(4562));
    layer3_outputs(336) <= layer2_outputs(3842);
    layer3_outputs(337) <= not(layer2_outputs(3235)) or (layer2_outputs(3043));
    layer3_outputs(338) <= (layer2_outputs(4136)) or (layer2_outputs(3420));
    layer3_outputs(339) <= layer2_outputs(2072);
    layer3_outputs(340) <= (layer2_outputs(3707)) and not (layer2_outputs(940));
    layer3_outputs(341) <= layer2_outputs(2581);
    layer3_outputs(342) <= (layer2_outputs(3797)) and (layer2_outputs(4499));
    layer3_outputs(343) <= (layer2_outputs(1607)) and not (layer2_outputs(3412));
    layer3_outputs(344) <= not(layer2_outputs(1610)) or (layer2_outputs(2335));
    layer3_outputs(345) <= not(layer2_outputs(674)) or (layer2_outputs(699));
    layer3_outputs(346) <= layer2_outputs(1243);
    layer3_outputs(347) <= layer2_outputs(3725);
    layer3_outputs(348) <= not(layer2_outputs(1668));
    layer3_outputs(349) <= not((layer2_outputs(211)) and (layer2_outputs(268)));
    layer3_outputs(350) <= not(layer2_outputs(3979));
    layer3_outputs(351) <= not(layer2_outputs(5049)) or (layer2_outputs(123));
    layer3_outputs(352) <= not(layer2_outputs(3397)) or (layer2_outputs(3628));
    layer3_outputs(353) <= (layer2_outputs(836)) or (layer2_outputs(2507));
    layer3_outputs(354) <= '1';
    layer3_outputs(355) <= not(layer2_outputs(4175));
    layer3_outputs(356) <= not(layer2_outputs(4727)) or (layer2_outputs(1078));
    layer3_outputs(357) <= not(layer2_outputs(1698)) or (layer2_outputs(2953));
    layer3_outputs(358) <= layer2_outputs(2718);
    layer3_outputs(359) <= '1';
    layer3_outputs(360) <= (layer2_outputs(606)) and not (layer2_outputs(114));
    layer3_outputs(361) <= '1';
    layer3_outputs(362) <= not(layer2_outputs(894));
    layer3_outputs(363) <= '1';
    layer3_outputs(364) <= not(layer2_outputs(2074));
    layer3_outputs(365) <= (layer2_outputs(5082)) and (layer2_outputs(2436));
    layer3_outputs(366) <= not(layer2_outputs(742));
    layer3_outputs(367) <= (layer2_outputs(3648)) or (layer2_outputs(4972));
    layer3_outputs(368) <= '0';
    layer3_outputs(369) <= (layer2_outputs(1664)) and not (layer2_outputs(2561));
    layer3_outputs(370) <= not((layer2_outputs(3919)) xor (layer2_outputs(1667)));
    layer3_outputs(371) <= not(layer2_outputs(31)) or (layer2_outputs(5079));
    layer3_outputs(372) <= layer2_outputs(513);
    layer3_outputs(373) <= (layer2_outputs(3460)) or (layer2_outputs(442));
    layer3_outputs(374) <= not((layer2_outputs(1649)) or (layer2_outputs(460)));
    layer3_outputs(375) <= not((layer2_outputs(80)) or (layer2_outputs(850)));
    layer3_outputs(376) <= layer2_outputs(4145);
    layer3_outputs(377) <= (layer2_outputs(4255)) and not (layer2_outputs(511));
    layer3_outputs(378) <= not(layer2_outputs(832));
    layer3_outputs(379) <= (layer2_outputs(2857)) and not (layer2_outputs(3426));
    layer3_outputs(380) <= (layer2_outputs(1484)) and not (layer2_outputs(3133));
    layer3_outputs(381) <= '0';
    layer3_outputs(382) <= not((layer2_outputs(1525)) or (layer2_outputs(3110)));
    layer3_outputs(383) <= '1';
    layer3_outputs(384) <= (layer2_outputs(4508)) and not (layer2_outputs(487));
    layer3_outputs(385) <= not(layer2_outputs(2994));
    layer3_outputs(386) <= '0';
    layer3_outputs(387) <= not((layer2_outputs(5011)) and (layer2_outputs(4081)));
    layer3_outputs(388) <= '1';
    layer3_outputs(389) <= '1';
    layer3_outputs(390) <= layer2_outputs(587);
    layer3_outputs(391) <= (layer2_outputs(3634)) and not (layer2_outputs(1463));
    layer3_outputs(392) <= layer2_outputs(4133);
    layer3_outputs(393) <= '0';
    layer3_outputs(394) <= not(layer2_outputs(3616)) or (layer2_outputs(602));
    layer3_outputs(395) <= not(layer2_outputs(3255)) or (layer2_outputs(2046));
    layer3_outputs(396) <= not((layer2_outputs(2033)) or (layer2_outputs(115)));
    layer3_outputs(397) <= '1';
    layer3_outputs(398) <= not((layer2_outputs(4611)) or (layer2_outputs(1246)));
    layer3_outputs(399) <= not(layer2_outputs(4953));
    layer3_outputs(400) <= not(layer2_outputs(2382)) or (layer2_outputs(2013));
    layer3_outputs(401) <= not((layer2_outputs(526)) or (layer2_outputs(179)));
    layer3_outputs(402) <= '0';
    layer3_outputs(403) <= (layer2_outputs(1123)) and (layer2_outputs(1008));
    layer3_outputs(404) <= not(layer2_outputs(4880)) or (layer2_outputs(4592));
    layer3_outputs(405) <= (layer2_outputs(4327)) or (layer2_outputs(231));
    layer3_outputs(406) <= (layer2_outputs(1754)) and not (layer2_outputs(3014));
    layer3_outputs(407) <= not(layer2_outputs(2505));
    layer3_outputs(408) <= layer2_outputs(3637);
    layer3_outputs(409) <= layer2_outputs(2141);
    layer3_outputs(410) <= (layer2_outputs(1380)) and (layer2_outputs(4684));
    layer3_outputs(411) <= not(layer2_outputs(567));
    layer3_outputs(412) <= not((layer2_outputs(1619)) and (layer2_outputs(4170)));
    layer3_outputs(413) <= not((layer2_outputs(4360)) or (layer2_outputs(4750)));
    layer3_outputs(414) <= '1';
    layer3_outputs(415) <= layer2_outputs(204);
    layer3_outputs(416) <= (layer2_outputs(2531)) or (layer2_outputs(316));
    layer3_outputs(417) <= (layer2_outputs(3602)) and not (layer2_outputs(59));
    layer3_outputs(418) <= not(layer2_outputs(1759)) or (layer2_outputs(1584));
    layer3_outputs(419) <= (layer2_outputs(2064)) and not (layer2_outputs(854));
    layer3_outputs(420) <= not(layer2_outputs(169)) or (layer2_outputs(4888));
    layer3_outputs(421) <= layer2_outputs(5054);
    layer3_outputs(422) <= (layer2_outputs(4161)) and not (layer2_outputs(4445));
    layer3_outputs(423) <= '1';
    layer3_outputs(424) <= not((layer2_outputs(2834)) or (layer2_outputs(941)));
    layer3_outputs(425) <= (layer2_outputs(1599)) and (layer2_outputs(3225));
    layer3_outputs(426) <= not(layer2_outputs(1635));
    layer3_outputs(427) <= layer2_outputs(1307);
    layer3_outputs(428) <= '1';
    layer3_outputs(429) <= not(layer2_outputs(3100)) or (layer2_outputs(798));
    layer3_outputs(430) <= not(layer2_outputs(1012)) or (layer2_outputs(3754));
    layer3_outputs(431) <= layer2_outputs(1790);
    layer3_outputs(432) <= '0';
    layer3_outputs(433) <= '1';
    layer3_outputs(434) <= not(layer2_outputs(1735));
    layer3_outputs(435) <= layer2_outputs(958);
    layer3_outputs(436) <= (layer2_outputs(355)) and (layer2_outputs(4920));
    layer3_outputs(437) <= (layer2_outputs(4919)) and not (layer2_outputs(3321));
    layer3_outputs(438) <= not((layer2_outputs(4135)) and (layer2_outputs(249)));
    layer3_outputs(439) <= layer2_outputs(2561);
    layer3_outputs(440) <= (layer2_outputs(1186)) and (layer2_outputs(4647));
    layer3_outputs(441) <= (layer2_outputs(2734)) and (layer2_outputs(999));
    layer3_outputs(442) <= (layer2_outputs(399)) and not (layer2_outputs(3701));
    layer3_outputs(443) <= layer2_outputs(4248);
    layer3_outputs(444) <= not(layer2_outputs(469)) or (layer2_outputs(817));
    layer3_outputs(445) <= not(layer2_outputs(1930)) or (layer2_outputs(2553));
    layer3_outputs(446) <= (layer2_outputs(4410)) or (layer2_outputs(4083));
    layer3_outputs(447) <= (layer2_outputs(1936)) and (layer2_outputs(2595));
    layer3_outputs(448) <= (layer2_outputs(384)) and not (layer2_outputs(1283));
    layer3_outputs(449) <= (layer2_outputs(495)) or (layer2_outputs(289));
    layer3_outputs(450) <= not((layer2_outputs(2728)) or (layer2_outputs(3185)));
    layer3_outputs(451) <= not((layer2_outputs(3988)) or (layer2_outputs(46)));
    layer3_outputs(452) <= '0';
    layer3_outputs(453) <= not((layer2_outputs(2761)) or (layer2_outputs(4522)));
    layer3_outputs(454) <= (layer2_outputs(1396)) and not (layer2_outputs(3958));
    layer3_outputs(455) <= not(layer2_outputs(2533));
    layer3_outputs(456) <= not(layer2_outputs(354));
    layer3_outputs(457) <= (layer2_outputs(1947)) and not (layer2_outputs(1592));
    layer3_outputs(458) <= layer2_outputs(5039);
    layer3_outputs(459) <= (layer2_outputs(2848)) or (layer2_outputs(4093));
    layer3_outputs(460) <= layer2_outputs(3875);
    layer3_outputs(461) <= layer2_outputs(2834);
    layer3_outputs(462) <= layer2_outputs(2306);
    layer3_outputs(463) <= (layer2_outputs(474)) and not (layer2_outputs(1385));
    layer3_outputs(464) <= not(layer2_outputs(2803)) or (layer2_outputs(4437));
    layer3_outputs(465) <= not(layer2_outputs(4536));
    layer3_outputs(466) <= '1';
    layer3_outputs(467) <= (layer2_outputs(3411)) and not (layer2_outputs(2324));
    layer3_outputs(468) <= layer2_outputs(1104);
    layer3_outputs(469) <= (layer2_outputs(2360)) and not (layer2_outputs(4778));
    layer3_outputs(470) <= (layer2_outputs(1498)) or (layer2_outputs(3336));
    layer3_outputs(471) <= not((layer2_outputs(2038)) or (layer2_outputs(5036)));
    layer3_outputs(472) <= not(layer2_outputs(1733));
    layer3_outputs(473) <= not((layer2_outputs(4097)) or (layer2_outputs(5031)));
    layer3_outputs(474) <= (layer2_outputs(2453)) and not (layer2_outputs(4264));
    layer3_outputs(475) <= layer2_outputs(3657);
    layer3_outputs(476) <= (layer2_outputs(2241)) and not (layer2_outputs(3457));
    layer3_outputs(477) <= layer2_outputs(4997);
    layer3_outputs(478) <= (layer2_outputs(4978)) and (layer2_outputs(3966));
    layer3_outputs(479) <= (layer2_outputs(662)) and not (layer2_outputs(2516));
    layer3_outputs(480) <= (layer2_outputs(3295)) and not (layer2_outputs(1460));
    layer3_outputs(481) <= not(layer2_outputs(3056)) or (layer2_outputs(2960));
    layer3_outputs(482) <= '0';
    layer3_outputs(483) <= not(layer2_outputs(795));
    layer3_outputs(484) <= '1';
    layer3_outputs(485) <= '0';
    layer3_outputs(486) <= (layer2_outputs(2904)) or (layer2_outputs(3837));
    layer3_outputs(487) <= layer2_outputs(2100);
    layer3_outputs(488) <= (layer2_outputs(1877)) and not (layer2_outputs(5066));
    layer3_outputs(489) <= not(layer2_outputs(1656)) or (layer2_outputs(2254));
    layer3_outputs(490) <= (layer2_outputs(951)) and not (layer2_outputs(3848));
    layer3_outputs(491) <= not(layer2_outputs(2193));
    layer3_outputs(492) <= '0';
    layer3_outputs(493) <= '1';
    layer3_outputs(494) <= '1';
    layer3_outputs(495) <= '1';
    layer3_outputs(496) <= (layer2_outputs(4074)) and not (layer2_outputs(5044));
    layer3_outputs(497) <= not(layer2_outputs(1146));
    layer3_outputs(498) <= (layer2_outputs(3489)) and (layer2_outputs(1495));
    layer3_outputs(499) <= (layer2_outputs(2878)) or (layer2_outputs(1910));
    layer3_outputs(500) <= (layer2_outputs(4853)) and not (layer2_outputs(1653));
    layer3_outputs(501) <= not(layer2_outputs(1696)) or (layer2_outputs(2913));
    layer3_outputs(502) <= layer2_outputs(4601);
    layer3_outputs(503) <= not(layer2_outputs(3767));
    layer3_outputs(504) <= layer2_outputs(2949);
    layer3_outputs(505) <= (layer2_outputs(2747)) xor (layer2_outputs(4367));
    layer3_outputs(506) <= not(layer2_outputs(467)) or (layer2_outputs(273));
    layer3_outputs(507) <= layer2_outputs(4224);
    layer3_outputs(508) <= not((layer2_outputs(4898)) or (layer2_outputs(3420)));
    layer3_outputs(509) <= not(layer2_outputs(4529)) or (layer2_outputs(3305));
    layer3_outputs(510) <= not(layer2_outputs(4709));
    layer3_outputs(511) <= not(layer2_outputs(2977)) or (layer2_outputs(4430));
    layer3_outputs(512) <= (layer2_outputs(3595)) xor (layer2_outputs(933));
    layer3_outputs(513) <= layer2_outputs(1727);
    layer3_outputs(514) <= '0';
    layer3_outputs(515) <= not((layer2_outputs(1755)) and (layer2_outputs(3615)));
    layer3_outputs(516) <= layer2_outputs(1873);
    layer3_outputs(517) <= '0';
    layer3_outputs(518) <= '1';
    layer3_outputs(519) <= (layer2_outputs(247)) and (layer2_outputs(3888));
    layer3_outputs(520) <= '1';
    layer3_outputs(521) <= not(layer2_outputs(1367));
    layer3_outputs(522) <= not(layer2_outputs(275));
    layer3_outputs(523) <= '0';
    layer3_outputs(524) <= not(layer2_outputs(4125)) or (layer2_outputs(4794));
    layer3_outputs(525) <= (layer2_outputs(1727)) and (layer2_outputs(2954));
    layer3_outputs(526) <= (layer2_outputs(1926)) and not (layer2_outputs(4703));
    layer3_outputs(527) <= not(layer2_outputs(3398)) or (layer2_outputs(1426));
    layer3_outputs(528) <= not(layer2_outputs(4756));
    layer3_outputs(529) <= '1';
    layer3_outputs(530) <= not(layer2_outputs(1874)) or (layer2_outputs(3836));
    layer3_outputs(531) <= (layer2_outputs(4976)) and not (layer2_outputs(4943));
    layer3_outputs(532) <= layer2_outputs(133);
    layer3_outputs(533) <= (layer2_outputs(2591)) and (layer2_outputs(561));
    layer3_outputs(534) <= '0';
    layer3_outputs(535) <= (layer2_outputs(635)) and not (layer2_outputs(3043));
    layer3_outputs(536) <= (layer2_outputs(1674)) or (layer2_outputs(3801));
    layer3_outputs(537) <= '1';
    layer3_outputs(538) <= (layer2_outputs(106)) or (layer2_outputs(4146));
    layer3_outputs(539) <= not(layer2_outputs(1903)) or (layer2_outputs(1946));
    layer3_outputs(540) <= '1';
    layer3_outputs(541) <= (layer2_outputs(1719)) xor (layer2_outputs(1229));
    layer3_outputs(542) <= not((layer2_outputs(3066)) and (layer2_outputs(3761)));
    layer3_outputs(543) <= (layer2_outputs(558)) and not (layer2_outputs(577));
    layer3_outputs(544) <= (layer2_outputs(850)) and not (layer2_outputs(1657));
    layer3_outputs(545) <= not(layer2_outputs(517)) or (layer2_outputs(3655));
    layer3_outputs(546) <= '0';
    layer3_outputs(547) <= not(layer2_outputs(522)) or (layer2_outputs(2763));
    layer3_outputs(548) <= not(layer2_outputs(1097));
    layer3_outputs(549) <= '1';
    layer3_outputs(550) <= (layer2_outputs(4158)) and (layer2_outputs(4946));
    layer3_outputs(551) <= layer2_outputs(4587);
    layer3_outputs(552) <= not(layer2_outputs(3685)) or (layer2_outputs(3385));
    layer3_outputs(553) <= not(layer2_outputs(4433)) or (layer2_outputs(3591));
    layer3_outputs(554) <= not((layer2_outputs(1250)) and (layer2_outputs(99)));
    layer3_outputs(555) <= '1';
    layer3_outputs(556) <= layer2_outputs(289);
    layer3_outputs(557) <= '0';
    layer3_outputs(558) <= (layer2_outputs(2005)) or (layer2_outputs(3509));
    layer3_outputs(559) <= '0';
    layer3_outputs(560) <= not((layer2_outputs(4082)) and (layer2_outputs(4084)));
    layer3_outputs(561) <= (layer2_outputs(2692)) and (layer2_outputs(4882));
    layer3_outputs(562) <= (layer2_outputs(4071)) and not (layer2_outputs(434));
    layer3_outputs(563) <= (layer2_outputs(2515)) and not (layer2_outputs(220));
    layer3_outputs(564) <= not((layer2_outputs(4060)) and (layer2_outputs(2159)));
    layer3_outputs(565) <= '0';
    layer3_outputs(566) <= (layer2_outputs(2221)) and not (layer2_outputs(3812));
    layer3_outputs(567) <= not(layer2_outputs(1394));
    layer3_outputs(568) <= (layer2_outputs(1712)) and not (layer2_outputs(2290));
    layer3_outputs(569) <= not(layer2_outputs(4522)) or (layer2_outputs(1548));
    layer3_outputs(570) <= not((layer2_outputs(4330)) or (layer2_outputs(4415)));
    layer3_outputs(571) <= not(layer2_outputs(3548)) or (layer2_outputs(4839));
    layer3_outputs(572) <= (layer2_outputs(3814)) and (layer2_outputs(1133));
    layer3_outputs(573) <= layer2_outputs(1773);
    layer3_outputs(574) <= (layer2_outputs(3796)) and not (layer2_outputs(287));
    layer3_outputs(575) <= (layer2_outputs(797)) and not (layer2_outputs(2616));
    layer3_outputs(576) <= not(layer2_outputs(545)) or (layer2_outputs(4027));
    layer3_outputs(577) <= '0';
    layer3_outputs(578) <= not((layer2_outputs(1266)) and (layer2_outputs(3946)));
    layer3_outputs(579) <= layer2_outputs(1678);
    layer3_outputs(580) <= (layer2_outputs(3634)) or (layer2_outputs(274));
    layer3_outputs(581) <= '0';
    layer3_outputs(582) <= not((layer2_outputs(3029)) xor (layer2_outputs(2296)));
    layer3_outputs(583) <= layer2_outputs(4887);
    layer3_outputs(584) <= (layer2_outputs(1235)) and not (layer2_outputs(1391));
    layer3_outputs(585) <= (layer2_outputs(787)) and (layer2_outputs(4314));
    layer3_outputs(586) <= not(layer2_outputs(5000));
    layer3_outputs(587) <= (layer2_outputs(1989)) and (layer2_outputs(357));
    layer3_outputs(588) <= (layer2_outputs(3112)) or (layer2_outputs(5056));
    layer3_outputs(589) <= (layer2_outputs(1705)) or (layer2_outputs(4667));
    layer3_outputs(590) <= not((layer2_outputs(1898)) and (layer2_outputs(2978)));
    layer3_outputs(591) <= '1';
    layer3_outputs(592) <= layer2_outputs(4184);
    layer3_outputs(593) <= not(layer2_outputs(2642));
    layer3_outputs(594) <= (layer2_outputs(129)) or (layer2_outputs(915));
    layer3_outputs(595) <= '1';
    layer3_outputs(596) <= (layer2_outputs(3790)) and not (layer2_outputs(1865));
    layer3_outputs(597) <= (layer2_outputs(3028)) and not (layer2_outputs(4418));
    layer3_outputs(598) <= (layer2_outputs(4990)) and not (layer2_outputs(2875));
    layer3_outputs(599) <= layer2_outputs(19);
    layer3_outputs(600) <= (layer2_outputs(1260)) and not (layer2_outputs(1832));
    layer3_outputs(601) <= '0';
    layer3_outputs(602) <= layer2_outputs(2011);
    layer3_outputs(603) <= (layer2_outputs(2094)) and not (layer2_outputs(4694));
    layer3_outputs(604) <= not(layer2_outputs(176));
    layer3_outputs(605) <= layer2_outputs(2138);
    layer3_outputs(606) <= layer2_outputs(3430);
    layer3_outputs(607) <= '1';
    layer3_outputs(608) <= not(layer2_outputs(2874)) or (layer2_outputs(2238));
    layer3_outputs(609) <= '1';
    layer3_outputs(610) <= (layer2_outputs(1509)) and (layer2_outputs(2979));
    layer3_outputs(611) <= (layer2_outputs(3503)) or (layer2_outputs(3921));
    layer3_outputs(612) <= layer2_outputs(4240);
    layer3_outputs(613) <= (layer2_outputs(2911)) and not (layer2_outputs(3138));
    layer3_outputs(614) <= '1';
    layer3_outputs(615) <= not(layer2_outputs(779));
    layer3_outputs(616) <= '0';
    layer3_outputs(617) <= '0';
    layer3_outputs(618) <= (layer2_outputs(2939)) and (layer2_outputs(5016));
    layer3_outputs(619) <= (layer2_outputs(738)) and not (layer2_outputs(4824));
    layer3_outputs(620) <= not((layer2_outputs(3869)) and (layer2_outputs(447)));
    layer3_outputs(621) <= not((layer2_outputs(1079)) xor (layer2_outputs(1926)));
    layer3_outputs(622) <= (layer2_outputs(4380)) or (layer2_outputs(3914));
    layer3_outputs(623) <= '0';
    layer3_outputs(624) <= (layer2_outputs(668)) and not (layer2_outputs(4300));
    layer3_outputs(625) <= not(layer2_outputs(561)) or (layer2_outputs(23));
    layer3_outputs(626) <= layer2_outputs(3149);
    layer3_outputs(627) <= (layer2_outputs(2293)) and not (layer2_outputs(2006));
    layer3_outputs(628) <= not(layer2_outputs(874)) or (layer2_outputs(4668));
    layer3_outputs(629) <= (layer2_outputs(3841)) xor (layer2_outputs(806));
    layer3_outputs(630) <= layer2_outputs(463);
    layer3_outputs(631) <= not((layer2_outputs(3524)) and (layer2_outputs(575)));
    layer3_outputs(632) <= (layer2_outputs(1545)) and (layer2_outputs(1348));
    layer3_outputs(633) <= layer2_outputs(2703);
    layer3_outputs(634) <= '1';
    layer3_outputs(635) <= (layer2_outputs(2324)) or (layer2_outputs(2012));
    layer3_outputs(636) <= not(layer2_outputs(4910)) or (layer2_outputs(2405));
    layer3_outputs(637) <= layer2_outputs(1779);
    layer3_outputs(638) <= '0';
    layer3_outputs(639) <= '1';
    layer3_outputs(640) <= not((layer2_outputs(977)) and (layer2_outputs(3493)));
    layer3_outputs(641) <= not((layer2_outputs(4906)) and (layer2_outputs(4441)));
    layer3_outputs(642) <= layer2_outputs(2390);
    layer3_outputs(643) <= layer2_outputs(1533);
    layer3_outputs(644) <= (layer2_outputs(2040)) and not (layer2_outputs(2807));
    layer3_outputs(645) <= '1';
    layer3_outputs(646) <= layer2_outputs(4868);
    layer3_outputs(647) <= not(layer2_outputs(2101)) or (layer2_outputs(4250));
    layer3_outputs(648) <= (layer2_outputs(606)) and not (layer2_outputs(5106));
    layer3_outputs(649) <= (layer2_outputs(3102)) and (layer2_outputs(2638));
    layer3_outputs(650) <= (layer2_outputs(3651)) or (layer2_outputs(3572));
    layer3_outputs(651) <= layer2_outputs(1428);
    layer3_outputs(652) <= not((layer2_outputs(4009)) or (layer2_outputs(885)));
    layer3_outputs(653) <= '1';
    layer3_outputs(654) <= (layer2_outputs(2034)) and not (layer2_outputs(3894));
    layer3_outputs(655) <= not((layer2_outputs(3729)) or (layer2_outputs(1505)));
    layer3_outputs(656) <= '1';
    layer3_outputs(657) <= (layer2_outputs(3425)) and not (layer2_outputs(3915));
    layer3_outputs(658) <= not(layer2_outputs(3302)) or (layer2_outputs(1209));
    layer3_outputs(659) <= not(layer2_outputs(1985));
    layer3_outputs(660) <= not(layer2_outputs(1517));
    layer3_outputs(661) <= not(layer2_outputs(3298));
    layer3_outputs(662) <= (layer2_outputs(1336)) or (layer2_outputs(4053));
    layer3_outputs(663) <= '1';
    layer3_outputs(664) <= (layer2_outputs(1212)) and (layer2_outputs(338));
    layer3_outputs(665) <= not(layer2_outputs(4775));
    layer3_outputs(666) <= not(layer2_outputs(1));
    layer3_outputs(667) <= '1';
    layer3_outputs(668) <= (layer2_outputs(4226)) or (layer2_outputs(2775));
    layer3_outputs(669) <= layer2_outputs(278);
    layer3_outputs(670) <= layer2_outputs(629);
    layer3_outputs(671) <= '0';
    layer3_outputs(672) <= '0';
    layer3_outputs(673) <= (layer2_outputs(1976)) and not (layer2_outputs(2277));
    layer3_outputs(674) <= (layer2_outputs(164)) and not (layer2_outputs(4920));
    layer3_outputs(675) <= not((layer2_outputs(4433)) and (layer2_outputs(3550)));
    layer3_outputs(676) <= not((layer2_outputs(4845)) and (layer2_outputs(645)));
    layer3_outputs(677) <= not((layer2_outputs(1613)) and (layer2_outputs(1170)));
    layer3_outputs(678) <= not(layer2_outputs(2395));
    layer3_outputs(679) <= not(layer2_outputs(209));
    layer3_outputs(680) <= not((layer2_outputs(2406)) and (layer2_outputs(5005)));
    layer3_outputs(681) <= not(layer2_outputs(4411)) or (layer2_outputs(3200));
    layer3_outputs(682) <= not(layer2_outputs(3147));
    layer3_outputs(683) <= not(layer2_outputs(1195));
    layer3_outputs(684) <= not(layer2_outputs(4815));
    layer3_outputs(685) <= (layer2_outputs(3283)) and (layer2_outputs(485));
    layer3_outputs(686) <= not(layer2_outputs(3855)) or (layer2_outputs(2933));
    layer3_outputs(687) <= (layer2_outputs(3366)) and not (layer2_outputs(3116));
    layer3_outputs(688) <= (layer2_outputs(2846)) or (layer2_outputs(776));
    layer3_outputs(689) <= not(layer2_outputs(2264));
    layer3_outputs(690) <= layer2_outputs(4175);
    layer3_outputs(691) <= not(layer2_outputs(892));
    layer3_outputs(692) <= not(layer2_outputs(74)) or (layer2_outputs(767));
    layer3_outputs(693) <= layer2_outputs(1873);
    layer3_outputs(694) <= '0';
    layer3_outputs(695) <= (layer2_outputs(1856)) xor (layer2_outputs(1615));
    layer3_outputs(696) <= not((layer2_outputs(461)) and (layer2_outputs(427)));
    layer3_outputs(697) <= not((layer2_outputs(762)) or (layer2_outputs(242)));
    layer3_outputs(698) <= layer2_outputs(1454);
    layer3_outputs(699) <= layer2_outputs(3496);
    layer3_outputs(700) <= not((layer2_outputs(2847)) and (layer2_outputs(2188)));
    layer3_outputs(701) <= (layer2_outputs(587)) or (layer2_outputs(1496));
    layer3_outputs(702) <= '1';
    layer3_outputs(703) <= not(layer2_outputs(538)) or (layer2_outputs(5042));
    layer3_outputs(704) <= not(layer2_outputs(4619));
    layer3_outputs(705) <= '1';
    layer3_outputs(706) <= layer2_outputs(1943);
    layer3_outputs(707) <= not(layer2_outputs(1777)) or (layer2_outputs(1027));
    layer3_outputs(708) <= '1';
    layer3_outputs(709) <= not((layer2_outputs(216)) and (layer2_outputs(4221)));
    layer3_outputs(710) <= '1';
    layer3_outputs(711) <= layer2_outputs(1104);
    layer3_outputs(712) <= not(layer2_outputs(3027));
    layer3_outputs(713) <= '1';
    layer3_outputs(714) <= (layer2_outputs(3993)) and not (layer2_outputs(3911));
    layer3_outputs(715) <= not(layer2_outputs(2066));
    layer3_outputs(716) <= (layer2_outputs(5020)) and (layer2_outputs(1939));
    layer3_outputs(717) <= (layer2_outputs(2503)) and (layer2_outputs(2094));
    layer3_outputs(718) <= '0';
    layer3_outputs(719) <= not(layer2_outputs(2582)) or (layer2_outputs(2259));
    layer3_outputs(720) <= not((layer2_outputs(1862)) and (layer2_outputs(977)));
    layer3_outputs(721) <= '0';
    layer3_outputs(722) <= '0';
    layer3_outputs(723) <= (layer2_outputs(4152)) or (layer2_outputs(1842));
    layer3_outputs(724) <= (layer2_outputs(2498)) and not (layer2_outputs(2262));
    layer3_outputs(725) <= (layer2_outputs(2106)) and not (layer2_outputs(1869));
    layer3_outputs(726) <= not(layer2_outputs(3662));
    layer3_outputs(727) <= not((layer2_outputs(987)) or (layer2_outputs(2164)));
    layer3_outputs(728) <= (layer2_outputs(1143)) and not (layer2_outputs(1476));
    layer3_outputs(729) <= (layer2_outputs(4707)) and not (layer2_outputs(2581));
    layer3_outputs(730) <= not(layer2_outputs(1994));
    layer3_outputs(731) <= (layer2_outputs(3094)) and not (layer2_outputs(2421));
    layer3_outputs(732) <= '1';
    layer3_outputs(733) <= not(layer2_outputs(5046));
    layer3_outputs(734) <= (layer2_outputs(4295)) or (layer2_outputs(2620));
    layer3_outputs(735) <= layer2_outputs(1423);
    layer3_outputs(736) <= '1';
    layer3_outputs(737) <= not(layer2_outputs(1982)) or (layer2_outputs(3554));
    layer3_outputs(738) <= (layer2_outputs(3053)) or (layer2_outputs(4279));
    layer3_outputs(739) <= (layer2_outputs(4059)) or (layer2_outputs(5104));
    layer3_outputs(740) <= (layer2_outputs(1473)) and not (layer2_outputs(4187));
    layer3_outputs(741) <= not((layer2_outputs(1252)) and (layer2_outputs(3057)));
    layer3_outputs(742) <= (layer2_outputs(2120)) and (layer2_outputs(4140));
    layer3_outputs(743) <= (layer2_outputs(1239)) and not (layer2_outputs(1305));
    layer3_outputs(744) <= (layer2_outputs(2312)) or (layer2_outputs(3180));
    layer3_outputs(745) <= not((layer2_outputs(300)) and (layer2_outputs(1515)));
    layer3_outputs(746) <= not((layer2_outputs(2643)) and (layer2_outputs(3253)));
    layer3_outputs(747) <= '1';
    layer3_outputs(748) <= not(layer2_outputs(2902)) or (layer2_outputs(2261));
    layer3_outputs(749) <= (layer2_outputs(4651)) and not (layer2_outputs(4629));
    layer3_outputs(750) <= (layer2_outputs(3332)) and not (layer2_outputs(1327));
    layer3_outputs(751) <= layer2_outputs(2667);
    layer3_outputs(752) <= '1';
    layer3_outputs(753) <= '0';
    layer3_outputs(754) <= (layer2_outputs(2712)) and not (layer2_outputs(1024));
    layer3_outputs(755) <= (layer2_outputs(618)) and not (layer2_outputs(3908));
    layer3_outputs(756) <= (layer2_outputs(1799)) xor (layer2_outputs(4633));
    layer3_outputs(757) <= not((layer2_outputs(3819)) or (layer2_outputs(2429)));
    layer3_outputs(758) <= (layer2_outputs(4518)) and not (layer2_outputs(3868));
    layer3_outputs(759) <= not(layer2_outputs(3847));
    layer3_outputs(760) <= layer2_outputs(3144);
    layer3_outputs(761) <= '1';
    layer3_outputs(762) <= layer2_outputs(2495);
    layer3_outputs(763) <= '0';
    layer3_outputs(764) <= '0';
    layer3_outputs(765) <= not(layer2_outputs(3005));
    layer3_outputs(766) <= '1';
    layer3_outputs(767) <= '0';
    layer3_outputs(768) <= '0';
    layer3_outputs(769) <= (layer2_outputs(623)) and not (layer2_outputs(2449));
    layer3_outputs(770) <= '1';
    layer3_outputs(771) <= layer2_outputs(883);
    layer3_outputs(772) <= not((layer2_outputs(2701)) xor (layer2_outputs(2992)));
    layer3_outputs(773) <= '1';
    layer3_outputs(774) <= (layer2_outputs(665)) and (layer2_outputs(4356));
    layer3_outputs(775) <= '0';
    layer3_outputs(776) <= not(layer2_outputs(1221)) or (layer2_outputs(3371));
    layer3_outputs(777) <= not((layer2_outputs(2375)) or (layer2_outputs(2543)));
    layer3_outputs(778) <= (layer2_outputs(1507)) and not (layer2_outputs(3317));
    layer3_outputs(779) <= not(layer2_outputs(3009)) or (layer2_outputs(498));
    layer3_outputs(780) <= '1';
    layer3_outputs(781) <= not(layer2_outputs(5088));
    layer3_outputs(782) <= (layer2_outputs(4895)) and not (layer2_outputs(4975));
    layer3_outputs(783) <= (layer2_outputs(1214)) or (layer2_outputs(2469));
    layer3_outputs(784) <= not((layer2_outputs(1203)) and (layer2_outputs(4966)));
    layer3_outputs(785) <= (layer2_outputs(3985)) and (layer2_outputs(4308));
    layer3_outputs(786) <= (layer2_outputs(3258)) and (layer2_outputs(1483));
    layer3_outputs(787) <= '0';
    layer3_outputs(788) <= layer2_outputs(2114);
    layer3_outputs(789) <= layer2_outputs(523);
    layer3_outputs(790) <= (layer2_outputs(499)) and not (layer2_outputs(3869));
    layer3_outputs(791) <= layer2_outputs(1614);
    layer3_outputs(792) <= (layer2_outputs(1505)) and not (layer2_outputs(3102));
    layer3_outputs(793) <= (layer2_outputs(1036)) and not (layer2_outputs(1154));
    layer3_outputs(794) <= (layer2_outputs(65)) and (layer2_outputs(376));
    layer3_outputs(795) <= (layer2_outputs(3568)) and not (layer2_outputs(2695));
    layer3_outputs(796) <= (layer2_outputs(1619)) or (layer2_outputs(1219));
    layer3_outputs(797) <= (layer2_outputs(1244)) and not (layer2_outputs(3793));
    layer3_outputs(798) <= (layer2_outputs(2753)) and not (layer2_outputs(2919));
    layer3_outputs(799) <= (layer2_outputs(1969)) and not (layer2_outputs(4137));
    layer3_outputs(800) <= (layer2_outputs(788)) and not (layer2_outputs(4263));
    layer3_outputs(801) <= (layer2_outputs(1295)) and not (layer2_outputs(1503));
    layer3_outputs(802) <= not(layer2_outputs(4646));
    layer3_outputs(803) <= not((layer2_outputs(3657)) or (layer2_outputs(564)));
    layer3_outputs(804) <= not((layer2_outputs(263)) or (layer2_outputs(3490)));
    layer3_outputs(805) <= not(layer2_outputs(462)) or (layer2_outputs(1840));
    layer3_outputs(806) <= not(layer2_outputs(2545)) or (layer2_outputs(4292));
    layer3_outputs(807) <= not((layer2_outputs(3644)) or (layer2_outputs(1072)));
    layer3_outputs(808) <= (layer2_outputs(1039)) and not (layer2_outputs(737));
    layer3_outputs(809) <= (layer2_outputs(101)) and not (layer2_outputs(1787));
    layer3_outputs(810) <= layer2_outputs(135);
    layer3_outputs(811) <= not(layer2_outputs(781)) or (layer2_outputs(2945));
    layer3_outputs(812) <= not(layer2_outputs(284)) or (layer2_outputs(1486));
    layer3_outputs(813) <= not((layer2_outputs(3203)) and (layer2_outputs(5108)));
    layer3_outputs(814) <= layer2_outputs(4135);
    layer3_outputs(815) <= '1';
    layer3_outputs(816) <= '0';
    layer3_outputs(817) <= '1';
    layer3_outputs(818) <= (layer2_outputs(2363)) and (layer2_outputs(173));
    layer3_outputs(819) <= layer2_outputs(2852);
    layer3_outputs(820) <= (layer2_outputs(2571)) and not (layer2_outputs(1928));
    layer3_outputs(821) <= (layer2_outputs(1472)) and not (layer2_outputs(3279));
    layer3_outputs(822) <= layer2_outputs(3125);
    layer3_outputs(823) <= (layer2_outputs(2584)) or (layer2_outputs(1527));
    layer3_outputs(824) <= (layer2_outputs(559)) and not (layer2_outputs(3293));
    layer3_outputs(825) <= (layer2_outputs(4237)) and (layer2_outputs(4432));
    layer3_outputs(826) <= (layer2_outputs(3395)) and (layer2_outputs(3796));
    layer3_outputs(827) <= not((layer2_outputs(2924)) and (layer2_outputs(4637)));
    layer3_outputs(828) <= not(layer2_outputs(2600));
    layer3_outputs(829) <= '1';
    layer3_outputs(830) <= (layer2_outputs(230)) and not (layer2_outputs(689));
    layer3_outputs(831) <= (layer2_outputs(1499)) and (layer2_outputs(2347));
    layer3_outputs(832) <= not((layer2_outputs(1810)) xor (layer2_outputs(4873)));
    layer3_outputs(833) <= not((layer2_outputs(4435)) or (layer2_outputs(112)));
    layer3_outputs(834) <= (layer2_outputs(3706)) and not (layer2_outputs(2959));
    layer3_outputs(835) <= (layer2_outputs(994)) and not (layer2_outputs(1065));
    layer3_outputs(836) <= layer2_outputs(3466);
    layer3_outputs(837) <= (layer2_outputs(1970)) or (layer2_outputs(3727));
    layer3_outputs(838) <= not(layer2_outputs(2392)) or (layer2_outputs(1929));
    layer3_outputs(839) <= layer2_outputs(3360);
    layer3_outputs(840) <= '0';
    layer3_outputs(841) <= (layer2_outputs(3538)) and not (layer2_outputs(866));
    layer3_outputs(842) <= not(layer2_outputs(4535)) or (layer2_outputs(3017));
    layer3_outputs(843) <= '1';
    layer3_outputs(844) <= not(layer2_outputs(2433));
    layer3_outputs(845) <= not((layer2_outputs(3124)) and (layer2_outputs(3686)));
    layer3_outputs(846) <= layer2_outputs(1485);
    layer3_outputs(847) <= '1';
    layer3_outputs(848) <= not(layer2_outputs(2918)) or (layer2_outputs(3759));
    layer3_outputs(849) <= '0';
    layer3_outputs(850) <= (layer2_outputs(4759)) and not (layer2_outputs(975));
    layer3_outputs(851) <= not((layer2_outputs(487)) and (layer2_outputs(4474)));
    layer3_outputs(852) <= not(layer2_outputs(2883));
    layer3_outputs(853) <= not((layer2_outputs(3429)) and (layer2_outputs(4427)));
    layer3_outputs(854) <= (layer2_outputs(3223)) and not (layer2_outputs(2368));
    layer3_outputs(855) <= (layer2_outputs(4758)) or (layer2_outputs(503));
    layer3_outputs(856) <= not((layer2_outputs(5024)) and (layer2_outputs(4484)));
    layer3_outputs(857) <= (layer2_outputs(1697)) xor (layer2_outputs(2739));
    layer3_outputs(858) <= not(layer2_outputs(2817)) or (layer2_outputs(2679));
    layer3_outputs(859) <= (layer2_outputs(491)) and not (layer2_outputs(4460));
    layer3_outputs(860) <= '1';
    layer3_outputs(861) <= (layer2_outputs(1363)) or (layer2_outputs(4686));
    layer3_outputs(862) <= not(layer2_outputs(4434)) or (layer2_outputs(4642));
    layer3_outputs(863) <= (layer2_outputs(2545)) and not (layer2_outputs(281));
    layer3_outputs(864) <= (layer2_outputs(1232)) and (layer2_outputs(25));
    layer3_outputs(865) <= '0';
    layer3_outputs(866) <= '0';
    layer3_outputs(867) <= (layer2_outputs(2146)) or (layer2_outputs(1627));
    layer3_outputs(868) <= not((layer2_outputs(2781)) or (layer2_outputs(3441)));
    layer3_outputs(869) <= not(layer2_outputs(329));
    layer3_outputs(870) <= layer2_outputs(217);
    layer3_outputs(871) <= not((layer2_outputs(1024)) xor (layer2_outputs(3016)));
    layer3_outputs(872) <= (layer2_outputs(2974)) and not (layer2_outputs(760));
    layer3_outputs(873) <= (layer2_outputs(2145)) and not (layer2_outputs(5038));
    layer3_outputs(874) <= (layer2_outputs(3174)) xor (layer2_outputs(1443));
    layer3_outputs(875) <= (layer2_outputs(1077)) and not (layer2_outputs(1367));
    layer3_outputs(876) <= not(layer2_outputs(2620)) or (layer2_outputs(323));
    layer3_outputs(877) <= not(layer2_outputs(1629));
    layer3_outputs(878) <= '0';
    layer3_outputs(879) <= (layer2_outputs(2361)) and not (layer2_outputs(2786));
    layer3_outputs(880) <= not(layer2_outputs(1447)) or (layer2_outputs(936));
    layer3_outputs(881) <= layer2_outputs(648);
    layer3_outputs(882) <= (layer2_outputs(4624)) and not (layer2_outputs(5024));
    layer3_outputs(883) <= (layer2_outputs(3087)) and (layer2_outputs(646));
    layer3_outputs(884) <= not(layer2_outputs(3560));
    layer3_outputs(885) <= '1';
    layer3_outputs(886) <= not(layer2_outputs(1023)) or (layer2_outputs(4051));
    layer3_outputs(887) <= not(layer2_outputs(1784));
    layer3_outputs(888) <= not(layer2_outputs(4606));
    layer3_outputs(889) <= (layer2_outputs(3571)) and not (layer2_outputs(2225));
    layer3_outputs(890) <= '0';
    layer3_outputs(891) <= not(layer2_outputs(4129));
    layer3_outputs(892) <= not(layer2_outputs(56)) or (layer2_outputs(1804));
    layer3_outputs(893) <= layer2_outputs(1007);
    layer3_outputs(894) <= (layer2_outputs(3106)) or (layer2_outputs(4542));
    layer3_outputs(895) <= layer2_outputs(187);
    layer3_outputs(896) <= (layer2_outputs(1531)) and not (layer2_outputs(2335));
    layer3_outputs(897) <= not((layer2_outputs(4194)) or (layer2_outputs(4366)));
    layer3_outputs(898) <= layer2_outputs(1355);
    layer3_outputs(899) <= layer2_outputs(3252);
    layer3_outputs(900) <= (layer2_outputs(1037)) or (layer2_outputs(1009));
    layer3_outputs(901) <= '0';
    layer3_outputs(902) <= not(layer2_outputs(4743)) or (layer2_outputs(3856));
    layer3_outputs(903) <= (layer2_outputs(718)) and (layer2_outputs(2900));
    layer3_outputs(904) <= '0';
    layer3_outputs(905) <= '0';
    layer3_outputs(906) <= (layer2_outputs(4803)) or (layer2_outputs(155));
    layer3_outputs(907) <= '1';
    layer3_outputs(908) <= (layer2_outputs(1625)) and not (layer2_outputs(137));
    layer3_outputs(909) <= '1';
    layer3_outputs(910) <= not(layer2_outputs(265)) or (layer2_outputs(1048));
    layer3_outputs(911) <= '1';
    layer3_outputs(912) <= not(layer2_outputs(2894));
    layer3_outputs(913) <= '1';
    layer3_outputs(914) <= '1';
    layer3_outputs(915) <= not(layer2_outputs(3692));
    layer3_outputs(916) <= not((layer2_outputs(1318)) and (layer2_outputs(2256)));
    layer3_outputs(917) <= (layer2_outputs(1931)) and (layer2_outputs(2771));
    layer3_outputs(918) <= (layer2_outputs(3513)) and (layer2_outputs(681));
    layer3_outputs(919) <= (layer2_outputs(4498)) and not (layer2_outputs(2996));
    layer3_outputs(920) <= (layer2_outputs(824)) and (layer2_outputs(2817));
    layer3_outputs(921) <= layer2_outputs(3889);
    layer3_outputs(922) <= (layer2_outputs(1502)) or (layer2_outputs(2237));
    layer3_outputs(923) <= not((layer2_outputs(4702)) and (layer2_outputs(292)));
    layer3_outputs(924) <= layer2_outputs(4119);
    layer3_outputs(925) <= (layer2_outputs(922)) and (layer2_outputs(1353));
    layer3_outputs(926) <= '1';
    layer3_outputs(927) <= not(layer2_outputs(3027));
    layer3_outputs(928) <= (layer2_outputs(1343)) and (layer2_outputs(28));
    layer3_outputs(929) <= '0';
    layer3_outputs(930) <= not(layer2_outputs(3065));
    layer3_outputs(931) <= layer2_outputs(1514);
    layer3_outputs(932) <= (layer2_outputs(644)) and not (layer2_outputs(3042));
    layer3_outputs(933) <= not(layer2_outputs(2932));
    layer3_outputs(934) <= '0';
    layer3_outputs(935) <= '1';
    layer3_outputs(936) <= (layer2_outputs(1105)) and not (layer2_outputs(5100));
    layer3_outputs(937) <= (layer2_outputs(4134)) or (layer2_outputs(1900));
    layer3_outputs(938) <= (layer2_outputs(3066)) and not (layer2_outputs(1852));
    layer3_outputs(939) <= '1';
    layer3_outputs(940) <= (layer2_outputs(4128)) and not (layer2_outputs(2113));
    layer3_outputs(941) <= (layer2_outputs(2968)) and (layer2_outputs(1899));
    layer3_outputs(942) <= not(layer2_outputs(2611)) or (layer2_outputs(4054));
    layer3_outputs(943) <= not(layer2_outputs(2580)) or (layer2_outputs(2348));
    layer3_outputs(944) <= (layer2_outputs(4005)) and not (layer2_outputs(1973));
    layer3_outputs(945) <= not(layer2_outputs(2475)) or (layer2_outputs(3862));
    layer3_outputs(946) <= layer2_outputs(3721);
    layer3_outputs(947) <= not(layer2_outputs(4626));
    layer3_outputs(948) <= layer2_outputs(4131);
    layer3_outputs(949) <= not((layer2_outputs(884)) or (layer2_outputs(1450)));
    layer3_outputs(950) <= not(layer2_outputs(3060)) or (layer2_outputs(4482));
    layer3_outputs(951) <= not(layer2_outputs(530)) or (layer2_outputs(2638));
    layer3_outputs(952) <= '0';
    layer3_outputs(953) <= not(layer2_outputs(3116)) or (layer2_outputs(3300));
    layer3_outputs(954) <= not((layer2_outputs(4756)) or (layer2_outputs(4690)));
    layer3_outputs(955) <= (layer2_outputs(4183)) and (layer2_outputs(3159));
    layer3_outputs(956) <= layer2_outputs(3685);
    layer3_outputs(957) <= not(layer2_outputs(2459));
    layer3_outputs(958) <= (layer2_outputs(2443)) or (layer2_outputs(1963));
    layer3_outputs(959) <= '1';
    layer3_outputs(960) <= not(layer2_outputs(808));
    layer3_outputs(961) <= '0';
    layer3_outputs(962) <= '1';
    layer3_outputs(963) <= '0';
    layer3_outputs(964) <= (layer2_outputs(1011)) and not (layer2_outputs(2412));
    layer3_outputs(965) <= not(layer2_outputs(2319)) or (layer2_outputs(3105));
    layer3_outputs(966) <= '0';
    layer3_outputs(967) <= not(layer2_outputs(1933));
    layer3_outputs(968) <= not(layer2_outputs(2542)) or (layer2_outputs(4229));
    layer3_outputs(969) <= not(layer2_outputs(1304)) or (layer2_outputs(4554));
    layer3_outputs(970) <= not(layer2_outputs(2560));
    layer3_outputs(971) <= not(layer2_outputs(3748)) or (layer2_outputs(3190));
    layer3_outputs(972) <= layer2_outputs(1984);
    layer3_outputs(973) <= '1';
    layer3_outputs(974) <= not(layer2_outputs(3167)) or (layer2_outputs(5029));
    layer3_outputs(975) <= layer2_outputs(1693);
    layer3_outputs(976) <= '1';
    layer3_outputs(977) <= (layer2_outputs(155)) or (layer2_outputs(2244));
    layer3_outputs(978) <= not(layer2_outputs(1419));
    layer3_outputs(979) <= '0';
    layer3_outputs(980) <= '1';
    layer3_outputs(981) <= layer2_outputs(1843);
    layer3_outputs(982) <= '0';
    layer3_outputs(983) <= not(layer2_outputs(2806)) or (layer2_outputs(2777));
    layer3_outputs(984) <= not(layer2_outputs(447));
    layer3_outputs(985) <= (layer2_outputs(1296)) and (layer2_outputs(3582));
    layer3_outputs(986) <= not((layer2_outputs(2352)) and (layer2_outputs(4056)));
    layer3_outputs(987) <= not(layer2_outputs(1117));
    layer3_outputs(988) <= '1';
    layer3_outputs(989) <= '1';
    layer3_outputs(990) <= not(layer2_outputs(598));
    layer3_outputs(991) <= '0';
    layer3_outputs(992) <= not(layer2_outputs(144));
    layer3_outputs(993) <= (layer2_outputs(1008)) and (layer2_outputs(873));
    layer3_outputs(994) <= '1';
    layer3_outputs(995) <= not((layer2_outputs(4812)) and (layer2_outputs(1028)));
    layer3_outputs(996) <= (layer2_outputs(1915)) or (layer2_outputs(497));
    layer3_outputs(997) <= '0';
    layer3_outputs(998) <= (layer2_outputs(1816)) and (layer2_outputs(91));
    layer3_outputs(999) <= '1';
    layer3_outputs(1000) <= (layer2_outputs(2450)) and not (layer2_outputs(2562));
    layer3_outputs(1001) <= not(layer2_outputs(4264)) or (layer2_outputs(784));
    layer3_outputs(1002) <= (layer2_outputs(2482)) and not (layer2_outputs(4523));
    layer3_outputs(1003) <= not(layer2_outputs(1238));
    layer3_outputs(1004) <= layer2_outputs(4248);
    layer3_outputs(1005) <= not(layer2_outputs(3098));
    layer3_outputs(1006) <= layer2_outputs(1057);
    layer3_outputs(1007) <= (layer2_outputs(1032)) and not (layer2_outputs(2036));
    layer3_outputs(1008) <= '1';
    layer3_outputs(1009) <= not(layer2_outputs(255)) or (layer2_outputs(1517));
    layer3_outputs(1010) <= not(layer2_outputs(235)) or (layer2_outputs(285));
    layer3_outputs(1011) <= not(layer2_outputs(4198)) or (layer2_outputs(2351));
    layer3_outputs(1012) <= not((layer2_outputs(3307)) xor (layer2_outputs(4784)));
    layer3_outputs(1013) <= (layer2_outputs(4797)) and (layer2_outputs(790));
    layer3_outputs(1014) <= (layer2_outputs(3587)) and (layer2_outputs(4545));
    layer3_outputs(1015) <= not((layer2_outputs(4408)) and (layer2_outputs(2731)));
    layer3_outputs(1016) <= (layer2_outputs(4400)) and (layer2_outputs(1311));
    layer3_outputs(1017) <= not((layer2_outputs(3677)) and (layer2_outputs(279)));
    layer3_outputs(1018) <= (layer2_outputs(1806)) and (layer2_outputs(2484));
    layer3_outputs(1019) <= not(layer2_outputs(3034));
    layer3_outputs(1020) <= (layer2_outputs(727)) and (layer2_outputs(4930));
    layer3_outputs(1021) <= '0';
    layer3_outputs(1022) <= '0';
    layer3_outputs(1023) <= '1';
    layer3_outputs(1024) <= not(layer2_outputs(2010));
    layer3_outputs(1025) <= (layer2_outputs(3427)) and (layer2_outputs(169));
    layer3_outputs(1026) <= not(layer2_outputs(2268));
    layer3_outputs(1027) <= not(layer2_outputs(2530)) or (layer2_outputs(3498));
    layer3_outputs(1028) <= not(layer2_outputs(2166));
    layer3_outputs(1029) <= layer2_outputs(360);
    layer3_outputs(1030) <= '1';
    layer3_outputs(1031) <= not(layer2_outputs(2982)) or (layer2_outputs(2478));
    layer3_outputs(1032) <= (layer2_outputs(2647)) or (layer2_outputs(134));
    layer3_outputs(1033) <= (layer2_outputs(4162)) and not (layer2_outputs(4905));
    layer3_outputs(1034) <= not(layer2_outputs(4088)) or (layer2_outputs(4507));
    layer3_outputs(1035) <= not(layer2_outputs(277));
    layer3_outputs(1036) <= layer2_outputs(2821);
    layer3_outputs(1037) <= (layer2_outputs(3404)) xor (layer2_outputs(5081));
    layer3_outputs(1038) <= not((layer2_outputs(3999)) or (layer2_outputs(868)));
    layer3_outputs(1039) <= not(layer2_outputs(3143));
    layer3_outputs(1040) <= '1';
    layer3_outputs(1041) <= '0';
    layer3_outputs(1042) <= not(layer2_outputs(2149));
    layer3_outputs(1043) <= '1';
    layer3_outputs(1044) <= '1';
    layer3_outputs(1045) <= not(layer2_outputs(3674)) or (layer2_outputs(188));
    layer3_outputs(1046) <= not((layer2_outputs(458)) or (layer2_outputs(2566)));
    layer3_outputs(1047) <= layer2_outputs(4701);
    layer3_outputs(1048) <= layer2_outputs(296);
    layer3_outputs(1049) <= '0';
    layer3_outputs(1050) <= (layer2_outputs(2842)) and (layer2_outputs(4741));
    layer3_outputs(1051) <= '0';
    layer3_outputs(1052) <= (layer2_outputs(4727)) and not (layer2_outputs(3952));
    layer3_outputs(1053) <= not(layer2_outputs(3238));
    layer3_outputs(1054) <= (layer2_outputs(4189)) and not (layer2_outputs(1219));
    layer3_outputs(1055) <= (layer2_outputs(3581)) and not (layer2_outputs(4640));
    layer3_outputs(1056) <= not(layer2_outputs(1262));
    layer3_outputs(1057) <= (layer2_outputs(2304)) or (layer2_outputs(3465));
    layer3_outputs(1058) <= (layer2_outputs(362)) xor (layer2_outputs(4126));
    layer3_outputs(1059) <= (layer2_outputs(3828)) and (layer2_outputs(624));
    layer3_outputs(1060) <= layer2_outputs(1773);
    layer3_outputs(1061) <= (layer2_outputs(1726)) and (layer2_outputs(3235));
    layer3_outputs(1062) <= not(layer2_outputs(4078));
    layer3_outputs(1063) <= (layer2_outputs(412)) and not (layer2_outputs(764));
    layer3_outputs(1064) <= not(layer2_outputs(2071)) or (layer2_outputs(1425));
    layer3_outputs(1065) <= (layer2_outputs(111)) and not (layer2_outputs(856));
    layer3_outputs(1066) <= not((layer2_outputs(4186)) or (layer2_outputs(4721)));
    layer3_outputs(1067) <= not((layer2_outputs(4344)) and (layer2_outputs(4640)));
    layer3_outputs(1068) <= not(layer2_outputs(2795)) or (layer2_outputs(4554));
    layer3_outputs(1069) <= not(layer2_outputs(4170)) or (layer2_outputs(2622));
    layer3_outputs(1070) <= not((layer2_outputs(1868)) or (layer2_outputs(1564)));
    layer3_outputs(1071) <= layer2_outputs(3937);
    layer3_outputs(1072) <= '0';
    layer3_outputs(1073) <= not(layer2_outputs(42)) or (layer2_outputs(3921));
    layer3_outputs(1074) <= not((layer2_outputs(1328)) xor (layer2_outputs(4921)));
    layer3_outputs(1075) <= '0';
    layer3_outputs(1076) <= not(layer2_outputs(2766)) or (layer2_outputs(2528));
    layer3_outputs(1077) <= layer2_outputs(1235);
    layer3_outputs(1078) <= not(layer2_outputs(646));
    layer3_outputs(1079) <= (layer2_outputs(2067)) or (layer2_outputs(2920));
    layer3_outputs(1080) <= '1';
    layer3_outputs(1081) <= layer2_outputs(1030);
    layer3_outputs(1082) <= (layer2_outputs(4335)) and (layer2_outputs(1933));
    layer3_outputs(1083) <= not((layer2_outputs(2111)) or (layer2_outputs(3381)));
    layer3_outputs(1084) <= (layer2_outputs(1009)) or (layer2_outputs(4576));
    layer3_outputs(1085) <= layer2_outputs(2612);
    layer3_outputs(1086) <= (layer2_outputs(306)) and (layer2_outputs(2588));
    layer3_outputs(1087) <= (layer2_outputs(1830)) and (layer2_outputs(1586));
    layer3_outputs(1088) <= (layer2_outputs(2485)) and (layer2_outputs(2625));
    layer3_outputs(1089) <= layer2_outputs(4305);
    layer3_outputs(1090) <= not(layer2_outputs(1308));
    layer3_outputs(1091) <= (layer2_outputs(1539)) or (layer2_outputs(4271));
    layer3_outputs(1092) <= not(layer2_outputs(488));
    layer3_outputs(1093) <= not(layer2_outputs(4046)) or (layer2_outputs(3234));
    layer3_outputs(1094) <= '0';
    layer3_outputs(1095) <= (layer2_outputs(4029)) or (layer2_outputs(3482));
    layer3_outputs(1096) <= (layer2_outputs(1075)) and not (layer2_outputs(2326));
    layer3_outputs(1097) <= not((layer2_outputs(5114)) or (layer2_outputs(3990)));
    layer3_outputs(1098) <= (layer2_outputs(3778)) and not (layer2_outputs(1336));
    layer3_outputs(1099) <= (layer2_outputs(4835)) and not (layer2_outputs(1094));
    layer3_outputs(1100) <= not(layer2_outputs(899));
    layer3_outputs(1101) <= layer2_outputs(3737);
    layer3_outputs(1102) <= layer2_outputs(3599);
    layer3_outputs(1103) <= layer2_outputs(4212);
    layer3_outputs(1104) <= layer2_outputs(733);
    layer3_outputs(1105) <= (layer2_outputs(3221)) and not (layer2_outputs(886));
    layer3_outputs(1106) <= not(layer2_outputs(1620));
    layer3_outputs(1107) <= '1';
    layer3_outputs(1108) <= layer2_outputs(1040);
    layer3_outputs(1109) <= '1';
    layer3_outputs(1110) <= '1';
    layer3_outputs(1111) <= (layer2_outputs(3570)) and not (layer2_outputs(1404));
    layer3_outputs(1112) <= not(layer2_outputs(3650));
    layer3_outputs(1113) <= '0';
    layer3_outputs(1114) <= '1';
    layer3_outputs(1115) <= not(layer2_outputs(3975)) or (layer2_outputs(2006));
    layer3_outputs(1116) <= (layer2_outputs(2073)) or (layer2_outputs(1381));
    layer3_outputs(1117) <= not((layer2_outputs(2840)) and (layer2_outputs(694)));
    layer3_outputs(1118) <= (layer2_outputs(2153)) and (layer2_outputs(1053));
    layer3_outputs(1119) <= (layer2_outputs(4160)) and not (layer2_outputs(4525));
    layer3_outputs(1120) <= (layer2_outputs(3401)) and not (layer2_outputs(352));
    layer3_outputs(1121) <= not(layer2_outputs(590)) or (layer2_outputs(3269));
    layer3_outputs(1122) <= '1';
    layer3_outputs(1123) <= (layer2_outputs(1346)) and not (layer2_outputs(5105));
    layer3_outputs(1124) <= '0';
    layer3_outputs(1125) <= '1';
    layer3_outputs(1126) <= layer2_outputs(460);
    layer3_outputs(1127) <= not(layer2_outputs(2836));
    layer3_outputs(1128) <= not((layer2_outputs(49)) and (layer2_outputs(3380)));
    layer3_outputs(1129) <= not(layer2_outputs(3416));
    layer3_outputs(1130) <= not(layer2_outputs(4145));
    layer3_outputs(1131) <= (layer2_outputs(2474)) xor (layer2_outputs(622));
    layer3_outputs(1132) <= (layer2_outputs(766)) and (layer2_outputs(3099));
    layer3_outputs(1133) <= (layer2_outputs(5040)) and (layer2_outputs(394));
    layer3_outputs(1134) <= not((layer2_outputs(2009)) and (layer2_outputs(1119)));
    layer3_outputs(1135) <= layer2_outputs(1207);
    layer3_outputs(1136) <= (layer2_outputs(386)) and not (layer2_outputs(2397));
    layer3_outputs(1137) <= '1';
    layer3_outputs(1138) <= not((layer2_outputs(4632)) or (layer2_outputs(4774)));
    layer3_outputs(1139) <= (layer2_outputs(1388)) and not (layer2_outputs(3362));
    layer3_outputs(1140) <= not(layer2_outputs(1662));
    layer3_outputs(1141) <= not(layer2_outputs(3907)) or (layer2_outputs(1390));
    layer3_outputs(1142) <= not(layer2_outputs(3109));
    layer3_outputs(1143) <= (layer2_outputs(553)) or (layer2_outputs(4153));
    layer3_outputs(1144) <= not((layer2_outputs(599)) xor (layer2_outputs(2146)));
    layer3_outputs(1145) <= not(layer2_outputs(5053));
    layer3_outputs(1146) <= (layer2_outputs(3205)) and not (layer2_outputs(1134));
    layer3_outputs(1147) <= layer2_outputs(2631);
    layer3_outputs(1148) <= '0';
    layer3_outputs(1149) <= (layer2_outputs(1883)) or (layer2_outputs(602));
    layer3_outputs(1150) <= (layer2_outputs(942)) and not (layer2_outputs(4968));
    layer3_outputs(1151) <= not(layer2_outputs(1089)) or (layer2_outputs(3633));
    layer3_outputs(1152) <= (layer2_outputs(4559)) or (layer2_outputs(3850));
    layer3_outputs(1153) <= '0';
    layer3_outputs(1154) <= layer2_outputs(3808);
    layer3_outputs(1155) <= not(layer2_outputs(4712)) or (layer2_outputs(2223));
    layer3_outputs(1156) <= layer2_outputs(1155);
    layer3_outputs(1157) <= not((layer2_outputs(2858)) or (layer2_outputs(1063)));
    layer3_outputs(1158) <= (layer2_outputs(4568)) and not (layer2_outputs(14));
    layer3_outputs(1159) <= '1';
    layer3_outputs(1160) <= not((layer2_outputs(3576)) xor (layer2_outputs(3809)));
    layer3_outputs(1161) <= layer2_outputs(2726);
    layer3_outputs(1162) <= layer2_outputs(4597);
    layer3_outputs(1163) <= (layer2_outputs(4551)) and not (layer2_outputs(2206));
    layer3_outputs(1164) <= (layer2_outputs(3532)) and not (layer2_outputs(2212));
    layer3_outputs(1165) <= layer2_outputs(3714);
    layer3_outputs(1166) <= '0';
    layer3_outputs(1167) <= (layer2_outputs(4478)) and not (layer2_outputs(1516));
    layer3_outputs(1168) <= '1';
    layer3_outputs(1169) <= not(layer2_outputs(4407)) or (layer2_outputs(2550));
    layer3_outputs(1170) <= '1';
    layer3_outputs(1171) <= not(layer2_outputs(1417)) or (layer2_outputs(1448));
    layer3_outputs(1172) <= (layer2_outputs(2236)) and not (layer2_outputs(3297));
    layer3_outputs(1173) <= (layer2_outputs(519)) and not (layer2_outputs(1202));
    layer3_outputs(1174) <= '0';
    layer3_outputs(1175) <= (layer2_outputs(3538)) and not (layer2_outputs(3259));
    layer3_outputs(1176) <= (layer2_outputs(2484)) and (layer2_outputs(1795));
    layer3_outputs(1177) <= not((layer2_outputs(4076)) and (layer2_outputs(4914)));
    layer3_outputs(1178) <= not((layer2_outputs(4572)) and (layer2_outputs(221)));
    layer3_outputs(1179) <= (layer2_outputs(2783)) or (layer2_outputs(88));
    layer3_outputs(1180) <= not(layer2_outputs(1997));
    layer3_outputs(1181) <= '1';
    layer3_outputs(1182) <= (layer2_outputs(953)) or (layer2_outputs(3183));
    layer3_outputs(1183) <= not(layer2_outputs(65));
    layer3_outputs(1184) <= layer2_outputs(2708);
    layer3_outputs(1185) <= '0';
    layer3_outputs(1186) <= not((layer2_outputs(3499)) and (layer2_outputs(4939)));
    layer3_outputs(1187) <= (layer2_outputs(787)) and (layer2_outputs(4859));
    layer3_outputs(1188) <= not(layer2_outputs(3177)) or (layer2_outputs(4045));
    layer3_outputs(1189) <= not(layer2_outputs(2792)) or (layer2_outputs(998));
    layer3_outputs(1190) <= not(layer2_outputs(418));
    layer3_outputs(1191) <= layer2_outputs(4581);
    layer3_outputs(1192) <= not(layer2_outputs(4254));
    layer3_outputs(1193) <= layer2_outputs(3074);
    layer3_outputs(1194) <= (layer2_outputs(4710)) and not (layer2_outputs(2816));
    layer3_outputs(1195) <= (layer2_outputs(1720)) or (layer2_outputs(500));
    layer3_outputs(1196) <= '0';
    layer3_outputs(1197) <= not(layer2_outputs(313)) or (layer2_outputs(1426));
    layer3_outputs(1198) <= (layer2_outputs(1702)) and not (layer2_outputs(636));
    layer3_outputs(1199) <= layer2_outputs(3263);
    layer3_outputs(1200) <= layer2_outputs(2984);
    layer3_outputs(1201) <= not(layer2_outputs(3484));
    layer3_outputs(1202) <= not((layer2_outputs(374)) or (layer2_outputs(1410)));
    layer3_outputs(1203) <= layer2_outputs(2339);
    layer3_outputs(1204) <= (layer2_outputs(4102)) and (layer2_outputs(90));
    layer3_outputs(1205) <= not((layer2_outputs(1747)) or (layer2_outputs(456)));
    layer3_outputs(1206) <= '1';
    layer3_outputs(1207) <= not(layer2_outputs(4385)) or (layer2_outputs(3669));
    layer3_outputs(1208) <= '0';
    layer3_outputs(1209) <= (layer2_outputs(3345)) and not (layer2_outputs(1073));
    layer3_outputs(1210) <= (layer2_outputs(531)) and not (layer2_outputs(1720));
    layer3_outputs(1211) <= not(layer2_outputs(1992));
    layer3_outputs(1212) <= (layer2_outputs(4628)) and not (layer2_outputs(4172));
    layer3_outputs(1213) <= not(layer2_outputs(1612));
    layer3_outputs(1214) <= not(layer2_outputs(522)) or (layer2_outputs(4591));
    layer3_outputs(1215) <= not(layer2_outputs(149)) or (layer2_outputs(605));
    layer3_outputs(1216) <= not(layer2_outputs(1412)) or (layer2_outputs(3977));
    layer3_outputs(1217) <= not((layer2_outputs(2468)) and (layer2_outputs(2717)));
    layer3_outputs(1218) <= (layer2_outputs(4267)) xor (layer2_outputs(4067));
    layer3_outputs(1219) <= not((layer2_outputs(3722)) or (layer2_outputs(1094)));
    layer3_outputs(1220) <= not(layer2_outputs(2539));
    layer3_outputs(1221) <= not((layer2_outputs(4496)) or (layer2_outputs(1844)));
    layer3_outputs(1222) <= not(layer2_outputs(834));
    layer3_outputs(1223) <= '1';
    layer3_outputs(1224) <= layer2_outputs(3585);
    layer3_outputs(1225) <= not((layer2_outputs(4598)) and (layer2_outputs(2267)));
    layer3_outputs(1226) <= not(layer2_outputs(445)) or (layer2_outputs(4703));
    layer3_outputs(1227) <= '1';
    layer3_outputs(1228) <= (layer2_outputs(4510)) or (layer2_outputs(1891));
    layer3_outputs(1229) <= layer2_outputs(1579);
    layer3_outputs(1230) <= (layer2_outputs(912)) xor (layer2_outputs(2377));
    layer3_outputs(1231) <= '1';
    layer3_outputs(1232) <= (layer2_outputs(136)) and not (layer2_outputs(3604));
    layer3_outputs(1233) <= (layer2_outputs(4753)) and not (layer2_outputs(2434));
    layer3_outputs(1234) <= layer2_outputs(372);
    layer3_outputs(1235) <= (layer2_outputs(3071)) or (layer2_outputs(4531));
    layer3_outputs(1236) <= '1';
    layer3_outputs(1237) <= not(layer2_outputs(4878)) or (layer2_outputs(973));
    layer3_outputs(1238) <= not((layer2_outputs(594)) and (layer2_outputs(3865)));
    layer3_outputs(1239) <= (layer2_outputs(2837)) and not (layer2_outputs(1798));
    layer3_outputs(1240) <= '0';
    layer3_outputs(1241) <= (layer2_outputs(1344)) or (layer2_outputs(1506));
    layer3_outputs(1242) <= not(layer2_outputs(1995));
    layer3_outputs(1243) <= '1';
    layer3_outputs(1244) <= layer2_outputs(1467);
    layer3_outputs(1245) <= '0';
    layer3_outputs(1246) <= (layer2_outputs(4992)) and (layer2_outputs(4317));
    layer3_outputs(1247) <= (layer2_outputs(4541)) or (layer2_outputs(4365));
    layer3_outputs(1248) <= not((layer2_outputs(3688)) and (layer2_outputs(465)));
    layer3_outputs(1249) <= layer2_outputs(3285);
    layer3_outputs(1250) <= not((layer2_outputs(3340)) or (layer2_outputs(2900)));
    layer3_outputs(1251) <= (layer2_outputs(563)) and not (layer2_outputs(4098));
    layer3_outputs(1252) <= (layer2_outputs(4947)) and not (layer2_outputs(1968));
    layer3_outputs(1253) <= '1';
    layer3_outputs(1254) <= layer2_outputs(182);
    layer3_outputs(1255) <= (layer2_outputs(1107)) or (layer2_outputs(3847));
    layer3_outputs(1256) <= (layer2_outputs(2521)) and (layer2_outputs(271));
    layer3_outputs(1257) <= '0';
    layer3_outputs(1258) <= '0';
    layer3_outputs(1259) <= '1';
    layer3_outputs(1260) <= not((layer2_outputs(3905)) or (layer2_outputs(1274)));
    layer3_outputs(1261) <= not((layer2_outputs(905)) and (layer2_outputs(1665)));
    layer3_outputs(1262) <= not(layer2_outputs(3511)) or (layer2_outputs(3324));
    layer3_outputs(1263) <= not((layer2_outputs(3055)) and (layer2_outputs(1512)));
    layer3_outputs(1264) <= '0';
    layer3_outputs(1265) <= not((layer2_outputs(1250)) and (layer2_outputs(858)));
    layer3_outputs(1266) <= '1';
    layer3_outputs(1267) <= not((layer2_outputs(4343)) and (layer2_outputs(1919)));
    layer3_outputs(1268) <= not(layer2_outputs(4817)) or (layer2_outputs(1838));
    layer3_outputs(1269) <= not(layer2_outputs(4028)) or (layer2_outputs(4063));
    layer3_outputs(1270) <= not(layer2_outputs(5043)) or (layer2_outputs(4210));
    layer3_outputs(1271) <= not(layer2_outputs(2820));
    layer3_outputs(1272) <= (layer2_outputs(1264)) or (layer2_outputs(508));
    layer3_outputs(1273) <= (layer2_outputs(2422)) and (layer2_outputs(948));
    layer3_outputs(1274) <= layer2_outputs(1198);
    layer3_outputs(1275) <= not((layer2_outputs(2353)) and (layer2_outputs(3951)));
    layer3_outputs(1276) <= not(layer2_outputs(743));
    layer3_outputs(1277) <= (layer2_outputs(1841)) and not (layer2_outputs(4579));
    layer3_outputs(1278) <= (layer2_outputs(1097)) xor (layer2_outputs(4272));
    layer3_outputs(1279) <= not(layer2_outputs(4246));
    layer3_outputs(1280) <= '1';
    layer3_outputs(1281) <= (layer2_outputs(3765)) xor (layer2_outputs(1082));
    layer3_outputs(1282) <= (layer2_outputs(925)) or (layer2_outputs(600));
    layer3_outputs(1283) <= not(layer2_outputs(1060)) or (layer2_outputs(3157));
    layer3_outputs(1284) <= not(layer2_outputs(628)) or (layer2_outputs(2833));
    layer3_outputs(1285) <= (layer2_outputs(3980)) and (layer2_outputs(2316));
    layer3_outputs(1286) <= not((layer2_outputs(2497)) and (layer2_outputs(3915)));
    layer3_outputs(1287) <= '1';
    layer3_outputs(1288) <= '0';
    layer3_outputs(1289) <= (layer2_outputs(2023)) and (layer2_outputs(22));
    layer3_outputs(1290) <= not(layer2_outputs(3074)) or (layer2_outputs(4093));
    layer3_outputs(1291) <= (layer2_outputs(3291)) and not (layer2_outputs(4144));
    layer3_outputs(1292) <= layer2_outputs(2275);
    layer3_outputs(1293) <= (layer2_outputs(1171)) and not (layer2_outputs(797));
    layer3_outputs(1294) <= (layer2_outputs(2488)) or (layer2_outputs(3939));
    layer3_outputs(1295) <= (layer2_outputs(4269)) and (layer2_outputs(1312));
    layer3_outputs(1296) <= not(layer2_outputs(4459)) or (layer2_outputs(771));
    layer3_outputs(1297) <= not((layer2_outputs(3089)) or (layer2_outputs(2859)));
    layer3_outputs(1298) <= layer2_outputs(3820);
    layer3_outputs(1299) <= not(layer2_outputs(2521)) or (layer2_outputs(2019));
    layer3_outputs(1300) <= not((layer2_outputs(3517)) or (layer2_outputs(2326)));
    layer3_outputs(1301) <= '0';
    layer3_outputs(1302) <= '1';
    layer3_outputs(1303) <= not(layer2_outputs(1282)) or (layer2_outputs(1695));
    layer3_outputs(1304) <= (layer2_outputs(4238)) and not (layer2_outputs(2450));
    layer3_outputs(1305) <= layer2_outputs(2736);
    layer3_outputs(1306) <= (layer2_outputs(2283)) and (layer2_outputs(1039));
    layer3_outputs(1307) <= (layer2_outputs(4574)) and not (layer2_outputs(2674));
    layer3_outputs(1308) <= '0';
    layer3_outputs(1309) <= (layer2_outputs(1785)) or (layer2_outputs(3393));
    layer3_outputs(1310) <= not(layer2_outputs(761));
    layer3_outputs(1311) <= (layer2_outputs(3122)) xor (layer2_outputs(576));
    layer3_outputs(1312) <= not((layer2_outputs(3442)) or (layer2_outputs(1462)));
    layer3_outputs(1313) <= '1';
    layer3_outputs(1314) <= not(layer2_outputs(4192));
    layer3_outputs(1315) <= not(layer2_outputs(2045)) or (layer2_outputs(3270));
    layer3_outputs(1316) <= not(layer2_outputs(3476)) or (layer2_outputs(3040));
    layer3_outputs(1317) <= not((layer2_outputs(4354)) or (layer2_outputs(2080)));
    layer3_outputs(1318) <= (layer2_outputs(3382)) and not (layer2_outputs(1265));
    layer3_outputs(1319) <= '1';
    layer3_outputs(1320) <= not((layer2_outputs(1522)) or (layer2_outputs(368)));
    layer3_outputs(1321) <= not(layer2_outputs(1415));
    layer3_outputs(1322) <= '0';
    layer3_outputs(1323) <= (layer2_outputs(2051)) and not (layer2_outputs(2895));
    layer3_outputs(1324) <= not((layer2_outputs(4204)) and (layer2_outputs(4087)));
    layer3_outputs(1325) <= '1';
    layer3_outputs(1326) <= (layer2_outputs(298)) and (layer2_outputs(3858));
    layer3_outputs(1327) <= not(layer2_outputs(4608)) or (layer2_outputs(4048));
    layer3_outputs(1328) <= not((layer2_outputs(1335)) and (layer2_outputs(370)));
    layer3_outputs(1329) <= not(layer2_outputs(3296)) or (layer2_outputs(1701));
    layer3_outputs(1330) <= layer2_outputs(1941);
    layer3_outputs(1331) <= '0';
    layer3_outputs(1332) <= (layer2_outputs(1342)) and (layer2_outputs(2128));
    layer3_outputs(1333) <= not((layer2_outputs(2364)) and (layer2_outputs(4448)));
    layer3_outputs(1334) <= not(layer2_outputs(1420)) or (layer2_outputs(4733));
    layer3_outputs(1335) <= not(layer2_outputs(3486)) or (layer2_outputs(1633));
    layer3_outputs(1336) <= (layer2_outputs(871)) or (layer2_outputs(1217));
    layer3_outputs(1337) <= not(layer2_outputs(4232)) or (layer2_outputs(2449));
    layer3_outputs(1338) <= (layer2_outputs(2867)) and not (layer2_outputs(2714));
    layer3_outputs(1339) <= (layer2_outputs(3852)) and (layer2_outputs(1893));
    layer3_outputs(1340) <= not(layer2_outputs(907));
    layer3_outputs(1341) <= (layer2_outputs(2916)) and not (layer2_outputs(2611));
    layer3_outputs(1342) <= not(layer2_outputs(1437)) or (layer2_outputs(2458));
    layer3_outputs(1343) <= not(layer2_outputs(1187));
    layer3_outputs(1344) <= not(layer2_outputs(4399)) or (layer2_outputs(1126));
    layer3_outputs(1345) <= not((layer2_outputs(152)) or (layer2_outputs(700)));
    layer3_outputs(1346) <= layer2_outputs(4715);
    layer3_outputs(1347) <= (layer2_outputs(4660)) and not (layer2_outputs(1955));
    layer3_outputs(1348) <= (layer2_outputs(167)) and not (layer2_outputs(3294));
    layer3_outputs(1349) <= (layer2_outputs(1942)) or (layer2_outputs(1557));
    layer3_outputs(1350) <= not(layer2_outputs(3636));
    layer3_outputs(1351) <= not((layer2_outputs(3957)) and (layer2_outputs(4956)));
    layer3_outputs(1352) <= '1';
    layer3_outputs(1353) <= layer2_outputs(312);
    layer3_outputs(1354) <= '1';
    layer3_outputs(1355) <= (layer2_outputs(3986)) or (layer2_outputs(3541));
    layer3_outputs(1356) <= not(layer2_outputs(1598)) or (layer2_outputs(1341));
    layer3_outputs(1357) <= (layer2_outputs(3687)) and not (layer2_outputs(4329));
    layer3_outputs(1358) <= not(layer2_outputs(3567));
    layer3_outputs(1359) <= (layer2_outputs(3406)) and not (layer2_outputs(2200));
    layer3_outputs(1360) <= layer2_outputs(2791);
    layer3_outputs(1361) <= not(layer2_outputs(3549));
    layer3_outputs(1362) <= '0';
    layer3_outputs(1363) <= not(layer2_outputs(4174)) or (layer2_outputs(2142));
    layer3_outputs(1364) <= layer2_outputs(1142);
    layer3_outputs(1365) <= not(layer2_outputs(3682));
    layer3_outputs(1366) <= layer2_outputs(1659);
    layer3_outputs(1367) <= '1';
    layer3_outputs(1368) <= '0';
    layer3_outputs(1369) <= (layer2_outputs(4260)) and (layer2_outputs(1264));
    layer3_outputs(1370) <= (layer2_outputs(2847)) and not (layer2_outputs(2354));
    layer3_outputs(1371) <= not((layer2_outputs(479)) or (layer2_outputs(3868)));
    layer3_outputs(1372) <= (layer2_outputs(4422)) and not (layer2_outputs(1758));
    layer3_outputs(1373) <= not(layer2_outputs(2231)) or (layer2_outputs(1706));
    layer3_outputs(1374) <= '1';
    layer3_outputs(1375) <= '0';
    layer3_outputs(1376) <= not((layer2_outputs(422)) or (layer2_outputs(4873)));
    layer3_outputs(1377) <= not(layer2_outputs(21)) or (layer2_outputs(1713));
    layer3_outputs(1378) <= (layer2_outputs(2402)) and not (layer2_outputs(714));
    layer3_outputs(1379) <= not((layer2_outputs(1067)) and (layer2_outputs(1409)));
    layer3_outputs(1380) <= not((layer2_outputs(2844)) and (layer2_outputs(76)));
    layer3_outputs(1381) <= (layer2_outputs(350)) or (layer2_outputs(4348));
    layer3_outputs(1382) <= not((layer2_outputs(3375)) or (layer2_outputs(2623)));
    layer3_outputs(1383) <= '1';
    layer3_outputs(1384) <= not(layer2_outputs(3345)) or (layer2_outputs(480));
    layer3_outputs(1385) <= '0';
    layer3_outputs(1386) <= not((layer2_outputs(4550)) or (layer2_outputs(1293)));
    layer3_outputs(1387) <= not((layer2_outputs(2928)) or (layer2_outputs(2380)));
    layer3_outputs(1388) <= layer2_outputs(2789);
    layer3_outputs(1389) <= not((layer2_outputs(1767)) and (layer2_outputs(2888)));
    layer3_outputs(1390) <= (layer2_outputs(1562)) xor (layer2_outputs(1731));
    layer3_outputs(1391) <= layer2_outputs(1366);
    layer3_outputs(1392) <= '1';
    layer3_outputs(1393) <= (layer2_outputs(1335)) and not (layer2_outputs(2509));
    layer3_outputs(1394) <= (layer2_outputs(542)) and not (layer2_outputs(347));
    layer3_outputs(1395) <= (layer2_outputs(1083)) and not (layer2_outputs(1113));
    layer3_outputs(1396) <= (layer2_outputs(2584)) or (layer2_outputs(1558));
    layer3_outputs(1397) <= not((layer2_outputs(2539)) and (layer2_outputs(3542)));
    layer3_outputs(1398) <= not((layer2_outputs(3122)) and (layer2_outputs(4249)));
    layer3_outputs(1399) <= (layer2_outputs(3188)) and not (layer2_outputs(4294));
    layer3_outputs(1400) <= (layer2_outputs(2230)) or (layer2_outputs(559));
    layer3_outputs(1401) <= layer2_outputs(3845);
    layer3_outputs(1402) <= (layer2_outputs(5057)) and not (layer2_outputs(784));
    layer3_outputs(1403) <= layer2_outputs(2137);
    layer3_outputs(1404) <= '0';
    layer3_outputs(1405) <= (layer2_outputs(172)) and not (layer2_outputs(1896));
    layer3_outputs(1406) <= not((layer2_outputs(1073)) or (layer2_outputs(2757)));
    layer3_outputs(1407) <= (layer2_outputs(4249)) or (layer2_outputs(1431));
    layer3_outputs(1408) <= '0';
    layer3_outputs(1409) <= not(layer2_outputs(2724));
    layer3_outputs(1410) <= (layer2_outputs(2536)) and (layer2_outputs(634));
    layer3_outputs(1411) <= (layer2_outputs(2514)) or (layer2_outputs(1184));
    layer3_outputs(1412) <= not(layer2_outputs(3400)) or (layer2_outputs(3958));
    layer3_outputs(1413) <= (layer2_outputs(584)) and not (layer2_outputs(1817));
    layer3_outputs(1414) <= not(layer2_outputs(1487));
    layer3_outputs(1415) <= not(layer2_outputs(2336));
    layer3_outputs(1416) <= (layer2_outputs(3603)) and not (layer2_outputs(4667));
    layer3_outputs(1417) <= not(layer2_outputs(4823));
    layer3_outputs(1418) <= '1';
    layer3_outputs(1419) <= not(layer2_outputs(4003));
    layer3_outputs(1420) <= not((layer2_outputs(2889)) or (layer2_outputs(816)));
    layer3_outputs(1421) <= not(layer2_outputs(12)) or (layer2_outputs(4157));
    layer3_outputs(1422) <= not((layer2_outputs(817)) xor (layer2_outputs(2677)));
    layer3_outputs(1423) <= (layer2_outputs(4391)) xor (layer2_outputs(4124));
    layer3_outputs(1424) <= (layer2_outputs(2828)) or (layer2_outputs(40));
    layer3_outputs(1425) <= not(layer2_outputs(837)) or (layer2_outputs(3935));
    layer3_outputs(1426) <= not(layer2_outputs(3876)) or (layer2_outputs(1955));
    layer3_outputs(1427) <= (layer2_outputs(3950)) and (layer2_outputs(2983));
    layer3_outputs(1428) <= not(layer2_outputs(3743)) or (layer2_outputs(2289));
    layer3_outputs(1429) <= (layer2_outputs(4690)) xor (layer2_outputs(4725));
    layer3_outputs(1430) <= '1';
    layer3_outputs(1431) <= layer2_outputs(4230);
    layer3_outputs(1432) <= '1';
    layer3_outputs(1433) <= '1';
    layer3_outputs(1434) <= (layer2_outputs(2947)) and not (layer2_outputs(620));
    layer3_outputs(1435) <= not(layer2_outputs(2502)) or (layer2_outputs(2840));
    layer3_outputs(1436) <= '1';
    layer3_outputs(1437) <= layer2_outputs(381);
    layer3_outputs(1438) <= layer2_outputs(4547);
    layer3_outputs(1439) <= not(layer2_outputs(3044)) or (layer2_outputs(2343));
    layer3_outputs(1440) <= '0';
    layer3_outputs(1441) <= '1';
    layer3_outputs(1442) <= '0';
    layer3_outputs(1443) <= not(layer2_outputs(3500));
    layer3_outputs(1444) <= (layer2_outputs(4180)) and not (layer2_outputs(1413));
    layer3_outputs(1445) <= (layer2_outputs(3970)) and not (layer2_outputs(690));
    layer3_outputs(1446) <= '1';
    layer3_outputs(1447) <= (layer2_outputs(2717)) and (layer2_outputs(5101));
    layer3_outputs(1448) <= layer2_outputs(1178);
    layer3_outputs(1449) <= not(layer2_outputs(590)) or (layer2_outputs(3426));
    layer3_outputs(1450) <= layer2_outputs(68);
    layer3_outputs(1451) <= (layer2_outputs(725)) or (layer2_outputs(1825));
    layer3_outputs(1452) <= not((layer2_outputs(528)) or (layer2_outputs(3002)));
    layer3_outputs(1453) <= '0';
    layer3_outputs(1454) <= (layer2_outputs(4701)) or (layer2_outputs(1684));
    layer3_outputs(1455) <= (layer2_outputs(4879)) and not (layer2_outputs(5061));
    layer3_outputs(1456) <= layer2_outputs(1051);
    layer3_outputs(1457) <= '0';
    layer3_outputs(1458) <= not((layer2_outputs(4383)) xor (layer2_outputs(3209)));
    layer3_outputs(1459) <= (layer2_outputs(1165)) and not (layer2_outputs(305));
    layer3_outputs(1460) <= '0';
    layer3_outputs(1461) <= not((layer2_outputs(105)) or (layer2_outputs(4241)));
    layer3_outputs(1462) <= not(layer2_outputs(2565)) or (layer2_outputs(93));
    layer3_outputs(1463) <= layer2_outputs(4483);
    layer3_outputs(1464) <= not((layer2_outputs(4071)) or (layer2_outputs(1067)));
    layer3_outputs(1465) <= (layer2_outputs(2595)) and not (layer2_outputs(1150));
    layer3_outputs(1466) <= layer2_outputs(816);
    layer3_outputs(1467) <= '0';
    layer3_outputs(1468) <= (layer2_outputs(1551)) and not (layer2_outputs(2477));
    layer3_outputs(1469) <= (layer2_outputs(2497)) and not (layer2_outputs(4064));
    layer3_outputs(1470) <= (layer2_outputs(3931)) or (layer2_outputs(4594));
    layer3_outputs(1471) <= not((layer2_outputs(657)) or (layer2_outputs(2337)));
    layer3_outputs(1472) <= not(layer2_outputs(3153)) or (layer2_outputs(224));
    layer3_outputs(1473) <= (layer2_outputs(4590)) and not (layer2_outputs(3645));
    layer3_outputs(1474) <= not(layer2_outputs(4386));
    layer3_outputs(1475) <= not(layer2_outputs(3853)) or (layer2_outputs(2212));
    layer3_outputs(1476) <= layer2_outputs(3651);
    layer3_outputs(1477) <= '0';
    layer3_outputs(1478) <= (layer2_outputs(600)) and (layer2_outputs(2533));
    layer3_outputs(1479) <= not((layer2_outputs(789)) xor (layer2_outputs(2986)));
    layer3_outputs(1480) <= '1';
    layer3_outputs(1481) <= (layer2_outputs(2462)) and not (layer2_outputs(3567));
    layer3_outputs(1482) <= (layer2_outputs(1657)) or (layer2_outputs(1801));
    layer3_outputs(1483) <= (layer2_outputs(1673)) and not (layer2_outputs(4468));
    layer3_outputs(1484) <= layer2_outputs(4018);
    layer3_outputs(1485) <= not(layer2_outputs(1357)) or (layer2_outputs(3726));
    layer3_outputs(1486) <= not(layer2_outputs(116));
    layer3_outputs(1487) <= not(layer2_outputs(2807));
    layer3_outputs(1488) <= layer2_outputs(3911);
    layer3_outputs(1489) <= not(layer2_outputs(666));
    layer3_outputs(1490) <= not(layer2_outputs(814));
    layer3_outputs(1491) <= layer2_outputs(1016);
    layer3_outputs(1492) <= layer2_outputs(3146);
    layer3_outputs(1493) <= layer2_outputs(4713);
    layer3_outputs(1494) <= layer2_outputs(2052);
    layer3_outputs(1495) <= not(layer2_outputs(3954)) or (layer2_outputs(579));
    layer3_outputs(1496) <= (layer2_outputs(2651)) and (layer2_outputs(1077));
    layer3_outputs(1497) <= not(layer2_outputs(962)) or (layer2_outputs(3990));
    layer3_outputs(1498) <= not(layer2_outputs(3374));
    layer3_outputs(1499) <= layer2_outputs(4849);
    layer3_outputs(1500) <= '1';
    layer3_outputs(1501) <= not((layer2_outputs(2491)) or (layer2_outputs(1356)));
    layer3_outputs(1502) <= '0';
    layer3_outputs(1503) <= not(layer2_outputs(4035)) or (layer2_outputs(325));
    layer3_outputs(1504) <= (layer2_outputs(4355)) or (layer2_outputs(2253));
    layer3_outputs(1505) <= not(layer2_outputs(4197)) or (layer2_outputs(2839));
    layer3_outputs(1506) <= not(layer2_outputs(595));
    layer3_outputs(1507) <= '1';
    layer3_outputs(1508) <= not((layer2_outputs(3485)) and (layer2_outputs(5002)));
    layer3_outputs(1509) <= not((layer2_outputs(2199)) or (layer2_outputs(132)));
    layer3_outputs(1510) <= (layer2_outputs(1621)) xor (layer2_outputs(446));
    layer3_outputs(1511) <= '1';
    layer3_outputs(1512) <= (layer2_outputs(3585)) and not (layer2_outputs(4641));
    layer3_outputs(1513) <= (layer2_outputs(3871)) or (layer2_outputs(1284));
    layer3_outputs(1514) <= (layer2_outputs(2863)) and not (layer2_outputs(272));
    layer3_outputs(1515) <= layer2_outputs(1660);
    layer3_outputs(1516) <= not(layer2_outputs(3767)) or (layer2_outputs(2681));
    layer3_outputs(1517) <= (layer2_outputs(4441)) and not (layer2_outputs(3600));
    layer3_outputs(1518) <= not(layer2_outputs(1924)) or (layer2_outputs(1421));
    layer3_outputs(1519) <= not(layer2_outputs(3134)) or (layer2_outputs(2573));
    layer3_outputs(1520) <= not(layer2_outputs(3879));
    layer3_outputs(1521) <= '0';
    layer3_outputs(1522) <= not((layer2_outputs(60)) or (layer2_outputs(4543)));
    layer3_outputs(1523) <= not(layer2_outputs(2505)) or (layer2_outputs(3835));
    layer3_outputs(1524) <= not((layer2_outputs(2384)) and (layer2_outputs(31)));
    layer3_outputs(1525) <= (layer2_outputs(2546)) and not (layer2_outputs(871));
    layer3_outputs(1526) <= '0';
    layer3_outputs(1527) <= '0';
    layer3_outputs(1528) <= not(layer2_outputs(2950));
    layer3_outputs(1529) <= not((layer2_outputs(851)) and (layer2_outputs(442)));
    layer3_outputs(1530) <= '0';
    layer3_outputs(1531) <= (layer2_outputs(4940)) and (layer2_outputs(3954));
    layer3_outputs(1532) <= not(layer2_outputs(4358)) or (layer2_outputs(3393));
    layer3_outputs(1533) <= '1';
    layer3_outputs(1534) <= not(layer2_outputs(435)) or (layer2_outputs(463));
    layer3_outputs(1535) <= '0';
    layer3_outputs(1536) <= '0';
    layer3_outputs(1537) <= not(layer2_outputs(2399)) or (layer2_outputs(4352));
    layer3_outputs(1538) <= not(layer2_outputs(2856));
    layer3_outputs(1539) <= (layer2_outputs(1655)) and (layer2_outputs(156));
    layer3_outputs(1540) <= not((layer2_outputs(69)) and (layer2_outputs(2393)));
    layer3_outputs(1541) <= not(layer2_outputs(3892));
    layer3_outputs(1542) <= (layer2_outputs(4288)) and (layer2_outputs(3095));
    layer3_outputs(1543) <= layer2_outputs(1968);
    layer3_outputs(1544) <= '0';
    layer3_outputs(1545) <= (layer2_outputs(3695)) and not (layer2_outputs(4177));
    layer3_outputs(1546) <= not(layer2_outputs(601));
    layer3_outputs(1547) <= not(layer2_outputs(1633));
    layer3_outputs(1548) <= not(layer2_outputs(1766)) or (layer2_outputs(2756));
    layer3_outputs(1549) <= (layer2_outputs(1725)) and not (layer2_outputs(1103));
    layer3_outputs(1550) <= layer2_outputs(1632);
    layer3_outputs(1551) <= (layer2_outputs(4429)) or (layer2_outputs(3680));
    layer3_outputs(1552) <= layer2_outputs(1897);
    layer3_outputs(1553) <= (layer2_outputs(3136)) or (layer2_outputs(1472));
    layer3_outputs(1554) <= (layer2_outputs(3308)) and (layer2_outputs(3117));
    layer3_outputs(1555) <= layer2_outputs(2305);
    layer3_outputs(1556) <= '1';
    layer3_outputs(1557) <= layer2_outputs(914);
    layer3_outputs(1558) <= layer2_outputs(2291);
    layer3_outputs(1559) <= not((layer2_outputs(2302)) or (layer2_outputs(2565)));
    layer3_outputs(1560) <= '0';
    layer3_outputs(1561) <= not(layer2_outputs(2585)) or (layer2_outputs(513));
    layer3_outputs(1562) <= (layer2_outputs(4983)) or (layer2_outputs(3925));
    layer3_outputs(1563) <= '0';
    layer3_outputs(1564) <= (layer2_outputs(1494)) and not (layer2_outputs(237));
    layer3_outputs(1565) <= (layer2_outputs(3422)) and not (layer2_outputs(44));
    layer3_outputs(1566) <= not((layer2_outputs(5045)) and (layer2_outputs(2993)));
    layer3_outputs(1567) <= '0';
    layer3_outputs(1568) <= (layer2_outputs(1393)) or (layer2_outputs(474));
    layer3_outputs(1569) <= layer2_outputs(302);
    layer3_outputs(1570) <= not(layer2_outputs(10)) or (layer2_outputs(4185));
    layer3_outputs(1571) <= not(layer2_outputs(2487));
    layer3_outputs(1572) <= not((layer2_outputs(4949)) or (layer2_outputs(3025)));
    layer3_outputs(1573) <= layer2_outputs(453);
    layer3_outputs(1574) <= not(layer2_outputs(338)) or (layer2_outputs(5060));
    layer3_outputs(1575) <= '0';
    layer3_outputs(1576) <= not((layer2_outputs(1307)) xor (layer2_outputs(4167)));
    layer3_outputs(1577) <= (layer2_outputs(2790)) or (layer2_outputs(183));
    layer3_outputs(1578) <= layer2_outputs(529);
    layer3_outputs(1579) <= (layer2_outputs(4883)) and not (layer2_outputs(3872));
    layer3_outputs(1580) <= not(layer2_outputs(5109)) or (layer2_outputs(619));
    layer3_outputs(1581) <= not((layer2_outputs(1783)) and (layer2_outputs(2372)));
    layer3_outputs(1582) <= (layer2_outputs(1228)) and not (layer2_outputs(4961));
    layer3_outputs(1583) <= layer2_outputs(241);
    layer3_outputs(1584) <= not((layer2_outputs(5068)) xor (layer2_outputs(4862)));
    layer3_outputs(1585) <= '0';
    layer3_outputs(1586) <= not((layer2_outputs(367)) or (layer2_outputs(2130)));
    layer3_outputs(1587) <= not((layer2_outputs(2759)) and (layer2_outputs(3746)));
    layer3_outputs(1588) <= layer2_outputs(2765);
    layer3_outputs(1589) <= not(layer2_outputs(4956)) or (layer2_outputs(4253));
    layer3_outputs(1590) <= not((layer2_outputs(3268)) or (layer2_outputs(2901)));
    layer3_outputs(1591) <= not((layer2_outputs(1792)) or (layer2_outputs(3142)));
    layer3_outputs(1592) <= layer2_outputs(3376);
    layer3_outputs(1593) <= not(layer2_outputs(1847));
    layer3_outputs(1594) <= layer2_outputs(4463);
    layer3_outputs(1595) <= (layer2_outputs(324)) and not (layer2_outputs(2615));
    layer3_outputs(1596) <= (layer2_outputs(370)) and not (layer2_outputs(103));
    layer3_outputs(1597) <= not(layer2_outputs(2632)) or (layer2_outputs(4516));
    layer3_outputs(1598) <= not(layer2_outputs(5080)) or (layer2_outputs(426));
    layer3_outputs(1599) <= not(layer2_outputs(2828)) or (layer2_outputs(1309));
    layer3_outputs(1600) <= (layer2_outputs(3021)) and (layer2_outputs(3989));
    layer3_outputs(1601) <= (layer2_outputs(3071)) and (layer2_outputs(1382));
    layer3_outputs(1602) <= not((layer2_outputs(3920)) and (layer2_outputs(1640)));
    layer3_outputs(1603) <= '0';
    layer3_outputs(1604) <= '0';
    layer3_outputs(1605) <= not(layer2_outputs(4306)) or (layer2_outputs(2963));
    layer3_outputs(1606) <= (layer2_outputs(2548)) and not (layer2_outputs(3821));
    layer3_outputs(1607) <= not(layer2_outputs(1198));
    layer3_outputs(1608) <= not(layer2_outputs(209));
    layer3_outputs(1609) <= not(layer2_outputs(379));
    layer3_outputs(1610) <= (layer2_outputs(2783)) or (layer2_outputs(3533));
    layer3_outputs(1611) <= (layer2_outputs(4901)) and not (layer2_outputs(3974));
    layer3_outputs(1612) <= layer2_outputs(1845);
    layer3_outputs(1613) <= '1';
    layer3_outputs(1614) <= '1';
    layer3_outputs(1615) <= (layer2_outputs(2279)) and (layer2_outputs(60));
    layer3_outputs(1616) <= layer2_outputs(2156);
    layer3_outputs(1617) <= not((layer2_outputs(4417)) and (layer2_outputs(3605)));
    layer3_outputs(1618) <= layer2_outputs(2155);
    layer3_outputs(1619) <= (layer2_outputs(1317)) and (layer2_outputs(4643));
    layer3_outputs(1620) <= layer2_outputs(4423);
    layer3_outputs(1621) <= not((layer2_outputs(3128)) and (layer2_outputs(2604)));
    layer3_outputs(1622) <= not(layer2_outputs(2636)) or (layer2_outputs(715));
    layer3_outputs(1623) <= not(layer2_outputs(3976)) or (layer2_outputs(3407));
    layer3_outputs(1624) <= (layer2_outputs(3734)) or (layer2_outputs(4434));
    layer3_outputs(1625) <= (layer2_outputs(1289)) and (layer2_outputs(1778));
    layer3_outputs(1626) <= not(layer2_outputs(2353));
    layer3_outputs(1627) <= (layer2_outputs(4026)) and not (layer2_outputs(1125));
    layer3_outputs(1628) <= layer2_outputs(3525);
    layer3_outputs(1629) <= '1';
    layer3_outputs(1630) <= not(layer2_outputs(3151));
    layer3_outputs(1631) <= '0';
    layer3_outputs(1632) <= (layer2_outputs(524)) and (layer2_outputs(2851));
    layer3_outputs(1633) <= layer2_outputs(4520);
    layer3_outputs(1634) <= layer2_outputs(2949);
    layer3_outputs(1635) <= (layer2_outputs(3786)) or (layer2_outputs(2177));
    layer3_outputs(1636) <= not(layer2_outputs(3462)) or (layer2_outputs(2559));
    layer3_outputs(1637) <= not(layer2_outputs(2091));
    layer3_outputs(1638) <= layer2_outputs(2091);
    layer3_outputs(1639) <= not(layer2_outputs(3715));
    layer3_outputs(1640) <= '0';
    layer3_outputs(1641) <= '0';
    layer3_outputs(1642) <= '1';
    layer3_outputs(1643) <= (layer2_outputs(4831)) and (layer2_outputs(2985));
    layer3_outputs(1644) <= not((layer2_outputs(3449)) and (layer2_outputs(1612)));
    layer3_outputs(1645) <= layer2_outputs(1369);
    layer3_outputs(1646) <= (layer2_outputs(2371)) and not (layer2_outputs(2776));
    layer3_outputs(1647) <= (layer2_outputs(2217)) and not (layer2_outputs(1150));
    layer3_outputs(1648) <= (layer2_outputs(2794)) or (layer2_outputs(2470));
    layer3_outputs(1649) <= layer2_outputs(3698);
    layer3_outputs(1650) <= not(layer2_outputs(2775));
    layer3_outputs(1651) <= (layer2_outputs(3021)) and (layer2_outputs(1882));
    layer3_outputs(1652) <= not(layer2_outputs(1047));
    layer3_outputs(1653) <= (layer2_outputs(3602)) or (layer2_outputs(4364));
    layer3_outputs(1654) <= not((layer2_outputs(1059)) and (layer2_outputs(3633)));
    layer3_outputs(1655) <= '0';
    layer3_outputs(1656) <= layer2_outputs(832);
    layer3_outputs(1657) <= (layer2_outputs(2506)) or (layer2_outputs(2886));
    layer3_outputs(1658) <= layer2_outputs(45);
    layer3_outputs(1659) <= not(layer2_outputs(2186));
    layer3_outputs(1660) <= '1';
    layer3_outputs(1661) <= not(layer2_outputs(1127)) or (layer2_outputs(925));
    layer3_outputs(1662) <= (layer2_outputs(4755)) and not (layer2_outputs(3639));
    layer3_outputs(1663) <= (layer2_outputs(3482)) xor (layer2_outputs(1868));
    layer3_outputs(1664) <= not((layer2_outputs(464)) xor (layer2_outputs(1834)));
    layer3_outputs(1665) <= not(layer2_outputs(1805)) or (layer2_outputs(4595));
    layer3_outputs(1666) <= (layer2_outputs(3)) and not (layer2_outputs(314));
    layer3_outputs(1667) <= (layer2_outputs(1525)) and (layer2_outputs(3659));
    layer3_outputs(1668) <= not(layer2_outputs(749)) or (layer2_outputs(3058));
    layer3_outputs(1669) <= (layer2_outputs(2001)) and not (layer2_outputs(3917));
    layer3_outputs(1670) <= (layer2_outputs(3891)) and not (layer2_outputs(2381));
    layer3_outputs(1671) <= (layer2_outputs(4768)) and not (layer2_outputs(3176));
    layer3_outputs(1672) <= (layer2_outputs(2682)) or (layer2_outputs(2370));
    layer3_outputs(1673) <= (layer2_outputs(4568)) and not (layer2_outputs(4866));
    layer3_outputs(1674) <= (layer2_outputs(3889)) and not (layer2_outputs(3703));
    layer3_outputs(1675) <= '0';
    layer3_outputs(1676) <= layer2_outputs(3443);
    layer3_outputs(1677) <= not((layer2_outputs(4514)) and (layer2_outputs(1979)));
    layer3_outputs(1678) <= not(layer2_outputs(3640));
    layer3_outputs(1679) <= layer2_outputs(1893);
    layer3_outputs(1680) <= layer2_outputs(3800);
    layer3_outputs(1681) <= not(layer2_outputs(4511));
    layer3_outputs(1682) <= (layer2_outputs(1081)) and (layer2_outputs(4995));
    layer3_outputs(1683) <= not((layer2_outputs(2269)) and (layer2_outputs(1538)));
    layer3_outputs(1684) <= (layer2_outputs(4763)) xor (layer2_outputs(4630));
    layer3_outputs(1685) <= (layer2_outputs(1006)) and not (layer2_outputs(2730));
    layer3_outputs(1686) <= layer2_outputs(2233);
    layer3_outputs(1687) <= not(layer2_outputs(2427));
    layer3_outputs(1688) <= not((layer2_outputs(2564)) or (layer2_outputs(125)));
    layer3_outputs(1689) <= (layer2_outputs(3339)) and not (layer2_outputs(1867));
    layer3_outputs(1690) <= (layer2_outputs(4884)) and not (layer2_outputs(1704));
    layer3_outputs(1691) <= not((layer2_outputs(394)) and (layer2_outputs(676)));
    layer3_outputs(1692) <= (layer2_outputs(3596)) and not (layer2_outputs(934));
    layer3_outputs(1693) <= not(layer2_outputs(2116)) or (layer2_outputs(1520));
    layer3_outputs(1694) <= not(layer2_outputs(3033));
    layer3_outputs(1695) <= not(layer2_outputs(1325));
    layer3_outputs(1696) <= '0';
    layer3_outputs(1697) <= '0';
    layer3_outputs(1698) <= not((layer2_outputs(4321)) xor (layer2_outputs(3374)));
    layer3_outputs(1699) <= (layer2_outputs(1087)) and (layer2_outputs(4801));
    layer3_outputs(1700) <= '1';
    layer3_outputs(1701) <= not(layer2_outputs(583));
    layer3_outputs(1702) <= (layer2_outputs(4438)) and not (layer2_outputs(3096));
    layer3_outputs(1703) <= layer2_outputs(1055);
    layer3_outputs(1704) <= layer2_outputs(346);
    layer3_outputs(1705) <= (layer2_outputs(2400)) and not (layer2_outputs(3719));
    layer3_outputs(1706) <= not(layer2_outputs(2939)) or (layer2_outputs(3075));
    layer3_outputs(1707) <= not(layer2_outputs(3450));
    layer3_outputs(1708) <= '0';
    layer3_outputs(1709) <= layer2_outputs(2168);
    layer3_outputs(1710) <= not(layer2_outputs(4652));
    layer3_outputs(1711) <= not(layer2_outputs(315)) or (layer2_outputs(1002));
    layer3_outputs(1712) <= '1';
    layer3_outputs(1713) <= not(layer2_outputs(4623)) or (layer2_outputs(2782));
    layer3_outputs(1714) <= layer2_outputs(3923);
    layer3_outputs(1715) <= '1';
    layer3_outputs(1716) <= (layer2_outputs(4941)) and not (layer2_outputs(552));
    layer3_outputs(1717) <= (layer2_outputs(759)) and not (layer2_outputs(1064));
    layer3_outputs(1718) <= not((layer2_outputs(4943)) and (layer2_outputs(4288)));
    layer3_outputs(1719) <= (layer2_outputs(629)) and not (layer2_outputs(3119));
    layer3_outputs(1720) <= not(layer2_outputs(2069)) or (layer2_outputs(4130));
    layer3_outputs(1721) <= layer2_outputs(77);
    layer3_outputs(1722) <= (layer2_outputs(406)) or (layer2_outputs(1770));
    layer3_outputs(1723) <= layer2_outputs(1302);
    layer3_outputs(1724) <= not((layer2_outputs(4683)) or (layer2_outputs(501)));
    layer3_outputs(1725) <= (layer2_outputs(1465)) and (layer2_outputs(3577));
    layer3_outputs(1726) <= (layer2_outputs(1686)) and (layer2_outputs(465));
    layer3_outputs(1727) <= '1';
    layer3_outputs(1728) <= (layer2_outputs(676)) xor (layer2_outputs(4262));
    layer3_outputs(1729) <= not((layer2_outputs(3227)) or (layer2_outputs(4797)));
    layer3_outputs(1730) <= not(layer2_outputs(1562));
    layer3_outputs(1731) <= (layer2_outputs(3161)) xor (layer2_outputs(3222));
    layer3_outputs(1732) <= not(layer2_outputs(1560));
    layer3_outputs(1733) <= not(layer2_outputs(1248));
    layer3_outputs(1734) <= not(layer2_outputs(3761));
    layer3_outputs(1735) <= not(layer2_outputs(1858));
    layer3_outputs(1736) <= not(layer2_outputs(617));
    layer3_outputs(1737) <= '1';
    layer3_outputs(1738) <= (layer2_outputs(4054)) and (layer2_outputs(4163));
    layer3_outputs(1739) <= '1';
    layer3_outputs(1740) <= layer2_outputs(429);
    layer3_outputs(1741) <= not((layer2_outputs(3561)) or (layer2_outputs(2769)));
    layer3_outputs(1742) <= '0';
    layer3_outputs(1743) <= (layer2_outputs(1888)) or (layer2_outputs(3575));
    layer3_outputs(1744) <= not((layer2_outputs(3994)) or (layer2_outputs(3642)));
    layer3_outputs(1745) <= (layer2_outputs(2322)) and not (layer2_outputs(2752));
    layer3_outputs(1746) <= not((layer2_outputs(1143)) or (layer2_outputs(540)));
    layer3_outputs(1747) <= layer2_outputs(2938);
    layer3_outputs(1748) <= (layer2_outputs(3537)) and not (layer2_outputs(3896));
    layer3_outputs(1749) <= (layer2_outputs(3079)) and not (layer2_outputs(336));
    layer3_outputs(1750) <= layer2_outputs(2292);
    layer3_outputs(1751) <= not((layer2_outputs(4398)) and (layer2_outputs(1596)));
    layer3_outputs(1752) <= not(layer2_outputs(1544)) or (layer2_outputs(3314));
    layer3_outputs(1753) <= not((layer2_outputs(997)) and (layer2_outputs(3428)));
    layer3_outputs(1754) <= (layer2_outputs(912)) and not (layer2_outputs(227));
    layer3_outputs(1755) <= not((layer2_outputs(3854)) or (layer2_outputs(2709)));
    layer3_outputs(1756) <= (layer2_outputs(2853)) xor (layer2_outputs(904));
    layer3_outputs(1757) <= not((layer2_outputs(3997)) or (layer2_outputs(2969)));
    layer3_outputs(1758) <= not(layer2_outputs(3204)) or (layer2_outputs(4942));
    layer3_outputs(1759) <= '0';
    layer3_outputs(1760) <= not(layer2_outputs(4730)) or (layer2_outputs(167));
    layer3_outputs(1761) <= '1';
    layer3_outputs(1762) <= not(layer2_outputs(1961)) or (layer2_outputs(2123));
    layer3_outputs(1763) <= (layer2_outputs(4326)) and (layer2_outputs(2909));
    layer3_outputs(1764) <= layer2_outputs(3369);
    layer3_outputs(1765) <= (layer2_outputs(539)) or (layer2_outputs(3598));
    layer3_outputs(1766) <= not(layer2_outputs(4296)) or (layer2_outputs(2551));
    layer3_outputs(1767) <= '1';
    layer3_outputs(1768) <= not(layer2_outputs(5111));
    layer3_outputs(1769) <= layer2_outputs(1442);
    layer3_outputs(1770) <= '0';
    layer3_outputs(1771) <= not(layer2_outputs(3154)) or (layer2_outputs(4586));
    layer3_outputs(1772) <= (layer2_outputs(3993)) and not (layer2_outputs(206));
    layer3_outputs(1773) <= (layer2_outputs(2081)) and not (layer2_outputs(4439));
    layer3_outputs(1774) <= (layer2_outputs(3884)) or (layer2_outputs(157));
    layer3_outputs(1775) <= layer2_outputs(30);
    layer3_outputs(1776) <= '1';
    layer3_outputs(1777) <= not(layer2_outputs(4495));
    layer3_outputs(1778) <= not(layer2_outputs(3036)) or (layer2_outputs(1522));
    layer3_outputs(1779) <= layer2_outputs(3168);
    layer3_outputs(1780) <= not(layer2_outputs(2644));
    layer3_outputs(1781) <= not((layer2_outputs(1114)) or (layer2_outputs(3806)));
    layer3_outputs(1782) <= not((layer2_outputs(774)) xor (layer2_outputs(2678)));
    layer3_outputs(1783) <= '1';
    layer3_outputs(1784) <= (layer2_outputs(4617)) and not (layer2_outputs(396));
    layer3_outputs(1785) <= '0';
    layer3_outputs(1786) <= (layer2_outputs(2164)) and (layer2_outputs(2180));
    layer3_outputs(1787) <= '1';
    layer3_outputs(1788) <= not(layer2_outputs(162)) or (layer2_outputs(1625));
    layer3_outputs(1789) <= (layer2_outputs(1074)) and (layer2_outputs(642));
    layer3_outputs(1790) <= '1';
    layer3_outputs(1791) <= (layer2_outputs(2144)) and not (layer2_outputs(5023));
    layer3_outputs(1792) <= '0';
    layer3_outputs(1793) <= '0';
    layer3_outputs(1794) <= not(layer2_outputs(4440));
    layer3_outputs(1795) <= not(layer2_outputs(4776));
    layer3_outputs(1796) <= (layer2_outputs(2970)) and not (layer2_outputs(3495));
    layer3_outputs(1797) <= layer2_outputs(4456);
    layer3_outputs(1798) <= not(layer2_outputs(506)) or (layer2_outputs(74));
    layer3_outputs(1799) <= (layer2_outputs(3271)) and not (layer2_outputs(3408));
    layer3_outputs(1800) <= layer2_outputs(2110);
    layer3_outputs(1801) <= layer2_outputs(3316);
    layer3_outputs(1802) <= (layer2_outputs(1756)) and (layer2_outputs(2093));
    layer3_outputs(1803) <= not(layer2_outputs(3984)) or (layer2_outputs(2525));
    layer3_outputs(1804) <= layer2_outputs(2203);
    layer3_outputs(1805) <= layer2_outputs(4730);
    layer3_outputs(1806) <= not(layer2_outputs(178)) or (layer2_outputs(865));
    layer3_outputs(1807) <= not((layer2_outputs(3906)) or (layer2_outputs(124)));
    layer3_outputs(1808) <= '0';
    layer3_outputs(1809) <= not(layer2_outputs(4622)) or (layer2_outputs(2441));
    layer3_outputs(1810) <= not(layer2_outputs(3609)) or (layer2_outputs(1056));
    layer3_outputs(1811) <= not(layer2_outputs(365));
    layer3_outputs(1812) <= layer2_outputs(2858);
    layer3_outputs(1813) <= not(layer2_outputs(3544));
    layer3_outputs(1814) <= layer2_outputs(4177);
    layer3_outputs(1815) <= layer2_outputs(3173);
    layer3_outputs(1816) <= not(layer2_outputs(3899));
    layer3_outputs(1817) <= not(layer2_outputs(390)) or (layer2_outputs(3901));
    layer3_outputs(1818) <= not(layer2_outputs(1279));
    layer3_outputs(1819) <= layer2_outputs(2227);
    layer3_outputs(1820) <= not((layer2_outputs(2142)) or (layer2_outputs(3387)));
    layer3_outputs(1821) <= (layer2_outputs(4355)) and not (layer2_outputs(4931));
    layer3_outputs(1822) <= (layer2_outputs(2898)) and (layer2_outputs(2739));
    layer3_outputs(1823) <= not((layer2_outputs(4286)) and (layer2_outputs(2183)));
    layer3_outputs(1824) <= '0';
    layer3_outputs(1825) <= not(layer2_outputs(4217)) or (layer2_outputs(3611));
    layer3_outputs(1826) <= '0';
    layer3_outputs(1827) <= (layer2_outputs(4447)) and not (layer2_outputs(1563));
    layer3_outputs(1828) <= not(layer2_outputs(3231));
    layer3_outputs(1829) <= layer2_outputs(3178);
    layer3_outputs(1830) <= '0';
    layer3_outputs(1831) <= (layer2_outputs(4818)) and not (layer2_outputs(3050));
    layer3_outputs(1832) <= '0';
    layer3_outputs(1833) <= layer2_outputs(1018);
    layer3_outputs(1834) <= layer2_outputs(4977);
    layer3_outputs(1835) <= layer2_outputs(6);
    layer3_outputs(1836) <= '0';
    layer3_outputs(1837) <= not(layer2_outputs(3113)) or (layer2_outputs(4283));
    layer3_outputs(1838) <= not(layer2_outputs(1478));
    layer3_outputs(1839) <= '0';
    layer3_outputs(1840) <= (layer2_outputs(2291)) and (layer2_outputs(578));
    layer3_outputs(1841) <= not(layer2_outputs(4406));
    layer3_outputs(1842) <= '1';
    layer3_outputs(1843) <= '0';
    layer3_outputs(1844) <= layer2_outputs(1756);
    layer3_outputs(1845) <= not((layer2_outputs(2483)) xor (layer2_outputs(4921)));
    layer3_outputs(1846) <= not(layer2_outputs(4617));
    layer3_outputs(1847) <= layer2_outputs(4198);
    layer3_outputs(1848) <= '1';
    layer3_outputs(1849) <= not(layer2_outputs(4674));
    layer3_outputs(1850) <= layer2_outputs(493);
    layer3_outputs(1851) <= layer2_outputs(740);
    layer3_outputs(1852) <= not(layer2_outputs(3364));
    layer3_outputs(1853) <= (layer2_outputs(2172)) and not (layer2_outputs(3483));
    layer3_outputs(1854) <= not(layer2_outputs(3758));
    layer3_outputs(1855) <= (layer2_outputs(869)) and (layer2_outputs(2788));
    layer3_outputs(1856) <= layer2_outputs(273);
    layer3_outputs(1857) <= (layer2_outputs(1171)) and not (layer2_outputs(803));
    layer3_outputs(1858) <= not(layer2_outputs(4998));
    layer3_outputs(1859) <= (layer2_outputs(2255)) and (layer2_outputs(377));
    layer3_outputs(1860) <= not(layer2_outputs(2271));
    layer3_outputs(1861) <= '0';
    layer3_outputs(1862) <= (layer2_outputs(3471)) or (layer2_outputs(79));
    layer3_outputs(1863) <= layer2_outputs(4028);
    layer3_outputs(1864) <= not(layer2_outputs(4792)) or (layer2_outputs(3527));
    layer3_outputs(1865) <= (layer2_outputs(1272)) and (layer2_outputs(1184));
    layer3_outputs(1866) <= not((layer2_outputs(3306)) or (layer2_outputs(893)));
    layer3_outputs(1867) <= '1';
    layer3_outputs(1868) <= (layer2_outputs(2059)) and not (layer2_outputs(451));
    layer3_outputs(1869) <= '0';
    layer3_outputs(1870) <= (layer2_outputs(1745)) or (layer2_outputs(3817));
    layer3_outputs(1871) <= layer2_outputs(3322);
    layer3_outputs(1872) <= '0';
    layer3_outputs(1873) <= (layer2_outputs(4202)) and not (layer2_outputs(1378));
    layer3_outputs(1874) <= not(layer2_outputs(1716)) or (layer2_outputs(2757));
    layer3_outputs(1875) <= layer2_outputs(2915);
    layer3_outputs(1876) <= (layer2_outputs(728)) and (layer2_outputs(3855));
    layer3_outputs(1877) <= (layer2_outputs(3328)) and not (layer2_outputs(4719));
    layer3_outputs(1878) <= '1';
    layer3_outputs(1879) <= not((layer2_outputs(2951)) or (layer2_outputs(2728)));
    layer3_outputs(1880) <= '1';
    layer3_outputs(1881) <= not((layer2_outputs(913)) and (layer2_outputs(3530)));
    layer3_outputs(1882) <= (layer2_outputs(1978)) and not (layer2_outputs(1978));
    layer3_outputs(1883) <= (layer2_outputs(2248)) or (layer2_outputs(4019));
    layer3_outputs(1884) <= (layer2_outputs(2397)) and not (layer2_outputs(3182));
    layer3_outputs(1885) <= not((layer2_outputs(5063)) and (layer2_outputs(5076)));
    layer3_outputs(1886) <= layer2_outputs(650);
    layer3_outputs(1887) <= '1';
    layer3_outputs(1888) <= (layer2_outputs(1889)) or (layer2_outputs(4842));
    layer3_outputs(1889) <= not(layer2_outputs(3631));
    layer3_outputs(1890) <= layer2_outputs(1709);
    layer3_outputs(1891) <= '0';
    layer3_outputs(1892) <= layer2_outputs(3228);
    layer3_outputs(1893) <= (layer2_outputs(4632)) and not (layer2_outputs(122));
    layer3_outputs(1894) <= not((layer2_outputs(3520)) or (layer2_outputs(454)));
    layer3_outputs(1895) <= (layer2_outputs(4762)) and not (layer2_outputs(3106));
    layer3_outputs(1896) <= (layer2_outputs(1947)) and (layer2_outputs(3090));
    layer3_outputs(1897) <= layer2_outputs(3145);
    layer3_outputs(1898) <= (layer2_outputs(251)) and not (layer2_outputs(3546));
    layer3_outputs(1899) <= (layer2_outputs(4263)) and (layer2_outputs(890));
    layer3_outputs(1900) <= not((layer2_outputs(993)) and (layer2_outputs(202)));
    layer3_outputs(1901) <= (layer2_outputs(369)) or (layer2_outputs(2547));
    layer3_outputs(1902) <= not(layer2_outputs(1534));
    layer3_outputs(1903) <= (layer2_outputs(1761)) and not (layer2_outputs(2942));
    layer3_outputs(1904) <= '1';
    layer3_outputs(1905) <= layer2_outputs(3679);
    layer3_outputs(1906) <= layer2_outputs(626);
    layer3_outputs(1907) <= layer2_outputs(3661);
    layer3_outputs(1908) <= '1';
    layer3_outputs(1909) <= not((layer2_outputs(1609)) or (layer2_outputs(2668)));
    layer3_outputs(1910) <= '0';
    layer3_outputs(1911) <= (layer2_outputs(785)) and not (layer2_outputs(2969));
    layer3_outputs(1912) <= (layer2_outputs(1624)) and not (layer2_outputs(2480));
    layer3_outputs(1913) <= not(layer2_outputs(4163));
    layer3_outputs(1914) <= not(layer2_outputs(4232));
    layer3_outputs(1915) <= (layer2_outputs(3699)) or (layer2_outputs(2182));
    layer3_outputs(1916) <= not((layer2_outputs(1878)) and (layer2_outputs(4765)));
    layer3_outputs(1917) <= (layer2_outputs(2951)) or (layer2_outputs(2055));
    layer3_outputs(1918) <= (layer2_outputs(4365)) and not (layer2_outputs(232));
    layer3_outputs(1919) <= not(layer2_outputs(2557));
    layer3_outputs(1920) <= '1';
    layer3_outputs(1921) <= not((layer2_outputs(1329)) and (layer2_outputs(2305)));
    layer3_outputs(1922) <= (layer2_outputs(3728)) and not (layer2_outputs(3977));
    layer3_outputs(1923) <= '0';
    layer3_outputs(1924) <= not(layer2_outputs(4477));
    layer3_outputs(1925) <= not(layer2_outputs(4488)) or (layer2_outputs(664));
    layer3_outputs(1926) <= '0';
    layer3_outputs(1927) <= (layer2_outputs(3234)) and not (layer2_outputs(4195));
    layer3_outputs(1928) <= not(layer2_outputs(1257));
    layer3_outputs(1929) <= '0';
    layer3_outputs(1930) <= '1';
    layer3_outputs(1931) <= (layer2_outputs(2028)) or (layer2_outputs(1860));
    layer3_outputs(1932) <= not((layer2_outputs(4479)) and (layer2_outputs(4324)));
    layer3_outputs(1933) <= '0';
    layer3_outputs(1934) <= '0';
    layer3_outputs(1935) <= '1';
    layer3_outputs(1936) <= not(layer2_outputs(4917));
    layer3_outputs(1937) <= '1';
    layer3_outputs(1938) <= '1';
    layer3_outputs(1939) <= not((layer2_outputs(4425)) xor (layer2_outputs(4033)));
    layer3_outputs(1940) <= (layer2_outputs(3682)) and not (layer2_outputs(4009));
    layer3_outputs(1941) <= layer2_outputs(192);
    layer3_outputs(1942) <= not((layer2_outputs(277)) or (layer2_outputs(4220)));
    layer3_outputs(1943) <= not(layer2_outputs(1036));
    layer3_outputs(1944) <= '1';
    layer3_outputs(1945) <= '0';
    layer3_outputs(1946) <= (layer2_outputs(519)) or (layer2_outputs(3470));
    layer3_outputs(1947) <= (layer2_outputs(4964)) and not (layer2_outputs(208));
    layer3_outputs(1948) <= not(layer2_outputs(4161)) or (layer2_outputs(4261));
    layer3_outputs(1949) <= not((layer2_outputs(659)) or (layer2_outputs(4869)));
    layer3_outputs(1950) <= '1';
    layer3_outputs(1951) <= '0';
    layer3_outputs(1952) <= not((layer2_outputs(2375)) or (layer2_outputs(4446)));
    layer3_outputs(1953) <= '0';
    layer3_outputs(1954) <= (layer2_outputs(3861)) and not (layer2_outputs(2784));
    layer3_outputs(1955) <= '0';
    layer3_outputs(1956) <= (layer2_outputs(2387)) and (layer2_outputs(3777));
    layer3_outputs(1957) <= layer2_outputs(3048);
    layer3_outputs(1958) <= (layer2_outputs(3738)) and not (layer2_outputs(5019));
    layer3_outputs(1959) <= (layer2_outputs(1931)) or (layer2_outputs(385));
    layer3_outputs(1960) <= layer2_outputs(4539);
    layer3_outputs(1961) <= not((layer2_outputs(4031)) and (layer2_outputs(4430)));
    layer3_outputs(1962) <= (layer2_outputs(801)) or (layer2_outputs(5061));
    layer3_outputs(1963) <= not(layer2_outputs(2671));
    layer3_outputs(1964) <= not(layer2_outputs(4010));
    layer3_outputs(1965) <= layer2_outputs(3107);
    layer3_outputs(1966) <= not(layer2_outputs(3771)) or (layer2_outputs(3527));
    layer3_outputs(1967) <= (layer2_outputs(2144)) and not (layer2_outputs(3649));
    layer3_outputs(1968) <= '1';
    layer3_outputs(1969) <= (layer2_outputs(2323)) or (layer2_outputs(2234));
    layer3_outputs(1970) <= not(layer2_outputs(3048)) or (layer2_outputs(4082));
    layer3_outputs(1971) <= '1';
    layer3_outputs(1972) <= (layer2_outputs(1392)) and (layer2_outputs(4099));
    layer3_outputs(1973) <= layer2_outputs(4256);
    layer3_outputs(1974) <= (layer2_outputs(578)) and (layer2_outputs(2530));
    layer3_outputs(1975) <= not(layer2_outputs(3729)) or (layer2_outputs(4670));
    layer3_outputs(1976) <= (layer2_outputs(4648)) xor (layer2_outputs(3751));
    layer3_outputs(1977) <= not((layer2_outputs(5081)) and (layer2_outputs(2742)));
    layer3_outputs(1978) <= not(layer2_outputs(2849));
    layer3_outputs(1979) <= not(layer2_outputs(3000));
    layer3_outputs(1980) <= '0';
    layer3_outputs(1981) <= '0';
    layer3_outputs(1982) <= (layer2_outputs(2043)) or (layer2_outputs(3837));
    layer3_outputs(1983) <= layer2_outputs(2116);
    layer3_outputs(1984) <= (layer2_outputs(772)) and (layer2_outputs(2179));
    layer3_outputs(1985) <= not((layer2_outputs(75)) or (layer2_outputs(2835)));
    layer3_outputs(1986) <= not((layer2_outputs(1291)) xor (layer2_outputs(2683)));
    layer3_outputs(1987) <= layer2_outputs(2665);
    layer3_outputs(1988) <= layer2_outputs(3358);
    layer3_outputs(1989) <= not(layer2_outputs(783)) or (layer2_outputs(4804));
    layer3_outputs(1990) <= not(layer2_outputs(3243));
    layer3_outputs(1991) <= layer2_outputs(1058);
    layer3_outputs(1992) <= (layer2_outputs(3867)) and (layer2_outputs(2696));
    layer3_outputs(1993) <= '0';
    layer3_outputs(1994) <= not((layer2_outputs(2084)) or (layer2_outputs(190)));
    layer3_outputs(1995) <= not((layer2_outputs(3849)) or (layer2_outputs(1912)));
    layer3_outputs(1996) <= not(layer2_outputs(3813));
    layer3_outputs(1997) <= not((layer2_outputs(982)) and (layer2_outputs(4277)));
    layer3_outputs(1998) <= not((layer2_outputs(97)) and (layer2_outputs(4017)));
    layer3_outputs(1999) <= (layer2_outputs(5013)) or (layer2_outputs(4650));
    layer3_outputs(2000) <= (layer2_outputs(2676)) or (layer2_outputs(4124));
    layer3_outputs(2001) <= layer2_outputs(1535);
    layer3_outputs(2002) <= not((layer2_outputs(4758)) or (layer2_outputs(1950)));
    layer3_outputs(2003) <= (layer2_outputs(2473)) or (layer2_outputs(2785));
    layer3_outputs(2004) <= '0';
    layer3_outputs(2005) <= not(layer2_outputs(5094));
    layer3_outputs(2006) <= not(layer2_outputs(3654));
    layer3_outputs(2007) <= '0';
    layer3_outputs(2008) <= (layer2_outputs(2247)) and not (layer2_outputs(4599));
    layer3_outputs(2009) <= '1';
    layer3_outputs(2010) <= (layer2_outputs(3985)) and not (layer2_outputs(4584));
    layer3_outputs(2011) <= '1';
    layer3_outputs(2012) <= not((layer2_outputs(3815)) or (layer2_outputs(923)));
    layer3_outputs(2013) <= (layer2_outputs(2357)) or (layer2_outputs(248));
    layer3_outputs(2014) <= not(layer2_outputs(1083));
    layer3_outputs(2015) <= not(layer2_outputs(4421));
    layer3_outputs(2016) <= not(layer2_outputs(3278));
    layer3_outputs(2017) <= not(layer2_outputs(300));
    layer3_outputs(2018) <= layer2_outputs(2289);
    layer3_outputs(2019) <= not((layer2_outputs(3187)) and (layer2_outputs(1137)));
    layer3_outputs(2020) <= '0';
    layer3_outputs(2021) <= '1';
    layer3_outputs(2022) <= layer2_outputs(4680);
    layer3_outputs(2023) <= not(layer2_outputs(3409));
    layer3_outputs(2024) <= not(layer2_outputs(12)) or (layer2_outputs(70));
    layer3_outputs(2025) <= (layer2_outputs(661)) and (layer2_outputs(1682));
    layer3_outputs(2026) <= layer2_outputs(911);
    layer3_outputs(2027) <= not(layer2_outputs(3635));
    layer3_outputs(2028) <= not((layer2_outputs(2891)) and (layer2_outputs(4800)));
    layer3_outputs(2029) <= (layer2_outputs(1699)) or (layer2_outputs(2210));
    layer3_outputs(2030) <= (layer2_outputs(2175)) and not (layer2_outputs(3562));
    layer3_outputs(2031) <= layer2_outputs(345);
    layer3_outputs(2032) <= not((layer2_outputs(2391)) and (layer2_outputs(468)));
    layer3_outputs(2033) <= not((layer2_outputs(3146)) or (layer2_outputs(1735)));
    layer3_outputs(2034) <= (layer2_outputs(4936)) and not (layer2_outputs(4704));
    layer3_outputs(2035) <= (layer2_outputs(402)) and not (layer2_outputs(2150));
    layer3_outputs(2036) <= '0';
    layer3_outputs(2037) <= not(layer2_outputs(4193));
    layer3_outputs(2038) <= not((layer2_outputs(1350)) and (layer2_outputs(470)));
    layer3_outputs(2039) <= '0';
    layer3_outputs(2040) <= '0';
    layer3_outputs(2041) <= not(layer2_outputs(1761));
    layer3_outputs(2042) <= '1';
    layer3_outputs(2043) <= '0';
    layer3_outputs(2044) <= layer2_outputs(1359);
    layer3_outputs(2045) <= '1';
    layer3_outputs(2046) <= '1';
    layer3_outputs(2047) <= not(layer2_outputs(4149)) or (layer2_outputs(3184));
    layer3_outputs(2048) <= '1';
    layer3_outputs(2049) <= not(layer2_outputs(1103));
    layer3_outputs(2050) <= (layer2_outputs(1124)) and not (layer2_outputs(1452));
    layer3_outputs(2051) <= '0';
    layer3_outputs(2052) <= not(layer2_outputs(1683)) or (layer2_outputs(2759));
    layer3_outputs(2053) <= not(layer2_outputs(1567)) or (layer2_outputs(1826));
    layer3_outputs(2054) <= not((layer2_outputs(2197)) and (layer2_outputs(931)));
    layer3_outputs(2055) <= (layer2_outputs(1957)) or (layer2_outputs(2216));
    layer3_outputs(2056) <= not(layer2_outputs(1751));
    layer3_outputs(2057) <= (layer2_outputs(2022)) and (layer2_outputs(1513));
    layer3_outputs(2058) <= (layer2_outputs(5010)) and not (layer2_outputs(3979));
    layer3_outputs(2059) <= not(layer2_outputs(649)) or (layer2_outputs(4383));
    layer3_outputs(2060) <= not((layer2_outputs(3696)) or (layer2_outputs(2049)));
    layer3_outputs(2061) <= layer2_outputs(2409);
    layer3_outputs(2062) <= not(layer2_outputs(3214));
    layer3_outputs(2063) <= not((layer2_outputs(4960)) or (layer2_outputs(4614)));
    layer3_outputs(2064) <= (layer2_outputs(1956)) xor (layer2_outputs(433));
    layer3_outputs(2065) <= (layer2_outputs(2419)) or (layer2_outputs(1284));
    layer3_outputs(2066) <= layer2_outputs(3172);
    layer3_outputs(2067) <= (layer2_outputs(4809)) xor (layer2_outputs(2050));
    layer3_outputs(2068) <= layer2_outputs(3843);
    layer3_outputs(2069) <= '0';
    layer3_outputs(2070) <= (layer2_outputs(4593)) and not (layer2_outputs(2373));
    layer3_outputs(2071) <= (layer2_outputs(3938)) or (layer2_outputs(411));
    layer3_outputs(2072) <= layer2_outputs(3472);
    layer3_outputs(2073) <= not(layer2_outputs(2260)) or (layer2_outputs(158));
    layer3_outputs(2074) <= not(layer2_outputs(373)) or (layer2_outputs(3710));
    layer3_outputs(2075) <= layer2_outputs(4276);
    layer3_outputs(2076) <= not(layer2_outputs(4988));
    layer3_outputs(2077) <= (layer2_outputs(2698)) or (layer2_outputs(539));
    layer3_outputs(2078) <= not((layer2_outputs(20)) and (layer2_outputs(1872)));
    layer3_outputs(2079) <= not((layer2_outputs(4612)) xor (layer2_outputs(3552)));
    layer3_outputs(2080) <= (layer2_outputs(1972)) and not (layer2_outputs(184));
    layer3_outputs(2081) <= '1';
    layer3_outputs(2082) <= (layer2_outputs(294)) and not (layer2_outputs(3686));
    layer3_outputs(2083) <= (layer2_outputs(1032)) or (layer2_outputs(1435));
    layer3_outputs(2084) <= layer2_outputs(4111);
    layer3_outputs(2085) <= (layer2_outputs(131)) or (layer2_outputs(4287));
    layer3_outputs(2086) <= layer2_outputs(210);
    layer3_outputs(2087) <= (layer2_outputs(585)) and (layer2_outputs(944));
    layer3_outputs(2088) <= not((layer2_outputs(2872)) and (layer2_outputs(2272)));
    layer3_outputs(2089) <= not(layer2_outputs(795));
    layer3_outputs(2090) <= (layer2_outputs(11)) and not (layer2_outputs(4174));
    layer3_outputs(2091) <= '1';
    layer3_outputs(2092) <= not((layer2_outputs(3940)) or (layer2_outputs(2232)));
    layer3_outputs(2093) <= '1';
    layer3_outputs(2094) <= (layer2_outputs(686)) or (layer2_outputs(1679));
    layer3_outputs(2095) <= '0';
    layer3_outputs(2096) <= '0';
    layer3_outputs(2097) <= not(layer2_outputs(746)) or (layer2_outputs(4016));
    layer3_outputs(2098) <= not((layer2_outputs(1405)) or (layer2_outputs(1362)));
    layer3_outputs(2099) <= '1';
    layer3_outputs(2100) <= '0';
    layer3_outputs(2101) <= '1';
    layer3_outputs(2102) <= (layer2_outputs(3510)) and (layer2_outputs(3292));
    layer3_outputs(2103) <= '1';
    layer3_outputs(2104) <= layer2_outputs(4611);
    layer3_outputs(2105) <= not(layer2_outputs(592)) or (layer2_outputs(2814));
    layer3_outputs(2106) <= '0';
    layer3_outputs(2107) <= '1';
    layer3_outputs(2108) <= not((layer2_outputs(2583)) or (layer2_outputs(262)));
    layer3_outputs(2109) <= not(layer2_outputs(1453));
    layer3_outputs(2110) <= not((layer2_outputs(4607)) and (layer2_outputs(2175)));
    layer3_outputs(2111) <= layer2_outputs(288);
    layer3_outputs(2112) <= '1';
    layer3_outputs(2113) <= layer2_outputs(3846);
    layer3_outputs(2114) <= '1';
    layer3_outputs(2115) <= not((layer2_outputs(3183)) xor (layer2_outputs(2607)));
    layer3_outputs(2116) <= (layer2_outputs(1704)) and not (layer2_outputs(1715));
    layer3_outputs(2117) <= not(layer2_outputs(4346)) or (layer2_outputs(3498));
    layer3_outputs(2118) <= (layer2_outputs(3857)) and not (layer2_outputs(3666));
    layer3_outputs(2119) <= not(layer2_outputs(1577)) or (layer2_outputs(194));
    layer3_outputs(2120) <= (layer2_outputs(2165)) and (layer2_outputs(1399));
    layer3_outputs(2121) <= not((layer2_outputs(1213)) or (layer2_outputs(3968)));
    layer3_outputs(2122) <= not(layer2_outputs(2911));
    layer3_outputs(2123) <= layer2_outputs(1361);
    layer3_outputs(2124) <= layer2_outputs(1414);
    layer3_outputs(2125) <= not(layer2_outputs(121)) or (layer2_outputs(751));
    layer3_outputs(2126) <= '0';
    layer3_outputs(2127) <= layer2_outputs(2923);
    layer3_outputs(2128) <= not(layer2_outputs(2791)) or (layer2_outputs(137));
    layer3_outputs(2129) <= not((layer2_outputs(2041)) and (layer2_outputs(4569)));
    layer3_outputs(2130) <= '0';
    layer3_outputs(2131) <= '1';
    layer3_outputs(2132) <= layer2_outputs(2526);
    layer3_outputs(2133) <= (layer2_outputs(4975)) or (layer2_outputs(4302));
    layer3_outputs(2134) <= (layer2_outputs(1975)) and (layer2_outputs(361));
    layer3_outputs(2135) <= (layer2_outputs(3998)) and not (layer2_outputs(4481));
    layer3_outputs(2136) <= not(layer2_outputs(2266));
    layer3_outputs(2137) <= not(layer2_outputs(4285)) or (layer2_outputs(721));
    layer3_outputs(2138) <= layer2_outputs(4830);
    layer3_outputs(2139) <= '0';
    layer3_outputs(2140) <= not(layer2_outputs(663));
    layer3_outputs(2141) <= '1';
    layer3_outputs(2142) <= not((layer2_outputs(4837)) and (layer2_outputs(4116)));
    layer3_outputs(2143) <= not((layer2_outputs(494)) and (layer2_outputs(4042)));
    layer3_outputs(2144) <= '0';
    layer3_outputs(2145) <= not(layer2_outputs(5055)) or (layer2_outputs(3452));
    layer3_outputs(2146) <= '1';
    layer3_outputs(2147) <= not((layer2_outputs(991)) and (layer2_outputs(2488)));
    layer3_outputs(2148) <= (layer2_outputs(3955)) or (layer2_outputs(2396));
    layer3_outputs(2149) <= not(layer2_outputs(2481)) or (layer2_outputs(1531));
    layer3_outputs(2150) <= (layer2_outputs(5056)) and not (layer2_outputs(1383));
    layer3_outputs(2151) <= not(layer2_outputs(2916)) or (layer2_outputs(4962));
    layer3_outputs(2152) <= (layer2_outputs(2745)) and not (layer2_outputs(4469));
    layer3_outputs(2153) <= not(layer2_outputs(4810)) or (layer2_outputs(64));
    layer3_outputs(2154) <= not(layer2_outputs(4470));
    layer3_outputs(2155) <= not(layer2_outputs(3003));
    layer3_outputs(2156) <= not((layer2_outputs(1965)) xor (layer2_outputs(1786)));
    layer3_outputs(2157) <= (layer2_outputs(177)) and not (layer2_outputs(3829));
    layer3_outputs(2158) <= not(layer2_outputs(514)) or (layer2_outputs(2351));
    layer3_outputs(2159) <= not((layer2_outputs(3070)) and (layer2_outputs(4882)));
    layer3_outputs(2160) <= not(layer2_outputs(4100)) or (layer2_outputs(258));
    layer3_outputs(2161) <= '0';
    layer3_outputs(2162) <= (layer2_outputs(552)) and (layer2_outputs(3201));
    layer3_outputs(2163) <= not(layer2_outputs(3597));
    layer3_outputs(2164) <= '0';
    layer3_outputs(2165) <= not(layer2_outputs(1057));
    layer3_outputs(2166) <= (layer2_outputs(4871)) and not (layer2_outputs(40));
    layer3_outputs(2167) <= '0';
    layer3_outputs(2168) <= not((layer2_outputs(731)) and (layer2_outputs(3458)));
    layer3_outputs(2169) <= (layer2_outputs(2869)) or (layer2_outputs(5010));
    layer3_outputs(2170) <= (layer2_outputs(4833)) or (layer2_outputs(4897));
    layer3_outputs(2171) <= '0';
    layer3_outputs(2172) <= layer2_outputs(2282);
    layer3_outputs(2173) <= (layer2_outputs(2535)) and not (layer2_outputs(3641));
    layer3_outputs(2174) <= layer2_outputs(3723);
    layer3_outputs(2175) <= (layer2_outputs(621)) and not (layer2_outputs(3244));
    layer3_outputs(2176) <= layer2_outputs(392);
    layer3_outputs(2177) <= not((layer2_outputs(2778)) or (layer2_outputs(1794)));
    layer3_outputs(2178) <= (layer2_outputs(5087)) and not (layer2_outputs(1846));
    layer3_outputs(2179) <= '0';
    layer3_outputs(2180) <= layer2_outputs(335);
    layer3_outputs(2181) <= not(layer2_outputs(5033));
    layer3_outputs(2182) <= not(layer2_outputs(1901)) or (layer2_outputs(2889));
    layer3_outputs(2183) <= not(layer2_outputs(2756));
    layer3_outputs(2184) <= not(layer2_outputs(166)) or (layer2_outputs(4004));
    layer3_outputs(2185) <= '1';
    layer3_outputs(2186) <= not(layer2_outputs(978));
    layer3_outputs(2187) <= not(layer2_outputs(1701));
    layer3_outputs(2188) <= not(layer2_outputs(4489)) or (layer2_outputs(1789));
    layer3_outputs(2189) <= (layer2_outputs(80)) or (layer2_outputs(652));
    layer3_outputs(2190) <= (layer2_outputs(1804)) and not (layer2_outputs(4442));
    layer3_outputs(2191) <= (layer2_outputs(3283)) and not (layer2_outputs(2760));
    layer3_outputs(2192) <= layer2_outputs(4162);
    layer3_outputs(2193) <= not((layer2_outputs(788)) or (layer2_outputs(2446)));
    layer3_outputs(2194) <= (layer2_outputs(809)) and (layer2_outputs(1222));
    layer3_outputs(2195) <= (layer2_outputs(2864)) and not (layer2_outputs(4034));
    layer3_outputs(2196) <= not((layer2_outputs(2431)) or (layer2_outputs(935)));
    layer3_outputs(2197) <= not((layer2_outputs(109)) and (layer2_outputs(402)));
    layer3_outputs(2198) <= layer2_outputs(1155);
    layer3_outputs(2199) <= not(layer2_outputs(4801)) or (layer2_outputs(303));
    layer3_outputs(2200) <= not(layer2_outputs(3897));
    layer3_outputs(2201) <= not((layer2_outputs(625)) or (layer2_outputs(1602)));
    layer3_outputs(2202) <= not((layer2_outputs(84)) and (layer2_outputs(4796)));
    layer3_outputs(2203) <= (layer2_outputs(2009)) xor (layer2_outputs(3199));
    layer3_outputs(2204) <= '1';
    layer3_outputs(2205) <= not(layer2_outputs(5107)) or (layer2_outputs(1556));
    layer3_outputs(2206) <= not(layer2_outputs(3843)) or (layer2_outputs(4157));
    layer3_outputs(2207) <= (layer2_outputs(5007)) and not (layer2_outputs(792));
    layer3_outputs(2208) <= not((layer2_outputs(2239)) and (layer2_outputs(3601)));
    layer3_outputs(2209) <= (layer2_outputs(1314)) and (layer2_outputs(4101));
    layer3_outputs(2210) <= '1';
    layer3_outputs(2211) <= not(layer2_outputs(3349)) or (layer2_outputs(3344));
    layer3_outputs(2212) <= (layer2_outputs(3385)) or (layer2_outputs(2010));
    layer3_outputs(2213) <= not((layer2_outputs(2183)) and (layer2_outputs(3221)));
    layer3_outputs(2214) <= (layer2_outputs(741)) and not (layer2_outputs(4268));
    layer3_outputs(2215) <= '0';
    layer3_outputs(2216) <= not((layer2_outputs(1971)) or (layer2_outputs(2451)));
    layer3_outputs(2217) <= (layer2_outputs(2050)) and not (layer2_outputs(775));
    layer3_outputs(2218) <= '1';
    layer3_outputs(2219) <= (layer2_outputs(3891)) and (layer2_outputs(2017));
    layer3_outputs(2220) <= (layer2_outputs(1853)) and not (layer2_outputs(1060));
    layer3_outputs(2221) <= (layer2_outputs(2246)) xor (layer2_outputs(319));
    layer3_outputs(2222) <= not((layer2_outputs(1960)) and (layer2_outputs(104)));
    layer3_outputs(2223) <= not(layer2_outputs(867));
    layer3_outputs(2224) <= not(layer2_outputs(1593)) or (layer2_outputs(767));
    layer3_outputs(2225) <= '1';
    layer3_outputs(2226) <= not(layer2_outputs(3239)) or (layer2_outputs(5062));
    layer3_outputs(2227) <= (layer2_outputs(1439)) and not (layer2_outputs(4144));
    layer3_outputs(2228) <= '1';
    layer3_outputs(2229) <= (layer2_outputs(315)) and not (layer2_outputs(4980));
    layer3_outputs(2230) <= not(layer2_outputs(2151));
    layer3_outputs(2231) <= not(layer2_outputs(108)) or (layer2_outputs(2294));
    layer3_outputs(2232) <= not((layer2_outputs(2184)) and (layer2_outputs(1915)));
    layer3_outputs(2233) <= (layer2_outputs(1639)) and (layer2_outputs(975));
    layer3_outputs(2234) <= not((layer2_outputs(571)) and (layer2_outputs(964)));
    layer3_outputs(2235) <= (layer2_outputs(4818)) and not (layer2_outputs(1098));
    layer3_outputs(2236) <= (layer2_outputs(4132)) xor (layer2_outputs(605));
    layer3_outputs(2237) <= not(layer2_outputs(4005)) or (layer2_outputs(1703));
    layer3_outputs(2238) <= not(layer2_outputs(1784));
    layer3_outputs(2239) <= (layer2_outputs(4225)) and not (layer2_outputs(3664));
    layer3_outputs(2240) <= not((layer2_outputs(33)) and (layer2_outputs(2626)));
    layer3_outputs(2241) <= layer2_outputs(480);
    layer3_outputs(2242) <= (layer2_outputs(256)) and not (layer2_outputs(625));
    layer3_outputs(2243) <= not(layer2_outputs(4771)) or (layer2_outputs(2835));
    layer3_outputs(2244) <= not(layer2_outputs(3752)) or (layer2_outputs(2454));
    layer3_outputs(2245) <= layer2_outputs(657);
    layer3_outputs(2246) <= not(layer2_outputs(2825));
    layer3_outputs(2247) <= not(layer2_outputs(19)) or (layer2_outputs(401));
    layer3_outputs(2248) <= not(layer2_outputs(2824)) or (layer2_outputs(3076));
    layer3_outputs(2249) <= (layer2_outputs(3948)) and not (layer2_outputs(4600));
    layer3_outputs(2250) <= not(layer2_outputs(1245));
    layer3_outputs(2251) <= not(layer2_outputs(3929)) or (layer2_outputs(4654));
    layer3_outputs(2252) <= not(layer2_outputs(1175)) or (layer2_outputs(943));
    layer3_outputs(2253) <= (layer2_outputs(4051)) and (layer2_outputs(2263));
    layer3_outputs(2254) <= layer2_outputs(3676);
    layer3_outputs(2255) <= (layer2_outputs(3329)) and not (layer2_outputs(3444));
    layer3_outputs(2256) <= (layer2_outputs(2316)) and not (layer2_outputs(5036));
    layer3_outputs(2257) <= not(layer2_outputs(3683));
    layer3_outputs(2258) <= '1';
    layer3_outputs(2259) <= '0';
    layer3_outputs(2260) <= '1';
    layer3_outputs(2261) <= (layer2_outputs(5095)) and (layer2_outputs(375));
    layer3_outputs(2262) <= not((layer2_outputs(2002)) and (layer2_outputs(2513)));
    layer3_outputs(2263) <= (layer2_outputs(3980)) and (layer2_outputs(2554));
    layer3_outputs(2264) <= not(layer2_outputs(1820)) or (layer2_outputs(5046));
    layer3_outputs(2265) <= (layer2_outputs(4)) or (layer2_outputs(4598));
    layer3_outputs(2266) <= not(layer2_outputs(4691)) or (layer2_outputs(2596));
    layer3_outputs(2267) <= not(layer2_outputs(2955)) or (layer2_outputs(3881));
    layer3_outputs(2268) <= not(layer2_outputs(215)) or (layer2_outputs(1441));
    layer3_outputs(2269) <= layer2_outputs(4256);
    layer3_outputs(2270) <= not((layer2_outputs(608)) or (layer2_outputs(3830)));
    layer3_outputs(2271) <= layer2_outputs(3748);
    layer3_outputs(2272) <= (layer2_outputs(4672)) and not (layer2_outputs(1927));
    layer3_outputs(2273) <= '1';
    layer3_outputs(2274) <= '0';
    layer3_outputs(2275) <= not((layer2_outputs(4348)) or (layer2_outputs(937)));
    layer3_outputs(2276) <= not(layer2_outputs(3927));
    layer3_outputs(2277) <= (layer2_outputs(2196)) and (layer2_outputs(4077));
    layer3_outputs(2278) <= not((layer2_outputs(171)) or (layer2_outputs(4749)));
    layer3_outputs(2279) <= (layer2_outputs(66)) and not (layer2_outputs(4218));
    layer3_outputs(2280) <= not(layer2_outputs(2325)) or (layer2_outputs(1771));
    layer3_outputs(2281) <= not(layer2_outputs(4494));
    layer3_outputs(2282) <= '1';
    layer3_outputs(2283) <= layer2_outputs(4528);
    layer3_outputs(2284) <= (layer2_outputs(530)) and not (layer2_outputs(776));
    layer3_outputs(2285) <= '1';
    layer3_outputs(2286) <= (layer2_outputs(4034)) and not (layer2_outputs(763));
    layer3_outputs(2287) <= (layer2_outputs(4695)) or (layer2_outputs(3670));
    layer3_outputs(2288) <= '1';
    layer3_outputs(2289) <= '1';
    layer3_outputs(2290) <= not((layer2_outputs(4155)) and (layer2_outputs(4770)));
    layer3_outputs(2291) <= (layer2_outputs(5097)) and (layer2_outputs(604));
    layer3_outputs(2292) <= not(layer2_outputs(2718));
    layer3_outputs(2293) <= not((layer2_outputs(2760)) and (layer2_outputs(2602)));
    layer3_outputs(2294) <= '0';
    layer3_outputs(2295) <= not(layer2_outputs(4822));
    layer3_outputs(2296) <= not((layer2_outputs(310)) and (layer2_outputs(2677)));
    layer3_outputs(2297) <= not(layer2_outputs(909));
    layer3_outputs(2298) <= not(layer2_outputs(4512)) or (layer2_outputs(848));
    layer3_outputs(2299) <= layer2_outputs(3363);
    layer3_outputs(2300) <= layer2_outputs(4155);
    layer3_outputs(2301) <= not((layer2_outputs(1714)) or (layer2_outputs(1332)));
    layer3_outputs(2302) <= not((layer2_outputs(3127)) or (layer2_outputs(3574)));
    layer3_outputs(2303) <= layer2_outputs(3995);
    layer3_outputs(2304) <= (layer2_outputs(120)) and not (layer2_outputs(4899));
    layer3_outputs(2305) <= not(layer2_outputs(1396));
    layer3_outputs(2306) <= layer2_outputs(3675);
    layer3_outputs(2307) <= not(layer2_outputs(1687)) or (layer2_outputs(405));
    layer3_outputs(2308) <= (layer2_outputs(2676)) and not (layer2_outputs(4490));
    layer3_outputs(2309) <= (layer2_outputs(2905)) and not (layer2_outputs(4739));
    layer3_outputs(2310) <= (layer2_outputs(264)) and not (layer2_outputs(2998));
    layer3_outputs(2311) <= '1';
    layer3_outputs(2312) <= not(layer2_outputs(308));
    layer3_outputs(2313) <= layer2_outputs(2818);
    layer3_outputs(2314) <= layer2_outputs(3458);
    layer3_outputs(2315) <= not(layer2_outputs(908)) or (layer2_outputs(4515));
    layer3_outputs(2316) <= (layer2_outputs(340)) and (layer2_outputs(1314));
    layer3_outputs(2317) <= not(layer2_outputs(3020)) or (layer2_outputs(3874));
    layer3_outputs(2318) <= not((layer2_outputs(2954)) and (layer2_outputs(2963)));
    layer3_outputs(2319) <= '0';
    layer3_outputs(2320) <= not((layer2_outputs(971)) and (layer2_outputs(2403)));
    layer3_outputs(2321) <= not(layer2_outputs(988)) or (layer2_outputs(3819));
    layer3_outputs(2322) <= (layer2_outputs(4824)) and (layer2_outputs(67));
    layer3_outputs(2323) <= not(layer2_outputs(461)) or (layer2_outputs(1056));
    layer3_outputs(2324) <= layer2_outputs(3256);
    layer3_outputs(2325) <= (layer2_outputs(1014)) and not (layer2_outputs(1710));
    layer3_outputs(2326) <= (layer2_outputs(4257)) or (layer2_outputs(547));
    layer3_outputs(2327) <= layer2_outputs(438);
    layer3_outputs(2328) <= not(layer2_outputs(3675));
    layer3_outputs(2329) <= '1';
    layer3_outputs(2330) <= not((layer2_outputs(4490)) or (layer2_outputs(493)));
    layer3_outputs(2331) <= not((layer2_outputs(3078)) or (layer2_outputs(1948)));
    layer3_outputs(2332) <= '1';
    layer3_outputs(2333) <= not((layer2_outputs(27)) or (layer2_outputs(395)));
    layer3_outputs(2334) <= (layer2_outputs(3620)) and (layer2_outputs(8));
    layer3_outputs(2335) <= layer2_outputs(42);
    layer3_outputs(2336) <= not((layer2_outputs(3937)) or (layer2_outputs(750)));
    layer3_outputs(2337) <= '1';
    layer3_outputs(2338) <= '0';
    layer3_outputs(2339) <= (layer2_outputs(4159)) or (layer2_outputs(757));
    layer3_outputs(2340) <= not((layer2_outputs(3829)) and (layer2_outputs(963)));
    layer3_outputs(2341) <= not(layer2_outputs(2990)) or (layer2_outputs(3750));
    layer3_outputs(2342) <= '0';
    layer3_outputs(2343) <= (layer2_outputs(4216)) and not (layer2_outputs(48));
    layer3_outputs(2344) <= (layer2_outputs(1110)) and not (layer2_outputs(1013));
    layer3_outputs(2345) <= (layer2_outputs(276)) xor (layer2_outputs(2932));
    layer3_outputs(2346) <= '1';
    layer3_outputs(2347) <= not(layer2_outputs(1753)) or (layer2_outputs(3895));
    layer3_outputs(2348) <= not((layer2_outputs(2691)) or (layer2_outputs(1785)));
    layer3_outputs(2349) <= not((layer2_outputs(3982)) or (layer2_outputs(3111)));
    layer3_outputs(2350) <= not((layer2_outputs(1038)) or (layer2_outputs(581)));
    layer3_outputs(2351) <= not((layer2_outputs(3561)) or (layer2_outputs(1563)));
    layer3_outputs(2352) <= '0';
    layer3_outputs(2353) <= (layer2_outputs(3150)) and (layer2_outputs(1768));
    layer3_outputs(2354) <= '1';
    layer3_outputs(2355) <= '0';
    layer3_outputs(2356) <= not((layer2_outputs(4569)) and (layer2_outputs(1423)));
    layer3_outputs(2357) <= not((layer2_outputs(2417)) and (layer2_outputs(3927)));
    layer3_outputs(2358) <= layer2_outputs(4901);
    layer3_outputs(2359) <= not(layer2_outputs(4517)) or (layer2_outputs(2541));
    layer3_outputs(2360) <= not((layer2_outputs(4916)) and (layer2_outputs(2208)));
    layer3_outputs(2361) <= not((layer2_outputs(1783)) xor (layer2_outputs(4165)));
    layer3_outputs(2362) <= not(layer2_outputs(1458));
    layer3_outputs(2363) <= not((layer2_outputs(875)) or (layer2_outputs(3156)));
    layer3_outputs(2364) <= not((layer2_outputs(4116)) or (layer2_outputs(2049)));
    layer3_outputs(2365) <= (layer2_outputs(698)) and not (layer2_outputs(4697));
    layer3_outputs(2366) <= '0';
    layer3_outputs(2367) <= layer2_outputs(5066);
    layer3_outputs(2368) <= (layer2_outputs(2110)) and (layer2_outputs(3440));
    layer3_outputs(2369) <= not((layer2_outputs(1707)) and (layer2_outputs(2070)));
    layer3_outputs(2370) <= (layer2_outputs(4156)) and not (layer2_outputs(2730));
    layer3_outputs(2371) <= (layer2_outputs(730)) and (layer2_outputs(2268));
    layer3_outputs(2372) <= (layer2_outputs(2873)) and not (layer2_outputs(1746));
    layer3_outputs(2373) <= '1';
    layer3_outputs(2374) <= not((layer2_outputs(1551)) or (layer2_outputs(2376)));
    layer3_outputs(2375) <= layer2_outputs(952);
    layer3_outputs(2376) <= '0';
    layer3_outputs(2377) <= (layer2_outputs(2331)) and not (layer2_outputs(305));
    layer3_outputs(2378) <= '0';
    layer3_outputs(2379) <= not(layer2_outputs(713)) or (layer2_outputs(3477));
    layer3_outputs(2380) <= '1';
    layer3_outputs(2381) <= (layer2_outputs(2118)) and not (layer2_outputs(3464));
    layer3_outputs(2382) <= (layer2_outputs(908)) and not (layer2_outputs(32));
    layer3_outputs(2383) <= not(layer2_outputs(2346)) or (layer2_outputs(4955));
    layer3_outputs(2384) <= '0';
    layer3_outputs(2385) <= not(layer2_outputs(950)) or (layer2_outputs(2508));
    layer3_outputs(2386) <= not((layer2_outputs(4552)) and (layer2_outputs(754)));
    layer3_outputs(2387) <= not((layer2_outputs(327)) and (layer2_outputs(1350)));
    layer3_outputs(2388) <= not(layer2_outputs(495));
    layer3_outputs(2389) <= (layer2_outputs(1047)) and not (layer2_outputs(16));
    layer3_outputs(2390) <= (layer2_outputs(1344)) or (layer2_outputs(3664));
    layer3_outputs(2391) <= not(layer2_outputs(4191));
    layer3_outputs(2392) <= not((layer2_outputs(4782)) and (layer2_outputs(1603)));
    layer3_outputs(2393) <= (layer2_outputs(2042)) and not (layer2_outputs(419));
    layer3_outputs(2394) <= not(layer2_outputs(1896));
    layer3_outputs(2395) <= not(layer2_outputs(4792));
    layer3_outputs(2396) <= '0';
    layer3_outputs(2397) <= (layer2_outputs(2985)) and (layer2_outputs(3140));
    layer3_outputs(2398) <= not((layer2_outputs(1581)) or (layer2_outputs(1839)));
    layer3_outputs(2399) <= not((layer2_outputs(3379)) and (layer2_outputs(3715)));
    layer3_outputs(2400) <= not((layer2_outputs(2119)) and (layer2_outputs(3983)));
    layer3_outputs(2401) <= '0';
    layer3_outputs(2402) <= not((layer2_outputs(3351)) or (layer2_outputs(670)));
    layer3_outputs(2403) <= '1';
    layer3_outputs(2404) <= (layer2_outputs(4274)) and not (layer2_outputs(4107));
    layer3_outputs(2405) <= '0';
    layer3_outputs(2406) <= not((layer2_outputs(3648)) and (layer2_outputs(593)));
    layer3_outputs(2407) <= not(layer2_outputs(5017));
    layer3_outputs(2408) <= not((layer2_outputs(4720)) and (layer2_outputs(3054)));
    layer3_outputs(2409) <= not(layer2_outputs(109));
    layer3_outputs(2410) <= not((layer2_outputs(1208)) and (layer2_outputs(2892)));
    layer3_outputs(2411) <= not(layer2_outputs(1951));
    layer3_outputs(2412) <= not(layer2_outputs(1760));
    layer3_outputs(2413) <= '0';
    layer3_outputs(2414) <= not(layer2_outputs(3343)) or (layer2_outputs(1005));
    layer3_outputs(2415) <= not((layer2_outputs(1454)) and (layer2_outputs(4030)));
    layer3_outputs(2416) <= '0';
    layer3_outputs(2417) <= '0';
    layer3_outputs(2418) <= not(layer2_outputs(1739));
    layer3_outputs(2419) <= (layer2_outputs(4507)) and not (layer2_outputs(3737));
    layer3_outputs(2420) <= (layer2_outputs(226)) or (layer2_outputs(3313));
    layer3_outputs(2421) <= not(layer2_outputs(3699));
    layer3_outputs(2422) <= not(layer2_outputs(4915)) or (layer2_outputs(3294));
    layer3_outputs(2423) <= not(layer2_outputs(3680));
    layer3_outputs(2424) <= layer2_outputs(3799);
    layer3_outputs(2425) <= '0';
    layer3_outputs(2426) <= '0';
    layer3_outputs(2427) <= not((layer2_outputs(4091)) and (layer2_outputs(2285)));
    layer3_outputs(2428) <= not(layer2_outputs(5086)) or (layer2_outputs(3162));
    layer3_outputs(2429) <= (layer2_outputs(3907)) and not (layer2_outputs(2067));
    layer3_outputs(2430) <= '0';
    layer3_outputs(2431) <= not(layer2_outputs(2613));
    layer3_outputs(2432) <= '1';
    layer3_outputs(2433) <= '0';
    layer3_outputs(2434) <= '0';
    layer3_outputs(2435) <= '0';
    layer3_outputs(2436) <= '1';
    layer3_outputs(2437) <= (layer2_outputs(344)) and (layer2_outputs(789));
    layer3_outputs(2438) <= not(layer2_outputs(3330)) or (layer2_outputs(3863));
    layer3_outputs(2439) <= not(layer2_outputs(225)) or (layer2_outputs(2194));
    layer3_outputs(2440) <= (layer2_outputs(2257)) and not (layer2_outputs(3720));
    layer3_outputs(2441) <= '1';
    layer3_outputs(2442) <= '1';
    layer3_outputs(2443) <= (layer2_outputs(2261)) or (layer2_outputs(896));
    layer3_outputs(2444) <= not((layer2_outputs(2622)) and (layer2_outputs(745)));
    layer3_outputs(2445) <= (layer2_outputs(2102)) and not (layer2_outputs(183));
    layer3_outputs(2446) <= layer2_outputs(236);
    layer3_outputs(2447) <= (layer2_outputs(4517)) and (layer2_outputs(239));
    layer3_outputs(2448) <= layer2_outputs(128);
    layer3_outputs(2449) <= not((layer2_outputs(1163)) or (layer2_outputs(4952)));
    layer3_outputs(2450) <= not(layer2_outputs(3695)) or (layer2_outputs(3554));
    layer3_outputs(2451) <= '0';
    layer3_outputs(2452) <= not((layer2_outputs(2574)) or (layer2_outputs(3061)));
    layer3_outputs(2453) <= not((layer2_outputs(4404)) and (layer2_outputs(3681)));
    layer3_outputs(2454) <= (layer2_outputs(2991)) and not (layer2_outputs(5026));
    layer3_outputs(2455) <= not(layer2_outputs(4935)) or (layer2_outputs(580));
    layer3_outputs(2456) <= (layer2_outputs(173)) and (layer2_outputs(3812));
    layer3_outputs(2457) <= not(layer2_outputs(3790)) or (layer2_outputs(3802));
    layer3_outputs(2458) <= '0';
    layer3_outputs(2459) <= '1';
    layer3_outputs(2460) <= (layer2_outputs(2768)) and not (layer2_outputs(2934));
    layer3_outputs(2461) <= '0';
    layer3_outputs(2462) <= (layer2_outputs(1374)) or (layer2_outputs(1980));
    layer3_outputs(2463) <= not(layer2_outputs(2057));
    layer3_outputs(2464) <= not(layer2_outputs(1846)) or (layer2_outputs(2327));
    layer3_outputs(2465) <= '1';
    layer3_outputs(2466) <= not((layer2_outputs(3011)) or (layer2_outputs(4771)));
    layer3_outputs(2467) <= not(layer2_outputs(4458)) or (layer2_outputs(4362));
    layer3_outputs(2468) <= not(layer2_outputs(2747)) or (layer2_outputs(4781));
    layer3_outputs(2469) <= not(layer2_outputs(2810)) or (layer2_outputs(4374));
    layer3_outputs(2470) <= layer2_outputs(3286);
    layer3_outputs(2471) <= (layer2_outputs(477)) or (layer2_outputs(3756));
    layer3_outputs(2472) <= not((layer2_outputs(1128)) xor (layer2_outputs(4989)));
    layer3_outputs(2473) <= '1';
    layer3_outputs(2474) <= not(layer2_outputs(244)) or (layer2_outputs(2883));
    layer3_outputs(2475) <= (layer2_outputs(1321)) and not (layer2_outputs(2064));
    layer3_outputs(2476) <= not(layer2_outputs(1445)) or (layer2_outputs(2957));
    layer3_outputs(2477) <= not((layer2_outputs(4470)) and (layer2_outputs(2572)));
    layer3_outputs(2478) <= (layer2_outputs(1684)) or (layer2_outputs(2725));
    layer3_outputs(2479) <= not((layer2_outputs(3261)) and (layer2_outputs(2485)));
    layer3_outputs(2480) <= not(layer2_outputs(1277)) or (layer2_outputs(5021));
    layer3_outputs(2481) <= not(layer2_outputs(4763));
    layer3_outputs(2482) <= (layer2_outputs(5026)) or (layer2_outputs(1182));
    layer3_outputs(2483) <= (layer2_outputs(1440)) or (layer2_outputs(3823));
    layer3_outputs(2484) <= '1';
    layer3_outputs(2485) <= not(layer2_outputs(1765)) or (layer2_outputs(1894));
    layer3_outputs(2486) <= (layer2_outputs(4773)) or (layer2_outputs(3422));
    layer3_outputs(2487) <= not(layer2_outputs(3211));
    layer3_outputs(2488) <= (layer2_outputs(2705)) and (layer2_outputs(1166));
    layer3_outputs(2489) <= not((layer2_outputs(248)) or (layer2_outputs(1140)));
    layer3_outputs(2490) <= (layer2_outputs(4842)) and not (layer2_outputs(1604));
    layer3_outputs(2491) <= '1';
    layer3_outputs(2492) <= layer2_outputs(730);
    layer3_outputs(2493) <= (layer2_outputs(4492)) and not (layer2_outputs(2048));
    layer3_outputs(2494) <= not((layer2_outputs(2226)) and (layer2_outputs(3791)));
    layer3_outputs(2495) <= not(layer2_outputs(383));
    layer3_outputs(2496) <= '0';
    layer3_outputs(2497) <= not(layer2_outputs(2751)) or (layer2_outputs(3722));
    layer3_outputs(2498) <= not((layer2_outputs(2257)) and (layer2_outputs(154)));
    layer3_outputs(2499) <= not((layer2_outputs(4782)) and (layer2_outputs(3624)));
    layer3_outputs(2500) <= (layer2_outputs(4304)) and not (layer2_outputs(1285));
    layer3_outputs(2501) <= not(layer2_outputs(2815));
    layer3_outputs(2502) <= not((layer2_outputs(653)) or (layer2_outputs(1424)));
    layer3_outputs(2503) <= (layer2_outputs(1908)) and (layer2_outputs(3092));
    layer3_outputs(2504) <= layer2_outputs(3564);
    layer3_outputs(2505) <= layer2_outputs(229);
    layer3_outputs(2506) <= '1';
    layer3_outputs(2507) <= not((layer2_outputs(2245)) and (layer2_outputs(4678)));
    layer3_outputs(2508) <= (layer2_outputs(640)) and not (layer2_outputs(3305));
    layer3_outputs(2509) <= not(layer2_outputs(2191)) or (layer2_outputs(3519));
    layer3_outputs(2510) <= '1';
    layer3_outputs(2511) <= (layer2_outputs(4844)) and not (layer2_outputs(786));
    layer3_outputs(2512) <= (layer2_outputs(4863)) and not (layer2_outputs(4246));
    layer3_outputs(2513) <= (layer2_outputs(4007)) or (layer2_outputs(1711));
    layer3_outputs(2514) <= not((layer2_outputs(2044)) and (layer2_outputs(3331)));
    layer3_outputs(2515) <= not(layer2_outputs(527)) or (layer2_outputs(4166));
    layer3_outputs(2516) <= '0';
    layer3_outputs(2517) <= not((layer2_outputs(1076)) and (layer2_outputs(572)));
    layer3_outputs(2518) <= (layer2_outputs(1398)) and not (layer2_outputs(437));
    layer3_outputs(2519) <= not(layer2_outputs(3072));
    layer3_outputs(2520) <= '0';
    layer3_outputs(2521) <= not(layer2_outputs(704));
    layer3_outputs(2522) <= not((layer2_outputs(89)) or (layer2_outputs(4834)));
    layer3_outputs(2523) <= not((layer2_outputs(144)) or (layer2_outputs(4711)));
    layer3_outputs(2524) <= not((layer2_outputs(1568)) and (layer2_outputs(3792)));
    layer3_outputs(2525) <= (layer2_outputs(3706)) and not (layer2_outputs(3775));
    layer3_outputs(2526) <= not((layer2_outputs(2163)) and (layer2_outputs(17)));
    layer3_outputs(2527) <= '1';
    layer3_outputs(2528) <= '0';
    layer3_outputs(2529) <= not(layer2_outputs(211));
    layer3_outputs(2530) <= not((layer2_outputs(3209)) or (layer2_outputs(2338)));
    layer3_outputs(2531) <= not(layer2_outputs(4195));
    layer3_outputs(2532) <= not(layer2_outputs(4967)) or (layer2_outputs(2167));
    layer3_outputs(2533) <= not((layer2_outputs(5118)) or (layer2_outputs(5047)));
    layer3_outputs(2534) <= not(layer2_outputs(1729));
    layer3_outputs(2535) <= (layer2_outputs(3387)) and not (layer2_outputs(1802));
    layer3_outputs(2536) <= not(layer2_outputs(3456)) or (layer2_outputs(2577));
    layer3_outputs(2537) <= not((layer2_outputs(95)) and (layer2_outputs(506)));
    layer3_outputs(2538) <= layer2_outputs(1034);
    layer3_outputs(2539) <= not(layer2_outputs(423)) or (layer2_outputs(2552));
    layer3_outputs(2540) <= not(layer2_outputs(1028)) or (layer2_outputs(3673));
    layer3_outputs(2541) <= not((layer2_outputs(2108)) or (layer2_outputs(257)));
    layer3_outputs(2542) <= layer2_outputs(4717);
    layer3_outputs(2543) <= (layer2_outputs(250)) and (layer2_outputs(382));
    layer3_outputs(2544) <= '0';
    layer3_outputs(2545) <= (layer2_outputs(2342)) xor (layer2_outputs(820));
    layer3_outputs(2546) <= (layer2_outputs(3202)) or (layer2_outputs(475));
    layer3_outputs(2547) <= not((layer2_outputs(3959)) and (layer2_outputs(3178)));
    layer3_outputs(2548) <= not((layer2_outputs(2177)) or (layer2_outputs(396)));
    layer3_outputs(2549) <= not(layer2_outputs(2682));
    layer3_outputs(2550) <= not(layer2_outputs(4993)) or (layer2_outputs(428));
    layer3_outputs(2551) <= '0';
    layer3_outputs(2552) <= (layer2_outputs(1366)) and (layer2_outputs(2929));
    layer3_outputs(2553) <= (layer2_outputs(4923)) and not (layer2_outputs(3504));
    layer3_outputs(2554) <= not(layer2_outputs(1772)) or (layer2_outputs(722));
    layer3_outputs(2555) <= '0';
    layer3_outputs(2556) <= not((layer2_outputs(1159)) or (layer2_outputs(5055)));
    layer3_outputs(2557) <= not(layer2_outputs(326));
    layer3_outputs(2558) <= '1';
    layer3_outputs(2559) <= not((layer2_outputs(3810)) or (layer2_outputs(4699)));
    layer3_outputs(2560) <= layer2_outputs(175);
    layer3_outputs(2561) <= (layer2_outputs(2237)) and (layer2_outputs(5093));
    layer3_outputs(2562) <= not((layer2_outputs(4712)) xor (layer2_outputs(1457)));
    layer3_outputs(2563) <= (layer2_outputs(3885)) xor (layer2_outputs(1652));
    layer3_outputs(2564) <= (layer2_outputs(5041)) or (layer2_outputs(356));
    layer3_outputs(2565) <= (layer2_outputs(4478)) and not (layer2_outputs(4297));
    layer3_outputs(2566) <= '1';
    layer3_outputs(2567) <= '0';
    layer3_outputs(2568) <= not(layer2_outputs(881)) or (layer2_outputs(1237));
    layer3_outputs(2569) <= (layer2_outputs(4322)) and not (layer2_outputs(4241));
    layer3_outputs(2570) <= (layer2_outputs(2135)) and (layer2_outputs(740));
    layer3_outputs(2571) <= (layer2_outputs(115)) and not (layer2_outputs(4030));
    layer3_outputs(2572) <= not(layer2_outputs(4189));
    layer3_outputs(2573) <= not((layer2_outputs(2918)) or (layer2_outputs(1193)));
    layer3_outputs(2574) <= (layer2_outputs(4622)) and not (layer2_outputs(2447));
    layer3_outputs(2575) <= not(layer2_outputs(1881));
    layer3_outputs(2576) <= not((layer2_outputs(4021)) or (layer2_outputs(3781)));
    layer3_outputs(2577) <= not(layer2_outputs(4306)) or (layer2_outputs(4038));
    layer3_outputs(2578) <= (layer2_outputs(73)) or (layer2_outputs(4235));
    layer3_outputs(2579) <= '0';
    layer3_outputs(2580) <= not((layer2_outputs(3886)) and (layer2_outputs(4612)));
    layer3_outputs(2581) <= (layer2_outputs(5067)) and not (layer2_outputs(4857));
    layer3_outputs(2582) <= (layer2_outputs(610)) or (layer2_outputs(3158));
    layer3_outputs(2583) <= '0';
    layer3_outputs(2584) <= '0';
    layer3_outputs(2585) <= (layer2_outputs(916)) and not (layer2_outputs(2956));
    layer3_outputs(2586) <= (layer2_outputs(2876)) and (layer2_outputs(2669));
    layer3_outputs(2587) <= layer2_outputs(747);
    layer3_outputs(2588) <= not(layer2_outputs(436)) or (layer2_outputs(3015));
    layer3_outputs(2589) <= '0';
    layer3_outputs(2590) <= (layer2_outputs(1937)) and (layer2_outputs(4301));
    layer3_outputs(2591) <= '0';
    layer3_outputs(2592) <= '1';
    layer3_outputs(2593) <= not((layer2_outputs(4851)) and (layer2_outputs(3014)));
    layer3_outputs(2594) <= not((layer2_outputs(4463)) xor (layer2_outputs(67)));
    layer3_outputs(2595) <= not((layer2_outputs(1579)) and (layer2_outputs(4903)));
    layer3_outputs(2596) <= layer2_outputs(3635);
    layer3_outputs(2597) <= not((layer2_outputs(2373)) and (layer2_outputs(2317)));
    layer3_outputs(2598) <= (layer2_outputs(895)) and not (layer2_outputs(1448));
    layer3_outputs(2599) <= not(layer2_outputs(1948));
    layer3_outputs(2600) <= not((layer2_outputs(1251)) or (layer2_outputs(1584)));
    layer3_outputs(2601) <= (layer2_outputs(4790)) or (layer2_outputs(2837));
    layer3_outputs(2602) <= not(layer2_outputs(4917));
    layer3_outputs(2603) <= (layer2_outputs(64)) and (layer2_outputs(1493));
    layer3_outputs(2604) <= layer2_outputs(2232);
    layer3_outputs(2605) <= (layer2_outputs(1180)) and not (layer2_outputs(3152));
    layer3_outputs(2606) <= layer2_outputs(1658);
    layer3_outputs(2607) <= '0';
    layer3_outputs(2608) <= not((layer2_outputs(4737)) and (layer2_outputs(1158)));
    layer3_outputs(2609) <= not((layer2_outputs(2813)) or (layer2_outputs(618)));
    layer3_outputs(2610) <= not(layer2_outputs(2690)) or (layer2_outputs(1904));
    layer3_outputs(2611) <= '0';
    layer3_outputs(2612) <= (layer2_outputs(2729)) and not (layer2_outputs(856));
    layer3_outputs(2613) <= not(layer2_outputs(3625)) or (layer2_outputs(3730));
    layer3_outputs(2614) <= (layer2_outputs(4649)) and not (layer2_outputs(1388));
    layer3_outputs(2615) <= layer2_outputs(2328);
    layer3_outputs(2616) <= (layer2_outputs(2607)) and (layer2_outputs(4415));
    layer3_outputs(2617) <= layer2_outputs(2687);
    layer3_outputs(2618) <= layer2_outputs(1669);
    layer3_outputs(2619) <= '1';
    layer3_outputs(2620) <= (layer2_outputs(2861)) xor (layer2_outputs(4659));
    layer3_outputs(2621) <= not(layer2_outputs(609)) or (layer2_outputs(4295));
    layer3_outputs(2622) <= (layer2_outputs(2524)) and not (layer2_outputs(756));
    layer3_outputs(2623) <= layer2_outputs(3383);
    layer3_outputs(2624) <= '1';
    layer3_outputs(2625) <= (layer2_outputs(2801)) and not (layer2_outputs(1209));
    layer3_outputs(2626) <= not((layer2_outputs(3631)) and (layer2_outputs(4334)));
    layer3_outputs(2627) <= '0';
    layer3_outputs(2628) <= '0';
    layer3_outputs(2629) <= '0';
    layer3_outputs(2630) <= (layer2_outputs(4224)) or (layer2_outputs(1636));
    layer3_outputs(2631) <= not((layer2_outputs(2401)) and (layer2_outputs(2447)));
    layer3_outputs(2632) <= (layer2_outputs(400)) and (layer2_outputs(1958));
    layer3_outputs(2633) <= (layer2_outputs(450)) or (layer2_outputs(1473));
    layer3_outputs(2634) <= (layer2_outputs(4740)) and (layer2_outputs(1564));
    layer3_outputs(2635) <= '0';
    layer3_outputs(2636) <= '0';
    layer3_outputs(2637) <= not(layer2_outputs(2034));
    layer3_outputs(2638) <= '0';
    layer3_outputs(2639) <= (layer2_outputs(1572)) and not (layer2_outputs(2945));
    layer3_outputs(2640) <= not((layer2_outputs(3042)) and (layer2_outputs(3341)));
    layer3_outputs(2641) <= not(layer2_outputs(3096)) or (layer2_outputs(3274));
    layer3_outputs(2642) <= not(layer2_outputs(1884)) or (layer2_outputs(1176));
    layer3_outputs(2643) <= (layer2_outputs(4386)) and (layer2_outputs(4089));
    layer3_outputs(2644) <= layer2_outputs(412);
    layer3_outputs(2645) <= (layer2_outputs(3900)) or (layer2_outputs(1236));
    layer3_outputs(2646) <= not(layer2_outputs(1455)) or (layer2_outputs(2263));
    layer3_outputs(2647) <= '1';
    layer3_outputs(2648) <= (layer2_outputs(2)) or (layer2_outputs(4750));
    layer3_outputs(2649) <= not((layer2_outputs(4208)) xor (layer2_outputs(1759)));
    layer3_outputs(2650) <= layer2_outputs(2609);
    layer3_outputs(2651) <= '1';
    layer3_outputs(2652) <= not(layer2_outputs(1123));
    layer3_outputs(2653) <= layer2_outputs(2339);
    layer3_outputs(2654) <= (layer2_outputs(1504)) and (layer2_outputs(3942));
    layer3_outputs(2655) <= '0';
    layer3_outputs(2656) <= not(layer2_outputs(4560));
    layer3_outputs(2657) <= (layer2_outputs(1451)) and (layer2_outputs(1135));
    layer3_outputs(2658) <= not((layer2_outputs(900)) or (layer2_outputs(2765)));
    layer3_outputs(2659) <= (layer2_outputs(4077)) and not (layer2_outputs(3873));
    layer3_outputs(2660) <= (layer2_outputs(2603)) and not (layer2_outputs(1675));
    layer3_outputs(2661) <= not((layer2_outputs(2575)) and (layer2_outputs(2347)));
    layer3_outputs(2662) <= '1';
    layer3_outputs(2663) <= layer2_outputs(1856);
    layer3_outputs(2664) <= not(layer2_outputs(3860));
    layer3_outputs(2665) <= not(layer2_outputs(4934));
    layer3_outputs(2666) <= (layer2_outputs(2366)) or (layer2_outputs(510));
    layer3_outputs(2667) <= '1';
    layer3_outputs(2668) <= '0';
    layer3_outputs(2669) <= not((layer2_outputs(638)) or (layer2_outputs(2809)));
    layer3_outputs(2670) <= '1';
    layer3_outputs(2671) <= (layer2_outputs(2995)) and (layer2_outputs(1397));
    layer3_outputs(2672) <= (layer2_outputs(688)) and not (layer2_outputs(118));
    layer3_outputs(2673) <= not((layer2_outputs(218)) or (layer2_outputs(4769)));
    layer3_outputs(2674) <= (layer2_outputs(4199)) and not (layer2_outputs(1013));
    layer3_outputs(2675) <= '1';
    layer3_outputs(2676) <= (layer2_outputs(2510)) and not (layer2_outputs(4328));
    layer3_outputs(2677) <= '0';
    layer3_outputs(2678) <= not((layer2_outputs(4973)) and (layer2_outputs(872)));
    layer3_outputs(2679) <= (layer2_outputs(2649)) or (layer2_outputs(3167));
    layer3_outputs(2680) <= (layer2_outputs(2138)) or (layer2_outputs(3736));
    layer3_outputs(2681) <= not(layer2_outputs(1987)) or (layer2_outputs(131));
    layer3_outputs(2682) <= '1';
    layer3_outputs(2683) <= not(layer2_outputs(3531)) or (layer2_outputs(2162));
    layer3_outputs(2684) <= '0';
    layer3_outputs(2685) <= '0';
    layer3_outputs(2686) <= (layer2_outputs(2705)) and (layer2_outputs(3803));
    layer3_outputs(2687) <= (layer2_outputs(4588)) and not (layer2_outputs(4631));
    layer3_outputs(2688) <= '0';
    layer3_outputs(2689) <= layer2_outputs(4837);
    layer3_outputs(2690) <= (layer2_outputs(3962)) and (layer2_outputs(916));
    layer3_outputs(2691) <= not((layer2_outputs(1588)) and (layer2_outputs(4417)));
    layer3_outputs(2692) <= '1';
    layer3_outputs(2693) <= not(layer2_outputs(2270)) or (layer2_outputs(1297));
    layer3_outputs(2694) <= not(layer2_outputs(3721)) or (layer2_outputs(2925));
    layer3_outputs(2695) <= '1';
    layer3_outputs(2696) <= (layer2_outputs(2290)) or (layer2_outputs(1080));
    layer3_outputs(2697) <= not(layer2_outputs(185));
    layer3_outputs(2698) <= (layer2_outputs(1561)) and not (layer2_outputs(2013));
    layer3_outputs(2699) <= (layer2_outputs(3867)) or (layer2_outputs(1168));
    layer3_outputs(2700) <= layer2_outputs(3447);
    layer3_outputs(2701) <= (layer2_outputs(2424)) and (layer2_outputs(3514));
    layer3_outputs(2702) <= (layer2_outputs(4377)) and (layer2_outputs(4326));
    layer3_outputs(2703) <= not(layer2_outputs(234)) or (layer2_outputs(5096));
    layer3_outputs(2704) <= '0';
    layer3_outputs(2705) <= not((layer2_outputs(783)) and (layer2_outputs(3160)));
    layer3_outputs(2706) <= not(layer2_outputs(4018));
    layer3_outputs(2707) <= not(layer2_outputs(793));
    layer3_outputs(2708) <= not(layer2_outputs(2247));
    layer3_outputs(2709) <= (layer2_outputs(174)) and (layer2_outputs(4656));
    layer3_outputs(2710) <= layer2_outputs(2158);
    layer3_outputs(2711) <= not((layer2_outputs(1644)) or (layer2_outputs(476)));
    layer3_outputs(2712) <= (layer2_outputs(2926)) or (layer2_outputs(3488));
    layer3_outputs(2713) <= not(layer2_outputs(3866));
    layer3_outputs(2714) <= layer2_outputs(2797);
    layer3_outputs(2715) <= not(layer2_outputs(4893)) or (layer2_outputs(4620));
    layer3_outputs(2716) <= '0';
    layer3_outputs(2717) <= '1';
    layer3_outputs(2718) <= not(layer2_outputs(4580));
    layer3_outputs(2719) <= (layer2_outputs(1807)) and not (layer2_outputs(3052));
    layer3_outputs(2720) <= not((layer2_outputs(827)) or (layer2_outputs(5075)));
    layer3_outputs(2721) <= not(layer2_outputs(4337));
    layer3_outputs(2722) <= not(layer2_outputs(2787)) or (layer2_outputs(1610));
    layer3_outputs(2723) <= layer2_outputs(4450);
    layer3_outputs(2724) <= '1';
    layer3_outputs(2725) <= layer2_outputs(5030);
    layer3_outputs(2726) <= layer2_outputs(213);
    layer3_outputs(2727) <= '1';
    layer3_outputs(2728) <= not(layer2_outputs(3118));
    layer3_outputs(2729) <= layer2_outputs(812);
    layer3_outputs(2730) <= (layer2_outputs(2085)) or (layer2_outputs(4676));
    layer3_outputs(2731) <= not(layer2_outputs(1834));
    layer3_outputs(2732) <= not((layer2_outputs(1623)) and (layer2_outputs(4877)));
    layer3_outputs(2733) <= not(layer2_outputs(2753));
    layer3_outputs(2734) <= '0';
    layer3_outputs(2735) <= (layer2_outputs(4668)) or (layer2_outputs(505));
    layer3_outputs(2736) <= '0';
    layer3_outputs(2737) <= not((layer2_outputs(2910)) or (layer2_outputs(3880)));
    layer3_outputs(2738) <= layer2_outputs(4955);
    layer3_outputs(2739) <= '0';
    layer3_outputs(2740) <= (layer2_outputs(3126)) and not (layer2_outputs(2077));
    layer3_outputs(2741) <= not(layer2_outputs(4891));
    layer3_outputs(2742) <= '1';
    layer3_outputs(2743) <= '0';
    layer3_outputs(2744) <= layer2_outputs(3457);
    layer3_outputs(2745) <= not((layer2_outputs(3788)) or (layer2_outputs(1114)));
    layer3_outputs(2746) <= not(layer2_outputs(1343));
    layer3_outputs(2747) <= layer2_outputs(2203);
    layer3_outputs(2748) <= not((layer2_outputs(2516)) and (layer2_outputs(2771)));
    layer3_outputs(2749) <= not(layer2_outputs(4062)) or (layer2_outputs(2131));
    layer3_outputs(2750) <= (layer2_outputs(4635)) and not (layer2_outputs(4095));
    layer3_outputs(2751) <= '1';
    layer3_outputs(2752) <= not((layer2_outputs(3315)) or (layer2_outputs(4685)));
    layer3_outputs(2753) <= not((layer2_outputs(4537)) xor (layer2_outputs(4436)));
    layer3_outputs(2754) <= (layer2_outputs(2398)) and (layer2_outputs(2580));
    layer3_outputs(2755) <= not(layer2_outputs(2416)) or (layer2_outputs(29));
    layer3_outputs(2756) <= '0';
    layer3_outputs(2757) <= '0';
    layer3_outputs(2758) <= not(layer2_outputs(3805));
    layer3_outputs(2759) <= not(layer2_outputs(4139)) or (layer2_outputs(3882));
    layer3_outputs(2760) <= not(layer2_outputs(2672));
    layer3_outputs(2761) <= '0';
    layer3_outputs(2762) <= not((layer2_outputs(3875)) or (layer2_outputs(454)));
    layer3_outputs(2763) <= layer2_outputs(2998);
    layer3_outputs(2764) <= layer2_outputs(351);
    layer3_outputs(2765) <= (layer2_outputs(3010)) and not (layer2_outputs(3097));
    layer3_outputs(2766) <= (layer2_outputs(613)) and not (layer2_outputs(99));
    layer3_outputs(2767) <= not(layer2_outputs(4560)) or (layer2_outputs(4227));
    layer3_outputs(2768) <= '0';
    layer3_outputs(2769) <= not((layer2_outputs(1803)) or (layer2_outputs(1822)));
    layer3_outputs(2770) <= not(layer2_outputs(2448));
    layer3_outputs(2771) <= layer2_outputs(2569);
    layer3_outputs(2772) <= not(layer2_outputs(4057));
    layer3_outputs(2773) <= layer2_outputs(1833);
    layer3_outputs(2774) <= '0';
    layer3_outputs(2775) <= layer2_outputs(3547);
    layer3_outputs(2776) <= not(layer2_outputs(3824));
    layer3_outputs(2777) <= layer2_outputs(1249);
    layer3_outputs(2778) <= not(layer2_outputs(3113)) or (layer2_outputs(2328));
    layer3_outputs(2779) <= (layer2_outputs(4543)) or (layer2_outputs(2986));
    layer3_outputs(2780) <= '0';
    layer3_outputs(2781) <= layer2_outputs(2984);
    layer3_outputs(2782) <= (layer2_outputs(4260)) and (layer2_outputs(2127));
    layer3_outputs(2783) <= '1';
    layer3_outputs(2784) <= (layer2_outputs(3262)) and not (layer2_outputs(2186));
    layer3_outputs(2785) <= '0';
    layer3_outputs(2786) <= '1';
    layer3_outputs(2787) <= not(layer2_outputs(4786)) or (layer2_outputs(4462));
    layer3_outputs(2788) <= not((layer2_outputs(4709)) and (layer2_outputs(364)));
    layer3_outputs(2789) <= layer2_outputs(4952);
    layer3_outputs(2790) <= not(layer2_outputs(4477)) or (layer2_outputs(2201));
    layer3_outputs(2791) <= not(layer2_outputs(3170)) or (layer2_outputs(2930));
    layer3_outputs(2792) <= not((layer2_outputs(4245)) and (layer2_outputs(1923)));
    layer3_outputs(2793) <= not((layer2_outputs(4839)) and (layer2_outputs(3035)));
    layer3_outputs(2794) <= not((layer2_outputs(4502)) and (layer2_outputs(4965)));
    layer3_outputs(2795) <= layer2_outputs(227);
    layer3_outputs(2796) <= layer2_outputs(378);
    layer3_outputs(2797) <= layer2_outputs(790);
    layer3_outputs(2798) <= not((layer2_outputs(4156)) and (layer2_outputs(1812)));
    layer3_outputs(2799) <= not(layer2_outputs(2046));
    layer3_outputs(2800) <= not(layer2_outputs(4581)) or (layer2_outputs(2124));
    layer3_outputs(2801) <= (layer2_outputs(2715)) and (layer2_outputs(4119));
    layer3_outputs(2802) <= '1';
    layer3_outputs(2803) <= '0';
    layer3_outputs(2804) <= (layer2_outputs(2921)) and (layer2_outputs(4454));
    layer3_outputs(2805) <= not(layer2_outputs(780)) or (layer2_outputs(3659));
    layer3_outputs(2806) <= '1';
    layer3_outputs(2807) <= (layer2_outputs(1120)) and not (layer2_outputs(1136));
    layer3_outputs(2808) <= '1';
    layer3_outputs(2809) <= not(layer2_outputs(2308));
    layer3_outputs(2810) <= not(layer2_outputs(900)) or (layer2_outputs(2893));
    layer3_outputs(2811) <= '1';
    layer3_outputs(2812) <= layer2_outputs(1469);
    layer3_outputs(2813) <= (layer2_outputs(3195)) or (layer2_outputs(2983));
    layer3_outputs(2814) <= layer2_outputs(5078);
    layer3_outputs(2815) <= (layer2_outputs(1764)) and not (layer2_outputs(3249));
    layer3_outputs(2816) <= '1';
    layer3_outputs(2817) <= '1';
    layer3_outputs(2818) <= not(layer2_outputs(1801));
    layer3_outputs(2819) <= '0';
    layer3_outputs(2820) <= (layer2_outputs(516)) and (layer2_outputs(2855));
    layer3_outputs(2821) <= (layer2_outputs(3438)) and not (layer2_outputs(2870));
    layer3_outputs(2822) <= (layer2_outputs(2303)) and not (layer2_outputs(4469));
    layer3_outputs(2823) <= (layer2_outputs(3595)) and not (layer2_outputs(2854));
    layer3_outputs(2824) <= layer2_outputs(3148);
    layer3_outputs(2825) <= (layer2_outputs(5032)) or (layer2_outputs(1211));
    layer3_outputs(2826) <= not(layer2_outputs(755)) or (layer2_outputs(1724));
    layer3_outputs(2827) <= not(layer2_outputs(3521)) or (layer2_outputs(3807));
    layer3_outputs(2828) <= not((layer2_outputs(4228)) and (layer2_outputs(1662)));
    layer3_outputs(2829) <= not((layer2_outputs(2709)) and (layer2_outputs(1247)));
    layer3_outputs(2830) <= (layer2_outputs(3953)) and (layer2_outputs(1414));
    layer3_outputs(2831) <= layer2_outputs(2300);
    layer3_outputs(2832) <= not(layer2_outputs(778));
    layer3_outputs(2833) <= layer2_outputs(1507);
    layer3_outputs(2834) <= not(layer2_outputs(4641)) or (layer2_outputs(2531));
    layer3_outputs(2835) <= '0';
    layer3_outputs(2836) <= not(layer2_outputs(2785));
    layer3_outputs(2837) <= (layer2_outputs(1227)) xor (layer2_outputs(1320));
    layer3_outputs(2838) <= not(layer2_outputs(4555));
    layer3_outputs(2839) <= not(layer2_outputs(3030));
    layer3_outputs(2840) <= (layer2_outputs(2602)) and not (layer2_outputs(83));
    layer3_outputs(2841) <= '0';
    layer3_outputs(2842) <= layer2_outputs(4111);
    layer3_outputs(2843) <= not(layer2_outputs(2145)) or (layer2_outputs(2687));
    layer3_outputs(2844) <= not(layer2_outputs(673));
    layer3_outputs(2845) <= not((layer2_outputs(1970)) or (layer2_outputs(3665)));
    layer3_outputs(2846) <= not(layer2_outputs(2455)) or (layer2_outputs(4561));
    layer3_outputs(2847) <= not(layer2_outputs(2655));
    layer3_outputs(2848) <= '1';
    layer3_outputs(2849) <= (layer2_outputs(3853)) and (layer2_outputs(4102));
    layer3_outputs(2850) <= not((layer2_outputs(738)) or (layer2_outputs(4578)));
    layer3_outputs(2851) <= not(layer2_outputs(1814));
    layer3_outputs(2852) <= (layer2_outputs(4914)) or (layer2_outputs(2205));
    layer3_outputs(2853) <= (layer2_outputs(1272)) and (layer2_outputs(861));
    layer3_outputs(2854) <= layer2_outputs(1724);
    layer3_outputs(2855) <= not(layer2_outputs(4014)) or (layer2_outputs(3793));
    layer3_outputs(2856) <= '1';
    layer3_outputs(2857) <= not((layer2_outputs(2829)) or (layer2_outputs(518)));
    layer3_outputs(2858) <= '1';
    layer3_outputs(2859) <= (layer2_outputs(773)) and (layer2_outputs(5071));
    layer3_outputs(2860) <= layer2_outputs(142);
    layer3_outputs(2861) <= not((layer2_outputs(2192)) and (layer2_outputs(802)));
    layer3_outputs(2862) <= (layer2_outputs(416)) or (layer2_outputs(1826));
    layer3_outputs(2863) <= (layer2_outputs(4547)) or (layer2_outputs(2550));
    layer3_outputs(2864) <= not((layer2_outputs(390)) and (layer2_outputs(3481)));
    layer3_outputs(2865) <= '1';
    layer3_outputs(2866) <= not(layer2_outputs(3414));
    layer3_outputs(2867) <= layer2_outputs(1481);
    layer3_outputs(2868) <= layer2_outputs(4065);
    layer3_outputs(2869) <= layer2_outputs(3481);
    layer3_outputs(2870) <= '1';
    layer3_outputs(2871) <= (layer2_outputs(2359)) and (layer2_outputs(4574));
    layer3_outputs(2872) <= layer2_outputs(2713);
    layer3_outputs(2873) <= (layer2_outputs(1712)) or (layer2_outputs(825));
    layer3_outputs(2874) <= layer2_outputs(1001);
    layer3_outputs(2875) <= not((layer2_outputs(2075)) and (layer2_outputs(917)));
    layer3_outputs(2876) <= '1';
    layer3_outputs(2877) <= '0';
    layer3_outputs(2878) <= (layer2_outputs(596)) and not (layer2_outputs(3663));
    layer3_outputs(2879) <= not((layer2_outputs(197)) and (layer2_outputs(1858)));
    layer3_outputs(2880) <= layer2_outputs(2047);
    layer3_outputs(2881) <= '0';
    layer3_outputs(2882) <= not(layer2_outputs(1760));
    layer3_outputs(2883) <= not(layer2_outputs(507)) or (layer2_outputs(5092));
    layer3_outputs(2884) <= (layer2_outputs(280)) xor (layer2_outputs(3697));
    layer3_outputs(2885) <= (layer2_outputs(1630)) and (layer2_outputs(1726));
    layer3_outputs(2886) <= not(layer2_outputs(1578)) or (layer2_outputs(247));
    layer3_outputs(2887) <= (layer2_outputs(3285)) and (layer2_outputs(4284));
    layer3_outputs(2888) <= '0';
    layer3_outputs(2889) <= (layer2_outputs(1685)) and not (layer2_outputs(218));
    layer3_outputs(2890) <= not(layer2_outputs(4044));
    layer3_outputs(2891) <= (layer2_outputs(4877)) and (layer2_outputs(355));
    layer3_outputs(2892) <= not(layer2_outputs(2030)) or (layer2_outputs(3459));
    layer3_outputs(2893) <= (layer2_outputs(4500)) or (layer2_outputs(4830));
    layer3_outputs(2894) <= '0';
    layer3_outputs(2895) <= '0';
    layer3_outputs(2896) <= not(layer2_outputs(1112)) or (layer2_outputs(1863));
    layer3_outputs(2897) <= layer2_outputs(3395);
    layer3_outputs(2898) <= not(layer2_outputs(3140)) or (layer2_outputs(1639));
    layer3_outputs(2899) <= not((layer2_outputs(1969)) or (layer2_outputs(1634)));
    layer3_outputs(2900) <= not(layer2_outputs(2418)) or (layer2_outputs(2062));
    layer3_outputs(2901) <= layer2_outputs(715);
    layer3_outputs(2902) <= '0';
    layer3_outputs(2903) <= not(layer2_outputs(1190)) or (layer2_outputs(2546));
    layer3_outputs(2904) <= not(layer2_outputs(358)) or (layer2_outputs(1185));
    layer3_outputs(2905) <= (layer2_outputs(3342)) and not (layer2_outputs(4969));
    layer3_outputs(2906) <= (layer2_outputs(4222)) and not (layer2_outputs(3278));
    layer3_outputs(2907) <= not((layer2_outputs(909)) or (layer2_outputs(736)));
    layer3_outputs(2908) <= not((layer2_outputs(622)) or (layer2_outputs(1728)));
    layer3_outputs(2909) <= layer2_outputs(295);
    layer3_outputs(2910) <= layer2_outputs(149);
    layer3_outputs(2911) <= not(layer2_outputs(3467));
    layer3_outputs(2912) <= not(layer2_outputs(3370)) or (layer2_outputs(4506));
    layer3_outputs(2913) <= layer2_outputs(1626);
    layer3_outputs(2914) <= '0';
    layer3_outputs(2915) <= not(layer2_outputs(1914)) or (layer2_outputs(1164));
    layer3_outputs(2916) <= not((layer2_outputs(1197)) or (layer2_outputs(2699)));
    layer3_outputs(2917) <= (layer2_outputs(1627)) and not (layer2_outputs(330));
    layer3_outputs(2918) <= not(layer2_outputs(926)) or (layer2_outputs(3371));
    layer3_outputs(2919) <= (layer2_outputs(3835)) and (layer2_outputs(4101));
    layer3_outputs(2920) <= not(layer2_outputs(3215));
    layer3_outputs(2921) <= (layer2_outputs(3509)) and not (layer2_outputs(3613));
    layer3_outputs(2922) <= '1';
    layer3_outputs(2923) <= not(layer2_outputs(1529));
    layer3_outputs(2924) <= not(layer2_outputs(2318)) or (layer2_outputs(809));
    layer3_outputs(2925) <= layer2_outputs(233);
    layer3_outputs(2926) <= layer2_outputs(933);
    layer3_outputs(2927) <= layer2_outputs(3798);
    layer3_outputs(2928) <= not((layer2_outputs(4913)) or (layer2_outputs(3802)));
    layer3_outputs(2929) <= (layer2_outputs(3238)) or (layer2_outputs(3474));
    layer3_outputs(2930) <= not(layer2_outputs(87)) or (layer2_outputs(1446));
    layer3_outputs(2931) <= not((layer2_outputs(283)) and (layer2_outputs(3331)));
    layer3_outputs(2932) <= not((layer2_outputs(985)) or (layer2_outputs(4789)));
    layer3_outputs(2933) <= not(layer2_outputs(4510));
    layer3_outputs(2934) <= layer2_outputs(1449);
    layer3_outputs(2935) <= not((layer2_outputs(4860)) xor (layer2_outputs(1791)));
    layer3_outputs(2936) <= '0';
    layer3_outputs(2937) <= layer2_outputs(251);
    layer3_outputs(2938) <= (layer2_outputs(4423)) and not (layer2_outputs(2583));
    layer3_outputs(2939) <= (layer2_outputs(2191)) and not (layer2_outputs(3218));
    layer3_outputs(2940) <= (layer2_outputs(2058)) and not (layer2_outputs(554));
    layer3_outputs(2941) <= '1';
    layer3_outputs(2942) <= (layer2_outputs(1542)) and not (layer2_outputs(882));
    layer3_outputs(2943) <= not((layer2_outputs(2276)) and (layer2_outputs(3368)));
    layer3_outputs(2944) <= not(layer2_outputs(3479)) or (layer2_outputs(2358));
    layer3_outputs(2945) <= (layer2_outputs(1296)) and not (layer2_outputs(2194));
    layer3_outputs(2946) <= not(layer2_outputs(3219));
    layer3_outputs(2947) <= '0';
    layer3_outputs(2948) <= (layer2_outputs(3088)) and not (layer2_outputs(4055));
    layer3_outputs(2949) <= (layer2_outputs(1528)) and not (layer2_outputs(4867));
    layer3_outputs(2950) <= (layer2_outputs(241)) xor (layer2_outputs(37));
    layer3_outputs(2951) <= not(layer2_outputs(293)) or (layer2_outputs(2780));
    layer3_outputs(2952) <= not(layer2_outputs(800)) or (layer2_outputs(3563));
    layer3_outputs(2953) <= layer2_outputs(1365);
    layer3_outputs(2954) <= layer2_outputs(4269);
    layer3_outputs(2955) <= not((layer2_outputs(4409)) and (layer2_outputs(165)));
    layer3_outputs(2956) <= not((layer2_outputs(2063)) or (layer2_outputs(2459)));
    layer3_outputs(2957) <= not((layer2_outputs(1098)) or (layer2_outputs(1363)));
    layer3_outputs(2958) <= not(layer2_outputs(483));
    layer3_outputs(2959) <= not(layer2_outputs(3903)) or (layer2_outputs(2515));
    layer3_outputs(2960) <= not(layer2_outputs(746));
    layer3_outputs(2961) <= (layer2_outputs(2540)) or (layer2_outputs(549));
    layer3_outputs(2962) <= not((layer2_outputs(1259)) and (layer2_outputs(4571)));
    layer3_outputs(2963) <= layer2_outputs(1066);
    layer3_outputs(2964) <= (layer2_outputs(3244)) or (layer2_outputs(2172));
    layer3_outputs(2965) <= '0';
    layer3_outputs(2966) <= (layer2_outputs(1709)) and not (layer2_outputs(503));
    layer3_outputs(2967) <= (layer2_outputs(970)) and (layer2_outputs(3079));
    layer3_outputs(2968) <= (layer2_outputs(3000)) and not (layer2_outputs(4171));
    layer3_outputs(2969) <= (layer2_outputs(1429)) and (layer2_outputs(729));
    layer3_outputs(2970) <= '0';
    layer3_outputs(2971) <= '1';
    layer3_outputs(2972) <= layer2_outputs(2171);
    layer3_outputs(2973) <= (layer2_outputs(1521)) and (layer2_outputs(3694));
    layer3_outputs(2974) <= '1';
    layer3_outputs(2975) <= not((layer2_outputs(3731)) and (layer2_outputs(62)));
    layer3_outputs(2976) <= layer2_outputs(1810);
    layer3_outputs(2977) <= not(layer2_outputs(4999));
    layer3_outputs(2978) <= layer2_outputs(2044);
    layer3_outputs(2979) <= not((layer2_outputs(4323)) xor (layer2_outputs(3080)));
    layer3_outputs(2980) <= (layer2_outputs(927)) and not (layer2_outputs(129));
    layer3_outputs(2981) <= layer2_outputs(2639);
    layer3_outputs(2982) <= not((layer2_outputs(2439)) xor (layer2_outputs(3045)));
    layer3_outputs(2983) <= not(layer2_outputs(33));
    layer3_outputs(2984) <= not((layer2_outputs(363)) or (layer2_outputs(3626)));
    layer3_outputs(2985) <= not(layer2_outputs(4206));
    layer3_outputs(2986) <= (layer2_outputs(4192)) and (layer2_outputs(2021));
    layer3_outputs(2987) <= (layer2_outputs(4347)) xor (layer2_outputs(2666));
    layer3_outputs(2988) <= not(layer2_outputs(2829)) or (layer2_outputs(4318));
    layer3_outputs(2989) <= '0';
    layer3_outputs(2990) <= not((layer2_outputs(1455)) or (layer2_outputs(4665)));
    layer3_outputs(2991) <= layer2_outputs(4513);
    layer3_outputs(2992) <= (layer2_outputs(2654)) and not (layer2_outputs(3454));
    layer3_outputs(2993) <= not(layer2_outputs(4467)) or (layer2_outputs(3492));
    layer3_outputs(2994) <= not(layer2_outputs(2921)) or (layer2_outputs(724));
    layer3_outputs(2995) <= (layer2_outputs(529)) and not (layer2_outputs(732));
    layer3_outputs(2996) <= layer2_outputs(4883);
    layer3_outputs(2997) <= not(layer2_outputs(1202));
    layer3_outputs(2998) <= not((layer2_outputs(761)) xor (layer2_outputs(1107)));
    layer3_outputs(2999) <= not((layer2_outputs(2438)) and (layer2_outputs(1443)));
    layer3_outputs(3000) <= not((layer2_outputs(467)) or (layer2_outputs(214)));
    layer3_outputs(3001) <= not(layer2_outputs(1068));
    layer3_outputs(3002) <= layer2_outputs(1958);
    layer3_outputs(3003) <= (layer2_outputs(2282)) or (layer2_outputs(1890));
    layer3_outputs(3004) <= not((layer2_outputs(3757)) and (layer2_outputs(32)));
    layer3_outputs(3005) <= not(layer2_outputs(376)) or (layer2_outputs(2494));
    layer3_outputs(3006) <= (layer2_outputs(1043)) and not (layer2_outputs(3198));
    layer3_outputs(3007) <= layer2_outputs(555);
    layer3_outputs(3008) <= not((layer2_outputs(541)) xor (layer2_outputs(3444)));
    layer3_outputs(3009) <= layer2_outputs(3717);
    layer3_outputs(3010) <= layer2_outputs(1717);
    layer3_outputs(3011) <= not(layer2_outputs(3019)) or (layer2_outputs(1498));
    layer3_outputs(3012) <= '0';
    layer3_outputs(3013) <= (layer2_outputs(3019)) and (layer2_outputs(591));
    layer3_outputs(3014) <= '0';
    layer3_outputs(3015) <= not((layer2_outputs(3902)) xor (layer2_outputs(3282)));
    layer3_outputs(3016) <= (layer2_outputs(4826)) and (layer2_outputs(3476));
    layer3_outputs(3017) <= not((layer2_outputs(631)) and (layer2_outputs(4373)));
    layer3_outputs(3018) <= (layer2_outputs(4982)) and not (layer2_outputs(54));
    layer3_outputs(3019) <= '0';
    layer3_outputs(3020) <= (layer2_outputs(259)) and not (layer2_outputs(3369));
    layer3_outputs(3021) <= '0';
    layer3_outputs(3022) <= not(layer2_outputs(2744));
    layer3_outputs(3023) <= (layer2_outputs(2267)) xor (layer2_outputs(3540));
    layer3_outputs(3024) <= not((layer2_outputs(2563)) and (layer2_outputs(3665)));
    layer3_outputs(3025) <= not(layer2_outputs(2955));
    layer3_outputs(3026) <= (layer2_outputs(4384)) and (layer2_outputs(1822));
    layer3_outputs(3027) <= (layer2_outputs(3008)) and not (layer2_outputs(4485));
    layer3_outputs(3028) <= (layer2_outputs(1590)) or (layer2_outputs(4299));
    layer3_outputs(3029) <= not((layer2_outputs(2884)) or (layer2_outputs(3475)));
    layer3_outputs(3030) <= '1';
    layer3_outputs(3031) <= not(layer2_outputs(1918));
    layer3_outputs(3032) <= not(layer2_outputs(3129)) or (layer2_outputs(4172));
    layer3_outputs(3033) <= not((layer2_outputs(3123)) or (layer2_outputs(2599)));
    layer3_outputs(3034) <= not(layer2_outputs(1897)) or (layer2_outputs(601));
    layer3_outputs(3035) <= '1';
    layer3_outputs(3036) <= not(layer2_outputs(2906)) or (layer2_outputs(780));
    layer3_outputs(3037) <= '1';
    layer3_outputs(3038) <= not(layer2_outputs(1802)) or (layer2_outputs(82));
    layer3_outputs(3039) <= (layer2_outputs(947)) or (layer2_outputs(3936));
    layer3_outputs(3040) <= not(layer2_outputs(901));
    layer3_outputs(3041) <= (layer2_outputs(4981)) and not (layer2_outputs(3952));
    layer3_outputs(3042) <= (layer2_outputs(1382)) and not (layer2_outputs(2910));
    layer3_outputs(3043) <= (layer2_outputs(4401)) or (layer2_outputs(3629));
    layer3_outputs(3044) <= '1';
    layer3_outputs(3045) <= not((layer2_outputs(4886)) or (layer2_outputs(3512)));
    layer3_outputs(3046) <= not(layer2_outputs(2589)) or (layer2_outputs(3101));
    layer3_outputs(3047) <= not((layer2_outputs(2092)) or (layer2_outputs(1738)));
    layer3_outputs(3048) <= '0';
    layer3_outputs(3049) <= not(layer2_outputs(669));
    layer3_outputs(3050) <= not(layer2_outputs(3349)) or (layer2_outputs(3237));
    layer3_outputs(3051) <= layer2_outputs(1850);
    layer3_outputs(3052) <= '1';
    layer3_outputs(3053) <= not(layer2_outputs(3012)) or (layer2_outputs(2103));
    layer3_outputs(3054) <= (layer2_outputs(4991)) and (layer2_outputs(1070));
    layer3_outputs(3055) <= (layer2_outputs(410)) and not (layer2_outputs(4616));
    layer3_outputs(3056) <= (layer2_outputs(1064)) and not (layer2_outputs(3039));
    layer3_outputs(3057) <= not(layer2_outputs(3104)) or (layer2_outputs(2233));
    layer3_outputs(3058) <= not(layer2_outputs(4123)) or (layer2_outputs(219));
    layer3_outputs(3059) <= not((layer2_outputs(2931)) and (layer2_outputs(202)));
    layer3_outputs(3060) <= (layer2_outputs(2570)) or (layer2_outputs(4325));
    layer3_outputs(3061) <= (layer2_outputs(4117)) and (layer2_outputs(3354));
    layer3_outputs(3062) <= not(layer2_outputs(4689)) or (layer2_outputs(4203));
    layer3_outputs(3063) <= (layer2_outputs(5025)) and not (layer2_outputs(1157));
    layer3_outputs(3064) <= not(layer2_outputs(429)) or (layer2_outputs(2997));
    layer3_outputs(3065) <= layer2_outputs(2089);
    layer3_outputs(3066) <= (layer2_outputs(5027)) and not (layer2_outputs(1929));
    layer3_outputs(3067) <= (layer2_outputs(4988)) and not (layer2_outputs(1411));
    layer3_outputs(3068) <= not((layer2_outputs(4817)) and (layer2_outputs(1935)));
    layer3_outputs(3069) <= not(layer2_outputs(3955));
    layer3_outputs(3070) <= not(layer2_outputs(612));
    layer3_outputs(3071) <= not((layer2_outputs(3667)) or (layer2_outputs(1240)));
    layer3_outputs(3072) <= (layer2_outputs(1131)) and (layer2_outputs(4787));
    layer3_outputs(3073) <= not((layer2_outputs(3350)) or (layer2_outputs(4859)));
    layer3_outputs(3074) <= not(layer2_outputs(126)) or (layer2_outputs(2202));
    layer3_outputs(3075) <= (layer2_outputs(5044)) and (layer2_outputs(3830));
    layer3_outputs(3076) <= not(layer2_outputs(3258)) or (layer2_outputs(2774));
    layer3_outputs(3077) <= not(layer2_outputs(4435));
    layer3_outputs(3078) <= not(layer2_outputs(2774)) or (layer2_outputs(779));
    layer3_outputs(3079) <= '0';
    layer3_outputs(3080) <= '1';
    layer3_outputs(3081) <= '1';
    layer3_outputs(3082) <= not(layer2_outputs(3002));
    layer3_outputs(3083) <= (layer2_outputs(2940)) or (layer2_outputs(1911));
    layer3_outputs(3084) <= not((layer2_outputs(2184)) and (layer2_outputs(1589)));
    layer3_outputs(3085) <= not(layer2_outputs(967)) or (layer2_outputs(1378));
    layer3_outputs(3086) <= not(layer2_outputs(2950));
    layer3_outputs(3087) <= not((layer2_outputs(4644)) or (layer2_outputs(4474)));
    layer3_outputs(3088) <= '0';
    layer3_outputs(3089) <= (layer2_outputs(263)) or (layer2_outputs(3293));
    layer3_outputs(3090) <= not(layer2_outputs(1)) or (layer2_outputs(3933));
    layer3_outputs(3091) <= (layer2_outputs(1654)) and (layer2_outputs(3579));
    layer3_outputs(3092) <= (layer2_outputs(3417)) or (layer2_outputs(708));
    layer3_outputs(3093) <= '0';
    layer3_outputs(3094) <= layer2_outputs(2420);
    layer3_outputs(3095) <= '1';
    layer3_outputs(3096) <= not(layer2_outputs(4181)) or (layer2_outputs(3623));
    layer3_outputs(3097) <= '0';
    layer3_outputs(3098) <= not(layer2_outputs(4173)) or (layer2_outputs(1536));
    layer3_outputs(3099) <= (layer2_outputs(3810)) or (layer2_outputs(859));
    layer3_outputs(3100) <= (layer2_outputs(3776)) and not (layer2_outputs(3578));
    layer3_outputs(3101) <= layer2_outputs(1254);
    layer3_outputs(3102) <= (layer2_outputs(26)) or (layer2_outputs(1101));
    layer3_outputs(3103) <= '0';
    layer3_outputs(3104) <= (layer2_outputs(4566)) and not (layer2_outputs(281));
    layer3_outputs(3105) <= (layer2_outputs(1386)) and not (layer2_outputs(3924));
    layer3_outputs(3106) <= (layer2_outputs(2012)) and not (layer2_outputs(3658));
    layer3_outputs(3107) <= not(layer2_outputs(3132)) or (layer2_outputs(2135));
    layer3_outputs(3108) <= not(layer2_outputs(3791));
    layer3_outputs(3109) <= not(layer2_outputs(48)) or (layer2_outputs(346));
    layer3_outputs(3110) <= (layer2_outputs(417)) and (layer2_outputs(4179));
    layer3_outputs(3111) <= (layer2_outputs(1402)) and not (layer2_outputs(1170));
    layer3_outputs(3112) <= '0';
    layer3_outputs(3113) <= '1';
    layer3_outputs(3114) <= not((layer2_outputs(4244)) or (layer2_outputs(3742)));
    layer3_outputs(3115) <= layer2_outputs(2025);
    layer3_outputs(3116) <= '1';
    layer3_outputs(3117) <= (layer2_outputs(778)) and (layer2_outputs(541));
    layer3_outputs(3118) <= (layer2_outputs(1205)) and not (layer2_outputs(2752));
    layer3_outputs(3119) <= '1';
    layer3_outputs(3120) <= '0';
    layer3_outputs(3121) <= (layer2_outputs(2815)) and not (layer2_outputs(4485));
    layer3_outputs(3122) <= not((layer2_outputs(3472)) and (layer2_outputs(656)));
    layer3_outputs(3123) <= layer2_outputs(5078);
    layer3_outputs(3124) <= not((layer2_outputs(1989)) and (layer2_outputs(4472)));
    layer3_outputs(3125) <= (layer2_outputs(107)) and not (layer2_outputs(3224));
    layer3_outputs(3126) <= layer2_outputs(637);
    layer3_outputs(3127) <= not((layer2_outputs(5104)) or (layer2_outputs(4739)));
    layer3_outputs(3128) <= (layer2_outputs(948)) and (layer2_outputs(4090));
    layer3_outputs(3129) <= not(layer2_outputs(943));
    layer3_outputs(3130) <= not(layer2_outputs(3571));
    layer3_outputs(3131) <= not(layer2_outputs(78));
    layer3_outputs(3132) <= not((layer2_outputs(643)) or (layer2_outputs(492)));
    layer3_outputs(3133) <= not(layer2_outputs(4570)) or (layer2_outputs(4303));
    layer3_outputs(3134) <= layer2_outputs(3551);
    layer3_outputs(3135) <= (layer2_outputs(4340)) and not (layer2_outputs(1960));
    layer3_outputs(3136) <= '1';
    layer3_outputs(3137) <= layer2_outputs(1668);
    layer3_outputs(3138) <= (layer2_outputs(2797)) or (layer2_outputs(4699));
    layer3_outputs(3139) <= not(layer2_outputs(4559));
    layer3_outputs(3140) <= (layer2_outputs(3884)) and not (layer2_outputs(1110));
    layer3_outputs(3141) <= (layer2_outputs(3495)) or (layer2_outputs(2966));
    layer3_outputs(3142) <= not(layer2_outputs(3031));
    layer3_outputs(3143) <= not(layer2_outputs(1663)) or (layer2_outputs(1661));
    layer3_outputs(3144) <= '0';
    layer3_outputs(3145) <= not((layer2_outputs(196)) or (layer2_outputs(2510)));
    layer3_outputs(3146) <= (layer2_outputs(2080)) and not (layer2_outputs(3415));
    layer3_outputs(3147) <= (layer2_outputs(5008)) and not (layer2_outputs(3378));
    layer3_outputs(3148) <= not(layer2_outputs(3257));
    layer3_outputs(3149) <= not((layer2_outputs(3522)) or (layer2_outputs(4900)));
    layer3_outputs(3150) <= '1';
    layer3_outputs(3151) <= not(layer2_outputs(1529)) or (layer2_outputs(242));
    layer3_outputs(3152) <= (layer2_outputs(3584)) and not (layer2_outputs(3643));
    layer3_outputs(3153) <= not((layer2_outputs(3818)) or (layer2_outputs(889)));
    layer3_outputs(3154) <= not(layer2_outputs(4850)) or (layer2_outputs(2015));
    layer3_outputs(3155) <= layer2_outputs(4919);
    layer3_outputs(3156) <= '1';
    layer3_outputs(3157) <= not(layer2_outputs(4113));
    layer3_outputs(3158) <= (layer2_outputs(2206)) and not (layer2_outputs(139));
    layer3_outputs(3159) <= '1';
    layer3_outputs(3160) <= (layer2_outputs(1210)) xor (layer2_outputs(4375));
    layer3_outputs(3161) <= not(layer2_outputs(878));
    layer3_outputs(3162) <= layer2_outputs(4405);
    layer3_outputs(3163) <= '0';
    layer3_outputs(3164) <= not(layer2_outputs(2720)) or (layer2_outputs(589));
    layer3_outputs(3165) <= layer2_outputs(3200);
    layer3_outputs(3166) <= (layer2_outputs(347)) and (layer2_outputs(4150));
    layer3_outputs(3167) <= (layer2_outputs(298)) and not (layer2_outputs(697));
    layer3_outputs(3168) <= layer2_outputs(2593);
    layer3_outputs(3169) <= '1';
    layer3_outputs(3170) <= not(layer2_outputs(534));
    layer3_outputs(3171) <= (layer2_outputs(3310)) or (layer2_outputs(4363));
    layer3_outputs(3172) <= (layer2_outputs(1791)) or (layer2_outputs(1153));
    layer3_outputs(3173) <= (layer2_outputs(1696)) and not (layer2_outputs(3512));
    layer3_outputs(3174) <= '1';
    layer3_outputs(3175) <= not((layer2_outputs(3378)) and (layer2_outputs(2964)));
    layer3_outputs(3176) <= '0';
    layer3_outputs(3177) <= not(layer2_outputs(4396));
    layer3_outputs(3178) <= '0';
    layer3_outputs(3179) <= (layer2_outputs(4385)) and not (layer2_outputs(4895));
    layer3_outputs(3180) <= (layer2_outputs(397)) and not (layer2_outputs(3628));
    layer3_outputs(3181) <= (layer2_outputs(3326)) and not (layer2_outputs(4538));
    layer3_outputs(3182) <= layer2_outputs(3692);
    layer3_outputs(3183) <= not(layer2_outputs(682));
    layer3_outputs(3184) <= (layer2_outputs(2704)) and not (layer2_outputs(3880));
    layer3_outputs(3185) <= (layer2_outputs(4558)) or (layer2_outputs(2219));
    layer3_outputs(3186) <= '1';
    layer3_outputs(3187) <= not((layer2_outputs(201)) or (layer2_outputs(5053)));
    layer3_outputs(3188) <= (layer2_outputs(4099)) xor (layer2_outputs(3383));
    layer3_outputs(3189) <= not(layer2_outputs(2558));
    layer3_outputs(3190) <= (layer2_outputs(3676)) and not (layer2_outputs(4361));
    layer3_outputs(3191) <= (layer2_outputs(1916)) or (layer2_outputs(3252));
    layer3_outputs(3192) <= '0';
    layer3_outputs(3193) <= not((layer2_outputs(414)) and (layer2_outputs(2694)));
    layer3_outputs(3194) <= '0';
    layer3_outputs(3195) <= not((layer2_outputs(1371)) and (layer2_outputs(4020)));
    layer3_outputs(3196) <= not(layer2_outputs(1006)) or (layer2_outputs(2454));
    layer3_outputs(3197) <= layer2_outputs(4342);
    layer3_outputs(3198) <= (layer2_outputs(1049)) and not (layer2_outputs(477));
    layer3_outputs(3199) <= not((layer2_outputs(2869)) or (layer2_outputs(4823)));
    layer3_outputs(3200) <= (layer2_outputs(3418)) or (layer2_outputs(4225));
    layer3_outputs(3201) <= (layer2_outputs(3431)) and not (layer2_outputs(4368));
    layer3_outputs(3202) <= '1';
    layer3_outputs(3203) <= not(layer2_outputs(2608));
    layer3_outputs(3204) <= not(layer2_outputs(3587)) or (layer2_outputs(2003));
    layer3_outputs(3205) <= not(layer2_outputs(3974)) or (layer2_outputs(2471));
    layer3_outputs(3206) <= not(layer2_outputs(846)) or (layer2_outputs(2136));
    layer3_outputs(3207) <= not(layer2_outputs(3114)) or (layer2_outputs(4299));
    layer3_outputs(3208) <= (layer2_outputs(4228)) and not (layer2_outputs(2054));
    layer3_outputs(3209) <= not(layer2_outputs(4132));
    layer3_outputs(3210) <= not(layer2_outputs(2277)) or (layer2_outputs(1201));
    layer3_outputs(3211) <= (layer2_outputs(2340)) xor (layer2_outputs(2382));
    layer3_outputs(3212) <= (layer2_outputs(4176)) and not (layer2_outputs(3337));
    layer3_outputs(3213) <= '1';
    layer3_outputs(3214) <= '0';
    layer3_outputs(3215) <= not(layer2_outputs(3508)) or (layer2_outputs(1574));
    layer3_outputs(3216) <= '1';
    layer3_outputs(3217) <= not(layer2_outputs(4143)) or (layer2_outputs(4040));
    layer3_outputs(3218) <= '0';
    layer3_outputs(3219) <= (layer2_outputs(2721)) and not (layer2_outputs(154));
    layer3_outputs(3220) <= not(layer2_outputs(257));
    layer3_outputs(3221) <= '1';
    layer3_outputs(3222) <= not(layer2_outputs(1818)) or (layer2_outputs(568));
    layer3_outputs(3223) <= not((layer2_outputs(1286)) and (layer2_outputs(2057)));
    layer3_outputs(3224) <= layer2_outputs(3839);
    layer3_outputs(3225) <= not(layer2_outputs(4985)) or (layer2_outputs(1276));
    layer3_outputs(3226) <= not(layer2_outputs(3568));
    layer3_outputs(3227) <= not((layer2_outputs(805)) or (layer2_outputs(693)));
    layer3_outputs(3228) <= (layer2_outputs(2680)) and (layer2_outputs(660));
    layer3_outputs(3229) <= (layer2_outputs(1375)) and not (layer2_outputs(1673));
    layer3_outputs(3230) <= not(layer2_outputs(2220));
    layer3_outputs(3231) <= (layer2_outputs(3773)) and not (layer2_outputs(3117));
    layer3_outputs(3232) <= '1';
    layer3_outputs(3233) <= not((layer2_outputs(138)) or (layer2_outputs(1977)));
    layer3_outputs(3234) <= layer2_outputs(3103);
    layer3_outputs(3235) <= not(layer2_outputs(82));
    layer3_outputs(3236) <= not((layer2_outputs(526)) and (layer2_outputs(502)));
    layer3_outputs(3237) <= not((layer2_outputs(1274)) or (layer2_outputs(2378)));
    layer3_outputs(3238) <= (layer2_outputs(2630)) or (layer2_outputs(2839));
    layer3_outputs(3239) <= '1';
    layer3_outputs(3240) <= layer2_outputs(2137);
    layer3_outputs(3241) <= '0';
    layer3_outputs(3242) <= not(layer2_outputs(4280));
    layer3_outputs(3243) <= not((layer2_outputs(1889)) and (layer2_outputs(1778)));
    layer3_outputs(3244) <= not((layer2_outputs(3226)) or (layer2_outputs(2778)));
    layer3_outputs(3245) <= not(layer2_outputs(1635));
    layer3_outputs(3246) <= not((layer2_outputs(1023)) and (layer2_outputs(254)));
    layer3_outputs(3247) <= (layer2_outputs(753)) and (layer2_outputs(2241));
    layer3_outputs(3248) <= '0';
    layer3_outputs(3249) <= not(layer2_outputs(471)) or (layer2_outputs(3032));
    layer3_outputs(3250) <= not(layer2_outputs(4508));
    layer3_outputs(3251) <= not(layer2_outputs(2407));
    layer3_outputs(3252) <= not(layer2_outputs(2796)) or (layer2_outputs(4726));
    layer3_outputs(3253) <= '0';
    layer3_outputs(3254) <= '1';
    layer3_outputs(3255) <= (layer2_outputs(4514)) or (layer2_outputs(3589));
    layer3_outputs(3256) <= not((layer2_outputs(4660)) and (layer2_outputs(2475)));
    layer3_outputs(3257) <= (layer2_outputs(4039)) or (layer2_outputs(252));
    layer3_outputs(3258) <= '0';
    layer3_outputs(3259) <= not(layer2_outputs(2946)) or (layer2_outputs(3314));
    layer3_outputs(3260) <= layer2_outputs(4700);
    layer3_outputs(3261) <= '1';
    layer3_outputs(3262) <= (layer2_outputs(2861)) and not (layer2_outputs(3067));
    layer3_outputs(3263) <= not((layer2_outputs(4870)) or (layer2_outputs(2684)));
    layer3_outputs(3264) <= '0';
    layer3_outputs(3265) <= not(layer2_outputs(3712)) or (layer2_outputs(4447));
    layer3_outputs(3266) <= not(layer2_outputs(3820)) or (layer2_outputs(1827));
    layer3_outputs(3267) <= not(layer2_outputs(2734)) or (layer2_outputs(2076));
    layer3_outputs(3268) <= not(layer2_outputs(5103));
    layer3_outputs(3269) <= (layer2_outputs(1675)) and not (layer2_outputs(3131));
    layer3_outputs(3270) <= (layer2_outputs(1489)) or (layer2_outputs(3268));
    layer3_outputs(3271) <= not(layer2_outputs(3175));
    layer3_outputs(3272) <= not((layer2_outputs(2178)) and (layer2_outputs(339)));
    layer3_outputs(3273) <= (layer2_outputs(4481)) or (layer2_outputs(2011));
    layer3_outputs(3274) <= layer2_outputs(2136);
    layer3_outputs(3275) <= (layer2_outputs(2082)) and (layer2_outputs(4876));
    layer3_outputs(3276) <= (layer2_outputs(2476)) and not (layer2_outputs(2975));
    layer3_outputs(3277) <= not((layer2_outputs(4777)) or (layer2_outputs(3289)));
    layer3_outputs(3278) <= not(layer2_outputs(1911)) or (layer2_outputs(3206));
    layer3_outputs(3279) <= (layer2_outputs(3876)) and not (layer2_outputs(3017));
    layer3_outputs(3280) <= (layer2_outputs(1637)) and (layer2_outputs(2926));
    layer3_outputs(3281) <= (layer2_outputs(4822)) and not (layer2_outputs(2437));
    layer3_outputs(3282) <= (layer2_outputs(2979)) and not (layer2_outputs(2563));
    layer3_outputs(3283) <= '1';
    layer3_outputs(3284) <= not(layer2_outputs(2060));
    layer3_outputs(3285) <= not(layer2_outputs(2852));
    layer3_outputs(3286) <= '0';
    layer3_outputs(3287) <= layer2_outputs(1471);
    layer3_outputs(3288) <= layer2_outputs(5112);
    layer3_outputs(3289) <= '0';
    layer3_outputs(3290) <= (layer2_outputs(1043)) and not (layer2_outputs(2476));
    layer3_outputs(3291) <= layer2_outputs(415);
    layer3_outputs(3292) <= not(layer2_outputs(1136));
    layer3_outputs(3293) <= (layer2_outputs(2438)) and not (layer2_outputs(1648));
    layer3_outputs(3294) <= (layer2_outputs(4546)) and (layer2_outputs(2995));
    layer3_outputs(3295) <= (layer2_outputs(3996)) and not (layer2_outputs(2037));
    layer3_outputs(3296) <= layer2_outputs(4832);
    layer3_outputs(3297) <= (layer2_outputs(4724)) and (layer2_outputs(4204));
    layer3_outputs(3298) <= '1';
    layer3_outputs(3299) <= not((layer2_outputs(3983)) or (layer2_outputs(1401)));
    layer3_outputs(3300) <= not(layer2_outputs(535)) or (layer2_outputs(594));
    layer3_outputs(3301) <= (layer2_outputs(1611)) and (layer2_outputs(4436));
    layer3_outputs(3302) <= not((layer2_outputs(2357)) and (layer2_outputs(191)));
    layer3_outputs(3303) <= (layer2_outputs(3711)) and not (layer2_outputs(3987));
    layer3_outputs(3304) <= (layer2_outputs(891)) and (layer2_outputs(4377));
    layer3_outputs(3305) <= (layer2_outputs(1326)) and not (layer2_outputs(35));
    layer3_outputs(3306) <= not(layer2_outputs(4086));
    layer3_outputs(3307) <= (layer2_outputs(677)) and not (layer2_outputs(3716));
    layer3_outputs(3308) <= '0';
    layer3_outputs(3309) <= not(layer2_outputs(3580));
    layer3_outputs(3310) <= not(layer2_outputs(293));
    layer3_outputs(3311) <= (layer2_outputs(3479)) and (layer2_outputs(3731));
    layer3_outputs(3312) <= '0';
    layer3_outputs(3313) <= not(layer2_outputs(3672)) or (layer2_outputs(1055));
    layer3_outputs(3314) <= not(layer2_outputs(4944));
    layer3_outputs(3315) <= not((layer2_outputs(3636)) or (layer2_outputs(3942)));
    layer3_outputs(3316) <= '1';
    layer3_outputs(3317) <= layer2_outputs(3502);
    layer3_outputs(3318) <= not(layer2_outputs(133)) or (layer2_outputs(2924));
    layer3_outputs(3319) <= '0';
    layer3_outputs(3320) <= (layer2_outputs(2724)) and not (layer2_outputs(2965));
    layer3_outputs(3321) <= (layer2_outputs(2564)) or (layer2_outputs(3469));
    layer3_outputs(3322) <= not(layer2_outputs(2457));
    layer3_outputs(3323) <= (layer2_outputs(990)) and (layer2_outputs(4985));
    layer3_outputs(3324) <= not((layer2_outputs(4114)) or (layer2_outputs(1330)));
    layer3_outputs(3325) <= not(layer2_outputs(3390)) or (layer2_outputs(3501));
    layer3_outputs(3326) <= not((layer2_outputs(527)) and (layer2_outputs(1121)));
    layer3_outputs(3327) <= not(layer2_outputs(2716));
    layer3_outputs(3328) <= (layer2_outputs(1091)) and not (layer2_outputs(2669));
    layer3_outputs(3329) <= (layer2_outputs(4752)) and (layer2_outputs(2018));
    layer3_outputs(3330) <= layer2_outputs(800);
    layer3_outputs(3331) <= layer2_outputs(5019);
    layer3_outputs(3332) <= not(layer2_outputs(847));
    layer3_outputs(3333) <= not(layer2_outputs(2465));
    layer3_outputs(3334) <= not((layer2_outputs(1244)) and (layer2_outputs(4530)));
    layer3_outputs(3335) <= '0';
    layer3_outputs(3336) <= not((layer2_outputs(1164)) or (layer2_outputs(1381)));
    layer3_outputs(3337) <= (layer2_outputs(3435)) and not (layer2_outputs(941));
    layer3_outputs(3338) <= (layer2_outputs(4995)) or (layer2_outputs(2528));
    layer3_outputs(3339) <= not(layer2_outputs(860));
    layer3_outputs(3340) <= '1';
    layer3_outputs(3341) <= (layer2_outputs(1315)) and (layer2_outputs(4180));
    layer3_outputs(3342) <= (layer2_outputs(1833)) and not (layer2_outputs(399));
    layer3_outputs(3343) <= (layer2_outputs(1041)) and (layer2_outputs(1550));
    layer3_outputs(3344) <= '1';
    layer3_outputs(3345) <= not(layer2_outputs(4141));
    layer3_outputs(3346) <= (layer2_outputs(924)) and not (layer2_outputs(3559));
    layer3_outputs(3347) <= not(layer2_outputs(2117));
    layer3_outputs(3348) <= not(layer2_outputs(228));
    layer3_outputs(3349) <= not(layer2_outputs(4693));
    layer3_outputs(3350) <= '0';
    layer3_outputs(3351) <= (layer2_outputs(835)) and not (layer2_outputs(4307));
    layer3_outputs(3352) <= layer2_outputs(141);
    layer3_outputs(3353) <= (layer2_outputs(4852)) and not (layer2_outputs(4687));
    layer3_outputs(3354) <= layer2_outputs(4208);
    layer3_outputs(3355) <= not((layer2_outputs(1088)) or (layer2_outputs(4063)));
    layer3_outputs(3356) <= not(layer2_outputs(4414));
    layer3_outputs(3357) <= not(layer2_outputs(2323));
    layer3_outputs(3358) <= not(layer2_outputs(966));
    layer3_outputs(3359) <= not(layer2_outputs(2235));
    layer3_outputs(3360) <= (layer2_outputs(4207)) xor (layer2_outputs(3749));
    layer3_outputs(3361) <= '1';
    layer3_outputs(3362) <= '0';
    layer3_outputs(3363) <= not((layer2_outputs(328)) and (layer2_outputs(656)));
    layer3_outputs(3364) <= not((layer2_outputs(612)) or (layer2_outputs(1923)));
    layer3_outputs(3365) <= (layer2_outputs(2105)) and not (layer2_outputs(4654));
    layer3_outputs(3366) <= (layer2_outputs(2207)) or (layer2_outputs(1638));
    layer3_outputs(3367) <= not((layer2_outputs(3316)) and (layer2_outputs(1430)));
    layer3_outputs(3368) <= not(layer2_outputs(1819)) or (layer2_outputs(2149));
    layer3_outputs(3369) <= (layer2_outputs(4207)) and not (layer2_outputs(1734));
    layer3_outputs(3370) <= (layer2_outputs(2679)) or (layer2_outputs(1941));
    layer3_outputs(3371) <= (layer2_outputs(256)) or (layer2_outputs(3194));
    layer3_outputs(3372) <= '0';
    layer3_outputs(3373) <= not(layer2_outputs(2980));
    layer3_outputs(3374) <= not(layer2_outputs(546)) or (layer2_outputs(613));
    layer3_outputs(3375) <= not(layer2_outputs(4010));
    layer3_outputs(3376) <= '1';
    layer3_outputs(3377) <= (layer2_outputs(2578)) and (layer2_outputs(3401));
    layer3_outputs(3378) <= not(layer2_outputs(4266)) or (layer2_outputs(1268));
    layer3_outputs(3379) <= (layer2_outputs(1979)) xor (layer2_outputs(2952));
    layer3_outputs(3380) <= (layer2_outputs(2419)) and (layer2_outputs(1618));
    layer3_outputs(3381) <= (layer2_outputs(102)) and not (layer2_outputs(190));
    layer3_outputs(3382) <= not(layer2_outputs(3006));
    layer3_outputs(3383) <= (layer2_outputs(2657)) and (layer2_outputs(846));
    layer3_outputs(3384) <= (layer2_outputs(1765)) and (layer2_outputs(3461));
    layer3_outputs(3385) <= not(layer2_outputs(2880)) or (layer2_outputs(380));
    layer3_outputs(3386) <= '1';
    layer3_outputs(3387) <= layer2_outputs(2385);
    layer3_outputs(3388) <= (layer2_outputs(3579)) and not (layer2_outputs(864));
    layer3_outputs(3389) <= (layer2_outputs(4368)) or (layer2_outputs(2871));
    layer3_outputs(3390) <= not(layer2_outputs(1210));
    layer3_outputs(3391) <= not(layer2_outputs(830)) or (layer2_outputs(1249));
    layer3_outputs(3392) <= not((layer2_outputs(862)) or (layer2_outputs(24)));
    layer3_outputs(3393) <= (layer2_outputs(1504)) and not (layer2_outputs(1312));
    layer3_outputs(3394) <= '0';
    layer3_outputs(3395) <= (layer2_outputs(4692)) and not (layer2_outputs(3689));
    layer3_outputs(3396) <= '0';
    layer3_outputs(3397) <= (layer2_outputs(999)) and (layer2_outputs(3376));
    layer3_outputs(3398) <= not(layer2_outputs(1694)) or (layer2_outputs(430));
    layer3_outputs(3399) <= (layer2_outputs(3978)) and not (layer2_outputs(1113));
    layer3_outputs(3400) <= layer2_outputs(2644);
    layer3_outputs(3401) <= not((layer2_outputs(1582)) or (layer2_outputs(2170)));
    layer3_outputs(3402) <= layer2_outputs(1011);
    layer3_outputs(3403) <= (layer2_outputs(1749)) and not (layer2_outputs(5072));
    layer3_outputs(3404) <= (layer2_outputs(3681)) and not (layer2_outputs(1245));
    layer3_outputs(3405) <= '1';
    layer3_outputs(3406) <= (layer2_outputs(4582)) and (layer2_outputs(3543));
    layer3_outputs(3407) <= (layer2_outputs(3623)) and not (layer2_outputs(5077));
    layer3_outputs(3408) <= not((layer2_outputs(4770)) and (layer2_outputs(1640)));
    layer3_outputs(3409) <= not((layer2_outputs(5113)) xor (layer2_outputs(4055)));
    layer3_outputs(3410) <= (layer2_outputs(4012)) and not (layer2_outputs(3844));
    layer3_outputs(3411) <= layer2_outputs(68);
    layer3_outputs(3412) <= not(layer2_outputs(4947)) or (layer2_outputs(4169));
    layer3_outputs(3413) <= not(layer2_outputs(4986)) or (layer2_outputs(1124));
    layer3_outputs(3414) <= layer2_outputs(2943);
    layer3_outputs(3415) <= not((layer2_outputs(1495)) or (layer2_outputs(4502)));
    layer3_outputs(3416) <= layer2_outputs(4605);
    layer3_outputs(3417) <= not(layer2_outputs(3910)) or (layer2_outputs(2018));
    layer3_outputs(3418) <= not(layer2_outputs(1961)) or (layer2_outputs(3504));
    layer3_outputs(3419) <= (layer2_outputs(4275)) or (layer2_outputs(3039));
    layer3_outputs(3420) <= layer2_outputs(555);
    layer3_outputs(3421) <= (layer2_outputs(582)) and not (layer2_outputs(3317));
    layer3_outputs(3422) <= not((layer2_outputs(3646)) or (layer2_outputs(4902)));
    layer3_outputs(3423) <= layer2_outputs(1468);
    layer3_outputs(3424) <= not((layer2_outputs(744)) and (layer2_outputs(1380)));
    layer3_outputs(3425) <= not((layer2_outputs(4176)) and (layer2_outputs(1895)));
    layer3_outputs(3426) <= (layer2_outputs(5069)) and not (layer2_outputs(936));
    layer3_outputs(3427) <= not((layer2_outputs(3121)) and (layer2_outputs(1111)));
    layer3_outputs(3428) <= not(layer2_outputs(424)) or (layer2_outputs(4704));
    layer3_outputs(3429) <= not((layer2_outputs(739)) and (layer2_outputs(4624)));
    layer3_outputs(3430) <= not(layer2_outputs(5090)) or (layer2_outputs(4835));
    layer3_outputs(3431) <= '0';
    layer3_outputs(3432) <= layer2_outputs(2779);
    layer3_outputs(3433) <= (layer2_outputs(1319)) xor (layer2_outputs(4776));
    layer3_outputs(3434) <= not((layer2_outputs(4528)) and (layer2_outputs(791)));
    layer3_outputs(3435) <= '0';
    layer3_outputs(3436) <= not(layer2_outputs(1451)) or (layer2_outputs(4531));
    layer3_outputs(3437) <= not((layer2_outputs(972)) or (layer2_outputs(3109)));
    layer3_outputs(3438) <= layer2_outputs(2901);
    layer3_outputs(3439) <= not(layer2_outputs(915));
    layer3_outputs(3440) <= (layer2_outputs(3225)) or (layer2_outputs(2384));
    layer3_outputs(3441) <= layer2_outputs(2095);
    layer3_outputs(3442) <= (layer2_outputs(1158)) and (layer2_outputs(3590));
    layer3_outputs(3443) <= '1';
    layer3_outputs(3444) <= '1';
    layer3_outputs(3445) <= '0';
    layer3_outputs(3446) <= not((layer2_outputs(1885)) or (layer2_outputs(4353)));
    layer3_outputs(3447) <= '0';
    layer3_outputs(3448) <= (layer2_outputs(2005)) or (layer2_outputs(4504));
    layer3_outputs(3449) <= not(layer2_outputs(5006)) or (layer2_outputs(5079));
    layer3_outputs(3450) <= layer2_outputs(2065);
    layer3_outputs(3451) <= '1';
    layer3_outputs(3452) <= (layer2_outputs(3120)) and not (layer2_outputs(4512));
    layer3_outputs(3453) <= not(layer2_outputs(4675)) or (layer2_outputs(1755));
    layer3_outputs(3454) <= not(layer2_outputs(2885)) or (layer2_outputs(4638));
    layer3_outputs(3455) <= (layer2_outputs(1597)) or (layer2_outputs(1233));
    layer3_outputs(3456) <= (layer2_outputs(4419)) and not (layer2_outputs(3640));
    layer3_outputs(3457) <= '0';
    layer3_outputs(3458) <= '1';
    layer3_outputs(3459) <= '1';
    layer3_outputs(3460) <= not(layer2_outputs(1719)) or (layer2_outputs(757));
    layer3_outputs(3461) <= not(layer2_outputs(119)) or (layer2_outputs(1349));
    layer3_outputs(3462) <= '0';
    layer3_outputs(3463) <= not((layer2_outputs(1740)) and (layer2_outputs(2101)));
    layer3_outputs(3464) <= not(layer2_outputs(1515)) or (layer2_outputs(26));
    layer3_outputs(3465) <= layer2_outputs(3147);
    layer3_outputs(3466) <= '1';
    layer3_outputs(3467) <= (layer2_outputs(4315)) and not (layer2_outputs(195));
    layer3_outputs(3468) <= not(layer2_outputs(2502)) or (layer2_outputs(974));
    layer3_outputs(3469) <= not((layer2_outputs(4239)) and (layer2_outputs(4861)));
    layer3_outputs(3470) <= '0';
    layer3_outputs(3471) <= (layer2_outputs(2914)) or (layer2_outputs(2472));
    layer3_outputs(3472) <= not((layer2_outputs(2610)) or (layer2_outputs(1559)));
    layer3_outputs(3473) <= not((layer2_outputs(798)) and (layer2_outputs(1594)));
    layer3_outputs(3474) <= layer2_outputs(444);
    layer3_outputs(3475) <= (layer2_outputs(4300)) or (layer2_outputs(2498));
    layer3_outputs(3476) <= '0';
    layer3_outputs(3477) <= not((layer2_outputs(2627)) and (layer2_outputs(304)));
    layer3_outputs(3478) <= '0';
    layer3_outputs(3479) <= (layer2_outputs(4881)) and not (layer2_outputs(3922));
    layer3_outputs(3480) <= not(layer2_outputs(3626)) or (layer2_outputs(969));
    layer3_outputs(3481) <= not(layer2_outputs(1467)) or (layer2_outputs(4353));
    layer3_outputs(3482) <= not(layer2_outputs(958));
    layer3_outputs(3483) <= (layer2_outputs(3671)) and (layer2_outputs(168));
    layer3_outputs(3484) <= not((layer2_outputs(3864)) and (layer2_outputs(2863)));
    layer3_outputs(3485) <= (layer2_outputs(989)) and not (layer2_outputs(1004));
    layer3_outputs(3486) <= not(layer2_outputs(974));
    layer3_outputs(3487) <= not(layer2_outputs(1866)) or (layer2_outputs(1464));
    layer3_outputs(3488) <= '1';
    layer3_outputs(3489) <= not(layer2_outputs(4015));
    layer3_outputs(3490) <= (layer2_outputs(3333)) and not (layer2_outputs(308));
    layer3_outputs(3491) <= layer2_outputs(2887);
    layer3_outputs(3492) <= not((layer2_outputs(130)) and (layer2_outputs(3068)));
    layer3_outputs(3493) <= not((layer2_outputs(4688)) or (layer2_outputs(3303)));
    layer3_outputs(3494) <= (layer2_outputs(983)) and not (layer2_outputs(1145));
    layer3_outputs(3495) <= not(layer2_outputs(1781));
    layer3_outputs(3496) <= not(layer2_outputs(4573)) or (layer2_outputs(3735));
    layer3_outputs(3497) <= (layer2_outputs(2555)) and not (layer2_outputs(4840));
    layer3_outputs(3498) <= not((layer2_outputs(1327)) or (layer2_outputs(3321)));
    layer3_outputs(3499) <= layer2_outputs(1916);
    layer3_outputs(3500) <= layer2_outputs(4245);
    layer3_outputs(3501) <= (layer2_outputs(4557)) and not (layer2_outputs(2707));
    layer3_outputs(3502) <= (layer2_outputs(2614)) and not (layer2_outputs(714));
    layer3_outputs(3503) <= not((layer2_outputs(1142)) or (layer2_outputs(2202)));
    layer3_outputs(3504) <= not((layer2_outputs(4503)) or (layer2_outputs(426)));
    layer3_outputs(3505) <= not(layer2_outputs(4086)) or (layer2_outputs(855));
    layer3_outputs(3506) <= (layer2_outputs(3379)) and not (layer2_outputs(328));
    layer3_outputs(3507) <= '1';
    layer3_outputs(3508) <= layer2_outputs(1271);
    layer3_outputs(3509) <= not(layer2_outputs(2512)) or (layer2_outputs(1256));
    layer3_outputs(3510) <= not(layer2_outputs(2330));
    layer3_outputs(3511) <= (layer2_outputs(2379)) and (layer2_outputs(3013));
    layer3_outputs(3512) <= (layer2_outputs(382)) and not (layer2_outputs(1581));
    layer3_outputs(3513) <= not(layer2_outputs(704));
    layer3_outputs(3514) <= (layer2_outputs(2702)) and (layer2_outputs(2333));
    layer3_outputs(3515) <= '0';
    layer3_outputs(3516) <= layer2_outputs(2656);
    layer3_outputs(3517) <= (layer2_outputs(3151)) and not (layer2_outputs(1485));
    layer3_outputs(3518) <= not(layer2_outputs(2455));
    layer3_outputs(3519) <= (layer2_outputs(868)) and not (layer2_outputs(2301));
    layer3_outputs(3520) <= '0';
    layer3_outputs(3521) <= (layer2_outputs(1196)) or (layer2_outputs(3690));
    layer3_outputs(3522) <= not(layer2_outputs(2128)) or (layer2_outputs(150));
    layer3_outputs(3523) <= not(layer2_outputs(5029)) or (layer2_outputs(565));
    layer3_outputs(3524) <= layer2_outputs(1583);
    layer3_outputs(3525) <= '0';
    layer3_outputs(3526) <= '0';
    layer3_outputs(3527) <= '0';
    layer3_outputs(3528) <= not(layer2_outputs(430)) or (layer2_outputs(2990));
    layer3_outputs(3529) <= (layer2_outputs(568)) or (layer2_outputs(2355));
    layer3_outputs(3530) <= (layer2_outputs(1676)) and (layer2_outputs(57));
    layer3_outputs(3531) <= (layer2_outputs(1764)) and not (layer2_outputs(1775));
    layer3_outputs(3532) <= '0';
    layer3_outputs(3533) <= layer2_outputs(2470);
    layer3_outputs(3534) <= not((layer2_outputs(3286)) xor (layer2_outputs(1316)));
    layer3_outputs(3535) <= (layer2_outputs(2908)) and (layer2_outputs(4984));
    layer3_outputs(3536) <= not(layer2_outputs(4534)) or (layer2_outputs(4884));
    layer3_outputs(3537) <= '0';
    layer3_outputs(3538) <= '0';
    layer3_outputs(3539) <= not(layer2_outputs(2336));
    layer3_outputs(3540) <= not(layer2_outputs(810));
    layer3_outputs(3541) <= (layer2_outputs(2143)) and not (layer2_outputs(3690));
    layer3_outputs(3542) <= '1';
    layer3_outputs(3543) <= '0';
    layer3_outputs(3544) <= not(layer2_outputs(135)) or (layer2_outputs(16));
    layer3_outputs(3545) <= not(layer2_outputs(3545));
    layer3_outputs(3546) <= (layer2_outputs(1647)) and not (layer2_outputs(3287));
    layer3_outputs(3547) <= (layer2_outputs(3404)) and not (layer2_outputs(923));
    layer3_outputs(3548) <= (layer2_outputs(4201)) or (layer2_outputs(3388));
    layer3_outputs(3549) <= '1';
    layer3_outputs(3550) <= '1';
    layer3_outputs(3551) <= not(layer2_outputs(4808)) or (layer2_outputs(87));
    layer3_outputs(3552) <= not(layer2_outputs(2742));
    layer3_outputs(3553) <= layer2_outputs(2865);
    layer3_outputs(3554) <= (layer2_outputs(2905)) and not (layer2_outputs(1771));
    layer3_outputs(3555) <= layer2_outputs(2729);
    layer3_outputs(3556) <= (layer2_outputs(2873)) or (layer2_outputs(2746));
    layer3_outputs(3557) <= layer2_outputs(4728);
    layer3_outputs(3558) <= not(layer2_outputs(3093));
    layer3_outputs(3559) <= not(layer2_outputs(985));
    layer3_outputs(3560) <= not((layer2_outputs(747)) and (layer2_outputs(3423)));
    layer3_outputs(3561) <= '1';
    layer3_outputs(3562) <= not((layer2_outputs(1359)) or (layer2_outputs(1191)));
    layer3_outputs(3563) <= layer2_outputs(1116);
    layer3_outputs(3564) <= layer2_outputs(1990);
    layer3_outputs(3565) <= (layer2_outputs(3917)) and not (layer2_outputs(2641));
    layer3_outputs(3566) <= '1';
    layer3_outputs(3567) <= not((layer2_outputs(4610)) and (layer2_outputs(2033)));
    layer3_outputs(3568) <= '0';
    layer3_outputs(3569) <= (layer2_outputs(3605)) and (layer2_outputs(1702));
    layer3_outputs(3570) <= (layer2_outputs(3678)) and not (layer2_outputs(4403));
    layer3_outputs(3571) <= not((layer2_outputs(5073)) or (layer2_outputs(2258)));
    layer3_outputs(3572) <= (layer2_outputs(98)) or (layer2_outputs(3794));
    layer3_outputs(3573) <= '1';
    layer3_outputs(3574) <= (layer2_outputs(1033)) or (layer2_outputs(819));
    layer3_outputs(3575) <= not(layer2_outputs(5001));
    layer3_outputs(3576) <= not(layer2_outputs(1246)) or (layer2_outputs(3618));
    layer3_outputs(3577) <= '1';
    layer3_outputs(3578) <= layer2_outputs(1093);
    layer3_outputs(3579) <= '1';
    layer3_outputs(3580) <= not(layer2_outputs(2219));
    layer3_outputs(3581) <= not(layer2_outputs(411));
    layer3_outputs(3582) <= not(layer2_outputs(5060));
    layer3_outputs(3583) <= (layer2_outputs(4779)) or (layer2_outputs(3572));
    layer3_outputs(3584) <= '0';
    layer3_outputs(3585) <= (layer2_outputs(1300)) and not (layer2_outputs(4480));
    layer3_outputs(3586) <= not((layer2_outputs(4872)) and (layer2_outputs(4843)));
    layer3_outputs(3587) <= '0';
    layer3_outputs(3588) <= (layer2_outputs(1022)) or (layer2_outputs(4577));
    layer3_outputs(3589) <= layer2_outputs(2028);
    layer3_outputs(3590) <= '0';
    layer3_outputs(3591) <= (layer2_outputs(3097)) and not (layer2_outputs(4024));
    layer3_outputs(3592) <= (layer2_outputs(4025)) and (layer2_outputs(243));
    layer3_outputs(3593) <= '0';
    layer3_outputs(3594) <= '0';
    layer3_outputs(3595) <= not((layer2_outputs(2922)) or (layer2_outputs(473)));
    layer3_outputs(3596) <= '1';
    layer3_outputs(3597) <= not(layer2_outputs(2740));
    layer3_outputs(3598) <= not((layer2_outputs(2088)) or (layer2_outputs(2555)));
    layer3_outputs(3599) <= '1';
    layer3_outputs(3600) <= (layer2_outputs(2504)) and (layer2_outputs(2109));
    layer3_outputs(3601) <= (layer2_outputs(4268)) and not (layer2_outputs(140));
    layer3_outputs(3602) <= not(layer2_outputs(1179)) or (layer2_outputs(1352));
    layer3_outputs(3603) <= not(layer2_outputs(3862)) or (layer2_outputs(1174));
    layer3_outputs(3604) <= not(layer2_outputs(818)) or (layer2_outputs(2494));
    layer3_outputs(3605) <= '1';
    layer3_outputs(3606) <= '0';
    layer3_outputs(3607) <= (layer2_outputs(1351)) and not (layer2_outputs(946));
    layer3_outputs(3608) <= not((layer2_outputs(4243)) or (layer2_outputs(2400)));
    layer3_outputs(3609) <= layer2_outputs(2586);
    layer3_outputs(3610) <= (layer2_outputs(2332)) and not (layer2_outputs(2349));
    layer3_outputs(3611) <= not((layer2_outputs(3080)) xor (layer2_outputs(2188)));
    layer3_outputs(3612) <= not(layer2_outputs(3725));
    layer3_outputs(3613) <= layer2_outputs(3289);
    layer3_outputs(3614) <= not(layer2_outputs(4946)) or (layer2_outputs(1524));
    layer3_outputs(3615) <= not((layer2_outputs(2075)) and (layer2_outputs(1660)));
    layer3_outputs(3616) <= (layer2_outputs(3507)) xor (layer2_outputs(5069));
    layer3_outputs(3617) <= not(layer2_outputs(1570));
    layer3_outputs(3618) <= '0';
    layer3_outputs(3619) <= layer2_outputs(794);
    layer3_outputs(3620) <= '1';
    layer3_outputs(3621) <= layer2_outputs(2710);
    layer3_outputs(3622) <= (layer2_outputs(3135)) and not (layer2_outputs(642));
    layer3_outputs(3623) <= not(layer2_outputs(2004));
    layer3_outputs(3624) <= '1';
    layer3_outputs(3625) <= '1';
    layer3_outputs(3626) <= (layer2_outputs(2369)) and not (layer2_outputs(538));
    layer3_outputs(3627) <= not(layer2_outputs(1497));
    layer3_outputs(3628) <= not(layer2_outputs(3609)) or (layer2_outputs(1025));
    layer3_outputs(3629) <= (layer2_outputs(4200)) and not (layer2_outputs(4322));
    layer3_outputs(3630) <= not((layer2_outputs(4810)) and (layer2_outputs(3924)));
    layer3_outputs(3631) <= not(layer2_outputs(50)) or (layer2_outputs(672));
    layer3_outputs(3632) <= '1';
    layer3_outputs(3633) <= layer2_outputs(3304);
    layer3_outputs(3634) <= (layer2_outputs(3443)) or (layer2_outputs(2596));
    layer3_outputs(3635) <= (layer2_outputs(3284)) and not (layer2_outputs(4338));
    layer3_outputs(3636) <= (layer2_outputs(2655)) xor (layer2_outputs(4550));
    layer3_outputs(3637) <= layer2_outputs(2517);
    layer3_outputs(3638) <= '0';
    layer3_outputs(3639) <= '0';
    layer3_outputs(3640) <= '0';
    layer3_outputs(3641) <= layer2_outputs(2569);
    layer3_outputs(3642) <= (layer2_outputs(2743)) and not (layer2_outputs(1253));
    layer3_outputs(3643) <= not(layer2_outputs(1798));
    layer3_outputs(3644) <= not((layer2_outputs(711)) or (layer2_outputs(1540)));
    layer3_outputs(3645) <= (layer2_outputs(2962)) and (layer2_outputs(3185));
    layer3_outputs(3646) <= not(layer2_outputs(1890)) or (layer2_outputs(543));
    layer3_outputs(3647) <= '0';
    layer3_outputs(3648) <= not(layer2_outputs(2432)) or (layer2_outputs(3001));
    layer3_outputs(3649) <= layer2_outputs(7);
    layer3_outputs(3650) <= not(layer2_outputs(3155)) or (layer2_outputs(4301));
    layer3_outputs(3651) <= (layer2_outputs(2832)) and (layer2_outputs(883));
    layer3_outputs(3652) <= (layer2_outputs(2446)) or (layer2_outputs(1042));
    layer3_outputs(3653) <= layer2_outputs(1444);
    layer3_outputs(3654) <= not(layer2_outputs(4649)) or (layer2_outputs(2600));
    layer3_outputs(3655) <= not(layer2_outputs(782));
    layer3_outputs(3656) <= (layer2_outputs(1429)) and not (layer2_outputs(965));
    layer3_outputs(3657) <= '1';
    layer3_outputs(3658) <= (layer2_outputs(4910)) and not (layer2_outputs(1303));
    layer3_outputs(3659) <= (layer2_outputs(4521)) or (layer2_outputs(1547));
    layer3_outputs(3660) <= not(layer2_outputs(5093)) or (layer2_outputs(3688));
    layer3_outputs(3661) <= (layer2_outputs(562)) and not (layer2_outputs(514));
    layer3_outputs(3662) <= not((layer2_outputs(3346)) and (layer2_outputs(4118)));
    layer3_outputs(3663) <= (layer2_outputs(1052)) and not (layer2_outputs(716));
    layer3_outputs(3664) <= '0';
    layer3_outputs(3665) <= '0';
    layer3_outputs(3666) <= not(layer2_outputs(2880));
    layer3_outputs(3667) <= not(layer2_outputs(174)) or (layer2_outputs(4971));
    layer3_outputs(3668) <= not((layer2_outputs(3433)) or (layer2_outputs(1225)));
    layer3_outputs(3669) <= '0';
    layer3_outputs(3670) <= '0';
    layer3_outputs(3671) <= layer2_outputs(4500);
    layer3_outputs(3672) <= (layer2_outputs(1090)) and not (layer2_outputs(4661));
    layer3_outputs(3673) <= layer2_outputs(2068);
    layer3_outputs(3674) <= (layer2_outputs(2386)) and (layer2_outputs(4317));
    layer3_outputs(3675) <= layer2_outputs(4983);
    layer3_outputs(3676) <= '1';
    layer3_outputs(3677) <= '1';
    layer3_outputs(3678) <= layer2_outputs(482);
    layer3_outputs(3679) <= layer2_outputs(2536);
    layer3_outputs(3680) <= not(layer2_outputs(621)) or (layer2_outputs(1217));
    layer3_outputs(3681) <= (layer2_outputs(3583)) and (layer2_outputs(987));
    layer3_outputs(3682) <= not(layer2_outputs(1316)) or (layer2_outputs(4896));
    layer3_outputs(3683) <= not((layer2_outputs(193)) or (layer2_outputs(2820)));
    layer3_outputs(3684) <= not((layer2_outputs(3768)) or (layer2_outputs(521)));
    layer3_outputs(3685) <= not(layer2_outputs(751));
    layer3_outputs(3686) <= (layer2_outputs(1358)) and not (layer2_outputs(3347));
    layer3_outputs(3687) <= (layer2_outputs(193)) and not (layer2_outputs(5072));
    layer3_outputs(3688) <= (layer2_outputs(1762)) or (layer2_outputs(1945));
    layer3_outputs(3689) <= '0';
    layer3_outputs(3690) <= not(layer2_outputs(3778));
    layer3_outputs(3691) <= (layer2_outputs(2658)) and not (layer2_outputs(3062));
    layer3_outputs(3692) <= not((layer2_outputs(2299)) and (layer2_outputs(3879)));
    layer3_outputs(3693) <= not(layer2_outputs(3898));
    layer3_outputs(3694) <= (layer2_outputs(2214)) and not (layer2_outputs(2174));
    layer3_outputs(3695) <= not((layer2_outputs(1010)) or (layer2_outputs(939)));
    layer3_outputs(3696) <= layer2_outputs(1556);
    layer3_outputs(3697) <= layer2_outputs(3987);
    layer3_outputs(3698) <= (layer2_outputs(2266)) and not (layer2_outputs(4112));
    layer3_outputs(3699) <= not((layer2_outputs(269)) and (layer2_outputs(72)));
    layer3_outputs(3700) <= not(layer2_outputs(2632));
    layer3_outputs(3701) <= not(layer2_outputs(406)) or (layer2_outputs(1518));
    layer3_outputs(3702) <= (layer2_outputs(3468)) xor (layer2_outputs(22));
    layer3_outputs(3703) <= '0';
    layer3_outputs(3704) <= not((layer2_outputs(4666)) xor (layer2_outputs(4466)));
    layer3_outputs(3705) <= not((layer2_outputs(2377)) and (layer2_outputs(4285)));
    layer3_outputs(3706) <= (layer2_outputs(4497)) xor (layer2_outputs(2831));
    layer3_outputs(3707) <= not(layer2_outputs(4233)) or (layer2_outputs(5115));
    layer3_outputs(3708) <= not((layer2_outputs(607)) and (layer2_outputs(1000)));
    layer3_outputs(3709) <= (layer2_outputs(980)) and (layer2_outputs(1588));
    layer3_outputs(3710) <= not(layer2_outputs(1260));
    layer3_outputs(3711) <= layer2_outputs(4870);
    layer3_outputs(3712) <= not((layer2_outputs(1776)) or (layer2_outputs(3026)));
    layer3_outputs(3713) <= not(layer2_outputs(953));
    layer3_outputs(3714) <= (layer2_outputs(614)) and (layer2_outputs(1901));
    layer3_outputs(3715) <= not(layer2_outputs(4777));
    layer3_outputs(3716) <= not((layer2_outputs(584)) and (layer2_outputs(3966)));
    layer3_outputs(3717) <= '0';
    layer3_outputs(3718) <= '0';
    layer3_outputs(3719) <= not((layer2_outputs(435)) and (layer2_outputs(2070)));
    layer3_outputs(3720) <= '1';
    layer3_outputs(3721) <= (layer2_outputs(4626)) and not (layer2_outputs(964));
    layer3_outputs(3722) <= not(layer2_outputs(4889));
    layer3_outputs(3723) <= not(layer2_outputs(366));
    layer3_outputs(3724) <= '0';
    layer3_outputs(3725) <= not((layer2_outputs(1851)) or (layer2_outputs(3733)));
    layer3_outputs(3726) <= layer2_outputs(175);
    layer3_outputs(3727) <= (layer2_outputs(3795)) or (layer2_outputs(222));
    layer3_outputs(3728) <= (layer2_outputs(208)) xor (layer2_outputs(441));
    layer3_outputs(3729) <= not((layer2_outputs(2112)) xor (layer2_outputs(3137)));
    layer3_outputs(3730) <= (layer2_outputs(3492)) and not (layer2_outputs(1940));
    layer3_outputs(3731) <= not(layer2_outputs(1105)) or (layer2_outputs(3615));
    layer3_outputs(3732) <= not(layer2_outputs(3735)) or (layer2_outputs(4041));
    layer3_outputs(3733) <= (layer2_outputs(4940)) and not (layer2_outputs(2187));
    layer3_outputs(3734) <= (layer2_outputs(3473)) and not (layer2_outputs(2589));
    layer3_outputs(3735) <= (layer2_outputs(410)) and not (layer2_outputs(2253));
    layer3_outputs(3736) <= layer2_outputs(4585);
    layer3_outputs(3737) <= '0';
    layer3_outputs(3738) <= (layer2_outputs(2229)) or (layer2_outputs(3191));
    layer3_outputs(3739) <= '0';
    layer3_outputs(3740) <= (layer2_outputs(1085)) and not (layer2_outputs(1407));
    layer3_outputs(3741) <= not(layer2_outputs(5115)) or (layer2_outputs(4925));
    layer3_outputs(3742) <= not((layer2_outputs(3414)) or (layer2_outputs(4764)));
    layer3_outputs(3743) <= '1';
    layer3_outputs(3744) <= not(layer2_outputs(4168)) or (layer2_outputs(2882));
    layer3_outputs(3745) <= '1';
    layer3_outputs(3746) <= not(layer2_outputs(145)) or (layer2_outputs(1236));
    layer3_outputs(3747) <= not((layer2_outputs(4751)) xor (layer2_outputs(361)));
    layer3_outputs(3748) <= (layer2_outputs(5017)) and not (layer2_outputs(1821));
    layer3_outputs(3749) <= (layer2_outputs(2974)) and not (layer2_outputs(1981));
    layer3_outputs(3750) <= layer2_outputs(2155);
    layer3_outputs(3751) <= not(layer2_outputs(2929));
    layer3_outputs(3752) <= not((layer2_outputs(4060)) and (layer2_outputs(3049)));
    layer3_outputs(3753) <= not((layer2_outputs(4206)) and (layer2_outputs(5099)));
    layer3_outputs(3754) <= not((layer2_outputs(319)) and (layer2_outputs(3247)));
    layer3_outputs(3755) <= layer2_outputs(2914);
    layer3_outputs(3756) <= not(layer2_outputs(4773)) or (layer2_outputs(3297));
    layer3_outputs(3757) <= not(layer2_outputs(4609));
    layer3_outputs(3758) <= not(layer2_outputs(585));
    layer3_outputs(3759) <= not(layer2_outputs(1168)) or (layer2_outputs(940));
    layer3_outputs(3760) <= not((layer2_outputs(4515)) or (layer2_outputs(4128)));
    layer3_outputs(3761) <= '0';
    layer3_outputs(3762) <= layer2_outputs(3478);
    layer3_outputs(3763) <= layer2_outputs(2712);
    layer3_outputs(3764) <= not(layer2_outputs(3652));
    layer3_outputs(3765) <= layer2_outputs(4532);
    layer3_outputs(3766) <= not(layer2_outputs(1829)) or (layer2_outputs(1029));
    layer3_outputs(3767) <= layer2_outputs(466);
    layer3_outputs(3768) <= (layer2_outputs(1736)) and not (layer2_outputs(3165));
    layer3_outputs(3769) <= (layer2_outputs(3887)) and not (layer2_outputs(2458));
    layer3_outputs(3770) <= (layer2_outputs(4698)) and not (layer2_outputs(2141));
    layer3_outputs(3771) <= not(layer2_outputs(5041));
    layer3_outputs(3772) <= layer2_outputs(320);
    layer3_outputs(3773) <= not(layer2_outputs(649)) or (layer2_outputs(712));
    layer3_outputs(3774) <= layer2_outputs(696);
    layer3_outputs(3775) <= layer2_outputs(3845);
    layer3_outputs(3776) <= not(layer2_outputs(182));
    layer3_outputs(3777) <= (layer2_outputs(3123)) and not (layer2_outputs(1477));
    layer3_outputs(3778) <= not(layer2_outputs(1360));
    layer3_outputs(3779) <= not(layer2_outputs(2781)) or (layer2_outputs(1797));
    layer3_outputs(3780) <= '0';
    layer3_outputs(3781) <= '1';
    layer3_outputs(3782) <= not(layer2_outputs(684));
    layer3_outputs(3783) <= (layer2_outputs(4658)) and (layer2_outputs(1855));
    layer3_outputs(3784) <= '0';
    layer3_outputs(3785) <= (layer2_outputs(2078)) and not (layer2_outputs(4080));
    layer3_outputs(3786) <= not((layer2_outputs(4014)) or (layer2_outputs(758)));
    layer3_outputs(3787) <= (layer2_outputs(2612)) or (layer2_outputs(765));
    layer3_outputs(3788) <= (layer2_outputs(791)) and not (layer2_outputs(5012));
    layer3_outputs(3789) <= '0';
    layer3_outputs(3790) <= not(layer2_outputs(4196)) or (layer2_outputs(603));
    layer3_outputs(3791) <= (layer2_outputs(1340)) or (layer2_outputs(979));
    layer3_outputs(3792) <= layer2_outputs(1607);
    layer3_outputs(3793) <= layer2_outputs(2432);
    layer3_outputs(3794) <= not((layer2_outputs(5048)) or (layer2_outputs(848)));
    layer3_outputs(3795) <= (layer2_outputs(5084)) or (layer2_outputs(393));
    layer3_outputs(3796) <= layer2_outputs(5062);
    layer3_outputs(3797) <= not(layer2_outputs(216));
    layer3_outputs(3798) <= (layer2_outputs(3035)) or (layer2_outputs(3392));
    layer3_outputs(3799) <= (layer2_outputs(537)) and (layer2_outputs(2174));
    layer3_outputs(3800) <= not((layer2_outputs(4112)) or (layer2_outputs(3265)));
    layer3_outputs(3801) <= layer2_outputs(3410);
    layer3_outputs(3802) <= (layer2_outputs(130)) and not (layer2_outputs(2859));
    layer3_outputs(3803) <= '1';
    layer3_outputs(3804) <= not(layer2_outputs(4397));
    layer3_outputs(3805) <= (layer2_outputs(2288)) and (layer2_outputs(2594));
    layer3_outputs(3806) <= not(layer2_outputs(3463)) or (layer2_outputs(1432));
    layer3_outputs(3807) <= not(layer2_outputs(4767)) or (layer2_outputs(1352));
    layer3_outputs(3808) <= '0';
    layer3_outputs(3809) <= not(layer2_outputs(699));
    layer3_outputs(3810) <= '0';
    layer3_outputs(3811) <= '1';
    layer3_outputs(3812) <= (layer2_outputs(4323)) and (layer2_outputs(1991));
    layer3_outputs(3813) <= not(layer2_outputs(1683));
    layer3_outputs(3814) <= not(layer2_outputs(4696));
    layer3_outputs(3815) <= layer2_outputs(712);
    layer3_outputs(3816) <= layer2_outputs(4931);
    layer3_outputs(3817) <= (layer2_outputs(86)) or (layer2_outputs(5070));
    layer3_outputs(3818) <= not(layer2_outputs(4476));
    layer3_outputs(3819) <= not(layer2_outputs(2465)) or (layer2_outputs(2737));
    layer3_outputs(3820) <= layer2_outputs(3196);
    layer3_outputs(3821) <= not((layer2_outputs(419)) and (layer2_outputs(2279)));
    layer3_outputs(3822) <= not((layer2_outputs(4572)) and (layer2_outputs(424)));
    layer3_outputs(3823) <= (layer2_outputs(4297)) and (layer2_outputs(55));
    layer3_outputs(3824) <= not(layer2_outputs(3006));
    layer3_outputs(3825) <= not(layer2_outputs(2472)) or (layer2_outputs(3637));
    layer3_outputs(3826) <= (layer2_outputs(3077)) and not (layer2_outputs(459));
    layer3_outputs(3827) <= '1';
    layer3_outputs(3828) <= layer2_outputs(1459);
    layer3_outputs(3829) <= layer2_outputs(2471);
    layer3_outputs(3830) <= not((layer2_outputs(4359)) or (layer2_outputs(1370)));
    layer3_outputs(3831) <= not(layer2_outputs(3104)) or (layer2_outputs(4666));
    layer3_outputs(3832) <= '0';
    layer3_outputs(3833) <= not(layer2_outputs(4505)) or (layer2_outputs(833));
    layer3_outputs(3834) <= (layer2_outputs(957)) and not (layer2_outputs(1339));
    layer3_outputs(3835) <= (layer2_outputs(4064)) and (layer2_outputs(4862));
    layer3_outputs(3836) <= layer2_outputs(1387);
    layer3_outputs(3837) <= (layer2_outputs(2496)) or (layer2_outputs(4715));
    layer3_outputs(3838) <= (layer2_outputs(726)) and (layer2_outputs(101));
    layer3_outputs(3839) <= not((layer2_outputs(3848)) or (layer2_outputs(845)));
    layer3_outputs(3840) <= (layer2_outputs(516)) and (layer2_outputs(4125));
    layer3_outputs(3841) <= (layer2_outputs(579)) and (layer2_outputs(3883));
    layer3_outputs(3842) <= not(layer2_outputs(4981)) or (layer2_outputs(4503));
    layer3_outputs(3843) <= layer2_outputs(2675);
    layer3_outputs(3844) <= (layer2_outputs(4602)) and not (layer2_outputs(4374));
    layer3_outputs(3845) <= not(layer2_outputs(697)) or (layer2_outputs(1461));
    layer3_outputs(3846) <= '0';
    layer3_outputs(3847) <= not((layer2_outputs(2562)) or (layer2_outputs(4957)));
    layer3_outputs(3848) <= '0';
    layer3_outputs(3849) <= '1';
    layer3_outputs(3850) <= not(layer2_outputs(1843)) or (layer2_outputs(4772));
    layer3_outputs(3851) <= '1';
    layer3_outputs(3852) <= (layer2_outputs(1669)) or (layer2_outputs(3555));
    layer3_outputs(3853) <= not(layer2_outputs(2217)) or (layer2_outputs(3732));
    layer3_outputs(3854) <= '1';
    layer3_outputs(3855) <= (layer2_outputs(4780)) and (layer2_outputs(1959));
    layer3_outputs(3856) <= not((layer2_outputs(421)) and (layer2_outputs(39)));
    layer3_outputs(3857) <= (layer2_outputs(1345)) or (layer2_outputs(2346));
    layer3_outputs(3858) <= not(layer2_outputs(2716));
    layer3_outputs(3859) <= layer2_outputs(766);
    layer3_outputs(3860) <= not(layer2_outputs(3601)) or (layer2_outputs(2404));
    layer3_outputs(3861) <= not(layer2_outputs(2549));
    layer3_outputs(3862) <= not(layer2_outputs(2431));
    layer3_outputs(3863) <= '0';
    layer3_outputs(3864) <= layer2_outputs(566);
    layer3_outputs(3865) <= (layer2_outputs(3714)) and not (layer2_outputs(3357));
    layer3_outputs(3866) <= (layer2_outputs(1641)) or (layer2_outputs(3717));
    layer3_outputs(3867) <= layer2_outputs(659);
    layer3_outputs(3868) <= (layer2_outputs(968)) and not (layer2_outputs(4918));
    layer3_outputs(3869) <= not(layer2_outputs(1357));
    layer3_outputs(3870) <= layer2_outputs(3945);
    layer3_outputs(3871) <= not(layer2_outputs(1543)) or (layer2_outputs(2410));
    layer3_outputs(3872) <= '0';
    layer3_outputs(3873) <= (layer2_outputs(2313)) and (layer2_outputs(5047));
    layer3_outputs(3874) <= '0';
    layer3_outputs(3875) <= layer2_outputs(4753);
    layer3_outputs(3876) <= not(layer2_outputs(2366));
    layer3_outputs(3877) <= layer2_outputs(4378);
    layer3_outputs(3878) <= '0';
    layer3_outputs(3879) <= not(layer2_outputs(2962)) or (layer2_outputs(1002));
    layer3_outputs(3880) <= layer2_outputs(5013);
    layer3_outputs(3881) <= '0';
    layer3_outputs(3882) <= (layer2_outputs(3065)) or (layer2_outputs(138));
    layer3_outputs(3883) <= (layer2_outputs(4202)) and (layer2_outputs(4178));
    layer3_outputs(3884) <= '0';
    layer3_outputs(3885) <= '1';
    layer3_outputs(3886) <= (layer2_outputs(3741)) and not (layer2_outputs(4084));
    layer3_outputs(3887) <= layer2_outputs(2125);
    layer3_outputs(3888) <= '1';
    layer3_outputs(3889) <= '1';
    layer3_outputs(3890) <= layer2_outputs(3230);
    layer3_outputs(3891) <= '1';
    layer3_outputs(3892) <= not(layer2_outputs(5030)) or (layer2_outputs(381));
    layer3_outputs(3893) <= not((layer2_outputs(1276)) or (layer2_outputs(3288)));
    layer3_outputs(3894) <= '1';
    layer3_outputs(3895) <= not(layer2_outputs(655));
    layer3_outputs(3896) <= '0';
    layer3_outputs(3897) <= layer2_outputs(4427);
    layer3_outputs(3898) <= (layer2_outputs(1120)) and not (layer2_outputs(455));
    layer3_outputs(3899) <= (layer2_outputs(917)) and not (layer2_outputs(3372));
    layer3_outputs(3900) <= (layer2_outputs(515)) and not (layer2_outputs(222));
    layer3_outputs(3901) <= (layer2_outputs(1279)) or (layer2_outputs(325));
    layer3_outputs(3902) <= not(layer2_outputs(1672));
    layer3_outputs(3903) <= not(layer2_outputs(2831));
    layer3_outputs(3904) <= layer2_outputs(3372);
    layer3_outputs(3905) <= '1';
    layer3_outputs(3906) <= '1';
    layer3_outputs(3907) <= layer2_outputs(3358);
    layer3_outputs(3908) <= not(layer2_outputs(4115)) or (layer2_outputs(5110));
    layer3_outputs(3909) <= not(layer2_outputs(1189));
    layer3_outputs(3910) <= layer2_outputs(326);
    layer3_outputs(3911) <= not(layer2_outputs(3947)) or (layer2_outputs(1462));
    layer3_outputs(3912) <= not(layer2_outputs(125));
    layer3_outputs(3913) <= not(layer2_outputs(792));
    layer3_outputs(3914) <= not((layer2_outputs(3384)) and (layer2_outputs(3455)));
    layer3_outputs(3915) <= not((layer2_outputs(400)) and (layer2_outputs(2492)));
    layer3_outputs(3916) <= '0';
    layer3_outputs(3917) <= not(layer2_outputs(2597)) or (layer2_outputs(3417));
    layer3_outputs(3918) <= (layer2_outputs(161)) and not (layer2_outputs(1689));
    layer3_outputs(3919) <= layer2_outputs(2227);
    layer3_outputs(3920) <= not(layer2_outputs(919)) or (layer2_outputs(701));
    layer3_outputs(3921) <= not(layer2_outputs(236)) or (layer2_outputs(2386));
    layer3_outputs(3922) <= not(layer2_outputs(3188));
    layer3_outputs(3923) <= (layer2_outputs(2156)) and not (layer2_outputs(2265));
    layer3_outputs(3924) <= (layer2_outputs(1642)) and (layer2_outputs(3702));
    layer3_outputs(3925) <= layer2_outputs(1139);
    layer3_outputs(3926) <= '1';
    layer3_outputs(3927) <= (layer2_outputs(2430)) or (layer2_outputs(61));
    layer3_outputs(3928) <= layer2_outputs(1076);
    layer3_outputs(3929) <= not((layer2_outputs(2934)) or (layer2_outputs(71)));
    layer3_outputs(3930) <= '0';
    layer3_outputs(3931) <= not(layer2_outputs(3375));
    layer3_outputs(3932) <= not(layer2_outputs(2157)) or (layer2_outputs(2524));
    layer3_outputs(3933) <= not((layer2_outputs(2190)) and (layer2_outputs(929)));
    layer3_outputs(3934) <= not(layer2_outputs(2833)) or (layer2_outputs(569));
    layer3_outputs(3935) <= '1';
    layer3_outputs(3936) <= not(layer2_outputs(4024));
    layer3_outputs(3937) <= not(layer2_outputs(4209)) or (layer2_outputs(3169));
    layer3_outputs(3938) <= '0';
    layer3_outputs(3939) <= '0';
    layer3_outputs(3940) <= (layer2_outputs(733)) and (layer2_outputs(1698));
    layer3_outputs(3941) <= '1';
    layer3_outputs(3942) <= not(layer2_outputs(3259));
    layer3_outputs(3943) <= '0';
    layer3_outputs(3944) <= not(layer2_outputs(4798));
    layer3_outputs(3945) <= (layer2_outputs(2981)) and not (layer2_outputs(5116));
    layer3_outputs(3946) <= not(layer2_outputs(1362));
    layer3_outputs(3947) <= '1';
    layer3_outputs(3948) <= '0';
    layer3_outputs(3949) <= (layer2_outputs(1807)) and (layer2_outputs(4080));
    layer3_outputs(3950) <= layer2_outputs(3528);
    layer3_outputs(3951) <= '0';
    layer3_outputs(3952) <= '0';
    layer3_outputs(3953) <= not(layer2_outputs(2071)) or (layer2_outputs(3242));
    layer3_outputs(3954) <= not((layer2_outputs(1347)) or (layer2_outputs(986)));
    layer3_outputs(3955) <= layer2_outputs(3179);
    layer3_outputs(3956) <= not((layer2_outputs(887)) or (layer2_outputs(1258)));
    layer3_outputs(3957) <= (layer2_outputs(3606)) or (layer2_outputs(4676));
    layer3_outputs(3958) <= layer2_outputs(3752);
    layer3_outputs(3959) <= (layer2_outputs(1132)) and not (layer2_outputs(407));
    layer3_outputs(3960) <= not(layer2_outputs(4888));
    layer3_outputs(3961) <= '1';
    layer3_outputs(3962) <= not((layer2_outputs(343)) and (layer2_outputs(3804)));
    layer3_outputs(3963) <= (layer2_outputs(2095)) and not (layer2_outputs(2456));
    layer3_outputs(3964) <= layer2_outputs(2896);
    layer3_outputs(3965) <= '1';
    layer3_outputs(3966) <= not(layer2_outputs(5015)) or (layer2_outputs(3438));
    layer3_outputs(3967) <= (layer2_outputs(4869)) and not (layer2_outputs(4310));
    layer3_outputs(3968) <= (layer2_outputs(627)) or (layer2_outputs(5116));
    layer3_outputs(3969) <= layer2_outputs(949);
    layer3_outputs(3970) <= not((layer2_outputs(1450)) or (layer2_outputs(1147)));
    layer3_outputs(3971) <= layer2_outputs(2711);
    layer3_outputs(3972) <= '0';
    layer3_outputs(3973) <= (layer2_outputs(4580)) and (layer2_outputs(1222));
    layer3_outputs(3974) <= '0';
    layer3_outputs(3975) <= (layer2_outputs(1763)) and not (layer2_outputs(2649));
    layer3_outputs(3976) <= layer2_outputs(4814);
    layer3_outputs(3977) <= (layer2_outputs(4746)) and not (layer2_outputs(5034));
    layer3_outputs(3978) <= (layer2_outputs(4930)) and not (layer2_outputs(4265));
    layer3_outputs(3979) <= '0';
    layer3_outputs(3980) <= layer2_outputs(1294);
    layer3_outputs(3981) <= not(layer2_outputs(2802));
    layer3_outputs(3982) <= '0';
    layer3_outputs(3983) <= (layer2_outputs(3922)) or (layer2_outputs(212));
    layer3_outputs(3984) <= (layer2_outputs(3256)) and not (layer2_outputs(2736));
    layer3_outputs(3985) <= '1';
    layer3_outputs(3986) <= '1';
    layer3_outputs(3987) <= not(layer2_outputs(4577)) or (layer2_outputs(1071));
    layer3_outputs(3988) <= not(layer2_outputs(2697));
    layer3_outputs(3989) <= not(layer2_outputs(4251)) or (layer2_outputs(1869));
    layer3_outputs(3990) <= not((layer2_outputs(2278)) and (layer2_outputs(4634)));
    layer3_outputs(3991) <= not(layer2_outputs(4907)) or (layer2_outputs(4127));
    layer3_outputs(3992) <= layer2_outputs(290);
    layer3_outputs(3993) <= not((layer2_outputs(3930)) and (layer2_outputs(2913)));
    layer3_outputs(3994) <= not(layer2_outputs(194)) or (layer2_outputs(534));
    layer3_outputs(3995) <= not(layer2_outputs(2789));
    layer3_outputs(3996) <= (layer2_outputs(4011)) and not (layer2_outputs(2618));
    layer3_outputs(3997) <= (layer2_outputs(2412)) and (layer2_outputs(434));
    layer3_outputs(3998) <= layer2_outputs(4565);
    layer3_outputs(3999) <= '0';
    layer3_outputs(4000) <= layer2_outputs(3319);
    layer3_outputs(4001) <= (layer2_outputs(2648)) and not (layer2_outputs(2856));
    layer3_outputs(4002) <= layer2_outputs(1543);
    layer3_outputs(4003) <= (layer2_outputs(5080)) and not (layer2_outputs(3020));
    layer3_outputs(4004) <= '1';
    layer3_outputs(4005) <= not((layer2_outputs(1211)) and (layer2_outputs(3673)));
    layer3_outputs(4006) <= not(layer2_outputs(3173));
    layer3_outputs(4007) <= layer2_outputs(2871);
    layer3_outputs(4008) <= layer2_outputs(807);
    layer3_outputs(4009) <= (layer2_outputs(3367)) or (layer2_outputs(4616));
    layer3_outputs(4010) <= layer2_outputs(1734);
    layer3_outputs(4011) <= not(layer2_outputs(667)) or (layer2_outputs(3586));
    layer3_outputs(4012) <= layer2_outputs(3318);
    layer3_outputs(4013) <= not(layer2_outputs(1205)) or (layer2_outputs(1188));
    layer3_outputs(4014) <= not(layer2_outputs(436));
    layer3_outputs(4015) <= not(layer2_outputs(1739));
    layer3_outputs(4016) <= '1';
    layer3_outputs(4017) <= (layer2_outputs(907)) and (layer2_outputs(403));
    layer3_outputs(4018) <= not(layer2_outputs(4488)) or (layer2_outputs(4661));
    layer3_outputs(4019) <= '1';
    layer3_outputs(4020) <= layer2_outputs(1017);
    layer3_outputs(4021) <= not((layer2_outputs(254)) and (layer2_outputs(94)));
    layer3_outputs(4022) <= '1';
    layer3_outputs(4023) <= (layer2_outputs(2811)) or (layer2_outputs(4472));
    layer3_outputs(4024) <= layer2_outputs(682);
    layer3_outputs(4025) <= not(layer2_outputs(4685)) or (layer2_outputs(2841));
    layer3_outputs(4026) <= layer2_outputs(4109);
    layer3_outputs(4027) <= (layer2_outputs(708)) xor (layer2_outputs(3141));
    layer3_outputs(4028) <= (layer2_outputs(1553)) and not (layer2_outputs(752));
    layer3_outputs(4029) <= '1';
    layer3_outputs(4030) <= '0';
    layer3_outputs(4031) <= '0';
    layer3_outputs(4032) <= not(layer2_outputs(1601));
    layer3_outputs(4033) <= '0';
    layer3_outputs(4034) <= layer2_outputs(2593);
    layer3_outputs(4035) <= (layer2_outputs(1304)) and not (layer2_outputs(1903));
    layer3_outputs(4036) <= not((layer2_outputs(134)) or (layer2_outputs(4558)));
    layer3_outputs(4037) <= (layer2_outputs(1108)) or (layer2_outputs(3674));
    layer3_outputs(4038) <= (layer2_outputs(3196)) and (layer2_outputs(1418));
    layer3_outputs(4039) <= layer2_outputs(1753);
    layer3_outputs(4040) <= (layer2_outputs(1049)) and not (layer2_outputs(4308));
    layer3_outputs(4041) <= not(layer2_outputs(3448)) or (layer2_outputs(1165));
    layer3_outputs(4042) <= '1';
    layer3_outputs(4043) <= (layer2_outputs(1216)) or (layer2_outputs(2790));
    layer3_outputs(4044) <= not((layer2_outputs(1922)) or (layer2_outputs(2688)));
    layer3_outputs(4045) <= (layer2_outputs(855)) or (layer2_outputs(2930));
    layer3_outputs(4046) <= (layer2_outputs(3381)) or (layer2_outputs(1714));
    layer3_outputs(4047) <= (layer2_outputs(4217)) and not (layer2_outputs(2297));
    layer3_outputs(4048) <= (layer2_outputs(968)) and (layer2_outputs(2500));
    layer3_outputs(4049) <= (layer2_outputs(2917)) and not (layer2_outputs(2733));
    layer3_outputs(4050) <= (layer2_outputs(1986)) and (layer2_outputs(180));
    layer3_outputs(4051) <= not((layer2_outputs(2452)) and (layer2_outputs(1331)));
    layer3_outputs(4052) <= not(layer2_outputs(5014));
    layer3_outputs(4053) <= (layer2_outputs(2537)) and not (layer2_outputs(2027));
    layer3_outputs(4054) <= not(layer2_outputs(2923));
    layer3_outputs(4055) <= (layer2_outputs(148)) or (layer2_outputs(560));
    layer3_outputs(4056) <= '0';
    layer3_outputs(4057) <= '0';
    layer3_outputs(4058) <= not((layer2_outputs(1620)) or (layer2_outputs(4872)));
    layer3_outputs(4059) <= (layer2_outputs(1886)) and not (layer2_outputs(2481));
    layer3_outputs(4060) <= not((layer2_outputs(765)) and (layer2_outputs(4341)));
    layer3_outputs(4061) <= layer2_outputs(3521);
    layer3_outputs(4062) <= '1';
    layer3_outputs(4063) <= (layer2_outputs(3588)) and not (layer2_outputs(3208));
    layer3_outputs(4064) <= '1';
    layer3_outputs(4065) <= (layer2_outputs(1408)) and not (layer2_outputs(4186));
    layer3_outputs(4066) <= not(layer2_outputs(4871));
    layer3_outputs(4067) <= not(layer2_outputs(4270));
    layer3_outputs(4068) <= not(layer2_outputs(1230)) or (layer2_outputs(4388));
    layer3_outputs(4069) <= (layer2_outputs(2230)) xor (layer2_outputs(1558));
    layer3_outputs(4070) <= (layer2_outputs(4419)) or (layer2_outputs(1658));
    layer3_outputs(4071) <= '0';
    layer3_outputs(4072) <= (layer2_outputs(2214)) and (layer2_outputs(5085));
    layer3_outputs(4073) <= (layer2_outputs(136)) and (layer2_outputs(3963));
    layer3_outputs(4074) <= '1';
    layer3_outputs(4075) <= not(layer2_outputs(3594)) or (layer2_outputs(3351));
    layer3_outputs(4076) <= not((layer2_outputs(3905)) or (layer2_outputs(5111)));
    layer3_outputs(4077) <= not(layer2_outputs(2773)) or (layer2_outputs(4592));
    layer3_outputs(4078) <= (layer2_outputs(3800)) and not (layer2_outputs(3337));
    layer3_outputs(4079) <= layer2_outputs(799);
    layer3_outputs(4080) <= not(layer2_outputs(658));
    layer3_outputs(4081) <= (layer2_outputs(4272)) and (layer2_outputs(1816));
    layer3_outputs(4082) <= layer2_outputs(1513);
    layer3_outputs(4083) <= layer2_outputs(946);
    layer3_outputs(4084) <= not(layer2_outputs(44)) or (layer2_outputs(3311));
    layer3_outputs(4085) <= not(layer2_outputs(1763)) or (layer2_outputs(4041));
    layer3_outputs(4086) <= (layer2_outputs(4614)) and not (layer2_outputs(3965));
    layer3_outputs(4087) <= not(layer2_outputs(3859)) or (layer2_outputs(3956));
    layer3_outputs(4088) <= (layer2_outputs(94)) and not (layer2_outputs(4781));
    layer3_outputs(4089) <= layer2_outputs(245);
    layer3_outputs(4090) <= (layer2_outputs(3201)) and not (layer2_outputs(3970));
    layer3_outputs(4091) <= (layer2_outputs(4431)) and not (layer2_outputs(3220));
    layer3_outputs(4092) <= layer2_outputs(1138);
    layer3_outputs(4093) <= layer2_outputs(2525);
    layer3_outputs(4094) <= layer2_outputs(1334);
    layer3_outputs(4095) <= (layer2_outputs(3589)) and not (layer2_outputs(1129));
    layer3_outputs(4096) <= not((layer2_outputs(457)) and (layer2_outputs(3272)));
    layer3_outputs(4097) <= not(layer2_outputs(2200));
    layer3_outputs(4098) <= '1';
    layer3_outputs(4099) <= (layer2_outputs(2867)) xor (layer2_outputs(1133));
    layer3_outputs(4100) <= '0';
    layer3_outputs(4101) <= not((layer2_outputs(4890)) and (layer2_outputs(1226)));
    layer3_outputs(4102) <= (layer2_outputs(4339)) and not (layer2_outputs(3280));
    layer3_outputs(4103) <= not(layer2_outputs(3471));
    layer3_outputs(4104) <= (layer2_outputs(4331)) and (layer2_outputs(1819));
    layer3_outputs(4105) <= layer2_outputs(1952);
    layer3_outputs(4106) <= '1';
    layer3_outputs(4107) <= '1';
    layer3_outputs(4108) <= not((layer2_outputs(3023)) and (layer2_outputs(1682)));
    layer3_outputs(4109) <= not(layer2_outputs(4339));
    layer3_outputs(4110) <= layer2_outputs(2723);
    layer3_outputs(4111) <= (layer2_outputs(4083)) and (layer2_outputs(283));
    layer3_outputs(4112) <= layer2_outputs(1998);
    layer3_outputs(4113) <= layer2_outputs(187);
    layer3_outputs(4114) <= not((layer2_outputs(2641)) or (layer2_outputs(2125)));
    layer3_outputs(4115) <= (layer2_outputs(3327)) and not (layer2_outputs(928));
    layer3_outputs(4116) <= not((layer2_outputs(2540)) or (layer2_outputs(1189)));
    layer3_outputs(4117) <= '0';
    layer3_outputs(4118) <= '1';
    layer3_outputs(4119) <= (layer2_outputs(839)) xor (layer2_outputs(489));
    layer3_outputs(4120) <= '1';
    layer3_outputs(4121) <= not(layer2_outputs(1949)) or (layer2_outputs(2107));
    layer3_outputs(4122) <= '1';
    layer3_outputs(4123) <= '1';
    layer3_outputs(4124) <= '0';
    layer3_outputs(4125) <= layer2_outputs(4854);
    layer3_outputs(4126) <= '0';
    layer3_outputs(4127) <= not(layer2_outputs(4426)) or (layer2_outputs(316));
    layer3_outputs(4128) <= not((layer2_outputs(1087)) and (layer2_outputs(873)));
    layer3_outputs(4129) <= not((layer2_outputs(1624)) xor (layer2_outputs(3277)));
    layer3_outputs(4130) <= (layer2_outputs(2762)) and not (layer2_outputs(1174));
    layer3_outputs(4131) <= not(layer2_outputs(4820)) or (layer2_outputs(2514));
    layer3_outputs(4132) <= '1';
    layer3_outputs(4133) <= not((layer2_outputs(2148)) xor (layer2_outputs(2024)));
    layer3_outputs(4134) <= layer2_outputs(1416);
    layer3_outputs(4135) <= '1';
    layer3_outputs(4136) <= not((layer2_outputs(332)) or (layer2_outputs(4432)));
    layer3_outputs(4137) <= (layer2_outputs(1705)) or (layer2_outputs(4369));
    layer3_outputs(4138) <= '1';
    layer3_outputs(4139) <= not((layer2_outputs(1952)) xor (layer2_outputs(73)));
    layer3_outputs(4140) <= (layer2_outputs(253)) or (layer2_outputs(2402));
    layer3_outputs(4141) <= not((layer2_outputs(3108)) or (layer2_outputs(4589)));
    layer3_outputs(4142) <= '1';
    layer3_outputs(4143) <= '1';
    layer3_outputs(4144) <= not(layer2_outputs(876)) or (layer2_outputs(4265));
    layer3_outputs(4145) <= '1';
    layer3_outputs(4146) <= (layer2_outputs(1377)) or (layer2_outputs(1750));
    layer3_outputs(4147) <= (layer2_outputs(2658)) and not (layer2_outputs(3766));
    layer3_outputs(4148) <= layer2_outputs(894);
    layer3_outputs(4149) <= (layer2_outputs(1148)) and (layer2_outputs(4315));
    layer3_outputs(4150) <= not(layer2_outputs(898)) or (layer2_outputs(1731));
    layer3_outputs(4151) <= not(layer2_outputs(162)) or (layer2_outputs(3026));
    layer3_outputs(4152) <= not((layer2_outputs(3556)) xor (layer2_outputs(5004)));
    layer3_outputs(4153) <= not(layer2_outputs(3677));
    layer3_outputs(4154) <= not(layer2_outputs(2103));
    layer3_outputs(4155) <= (layer2_outputs(558)) or (layer2_outputs(4509));
    layer3_outputs(4156) <= layer2_outputs(258);
    layer3_outputs(4157) <= (layer2_outputs(3557)) xor (layer2_outputs(1204));
    layer3_outputs(4158) <= (layer2_outputs(3453)) xor (layer2_outputs(4650));
    layer3_outputs(4159) <= (layer2_outputs(4740)) and (layer2_outputs(1934));
    layer3_outputs(4160) <= not(layer2_outputs(391));
    layer3_outputs(4161) <= not(layer2_outputs(2523));
    layer3_outputs(4162) <= (layer2_outputs(313)) and not (layer2_outputs(2073));
    layer3_outputs(4163) <= not(layer2_outputs(992));
    layer3_outputs(4164) <= not(layer2_outputs(3264));
    layer3_outputs(4165) <= '0';
    layer3_outputs(4166) <= '0';
    layer3_outputs(4167) <= (layer2_outputs(1742)) and not (layer2_outputs(748));
    layer3_outputs(4168) <= not(layer2_outputs(1934));
    layer3_outputs(4169) <= layer2_outputs(4294);
    layer3_outputs(4170) <= not(layer2_outputs(4538));
    layer3_outputs(4171) <= not(layer2_outputs(2642));
    layer3_outputs(4172) <= '1';
    layer3_outputs(4173) <= layer2_outputs(4282);
    layer3_outputs(4174) <= (layer2_outputs(2329)) or (layer2_outputs(3202));
    layer3_outputs(4175) <= not(layer2_outputs(4935)) or (layer2_outputs(1751));
    layer3_outputs(4176) <= not((layer2_outputs(1875)) or (layer2_outputs(711)));
    layer3_outputs(4177) <= (layer2_outputs(1599)) and not (layer2_outputs(158));
    layer3_outputs(4178) <= layer2_outputs(4373);
    layer3_outputs(4179) <= not((layer2_outputs(97)) and (layer2_outputs(2273)));
    layer3_outputs(4180) <= not((layer2_outputs(4309)) and (layer2_outputs(3720)));
    layer3_outputs(4181) <= (layer2_outputs(4757)) and (layer2_outputs(2394));
    layer3_outputs(4182) <= (layer2_outputs(680)) and not (layer2_outputs(2474));
    layer3_outputs(4183) <= (layer2_outputs(831)) and not (layer2_outputs(427));
    layer3_outputs(4184) <= not(layer2_outputs(1643));
    layer3_outputs(4185) <= '0';
    layer3_outputs(4186) <= '1';
    layer3_outputs(4187) <= (layer2_outputs(4043)) and (layer2_outputs(1175));
    layer3_outputs(4188) <= (layer2_outputs(683)) or (layer2_outputs(2331));
    layer3_outputs(4189) <= (layer2_outputs(3214)) and not (layer2_outputs(1757));
    layer3_outputs(4190) <= not(layer2_outputs(1185));
    layer3_outputs(4191) <= not(layer2_outputs(403));
    layer3_outputs(4192) <= (layer2_outputs(4139)) or (layer2_outputs(4342));
    layer3_outputs(4193) <= (layer2_outputs(2618)) xor (layer2_outputs(2092));
    layer3_outputs(4194) <= (layer2_outputs(2744)) and (layer2_outputs(2719));
    layer3_outputs(4195) <= layer2_outputs(3639);
    layer3_outputs(4196) <= '0';
    layer3_outputs(4197) <= '1';
    layer3_outputs(4198) <= not(layer2_outputs(3213)) or (layer2_outputs(4774));
    layer3_outputs(4199) <= not(layer2_outputs(5052)) or (layer2_outputs(268));
    layer3_outputs(4200) <= not(layer2_outputs(69));
    layer3_outputs(4201) <= not(layer2_outputs(4662)) or (layer2_outputs(4647));
    layer3_outputs(4202) <= (layer2_outputs(1565)) and not (layer2_outputs(5050));
    layer3_outputs(4203) <= '1';
    layer3_outputs(4204) <= not((layer2_outputs(231)) and (layer2_outputs(1849)));
    layer3_outputs(4205) <= (layer2_outputs(1318)) and not (layer2_outputs(1364));
    layer3_outputs(4206) <= not(layer2_outputs(1135)) or (layer2_outputs(2120));
    layer3_outputs(4207) <= '1';
    layer3_outputs(4208) <= (layer2_outputs(4402)) and not (layer2_outputs(1194));
    layer3_outputs(4209) <= layer2_outputs(4979);
    layer3_outputs(4210) <= not(layer2_outputs(353)) or (layer2_outputs(1130));
    layer3_outputs(4211) <= '0';
    layer3_outputs(4212) <= layer2_outputs(4392);
    layer3_outputs(4213) <= not(layer2_outputs(4516));
    layer3_outputs(4214) <= layer2_outputs(806);
    layer3_outputs(4215) <= not(layer2_outputs(4451));
    layer3_outputs(4216) <= (layer2_outputs(3159)) and not (layer2_outputs(1294));
    layer3_outputs(4217) <= not((layer2_outputs(4579)) and (layer2_outputs(4019)));
    layer3_outputs(4218) <= (layer2_outputs(842)) and not (layer2_outputs(3032));
    layer3_outputs(4219) <= not(layer2_outputs(3932));
    layer3_outputs(4220) <= (layer2_outputs(2140)) and not (layer2_outputs(1127));
    layer3_outputs(4221) <= not(layer2_outputs(2762));
    layer3_outputs(4222) <= layer2_outputs(4826);
    layer3_outputs(4223) <= not(layer2_outputs(4484)) or (layer2_outputs(3694));
    layer3_outputs(4224) <= (layer2_outputs(2436)) and not (layer2_outputs(1445));
    layer3_outputs(4225) <= not(layer2_outputs(3454));
    layer3_outputs(4226) <= layer2_outputs(4073);
    layer3_outputs(4227) <= not(layer2_outputs(543)) or (layer2_outputs(826));
    layer3_outputs(4228) <= '1';
    layer3_outputs(4229) <= not((layer2_outputs(3964)) and (layer2_outputs(992)));
    layer3_outputs(4230) <= layer2_outputs(1774);
    layer3_outputs(4231) <= '0';
    layer3_outputs(4232) <= not(layer2_outputs(2334));
    layer3_outputs(4233) <= not(layer2_outputs(2422));
    layer3_outputs(4234) <= '0';
    layer3_outputs(4235) <= (layer2_outputs(4856)) or (layer2_outputs(3912));
    layer3_outputs(4236) <= not(layer2_outputs(2621));
    layer3_outputs(4237) <= layer2_outputs(1980);
    layer3_outputs(4238) <= '0';
    layer3_outputs(4239) <= not(layer2_outputs(3260)) or (layer2_outputs(3678));
    layer3_outputs(4240) <= '1';
    layer3_outputs(4241) <= (layer2_outputs(4349)) and (layer2_outputs(3650));
    layer3_outputs(4242) <= (layer2_outputs(2842)) and (layer2_outputs(1758));
    layer3_outputs(4243) <= '0';
    layer3_outputs(4244) <= layer2_outputs(1711);
    layer3_outputs(4245) <= layer2_outputs(4865);
    layer3_outputs(4246) <= not((layer2_outputs(4813)) and (layer2_outputs(2352)));
    layer3_outputs(4247) <= not(layer2_outputs(1533)) or (layer2_outputs(408));
    layer3_outputs(4248) <= not((layer2_outputs(4960)) and (layer2_outputs(3781)));
    layer3_outputs(4249) <= not(layer2_outputs(837)) or (layer2_outputs(1377));
    layer3_outputs(4250) <= '0';
    layer3_outputs(4251) <= (layer2_outputs(2320)) or (layer2_outputs(3412));
    layer3_outputs(4252) <= not(layer2_outputs(581)) or (layer2_outputs(1565));
    layer3_outputs(4253) <= (layer2_outputs(4400)) and not (layer2_outputs(4636));
    layer3_outputs(4254) <= (layer2_outputs(678)) or (layer2_outputs(1167));
    layer3_outputs(4255) <= layer2_outputs(446);
    layer3_outputs(4256) <= '0';
    layer3_outputs(4257) <= '0';
    layer3_outputs(4258) <= not(layer2_outputs(5057)) or (layer2_outputs(2518));
    layer3_outputs(4259) <= '1';
    layer3_outputs(4260) <= (layer2_outputs(3211)) and not (layer2_outputs(1156));
    layer3_outputs(4261) <= layer2_outputs(4903);
    layer3_outputs(4262) <= not(layer2_outputs(952)) or (layer2_outputs(1780));
    layer3_outputs(4263) <= not(layer2_outputs(3124)) or (layer2_outputs(4815));
    layer3_outputs(4264) <= not((layer2_outputs(3944)) xor (layer2_outputs(1018)));
    layer3_outputs(4265) <= (layer2_outputs(2862)) and (layer2_outputs(2242));
    layer3_outputs(4266) <= (layer2_outputs(4799)) and not (layer2_outputs(4621));
    layer3_outputs(4267) <= not(layer2_outputs(1788));
    layer3_outputs(4268) <= '1';
    layer3_outputs(4269) <= (layer2_outputs(892)) and not (layer2_outputs(1408));
    layer3_outputs(4270) <= not(layer2_outputs(1944));
    layer3_outputs(4271) <= not(layer2_outputs(690));
    layer3_outputs(4272) <= '1';
    layer3_outputs(4273) <= not(layer2_outputs(4414)) or (layer2_outputs(2097));
    layer3_outputs(4274) <= (layer2_outputs(5077)) and (layer2_outputs(282));
    layer3_outputs(4275) <= '1';
    layer3_outputs(4276) <= (layer2_outputs(4832)) and not (layer2_outputs(1379));
    layer3_outputs(4277) <= (layer2_outputs(1166)) and not (layer2_outputs(3551));
    layer3_outputs(4278) <= layer2_outputs(3890);
    layer3_outputs(4279) <= not((layer2_outputs(2403)) and (layer2_outputs(4564)));
    layer3_outputs(4280) <= layer2_outputs(796);
    layer3_outputs(4281) <= not(layer2_outputs(3410)) or (layer2_outputs(4926));
    layer3_outputs(4282) <= (layer2_outputs(1645)) xor (layer2_outputs(4182));
    layer3_outputs(4283) <= '1';
    layer3_outputs(4284) <= (layer2_outputs(5063)) and (layer2_outputs(3164));
    layer3_outputs(4285) <= layer2_outputs(1908);
    layer3_outputs(4286) <= not((layer2_outputs(1251)) or (layer2_outputs(3779)));
    layer3_outputs(4287) <= layer2_outputs(2702);
    layer3_outputs(4288) <= not(layer2_outputs(636));
    layer3_outputs(4289) <= not(layer2_outputs(1106)) or (layer2_outputs(3728));
    layer3_outputs(4290) <= not(layer2_outputs(1411));
    layer3_outputs(4291) <= (layer2_outputs(764)) and (layer2_outputs(180));
    layer3_outputs(4292) <= '1';
    layer3_outputs(4293) <= '1';
    layer3_outputs(4294) <= not(layer2_outputs(78));
    layer3_outputs(4295) <= (layer2_outputs(4693)) and (layer2_outputs(2329));
    layer3_outputs(4296) <= (layer2_outputs(3643)) xor (layer2_outputs(1870));
    layer3_outputs(4297) <= not((layer2_outputs(4370)) and (layer2_outputs(58)));
    layer3_outputs(4298) <= (layer2_outputs(717)) and not (layer2_outputs(1566));
    layer3_outputs(4299) <= not((layer2_outputs(3009)) and (layer2_outputs(4705)));
    layer3_outputs(4300) <= not(layer2_outputs(1368));
    layer3_outputs(4301) <= not((layer2_outputs(1570)) or (layer2_outputs(4252)));
    layer3_outputs(4302) <= (layer2_outputs(2617)) and not (layer2_outputs(556));
    layer3_outputs(4303) <= '1';
    layer3_outputs(4304) <= layer2_outputs(3323);
    layer3_outputs(4305) <= (layer2_outputs(863)) and (layer2_outputs(4825));
    layer3_outputs(4306) <= (layer2_outputs(2700)) or (layer2_outputs(4146));
    layer3_outputs(4307) <= '0';
    layer3_outputs(4308) <= '0';
    layer3_outputs(4309) <= not(layer2_outputs(2746));
    layer3_outputs(4310) <= not((layer2_outputs(3826)) or (layer2_outputs(3613)));
    layer3_outputs(4311) <= '1';
    layer3_outputs(4312) <= layer2_outputs(38);
    layer3_outputs(4313) <= (layer2_outputs(1319)) and (layer2_outputs(2378));
    layer3_outputs(4314) <= '1';
    layer3_outputs(4315) <= (layer2_outputs(2967)) and not (layer2_outputs(1964));
    layer3_outputs(4316) <= not(layer2_outputs(2259)) or (layer2_outputs(2157));
    layer3_outputs(4317) <= layer2_outputs(3860);
    layer3_outputs(4318) <= (layer2_outputs(4913)) and not (layer2_outputs(1475));
    layer3_outputs(4319) <= (layer2_outputs(5092)) and (layer2_outputs(2566));
    layer3_outputs(4320) <= layer2_outputs(4814);
    layer3_outputs(4321) <= (layer2_outputs(2463)) and (layer2_outputs(4889));
    layer3_outputs(4322) <= '0';
    layer3_outputs(4323) <= (layer2_outputs(728)) or (layer2_outputs(1557));
    layer3_outputs(4324) <= (layer2_outputs(573)) and not (layer2_outputs(967));
    layer3_outputs(4325) <= '0';
    layer3_outputs(4326) <= '1';
    layer3_outputs(4327) <= (layer2_outputs(117)) or (layer2_outputs(1677));
    layer3_outputs(4328) <= (layer2_outputs(3851)) and (layer2_outputs(4215));
    layer3_outputs(4329) <= layer2_outputs(4540);
    layer3_outputs(4330) <= not(layer2_outputs(2464)) or (layer2_outputs(727));
    layer3_outputs(4331) <= not(layer2_outputs(1680));
    layer3_outputs(4332) <= (layer2_outputs(2041)) and not (layer2_outputs(2119));
    layer3_outputs(4333) <= not(layer2_outputs(2231));
    layer3_outputs(4334) <= (layer2_outputs(1437)) and (layer2_outputs(1859));
    layer3_outputs(4335) <= (layer2_outputs(4376)) and not (layer2_outputs(371));
    layer3_outputs(4336) <= not(layer2_outputs(3164)) or (layer2_outputs(2617));
    layer3_outputs(4337) <= (layer2_outputs(962)) and (layer2_outputs(2690));
    layer3_outputs(4338) <= '1';
    layer3_outputs(4339) <= not(layer2_outputs(4178));
    layer3_outputs(4340) <= not(layer2_outputs(45));
    layer3_outputs(4341) <= layer2_outputs(294);
    layer3_outputs(4342) <= not(layer2_outputs(1428)) or (layer2_outputs(1206));
    layer3_outputs(4343) <= '0';
    layer3_outputs(4344) <= '0';
    layer3_outputs(4345) <= (layer2_outputs(1052)) and (layer2_outputs(3439));
    layer3_outputs(4346) <= not(layer2_outputs(950));
    layer3_outputs(4347) <= (layer2_outputs(4236)) or (layer2_outputs(478));
    layer3_outputs(4348) <= (layer2_outputs(2864)) and not (layer2_outputs(4989));
    layer3_outputs(4349) <= not((layer2_outputs(3811)) and (layer2_outputs(1681)));
    layer3_outputs(4350) <= (layer2_outputs(1001)) or (layer2_outputs(650));
    layer3_outputs(4351) <= (layer2_outputs(3233)) and not (layer2_outputs(3036));
    layer3_outputs(4352) <= not((layer2_outputs(4894)) xor (layer2_outputs(2341)));
    layer3_outputs(4353) <= (layer2_outputs(1061)) and not (layer2_outputs(43));
    layer3_outputs(4354) <= (layer2_outputs(2499)) and (layer2_outputs(4048));
    layer3_outputs(4355) <= not((layer2_outputs(847)) and (layer2_outputs(2045)));
    layer3_outputs(4356) <= not(layer2_outputs(178)) or (layer2_outputs(1320));
    layer3_outputs(4357) <= '1';
    layer3_outputs(4358) <= (layer2_outputs(1757)) or (layer2_outputs(2928));
    layer3_outputs(4359) <= (layer2_outputs(1972)) and not (layer2_outputs(4662));
    layer3_outputs(4360) <= not(layer2_outputs(3439)) or (layer2_outputs(3497));
    layer3_outputs(4361) <= not((layer2_outputs(3446)) and (layer2_outputs(3704)));
    layer3_outputs(4362) <= not((layer2_outputs(4677)) xor (layer2_outputs(432)));
    layer3_outputs(4363) <= not((layer2_outputs(833)) or (layer2_outputs(1676)));
    layer3_outputs(4364) <= not(layer2_outputs(3038)) or (layer2_outputs(1631));
    layer3_outputs(4365) <= not(layer2_outputs(122)) or (layer2_outputs(4751));
    layer3_outputs(4366) <= not(layer2_outputs(2338));
    layer3_outputs(4367) <= not((layer2_outputs(3557)) and (layer2_outputs(3213)));
    layer3_outputs(4368) <= (layer2_outputs(2176)) and not (layer2_outputs(753));
    layer3_outputs(4369) <= (layer2_outputs(1053)) and not (layer2_outputs(3760));
    layer3_outputs(4370) <= '0';
    layer3_outputs(4371) <= '0';
    layer3_outputs(4372) <= not(layer2_outputs(24));
    layer3_outputs(4373) <= '0';
    layer3_outputs(4374) <= (layer2_outputs(1447)) and (layer2_outputs(4627));
    layer3_outputs(4375) <= '1';
    layer3_outputs(4376) <= not(layer2_outputs(3914));
    layer3_outputs(4377) <= '0';
    layer3_outputs(4378) <= not(layer2_outputs(574)) or (layer2_outputs(662));
    layer3_outputs(4379) <= layer2_outputs(2287);
    layer3_outputs(4380) <= '0';
    layer3_outputs(4381) <= not((layer2_outputs(839)) or (layer2_outputs(3181)));
    layer3_outputs(4382) <= (layer2_outputs(995)) and not (layer2_outputs(4600));
    layer3_outputs(4383) <= layer2_outputs(2819);
    layer3_outputs(4384) <= not(layer2_outputs(3154));
    layer3_outputs(4385) <= '1';
    layer3_outputs(4386) <= not(layer2_outputs(2461));
    layer3_outputs(4387) <= '1';
    layer3_outputs(4388) <= layer2_outputs(3764);
    layer3_outputs(4389) <= (layer2_outputs(2652)) xor (layer2_outputs(3095));
    layer3_outputs(4390) <= '0';
    layer3_outputs(4391) <= '1';
    layer3_outputs(4392) <= not((layer2_outputs(2534)) or (layer2_outputs(3753)));
    layer3_outputs(4393) <= (layer2_outputs(395)) and not (layer2_outputs(2506));
    layer3_outputs(4394) <= (layer2_outputs(2627)) or (layer2_outputs(2684));
    layer3_outputs(4395) <= not(layer2_outputs(2367));
    layer3_outputs(4396) <= not((layer2_outputs(4428)) or (layer2_outputs(2981)));
    layer3_outputs(4397) <= (layer2_outputs(3386)) and not (layer2_outputs(4987));
    layer3_outputs(4398) <= (layer2_outputs(2513)) and not (layer2_outputs(1095));
    layer3_outputs(4399) <= layer2_outputs(796);
    layer3_outputs(4400) <= not((layer2_outputs(1348)) xor (layer2_outputs(3774)));
    layer3_outputs(4401) <= (layer2_outputs(2715)) and (layer2_outputs(4210));
    layer3_outputs(4402) <= (layer2_outputs(3219)) or (layer2_outputs(4977));
    layer3_outputs(4403) <= not(layer2_outputs(4846)) or (layer2_outputs(3718));
    layer3_outputs(4404) <= '0';
    layer3_outputs(4405) <= (layer2_outputs(1883)) and (layer2_outputs(2619));
    layer3_outputs(4406) <= not(layer2_outputs(3192)) or (layer2_outputs(3711));
    layer3_outputs(4407) <= (layer2_outputs(4251)) and not (layer2_outputs(1601));
    layer3_outputs(4408) <= (layer2_outputs(2909)) or (layer2_outputs(1112));
    layer3_outputs(4409) <= not(layer2_outputs(2207));
    layer3_outputs(4410) <= not((layer2_outputs(2376)) and (layer2_outputs(651)));
    layer3_outputs(4411) <= not(layer2_outputs(3088));
    layer3_outputs(4412) <= not((layer2_outputs(1576)) or (layer2_outputs(4987)));
    layer3_outputs(4413) <= not((layer2_outputs(4247)) and (layer2_outputs(2876)));
    layer3_outputs(4414) <= layer2_outputs(2429);
    layer3_outputs(4415) <= (layer2_outputs(2767)) and (layer2_outputs(3764));
    layer3_outputs(4416) <= '0';
    layer3_outputs(4417) <= not((layer2_outputs(3828)) and (layer2_outputs(4094)));
    layer3_outputs(4418) <= '1';
    layer3_outputs(4419) <= (layer2_outputs(920)) or (layer2_outputs(4954));
    layer3_outputs(4420) <= not(layer2_outputs(3515)) or (layer2_outputs(3610));
    layer3_outputs(4421) <= (layer2_outputs(922)) and (layer2_outputs(1631));
    layer3_outputs(4422) <= (layer2_outputs(2704)) and (layer2_outputs(2489));
    layer3_outputs(4423) <= not(layer2_outputs(4091)) or (layer2_outputs(3841));
    layer3_outputs(4424) <= (layer2_outputs(1604)) or (layer2_outputs(2108));
    layer3_outputs(4425) <= not((layer2_outputs(1373)) and (layer2_outputs(825)));
    layer3_outputs(4426) <= layer2_outputs(4070);
    layer3_outputs(4427) <= layer2_outputs(4686);
    layer3_outputs(4428) <= not(layer2_outputs(1322));
    layer3_outputs(4429) <= not(layer2_outputs(417)) or (layer2_outputs(1609));
    layer3_outputs(4430) <= not(layer2_outputs(4716));
    layer3_outputs(4431) <= (layer2_outputs(5022)) or (layer2_outputs(5098));
    layer3_outputs(4432) <= not(layer2_outputs(1708));
    layer3_outputs(4433) <= (layer2_outputs(2311)) and not (layer2_outputs(3904));
    layer3_outputs(4434) <= not(layer2_outputs(1212)) or (layer2_outputs(1987));
    layer3_outputs(4435) <= (layer2_outputs(2577)) and not (layer2_outputs(710));
    layer3_outputs(4436) <= not(layer2_outputs(4438)) or (layer2_outputs(1546));
    layer3_outputs(4437) <= not(layer2_outputs(4069));
    layer3_outputs(4438) <= (layer2_outputs(1035)) xor (layer2_outputs(2166));
    layer3_outputs(4439) <= not(layer2_outputs(2030)) or (layer2_outputs(2973));
    layer3_outputs(4440) <= '0';
    layer3_outputs(4441) <= not(layer2_outputs(260));
    layer3_outputs(4442) <= not(layer2_outputs(3069)) or (layer2_outputs(1814));
    layer3_outputs(4443) <= '1';
    layer3_outputs(4444) <= (layer2_outputs(2285)) and (layer2_outputs(2772));
    layer3_outputs(4445) <= (layer2_outputs(2414)) and not (layer2_outputs(437));
    layer3_outputs(4446) <= not(layer2_outputs(4449)) or (layer2_outputs(3075));
    layer3_outputs(4447) <= layer2_outputs(4425);
    layer3_outputs(4448) <= (layer2_outputs(1116)) and not (layer2_outputs(965));
    layer3_outputs(4449) <= not(layer2_outputs(3655));
    layer3_outputs(4450) <= '0';
    layer3_outputs(4451) <= '1';
    layer3_outputs(4452) <= not(layer2_outputs(1754)) or (layer2_outputs(4892));
    layer3_outputs(4453) <= not(layer2_outputs(5023)) or (layer2_outputs(2249));
    layer3_outputs(4454) <= not((layer2_outputs(2038)) or (layer2_outputs(2457)));
    layer3_outputs(4455) <= '0';
    layer3_outputs(4456) <= not(layer2_outputs(723));
    layer3_outputs(4457) <= (layer2_outputs(3447)) or (layer2_outputs(2822));
    layer3_outputs(4458) <= '1';
    layer3_outputs(4459) <= (layer2_outputs(1963)) and not (layer2_outputs(2240));
    layer3_outputs(4460) <= (layer2_outputs(4575)) and (layer2_outputs(663));
    layer3_outputs(4461) <= (layer2_outputs(322)) xor (layer2_outputs(1997));
    layer3_outputs(4462) <= not(layer2_outputs(1482)) or (layer2_outputs(195));
    layer3_outputs(4463) <= not((layer2_outputs(930)) and (layer2_outputs(2140)));
    layer3_outputs(4464) <= (layer2_outputs(4346)) and not (layer2_outputs(1100));
    layer3_outputs(4465) <= '1';
    layer3_outputs(4466) <= not((layer2_outputs(4072)) or (layer2_outputs(4821)));
    layer3_outputs(4467) <= not(layer2_outputs(157)) or (layer2_outputs(270));
    layer3_outputs(4468) <= not((layer2_outputs(4201)) or (layer2_outputs(1976)));
    layer3_outputs(4469) <= '1';
    layer3_outputs(4470) <= not((layer2_outputs(70)) and (layer2_outputs(4108)));
    layer3_outputs(4471) <= layer2_outputs(2123);
    layer3_outputs(4472) <= not(layer2_outputs(5083)) or (layer2_outputs(4529));
    layer3_outputs(4473) <= (layer2_outputs(4861)) and (layer2_outputs(2453));
    layer3_outputs(4474) <= '0';
    layer3_outputs(4475) <= not(layer2_outputs(2961));
    layer3_outputs(4476) <= (layer2_outputs(4527)) and not (layer2_outputs(444));
    layer3_outputs(4477) <= '1';
    layer3_outputs(4478) <= (layer2_outputs(497)) or (layer2_outputs(3402));
    layer3_outputs(4479) <= (layer2_outputs(198)) and (layer2_outputs(1512));
    layer3_outputs(4480) <= (layer2_outputs(4627)) and not (layer2_outputs(1461));
    layer3_outputs(4481) <= (layer2_outputs(3161)) and (layer2_outputs(4760));
    layer3_outputs(4482) <= not(layer2_outputs(3130)) or (layer2_outputs(1823));
    layer3_outputs(4483) <= not(layer2_outputs(4130));
    layer3_outputs(4484) <= (layer2_outputs(1983)) and not (layer2_outputs(3415));
    layer3_outputs(4485) <= not(layer2_outputs(834));
    layer3_outputs(4486) <= '0';
    layer3_outputs(4487) <= not(layer2_outputs(3475)) or (layer2_outputs(804));
    layer3_outputs(4488) <= not(layer2_outputs(3903)) or (layer2_outputs(2571));
    layer3_outputs(4489) <= not((layer2_outputs(852)) and (layer2_outputs(667)));
    layer3_outputs(4490) <= not(layer2_outputs(3030));
    layer3_outputs(4491) <= not(layer2_outputs(1034));
    layer3_outputs(4492) <= not((layer2_outputs(1876)) and (layer2_outputs(2527)));
    layer3_outputs(4493) <= '0';
    layer3_outputs(4494) <= not((layer2_outputs(4455)) or (layer2_outputs(2274)));
    layer3_outputs(4495) <= not(layer2_outputs(4673)) or (layer2_outputs(830));
    layer3_outputs(4496) <= not(layer2_outputs(1007));
    layer3_outputs(4497) <= layer2_outputs(3261);
    layer3_outputs(4498) <= '0';
    layer3_outputs(4499) <= '1';
    layer3_outputs(4500) <= (layer2_outputs(4735)) or (layer2_outputs(170));
    layer3_outputs(4501) <= '0';
    layer3_outputs(4502) <= layer2_outputs(2053);
    layer3_outputs(4503) <= '1';
    layer3_outputs(4504) <= not(layer2_outputs(3058));
    layer3_outputs(4505) <= not(layer2_outputs(2264)) or (layer2_outputs(2872));
    layer3_outputs(4506) <= '1';
    layer3_outputs(4507) <= not(layer2_outputs(3886)) or (layer2_outputs(3257));
    layer3_outputs(4508) <= '1';
    layer3_outputs(4509) <= (layer2_outputs(1196)) and not (layer2_outputs(2276));
    layer3_outputs(4510) <= not((layer2_outputs(1722)) and (layer2_outputs(3960)));
    layer3_outputs(4511) <= (layer2_outputs(3949)) or (layer2_outputs(664));
    layer3_outputs(4512) <= (layer2_outputs(3503)) and not (layer2_outputs(2936));
    layer3_outputs(4513) <= not((layer2_outputs(351)) and (layer2_outputs(2118)));
    layer3_outputs(4514) <= not(layer2_outputs(2529));
    layer3_outputs(4515) <= layer2_outputs(3347);
    layer3_outputs(4516) <= not(layer2_outputs(691)) or (layer2_outputs(617));
    layer3_outputs(4517) <= not(layer2_outputs(695));
    layer3_outputs(4518) <= not((layer2_outputs(4638)) or (layer2_outputs(4367)));
    layer3_outputs(4519) <= (layer2_outputs(4179)) and not (layer2_outputs(4183));
    layer3_outputs(4520) <= not((layer2_outputs(2380)) or (layer2_outputs(114)));
    layer3_outputs(4521) <= (layer2_outputs(719)) xor (layer2_outputs(1655));
    layer3_outputs(4522) <= '0';
    layer3_outputs(4523) <= '1';
    layer3_outputs(4524) <= not((layer2_outputs(4360)) or (layer2_outputs(944)));
    layer3_outputs(4525) <= '0';
    layer3_outputs(4526) <= not(layer2_outputs(1805));
    layer3_outputs(4527) <= not((layer2_outputs(3573)) or (layer2_outputs(4594)));
    layer3_outputs(4528) <= (layer2_outputs(3246)) and (layer2_outputs(4679));
    layer3_outputs(4529) <= '0';
    layer3_outputs(4530) <= (layer2_outputs(4089)) and not (layer2_outputs(3704));
    layer3_outputs(4531) <= not(layer2_outputs(4291)) or (layer2_outputs(3324));
    layer3_outputs(4532) <= (layer2_outputs(3745)) or (layer2_outputs(3500));
    layer3_outputs(4533) <= not(layer2_outputs(2467));
    layer3_outputs(4534) <= '0';
    layer3_outputs(4535) <= (layer2_outputs(1434)) and (layer2_outputs(2735));
    layer3_outputs(4536) <= (layer2_outputs(4199)) or (layer2_outputs(4345));
    layer3_outputs(4537) <= (layer2_outputs(3100)) or (layer2_outputs(512));
    layer3_outputs(4538) <= layer2_outputs(4738);
    layer3_outputs(4539) <= not(layer2_outputs(2330));
    layer3_outputs(4540) <= layer2_outputs(1637);
    layer3_outputs(4541) <= (layer2_outputs(3280)) or (layer2_outputs(1242));
    layer3_outputs(4542) <= not((layer2_outputs(4437)) or (layer2_outputs(3961)));
    layer3_outputs(4543) <= (layer2_outputs(880)) and not (layer2_outputs(2665));
    layer3_outputs(4544) <= not(layer2_outputs(3281));
    layer3_outputs(4545) <= not(layer2_outputs(3399)) or (layer2_outputs(3491));
    layer3_outputs(4546) <= not(layer2_outputs(4068)) or (layer2_outputs(4350));
    layer3_outputs(4547) <= '0';
    layer3_outputs(4548) <= not(layer2_outputs(2211)) or (layer2_outputs(1884));
    layer3_outputs(4549) <= layer2_outputs(1356);
    layer3_outputs(4550) <= not((layer2_outputs(1247)) and (layer2_outputs(2104)));
    layer3_outputs(4551) <= not(layer2_outputs(1853)) or (layer2_outputs(4361));
    layer3_outputs(4552) <= not((layer2_outputs(1404)) or (layer2_outputs(4526)));
    layer3_outputs(4553) <= '0';
    layer3_outputs(4554) <= (layer2_outputs(201)) and not (layer2_outputs(1690));
    layer3_outputs(4555) <= not(layer2_outputs(1555)) or (layer2_outputs(4874));
    layer3_outputs(4556) <= '0';
    layer3_outputs(4557) <= layer2_outputs(324);
    layer3_outputs(4558) <= not((layer2_outputs(1959)) and (layer2_outputs(1200)));
    layer3_outputs(4559) <= not(layer2_outputs(2445));
    layer3_outputs(4560) <= layer2_outputs(458);
    layer3_outputs(4561) <= layer2_outputs(3712);
    layer3_outputs(4562) <= not(layer2_outputs(318));
    layer3_outputs(4563) <= '1';
    layer3_outputs(4564) <= not(layer2_outputs(2480));
    layer3_outputs(4565) <= layer2_outputs(3323);
    layer3_outputs(4566) <= '1';
    layer3_outputs(4567) <= not((layer2_outputs(3063)) or (layer2_outputs(2007)));
    layer3_outputs(4568) <= not((layer2_outputs(633)) and (layer2_outputs(1151)));
    layer3_outputs(4569) <= layer2_outputs(2799);
    layer3_outputs(4570) <= '0';
    layer3_outputs(4571) <= (layer2_outputs(744)) and not (layer2_outputs(2579));
    layer3_outputs(4572) <= '0';
    layer3_outputs(4573) <= layer2_outputs(4274);
    layer3_outputs(4574) <= not((layer2_outputs(5039)) or (layer2_outputs(4642)));
    layer3_outputs(4575) <= layer2_outputs(2309);
    layer3_outputs(4576) <= '0';
    layer3_outputs(4577) <= '0';
    layer3_outputs(4578) <= (layer2_outputs(198)) and (layer2_outputs(413));
    layer3_outputs(4579) <= layer2_outputs(5020);
    layer3_outputs(4580) <= (layer2_outputs(1044)) and not (layer2_outputs(1309));
    layer3_outputs(4581) <= not(layer2_outputs(4392));
    layer3_outputs(4582) <= '0';
    layer3_outputs(4583) <= (layer2_outputs(1258)) and not (layer2_outputs(4672));
    layer3_outputs(4584) <= layer2_outputs(904);
    layer3_outputs(4585) <= '0';
    layer3_outputs(4586) <= (layer2_outputs(687)) or (layer2_outputs(2884));
    layer3_outputs(4587) <= (layer2_outputs(2048)) and (layer2_outputs(3604));
    layer3_outputs(4588) <= layer2_outputs(1544);
    layer3_outputs(4589) <= (layer2_outputs(1541)) and not (layer2_outputs(4996));
    layer3_outputs(4590) <= (layer2_outputs(4393)) and (layer2_outputs(3455));
    layer3_outputs(4591) <= (layer2_outputs(4327)) and not (layer2_outputs(4829));
    layer3_outputs(4592) <= not((layer2_outputs(240)) and (layer2_outputs(2822)));
    layer3_outputs(4593) <= '0';
    layer3_outputs(4594) <= not((layer2_outputs(301)) or (layer2_outputs(2925)));
    layer3_outputs(4595) <= (layer2_outputs(107)) and (layer2_outputs(151));
    layer3_outputs(4596) <= not(layer2_outputs(2344)) or (layer2_outputs(1782));
    layer3_outputs(4597) <= (layer2_outputs(1917)) or (layer2_outputs(4129));
    layer3_outputs(4598) <= (layer2_outputs(1012)) xor (layer2_outputs(3394));
    layer3_outputs(4599) <= '0';
    layer3_outputs(4600) <= '0';
    layer3_outputs(4601) <= (layer2_outputs(1510)) or (layer2_outputs(822));
    layer3_outputs(4602) <= (layer2_outputs(5090)) and not (layer2_outputs(2899));
    layer3_outputs(4603) <= not((layer2_outputs(4475)) and (layer2_outputs(545)));
    layer3_outputs(4604) <= layer2_outputs(632);
    layer3_outputs(4605) <= layer2_outputs(3593);
    layer3_outputs(4606) <= '0';
    layer3_outputs(4607) <= (layer2_outputs(1466)) and not (layer2_outputs(3265));
    layer3_outputs(4608) <= (layer2_outputs(2361)) and not (layer2_outputs(939));
    layer3_outputs(4609) <= not((layer2_outputs(1555)) and (layer2_outputs(3945)));
    layer3_outputs(4610) <= not((layer2_outputs(3260)) and (layer2_outputs(4057)));
    layer3_outputs(4611) <= (layer2_outputs(2025)) or (layer2_outputs(984));
    layer3_outputs(4612) <= not(layer2_outputs(3957)) or (layer2_outputs(4644));
    layer3_outputs(4613) <= not(layer2_outputs(3175)) or (layer2_outputs(1566));
    layer3_outputs(4614) <= layer2_outputs(4970);
    layer3_outputs(4615) <= '0';
    layer3_outputs(4616) <= (layer2_outputs(3064)) xor (layer2_outputs(4605));
    layer3_outputs(4617) <= layer2_outputs(4714);
    layer3_outputs(4618) <= not(layer2_outputs(3562));
    layer3_outputs(4619) <= not(layer2_outputs(1026)) or (layer2_outputs(4188));
    layer3_outputs(4620) <= not(layer2_outputs(3887)) or (layer2_outputs(1084));
    layer3_outputs(4621) <= '1';
    layer3_outputs(4622) <= '0';
    layer3_outputs(4623) <= layer2_outputs(3524);
    layer3_outputs(4624) <= not(layer2_outputs(3971));
    layer3_outputs(4625) <= (layer2_outputs(4608)) and not (layer2_outputs(4603));
    layer3_outputs(4626) <= not(layer2_outputs(2825));
    layer3_outputs(4627) <= (layer2_outputs(4902)) or (layer2_outputs(5033));
    layer3_outputs(4628) <= (layer2_outputs(1650)) and (layer2_outputs(2590));
    layer3_outputs(4629) <= layer2_outputs(1666);
    layer3_outputs(4630) <= '1';
    layer3_outputs(4631) <= (layer2_outputs(4689)) and not (layer2_outputs(1608));
    layer3_outputs(4632) <= not(layer2_outputs(1054)) or (layer2_outputs(2039));
    layer3_outputs(4633) <= layer2_outputs(3909);
    layer3_outputs(4634) <= not(layer2_outputs(2364)) or (layer2_outputs(1130));
    layer3_outputs(4635) <= (layer2_outputs(3646)) and not (layer2_outputs(2959));
    layer3_outputs(4636) <= (layer2_outputs(3769)) and not (layer2_outputs(3825));
    layer3_outputs(4637) <= layer2_outputs(34);
    layer3_outputs(4638) <= not(layer2_outputs(1390)) or (layer2_outputs(1323));
    layer3_outputs(4639) <= not((layer2_outputs(2896)) or (layer2_outputs(3309)));
    layer3_outputs(4640) <= not(layer2_outputs(3758)) or (layer2_outputs(928));
    layer3_outputs(4641) <= not(layer2_outputs(2374)) or (layer2_outputs(4972));
    layer3_outputs(4642) <= (layer2_outputs(2732)) and (layer2_outputs(853));
    layer3_outputs(4643) <= not(layer2_outputs(4371)) or (layer2_outputs(2853));
    layer3_outputs(4644) <= '1';
    layer3_outputs(4645) <= (layer2_outputs(1857)) or (layer2_outputs(3834));
    layer3_outputs(4646) <= not(layer2_outputs(1280)) or (layer2_outputs(1590));
    layer3_outputs(4647) <= '1';
    layer3_outputs(4648) <= (layer2_outputs(428)) or (layer2_outputs(643));
    layer3_outputs(4649) <= (layer2_outputs(2270)) and (layer2_outputs(4439));
    layer3_outputs(4650) <= not((layer2_outputs(2054)) and (layer2_outputs(2784)));
    layer3_outputs(4651) <= '0';
    layer3_outputs(4652) <= (layer2_outputs(2796)) and not (layer2_outputs(153));
    layer3_outputs(4653) <= '0';
    layer3_outputs(4654) <= (layer2_outputs(2989)) or (layer2_outputs(2786));
    layer3_outputs(4655) <= layer2_outputs(4103);
    layer3_outputs(4656) <= '0';
    layer3_outputs(4657) <= layer2_outputs(4847);
    layer3_outputs(4658) <= '1';
    layer3_outputs(4659) <= not(layer2_outputs(1664)) or (layer2_outputs(3614));
    layer3_outputs(4660) <= (layer2_outputs(311)) and not (layer2_outputs(4656));
    layer3_outputs(4661) <= '1';
    layer3_outputs(4662) <= not((layer2_outputs(5049)) xor (layer2_outputs(748)));
    layer3_outputs(4663) <= (layer2_outputs(1927)) or (layer2_outputs(2072));
    layer3_outputs(4664) <= not(layer2_outputs(2630)) or (layer2_outputs(3028));
    layer3_outputs(4665) <= not((layer2_outputs(1905)) or (layer2_outputs(750)));
    layer3_outputs(4666) <= not(layer2_outputs(951)) or (layer2_outputs(2777));
    layer3_outputs(4667) <= (layer2_outputs(2917)) or (layer2_outputs(3270));
    layer3_outputs(4668) <= (layer2_outputs(4734)) or (layer2_outputs(2700));
    layer3_outputs(4669) <= (layer2_outputs(1310)) and not (layer2_outputs(3340));
    layer3_outputs(4670) <= not((layer2_outputs(4166)) xor (layer2_outputs(4576)));
    layer3_outputs(4671) <= (layer2_outputs(4079)) and (layer2_outputs(108));
    layer3_outputs(4672) <= (layer2_outputs(3359)) and (layer2_outputs(1106));
    layer3_outputs(4673) <= (layer2_outputs(630)) or (layer2_outputs(1957));
    layer3_outputs(4674) <= (layer2_outputs(1375)) and not (layer2_outputs(2848));
    layer3_outputs(4675) <= (layer2_outputs(675)) xor (layer2_outputs(1886));
    layer3_outputs(4676) <= layer2_outputs(3801);
    layer3_outputs(4677) <= (layer2_outputs(3614)) or (layer2_outputs(5070));
    layer3_outputs(4678) <= (layer2_outputs(2973)) and not (layer2_outputs(2362));
    layer3_outputs(4679) <= '1';
    layer3_outputs(4680) <= layer2_outputs(4276);
    layer3_outputs(4681) <= not(layer2_outputs(2371)) or (layer2_outputs(4744));
    layer3_outputs(4682) <= '0';
    layer3_outputs(4683) <= (layer2_outputs(3606)) or (layer2_outputs(1479));
    layer3_outputs(4684) <= not(layer2_outputs(2523));
    layer3_outputs(4685) <= not(layer2_outputs(1122));
    layer3_outputs(4686) <= not(layer2_outputs(2026)) or (layer2_outputs(2424));
    layer3_outputs(4687) <= not((layer2_outputs(3462)) and (layer2_outputs(1474)));
    layer3_outputs(4688) <= not(layer2_outputs(3400));
    layer3_outputs(4689) <= (layer2_outputs(2096)) and not (layer2_outputs(1750));
    layer3_outputs(4690) <= not(layer2_outputs(2008)) or (layer2_outputs(1930));
    layer3_outputs(4691) <= (layer2_outputs(2466)) and (layer2_outputs(5064));
    layer3_outputs(4692) <= not(layer2_outputs(1436));
    layer3_outputs(4693) <= '0';
    layer3_outputs(4694) <= (layer2_outputs(3515)) and not (layer2_outputs(2860));
    layer3_outputs(4695) <= not(layer2_outputs(472));
    layer3_outputs(4696) <= '0';
    layer3_outputs(4697) <= layer2_outputs(1305);
    layer3_outputs(4698) <= not(layer2_outputs(498));
    layer3_outputs(4699) <= (layer2_outputs(2321)) and not (layer2_outputs(3946));
    layer3_outputs(4700) <= (layer2_outputs(1623)) and (layer2_outputs(3537));
    layer3_outputs(4701) <= not(layer2_outputs(3918));
    layer3_outputs(4702) <= (layer2_outputs(1267)) and not (layer2_outputs(3798));
    layer3_outputs(4703) <= (layer2_outputs(1354)) or (layer2_outputs(3910));
    layer3_outputs(4704) <= not(layer2_outputs(1587));
    layer3_outputs(4705) <= not(layer2_outputs(4389)) or (layer2_outputs(296));
    layer3_outputs(4706) <= '1';
    layer3_outputs(4707) <= (layer2_outputs(159)) and not (layer2_outputs(3896));
    layer3_outputs(4708) <= not(layer2_outputs(861)) or (layer2_outputs(5074));
    layer3_outputs(4709) <= not(layer2_outputs(3348));
    layer3_outputs(4710) <= (layer2_outputs(2751)) or (layer2_outputs(1019));
    layer3_outputs(4711) <= (layer2_outputs(1263)) and not (layer2_outputs(5114));
    layer3_outputs(4712) <= '0';
    layer3_outputs(4713) <= (layer2_outputs(4639)) and not (layer2_outputs(3763));
    layer3_outputs(4714) <= layer2_outputs(1328);
    layer3_outputs(4715) <= (layer2_outputs(2794)) and (layer2_outputs(2890));
    layer3_outputs(4716) <= not(layer2_outputs(628)) or (layer2_outputs(1161));
    layer3_outputs(4717) <= '1';
    layer3_outputs(4718) <= not(layer2_outputs(4068));
    layer3_outputs(4719) <= (layer2_outputs(3429)) and not (layer2_outputs(1403));
    layer3_outputs(4720) <= layer2_outputs(3713);
    layer3_outputs(4721) <= (layer2_outputs(3405)) and not (layer2_outputs(2099));
    layer3_outputs(4722) <= not((layer2_outputs(3647)) and (layer2_outputs(1870)));
    layer3_outputs(4723) <= (layer2_outputs(4922)) and not (layer2_outputs(4933));
    layer3_outputs(4724) <= (layer2_outputs(4059)) xor (layer2_outputs(1346));
    layer3_outputs(4725) <= '1';
    layer3_outputs(4726) <= (layer2_outputs(4820)) or (layer2_outputs(3603));
    layer3_outputs(4727) <= '0';
    layer3_outputs(4728) <= (layer2_outputs(2309)) and not (layer2_outputs(3771));
    layer3_outputs(4729) <= (layer2_outputs(4408)) and not (layer2_outputs(1574));
    layer3_outputs(4730) <= not((layer2_outputs(4994)) and (layer2_outputs(3018)));
    layer3_outputs(4731) <= (layer2_outputs(4266)) and not (layer2_outputs(4879));
    layer3_outputs(4732) <= (layer2_outputs(2972)) and (layer2_outputs(2239));
    layer3_outputs(4733) <= not(layer2_outputs(2121)) or (layer2_outputs(4164));
    layer3_outputs(4734) <= '1';
    layer3_outputs(4735) <= not(layer2_outputs(4827));
    layer3_outputs(4736) <= not(layer2_outputs(3037));
    layer3_outputs(4737) <= (layer2_outputs(2435)) and not (layer2_outputs(3391));
    layer3_outputs(4738) <= (layer2_outputs(2935)) and not (layer2_outputs(286));
    layer3_outputs(4739) <= not(layer2_outputs(4270)) or (layer2_outputs(440));
    layer3_outputs(4740) <= not(layer2_outputs(1200));
    layer3_outputs(4741) <= (layer2_outputs(3928)) or (layer2_outputs(3882));
    layer3_outputs(4742) <= (layer2_outputs(2691)) xor (layer2_outputs(4332));
    layer3_outputs(4743) <= layer2_outputs(2906);
    layer3_outputs(4744) <= not((layer2_outputs(1292)) xor (layer2_outputs(3463)));
    layer3_outputs(4745) <= layer2_outputs(586);
    layer3_outputs(4746) <= not((layer2_outputs(811)) and (layer2_outputs(2592)));
    layer3_outputs(4747) <= not(layer2_outputs(1967));
    layer3_outputs(4748) <= (layer2_outputs(2764)) and (layer2_outputs(4378));
    layer3_outputs(4749) <= layer2_outputs(4825);
    layer3_outputs(4750) <= (layer2_outputs(5003)) and not (layer2_outputs(4711));
    layer3_outputs(4751) <= layer2_outputs(2023);
    layer3_outputs(4752) <= '0';
    layer3_outputs(4753) <= layer2_outputs(462);
    layer3_outputs(4754) <= '1';
    layer3_outputs(4755) <= '0';
    layer3_outputs(4756) <= '0';
    layer3_outputs(4757) <= not(layer2_outputs(4718)) or (layer2_outputs(5098));
    layer3_outputs(4758) <= (layer2_outputs(4122)) or (layer2_outputs(4095));
    layer3_outputs(4759) <= not(layer2_outputs(2314)) or (layer2_outputs(2881));
    layer3_outputs(4760) <= not((layer2_outputs(1792)) or (layer2_outputs(955)));
    layer3_outputs(4761) <= (layer2_outputs(4211)) and (layer2_outputs(3505));
    layer3_outputs(4762) <= not(layer2_outputs(741));
    layer3_outputs(4763) <= '0';
    layer3_outputs(4764) <= not(layer2_outputs(2748)) or (layer2_outputs(1697));
    layer3_outputs(4765) <= '0';
    layer3_outputs(4766) <= not((layer2_outputs(1774)) and (layer2_outputs(1440)));
    layer3_outputs(4767) <= (layer2_outputs(4252)) or (layer2_outputs(1876));
    layer3_outputs(4768) <= not(layer2_outputs(838));
    layer3_outputs(4769) <= (layer2_outputs(1015)) xor (layer2_outputs(696));
    layer3_outputs(4770) <= '1';
    layer3_outputs(4771) <= not((layer2_outputs(3740)) or (layer2_outputs(2868)));
    layer3_outputs(4772) <= not(layer2_outputs(1622));
    layer3_outputs(4773) <= (layer2_outputs(963)) xor (layer2_outputs(2448));
    layer3_outputs(4774) <= not(layer2_outputs(132));
    layer3_outputs(4775) <= '1';
    layer3_outputs(4776) <= (layer2_outputs(4848)) or (layer2_outputs(2686));
    layer3_outputs(4777) <= '1';
    layer3_outputs(4778) <= (layer2_outputs(4800)) and (layer2_outputs(4945));
    layer3_outputs(4779) <= not((layer2_outputs(2414)) xor (layer2_outputs(3105)));
    layer3_outputs(4780) <= not(layer2_outputs(4527)) or (layer2_outputs(710));
    layer3_outputs(4781) <= '1';
    layer3_outputs(4782) <= (layer2_outputs(3923)) and (layer2_outputs(50));
    layer3_outputs(4783) <= not((layer2_outputs(1977)) and (layer2_outputs(533)));
    layer3_outputs(4784) <= (layer2_outputs(919)) and not (layer2_outputs(2098));
    layer3_outputs(4785) <= '0';
    layer3_outputs(4786) <= (layer2_outputs(3365)) and not (layer2_outputs(365));
    layer3_outputs(4787) <= '1';
    layer3_outputs(4788) <= not((layer2_outputs(4486)) or (layer2_outputs(1794)));
    layer3_outputs(4789) <= (layer2_outputs(980)) and (layer2_outputs(2236));
    layer3_outputs(4790) <= not((layer2_outputs(4020)) and (layer2_outputs(841)));
    layer3_outputs(4791) <= (layer2_outputs(2952)) and (layer2_outputs(1715));
    layer3_outputs(4792) <= not(layer2_outputs(3534));
    layer3_outputs(4793) <= not(layer2_outputs(15));
    layer3_outputs(4794) <= (layer2_outputs(1285)) or (layer2_outputs(3086));
    layer3_outputs(4795) <= not(layer2_outputs(971)) or (layer2_outputs(4857));
    layer3_outputs(4796) <= (layer2_outputs(3707)) and (layer2_outputs(2077));
    layer3_outputs(4797) <= (layer2_outputs(1825)) or (layer2_outputs(857));
    layer3_outputs(4798) <= layer2_outputs(4457);
    layer3_outputs(4799) <= not((layer2_outputs(4493)) and (layer2_outputs(5042)));
    layer3_outputs(4800) <= layer2_outputs(1092);
    layer3_outputs(4801) <= layer2_outputs(3570);
    layer3_outputs(4802) <= (layer2_outputs(4104)) and not (layer2_outputs(4851));
    layer3_outputs(4803) <= layer2_outputs(3342);
    layer3_outputs(4804) <= layer2_outputs(4549);
    layer3_outputs(4805) <= layer2_outputs(1401);
    layer3_outputs(4806) <= '1';
    layer3_outputs(4807) <= not((layer2_outputs(4345)) or (layer2_outputs(1532)));
    layer3_outputs(4808) <= not(layer2_outputs(3576));
    layer3_outputs(4809) <= layer2_outputs(1925);
    layer3_outputs(4810) <= '1';
    layer3_outputs(4811) <= (layer2_outputs(3388)) and not (layer2_outputs(3656));
    layer3_outputs(4812) <= '0';
    layer3_outputs(4813) <= not((layer2_outputs(3703)) or (layer2_outputs(53)));
    layer3_outputs(4814) <= (layer2_outputs(1595)) and not (layer2_outputs(1281));
    layer3_outputs(4815) <= (layer2_outputs(2601)) and not (layer2_outputs(2460));
    layer3_outputs(4816) <= layer2_outputs(1733);
    layer3_outputs(4817) <= not(layer2_outputs(1214));
    layer3_outputs(4818) <= not(layer2_outputs(3766));
    layer3_outputs(4819) <= not(layer2_outputs(1594)) or (layer2_outputs(2443));
    layer3_outputs(4820) <= '0';
    layer3_outputs(4821) <= (layer2_outputs(4555)) and (layer2_outputs(3642));
    layer3_outputs(4822) <= not((layer2_outputs(1509)) or (layer2_outputs(1179)));
    layer3_outputs(4823) <= (layer2_outputs(3060)) and not (layer2_outputs(3480));
    layer3_outputs(4824) <= not((layer2_outputs(416)) or (layer2_outputs(4744)));
    layer3_outputs(4825) <= not(layer2_outputs(2722)) or (layer2_outputs(1102));
    layer3_outputs(4826) <= '0';
    layer3_outputs(4827) <= (layer2_outputs(820)) and not (layer2_outputs(4278));
    layer3_outputs(4828) <= (layer2_outputs(5068)) and not (layer2_outputs(96));
    layer3_outputs(4829) <= (layer2_outputs(4312)) and not (layer2_outputs(2653));
    layer3_outputs(4830) <= not((layer2_outputs(893)) or (layer2_outputs(2699)));
    layer3_outputs(4831) <= not(layer2_outputs(2846));
    layer3_outputs(4832) <= not(layer2_outputs(4330)) or (layer2_outputs(2663));
    layer3_outputs(4833) <= '1';
    layer3_outputs(4834) <= not(layer2_outputs(3076));
    layer3_outputs(4835) <= not(layer2_outputs(3596));
    layer3_outputs(4836) <= (layer2_outputs(1790)) and not (layer2_outputs(369));
    layer3_outputs(4837) <= layer2_outputs(782);
    layer3_outputs(4838) <= not(layer2_outputs(264));
    layer3_outputs(4839) <= not(layer2_outputs(4498)) or (layer2_outputs(2557));
    layer3_outputs(4840) <= layer2_outputs(5096);
    layer3_outputs(4841) <= '0';
    layer3_outputs(4842) <= not(layer2_outputs(1131));
    layer3_outputs(4843) <= not(layer2_outputs(4968)) or (layer2_outputs(956));
    layer3_outputs(4844) <= (layer2_outputs(4722)) and not (layer2_outputs(320));
    layer3_outputs(4845) <= not(layer2_outputs(1700)) or (layer2_outputs(4357));
    layer3_outputs(4846) <= (layer2_outputs(3840)) and not (layer2_outputs(309));
    layer3_outputs(4847) <= (layer2_outputs(4033)) and not (layer2_outputs(685));
    layer3_outputs(4848) <= not(layer2_outputs(840)) or (layer2_outputs(4230));
    layer3_outputs(4849) <= layer2_outputs(3719);
    layer3_outputs(4850) <= (layer2_outputs(344)) and (layer2_outputs(2851));
    layer3_outputs(4851) <= not(layer2_outputs(2572));
    layer3_outputs(4852) <= (layer2_outputs(695)) or (layer2_outputs(3031));
    layer3_outputs(4853) <= layer2_outputs(89);
    layer3_outputs(4854) <= '1';
    layer3_outputs(4855) <= (layer2_outputs(1045)) and not (layer2_outputs(520));
    layer3_outputs(4856) <= (layer2_outputs(3320)) xor (layer2_outputs(3747));
    layer3_outputs(4857) <= layer2_outputs(4836);
    layer3_outputs(4858) <= '0';
    layer3_outputs(4859) <= (layer2_outputs(1262)) and not (layer2_outputs(1691));
    layer3_outputs(4860) <= not(layer2_outputs(1528));
    layer3_outputs(4861) <= not((layer2_outputs(311)) and (layer2_outputs(4671)));
    layer3_outputs(4862) <= not((layer2_outputs(1585)) or (layer2_outputs(2579)));
    layer3_outputs(4863) <= '1';
    layer3_outputs(4864) <= not(layer2_outputs(2698)) or (layer2_outputs(443));
    layer3_outputs(4865) <= not(layer2_outputs(1456)) or (layer2_outputs(1653));
    layer3_outputs(4866) <= layer2_outputs(1535);
    layer3_outputs(4867) <= (layer2_outputs(1345)) and not (layer2_outputs(4092));
    layer3_outputs(4868) <= (layer2_outputs(3808)) and not (layer2_outputs(2139));
    layer3_outputs(4869) <= not(layer2_outputs(3789)) or (layer2_outputs(1456));
    layer3_outputs(4870) <= (layer2_outputs(3693)) xor (layer2_outputs(838));
    layer3_outputs(4871) <= (layer2_outputs(3004)) and not (layer2_outputs(745));
    layer3_outputs(4872) <= (layer2_outputs(4153)) and not (layer2_outputs(3535));
    layer3_outputs(4873) <= not((layer2_outputs(1988)) and (layer2_outputs(731)));
    layer3_outputs(4874) <= (layer2_outputs(3275)) xor (layer2_outputs(453));
    layer3_outputs(4875) <= layer2_outputs(2738);
    layer3_outputs(4876) <= (layer2_outputs(333)) and not (layer2_outputs(349));
    layer3_outputs(4877) <= (layer2_outputs(4394)) and (layer2_outputs(1146));
    layer3_outputs(4878) <= '0';
    layer3_outputs(4879) <= (layer2_outputs(2003)) and not (layer2_outputs(4491));
    layer3_outputs(4880) <= (layer2_outputs(3877)) and (layer2_outputs(2413));
    layer3_outputs(4881) <= '1';
    layer3_outputs(4882) <= '0';
    layer3_outputs(4883) <= not(layer2_outputs(3332)) or (layer2_outputs(4729));
    layer3_outputs(4884) <= layer2_outputs(71);
    layer3_outputs(4885) <= not(layer2_outputs(4741)) or (layer2_outputs(4804));
    layer3_outputs(4886) <= not(layer2_outputs(4540));
    layer3_outputs(4887) <= not(layer2_outputs(3679)) or (layer2_outputs(1206));
    layer3_outputs(4888) <= layer2_outputs(1466);
    layer3_outputs(4889) <= '0';
    layer3_outputs(4890) <= not(layer2_outputs(4964));
    layer3_outputs(4891) <= '1';
    layer3_outputs(4892) <= (layer2_outputs(4953)) and (layer2_outputs(3311));
    layer3_outputs(4893) <= layer2_outputs(4552);
    layer3_outputs(4894) <= layer2_outputs(5119);
    layer3_outputs(4895) <= '1';
    layer3_outputs(4896) <= layer2_outputs(1102);
    layer3_outputs(4897) <= not(layer2_outputs(384));
    layer3_outputs(4898) <= not(layer2_outputs(1224)) or (layer2_outputs(3240));
    layer3_outputs(4899) <= not(layer2_outputs(4480));
    layer3_outputs(4900) <= not((layer2_outputs(4234)) or (layer2_outputs(1035)));
    layer3_outputs(4901) <= layer2_outputs(4190);
    layer3_outputs(4902) <= not(layer2_outputs(4023)) or (layer2_outputs(3466));
    layer3_outputs(4903) <= (layer2_outputs(3241)) and not (layer2_outputs(2664));
    layer3_outputs(4904) <= layer2_outputs(2793);
    layer3_outputs(4905) <= not((layer2_outputs(1177)) and (layer2_outputs(3435)));
    layer3_outputs(4906) <= not(layer2_outputs(3991)) or (layer2_outputs(420));
    layer3_outputs(4907) <= '1';
    layer3_outputs(4908) <= layer2_outputs(2405);
    layer3_outputs(4909) <= '1';
    layer3_outputs(4910) <= not(layer2_outputs(1602)) or (layer2_outputs(1427));
    layer3_outputs(4911) <= not((layer2_outputs(4008)) and (layer2_outputs(448)));
    layer3_outputs(4912) <= (layer2_outputs(303)) and (layer2_outputs(4338));
    layer3_outputs(4913) <= not(layer2_outputs(3505)) or (layer2_outputs(3750));
    layer3_outputs(4914) <= not(layer2_outputs(4997)) or (layer2_outputs(1277));
    layer3_outputs(4915) <= not((layer2_outputs(549)) or (layer2_outputs(4185)));
    layer3_outputs(4916) <= (layer2_outputs(1248)) or (layer2_outputs(2860));
    layer3_outputs(4917) <= not((layer2_outputs(3171)) xor (layer2_outputs(2333)));
    layer3_outputs(4918) <= not(layer2_outputs(698)) or (layer2_outputs(5007));
    layer3_outputs(4919) <= (layer2_outputs(4290)) and not (layer2_outputs(986));
    layer3_outputs(4920) <= '1';
    layer3_outputs(4921) <= layer2_outputs(1665);
    layer3_outputs(4922) <= '0';
    layer3_outputs(4923) <= not((layer2_outputs(1743)) xor (layer2_outputs(3061)));
    layer3_outputs(4924) <= (layer2_outputs(2433)) and not (layer2_outputs(2661));
    layer3_outputs(4925) <= not((layer2_outputs(2489)) or (layer2_outputs(2804)));
    layer3_outputs(4926) <= (layer2_outputs(2303)) and not (layer2_outputs(4548));
    layer3_outputs(4927) <= (layer2_outputs(1780)) or (layer2_outputs(4669));
    layer3_outputs(4928) <= (layer2_outputs(3408)) and not (layer2_outputs(2504));
    layer3_outputs(4929) <= (layer2_outputs(4898)) and not (layer2_outputs(3148));
    layer3_outputs(4930) <= not(layer2_outputs(4259));
    layer3_outputs(4931) <= '1';
    layer3_outputs(4932) <= '0';
    layer3_outputs(4933) <= layer2_outputs(232);
    layer3_outputs(4934) <= not((layer2_outputs(544)) and (layer2_outputs(3526)));
    layer3_outputs(4935) <= (layer2_outputs(284)) or (layer2_outputs(1906));
    layer3_outputs(4936) <= not(layer2_outputs(3999)) or (layer2_outputs(4613));
    layer3_outputs(4937) <= not(layer2_outputs(4239));
    layer3_outputs(4938) <= not(layer2_outputs(4142));
    layer3_outputs(4939) <= layer2_outputs(1453);
    layer3_outputs(4940) <= not(layer2_outputs(3528)) or (layer2_outputs(3582));
    layer3_outputs(4941) <= not((layer2_outputs(2133)) or (layer2_outputs(1646)));
    layer3_outputs(4942) <= (layer2_outputs(2394)) and not (layer2_outputs(3705));
    layer3_outputs(4943) <= not(layer2_outputs(4347)) or (layer2_outputs(859));
    layer3_outputs(4944) <= layer2_outputs(3216);
    layer3_outputs(4945) <= (layer2_outputs(1560)) or (layer2_outputs(2131));
    layer3_outputs(4946) <= not((layer2_outputs(4000)) and (layer2_outputs(4293)));
    layer3_outputs(4947) <= (layer2_outputs(691)) and (layer2_outputs(4524));
    layer3_outputs(4948) <= not((layer2_outputs(577)) or (layer2_outputs(4194)));
    layer3_outputs(4949) <= not((layer2_outputs(2293)) and (layer2_outputs(1177)));
    layer3_outputs(4950) <= (layer2_outputs(3610)) or (layer2_outputs(4530));
    layer3_outputs(4951) <= not((layer2_outputs(4131)) and (layer2_outputs(3934)));
    layer3_outputs(4952) <= (layer2_outputs(3047)) and not (layer2_outputs(518));
    layer3_outputs(4953) <= layer2_outputs(3365);
    layer3_outputs(4954) <= not((layer2_outputs(2663)) or (layer2_outputs(3119)));
    layer3_outputs(4955) <= not(layer2_outputs(2737));
    layer3_outputs(4956) <= layer2_outputs(4310);
    layer3_outputs(4957) <= (layer2_outputs(1706)) or (layer2_outputs(4267));
    layer3_outputs(4958) <= not((layer2_outputs(1830)) and (layer2_outputs(3130)));
    layer3_outputs(4959) <= not(layer2_outputs(3574)) or (layer2_outputs(3461));
    layer3_outputs(4960) <= not((layer2_outputs(4416)) and (layer2_outputs(4325)));
    layer3_outputs(4961) <= '0';
    layer3_outputs(4962) <= (layer2_outputs(2647)) and (layer2_outputs(5011));
    layer3_outputs(4963) <= not((layer2_outputs(509)) and (layer2_outputs(1988)));
    layer3_outputs(4964) <= not(layer2_outputs(3051)) or (layer2_outputs(2197));
    layer3_outputs(4965) <= not(layer2_outputs(3488));
    layer3_outputs(4966) <= not(layer2_outputs(1420)) or (layer2_outputs(4891));
    layer3_outputs(4967) <= not(layer2_outputs(4043)) or (layer2_outputs(1648));
    layer3_outputs(4968) <= not(layer2_outputs(2652)) or (layer2_outputs(3403));
    layer3_outputs(4969) <= (layer2_outputs(4768)) xor (layer2_outputs(3434));
    layer3_outputs(4970) <= layer2_outputs(2307);
    layer3_outputs(4971) <= layer2_outputs(1656);
    layer3_outputs(4972) <= (layer2_outputs(1109)) and not (layer2_outputs(3226));
    layer3_outputs(4973) <= layer2_outputs(1493);
    layer3_outputs(4974) <= '0';
    layer3_outputs(4975) <= not(layer2_outputs(2787)) or (layer2_outputs(459));
    layer3_outputs(4976) <= '0';
    layer3_outputs(4977) <= not(layer2_outputs(4634)) or (layer2_outputs(768));
    layer3_outputs(4978) <= not(layer2_outputs(665)) or (layer2_outputs(237));
    layer3_outputs(4979) <= (layer2_outputs(1789)) and not (layer2_outputs(1900));
    layer3_outputs(4980) <= layer2_outputs(4573);
    layer3_outputs(4981) <= not(layer2_outputs(1645)) or (layer2_outputs(171));
    layer3_outputs(4982) <= (layer2_outputs(4223)) and (layer2_outputs(4311));
    layer3_outputs(4983) <= (layer2_outputs(4567)) and not (layer2_outputs(4653));
    layer3_outputs(4984) <= '0';
    layer3_outputs(4985) <= not(layer2_outputs(3760));
    layer3_outputs(4986) <= '1';
    layer3_outputs(4987) <= (layer2_outputs(1817)) or (layer2_outputs(4795));
    layer3_outputs(4988) <= not(layer2_outputs(2165));
    layer3_outputs(4989) <= '0';
    layer3_outputs(4990) <= layer2_outputs(2428);
    layer3_outputs(4991) <= not(layer2_outputs(4912)) or (layer2_outputs(3288));
    layer3_outputs(4992) <= not((layer2_outputs(1600)) or (layer2_outputs(2511)));
    layer3_outputs(4993) <= not((layer2_outputs(8)) and (layer2_outputs(3046)));
    layer3_outputs(4994) <= (layer2_outputs(1848)) or (layer2_outputs(2685));
    layer3_outputs(4995) <= (layer2_outputs(3251)) and not (layer2_outputs(359));
    layer3_outputs(4996) <= (layer2_outputs(3784)) and (layer2_outputs(3548));
    layer3_outputs(4997) <= layer2_outputs(1775);
    layer3_outputs(4998) <= layer2_outputs(3007);
    layer3_outputs(4999) <= '1';
    layer3_outputs(5000) <= '1';
    layer3_outputs(5001) <= (layer2_outputs(205)) and not (layer2_outputs(179));
    layer3_outputs(5002) <= (layer2_outputs(189)) or (layer2_outputs(2260));
    layer3_outputs(5003) <= not(layer2_outputs(2370));
    layer3_outputs(5004) <= layer2_outputs(2897);
    layer3_outputs(5005) <= not((layer2_outputs(0)) or (layer2_outputs(2631)));
    layer3_outputs(5006) <= (layer2_outputs(3436)) and not (layer2_outputs(4053));
    layer3_outputs(5007) <= not((layer2_outputs(63)) and (layer2_outputs(1596)));
    layer3_outputs(5008) <= not(layer2_outputs(1436));
    layer3_outputs(5009) <= (layer2_outputs(443)) and not (layer2_outputs(1583));
    layer3_outputs(5010) <= (layer2_outputs(4708)) and (layer2_outputs(3510));
    layer3_outputs(5011) <= (layer2_outputs(4700)) or (layer2_outputs(2886));
    layer3_outputs(5012) <= not(layer2_outputs(4218));
    layer3_outputs(5013) <= '1';
    layer3_outputs(5014) <= not(layer2_outputs(2213));
    layer3_outputs(5015) <= '1';
    layer3_outputs(5016) <= not((layer2_outputs(4049)) or (layer2_outputs(224)));
    layer3_outputs(5017) <= not(layer2_outputs(3182)) or (layer2_outputs(2941));
    layer3_outputs(5018) <= (layer2_outputs(163)) and (layer2_outputs(1181));
    layer3_outputs(5019) <= (layer2_outputs(808)) xor (layer2_outputs(3746));
    layer3_outputs(5020) <= not((layer2_outputs(304)) or (layer2_outputs(4726)));
    layer3_outputs(5021) <= (layer2_outputs(548)) and not (layer2_outputs(285));
    layer3_outputs(5022) <= '1';
    layer3_outputs(5023) <= (layer2_outputs(2161)) and not (layer2_outputs(2173));
    layer3_outputs(5024) <= (layer2_outputs(4513)) or (layer2_outputs(63));
    layer3_outputs(5025) <= not((layer2_outputs(1099)) and (layer2_outputs(3352)));
    layer3_outputs(5026) <= (layer2_outputs(1861)) and not (layer2_outputs(4670));
    layer3_outputs(5027) <= '0';
    layer3_outputs(5028) <= layer2_outputs(4922);
    layer3_outputs(5029) <= '1';
    layer3_outputs(5030) <= not((layer2_outputs(2021)) or (layer2_outputs(2205)));
    layer3_outputs(5031) <= (layer2_outputs(3307)) and (layer2_outputs(2898));
    layer3_outputs(5032) <= layer2_outputs(4831);
    layer3_outputs(5033) <= layer2_outputs(4445);
    layer3_outputs(5034) <= (layer2_outputs(1059)) and not (layer2_outputs(1628));
    layer3_outputs(5035) <= layer2_outputs(200);
    layer3_outputs(5036) <= layer2_outputs(3344);
    layer3_outputs(5037) <= not(layer2_outputs(1080));
    layer3_outputs(5038) <= not((layer2_outputs(841)) or (layer2_outputs(2994)));
    layer3_outputs(5039) <= layer2_outputs(1847);
    layer3_outputs(5040) <= '0';
    layer3_outputs(5041) <= '1';
    layer3_outputs(5042) <= '1';
    layer3_outputs(5043) <= not((layer2_outputs(3776)) and (layer2_outputs(3516)));
    layer3_outputs(5044) <= not((layer2_outputs(2210)) or (layer2_outputs(484)));
    layer3_outputs(5045) <= layer2_outputs(4748);
    layer3_outputs(5046) <= not(layer2_outputs(562)) or (layer2_outputs(3005));
    layer3_outputs(5047) <= not(layer2_outputs(4452)) or (layer2_outputs(1299));
    layer3_outputs(5048) <= not((layer2_outputs(890)) and (layer2_outputs(2411)));
    layer3_outputs(5049) <= not(layer2_outputs(4707)) or (layer2_outputs(2838));
    layer3_outputs(5050) <= (layer2_outputs(331)) and not (layer2_outputs(4258));
    layer3_outputs(5051) <= not((layer2_outputs(654)) or (layer2_outputs(2487)));
    layer3_outputs(5052) <= (layer2_outputs(3247)) and not (layer2_outputs(2683));
    layer3_outputs(5053) <= '1';
    layer3_outputs(5054) <= layer2_outputs(3988);
    layer3_outputs(5055) <= (layer2_outputs(4615)) and not (layer2_outputs(4203));
    layer3_outputs(5056) <= (layer2_outputs(4444)) xor (layer2_outputs(3804));
    layer3_outputs(5057) <= not((layer2_outputs(3081)) or (layer2_outputs(335)));
    layer3_outputs(5058) <= (layer2_outputs(4504)) and (layer2_outputs(641));
    layer3_outputs(5059) <= not(layer2_outputs(1965)) or (layer2_outputs(3236));
    layer3_outputs(5060) <= '0';
    layer3_outputs(5061) <= layer2_outputs(3220);
    layer3_outputs(5062) <= '0';
    layer3_outputs(5063) <= not(layer2_outputs(2980)) or (layer2_outputs(4243));
    layer3_outputs(5064) <= '1';
    layer3_outputs(5065) <= '1';
    layer3_outputs(5066) <= '0';
    layer3_outputs(5067) <= (layer2_outputs(4535)) and not (layer2_outputs(2849));
    layer3_outputs(5068) <= '1';
    layer3_outputs(5069) <= (layer2_outputs(3916)) and (layer2_outputs(4118));
    layer3_outputs(5070) <= (layer2_outputs(4854)) and not (layer2_outputs(1391));
    layer3_outputs(5071) <= not((layer2_outputs(1406)) xor (layer2_outputs(2862)));
    layer3_outputs(5072) <= (layer2_outputs(1632)) and not (layer2_outputs(596));
    layer3_outputs(5073) <= not(layer2_outputs(4466)) or (layer2_outputs(4791));
    layer3_outputs(5074) <= (layer2_outputs(544)) and (layer2_outputs(4407));
    layer3_outputs(5075) <= '0';
    layer3_outputs(5076) <= (layer2_outputs(981)) xor (layer2_outputs(1302));
    layer3_outputs(5077) <= (layer2_outputs(3362)) and not (layer2_outputs(1796));
    layer3_outputs(5078) <= (layer2_outputs(5082)) or (layer2_outputs(1747));
    layer3_outputs(5079) <= (layer2_outputs(295)) and (layer2_outputs(4562));
    layer3_outputs(5080) <= '0';
    layer3_outputs(5081) <= '1';
    layer3_outputs(5082) <= '0';
    layer3_outputs(5083) <= (layer2_outputs(4369)) or (layer2_outputs(405));
    layer3_outputs(5084) <= not(layer2_outputs(2));
    layer3_outputs(5085) <= '0';
    layer3_outputs(5086) <= not(layer2_outputs(2943)) or (layer2_outputs(4954));
    layer3_outputs(5087) <= layer2_outputs(2965);
    layer3_outputs(5088) <= (layer2_outputs(3859)) and not (layer2_outputs(1766));
    layer3_outputs(5089) <= not(layer2_outputs(3616)) or (layer2_outputs(96));
    layer3_outputs(5090) <= not(layer2_outputs(1659));
    layer3_outputs(5091) <= (layer2_outputs(1292)) or (layer2_outputs(1275));
    layer3_outputs(5092) <= not(layer2_outputs(4610)) or (layer2_outputs(3787));
    layer3_outputs(5093) <= layer2_outputs(2129);
    layer3_outputs(5094) <= not(layer2_outputs(386));
    layer3_outputs(5095) <= not(layer2_outputs(2225)) or (layer2_outputs(1907));
    layer3_outputs(5096) <= not(layer2_outputs(1569)) or (layer2_outputs(3112));
    layer3_outputs(5097) <= not((layer2_outputs(3057)) or (layer2_outputs(2332)));
    layer3_outputs(5098) <= not(layer2_outputs(3700)) or (layer2_outputs(5059));
    layer3_outputs(5099) <= (layer2_outputs(5107)) and not (layer2_outputs(3360));
    layer3_outputs(5100) <= (layer2_outputs(3751)) or (layer2_outputs(1820));
    layer3_outputs(5101) <= '0';
    layer3_outputs(5102) <= not((layer2_outputs(547)) or (layer2_outputs(147)));
    layer3_outputs(5103) <= layer2_outputs(2671);
    layer3_outputs(5104) <= layer2_outputs(3864);
    layer3_outputs(5105) <= layer2_outputs(4486);
    layer3_outputs(5106) <= not(layer2_outputs(3));
    layer3_outputs(5107) <= '1';
    layer3_outputs(5108) <= (layer2_outputs(4629)) and not (layer2_outputs(1894));
    layer3_outputs(5109) <= (layer2_outputs(1044)) or (layer2_outputs(3353));
    layer3_outputs(5110) <= not(layer2_outputs(4625));
    layer3_outputs(5111) <= (layer2_outputs(3709)) and not (layer2_outputs(2944));
    layer3_outputs(5112) <= not(layer2_outputs(2726)) or (layer2_outputs(4897));
    layer3_outputs(5113) <= (layer2_outputs(4687)) or (layer2_outputs(2486));
    layer3_outputs(5114) <= layer2_outputs(4148);
    layer3_outputs(5115) <= (layer2_outputs(2592)) or (layer2_outputs(1732));
    layer3_outputs(5116) <= not(layer2_outputs(213)) or (layer2_outputs(2325));
    layer3_outputs(5117) <= not(layer2_outputs(3115)) or (layer2_outputs(2154));
    layer3_outputs(5118) <= (layer2_outputs(4026)) and not (layer2_outputs(4168));
    layer3_outputs(5119) <= not(layer2_outputs(954));
    layer4_outputs(0) <= not(layer3_outputs(3140));
    layer4_outputs(1) <= (layer3_outputs(3063)) and (layer3_outputs(3869));
    layer4_outputs(2) <= layer3_outputs(1135);
    layer4_outputs(3) <= (layer3_outputs(597)) xor (layer3_outputs(4056));
    layer4_outputs(4) <= not(layer3_outputs(1448)) or (layer3_outputs(4960));
    layer4_outputs(5) <= '0';
    layer4_outputs(6) <= layer3_outputs(2293);
    layer4_outputs(7) <= not((layer3_outputs(3245)) and (layer3_outputs(2211)));
    layer4_outputs(8) <= not((layer3_outputs(3268)) or (layer3_outputs(3334)));
    layer4_outputs(9) <= (layer3_outputs(3166)) or (layer3_outputs(1763));
    layer4_outputs(10) <= '1';
    layer4_outputs(11) <= '1';
    layer4_outputs(12) <= (layer3_outputs(2830)) and not (layer3_outputs(2724));
    layer4_outputs(13) <= not((layer3_outputs(2970)) and (layer3_outputs(242)));
    layer4_outputs(14) <= not((layer3_outputs(3216)) or (layer3_outputs(1302)));
    layer4_outputs(15) <= (layer3_outputs(2982)) and not (layer3_outputs(3029));
    layer4_outputs(16) <= not((layer3_outputs(4481)) or (layer3_outputs(1804)));
    layer4_outputs(17) <= '0';
    layer4_outputs(18) <= not(layer3_outputs(1483));
    layer4_outputs(19) <= not(layer3_outputs(2841));
    layer4_outputs(20) <= (layer3_outputs(79)) and not (layer3_outputs(3265));
    layer4_outputs(21) <= (layer3_outputs(2671)) and not (layer3_outputs(4314));
    layer4_outputs(22) <= not(layer3_outputs(1361));
    layer4_outputs(23) <= '0';
    layer4_outputs(24) <= layer3_outputs(1117);
    layer4_outputs(25) <= not((layer3_outputs(881)) or (layer3_outputs(2829)));
    layer4_outputs(26) <= not(layer3_outputs(4216));
    layer4_outputs(27) <= not((layer3_outputs(810)) and (layer3_outputs(517)));
    layer4_outputs(28) <= not((layer3_outputs(4921)) and (layer3_outputs(1215)));
    layer4_outputs(29) <= (layer3_outputs(4261)) xor (layer3_outputs(1482));
    layer4_outputs(30) <= not(layer3_outputs(3157)) or (layer3_outputs(4670));
    layer4_outputs(31) <= (layer3_outputs(1694)) and not (layer3_outputs(2316));
    layer4_outputs(32) <= not((layer3_outputs(410)) or (layer3_outputs(2953)));
    layer4_outputs(33) <= '1';
    layer4_outputs(34) <= layer3_outputs(2564);
    layer4_outputs(35) <= (layer3_outputs(1784)) xor (layer3_outputs(431));
    layer4_outputs(36) <= layer3_outputs(2252);
    layer4_outputs(37) <= '0';
    layer4_outputs(38) <= not(layer3_outputs(1654));
    layer4_outputs(39) <= not((layer3_outputs(565)) and (layer3_outputs(2253)));
    layer4_outputs(40) <= not((layer3_outputs(1834)) or (layer3_outputs(4809)));
    layer4_outputs(41) <= not(layer3_outputs(1416)) or (layer3_outputs(4056));
    layer4_outputs(42) <= (layer3_outputs(4435)) and (layer3_outputs(293));
    layer4_outputs(43) <= (layer3_outputs(3707)) or (layer3_outputs(2890));
    layer4_outputs(44) <= not(layer3_outputs(3327));
    layer4_outputs(45) <= '0';
    layer4_outputs(46) <= (layer3_outputs(4917)) and not (layer3_outputs(290));
    layer4_outputs(47) <= '1';
    layer4_outputs(48) <= '0';
    layer4_outputs(49) <= '1';
    layer4_outputs(50) <= (layer3_outputs(2095)) and not (layer3_outputs(357));
    layer4_outputs(51) <= (layer3_outputs(74)) and not (layer3_outputs(4180));
    layer4_outputs(52) <= '0';
    layer4_outputs(53) <= layer3_outputs(2603);
    layer4_outputs(54) <= not(layer3_outputs(3749));
    layer4_outputs(55) <= (layer3_outputs(755)) and (layer3_outputs(135));
    layer4_outputs(56) <= not(layer3_outputs(4372));
    layer4_outputs(57) <= layer3_outputs(2923);
    layer4_outputs(58) <= (layer3_outputs(5082)) and not (layer3_outputs(4856));
    layer4_outputs(59) <= (layer3_outputs(801)) and not (layer3_outputs(1783));
    layer4_outputs(60) <= (layer3_outputs(3803)) and not (layer3_outputs(1216));
    layer4_outputs(61) <= (layer3_outputs(4429)) and (layer3_outputs(883));
    layer4_outputs(62) <= not(layer3_outputs(1628));
    layer4_outputs(63) <= layer3_outputs(233);
    layer4_outputs(64) <= not(layer3_outputs(961)) or (layer3_outputs(843));
    layer4_outputs(65) <= (layer3_outputs(437)) and (layer3_outputs(3545));
    layer4_outputs(66) <= not(layer3_outputs(1004));
    layer4_outputs(67) <= not(layer3_outputs(1808));
    layer4_outputs(68) <= '0';
    layer4_outputs(69) <= '0';
    layer4_outputs(70) <= not(layer3_outputs(1225)) or (layer3_outputs(4928));
    layer4_outputs(71) <= (layer3_outputs(4582)) and not (layer3_outputs(4376));
    layer4_outputs(72) <= layer3_outputs(1205);
    layer4_outputs(73) <= '0';
    layer4_outputs(74) <= '0';
    layer4_outputs(75) <= not((layer3_outputs(2884)) or (layer3_outputs(4649)));
    layer4_outputs(76) <= (layer3_outputs(2559)) and not (layer3_outputs(4441));
    layer4_outputs(77) <= layer3_outputs(946);
    layer4_outputs(78) <= not((layer3_outputs(2475)) or (layer3_outputs(365)));
    layer4_outputs(79) <= not(layer3_outputs(2949)) or (layer3_outputs(2112));
    layer4_outputs(80) <= (layer3_outputs(937)) and not (layer3_outputs(3730));
    layer4_outputs(81) <= (layer3_outputs(1152)) and (layer3_outputs(2891));
    layer4_outputs(82) <= (layer3_outputs(4973)) and (layer3_outputs(3057));
    layer4_outputs(83) <= (layer3_outputs(4874)) xor (layer3_outputs(2235));
    layer4_outputs(84) <= layer3_outputs(1892);
    layer4_outputs(85) <= '0';
    layer4_outputs(86) <= layer3_outputs(111);
    layer4_outputs(87) <= not(layer3_outputs(1805));
    layer4_outputs(88) <= (layer3_outputs(1142)) and (layer3_outputs(1801));
    layer4_outputs(89) <= (layer3_outputs(2605)) and not (layer3_outputs(300));
    layer4_outputs(90) <= layer3_outputs(2090);
    layer4_outputs(91) <= (layer3_outputs(174)) and (layer3_outputs(3554));
    layer4_outputs(92) <= (layer3_outputs(1742)) and not (layer3_outputs(2427));
    layer4_outputs(93) <= not(layer3_outputs(3670));
    layer4_outputs(94) <= layer3_outputs(30);
    layer4_outputs(95) <= not((layer3_outputs(3019)) and (layer3_outputs(63)));
    layer4_outputs(96) <= (layer3_outputs(5108)) and not (layer3_outputs(3554));
    layer4_outputs(97) <= not(layer3_outputs(1102));
    layer4_outputs(98) <= '0';
    layer4_outputs(99) <= not(layer3_outputs(1523));
    layer4_outputs(100) <= (layer3_outputs(117)) and not (layer3_outputs(667));
    layer4_outputs(101) <= layer3_outputs(2963);
    layer4_outputs(102) <= not(layer3_outputs(383));
    layer4_outputs(103) <= not(layer3_outputs(1491));
    layer4_outputs(104) <= not(layer3_outputs(4072));
    layer4_outputs(105) <= layer3_outputs(1033);
    layer4_outputs(106) <= not(layer3_outputs(4039));
    layer4_outputs(107) <= (layer3_outputs(3237)) and (layer3_outputs(592));
    layer4_outputs(108) <= layer3_outputs(3081);
    layer4_outputs(109) <= '0';
    layer4_outputs(110) <= not((layer3_outputs(1024)) and (layer3_outputs(3601)));
    layer4_outputs(111) <= (layer3_outputs(5080)) and not (layer3_outputs(1268));
    layer4_outputs(112) <= not(layer3_outputs(884)) or (layer3_outputs(2681));
    layer4_outputs(113) <= not((layer3_outputs(2874)) xor (layer3_outputs(1829)));
    layer4_outputs(114) <= (layer3_outputs(764)) and not (layer3_outputs(1229));
    layer4_outputs(115) <= not(layer3_outputs(3531));
    layer4_outputs(116) <= layer3_outputs(1033);
    layer4_outputs(117) <= not((layer3_outputs(4240)) or (layer3_outputs(247)));
    layer4_outputs(118) <= '0';
    layer4_outputs(119) <= layer3_outputs(4269);
    layer4_outputs(120) <= (layer3_outputs(1584)) or (layer3_outputs(509));
    layer4_outputs(121) <= (layer3_outputs(4061)) and (layer3_outputs(4488));
    layer4_outputs(122) <= not(layer3_outputs(4802)) or (layer3_outputs(1266));
    layer4_outputs(123) <= '0';
    layer4_outputs(124) <= '0';
    layer4_outputs(125) <= not(layer3_outputs(5058)) or (layer3_outputs(3256));
    layer4_outputs(126) <= '1';
    layer4_outputs(127) <= (layer3_outputs(3406)) and not (layer3_outputs(2546));
    layer4_outputs(128) <= not(layer3_outputs(175)) or (layer3_outputs(669));
    layer4_outputs(129) <= (layer3_outputs(1353)) and not (layer3_outputs(3209));
    layer4_outputs(130) <= (layer3_outputs(2346)) xor (layer3_outputs(2530));
    layer4_outputs(131) <= '0';
    layer4_outputs(132) <= layer3_outputs(4484);
    layer4_outputs(133) <= not(layer3_outputs(4810));
    layer4_outputs(134) <= layer3_outputs(440);
    layer4_outputs(135) <= not((layer3_outputs(2610)) xor (layer3_outputs(4956)));
    layer4_outputs(136) <= (layer3_outputs(1982)) or (layer3_outputs(4757));
    layer4_outputs(137) <= '0';
    layer4_outputs(138) <= '0';
    layer4_outputs(139) <= not(layer3_outputs(2142));
    layer4_outputs(140) <= (layer3_outputs(2648)) and not (layer3_outputs(3153));
    layer4_outputs(141) <= '1';
    layer4_outputs(142) <= not(layer3_outputs(1534));
    layer4_outputs(143) <= (layer3_outputs(3658)) and not (layer3_outputs(2029));
    layer4_outputs(144) <= not((layer3_outputs(436)) and (layer3_outputs(1399)));
    layer4_outputs(145) <= '1';
    layer4_outputs(146) <= not(layer3_outputs(324)) or (layer3_outputs(2257));
    layer4_outputs(147) <= layer3_outputs(327);
    layer4_outputs(148) <= not(layer3_outputs(2008)) or (layer3_outputs(137));
    layer4_outputs(149) <= layer3_outputs(608);
    layer4_outputs(150) <= not(layer3_outputs(2697)) or (layer3_outputs(3521));
    layer4_outputs(151) <= (layer3_outputs(3143)) and not (layer3_outputs(4982));
    layer4_outputs(152) <= '1';
    layer4_outputs(153) <= (layer3_outputs(197)) or (layer3_outputs(1023));
    layer4_outputs(154) <= not(layer3_outputs(4590));
    layer4_outputs(155) <= not((layer3_outputs(3927)) or (layer3_outputs(3505)));
    layer4_outputs(156) <= not(layer3_outputs(176));
    layer4_outputs(157) <= not(layer3_outputs(1865)) or (layer3_outputs(1813));
    layer4_outputs(158) <= not(layer3_outputs(3584)) or (layer3_outputs(118));
    layer4_outputs(159) <= not(layer3_outputs(2057));
    layer4_outputs(160) <= not((layer3_outputs(3469)) or (layer3_outputs(3466)));
    layer4_outputs(161) <= not(layer3_outputs(4161)) or (layer3_outputs(3206));
    layer4_outputs(162) <= layer3_outputs(350);
    layer4_outputs(163) <= (layer3_outputs(2736)) and (layer3_outputs(4949));
    layer4_outputs(164) <= layer3_outputs(107);
    layer4_outputs(165) <= not(layer3_outputs(3884));
    layer4_outputs(166) <= (layer3_outputs(4915)) and not (layer3_outputs(4204));
    layer4_outputs(167) <= layer3_outputs(2616);
    layer4_outputs(168) <= not(layer3_outputs(1417)) or (layer3_outputs(2208));
    layer4_outputs(169) <= (layer3_outputs(3007)) and not (layer3_outputs(4295));
    layer4_outputs(170) <= '1';
    layer4_outputs(171) <= layer3_outputs(730);
    layer4_outputs(172) <= (layer3_outputs(95)) or (layer3_outputs(3003));
    layer4_outputs(173) <= (layer3_outputs(3916)) and not (layer3_outputs(4951));
    layer4_outputs(174) <= (layer3_outputs(2018)) and (layer3_outputs(219));
    layer4_outputs(175) <= not(layer3_outputs(2425));
    layer4_outputs(176) <= not(layer3_outputs(783));
    layer4_outputs(177) <= not(layer3_outputs(1252)) or (layer3_outputs(2199));
    layer4_outputs(178) <= (layer3_outputs(3888)) and not (layer3_outputs(2001));
    layer4_outputs(179) <= not(layer3_outputs(2001));
    layer4_outputs(180) <= not(layer3_outputs(3223));
    layer4_outputs(181) <= not((layer3_outputs(3274)) or (layer3_outputs(3242)));
    layer4_outputs(182) <= layer3_outputs(3403);
    layer4_outputs(183) <= not((layer3_outputs(677)) and (layer3_outputs(2885)));
    layer4_outputs(184) <= '1';
    layer4_outputs(185) <= not((layer3_outputs(2904)) and (layer3_outputs(3199)));
    layer4_outputs(186) <= (layer3_outputs(2586)) and not (layer3_outputs(3425));
    layer4_outputs(187) <= layer3_outputs(2091);
    layer4_outputs(188) <= '0';
    layer4_outputs(189) <= layer3_outputs(4390);
    layer4_outputs(190) <= not(layer3_outputs(3188));
    layer4_outputs(191) <= not(layer3_outputs(4530));
    layer4_outputs(192) <= (layer3_outputs(763)) xor (layer3_outputs(3949));
    layer4_outputs(193) <= (layer3_outputs(4359)) and (layer3_outputs(990));
    layer4_outputs(194) <= (layer3_outputs(1475)) or (layer3_outputs(3983));
    layer4_outputs(195) <= not(layer3_outputs(79));
    layer4_outputs(196) <= not(layer3_outputs(109)) or (layer3_outputs(3197));
    layer4_outputs(197) <= not((layer3_outputs(3034)) xor (layer3_outputs(5009)));
    layer4_outputs(198) <= layer3_outputs(4050);
    layer4_outputs(199) <= '0';
    layer4_outputs(200) <= not((layer3_outputs(1652)) or (layer3_outputs(1283)));
    layer4_outputs(201) <= layer3_outputs(3234);
    layer4_outputs(202) <= (layer3_outputs(2791)) and not (layer3_outputs(950));
    layer4_outputs(203) <= (layer3_outputs(1727)) and not (layer3_outputs(4155));
    layer4_outputs(204) <= not(layer3_outputs(2381));
    layer4_outputs(205) <= '0';
    layer4_outputs(206) <= '0';
    layer4_outputs(207) <= not(layer3_outputs(4227)) or (layer3_outputs(4087));
    layer4_outputs(208) <= not(layer3_outputs(4205));
    layer4_outputs(209) <= (layer3_outputs(3739)) and (layer3_outputs(3158));
    layer4_outputs(210) <= '1';
    layer4_outputs(211) <= not(layer3_outputs(1771));
    layer4_outputs(212) <= (layer3_outputs(1465)) and not (layer3_outputs(58));
    layer4_outputs(213) <= not((layer3_outputs(736)) or (layer3_outputs(1739)));
    layer4_outputs(214) <= not((layer3_outputs(602)) or (layer3_outputs(1475)));
    layer4_outputs(215) <= layer3_outputs(1811);
    layer4_outputs(216) <= not((layer3_outputs(4306)) or (layer3_outputs(4544)));
    layer4_outputs(217) <= '1';
    layer4_outputs(218) <= not(layer3_outputs(3512)) or (layer3_outputs(5091));
    layer4_outputs(219) <= not(layer3_outputs(7));
    layer4_outputs(220) <= not(layer3_outputs(817)) or (layer3_outputs(1833));
    layer4_outputs(221) <= (layer3_outputs(3167)) and (layer3_outputs(3187));
    layer4_outputs(222) <= layer3_outputs(1889);
    layer4_outputs(223) <= '0';
    layer4_outputs(224) <= not(layer3_outputs(4596));
    layer4_outputs(225) <= not(layer3_outputs(912));
    layer4_outputs(226) <= (layer3_outputs(4772)) and not (layer3_outputs(305));
    layer4_outputs(227) <= (layer3_outputs(405)) and not (layer3_outputs(4388));
    layer4_outputs(228) <= (layer3_outputs(3647)) and (layer3_outputs(5075));
    layer4_outputs(229) <= layer3_outputs(4645);
    layer4_outputs(230) <= not((layer3_outputs(4615)) and (layer3_outputs(2145)));
    layer4_outputs(231) <= (layer3_outputs(1766)) and not (layer3_outputs(2928));
    layer4_outputs(232) <= (layer3_outputs(3464)) or (layer3_outputs(943));
    layer4_outputs(233) <= not((layer3_outputs(748)) or (layer3_outputs(3652)));
    layer4_outputs(234) <= not((layer3_outputs(1725)) and (layer3_outputs(2502)));
    layer4_outputs(235) <= (layer3_outputs(2734)) and not (layer3_outputs(749));
    layer4_outputs(236) <= not(layer3_outputs(2122)) or (layer3_outputs(3025));
    layer4_outputs(237) <= (layer3_outputs(2364)) and not (layer3_outputs(0));
    layer4_outputs(238) <= (layer3_outputs(895)) and (layer3_outputs(3636));
    layer4_outputs(239) <= not((layer3_outputs(407)) and (layer3_outputs(4754)));
    layer4_outputs(240) <= not(layer3_outputs(3493)) or (layer3_outputs(3876));
    layer4_outputs(241) <= (layer3_outputs(3501)) and (layer3_outputs(905));
    layer4_outputs(242) <= layer3_outputs(4961);
    layer4_outputs(243) <= layer3_outputs(927);
    layer4_outputs(244) <= (layer3_outputs(2688)) and (layer3_outputs(3132));
    layer4_outputs(245) <= not((layer3_outputs(1024)) and (layer3_outputs(1387)));
    layer4_outputs(246) <= not(layer3_outputs(3594)) or (layer3_outputs(3516));
    layer4_outputs(247) <= (layer3_outputs(3504)) and not (layer3_outputs(3779));
    layer4_outputs(248) <= not((layer3_outputs(2046)) or (layer3_outputs(1864)));
    layer4_outputs(249) <= (layer3_outputs(2674)) and (layer3_outputs(5030));
    layer4_outputs(250) <= not((layer3_outputs(972)) or (layer3_outputs(4885)));
    layer4_outputs(251) <= not(layer3_outputs(3348)) or (layer3_outputs(3178));
    layer4_outputs(252) <= (layer3_outputs(338)) or (layer3_outputs(3236));
    layer4_outputs(253) <= '1';
    layer4_outputs(254) <= not((layer3_outputs(4548)) or (layer3_outputs(2260)));
    layer4_outputs(255) <= (layer3_outputs(1651)) and not (layer3_outputs(662));
    layer4_outputs(256) <= layer3_outputs(2055);
    layer4_outputs(257) <= not(layer3_outputs(1098)) or (layer3_outputs(4767));
    layer4_outputs(258) <= not(layer3_outputs(1696));
    layer4_outputs(259) <= not(layer3_outputs(2135));
    layer4_outputs(260) <= (layer3_outputs(2574)) and not (layer3_outputs(3707));
    layer4_outputs(261) <= not(layer3_outputs(2233)) or (layer3_outputs(988));
    layer4_outputs(262) <= '0';
    layer4_outputs(263) <= not(layer3_outputs(4234)) or (layer3_outputs(4138));
    layer4_outputs(264) <= (layer3_outputs(2460)) and not (layer3_outputs(2825));
    layer4_outputs(265) <= layer3_outputs(2977);
    layer4_outputs(266) <= (layer3_outputs(1549)) and (layer3_outputs(996));
    layer4_outputs(267) <= (layer3_outputs(3562)) or (layer3_outputs(2222));
    layer4_outputs(268) <= (layer3_outputs(3715)) and (layer3_outputs(2938));
    layer4_outputs(269) <= not((layer3_outputs(2306)) and (layer3_outputs(96)));
    layer4_outputs(270) <= layer3_outputs(68);
    layer4_outputs(271) <= not((layer3_outputs(2099)) or (layer3_outputs(468)));
    layer4_outputs(272) <= not((layer3_outputs(2966)) and (layer3_outputs(3508)));
    layer4_outputs(273) <= not((layer3_outputs(3921)) xor (layer3_outputs(2795)));
    layer4_outputs(274) <= not(layer3_outputs(250));
    layer4_outputs(275) <= not((layer3_outputs(1543)) or (layer3_outputs(1266)));
    layer4_outputs(276) <= '0';
    layer4_outputs(277) <= (layer3_outputs(1422)) and not (layer3_outputs(1722));
    layer4_outputs(278) <= (layer3_outputs(3753)) and (layer3_outputs(1368));
    layer4_outputs(279) <= '1';
    layer4_outputs(280) <= not(layer3_outputs(2193)) or (layer3_outputs(2861));
    layer4_outputs(281) <= (layer3_outputs(3932)) or (layer3_outputs(3589));
    layer4_outputs(282) <= not(layer3_outputs(1615));
    layer4_outputs(283) <= not(layer3_outputs(4697));
    layer4_outputs(284) <= not(layer3_outputs(1918)) or (layer3_outputs(4128));
    layer4_outputs(285) <= not(layer3_outputs(3775));
    layer4_outputs(286) <= (layer3_outputs(657)) and (layer3_outputs(781));
    layer4_outputs(287) <= '1';
    layer4_outputs(288) <= not(layer3_outputs(3875)) or (layer3_outputs(2547));
    layer4_outputs(289) <= '1';
    layer4_outputs(290) <= '1';
    layer4_outputs(291) <= not(layer3_outputs(3655));
    layer4_outputs(292) <= not(layer3_outputs(2310)) or (layer3_outputs(3896));
    layer4_outputs(293) <= (layer3_outputs(1252)) and not (layer3_outputs(3696));
    layer4_outputs(294) <= not(layer3_outputs(1936)) or (layer3_outputs(3694));
    layer4_outputs(295) <= '1';
    layer4_outputs(296) <= not(layer3_outputs(2399));
    layer4_outputs(297) <= layer3_outputs(5021);
    layer4_outputs(298) <= (layer3_outputs(43)) and not (layer3_outputs(3474));
    layer4_outputs(299) <= layer3_outputs(2671);
    layer4_outputs(300) <= '0';
    layer4_outputs(301) <= '0';
    layer4_outputs(302) <= not(layer3_outputs(4672));
    layer4_outputs(303) <= not((layer3_outputs(1332)) or (layer3_outputs(3807)));
    layer4_outputs(304) <= not(layer3_outputs(3778));
    layer4_outputs(305) <= '1';
    layer4_outputs(306) <= layer3_outputs(2923);
    layer4_outputs(307) <= (layer3_outputs(4829)) or (layer3_outputs(2409));
    layer4_outputs(308) <= layer3_outputs(4241);
    layer4_outputs(309) <= (layer3_outputs(1234)) and not (layer3_outputs(2275));
    layer4_outputs(310) <= not(layer3_outputs(4076)) or (layer3_outputs(77));
    layer4_outputs(311) <= (layer3_outputs(4257)) and (layer3_outputs(1258));
    layer4_outputs(312) <= '0';
    layer4_outputs(313) <= not(layer3_outputs(3054)) or (layer3_outputs(4603));
    layer4_outputs(314) <= '0';
    layer4_outputs(315) <= layer3_outputs(4580);
    layer4_outputs(316) <= not(layer3_outputs(4643)) or (layer3_outputs(181));
    layer4_outputs(317) <= not((layer3_outputs(4119)) and (layer3_outputs(513)));
    layer4_outputs(318) <= (layer3_outputs(2616)) and not (layer3_outputs(3421));
    layer4_outputs(319) <= layer3_outputs(3407);
    layer4_outputs(320) <= '1';
    layer4_outputs(321) <= not(layer3_outputs(106));
    layer4_outputs(322) <= '0';
    layer4_outputs(323) <= '0';
    layer4_outputs(324) <= layer3_outputs(2183);
    layer4_outputs(325) <= (layer3_outputs(720)) or (layer3_outputs(4938));
    layer4_outputs(326) <= '0';
    layer4_outputs(327) <= (layer3_outputs(2573)) and not (layer3_outputs(5097));
    layer4_outputs(328) <= '1';
    layer4_outputs(329) <= not(layer3_outputs(398)) or (layer3_outputs(3248));
    layer4_outputs(330) <= (layer3_outputs(3303)) and not (layer3_outputs(1026));
    layer4_outputs(331) <= not((layer3_outputs(248)) and (layer3_outputs(1035)));
    layer4_outputs(332) <= not(layer3_outputs(1495));
    layer4_outputs(333) <= not(layer3_outputs(1863)) or (layer3_outputs(4374));
    layer4_outputs(334) <= not(layer3_outputs(4092));
    layer4_outputs(335) <= not(layer3_outputs(2660));
    layer4_outputs(336) <= (layer3_outputs(3607)) and not (layer3_outputs(1374));
    layer4_outputs(337) <= (layer3_outputs(3998)) and (layer3_outputs(771));
    layer4_outputs(338) <= not((layer3_outputs(4016)) and (layer3_outputs(4233)));
    layer4_outputs(339) <= (layer3_outputs(223)) and (layer3_outputs(1406));
    layer4_outputs(340) <= not(layer3_outputs(1498)) or (layer3_outputs(1710));
    layer4_outputs(341) <= (layer3_outputs(2060)) and not (layer3_outputs(2672));
    layer4_outputs(342) <= not(layer3_outputs(1606)) or (layer3_outputs(3841));
    layer4_outputs(343) <= not(layer3_outputs(3934));
    layer4_outputs(344) <= not((layer3_outputs(4244)) and (layer3_outputs(4796)));
    layer4_outputs(345) <= not(layer3_outputs(2731));
    layer4_outputs(346) <= (layer3_outputs(4084)) and (layer3_outputs(758));
    layer4_outputs(347) <= layer3_outputs(2063);
    layer4_outputs(348) <= (layer3_outputs(3287)) or (layer3_outputs(1668));
    layer4_outputs(349) <= not(layer3_outputs(4793));
    layer4_outputs(350) <= (layer3_outputs(3243)) and not (layer3_outputs(382));
    layer4_outputs(351) <= (layer3_outputs(3529)) xor (layer3_outputs(3085));
    layer4_outputs(352) <= (layer3_outputs(3271)) or (layer3_outputs(962));
    layer4_outputs(353) <= not((layer3_outputs(561)) and (layer3_outputs(2797)));
    layer4_outputs(354) <= not(layer3_outputs(154)) or (layer3_outputs(1040));
    layer4_outputs(355) <= (layer3_outputs(1891)) and not (layer3_outputs(3459));
    layer4_outputs(356) <= layer3_outputs(2996);
    layer4_outputs(357) <= (layer3_outputs(1263)) or (layer3_outputs(416));
    layer4_outputs(358) <= not(layer3_outputs(3444));
    layer4_outputs(359) <= not(layer3_outputs(4997));
    layer4_outputs(360) <= not(layer3_outputs(347));
    layer4_outputs(361) <= layer3_outputs(1066);
    layer4_outputs(362) <= (layer3_outputs(1309)) or (layer3_outputs(2114));
    layer4_outputs(363) <= not(layer3_outputs(4134)) or (layer3_outputs(3769));
    layer4_outputs(364) <= not((layer3_outputs(3349)) or (layer3_outputs(1850)));
    layer4_outputs(365) <= '0';
    layer4_outputs(366) <= (layer3_outputs(5072)) or (layer3_outputs(3007));
    layer4_outputs(367) <= '0';
    layer4_outputs(368) <= not(layer3_outputs(3790));
    layer4_outputs(369) <= (layer3_outputs(2628)) and not (layer3_outputs(2159));
    layer4_outputs(370) <= not(layer3_outputs(261));
    layer4_outputs(371) <= not(layer3_outputs(5010)) or (layer3_outputs(2717));
    layer4_outputs(372) <= '0';
    layer4_outputs(373) <= (layer3_outputs(1070)) and not (layer3_outputs(356));
    layer4_outputs(374) <= layer3_outputs(4185);
    layer4_outputs(375) <= '1';
    layer4_outputs(376) <= not(layer3_outputs(1620));
    layer4_outputs(377) <= layer3_outputs(1656);
    layer4_outputs(378) <= layer3_outputs(1215);
    layer4_outputs(379) <= not(layer3_outputs(832)) or (layer3_outputs(364));
    layer4_outputs(380) <= not(layer3_outputs(3881)) or (layer3_outputs(2886));
    layer4_outputs(381) <= not(layer3_outputs(256)) or (layer3_outputs(2248));
    layer4_outputs(382) <= (layer3_outputs(2749)) or (layer3_outputs(352));
    layer4_outputs(383) <= not((layer3_outputs(5023)) or (layer3_outputs(2760)));
    layer4_outputs(384) <= (layer3_outputs(4392)) and not (layer3_outputs(3562));
    layer4_outputs(385) <= (layer3_outputs(2376)) and not (layer3_outputs(4399));
    layer4_outputs(386) <= not((layer3_outputs(792)) and (layer3_outputs(3569)));
    layer4_outputs(387) <= not((layer3_outputs(3190)) and (layer3_outputs(4391)));
    layer4_outputs(388) <= (layer3_outputs(4237)) and not (layer3_outputs(4674));
    layer4_outputs(389) <= not((layer3_outputs(3681)) and (layer3_outputs(4945)));
    layer4_outputs(390) <= layer3_outputs(2308);
    layer4_outputs(391) <= (layer3_outputs(2373)) or (layer3_outputs(1913));
    layer4_outputs(392) <= not(layer3_outputs(2020)) or (layer3_outputs(4163));
    layer4_outputs(393) <= not(layer3_outputs(4492));
    layer4_outputs(394) <= (layer3_outputs(1754)) and (layer3_outputs(100));
    layer4_outputs(395) <= layer3_outputs(1494);
    layer4_outputs(396) <= layer3_outputs(2969);
    layer4_outputs(397) <= layer3_outputs(730);
    layer4_outputs(398) <= (layer3_outputs(390)) and not (layer3_outputs(3268));
    layer4_outputs(399) <= not(layer3_outputs(1331)) or (layer3_outputs(4946));
    layer4_outputs(400) <= layer3_outputs(3617);
    layer4_outputs(401) <= (layer3_outputs(2784)) and (layer3_outputs(3118));
    layer4_outputs(402) <= layer3_outputs(2509);
    layer4_outputs(403) <= '1';
    layer4_outputs(404) <= not(layer3_outputs(4129));
    layer4_outputs(405) <= not(layer3_outputs(4169));
    layer4_outputs(406) <= (layer3_outputs(4324)) and not (layer3_outputs(1158));
    layer4_outputs(407) <= not(layer3_outputs(3830)) or (layer3_outputs(1093));
    layer4_outputs(408) <= '0';
    layer4_outputs(409) <= not(layer3_outputs(4090)) or (layer3_outputs(2078));
    layer4_outputs(410) <= (layer3_outputs(2318)) or (layer3_outputs(545));
    layer4_outputs(411) <= (layer3_outputs(3843)) and not (layer3_outputs(3304));
    layer4_outputs(412) <= not((layer3_outputs(1610)) or (layer3_outputs(1175)));
    layer4_outputs(413) <= not(layer3_outputs(3550)) or (layer3_outputs(2373));
    layer4_outputs(414) <= not((layer3_outputs(3930)) or (layer3_outputs(710)));
    layer4_outputs(415) <= not((layer3_outputs(2542)) and (layer3_outputs(5116)));
    layer4_outputs(416) <= (layer3_outputs(1957)) or (layer3_outputs(3793));
    layer4_outputs(417) <= '1';
    layer4_outputs(418) <= layer3_outputs(1663);
    layer4_outputs(419) <= (layer3_outputs(1365)) and not (layer3_outputs(89));
    layer4_outputs(420) <= not(layer3_outputs(2128));
    layer4_outputs(421) <= (layer3_outputs(3792)) and not (layer3_outputs(5081));
    layer4_outputs(422) <= not(layer3_outputs(1891)) or (layer3_outputs(3099));
    layer4_outputs(423) <= (layer3_outputs(1316)) and (layer3_outputs(490));
    layer4_outputs(424) <= (layer3_outputs(5066)) and not (layer3_outputs(2951));
    layer4_outputs(425) <= not(layer3_outputs(2668));
    layer4_outputs(426) <= '0';
    layer4_outputs(427) <= not((layer3_outputs(4180)) or (layer3_outputs(3933)));
    layer4_outputs(428) <= not((layer3_outputs(2699)) or (layer3_outputs(1132)));
    layer4_outputs(429) <= '1';
    layer4_outputs(430) <= '1';
    layer4_outputs(431) <= (layer3_outputs(4450)) and not (layer3_outputs(4790));
    layer4_outputs(432) <= not((layer3_outputs(4047)) and (layer3_outputs(3532)));
    layer4_outputs(433) <= '0';
    layer4_outputs(434) <= (layer3_outputs(190)) or (layer3_outputs(2538));
    layer4_outputs(435) <= not(layer3_outputs(1384));
    layer4_outputs(436) <= not(layer3_outputs(4373)) or (layer3_outputs(2863));
    layer4_outputs(437) <= not(layer3_outputs(2816)) or (layer3_outputs(3656));
    layer4_outputs(438) <= '1';
    layer4_outputs(439) <= not(layer3_outputs(3612));
    layer4_outputs(440) <= (layer3_outputs(3984)) and not (layer3_outputs(2047));
    layer4_outputs(441) <= (layer3_outputs(1251)) and not (layer3_outputs(564));
    layer4_outputs(442) <= '1';
    layer4_outputs(443) <= not((layer3_outputs(4691)) or (layer3_outputs(5028)));
    layer4_outputs(444) <= layer3_outputs(876);
    layer4_outputs(445) <= '1';
    layer4_outputs(446) <= not(layer3_outputs(1934));
    layer4_outputs(447) <= '1';
    layer4_outputs(448) <= (layer3_outputs(3047)) and not (layer3_outputs(418));
    layer4_outputs(449) <= layer3_outputs(3020);
    layer4_outputs(450) <= layer3_outputs(1203);
    layer4_outputs(451) <= not(layer3_outputs(2121));
    layer4_outputs(452) <= not(layer3_outputs(1764)) or (layer3_outputs(616));
    layer4_outputs(453) <= not(layer3_outputs(183));
    layer4_outputs(454) <= not((layer3_outputs(2660)) xor (layer3_outputs(1443)));
    layer4_outputs(455) <= layer3_outputs(3014);
    layer4_outputs(456) <= not(layer3_outputs(1521)) or (layer3_outputs(47));
    layer4_outputs(457) <= (layer3_outputs(2948)) and not (layer3_outputs(3174));
    layer4_outputs(458) <= not(layer3_outputs(3353)) or (layer3_outputs(2107));
    layer4_outputs(459) <= '1';
    layer4_outputs(460) <= '0';
    layer4_outputs(461) <= (layer3_outputs(1702)) and not (layer3_outputs(4300));
    layer4_outputs(462) <= layer3_outputs(451);
    layer4_outputs(463) <= not(layer3_outputs(1901));
    layer4_outputs(464) <= '0';
    layer4_outputs(465) <= (layer3_outputs(3843)) xor (layer3_outputs(1856));
    layer4_outputs(466) <= not((layer3_outputs(1888)) or (layer3_outputs(4281)));
    layer4_outputs(467) <= not(layer3_outputs(2117));
    layer4_outputs(468) <= layer3_outputs(3485);
    layer4_outputs(469) <= (layer3_outputs(3336)) and (layer3_outputs(1231));
    layer4_outputs(470) <= not(layer3_outputs(5062));
    layer4_outputs(471) <= '1';
    layer4_outputs(472) <= not(layer3_outputs(1351));
    layer4_outputs(473) <= (layer3_outputs(525)) and (layer3_outputs(1666));
    layer4_outputs(474) <= not(layer3_outputs(4557));
    layer4_outputs(475) <= not(layer3_outputs(1318)) or (layer3_outputs(1041));
    layer4_outputs(476) <= not(layer3_outputs(2030)) or (layer3_outputs(2667));
    layer4_outputs(477) <= (layer3_outputs(1860)) or (layer3_outputs(3123));
    layer4_outputs(478) <= (layer3_outputs(2983)) and not (layer3_outputs(4058));
    layer4_outputs(479) <= '0';
    layer4_outputs(480) <= not((layer3_outputs(2654)) and (layer3_outputs(807)));
    layer4_outputs(481) <= (layer3_outputs(3318)) and not (layer3_outputs(2664));
    layer4_outputs(482) <= not(layer3_outputs(2937)) or (layer3_outputs(4489));
    layer4_outputs(483) <= '1';
    layer4_outputs(484) <= '1';
    layer4_outputs(485) <= layer3_outputs(4307);
    layer4_outputs(486) <= (layer3_outputs(558)) or (layer3_outputs(4687));
    layer4_outputs(487) <= not(layer3_outputs(3569));
    layer4_outputs(488) <= '0';
    layer4_outputs(489) <= layer3_outputs(2230);
    layer4_outputs(490) <= not((layer3_outputs(944)) xor (layer3_outputs(667)));
    layer4_outputs(491) <= (layer3_outputs(3452)) and not (layer3_outputs(2463));
    layer4_outputs(492) <= not(layer3_outputs(3267));
    layer4_outputs(493) <= not(layer3_outputs(2701));
    layer4_outputs(494) <= layer3_outputs(4366);
    layer4_outputs(495) <= not(layer3_outputs(663));
    layer4_outputs(496) <= not(layer3_outputs(2165));
    layer4_outputs(497) <= (layer3_outputs(2832)) and (layer3_outputs(3766));
    layer4_outputs(498) <= '1';
    layer4_outputs(499) <= (layer3_outputs(889)) and (layer3_outputs(4476));
    layer4_outputs(500) <= not(layer3_outputs(2284)) or (layer3_outputs(3492));
    layer4_outputs(501) <= layer3_outputs(4518);
    layer4_outputs(502) <= not(layer3_outputs(2043)) or (layer3_outputs(2780));
    layer4_outputs(503) <= (layer3_outputs(2623)) xor (layer3_outputs(3579));
    layer4_outputs(504) <= not((layer3_outputs(578)) or (layer3_outputs(1790)));
    layer4_outputs(505) <= not((layer3_outputs(2370)) and (layer3_outputs(2395)));
    layer4_outputs(506) <= not(layer3_outputs(1772));
    layer4_outputs(507) <= (layer3_outputs(1009)) and not (layer3_outputs(4816));
    layer4_outputs(508) <= (layer3_outputs(3030)) or (layer3_outputs(3922));
    layer4_outputs(509) <= not((layer3_outputs(1845)) xor (layer3_outputs(2960)));
    layer4_outputs(510) <= not(layer3_outputs(2236));
    layer4_outputs(511) <= (layer3_outputs(3786)) and (layer3_outputs(1542));
    layer4_outputs(512) <= (layer3_outputs(2567)) and not (layer3_outputs(591));
    layer4_outputs(513) <= (layer3_outputs(2969)) xor (layer3_outputs(2216));
    layer4_outputs(514) <= (layer3_outputs(3680)) xor (layer3_outputs(2998));
    layer4_outputs(515) <= not((layer3_outputs(3679)) and (layer3_outputs(5040)));
    layer4_outputs(516) <= not((layer3_outputs(2729)) and (layer3_outputs(2634)));
    layer4_outputs(517) <= not((layer3_outputs(4360)) or (layer3_outputs(645)));
    layer4_outputs(518) <= not(layer3_outputs(2025)) or (layer3_outputs(3475));
    layer4_outputs(519) <= not(layer3_outputs(1450));
    layer4_outputs(520) <= (layer3_outputs(1724)) and not (layer3_outputs(4981));
    layer4_outputs(521) <= not(layer3_outputs(4074));
    layer4_outputs(522) <= (layer3_outputs(930)) and not (layer3_outputs(4405));
    layer4_outputs(523) <= (layer3_outputs(1745)) and (layer3_outputs(1273));
    layer4_outputs(524) <= (layer3_outputs(1720)) or (layer3_outputs(3574));
    layer4_outputs(525) <= (layer3_outputs(875)) or (layer3_outputs(123));
    layer4_outputs(526) <= not(layer3_outputs(1975)) or (layer3_outputs(4521));
    layer4_outputs(527) <= '0';
    layer4_outputs(528) <= layer3_outputs(4485);
    layer4_outputs(529) <= not(layer3_outputs(4273));
    layer4_outputs(530) <= (layer3_outputs(1126)) or (layer3_outputs(802));
    layer4_outputs(531) <= (layer3_outputs(1163)) and (layer3_outputs(2313));
    layer4_outputs(532) <= layer3_outputs(853);
    layer4_outputs(533) <= (layer3_outputs(1819)) and not (layer3_outputs(3915));
    layer4_outputs(534) <= (layer3_outputs(2096)) and not (layer3_outputs(2727));
    layer4_outputs(535) <= not(layer3_outputs(267)) or (layer3_outputs(4171));
    layer4_outputs(536) <= not(layer3_outputs(3511)) or (layer3_outputs(13));
    layer4_outputs(537) <= (layer3_outputs(2441)) or (layer3_outputs(1472));
    layer4_outputs(538) <= (layer3_outputs(3377)) and (layer3_outputs(4344));
    layer4_outputs(539) <= not((layer3_outputs(4827)) xor (layer3_outputs(226)));
    layer4_outputs(540) <= (layer3_outputs(5060)) and not (layer3_outputs(1435));
    layer4_outputs(541) <= (layer3_outputs(419)) and not (layer3_outputs(3436));
    layer4_outputs(542) <= (layer3_outputs(4768)) or (layer3_outputs(743));
    layer4_outputs(543) <= (layer3_outputs(3724)) and (layer3_outputs(4390));
    layer4_outputs(544) <= not(layer3_outputs(992));
    layer4_outputs(545) <= not(layer3_outputs(2982)) or (layer3_outputs(428));
    layer4_outputs(546) <= (layer3_outputs(2966)) and (layer3_outputs(4190));
    layer4_outputs(547) <= not(layer3_outputs(3292)) or (layer3_outputs(4682));
    layer4_outputs(548) <= '0';
    layer4_outputs(549) <= (layer3_outputs(333)) and (layer3_outputs(3725));
    layer4_outputs(550) <= (layer3_outputs(102)) and not (layer3_outputs(1570));
    layer4_outputs(551) <= layer3_outputs(4052);
    layer4_outputs(552) <= not((layer3_outputs(2308)) or (layer3_outputs(642)));
    layer4_outputs(553) <= not(layer3_outputs(1357)) or (layer3_outputs(4067));
    layer4_outputs(554) <= '1';
    layer4_outputs(555) <= not(layer3_outputs(3437)) or (layer3_outputs(2900));
    layer4_outputs(556) <= (layer3_outputs(2794)) or (layer3_outputs(2539));
    layer4_outputs(557) <= not((layer3_outputs(723)) or (layer3_outputs(3288)));
    layer4_outputs(558) <= layer3_outputs(5100);
    layer4_outputs(559) <= (layer3_outputs(2234)) and not (layer3_outputs(1927));
    layer4_outputs(560) <= (layer3_outputs(4164)) or (layer3_outputs(3875));
    layer4_outputs(561) <= '0';
    layer4_outputs(562) <= (layer3_outputs(2484)) or (layer3_outputs(4523));
    layer4_outputs(563) <= '0';
    layer4_outputs(564) <= (layer3_outputs(3812)) and (layer3_outputs(3431));
    layer4_outputs(565) <= not(layer3_outputs(3433)) or (layer3_outputs(3032));
    layer4_outputs(566) <= not(layer3_outputs(3806));
    layer4_outputs(567) <= not(layer3_outputs(4591)) or (layer3_outputs(3620));
    layer4_outputs(568) <= (layer3_outputs(1219)) and not (layer3_outputs(465));
    layer4_outputs(569) <= not(layer3_outputs(2433));
    layer4_outputs(570) <= not(layer3_outputs(1365));
    layer4_outputs(571) <= (layer3_outputs(1462)) and (layer3_outputs(980));
    layer4_outputs(572) <= not((layer3_outputs(3865)) and (layer3_outputs(3685)));
    layer4_outputs(573) <= not(layer3_outputs(3042)) or (layer3_outputs(4097));
    layer4_outputs(574) <= (layer3_outputs(2723)) and not (layer3_outputs(788));
    layer4_outputs(575) <= layer3_outputs(1643);
    layer4_outputs(576) <= not((layer3_outputs(2499)) or (layer3_outputs(4291)));
    layer4_outputs(577) <= (layer3_outputs(332)) or (layer3_outputs(3507));
    layer4_outputs(578) <= (layer3_outputs(3705)) or (layer3_outputs(3382));
    layer4_outputs(579) <= '0';
    layer4_outputs(580) <= not((layer3_outputs(232)) or (layer3_outputs(5105)));
    layer4_outputs(581) <= not((layer3_outputs(1529)) or (layer3_outputs(580)));
    layer4_outputs(582) <= (layer3_outputs(2575)) xor (layer3_outputs(4931));
    layer4_outputs(583) <= not(layer3_outputs(1788));
    layer4_outputs(584) <= not(layer3_outputs(301));
    layer4_outputs(585) <= not(layer3_outputs(296)) or (layer3_outputs(1792));
    layer4_outputs(586) <= (layer3_outputs(5038)) and not (layer3_outputs(1755));
    layer4_outputs(587) <= not(layer3_outputs(4193));
    layer4_outputs(588) <= (layer3_outputs(3695)) and (layer3_outputs(53));
    layer4_outputs(589) <= layer3_outputs(3622);
    layer4_outputs(590) <= (layer3_outputs(524)) and not (layer3_outputs(3626));
    layer4_outputs(591) <= not((layer3_outputs(3918)) and (layer3_outputs(4716)));
    layer4_outputs(592) <= not(layer3_outputs(1897));
    layer4_outputs(593) <= layer3_outputs(2229);
    layer4_outputs(594) <= (layer3_outputs(1400)) and not (layer3_outputs(2510));
    layer4_outputs(595) <= not(layer3_outputs(3250)) or (layer3_outputs(4952));
    layer4_outputs(596) <= not((layer3_outputs(3125)) and (layer3_outputs(1205)));
    layer4_outputs(597) <= (layer3_outputs(4369)) and not (layer3_outputs(2071));
    layer4_outputs(598) <= (layer3_outputs(2917)) and (layer3_outputs(3672));
    layer4_outputs(599) <= layer3_outputs(116);
    layer4_outputs(600) <= '0';
    layer4_outputs(601) <= layer3_outputs(329);
    layer4_outputs(602) <= '0';
    layer4_outputs(603) <= not((layer3_outputs(2498)) and (layer3_outputs(3608)));
    layer4_outputs(604) <= not((layer3_outputs(2255)) and (layer3_outputs(2598)));
    layer4_outputs(605) <= (layer3_outputs(2646)) or (layer3_outputs(1533));
    layer4_outputs(606) <= (layer3_outputs(718)) and not (layer3_outputs(1439));
    layer4_outputs(607) <= '0';
    layer4_outputs(608) <= layer3_outputs(2089);
    layer4_outputs(609) <= (layer3_outputs(5073)) or (layer3_outputs(1084));
    layer4_outputs(610) <= (layer3_outputs(1300)) xor (layer3_outputs(1043));
    layer4_outputs(611) <= not((layer3_outputs(3341)) and (layer3_outputs(1689)));
    layer4_outputs(612) <= '0';
    layer4_outputs(613) <= layer3_outputs(1576);
    layer4_outputs(614) <= (layer3_outputs(2276)) and (layer3_outputs(4246));
    layer4_outputs(615) <= not(layer3_outputs(185));
    layer4_outputs(616) <= not(layer3_outputs(1569));
    layer4_outputs(617) <= (layer3_outputs(246)) or (layer3_outputs(4137));
    layer4_outputs(618) <= '1';
    layer4_outputs(619) <= layer3_outputs(2939);
    layer4_outputs(620) <= layer3_outputs(654);
    layer4_outputs(621) <= layer3_outputs(4353);
    layer4_outputs(622) <= (layer3_outputs(2872)) and not (layer3_outputs(4487));
    layer4_outputs(623) <= not(layer3_outputs(1158)) or (layer3_outputs(1426));
    layer4_outputs(624) <= layer3_outputs(3566);
    layer4_outputs(625) <= not((layer3_outputs(1157)) and (layer3_outputs(899)));
    layer4_outputs(626) <= layer3_outputs(1287);
    layer4_outputs(627) <= (layer3_outputs(141)) or (layer3_outputs(468));
    layer4_outputs(628) <= not(layer3_outputs(1132)) or (layer3_outputs(318));
    layer4_outputs(629) <= not(layer3_outputs(2503));
    layer4_outputs(630) <= layer3_outputs(938);
    layer4_outputs(631) <= (layer3_outputs(1893)) or (layer3_outputs(4436));
    layer4_outputs(632) <= layer3_outputs(4950);
    layer4_outputs(633) <= (layer3_outputs(1271)) and (layer3_outputs(4323));
    layer4_outputs(634) <= (layer3_outputs(2233)) and (layer3_outputs(683));
    layer4_outputs(635) <= (layer3_outputs(3734)) and (layer3_outputs(4374));
    layer4_outputs(636) <= layer3_outputs(1189);
    layer4_outputs(637) <= (layer3_outputs(4342)) and not (layer3_outputs(2850));
    layer4_outputs(638) <= (layer3_outputs(4094)) or (layer3_outputs(2027));
    layer4_outputs(639) <= not(layer3_outputs(705)) or (layer3_outputs(2472));
    layer4_outputs(640) <= not(layer3_outputs(2872));
    layer4_outputs(641) <= not((layer3_outputs(3207)) and (layer3_outputs(1569)));
    layer4_outputs(642) <= not(layer3_outputs(1816)) or (layer3_outputs(3637));
    layer4_outputs(643) <= layer3_outputs(3506);
    layer4_outputs(644) <= not(layer3_outputs(1923)) or (layer3_outputs(2341));
    layer4_outputs(645) <= (layer3_outputs(2783)) and (layer3_outputs(2637));
    layer4_outputs(646) <= '0';
    layer4_outputs(647) <= '0';
    layer4_outputs(648) <= (layer3_outputs(87)) and not (layer3_outputs(5092));
    layer4_outputs(649) <= layer3_outputs(2377);
    layer4_outputs(650) <= layer3_outputs(3224);
    layer4_outputs(651) <= not(layer3_outputs(4459)) or (layer3_outputs(2593));
    layer4_outputs(652) <= not(layer3_outputs(1561));
    layer4_outputs(653) <= not(layer3_outputs(3967)) or (layer3_outputs(1131));
    layer4_outputs(654) <= layer3_outputs(4377);
    layer4_outputs(655) <= not(layer3_outputs(768)) or (layer3_outputs(2081));
    layer4_outputs(656) <= not((layer3_outputs(741)) and (layer3_outputs(4105)));
    layer4_outputs(657) <= not(layer3_outputs(5048)) or (layer3_outputs(1473));
    layer4_outputs(658) <= not((layer3_outputs(4899)) and (layer3_outputs(1053)));
    layer4_outputs(659) <= not((layer3_outputs(3240)) or (layer3_outputs(4579)));
    layer4_outputs(660) <= layer3_outputs(4123);
    layer4_outputs(661) <= layer3_outputs(3091);
    layer4_outputs(662) <= layer3_outputs(1788);
    layer4_outputs(663) <= (layer3_outputs(4482)) and not (layer3_outputs(3960));
    layer4_outputs(664) <= (layer3_outputs(2955)) and not (layer3_outputs(1103));
    layer4_outputs(665) <= not((layer3_outputs(2215)) and (layer3_outputs(1124)));
    layer4_outputs(666) <= not(layer3_outputs(3467)) or (layer3_outputs(3136));
    layer4_outputs(667) <= not(layer3_outputs(2818)) or (layer3_outputs(235));
    layer4_outputs(668) <= not(layer3_outputs(5035)) or (layer3_outputs(170));
    layer4_outputs(669) <= not(layer3_outputs(1192)) or (layer3_outputs(2937));
    layer4_outputs(670) <= (layer3_outputs(2333)) or (layer3_outputs(3057));
    layer4_outputs(671) <= '1';
    layer4_outputs(672) <= not(layer3_outputs(4860)) or (layer3_outputs(967));
    layer4_outputs(673) <= layer3_outputs(4211);
    layer4_outputs(674) <= not(layer3_outputs(3387)) or (layer3_outputs(507));
    layer4_outputs(675) <= not((layer3_outputs(2169)) or (layer3_outputs(3424)));
    layer4_outputs(676) <= not(layer3_outputs(4476)) or (layer3_outputs(3434));
    layer4_outputs(677) <= not(layer3_outputs(2196));
    layer4_outputs(678) <= not((layer3_outputs(3956)) and (layer3_outputs(4351)));
    layer4_outputs(679) <= (layer3_outputs(3224)) and not (layer3_outputs(1144));
    layer4_outputs(680) <= (layer3_outputs(2739)) and (layer3_outputs(2659));
    layer4_outputs(681) <= '1';
    layer4_outputs(682) <= not(layer3_outputs(4670)) or (layer3_outputs(2839));
    layer4_outputs(683) <= (layer3_outputs(274)) and (layer3_outputs(869));
    layer4_outputs(684) <= not((layer3_outputs(604)) and (layer3_outputs(2948)));
    layer4_outputs(685) <= (layer3_outputs(1937)) or (layer3_outputs(298));
    layer4_outputs(686) <= not(layer3_outputs(1897));
    layer4_outputs(687) <= (layer3_outputs(4008)) and (layer3_outputs(742));
    layer4_outputs(688) <= (layer3_outputs(3107)) or (layer3_outputs(1899));
    layer4_outputs(689) <= layer3_outputs(3333);
    layer4_outputs(690) <= (layer3_outputs(4878)) and (layer3_outputs(3022));
    layer4_outputs(691) <= (layer3_outputs(4748)) or (layer3_outputs(4559));
    layer4_outputs(692) <= not(layer3_outputs(4192));
    layer4_outputs(693) <= (layer3_outputs(17)) and (layer3_outputs(4189));
    layer4_outputs(694) <= '0';
    layer4_outputs(695) <= layer3_outputs(1745);
    layer4_outputs(696) <= (layer3_outputs(1541)) and not (layer3_outputs(2292));
    layer4_outputs(697) <= layer3_outputs(2266);
    layer4_outputs(698) <= not(layer3_outputs(622));
    layer4_outputs(699) <= (layer3_outputs(2125)) or (layer3_outputs(4601));
    layer4_outputs(700) <= not(layer3_outputs(2687)) or (layer3_outputs(2760));
    layer4_outputs(701) <= layer3_outputs(2013);
    layer4_outputs(702) <= '1';
    layer4_outputs(703) <= (layer3_outputs(2067)) and (layer3_outputs(3000));
    layer4_outputs(704) <= not(layer3_outputs(4398)) or (layer3_outputs(2392));
    layer4_outputs(705) <= (layer3_outputs(4505)) or (layer3_outputs(3758));
    layer4_outputs(706) <= not((layer3_outputs(5063)) or (layer3_outputs(1559)));
    layer4_outputs(707) <= (layer3_outputs(1419)) and not (layer3_outputs(4025));
    layer4_outputs(708) <= (layer3_outputs(4996)) and not (layer3_outputs(3035));
    layer4_outputs(709) <= not(layer3_outputs(4098));
    layer4_outputs(710) <= not(layer3_outputs(55)) or (layer3_outputs(2617));
    layer4_outputs(711) <= layer3_outputs(42);
    layer4_outputs(712) <= (layer3_outputs(434)) or (layer3_outputs(4804));
    layer4_outputs(713) <= layer3_outputs(4621);
    layer4_outputs(714) <= not(layer3_outputs(876)) or (layer3_outputs(2127));
    layer4_outputs(715) <= not(layer3_outputs(4746)) or (layer3_outputs(1503));
    layer4_outputs(716) <= (layer3_outputs(2624)) or (layer3_outputs(3678));
    layer4_outputs(717) <= not(layer3_outputs(4749));
    layer4_outputs(718) <= layer3_outputs(172);
    layer4_outputs(719) <= not(layer3_outputs(1996));
    layer4_outputs(720) <= not(layer3_outputs(4188));
    layer4_outputs(721) <= layer3_outputs(1351);
    layer4_outputs(722) <= not(layer3_outputs(2423)) or (layer3_outputs(86));
    layer4_outputs(723) <= layer3_outputs(2094);
    layer4_outputs(724) <= (layer3_outputs(829)) and (layer3_outputs(3104));
    layer4_outputs(725) <= not((layer3_outputs(1122)) or (layer3_outputs(3403)));
    layer4_outputs(726) <= '1';
    layer4_outputs(727) <= (layer3_outputs(2160)) and not (layer3_outputs(796));
    layer4_outputs(728) <= (layer3_outputs(1413)) and (layer3_outputs(3407));
    layer4_outputs(729) <= not(layer3_outputs(3167)) or (layer3_outputs(796));
    layer4_outputs(730) <= (layer3_outputs(325)) and (layer3_outputs(2942));
    layer4_outputs(731) <= not((layer3_outputs(1247)) or (layer3_outputs(3766)));
    layer4_outputs(732) <= layer3_outputs(4788);
    layer4_outputs(733) <= layer3_outputs(4250);
    layer4_outputs(734) <= not(layer3_outputs(2442));
    layer4_outputs(735) <= not(layer3_outputs(2737)) or (layer3_outputs(4042));
    layer4_outputs(736) <= layer3_outputs(5084);
    layer4_outputs(737) <= '1';
    layer4_outputs(738) <= (layer3_outputs(1386)) and not (layer3_outputs(1179));
    layer4_outputs(739) <= layer3_outputs(2838);
    layer4_outputs(740) <= not((layer3_outputs(4591)) xor (layer3_outputs(3512)));
    layer4_outputs(741) <= not(layer3_outputs(3708));
    layer4_outputs(742) <= not(layer3_outputs(2056)) or (layer3_outputs(4401));
    layer4_outputs(743) <= not(layer3_outputs(4807));
    layer4_outputs(744) <= layer3_outputs(2052);
    layer4_outputs(745) <= layer3_outputs(2439);
    layer4_outputs(746) <= (layer3_outputs(121)) and not (layer3_outputs(426));
    layer4_outputs(747) <= (layer3_outputs(3725)) and not (layer3_outputs(3376));
    layer4_outputs(748) <= (layer3_outputs(3476)) and not (layer3_outputs(4352));
    layer4_outputs(749) <= not((layer3_outputs(4406)) or (layer3_outputs(1664)));
    layer4_outputs(750) <= not((layer3_outputs(1585)) and (layer3_outputs(27)));
    layer4_outputs(751) <= not((layer3_outputs(163)) and (layer3_outputs(4594)));
    layer4_outputs(752) <= not((layer3_outputs(1500)) xor (layer3_outputs(4299)));
    layer4_outputs(753) <= not((layer3_outputs(3963)) or (layer3_outputs(706)));
    layer4_outputs(754) <= (layer3_outputs(3528)) or (layer3_outputs(2836));
    layer4_outputs(755) <= '0';
    layer4_outputs(756) <= not(layer3_outputs(2348)) or (layer3_outputs(1032));
    layer4_outputs(757) <= layer3_outputs(4001);
    layer4_outputs(758) <= not(layer3_outputs(2033));
    layer4_outputs(759) <= not(layer3_outputs(4700));
    layer4_outputs(760) <= not(layer3_outputs(1436)) or (layer3_outputs(3357));
    layer4_outputs(761) <= not((layer3_outputs(4364)) or (layer3_outputs(2791)));
    layer4_outputs(762) <= (layer3_outputs(3360)) and not (layer3_outputs(4471));
    layer4_outputs(763) <= layer3_outputs(2467);
    layer4_outputs(764) <= (layer3_outputs(4652)) or (layer3_outputs(3583));
    layer4_outputs(765) <= not(layer3_outputs(4761)) or (layer3_outputs(4106));
    layer4_outputs(766) <= not(layer3_outputs(4969));
    layer4_outputs(767) <= not(layer3_outputs(3181)) or (layer3_outputs(2448));
    layer4_outputs(768) <= (layer3_outputs(923)) and not (layer3_outputs(2646));
    layer4_outputs(769) <= not(layer3_outputs(2150)) or (layer3_outputs(2861));
    layer4_outputs(770) <= not(layer3_outputs(3194));
    layer4_outputs(771) <= not(layer3_outputs(844));
    layer4_outputs(772) <= '0';
    layer4_outputs(773) <= not(layer3_outputs(3595)) or (layer3_outputs(664));
    layer4_outputs(774) <= not((layer3_outputs(5046)) or (layer3_outputs(4132)));
    layer4_outputs(775) <= (layer3_outputs(5035)) and (layer3_outputs(374));
    layer4_outputs(776) <= layer3_outputs(355);
    layer4_outputs(777) <= not(layer3_outputs(2003));
    layer4_outputs(778) <= layer3_outputs(5069);
    layer4_outputs(779) <= (layer3_outputs(4483)) and not (layer3_outputs(3964));
    layer4_outputs(780) <= '1';
    layer4_outputs(781) <= not(layer3_outputs(1068));
    layer4_outputs(782) <= layer3_outputs(2777);
    layer4_outputs(783) <= '1';
    layer4_outputs(784) <= (layer3_outputs(2205)) and (layer3_outputs(5111));
    layer4_outputs(785) <= '1';
    layer4_outputs(786) <= layer3_outputs(2191);
    layer4_outputs(787) <= layer3_outputs(4643);
    layer4_outputs(788) <= (layer3_outputs(2905)) and (layer3_outputs(4177));
    layer4_outputs(789) <= (layer3_outputs(1432)) or (layer3_outputs(3756));
    layer4_outputs(790) <= not(layer3_outputs(0));
    layer4_outputs(791) <= not((layer3_outputs(1551)) and (layer3_outputs(2650)));
    layer4_outputs(792) <= not((layer3_outputs(2927)) and (layer3_outputs(1960)));
    layer4_outputs(793) <= not(layer3_outputs(2528)) or (layer3_outputs(2322));
    layer4_outputs(794) <= layer3_outputs(3618);
    layer4_outputs(795) <= not((layer3_outputs(4383)) or (layer3_outputs(4144)));
    layer4_outputs(796) <= not((layer3_outputs(4086)) or (layer3_outputs(782)));
    layer4_outputs(797) <= not((layer3_outputs(3631)) or (layer3_outputs(4949)));
    layer4_outputs(798) <= (layer3_outputs(4315)) and (layer3_outputs(327));
    layer4_outputs(799) <= not((layer3_outputs(2124)) and (layer3_outputs(5053)));
    layer4_outputs(800) <= (layer3_outputs(3629)) or (layer3_outputs(2795));
    layer4_outputs(801) <= not(layer3_outputs(4332)) or (layer3_outputs(713));
    layer4_outputs(802) <= layer3_outputs(1937);
    layer4_outputs(803) <= (layer3_outputs(4924)) or (layer3_outputs(21));
    layer4_outputs(804) <= '1';
    layer4_outputs(805) <= (layer3_outputs(2686)) and (layer3_outputs(2022));
    layer4_outputs(806) <= (layer3_outputs(1272)) and (layer3_outputs(1452));
    layer4_outputs(807) <= not(layer3_outputs(1222));
    layer4_outputs(808) <= (layer3_outputs(2635)) and not (layer3_outputs(3862));
    layer4_outputs(809) <= layer3_outputs(347);
    layer4_outputs(810) <= (layer3_outputs(5018)) and not (layer3_outputs(640));
    layer4_outputs(811) <= layer3_outputs(4763);
    layer4_outputs(812) <= not((layer3_outputs(925)) and (layer3_outputs(1879)));
    layer4_outputs(813) <= '0';
    layer4_outputs(814) <= not(layer3_outputs(1082));
    layer4_outputs(815) <= (layer3_outputs(3898)) and (layer3_outputs(3780));
    layer4_outputs(816) <= not(layer3_outputs(1865));
    layer4_outputs(817) <= '1';
    layer4_outputs(818) <= not(layer3_outputs(3021)) or (layer3_outputs(3632));
    layer4_outputs(819) <= not((layer3_outputs(2087)) or (layer3_outputs(1466)));
    layer4_outputs(820) <= (layer3_outputs(215)) and (layer3_outputs(2364));
    layer4_outputs(821) <= (layer3_outputs(3997)) and not (layer3_outputs(4475));
    layer4_outputs(822) <= (layer3_outputs(4104)) or (layer3_outputs(349));
    layer4_outputs(823) <= not((layer3_outputs(449)) or (layer3_outputs(1171)));
    layer4_outputs(824) <= not(layer3_outputs(4937)) or (layer3_outputs(4797));
    layer4_outputs(825) <= (layer3_outputs(3750)) and (layer3_outputs(2238));
    layer4_outputs(826) <= not(layer3_outputs(3568));
    layer4_outputs(827) <= '1';
    layer4_outputs(828) <= not(layer3_outputs(4007));
    layer4_outputs(829) <= (layer3_outputs(4053)) and (layer3_outputs(381));
    layer4_outputs(830) <= (layer3_outputs(941)) and not (layer3_outputs(90));
    layer4_outputs(831) <= (layer3_outputs(2944)) or (layer3_outputs(4062));
    layer4_outputs(832) <= (layer3_outputs(3611)) or (layer3_outputs(3159));
    layer4_outputs(833) <= not((layer3_outputs(1939)) and (layer3_outputs(2255)));
    layer4_outputs(834) <= not((layer3_outputs(4210)) and (layer3_outputs(651)));
    layer4_outputs(835) <= (layer3_outputs(4601)) and not (layer3_outputs(1776));
    layer4_outputs(836) <= not((layer3_outputs(4368)) and (layer3_outputs(2466)));
    layer4_outputs(837) <= not(layer3_outputs(4257)) or (layer3_outputs(4832));
    layer4_outputs(838) <= layer3_outputs(3971);
    layer4_outputs(839) <= (layer3_outputs(1667)) or (layer3_outputs(3469));
    layer4_outputs(840) <= not(layer3_outputs(1391)) or (layer3_outputs(823));
    layer4_outputs(841) <= not(layer3_outputs(1560)) or (layer3_outputs(5025));
    layer4_outputs(842) <= not(layer3_outputs(4433));
    layer4_outputs(843) <= not((layer3_outputs(1173)) and (layer3_outputs(4655)));
    layer4_outputs(844) <= layer3_outputs(354);
    layer4_outputs(845) <= not(layer3_outputs(4184)) or (layer3_outputs(512));
    layer4_outputs(846) <= (layer3_outputs(14)) and not (layer3_outputs(1367));
    layer4_outputs(847) <= '1';
    layer4_outputs(848) <= (layer3_outputs(4558)) and not (layer3_outputs(4275));
    layer4_outputs(849) <= not(layer3_outputs(3115));
    layer4_outputs(850) <= not((layer3_outputs(4239)) or (layer3_outputs(3542)));
    layer4_outputs(851) <= (layer3_outputs(4874)) and (layer3_outputs(1841));
    layer4_outputs(852) <= (layer3_outputs(1896)) and (layer3_outputs(3509));
    layer4_outputs(853) <= not(layer3_outputs(4932));
    layer4_outputs(854) <= not(layer3_outputs(300));
    layer4_outputs(855) <= layer3_outputs(2750);
    layer4_outputs(856) <= (layer3_outputs(725)) and (layer3_outputs(901));
    layer4_outputs(857) <= (layer3_outputs(316)) xor (layer3_outputs(184));
    layer4_outputs(858) <= not((layer3_outputs(821)) and (layer3_outputs(353)));
    layer4_outputs(859) <= not(layer3_outputs(4115)) or (layer3_outputs(1970));
    layer4_outputs(860) <= (layer3_outputs(2880)) or (layer3_outputs(4106));
    layer4_outputs(861) <= not(layer3_outputs(4483)) or (layer3_outputs(3202));
    layer4_outputs(862) <= '1';
    layer4_outputs(863) <= (layer3_outputs(625)) or (layer3_outputs(841));
    layer4_outputs(864) <= layer3_outputs(2858);
    layer4_outputs(865) <= not(layer3_outputs(2625)) or (layer3_outputs(994));
    layer4_outputs(866) <= (layer3_outputs(2816)) or (layer3_outputs(805));
    layer4_outputs(867) <= not((layer3_outputs(1017)) or (layer3_outputs(1940)));
    layer4_outputs(868) <= not(layer3_outputs(1812)) or (layer3_outputs(3430));
    layer4_outputs(869) <= layer3_outputs(2416);
    layer4_outputs(870) <= (layer3_outputs(4551)) and not (layer3_outputs(1780));
    layer4_outputs(871) <= not((layer3_outputs(2662)) or (layer3_outputs(3455)));
    layer4_outputs(872) <= not(layer3_outputs(425));
    layer4_outputs(873) <= not(layer3_outputs(1742)) or (layer3_outputs(5079));
    layer4_outputs(874) <= layer3_outputs(2726);
    layer4_outputs(875) <= '0';
    layer4_outputs(876) <= not(layer3_outputs(3370)) or (layer3_outputs(2017));
    layer4_outputs(877) <= (layer3_outputs(3949)) and not (layer3_outputs(2470));
    layer4_outputs(878) <= not((layer3_outputs(1369)) or (layer3_outputs(4857)));
    layer4_outputs(879) <= not(layer3_outputs(2628)) or (layer3_outputs(1545));
    layer4_outputs(880) <= layer3_outputs(4086);
    layer4_outputs(881) <= layer3_outputs(4919);
    layer4_outputs(882) <= not(layer3_outputs(3144)) or (layer3_outputs(4358));
    layer4_outputs(883) <= layer3_outputs(4355);
    layer4_outputs(884) <= not(layer3_outputs(769)) or (layer3_outputs(1389));
    layer4_outputs(885) <= layer3_outputs(3552);
    layer4_outputs(886) <= (layer3_outputs(2842)) or (layer3_outputs(4913));
    layer4_outputs(887) <= '1';
    layer4_outputs(888) <= not(layer3_outputs(1889)) or (layer3_outputs(4447));
    layer4_outputs(889) <= not(layer3_outputs(2745));
    layer4_outputs(890) <= layer3_outputs(4102);
    layer4_outputs(891) <= (layer3_outputs(1987)) and not (layer3_outputs(1443));
    layer4_outputs(892) <= not(layer3_outputs(2058)) or (layer3_outputs(3627));
    layer4_outputs(893) <= not(layer3_outputs(3104)) or (layer3_outputs(4602));
    layer4_outputs(894) <= '1';
    layer4_outputs(895) <= not(layer3_outputs(2438));
    layer4_outputs(896) <= '1';
    layer4_outputs(897) <= not((layer3_outputs(1213)) and (layer3_outputs(1826)));
    layer4_outputs(898) <= layer3_outputs(4511);
    layer4_outputs(899) <= (layer3_outputs(1992)) and (layer3_outputs(1682));
    layer4_outputs(900) <= not(layer3_outputs(2678)) or (layer3_outputs(2601));
    layer4_outputs(901) <= layer3_outputs(1133);
    layer4_outputs(902) <= (layer3_outputs(1637)) or (layer3_outputs(199));
    layer4_outputs(903) <= not(layer3_outputs(1692));
    layer4_outputs(904) <= '1';
    layer4_outputs(905) <= (layer3_outputs(2735)) or (layer3_outputs(4799));
    layer4_outputs(906) <= not(layer3_outputs(3534));
    layer4_outputs(907) <= (layer3_outputs(3731)) or (layer3_outputs(4058));
    layer4_outputs(908) <= layer3_outputs(924);
    layer4_outputs(909) <= (layer3_outputs(1019)) and (layer3_outputs(3391));
    layer4_outputs(910) <= not(layer3_outputs(1919));
    layer4_outputs(911) <= not((layer3_outputs(1699)) or (layer3_outputs(4627)));
    layer4_outputs(912) <= not(layer3_outputs(1046)) or (layer3_outputs(921));
    layer4_outputs(913) <= not((layer3_outputs(417)) and (layer3_outputs(4030)));
    layer4_outputs(914) <= (layer3_outputs(4924)) and not (layer3_outputs(88));
    layer4_outputs(915) <= not(layer3_outputs(3952)) or (layer3_outputs(216));
    layer4_outputs(916) <= not(layer3_outputs(377));
    layer4_outputs(917) <= not((layer3_outputs(4659)) and (layer3_outputs(1820)));
    layer4_outputs(918) <= (layer3_outputs(3216)) xor (layer3_outputs(1146));
    layer4_outputs(919) <= '0';
    layer4_outputs(920) <= (layer3_outputs(1691)) or (layer3_outputs(1917));
    layer4_outputs(921) <= layer3_outputs(4818);
    layer4_outputs(922) <= not(layer3_outputs(401)) or (layer3_outputs(3209));
    layer4_outputs(923) <= (layer3_outputs(54)) and (layer3_outputs(2752));
    layer4_outputs(924) <= layer3_outputs(4270);
    layer4_outputs(925) <= (layer3_outputs(4095)) and (layer3_outputs(1697));
    layer4_outputs(926) <= '1';
    layer4_outputs(927) <= not(layer3_outputs(3978));
    layer4_outputs(928) <= not(layer3_outputs(596));
    layer4_outputs(929) <= not((layer3_outputs(4598)) or (layer3_outputs(3316)));
    layer4_outputs(930) <= layer3_outputs(1962);
    layer4_outputs(931) <= not((layer3_outputs(3465)) and (layer3_outputs(846)));
    layer4_outputs(932) <= not(layer3_outputs(728)) or (layer3_outputs(3043));
    layer4_outputs(933) <= (layer3_outputs(3561)) or (layer3_outputs(3657));
    layer4_outputs(934) <= layer3_outputs(4054);
    layer4_outputs(935) <= not(layer3_outputs(4901)) or (layer3_outputs(4293));
    layer4_outputs(936) <= layer3_outputs(4271);
    layer4_outputs(937) <= not(layer3_outputs(3397));
    layer4_outputs(938) <= layer3_outputs(82);
    layer4_outputs(939) <= not((layer3_outputs(1611)) and (layer3_outputs(2268)));
    layer4_outputs(940) <= (layer3_outputs(2721)) or (layer3_outputs(4237));
    layer4_outputs(941) <= '1';
    layer4_outputs(942) <= (layer3_outputs(2568)) and (layer3_outputs(2959));
    layer4_outputs(943) <= not(layer3_outputs(4205));
    layer4_outputs(944) <= not((layer3_outputs(181)) or (layer3_outputs(976)));
    layer4_outputs(945) <= not((layer3_outputs(3145)) xor (layer3_outputs(4929)));
    layer4_outputs(946) <= not(layer3_outputs(673));
    layer4_outputs(947) <= (layer3_outputs(3371)) or (layer3_outputs(669));
    layer4_outputs(948) <= (layer3_outputs(2589)) and (layer3_outputs(252));
    layer4_outputs(949) <= '0';
    layer4_outputs(950) <= '1';
    layer4_outputs(951) <= (layer3_outputs(1010)) and (layer3_outputs(772));
    layer4_outputs(952) <= (layer3_outputs(3874)) and not (layer3_outputs(3604));
    layer4_outputs(953) <= (layer3_outputs(479)) and not (layer3_outputs(2798));
    layer4_outputs(954) <= not((layer3_outputs(4103)) and (layer3_outputs(2247)));
    layer4_outputs(955) <= not(layer3_outputs(1907)) or (layer3_outputs(3440));
    layer4_outputs(956) <= not((layer3_outputs(697)) or (layer3_outputs(4994)));
    layer4_outputs(957) <= (layer3_outputs(4701)) and (layer3_outputs(3366));
    layer4_outputs(958) <= not(layer3_outputs(2600)) or (layer3_outputs(2817));
    layer4_outputs(959) <= '0';
    layer4_outputs(960) <= not((layer3_outputs(3139)) and (layer3_outputs(177)));
    layer4_outputs(961) <= layer3_outputs(1427);
    layer4_outputs(962) <= not(layer3_outputs(71)) or (layer3_outputs(2894));
    layer4_outputs(963) <= layer3_outputs(2411);
    layer4_outputs(964) <= not(layer3_outputs(4574)) or (layer3_outputs(3623));
    layer4_outputs(965) <= not((layer3_outputs(411)) xor (layer3_outputs(4276)));
    layer4_outputs(966) <= not(layer3_outputs(2197));
    layer4_outputs(967) <= not((layer3_outputs(1751)) or (layer3_outputs(5021)));
    layer4_outputs(968) <= (layer3_outputs(4900)) and not (layer3_outputs(1641));
    layer4_outputs(969) <= not((layer3_outputs(1724)) or (layer3_outputs(2985)));
    layer4_outputs(970) <= layer3_outputs(3846);
    layer4_outputs(971) <= (layer3_outputs(375)) and (layer3_outputs(1938));
    layer4_outputs(972) <= not(layer3_outputs(629));
    layer4_outputs(973) <= (layer3_outputs(3471)) or (layer3_outputs(4613));
    layer4_outputs(974) <= (layer3_outputs(4904)) and not (layer3_outputs(1961));
    layer4_outputs(975) <= '1';
    layer4_outputs(976) <= not(layer3_outputs(4376)) or (layer3_outputs(1224));
    layer4_outputs(977) <= '1';
    layer4_outputs(978) <= layer3_outputs(3081);
    layer4_outputs(979) <= (layer3_outputs(2302)) xor (layer3_outputs(4581));
    layer4_outputs(980) <= '1';
    layer4_outputs(981) <= not((layer3_outputs(3015)) xor (layer3_outputs(1212)));
    layer4_outputs(982) <= (layer3_outputs(2261)) and not (layer3_outputs(2188));
    layer4_outputs(983) <= (layer3_outputs(3667)) and (layer3_outputs(4939));
    layer4_outputs(984) <= '0';
    layer4_outputs(985) <= (layer3_outputs(2286)) and not (layer3_outputs(1887));
    layer4_outputs(986) <= '0';
    layer4_outputs(987) <= not(layer3_outputs(259));
    layer4_outputs(988) <= not(layer3_outputs(1919)) or (layer3_outputs(3313));
    layer4_outputs(989) <= (layer3_outputs(4364)) or (layer3_outputs(3326));
    layer4_outputs(990) <= '0';
    layer4_outputs(991) <= '1';
    layer4_outputs(992) <= '1';
    layer4_outputs(993) <= '0';
    layer4_outputs(994) <= not(layer3_outputs(4509));
    layer4_outputs(995) <= not((layer3_outputs(2790)) or (layer3_outputs(3129)));
    layer4_outputs(996) <= not(layer3_outputs(2408));
    layer4_outputs(997) <= layer3_outputs(4443);
    layer4_outputs(998) <= (layer3_outputs(188)) or (layer3_outputs(2014));
    layer4_outputs(999) <= '0';
    layer4_outputs(1000) <= (layer3_outputs(2184)) and not (layer3_outputs(4294));
    layer4_outputs(1001) <= (layer3_outputs(4751)) xor (layer3_outputs(1354));
    layer4_outputs(1002) <= not((layer3_outputs(2531)) and (layer3_outputs(5110)));
    layer4_outputs(1003) <= '0';
    layer4_outputs(1004) <= not(layer3_outputs(759));
    layer4_outputs(1005) <= '0';
    layer4_outputs(1006) <= not(layer3_outputs(4457)) or (layer3_outputs(3117));
    layer4_outputs(1007) <= not(layer3_outputs(2747)) or (layer3_outputs(2278));
    layer4_outputs(1008) <= not((layer3_outputs(1236)) and (layer3_outputs(2221)));
    layer4_outputs(1009) <= not(layer3_outputs(3091)) or (layer3_outputs(1661));
    layer4_outputs(1010) <= not((layer3_outputs(3446)) and (layer3_outputs(1663)));
    layer4_outputs(1011) <= not(layer3_outputs(3198));
    layer4_outputs(1012) <= layer3_outputs(3618);
    layer4_outputs(1013) <= '1';
    layer4_outputs(1014) <= not((layer3_outputs(2673)) xor (layer3_outputs(1954)));
    layer4_outputs(1015) <= '1';
    layer4_outputs(1016) <= (layer3_outputs(1118)) and not (layer3_outputs(4140));
    layer4_outputs(1017) <= not(layer3_outputs(4043));
    layer4_outputs(1018) <= not((layer3_outputs(3590)) and (layer3_outputs(221)));
    layer4_outputs(1019) <= not(layer3_outputs(2812));
    layer4_outputs(1020) <= (layer3_outputs(15)) and not (layer3_outputs(3391));
    layer4_outputs(1021) <= not(layer3_outputs(3330));
    layer4_outputs(1022) <= (layer3_outputs(343)) and (layer3_outputs(3232));
    layer4_outputs(1023) <= '1';
    layer4_outputs(1024) <= not(layer3_outputs(2342));
    layer4_outputs(1025) <= '1';
    layer4_outputs(1026) <= not((layer3_outputs(2348)) and (layer3_outputs(4190)));
    layer4_outputs(1027) <= (layer3_outputs(2776)) xor (layer3_outputs(2639));
    layer4_outputs(1028) <= (layer3_outputs(302)) and not (layer3_outputs(838));
    layer4_outputs(1029) <= not((layer3_outputs(1325)) xor (layer3_outputs(5015)));
    layer4_outputs(1030) <= layer3_outputs(94);
    layer4_outputs(1031) <= not(layer3_outputs(2618));
    layer4_outputs(1032) <= (layer3_outputs(4276)) and not (layer3_outputs(353));
    layer4_outputs(1033) <= not((layer3_outputs(761)) and (layer3_outputs(4331)));
    layer4_outputs(1034) <= '1';
    layer4_outputs(1035) <= not(layer3_outputs(1343));
    layer4_outputs(1036) <= not(layer3_outputs(3871)) or (layer3_outputs(3838));
    layer4_outputs(1037) <= not((layer3_outputs(4641)) xor (layer3_outputs(4127)));
    layer4_outputs(1038) <= not((layer3_outputs(725)) and (layer3_outputs(1699)));
    layer4_outputs(1039) <= not((layer3_outputs(3311)) and (layer3_outputs(3093)));
    layer4_outputs(1040) <= (layer3_outputs(952)) and not (layer3_outputs(3869));
    layer4_outputs(1041) <= not((layer3_outputs(4440)) xor (layer3_outputs(653)));
    layer4_outputs(1042) <= not(layer3_outputs(2845)) or (layer3_outputs(3576));
    layer4_outputs(1043) <= not(layer3_outputs(1401));
    layer4_outputs(1044) <= (layer3_outputs(4158)) and not (layer3_outputs(4386));
    layer4_outputs(1045) <= not(layer3_outputs(4589));
    layer4_outputs(1046) <= not((layer3_outputs(966)) and (layer3_outputs(3013)));
    layer4_outputs(1047) <= not(layer3_outputs(4081)) or (layer3_outputs(566));
    layer4_outputs(1048) <= not((layer3_outputs(3671)) xor (layer3_outputs(1195)));
    layer4_outputs(1049) <= not(layer3_outputs(4335)) or (layer3_outputs(4549));
    layer4_outputs(1050) <= not(layer3_outputs(1749));
    layer4_outputs(1051) <= (layer3_outputs(4687)) or (layer3_outputs(1370));
    layer4_outputs(1052) <= not((layer3_outputs(133)) or (layer3_outputs(3894)));
    layer4_outputs(1053) <= not((layer3_outputs(2072)) xor (layer3_outputs(4292)));
    layer4_outputs(1054) <= (layer3_outputs(3585)) and not (layer3_outputs(169));
    layer4_outputs(1055) <= not(layer3_outputs(4820)) or (layer3_outputs(2223));
    layer4_outputs(1056) <= '1';
    layer4_outputs(1057) <= '0';
    layer4_outputs(1058) <= (layer3_outputs(4461)) and not (layer3_outputs(357));
    layer4_outputs(1059) <= layer3_outputs(4248);
    layer4_outputs(1060) <= not((layer3_outputs(1716)) and (layer3_outputs(2076)));
    layer4_outputs(1061) <= '1';
    layer4_outputs(1062) <= (layer3_outputs(1380)) or (layer3_outputs(2000));
    layer4_outputs(1063) <= not(layer3_outputs(3877));
    layer4_outputs(1064) <= (layer3_outputs(4495)) and (layer3_outputs(1200));
    layer4_outputs(1065) <= not(layer3_outputs(511)) or (layer3_outputs(384));
    layer4_outputs(1066) <= not(layer3_outputs(2163));
    layer4_outputs(1067) <= '1';
    layer4_outputs(1068) <= '0';
    layer4_outputs(1069) <= not(layer3_outputs(4240));
    layer4_outputs(1070) <= not(layer3_outputs(1105)) or (layer3_outputs(3599));
    layer4_outputs(1071) <= '1';
    layer4_outputs(1072) <= (layer3_outputs(2843)) or (layer3_outputs(3609));
    layer4_outputs(1073) <= layer3_outputs(2312);
    layer4_outputs(1074) <= (layer3_outputs(2999)) and (layer3_outputs(1051));
    layer4_outputs(1075) <= not(layer3_outputs(2006));
    layer4_outputs(1076) <= not((layer3_outputs(4706)) and (layer3_outputs(3006)));
    layer4_outputs(1077) <= not(layer3_outputs(3760)) or (layer3_outputs(5087));
    layer4_outputs(1078) <= (layer3_outputs(3582)) and not (layer3_outputs(4395));
    layer4_outputs(1079) <= (layer3_outputs(903)) and (layer3_outputs(2844));
    layer4_outputs(1080) <= (layer3_outputs(4622)) and (layer3_outputs(4076));
    layer4_outputs(1081) <= not(layer3_outputs(1204));
    layer4_outputs(1082) <= not(layer3_outputs(4756));
    layer4_outputs(1083) <= layer3_outputs(3908);
    layer4_outputs(1084) <= layer3_outputs(1211);
    layer4_outputs(1085) <= not(layer3_outputs(2912));
    layer4_outputs(1086) <= layer3_outputs(2212);
    layer4_outputs(1087) <= (layer3_outputs(1851)) and not (layer3_outputs(3055));
    layer4_outputs(1088) <= not(layer3_outputs(4876));
    layer4_outputs(1089) <= not((layer3_outputs(573)) or (layer3_outputs(4343)));
    layer4_outputs(1090) <= (layer3_outputs(2247)) xor (layer3_outputs(2489));
    layer4_outputs(1091) <= (layer3_outputs(2352)) and not (layer3_outputs(2204));
    layer4_outputs(1092) <= (layer3_outputs(1957)) or (layer3_outputs(3701));
    layer4_outputs(1093) <= layer3_outputs(3199);
    layer4_outputs(1094) <= layer3_outputs(764);
    layer4_outputs(1095) <= not((layer3_outputs(408)) and (layer3_outputs(2545)));
    layer4_outputs(1096) <= layer3_outputs(648);
    layer4_outputs(1097) <= (layer3_outputs(2752)) and not (layer3_outputs(5007));
    layer4_outputs(1098) <= not((layer3_outputs(4721)) and (layer3_outputs(1899)));
    layer4_outputs(1099) <= '1';
    layer4_outputs(1100) <= not(layer3_outputs(2584)) or (layer3_outputs(261));
    layer4_outputs(1101) <= not(layer3_outputs(2908)) or (layer3_outputs(371));
    layer4_outputs(1102) <= not(layer3_outputs(1945));
    layer4_outputs(1103) <= (layer3_outputs(5061)) and not (layer3_outputs(4650));
    layer4_outputs(1104) <= layer3_outputs(4559);
    layer4_outputs(1105) <= '1';
    layer4_outputs(1106) <= not(layer3_outputs(679));
    layer4_outputs(1107) <= not(layer3_outputs(2973));
    layer4_outputs(1108) <= (layer3_outputs(2013)) or (layer3_outputs(4937));
    layer4_outputs(1109) <= '0';
    layer4_outputs(1110) <= layer3_outputs(2570);
    layer4_outputs(1111) <= not(layer3_outputs(859)) or (layer3_outputs(319));
    layer4_outputs(1112) <= not(layer3_outputs(585)) or (layer3_outputs(199));
    layer4_outputs(1113) <= (layer3_outputs(3932)) and (layer3_outputs(3313));
    layer4_outputs(1114) <= (layer3_outputs(2611)) xor (layer3_outputs(4314));
    layer4_outputs(1115) <= layer3_outputs(1844);
    layer4_outputs(1116) <= (layer3_outputs(2888)) and not (layer3_outputs(4971));
    layer4_outputs(1117) <= not((layer3_outputs(106)) and (layer3_outputs(502)));
    layer4_outputs(1118) <= (layer3_outputs(2931)) or (layer3_outputs(1705));
    layer4_outputs(1119) <= not(layer3_outputs(795));
    layer4_outputs(1120) <= not(layer3_outputs(1398));
    layer4_outputs(1121) <= (layer3_outputs(3105)) and not (layer3_outputs(3249));
    layer4_outputs(1122) <= not((layer3_outputs(2305)) or (layer3_outputs(4221)));
    layer4_outputs(1123) <= layer3_outputs(4329);
    layer4_outputs(1124) <= '0';
    layer4_outputs(1125) <= layer3_outputs(800);
    layer4_outputs(1126) <= not(layer3_outputs(2391));
    layer4_outputs(1127) <= not((layer3_outputs(2909)) or (layer3_outputs(675)));
    layer4_outputs(1128) <= layer3_outputs(415);
    layer4_outputs(1129) <= (layer3_outputs(3870)) and not (layer3_outputs(4137));
    layer4_outputs(1130) <= not(layer3_outputs(379));
    layer4_outputs(1131) <= (layer3_outputs(2514)) and not (layer3_outputs(2524));
    layer4_outputs(1132) <= not((layer3_outputs(566)) and (layer3_outputs(3397)));
    layer4_outputs(1133) <= '0';
    layer4_outputs(1134) <= not(layer3_outputs(2523)) or (layer3_outputs(3831));
    layer4_outputs(1135) <= not(layer3_outputs(173)) or (layer3_outputs(4894));
    layer4_outputs(1136) <= not(layer3_outputs(2612));
    layer4_outputs(1137) <= not(layer3_outputs(1768));
    layer4_outputs(1138) <= (layer3_outputs(4699)) and not (layer3_outputs(4635));
    layer4_outputs(1139) <= layer3_outputs(2295);
    layer4_outputs(1140) <= not(layer3_outputs(4274));
    layer4_outputs(1141) <= '0';
    layer4_outputs(1142) <= (layer3_outputs(4638)) or (layer3_outputs(2228));
    layer4_outputs(1143) <= not(layer3_outputs(143));
    layer4_outputs(1144) <= not(layer3_outputs(4813));
    layer4_outputs(1145) <= (layer3_outputs(735)) and not (layer3_outputs(2565));
    layer4_outputs(1146) <= '1';
    layer4_outputs(1147) <= not(layer3_outputs(4552));
    layer4_outputs(1148) <= not((layer3_outputs(1839)) and (layer3_outputs(4243)));
    layer4_outputs(1149) <= (layer3_outputs(2548)) and (layer3_outputs(473));
    layer4_outputs(1150) <= (layer3_outputs(436)) and (layer3_outputs(3231));
    layer4_outputs(1151) <= not(layer3_outputs(1396));
    layer4_outputs(1152) <= not(layer3_outputs(4844)) or (layer3_outputs(2779));
    layer4_outputs(1153) <= not(layer3_outputs(1340));
    layer4_outputs(1154) <= layer3_outputs(4958);
    layer4_outputs(1155) <= not((layer3_outputs(4612)) or (layer3_outputs(190)));
    layer4_outputs(1156) <= layer3_outputs(2211);
    layer4_outputs(1157) <= not((layer3_outputs(4713)) or (layer3_outputs(3783)));
    layer4_outputs(1158) <= layer3_outputs(1716);
    layer4_outputs(1159) <= not((layer3_outputs(1659)) and (layer3_outputs(2935)));
    layer4_outputs(1160) <= not(layer3_outputs(2543)) or (layer3_outputs(1449));
    layer4_outputs(1161) <= (layer3_outputs(2449)) and not (layer3_outputs(4745));
    layer4_outputs(1162) <= layer3_outputs(511);
    layer4_outputs(1163) <= not(layer3_outputs(3958));
    layer4_outputs(1164) <= '1';
    layer4_outputs(1165) <= not((layer3_outputs(1251)) and (layer3_outputs(3987)));
    layer4_outputs(1166) <= (layer3_outputs(5026)) and (layer3_outputs(4321));
    layer4_outputs(1167) <= not(layer3_outputs(1207)) or (layer3_outputs(1100));
    layer4_outputs(1168) <= (layer3_outputs(3483)) and (layer3_outputs(3441));
    layer4_outputs(1169) <= not((layer3_outputs(51)) or (layer3_outputs(2777)));
    layer4_outputs(1170) <= not((layer3_outputs(2130)) and (layer3_outputs(2589)));
    layer4_outputs(1171) <= (layer3_outputs(646)) and (layer3_outputs(2452));
    layer4_outputs(1172) <= not((layer3_outputs(2637)) and (layer3_outputs(3916)));
    layer4_outputs(1173) <= '0';
    layer4_outputs(1174) <= not(layer3_outputs(1143));
    layer4_outputs(1175) <= '1';
    layer4_outputs(1176) <= (layer3_outputs(3467)) and (layer3_outputs(2753));
    layer4_outputs(1177) <= (layer3_outputs(509)) or (layer3_outputs(550));
    layer4_outputs(1178) <= not(layer3_outputs(4575));
    layer4_outputs(1179) <= not(layer3_outputs(165)) or (layer3_outputs(2606));
    layer4_outputs(1180) <= layer3_outputs(4417);
    layer4_outputs(1181) <= (layer3_outputs(3924)) and not (layer3_outputs(3131));
    layer4_outputs(1182) <= (layer3_outputs(4204)) and (layer3_outputs(1462));
    layer4_outputs(1183) <= not(layer3_outputs(4938)) or (layer3_outputs(3621));
    layer4_outputs(1184) <= not(layer3_outputs(1526)) or (layer3_outputs(3891));
    layer4_outputs(1185) <= not(layer3_outputs(3102));
    layer4_outputs(1186) <= not((layer3_outputs(2401)) and (layer3_outputs(132)));
    layer4_outputs(1187) <= (layer3_outputs(2351)) and not (layer3_outputs(2864));
    layer4_outputs(1188) <= not(layer3_outputs(2340));
    layer4_outputs(1189) <= not(layer3_outputs(2804));
    layer4_outputs(1190) <= (layer3_outputs(2609)) and not (layer3_outputs(2904));
    layer4_outputs(1191) <= (layer3_outputs(1654)) and not (layer3_outputs(4146));
    layer4_outputs(1192) <= '1';
    layer4_outputs(1193) <= not(layer3_outputs(1929)) or (layer3_outputs(1869));
    layer4_outputs(1194) <= (layer3_outputs(266)) or (layer3_outputs(541));
    layer4_outputs(1195) <= (layer3_outputs(57)) and not (layer3_outputs(2959));
    layer4_outputs(1196) <= not(layer3_outputs(579));
    layer4_outputs(1197) <= not(layer3_outputs(1713)) or (layer3_outputs(4730));
    layer4_outputs(1198) <= (layer3_outputs(4339)) or (layer3_outputs(2604));
    layer4_outputs(1199) <= not(layer3_outputs(1431));
    layer4_outputs(1200) <= (layer3_outputs(4469)) or (layer3_outputs(323));
    layer4_outputs(1201) <= not(layer3_outputs(831));
    layer4_outputs(1202) <= (layer3_outputs(3545)) or (layer3_outputs(164));
    layer4_outputs(1203) <= layer3_outputs(2483);
    layer4_outputs(1204) <= not((layer3_outputs(3213)) xor (layer3_outputs(1679)));
    layer4_outputs(1205) <= layer3_outputs(1350);
    layer4_outputs(1206) <= (layer3_outputs(3096)) and (layer3_outputs(4162));
    layer4_outputs(1207) <= '0';
    layer4_outputs(1208) <= '1';
    layer4_outputs(1209) <= (layer3_outputs(4889)) and not (layer3_outputs(3417));
    layer4_outputs(1210) <= not(layer3_outputs(2857)) or (layer3_outputs(5037));
    layer4_outputs(1211) <= layer3_outputs(21);
    layer4_outputs(1212) <= not(layer3_outputs(4238)) or (layer3_outputs(3036));
    layer4_outputs(1213) <= '1';
    layer4_outputs(1214) <= '0';
    layer4_outputs(1215) <= '1';
    layer4_outputs(1216) <= layer3_outputs(1586);
    layer4_outputs(1217) <= not((layer3_outputs(3677)) or (layer3_outputs(2692)));
    layer4_outputs(1218) <= not(layer3_outputs(582)) or (layer3_outputs(3859));
    layer4_outputs(1219) <= (layer3_outputs(2172)) and not (layer3_outputs(4538));
    layer4_outputs(1220) <= not(layer3_outputs(3920));
    layer4_outputs(1221) <= not(layer3_outputs(1106));
    layer4_outputs(1222) <= not(layer3_outputs(4415));
    layer4_outputs(1223) <= not((layer3_outputs(630)) or (layer3_outputs(4176)));
    layer4_outputs(1224) <= not(layer3_outputs(2411));
    layer4_outputs(1225) <= (layer3_outputs(205)) and not (layer3_outputs(4900));
    layer4_outputs(1226) <= not(layer3_outputs(3072)) or (layer3_outputs(4186));
    layer4_outputs(1227) <= layer3_outputs(1238);
    layer4_outputs(1228) <= layer3_outputs(4605);
    layer4_outputs(1229) <= layer3_outputs(4739);
    layer4_outputs(1230) <= layer3_outputs(387);
    layer4_outputs(1231) <= '0';
    layer4_outputs(1232) <= not(layer3_outputs(4019));
    layer4_outputs(1233) <= '0';
    layer4_outputs(1234) <= (layer3_outputs(4675)) or (layer3_outputs(1524));
    layer4_outputs(1235) <= (layer3_outputs(4173)) xor (layer3_outputs(945));
    layer4_outputs(1236) <= not(layer3_outputs(1634));
    layer4_outputs(1237) <= layer3_outputs(1671);
    layer4_outputs(1238) <= (layer3_outputs(4100)) and not (layer3_outputs(1711));
    layer4_outputs(1239) <= not(layer3_outputs(4018));
    layer4_outputs(1240) <= not((layer3_outputs(3259)) or (layer3_outputs(4560)));
    layer4_outputs(1241) <= '0';
    layer4_outputs(1242) <= layer3_outputs(3097);
    layer4_outputs(1243) <= not(layer3_outputs(835)) or (layer3_outputs(3593));
    layer4_outputs(1244) <= not(layer3_outputs(3038)) or (layer3_outputs(4805));
    layer4_outputs(1245) <= not((layer3_outputs(3296)) and (layer3_outputs(734)));
    layer4_outputs(1246) <= (layer3_outputs(3039)) and (layer3_outputs(1270));
    layer4_outputs(1247) <= '1';
    layer4_outputs(1248) <= '1';
    layer4_outputs(1249) <= not((layer3_outputs(2004)) and (layer3_outputs(1467)));
    layer4_outputs(1250) <= (layer3_outputs(4219)) or (layer3_outputs(995));
    layer4_outputs(1251) <= not(layer3_outputs(652)) or (layer3_outputs(1316));
    layer4_outputs(1252) <= (layer3_outputs(4880)) and not (layer3_outputs(4424));
    layer4_outputs(1253) <= layer3_outputs(4923);
    layer4_outputs(1254) <= '0';
    layer4_outputs(1255) <= '1';
    layer4_outputs(1256) <= not(layer3_outputs(251)) or (layer3_outputs(4231));
    layer4_outputs(1257) <= (layer3_outputs(2070)) and not (layer3_outputs(1630));
    layer4_outputs(1258) <= (layer3_outputs(4583)) and not (layer3_outputs(1985));
    layer4_outputs(1259) <= layer3_outputs(497);
    layer4_outputs(1260) <= not((layer3_outputs(1466)) and (layer3_outputs(4353)));
    layer4_outputs(1261) <= not((layer3_outputs(4817)) or (layer3_outputs(606)));
    layer4_outputs(1262) <= not(layer3_outputs(4518)) or (layer3_outputs(1190));
    layer4_outputs(1263) <= layer3_outputs(3069);
    layer4_outputs(1264) <= layer3_outputs(1220);
    layer4_outputs(1265) <= not(layer3_outputs(3815));
    layer4_outputs(1266) <= not((layer3_outputs(4910)) and (layer3_outputs(3742)));
    layer4_outputs(1267) <= (layer3_outputs(722)) and not (layer3_outputs(2876));
    layer4_outputs(1268) <= (layer3_outputs(1961)) or (layer3_outputs(50));
    layer4_outputs(1269) <= not(layer3_outputs(3066)) or (layer3_outputs(3468));
    layer4_outputs(1270) <= layer3_outputs(3972);
    layer4_outputs(1271) <= '0';
    layer4_outputs(1272) <= (layer3_outputs(1927)) xor (layer3_outputs(2607));
    layer4_outputs(1273) <= (layer3_outputs(1966)) or (layer3_outputs(3660));
    layer4_outputs(1274) <= not((layer3_outputs(1021)) and (layer3_outputs(478)));
    layer4_outputs(1275) <= not((layer3_outputs(3064)) or (layer3_outputs(2079)));
    layer4_outputs(1276) <= '0';
    layer4_outputs(1277) <= layer3_outputs(1588);
    layer4_outputs(1278) <= '0';
    layer4_outputs(1279) <= layer3_outputs(4214);
    layer4_outputs(1280) <= '0';
    layer4_outputs(1281) <= not(layer3_outputs(4979));
    layer4_outputs(1282) <= (layer3_outputs(4622)) and not (layer3_outputs(641));
    layer4_outputs(1283) <= '1';
    layer4_outputs(1284) <= not(layer3_outputs(196)) or (layer3_outputs(2986));
    layer4_outputs(1285) <= '1';
    layer4_outputs(1286) <= (layer3_outputs(524)) xor (layer3_outputs(557));
    layer4_outputs(1287) <= '1';
    layer4_outputs(1288) <= not(layer3_outputs(3336)) or (layer3_outputs(3534));
    layer4_outputs(1289) <= (layer3_outputs(693)) and (layer3_outputs(2522));
    layer4_outputs(1290) <= not((layer3_outputs(119)) and (layer3_outputs(3850)));
    layer4_outputs(1291) <= layer3_outputs(1625);
    layer4_outputs(1292) <= not(layer3_outputs(3880)) or (layer3_outputs(1479));
    layer4_outputs(1293) <= '0';
    layer4_outputs(1294) <= (layer3_outputs(2640)) and not (layer3_outputs(983));
    layer4_outputs(1295) <= not(layer3_outputs(4509)) or (layer3_outputs(4013));
    layer4_outputs(1296) <= '1';
    layer4_outputs(1297) <= not(layer3_outputs(1194)) or (layer3_outputs(4464));
    layer4_outputs(1298) <= (layer3_outputs(4417)) or (layer3_outputs(2730));
    layer4_outputs(1299) <= not(layer3_outputs(3663)) or (layer3_outputs(746));
    layer4_outputs(1300) <= not((layer3_outputs(3969)) and (layer3_outputs(372)));
    layer4_outputs(1301) <= not(layer3_outputs(2225));
    layer4_outputs(1302) <= not(layer3_outputs(3098));
    layer4_outputs(1303) <= (layer3_outputs(934)) or (layer3_outputs(3580));
    layer4_outputs(1304) <= not(layer3_outputs(2461)) or (layer3_outputs(48));
    layer4_outputs(1305) <= not(layer3_outputs(1088)) or (layer3_outputs(2916));
    layer4_outputs(1306) <= not(layer3_outputs(1738));
    layer4_outputs(1307) <= not(layer3_outputs(3008)) or (layer3_outputs(1349));
    layer4_outputs(1308) <= '0';
    layer4_outputs(1309) <= layer3_outputs(4328);
    layer4_outputs(1310) <= '1';
    layer4_outputs(1311) <= '0';
    layer4_outputs(1312) <= (layer3_outputs(3446)) and (layer3_outputs(4020));
    layer4_outputs(1313) <= (layer3_outputs(1832)) and (layer3_outputs(5050));
    layer4_outputs(1314) <= not(layer3_outputs(974));
    layer4_outputs(1315) <= '0';
    layer4_outputs(1316) <= not((layer3_outputs(2707)) and (layer3_outputs(3181)));
    layer4_outputs(1317) <= (layer3_outputs(3782)) and not (layer3_outputs(4568));
    layer4_outputs(1318) <= not(layer3_outputs(2703)) or (layer3_outputs(3727));
    layer4_outputs(1319) <= not((layer3_outputs(4375)) xor (layer3_outputs(1104)));
    layer4_outputs(1320) <= '0';
    layer4_outputs(1321) <= (layer3_outputs(2326)) and not (layer3_outputs(702));
    layer4_outputs(1322) <= '1';
    layer4_outputs(1323) <= layer3_outputs(632);
    layer4_outputs(1324) <= not(layer3_outputs(4201));
    layer4_outputs(1325) <= not(layer3_outputs(3022));
    layer4_outputs(1326) <= (layer3_outputs(1892)) and (layer3_outputs(230));
    layer4_outputs(1327) <= layer3_outputs(627);
    layer4_outputs(1328) <= (layer3_outputs(1831)) and (layer3_outputs(1632));
    layer4_outputs(1329) <= not(layer3_outputs(600));
    layer4_outputs(1330) <= (layer3_outputs(2540)) and not (layer3_outputs(1804));
    layer4_outputs(1331) <= layer3_outputs(771);
    layer4_outputs(1332) <= layer3_outputs(861);
    layer4_outputs(1333) <= layer3_outputs(4851);
    layer4_outputs(1334) <= not(layer3_outputs(2490));
    layer4_outputs(1335) <= layer3_outputs(2896);
    layer4_outputs(1336) <= layer3_outputs(3688);
    layer4_outputs(1337) <= (layer3_outputs(981)) and (layer3_outputs(3264));
    layer4_outputs(1338) <= '0';
    layer4_outputs(1339) <= not(layer3_outputs(3284)) or (layer3_outputs(4822));
    layer4_outputs(1340) <= layer3_outputs(4731);
    layer4_outputs(1341) <= not(layer3_outputs(4170));
    layer4_outputs(1342) <= not(layer3_outputs(2315));
    layer4_outputs(1343) <= not(layer3_outputs(4929)) or (layer3_outputs(222));
    layer4_outputs(1344) <= not(layer3_outputs(2767));
    layer4_outputs(1345) <= layer3_outputs(447);
    layer4_outputs(1346) <= layer3_outputs(1373);
    layer4_outputs(1347) <= layer3_outputs(1690);
    layer4_outputs(1348) <= not((layer3_outputs(3785)) or (layer3_outputs(1423)));
    layer4_outputs(1349) <= (layer3_outputs(4760)) and (layer3_outputs(3526));
    layer4_outputs(1350) <= (layer3_outputs(2155)) or (layer3_outputs(2356));
    layer4_outputs(1351) <= not(layer3_outputs(1355));
    layer4_outputs(1352) <= (layer3_outputs(191)) and (layer3_outputs(1910));
    layer4_outputs(1353) <= '0';
    layer4_outputs(1354) <= not(layer3_outputs(507));
    layer4_outputs(1355) <= (layer3_outputs(871)) or (layer3_outputs(3996));
    layer4_outputs(1356) <= (layer3_outputs(2096)) and not (layer3_outputs(3581));
    layer4_outputs(1357) <= (layer3_outputs(3432)) and not (layer3_outputs(2758));
    layer4_outputs(1358) <= not((layer3_outputs(1924)) xor (layer3_outputs(4468)));
    layer4_outputs(1359) <= not(layer3_outputs(1126));
    layer4_outputs(1360) <= (layer3_outputs(272)) and not (layer3_outputs(1712));
    layer4_outputs(1361) <= (layer3_outputs(2073)) or (layer3_outputs(2631));
    layer4_outputs(1362) <= not(layer3_outputs(1737)) or (layer3_outputs(4545));
    layer4_outputs(1363) <= not((layer3_outputs(3901)) or (layer3_outputs(2695)));
    layer4_outputs(1364) <= (layer3_outputs(806)) and (layer3_outputs(3418));
    layer4_outputs(1365) <= not(layer3_outputs(2644)) or (layer3_outputs(76));
    layer4_outputs(1366) <= '0';
    layer4_outputs(1367) <= (layer3_outputs(3062)) and not (layer3_outputs(2116));
    layer4_outputs(1368) <= not(layer3_outputs(1123));
    layer4_outputs(1369) <= layer3_outputs(2583);
    layer4_outputs(1370) <= not((layer3_outputs(4192)) or (layer3_outputs(1294)));
    layer4_outputs(1371) <= not(layer3_outputs(2242));
    layer4_outputs(1372) <= not(layer3_outputs(2242)) or (layer3_outputs(3781));
    layer4_outputs(1373) <= not(layer3_outputs(4726));
    layer4_outputs(1374) <= layer3_outputs(3904);
    layer4_outputs(1375) <= not((layer3_outputs(122)) and (layer3_outputs(452)));
    layer4_outputs(1376) <= (layer3_outputs(2619)) and not (layer3_outputs(4032));
    layer4_outputs(1377) <= (layer3_outputs(3323)) and not (layer3_outputs(538));
    layer4_outputs(1378) <= (layer3_outputs(1728)) and not (layer3_outputs(3306));
    layer4_outputs(1379) <= layer3_outputs(1582);
    layer4_outputs(1380) <= (layer3_outputs(4110)) and (layer3_outputs(4983));
    layer4_outputs(1381) <= (layer3_outputs(2567)) and not (layer3_outputs(3340));
    layer4_outputs(1382) <= not((layer3_outputs(4246)) or (layer3_outputs(2755)));
    layer4_outputs(1383) <= '1';
    layer4_outputs(1384) <= (layer3_outputs(1614)) and not (layer3_outputs(3552));
    layer4_outputs(1385) <= (layer3_outputs(2325)) and not (layer3_outputs(1087));
    layer4_outputs(1386) <= (layer3_outputs(607)) or (layer3_outputs(3538));
    layer4_outputs(1387) <= not(layer3_outputs(1839)) or (layer3_outputs(359));
    layer4_outputs(1388) <= not((layer3_outputs(4380)) and (layer3_outputs(1022)));
    layer4_outputs(1389) <= '0';
    layer4_outputs(1390) <= layer3_outputs(712);
    layer4_outputs(1391) <= not(layer3_outputs(2838)) or (layer3_outputs(4745));
    layer4_outputs(1392) <= not((layer3_outputs(5077)) and (layer3_outputs(2275)));
    layer4_outputs(1393) <= not((layer3_outputs(2501)) or (layer3_outputs(573)));
    layer4_outputs(1394) <= not((layer3_outputs(3379)) xor (layer3_outputs(4227)));
    layer4_outputs(1395) <= layer3_outputs(2950);
    layer4_outputs(1396) <= not(layer3_outputs(577));
    layer4_outputs(1397) <= not(layer3_outputs(4998));
    layer4_outputs(1398) <= not(layer3_outputs(2847));
    layer4_outputs(1399) <= (layer3_outputs(2377)) or (layer3_outputs(4801));
    layer4_outputs(1400) <= '0';
    layer4_outputs(1401) <= not(layer3_outputs(1682)) or (layer3_outputs(4775));
    layer4_outputs(1402) <= (layer3_outputs(2947)) and not (layer3_outputs(2403));
    layer4_outputs(1403) <= layer3_outputs(2106);
    layer4_outputs(1404) <= layer3_outputs(303);
    layer4_outputs(1405) <= not(layer3_outputs(3163)) or (layer3_outputs(3533));
    layer4_outputs(1406) <= (layer3_outputs(3504)) and (layer3_outputs(4522));
    layer4_outputs(1407) <= not(layer3_outputs(1854));
    layer4_outputs(1408) <= layer3_outputs(2765);
    layer4_outputs(1409) <= not(layer3_outputs(2246));
    layer4_outputs(1410) <= layer3_outputs(3819);
    layer4_outputs(1411) <= not(layer3_outputs(1114));
    layer4_outputs(1412) <= (layer3_outputs(1851)) and not (layer3_outputs(1748));
    layer4_outputs(1413) <= (layer3_outputs(3347)) or (layer3_outputs(2469));
    layer4_outputs(1414) <= (layer3_outputs(4546)) and not (layer3_outputs(3192));
    layer4_outputs(1415) <= layer3_outputs(1152);
    layer4_outputs(1416) <= not(layer3_outputs(3836));
    layer4_outputs(1417) <= not(layer3_outputs(3061)) or (layer3_outputs(2038));
    layer4_outputs(1418) <= (layer3_outputs(1260)) and not (layer3_outputs(2155));
    layer4_outputs(1419) <= '0';
    layer4_outputs(1420) <= (layer3_outputs(1921)) and (layer3_outputs(1518));
    layer4_outputs(1421) <= (layer3_outputs(1986)) and not (layer3_outputs(4767));
    layer4_outputs(1422) <= not((layer3_outputs(1685)) and (layer3_outputs(2156)));
    layer4_outputs(1423) <= '1';
    layer4_outputs(1424) <= '0';
    layer4_outputs(1425) <= not(layer3_outputs(1866));
    layer4_outputs(1426) <= not((layer3_outputs(2622)) and (layer3_outputs(3069)));
    layer4_outputs(1427) <= layer3_outputs(4631);
    layer4_outputs(1428) <= layer3_outputs(4886);
    layer4_outputs(1429) <= not((layer3_outputs(2042)) or (layer3_outputs(218)));
    layer4_outputs(1430) <= (layer3_outputs(984)) or (layer3_outputs(3929));
    layer4_outputs(1431) <= not(layer3_outputs(526)) or (layer3_outputs(3150));
    layer4_outputs(1432) <= not((layer3_outputs(3310)) or (layer3_outputs(3723)));
    layer4_outputs(1433) <= not(layer3_outputs(1816));
    layer4_outputs(1434) <= not((layer3_outputs(1521)) and (layer3_outputs(619)));
    layer4_outputs(1435) <= '1';
    layer4_outputs(1436) <= not(layer3_outputs(1538));
    layer4_outputs(1437) <= not((layer3_outputs(2528)) and (layer3_outputs(650)));
    layer4_outputs(1438) <= layer3_outputs(708);
    layer4_outputs(1439) <= (layer3_outputs(4636)) and not (layer3_outputs(2543));
    layer4_outputs(1440) <= not((layer3_outputs(665)) and (layer3_outputs(4822)));
    layer4_outputs(1441) <= (layer3_outputs(4991)) and (layer3_outputs(2174));
    layer4_outputs(1442) <= '0';
    layer4_outputs(1443) <= not(layer3_outputs(3535));
    layer4_outputs(1444) <= (layer3_outputs(4012)) and not (layer3_outputs(2015));
    layer4_outputs(1445) <= '1';
    layer4_outputs(1446) <= layer3_outputs(3110);
    layer4_outputs(1447) <= (layer3_outputs(498)) and not (layer3_outputs(4794));
    layer4_outputs(1448) <= layer3_outputs(1366);
    layer4_outputs(1449) <= (layer3_outputs(2438)) and not (layer3_outputs(2264));
    layer4_outputs(1450) <= (layer3_outputs(4466)) and (layer3_outputs(3585));
    layer4_outputs(1451) <= '0';
    layer4_outputs(1452) <= not(layer3_outputs(1072)) or (layer3_outputs(2015));
    layer4_outputs(1453) <= not((layer3_outputs(886)) and (layer3_outputs(151)));
    layer4_outputs(1454) <= not(layer3_outputs(2369));
    layer4_outputs(1455) <= layer3_outputs(3666);
    layer4_outputs(1456) <= (layer3_outputs(4038)) and not (layer3_outputs(3149));
    layer4_outputs(1457) <= not((layer3_outputs(1757)) and (layer3_outputs(3388)));
    layer4_outputs(1458) <= '0';
    layer4_outputs(1459) <= not(layer3_outputs(3523)) or (layer3_outputs(338));
    layer4_outputs(1460) <= (layer3_outputs(919)) or (layer3_outputs(4664));
    layer4_outputs(1461) <= (layer3_outputs(4310)) or (layer3_outputs(2379));
    layer4_outputs(1462) <= not(layer3_outputs(502));
    layer4_outputs(1463) <= not(layer3_outputs(4088));
    layer4_outputs(1464) <= (layer3_outputs(4955)) or (layer3_outputs(1241));
    layer4_outputs(1465) <= (layer3_outputs(3015)) and not (layer3_outputs(3623));
    layer4_outputs(1466) <= '0';
    layer4_outputs(1467) <= (layer3_outputs(2829)) or (layer3_outputs(5032));
    layer4_outputs(1468) <= not(layer3_outputs(4660)) or (layer3_outputs(595));
    layer4_outputs(1469) <= not((layer3_outputs(2248)) or (layer3_outputs(380)));
    layer4_outputs(1470) <= (layer3_outputs(1527)) and not (layer3_outputs(4555));
    layer4_outputs(1471) <= (layer3_outputs(1134)) xor (layer3_outputs(3422));
    layer4_outputs(1472) <= not(layer3_outputs(1135));
    layer4_outputs(1473) <= (layer3_outputs(1127)) and not (layer3_outputs(3723));
    layer4_outputs(1474) <= layer3_outputs(1980);
    layer4_outputs(1475) <= (layer3_outputs(3648)) or (layer3_outputs(2929));
    layer4_outputs(1476) <= not((layer3_outputs(4236)) or (layer3_outputs(1650)));
    layer4_outputs(1477) <= (layer3_outputs(4155)) and not (layer3_outputs(441));
    layer4_outputs(1478) <= (layer3_outputs(1304)) or (layer3_outputs(1925));
    layer4_outputs(1479) <= layer3_outputs(3608);
    layer4_outputs(1480) <= not(layer3_outputs(169));
    layer4_outputs(1481) <= (layer3_outputs(3494)) and not (layer3_outputs(3141));
    layer4_outputs(1482) <= '0';
    layer4_outputs(1483) <= not((layer3_outputs(4280)) and (layer3_outputs(2614)));
    layer4_outputs(1484) <= (layer3_outputs(4779)) and not (layer3_outputs(344));
    layer4_outputs(1485) <= (layer3_outputs(2265)) and not (layer3_outputs(1949));
    layer4_outputs(1486) <= not(layer3_outputs(1063));
    layer4_outputs(1487) <= (layer3_outputs(4003)) and not (layer3_outputs(4342));
    layer4_outputs(1488) <= not((layer3_outputs(1570)) or (layer3_outputs(3781)));
    layer4_outputs(1489) <= '0';
    layer4_outputs(1490) <= layer3_outputs(4055);
    layer4_outputs(1491) <= not(layer3_outputs(3972)) or (layer3_outputs(3419));
    layer4_outputs(1492) <= not(layer3_outputs(4880)) or (layer3_outputs(4714));
    layer4_outputs(1493) <= (layer3_outputs(649)) and not (layer3_outputs(3289));
    layer4_outputs(1494) <= not((layer3_outputs(5037)) and (layer3_outputs(2933)));
    layer4_outputs(1495) <= not(layer3_outputs(122));
    layer4_outputs(1496) <= layer3_outputs(716);
    layer4_outputs(1497) <= not(layer3_outputs(4878));
    layer4_outputs(1498) <= layer3_outputs(655);
    layer4_outputs(1499) <= (layer3_outputs(4954)) and not (layer3_outputs(5025));
    layer4_outputs(1500) <= not(layer3_outputs(4148));
    layer4_outputs(1501) <= (layer3_outputs(3332)) or (layer3_outputs(4402));
    layer4_outputs(1502) <= not(layer3_outputs(4354)) or (layer3_outputs(1675));
    layer4_outputs(1503) <= not((layer3_outputs(2205)) or (layer3_outputs(1334)));
    layer4_outputs(1504) <= '1';
    layer4_outputs(1505) <= (layer3_outputs(1656)) and not (layer3_outputs(2649));
    layer4_outputs(1506) <= (layer3_outputs(4049)) or (layer3_outputs(378));
    layer4_outputs(1507) <= layer3_outputs(1512);
    layer4_outputs(1508) <= (layer3_outputs(2139)) xor (layer3_outputs(421));
    layer4_outputs(1509) <= layer3_outputs(3294);
    layer4_outputs(1510) <= layer3_outputs(1974);
    layer4_outputs(1511) <= not(layer3_outputs(3393)) or (layer3_outputs(1997));
    layer4_outputs(1512) <= '1';
    layer4_outputs(1513) <= layer3_outputs(3647);
    layer4_outputs(1514) <= '1';
    layer4_outputs(1515) <= '0';
    layer4_outputs(1516) <= '1';
    layer4_outputs(1517) <= not(layer3_outputs(440));
    layer4_outputs(1518) <= (layer3_outputs(2222)) xor (layer3_outputs(2765));
    layer4_outputs(1519) <= (layer3_outputs(497)) and not (layer3_outputs(4620));
    layer4_outputs(1520) <= not(layer3_outputs(3026));
    layer4_outputs(1521) <= (layer3_outputs(3860)) and (layer3_outputs(3797));
    layer4_outputs(1522) <= (layer3_outputs(3153)) and not (layer3_outputs(1090));
    layer4_outputs(1523) <= not(layer3_outputs(3355)) or (layer3_outputs(3591));
    layer4_outputs(1524) <= layer3_outputs(4495);
    layer4_outputs(1525) <= (layer3_outputs(4958)) or (layer3_outputs(2675));
    layer4_outputs(1526) <= (layer3_outputs(65)) xor (layer3_outputs(3659));
    layer4_outputs(1527) <= (layer3_outputs(4783)) and not (layer3_outputs(1359));
    layer4_outputs(1528) <= (layer3_outputs(4456)) and not (layer3_outputs(4887));
    layer4_outputs(1529) <= not(layer3_outputs(1378)) or (layer3_outputs(2689));
    layer4_outputs(1530) <= '0';
    layer4_outputs(1531) <= not((layer3_outputs(2421)) and (layer3_outputs(4723)));
    layer4_outputs(1532) <= '0';
    layer4_outputs(1533) <= '0';
    layer4_outputs(1534) <= (layer3_outputs(3401)) and (layer3_outputs(1696));
    layer4_outputs(1535) <= not(layer3_outputs(3331));
    layer4_outputs(1536) <= not(layer3_outputs(1441));
    layer4_outputs(1537) <= layer3_outputs(2673);
    layer4_outputs(1538) <= (layer3_outputs(4336)) or (layer3_outputs(988));
    layer4_outputs(1539) <= (layer3_outputs(1635)) or (layer3_outputs(611));
    layer4_outputs(1540) <= not((layer3_outputs(1296)) or (layer3_outputs(2924)));
    layer4_outputs(1541) <= not(layer3_outputs(320));
    layer4_outputs(1542) <= (layer3_outputs(240)) and (layer3_outputs(2949));
    layer4_outputs(1543) <= not(layer3_outputs(4131)) or (layer3_outputs(2123));
    layer4_outputs(1544) <= layer3_outputs(2151);
    layer4_outputs(1545) <= layer3_outputs(4753);
    layer4_outputs(1546) <= (layer3_outputs(1318)) and not (layer3_outputs(2598));
    layer4_outputs(1547) <= not(layer3_outputs(3185)) or (layer3_outputs(1315));
    layer4_outputs(1548) <= not(layer3_outputs(1602)) or (layer3_outputs(3557));
    layer4_outputs(1549) <= '1';
    layer4_outputs(1550) <= layer3_outputs(2767);
    layer4_outputs(1551) <= not(layer3_outputs(3005));
    layer4_outputs(1552) <= '1';
    layer4_outputs(1553) <= not(layer3_outputs(2971)) or (layer3_outputs(162));
    layer4_outputs(1554) <= not((layer3_outputs(596)) and (layer3_outputs(661)));
    layer4_outputs(1555) <= (layer3_outputs(4120)) or (layer3_outputs(4462));
    layer4_outputs(1556) <= (layer3_outputs(4379)) and (layer3_outputs(2218));
    layer4_outputs(1557) <= not((layer3_outputs(1917)) or (layer3_outputs(2480)));
    layer4_outputs(1558) <= not((layer3_outputs(231)) and (layer3_outputs(2849)));
    layer4_outputs(1559) <= layer3_outputs(1433);
    layer4_outputs(1560) <= not((layer3_outputs(3777)) or (layer3_outputs(3344)));
    layer4_outputs(1561) <= not((layer3_outputs(2984)) and (layer3_outputs(2569)));
    layer4_outputs(1562) <= '0';
    layer4_outputs(1563) <= (layer3_outputs(2147)) and not (layer3_outputs(4453));
    layer4_outputs(1564) <= not(layer3_outputs(2342));
    layer4_outputs(1565) <= not((layer3_outputs(4159)) and (layer3_outputs(2142)));
    layer4_outputs(1566) <= layer3_outputs(4915);
    layer4_outputs(1567) <= not((layer3_outputs(2706)) or (layer3_outputs(3281)));
    layer4_outputs(1568) <= not(layer3_outputs(2976)) or (layer3_outputs(548));
    layer4_outputs(1569) <= (layer3_outputs(1101)) and not (layer3_outputs(5102));
    layer4_outputs(1570) <= not(layer3_outputs(4843));
    layer4_outputs(1571) <= '1';
    layer4_outputs(1572) <= not((layer3_outputs(2782)) and (layer3_outputs(4366)));
    layer4_outputs(1573) <= not(layer3_outputs(4200));
    layer4_outputs(1574) <= (layer3_outputs(4903)) and not (layer3_outputs(3329));
    layer4_outputs(1575) <= (layer3_outputs(2599)) and not (layer3_outputs(2521));
    layer4_outputs(1576) <= not(layer3_outputs(4971));
    layer4_outputs(1577) <= not(layer3_outputs(1490)) or (layer3_outputs(3521));
    layer4_outputs(1578) <= not((layer3_outputs(4166)) or (layer3_outputs(1141)));
    layer4_outputs(1579) <= layer3_outputs(120);
    layer4_outputs(1580) <= (layer3_outputs(1454)) or (layer3_outputs(2464));
    layer4_outputs(1581) <= (layer3_outputs(4091)) or (layer3_outputs(2124));
    layer4_outputs(1582) <= not(layer3_outputs(3924)) or (layer3_outputs(1933));
    layer4_outputs(1583) <= (layer3_outputs(4553)) and not (layer3_outputs(2856));
    layer4_outputs(1584) <= '1';
    layer4_outputs(1585) <= not(layer3_outputs(4993));
    layer4_outputs(1586) <= (layer3_outputs(4948)) and not (layer3_outputs(3578));
    layer4_outputs(1587) <= not(layer3_outputs(700));
    layer4_outputs(1588) <= (layer3_outputs(2508)) and (layer3_outputs(3675));
    layer4_outputs(1589) <= (layer3_outputs(3038)) and not (layer3_outputs(4027));
    layer4_outputs(1590) <= '0';
    layer4_outputs(1591) <= (layer3_outputs(1375)) and not (layer3_outputs(2776));
    layer4_outputs(1592) <= layer3_outputs(3622);
    layer4_outputs(1593) <= '1';
    layer4_outputs(1594) <= not(layer3_outputs(3692));
    layer4_outputs(1595) <= not(layer3_outputs(3619));
    layer4_outputs(1596) <= not(layer3_outputs(3012)) or (layer3_outputs(3089));
    layer4_outputs(1597) <= not(layer3_outputs(1574));
    layer4_outputs(1598) <= not((layer3_outputs(1509)) and (layer3_outputs(1662)));
    layer4_outputs(1599) <= (layer3_outputs(4593)) and not (layer3_outputs(2136));
    layer4_outputs(1600) <= layer3_outputs(1206);
    layer4_outputs(1601) <= not(layer3_outputs(516));
    layer4_outputs(1602) <= not((layer3_outputs(149)) and (layer3_outputs(3774)));
    layer4_outputs(1603) <= not((layer3_outputs(2002)) or (layer3_outputs(2758)));
    layer4_outputs(1604) <= not(layer3_outputs(804));
    layer4_outputs(1605) <= not((layer3_outputs(1787)) or (layer3_outputs(367)));
    layer4_outputs(1606) <= not((layer3_outputs(208)) and (layer3_outputs(3337)));
    layer4_outputs(1607) <= (layer3_outputs(1067)) and not (layer3_outputs(1004));
    layer4_outputs(1608) <= (layer3_outputs(5088)) or (layer3_outputs(4967));
    layer4_outputs(1609) <= not(layer3_outputs(964)) or (layer3_outputs(44));
    layer4_outputs(1610) <= not((layer3_outputs(1067)) or (layer3_outputs(1790)));
    layer4_outputs(1611) <= layer3_outputs(4970);
    layer4_outputs(1612) <= (layer3_outputs(461)) or (layer3_outputs(4933));
    layer4_outputs(1613) <= '0';
    layer4_outputs(1614) <= layer3_outputs(1527);
    layer4_outputs(1615) <= (layer3_outputs(2179)) and not (layer3_outputs(3553));
    layer4_outputs(1616) <= not(layer3_outputs(3319)) or (layer3_outputs(4943));
    layer4_outputs(1617) <= not(layer3_outputs(87));
    layer4_outputs(1618) <= layer3_outputs(1580);
    layer4_outputs(1619) <= layer3_outputs(156);
    layer4_outputs(1620) <= not(layer3_outputs(2054)) or (layer3_outputs(3221));
    layer4_outputs(1621) <= (layer3_outputs(3885)) or (layer3_outputs(129));
    layer4_outputs(1622) <= (layer3_outputs(2974)) and not (layer3_outputs(2593));
    layer4_outputs(1623) <= '0';
    layer4_outputs(1624) <= not(layer3_outputs(2790)) or (layer3_outputs(4012));
    layer4_outputs(1625) <= not((layer3_outputs(3398)) xor (layer3_outputs(4288)));
    layer4_outputs(1626) <= layer3_outputs(5090);
    layer4_outputs(1627) <= (layer3_outputs(1015)) and not (layer3_outputs(1586));
    layer4_outputs(1628) <= (layer3_outputs(2868)) and (layer3_outputs(3864));
    layer4_outputs(1629) <= not((layer3_outputs(793)) and (layer3_outputs(4812)));
    layer4_outputs(1630) <= not(layer3_outputs(620));
    layer4_outputs(1631) <= not(layer3_outputs(2074));
    layer4_outputs(1632) <= not(layer3_outputs(3074));
    layer4_outputs(1633) <= '1';
    layer4_outputs(1634) <= not(layer3_outputs(54)) or (layer3_outputs(1587));
    layer4_outputs(1635) <= not(layer3_outputs(1312));
    layer4_outputs(1636) <= not((layer3_outputs(3656)) and (layer3_outputs(2353)));
    layer4_outputs(1637) <= layer3_outputs(708);
    layer4_outputs(1638) <= not(layer3_outputs(2619));
    layer4_outputs(1639) <= (layer3_outputs(1873)) and not (layer3_outputs(1012));
    layer4_outputs(1640) <= not((layer3_outputs(1599)) xor (layer3_outputs(4747)));
    layer4_outputs(1641) <= (layer3_outputs(5057)) xor (layer3_outputs(1453));
    layer4_outputs(1642) <= (layer3_outputs(3851)) and not (layer3_outputs(1962));
    layer4_outputs(1643) <= layer3_outputs(3130);
    layer4_outputs(1644) <= (layer3_outputs(1077)) and not (layer3_outputs(119));
    layer4_outputs(1645) <= not(layer3_outputs(717)) or (layer3_outputs(3468));
    layer4_outputs(1646) <= not(layer3_outputs(1078));
    layer4_outputs(1647) <= (layer3_outputs(3118)) and not (layer3_outputs(1867));
    layer4_outputs(1648) <= layer3_outputs(1411);
    layer4_outputs(1649) <= (layer3_outputs(2398)) and (layer3_outputs(2175));
    layer4_outputs(1650) <= not(layer3_outputs(232)) or (layer3_outputs(1076));
    layer4_outputs(1651) <= not(layer3_outputs(4423));
    layer4_outputs(1652) <= layer3_outputs(160);
    layer4_outputs(1653) <= not((layer3_outputs(4917)) and (layer3_outputs(2132)));
    layer4_outputs(1654) <= not(layer3_outputs(4637));
    layer4_outputs(1655) <= not((layer3_outputs(777)) xor (layer3_outputs(3910)));
    layer4_outputs(1656) <= not((layer3_outputs(2176)) or (layer3_outputs(2350)));
    layer4_outputs(1657) <= (layer3_outputs(3021)) and (layer3_outputs(1799));
    layer4_outputs(1658) <= (layer3_outputs(1857)) and (layer3_outputs(3992));
    layer4_outputs(1659) <= layer3_outputs(4925);
    layer4_outputs(1660) <= layer3_outputs(3412);
    layer4_outputs(1661) <= layer3_outputs(1488);
    layer4_outputs(1662) <= not(layer3_outputs(401)) or (layer3_outputs(4008));
    layer4_outputs(1663) <= '0';
    layer4_outputs(1664) <= not(layer3_outputs(4147)) or (layer3_outputs(1756));
    layer4_outputs(1665) <= not((layer3_outputs(4794)) or (layer3_outputs(2054)));
    layer4_outputs(1666) <= '0';
    layer4_outputs(1667) <= (layer3_outputs(3962)) xor (layer3_outputs(1444));
    layer4_outputs(1668) <= layer3_outputs(2080);
    layer4_outputs(1669) <= not((layer3_outputs(2587)) or (layer3_outputs(522)));
    layer4_outputs(1670) <= not((layer3_outputs(1759)) and (layer3_outputs(769)));
    layer4_outputs(1671) <= not(layer3_outputs(4829)) or (layer3_outputs(2309));
    layer4_outputs(1672) <= not((layer3_outputs(3095)) xor (layer3_outputs(1802)));
    layer4_outputs(1673) <= (layer3_outputs(2920)) and not (layer3_outputs(3077));
    layer4_outputs(1674) <= (layer3_outputs(3490)) and (layer3_outputs(3582));
    layer4_outputs(1675) <= (layer3_outputs(1456)) or (layer3_outputs(4412));
    layer4_outputs(1676) <= not((layer3_outputs(3665)) and (layer3_outputs(2945)));
    layer4_outputs(1677) <= (layer3_outputs(2050)) and (layer3_outputs(4562));
    layer4_outputs(1678) <= '1';
    layer4_outputs(1679) <= (layer3_outputs(1387)) and (layer3_outputs(3698));
    layer4_outputs(1680) <= layer3_outputs(3976);
    layer4_outputs(1681) <= (layer3_outputs(5033)) and not (layer3_outputs(1101));
    layer4_outputs(1682) <= (layer3_outputs(4658)) or (layer3_outputs(3084));
    layer4_outputs(1683) <= not((layer3_outputs(3373)) and (layer3_outputs(3372)));
    layer4_outputs(1684) <= layer3_outputs(3566);
    layer4_outputs(1685) <= not(layer3_outputs(704));
    layer4_outputs(1686) <= not((layer3_outputs(3820)) and (layer3_outputs(273)));
    layer4_outputs(1687) <= not((layer3_outputs(4399)) and (layer3_outputs(4005)));
    layer4_outputs(1688) <= (layer3_outputs(2320)) and not (layer3_outputs(2696));
    layer4_outputs(1689) <= (layer3_outputs(793)) and not (layer3_outputs(184));
    layer4_outputs(1690) <= '1';
    layer4_outputs(1691) <= layer3_outputs(3389);
    layer4_outputs(1692) <= layer3_outputs(750);
    layer4_outputs(1693) <= '0';
    layer4_outputs(1694) <= not(layer3_outputs(1882)) or (layer3_outputs(1149));
    layer4_outputs(1695) <= layer3_outputs(340);
    layer4_outputs(1696) <= (layer3_outputs(4141)) or (layer3_outputs(3027));
    layer4_outputs(1697) <= not((layer3_outputs(635)) xor (layer3_outputs(1619)));
    layer4_outputs(1698) <= '0';
    layer4_outputs(1699) <= '0';
    layer4_outputs(1700) <= not(layer3_outputs(2863));
    layer4_outputs(1701) <= '1';
    layer4_outputs(1702) <= '0';
    layer4_outputs(1703) <= (layer3_outputs(1226)) or (layer3_outputs(2185));
    layer4_outputs(1704) <= (layer3_outputs(3257)) and (layer3_outputs(1545));
    layer4_outputs(1705) <= (layer3_outputs(842)) and (layer3_outputs(3872));
    layer4_outputs(1706) <= not(layer3_outputs(3883));
    layer4_outputs(1707) <= (layer3_outputs(4544)) or (layer3_outputs(611));
    layer4_outputs(1708) <= layer3_outputs(1312);
    layer4_outputs(1709) <= layer3_outputs(4083);
    layer4_outputs(1710) <= (layer3_outputs(203)) and not (layer3_outputs(342));
    layer4_outputs(1711) <= not(layer3_outputs(1446));
    layer4_outputs(1712) <= layer3_outputs(1125);
    layer4_outputs(1713) <= not(layer3_outputs(3663));
    layer4_outputs(1714) <= not((layer3_outputs(2018)) or (layer3_outputs(4960)));
    layer4_outputs(1715) <= (layer3_outputs(806)) or (layer3_outputs(209));
    layer4_outputs(1716) <= '1';
    layer4_outputs(1717) <= not(layer3_outputs(1624)) or (layer3_outputs(934));
    layer4_outputs(1718) <= not((layer3_outputs(1238)) or (layer3_outputs(445)));
    layer4_outputs(1719) <= '1';
    layer4_outputs(1720) <= not(layer3_outputs(1972)) or (layer3_outputs(3454));
    layer4_outputs(1721) <= '0';
    layer4_outputs(1722) <= not(layer3_outputs(3544));
    layer4_outputs(1723) <= '1';
    layer4_outputs(1724) <= not((layer3_outputs(1878)) and (layer3_outputs(264)));
    layer4_outputs(1725) <= (layer3_outputs(386)) and not (layer3_outputs(273));
    layer4_outputs(1726) <= (layer3_outputs(2118)) and not (layer3_outputs(1931));
    layer4_outputs(1727) <= not(layer3_outputs(3449)) or (layer3_outputs(4487));
    layer4_outputs(1728) <= (layer3_outputs(2371)) and (layer3_outputs(2710));
    layer4_outputs(1729) <= not(layer3_outputs(1284));
    layer4_outputs(1730) <= layer3_outputs(3839);
    layer4_outputs(1731) <= not(layer3_outputs(2822));
    layer4_outputs(1732) <= not(layer3_outputs(4675)) or (layer3_outputs(2019));
    layer4_outputs(1733) <= not(layer3_outputs(1595)) or (layer3_outputs(2153));
    layer4_outputs(1734) <= layer3_outputs(1597);
    layer4_outputs(1735) <= layer3_outputs(2459);
    layer4_outputs(1736) <= not(layer3_outputs(339)) or (layer3_outputs(838));
    layer4_outputs(1737) <= layer3_outputs(4789);
    layer4_outputs(1738) <= not(layer3_outputs(1332));
    layer4_outputs(1739) <= layer3_outputs(2869);
    layer4_outputs(1740) <= not(layer3_outputs(4627));
    layer4_outputs(1741) <= layer3_outputs(4729);
    layer4_outputs(1742) <= layer3_outputs(1474);
    layer4_outputs(1743) <= '1';
    layer4_outputs(1744) <= (layer3_outputs(2563)) and (layer3_outputs(5106));
    layer4_outputs(1745) <= (layer3_outputs(1531)) and not (layer3_outputs(3624));
    layer4_outputs(1746) <= (layer3_outputs(830)) and not (layer3_outputs(564));
    layer4_outputs(1747) <= '0';
    layer4_outputs(1748) <= not(layer3_outputs(2510)) or (layer3_outputs(747));
    layer4_outputs(1749) <= layer3_outputs(4754);
    layer4_outputs(1750) <= not(layer3_outputs(188));
    layer4_outputs(1751) <= '1';
    layer4_outputs(1752) <= layer3_outputs(2174);
    layer4_outputs(1753) <= (layer3_outputs(164)) or (layer3_outputs(4001));
    layer4_outputs(1754) <= not((layer3_outputs(2246)) and (layer3_outputs(1735)));
    layer4_outputs(1755) <= not(layer3_outputs(891)) or (layer3_outputs(4413));
    layer4_outputs(1756) <= layer3_outputs(2558);
    layer4_outputs(1757) <= not((layer3_outputs(314)) and (layer3_outputs(1007)));
    layer4_outputs(1758) <= (layer3_outputs(2605)) and not (layer3_outputs(1977));
    layer4_outputs(1759) <= '1';
    layer4_outputs(1760) <= not(layer3_outputs(1948));
    layer4_outputs(1761) <= not(layer3_outputs(4524));
    layer4_outputs(1762) <= not(layer3_outputs(308));
    layer4_outputs(1763) <= layer3_outputs(2804);
    layer4_outputs(1764) <= (layer3_outputs(4393)) and (layer3_outputs(2351));
    layer4_outputs(1765) <= not(layer3_outputs(1491)) or (layer3_outputs(2170));
    layer4_outputs(1766) <= (layer3_outputs(1514)) and not (layer3_outputs(1281));
    layer4_outputs(1767) <= layer3_outputs(306);
    layer4_outputs(1768) <= '1';
    layer4_outputs(1769) <= not((layer3_outputs(1798)) or (layer3_outputs(4647)));
    layer4_outputs(1770) <= layer3_outputs(42);
    layer4_outputs(1771) <= (layer3_outputs(5050)) and not (layer3_outputs(527));
    layer4_outputs(1772) <= not(layer3_outputs(3277));
    layer4_outputs(1773) <= '0';
    layer4_outputs(1774) <= not(layer3_outputs(2367));
    layer4_outputs(1775) <= (layer3_outputs(3226)) and not (layer3_outputs(2407));
    layer4_outputs(1776) <= '0';
    layer4_outputs(1777) <= '0';
    layer4_outputs(1778) <= layer3_outputs(1653);
    layer4_outputs(1779) <= not(layer3_outputs(1038)) or (layer3_outputs(3196));
    layer4_outputs(1780) <= not((layer3_outputs(2290)) or (layer3_outputs(140)));
    layer4_outputs(1781) <= '0';
    layer4_outputs(1782) <= not(layer3_outputs(1635)) or (layer3_outputs(3737));
    layer4_outputs(1783) <= not(layer3_outputs(681)) or (layer3_outputs(704));
    layer4_outputs(1784) <= not(layer3_outputs(3088)) or (layer3_outputs(4609));
    layer4_outputs(1785) <= not(layer3_outputs(2127));
    layer4_outputs(1786) <= not(layer3_outputs(3474));
    layer4_outputs(1787) <= not(layer3_outputs(1945)) or (layer3_outputs(3389));
    layer4_outputs(1788) <= (layer3_outputs(5065)) and not (layer3_outputs(4108));
    layer4_outputs(1789) <= (layer3_outputs(5085)) and not (layer3_outputs(911));
    layer4_outputs(1790) <= (layer3_outputs(1220)) or (layer3_outputs(1820));
    layer4_outputs(1791) <= (layer3_outputs(2087)) and not (layer3_outputs(5103));
    layer4_outputs(1792) <= not(layer3_outputs(3475)) or (layer3_outputs(4440));
    layer4_outputs(1793) <= not(layer3_outputs(4985));
    layer4_outputs(1794) <= not(layer3_outputs(3513));
    layer4_outputs(1795) <= not((layer3_outputs(4792)) or (layer3_outputs(3559)));
    layer4_outputs(1796) <= not(layer3_outputs(4621));
    layer4_outputs(1797) <= (layer3_outputs(2603)) and not (layer3_outputs(3270));
    layer4_outputs(1798) <= not((layer3_outputs(2482)) and (layer3_outputs(356)));
    layer4_outputs(1799) <= '1';
    layer4_outputs(1800) <= (layer3_outputs(3683)) and (layer3_outputs(4357));
    layer4_outputs(1801) <= (layer3_outputs(1913)) and (layer3_outputs(2978));
    layer4_outputs(1802) <= layer3_outputs(3495);
    layer4_outputs(1803) <= (layer3_outputs(2025)) and not (layer3_outputs(3835));
    layer4_outputs(1804) <= not(layer3_outputs(2462));
    layer4_outputs(1805) <= not(layer3_outputs(3235));
    layer4_outputs(1806) <= '0';
    layer4_outputs(1807) <= layer3_outputs(5100);
    layer4_outputs(1808) <= '1';
    layer4_outputs(1809) <= '0';
    layer4_outputs(1810) <= (layer3_outputs(3305)) and not (layer3_outputs(2180));
    layer4_outputs(1811) <= (layer3_outputs(2954)) and (layer3_outputs(402));
    layer4_outputs(1812) <= layer3_outputs(3655);
    layer4_outputs(1813) <= not(layer3_outputs(3684)) or (layer3_outputs(4222));
    layer4_outputs(1814) <= not(layer3_outputs(161));
    layer4_outputs(1815) <= (layer3_outputs(336)) and (layer3_outputs(1753));
    layer4_outputs(1816) <= layer3_outputs(738);
    layer4_outputs(1817) <= (layer3_outputs(3124)) and not (layer3_outputs(823));
    layer4_outputs(1818) <= layer3_outputs(2052);
    layer4_outputs(1819) <= (layer3_outputs(2599)) and not (layer3_outputs(2527));
    layer4_outputs(1820) <= not((layer3_outputs(3842)) or (layer3_outputs(3649)));
    layer4_outputs(1821) <= not(layer3_outputs(4065)) or (layer3_outputs(4128));
    layer4_outputs(1822) <= (layer3_outputs(4368)) and (layer3_outputs(2575));
    layer4_outputs(1823) <= not(layer3_outputs(3087));
    layer4_outputs(1824) <= '1';
    layer4_outputs(1825) <= (layer3_outputs(664)) and not (layer3_outputs(5043));
    layer4_outputs(1826) <= layer3_outputs(4491);
    layer4_outputs(1827) <= (layer3_outputs(4788)) and not (layer3_outputs(1818));
    layer4_outputs(1828) <= not(layer3_outputs(3638)) or (layer3_outputs(2065));
    layer4_outputs(1829) <= layer3_outputs(974);
    layer4_outputs(1830) <= not((layer3_outputs(4263)) or (layer3_outputs(833)));
    layer4_outputs(1831) <= (layer3_outputs(121)) and (layer3_outputs(1304));
    layer4_outputs(1832) <= '1';
    layer4_outputs(1833) <= (layer3_outputs(1040)) or (layer3_outputs(2550));
    layer4_outputs(1834) <= (layer3_outputs(396)) and not (layer3_outputs(3577));
    layer4_outputs(1835) <= '0';
    layer4_outputs(1836) <= not((layer3_outputs(4811)) or (layer3_outputs(2177)));
    layer4_outputs(1837) <= layer3_outputs(4206);
    layer4_outputs(1838) <= '1';
    layer4_outputs(1839) <= '0';
    layer4_outputs(1840) <= not(layer3_outputs(3040)) or (layer3_outputs(595));
    layer4_outputs(1841) <= layer3_outputs(1625);
    layer4_outputs(1842) <= not((layer3_outputs(2423)) and (layer3_outputs(3370)));
    layer4_outputs(1843) <= not(layer3_outputs(5070));
    layer4_outputs(1844) <= layer3_outputs(3413);
    layer4_outputs(1845) <= not(layer3_outputs(4449));
    layer4_outputs(1846) <= '0';
    layer4_outputs(1847) <= not(layer3_outputs(4533));
    layer4_outputs(1848) <= not(layer3_outputs(1559));
    layer4_outputs(1849) <= (layer3_outputs(93)) and not (layer3_outputs(295));
    layer4_outputs(1850) <= not(layer3_outputs(545));
    layer4_outputs(1851) <= (layer3_outputs(2393)) and not (layer3_outputs(569));
    layer4_outputs(1852) <= (layer3_outputs(3254)) or (layer3_outputs(3102));
    layer4_outputs(1853) <= not(layer3_outputs(1964));
    layer4_outputs(1854) <= (layer3_outputs(3070)) and not (layer3_outputs(2375));
    layer4_outputs(1855) <= not((layer3_outputs(1155)) or (layer3_outputs(2224)));
    layer4_outputs(1856) <= layer3_outputs(2026);
    layer4_outputs(1857) <= (layer3_outputs(4245)) or (layer3_outputs(4945));
    layer4_outputs(1858) <= not((layer3_outputs(1732)) and (layer3_outputs(2299)));
    layer4_outputs(1859) <= not((layer3_outputs(459)) or (layer3_outputs(4861)));
    layer4_outputs(1860) <= layer3_outputs(3123);
    layer4_outputs(1861) <= not((layer3_outputs(1781)) or (layer3_outputs(3644)));
    layer4_outputs(1862) <= not((layer3_outputs(4397)) and (layer3_outputs(800)));
    layer4_outputs(1863) <= not(layer3_outputs(1210));
    layer4_outputs(1864) <= not(layer3_outputs(865));
    layer4_outputs(1865) <= (layer3_outputs(4562)) xor (layer3_outputs(2855));
    layer4_outputs(1866) <= '1';
    layer4_outputs(1867) <= not(layer3_outputs(3246));
    layer4_outputs(1868) <= not(layer3_outputs(2741)) or (layer3_outputs(4935));
    layer4_outputs(1869) <= (layer3_outputs(216)) and not (layer3_outputs(4977));
    layer4_outputs(1870) <= layer3_outputs(2560);
    layer4_outputs(1871) <= not(layer3_outputs(1083));
    layer4_outputs(1872) <= layer3_outputs(2343);
    layer4_outputs(1873) <= '0';
    layer4_outputs(1874) <= not(layer3_outputs(4450));
    layer4_outputs(1875) <= (layer3_outputs(2913)) and not (layer3_outputs(2484));
    layer4_outputs(1876) <= not((layer3_outputs(129)) xor (layer3_outputs(897)));
    layer4_outputs(1877) <= not(layer3_outputs(314)) or (layer3_outputs(1869));
    layer4_outputs(1878) <= not(layer3_outputs(2661));
    layer4_outputs(1879) <= not(layer3_outputs(3840)) or (layer3_outputs(3259));
    layer4_outputs(1880) <= '0';
    layer4_outputs(1881) <= layer3_outputs(776);
    layer4_outputs(1882) <= not(layer3_outputs(5013)) or (layer3_outputs(4500));
    layer4_outputs(1883) <= not(layer3_outputs(4854));
    layer4_outputs(1884) <= not(layer3_outputs(350)) or (layer3_outputs(5107));
    layer4_outputs(1885) <= (layer3_outputs(1562)) or (layer3_outputs(234));
    layer4_outputs(1886) <= not(layer3_outputs(448)) or (layer3_outputs(1529));
    layer4_outputs(1887) <= (layer3_outputs(1310)) and not (layer3_outputs(5074));
    layer4_outputs(1888) <= not(layer3_outputs(3293));
    layer4_outputs(1889) <= not(layer3_outputs(2939)) or (layer3_outputs(4512));
    layer4_outputs(1890) <= (layer3_outputs(144)) and not (layer3_outputs(2821));
    layer4_outputs(1891) <= not(layer3_outputs(1496));
    layer4_outputs(1892) <= not(layer3_outputs(1049)) or (layer3_outputs(2091));
    layer4_outputs(1893) <= not((layer3_outputs(3182)) xor (layer3_outputs(4019)));
    layer4_outputs(1894) <= (layer3_outputs(380)) and not (layer3_outputs(3773));
    layer4_outputs(1895) <= '1';
    layer4_outputs(1896) <= not(layer3_outputs(2195)) or (layer3_outputs(3889));
    layer4_outputs(1897) <= not(layer3_outputs(4849)) or (layer3_outputs(4291));
    layer4_outputs(1898) <= (layer3_outputs(2919)) and not (layer3_outputs(1771));
    layer4_outputs(1899) <= not(layer3_outputs(966)) or (layer3_outputs(1568));
    layer4_outputs(1900) <= (layer3_outputs(4403)) or (layer3_outputs(4845));
    layer4_outputs(1901) <= (layer3_outputs(4844)) and not (layer3_outputs(4083));
    layer4_outputs(1902) <= (layer3_outputs(325)) xor (layer3_outputs(4381));
    layer4_outputs(1903) <= layer3_outputs(4502);
    layer4_outputs(1904) <= not((layer3_outputs(457)) and (layer3_outputs(1309)));
    layer4_outputs(1905) <= (layer3_outputs(4726)) or (layer3_outputs(3460));
    layer4_outputs(1906) <= '0';
    layer4_outputs(1907) <= (layer3_outputs(2722)) or (layer3_outputs(331));
    layer4_outputs(1908) <= (layer3_outputs(605)) or (layer3_outputs(2621));
    layer4_outputs(1909) <= not((layer3_outputs(1229)) and (layer3_outputs(851)));
    layer4_outputs(1910) <= not(layer3_outputs(3651)) or (layer3_outputs(1629));
    layer4_outputs(1911) <= (layer3_outputs(4608)) and not (layer3_outputs(3830));
    layer4_outputs(1912) <= layer3_outputs(3564);
    layer4_outputs(1913) <= not((layer3_outputs(120)) or (layer3_outputs(2038)));
    layer4_outputs(1914) <= not((layer3_outputs(1026)) xor (layer3_outputs(4282)));
    layer4_outputs(1915) <= layer3_outputs(2262);
    layer4_outputs(1916) <= '0';
    layer4_outputs(1917) <= (layer3_outputs(4625)) and (layer3_outputs(3179));
    layer4_outputs(1918) <= '1';
    layer4_outputs(1919) <= not((layer3_outputs(1907)) and (layer3_outputs(527)));
    layer4_outputs(1920) <= not((layer3_outputs(4710)) or (layer3_outputs(4555)));
    layer4_outputs(1921) <= not(layer3_outputs(4295));
    layer4_outputs(1922) <= not((layer3_outputs(2181)) or (layer3_outputs(4419)));
    layer4_outputs(1923) <= not(layer3_outputs(3182)) or (layer3_outputs(3637));
    layer4_outputs(1924) <= not(layer3_outputs(4990)) or (layer3_outputs(3854));
    layer4_outputs(1925) <= layer3_outputs(3497);
    layer4_outputs(1926) <= '0';
    layer4_outputs(1927) <= (layer3_outputs(1593)) or (layer3_outputs(2319));
    layer4_outputs(1928) <= '0';
    layer4_outputs(1929) <= not(layer3_outputs(4930)) or (layer3_outputs(1377));
    layer4_outputs(1930) <= (layer3_outputs(1279)) and not (layer3_outputs(284));
    layer4_outputs(1931) <= '0';
    layer4_outputs(1932) <= layer3_outputs(2653);
    layer4_outputs(1933) <= not((layer3_outputs(4320)) and (layer3_outputs(4753)));
    layer4_outputs(1934) <= (layer3_outputs(3448)) or (layer3_outputs(880));
    layer4_outputs(1935) <= not(layer3_outputs(294)) or (layer3_outputs(2258));
    layer4_outputs(1936) <= layer3_outputs(3897);
    layer4_outputs(1937) <= layer3_outputs(220);
    layer4_outputs(1938) <= not(layer3_outputs(3045));
    layer4_outputs(1939) <= not(layer3_outputs(1485));
    layer4_outputs(1940) <= '0';
    layer4_outputs(1941) <= layer3_outputs(505);
    layer4_outputs(1942) <= (layer3_outputs(4228)) xor (layer3_outputs(4344));
    layer4_outputs(1943) <= not(layer3_outputs(2063)) or (layer3_outputs(638));
    layer4_outputs(1944) <= not(layer3_outputs(1760));
    layer4_outputs(1945) <= not(layer3_outputs(4100));
    layer4_outputs(1946) <= not((layer3_outputs(1468)) or (layer3_outputs(1060)));
    layer4_outputs(1947) <= not((layer3_outputs(2980)) and (layer3_outputs(3848)));
    layer4_outputs(1948) <= layer3_outputs(2706);
    layer4_outputs(1949) <= (layer3_outputs(666)) and (layer3_outputs(1573));
    layer4_outputs(1950) <= layer3_outputs(1941);
    layer4_outputs(1951) <= not((layer3_outputs(3328)) or (layer3_outputs(576)));
    layer4_outputs(1952) <= not(layer3_outputs(2681));
    layer4_outputs(1953) <= not(layer3_outputs(479));
    layer4_outputs(1954) <= layer3_outputs(4738);
    layer4_outputs(1955) <= (layer3_outputs(2985)) and not (layer3_outputs(3342));
    layer4_outputs(1956) <= not(layer3_outputs(670)) or (layer3_outputs(4051));
    layer4_outputs(1957) <= '1';
    layer4_outputs(1958) <= layer3_outputs(2488);
    layer4_outputs(1959) <= '0';
    layer4_outputs(1960) <= layer3_outputs(2158);
    layer4_outputs(1961) <= not(layer3_outputs(3078));
    layer4_outputs(1962) <= layer3_outputs(4635);
    layer4_outputs(1963) <= not((layer3_outputs(1825)) or (layer3_outputs(1122)));
    layer4_outputs(1964) <= '1';
    layer4_outputs(1965) <= (layer3_outputs(682)) and not (layer3_outputs(3925));
    layer4_outputs(1966) <= (layer3_outputs(1188)) xor (layer3_outputs(1165));
    layer4_outputs(1967) <= not((layer3_outputs(4746)) and (layer3_outputs(3824)));
    layer4_outputs(1968) <= not(layer3_outputs(3928)) or (layer3_outputs(3378));
    layer4_outputs(1969) <= not(layer3_outputs(489));
    layer4_outputs(1970) <= (layer3_outputs(2454)) and (layer3_outputs(3669));
    layer4_outputs(1971) <= (layer3_outputs(1262)) and (layer3_outputs(1860));
    layer4_outputs(1972) <= not(layer3_outputs(5016));
    layer4_outputs(1973) <= layer3_outputs(124);
    layer4_outputs(1974) <= (layer3_outputs(2585)) and not (layer3_outputs(1496));
    layer4_outputs(1975) <= (layer3_outputs(4152)) and not (layer3_outputs(118));
    layer4_outputs(1976) <= not(layer3_outputs(3036)) or (layer3_outputs(2808));
    layer4_outputs(1977) <= not(layer3_outputs(1633));
    layer4_outputs(1978) <= (layer3_outputs(4519)) and not (layer3_outputs(1392));
    layer4_outputs(1979) <= not(layer3_outputs(3486)) or (layer3_outputs(3796));
    layer4_outputs(1980) <= layer3_outputs(3755);
    layer4_outputs(1981) <= not(layer3_outputs(2405)) or (layer3_outputs(3611));
    layer4_outputs(1982) <= '0';
    layer4_outputs(1983) <= '0';
    layer4_outputs(1984) <= not(layer3_outputs(4696));
    layer4_outputs(1985) <= '0';
    layer4_outputs(1986) <= layer3_outputs(809);
    layer4_outputs(1987) <= not(layer3_outputs(4876));
    layer4_outputs(1988) <= (layer3_outputs(1852)) and (layer3_outputs(3565));
    layer4_outputs(1989) <= (layer3_outputs(523)) and (layer3_outputs(1673));
    layer4_outputs(1990) <= not((layer3_outputs(4616)) or (layer3_outputs(45)));
    layer4_outputs(1991) <= not(layer3_outputs(3342));
    layer4_outputs(1992) <= layer3_outputs(4084);
    layer4_outputs(1993) <= not((layer3_outputs(2069)) xor (layer3_outputs(456)));
    layer4_outputs(1994) <= layer3_outputs(619);
    layer4_outputs(1995) <= not(layer3_outputs(2729)) or (layer3_outputs(799));
    layer4_outputs(1996) <= layer3_outputs(1193);
    layer4_outputs(1997) <= not(layer3_outputs(2101));
    layer4_outputs(1998) <= '0';
    layer4_outputs(1999) <= layer3_outputs(253);
    layer4_outputs(2000) <= not((layer3_outputs(58)) or (layer3_outputs(3758)));
    layer4_outputs(2001) <= (layer3_outputs(2906)) and not (layer3_outputs(4692));
    layer4_outputs(2002) <= (layer3_outputs(1417)) and (layer3_outputs(3131));
    layer4_outputs(2003) <= (layer3_outputs(5027)) and not (layer3_outputs(3316));
    layer4_outputs(2004) <= not(layer3_outputs(2022)) or (layer3_outputs(2700));
    layer4_outputs(2005) <= (layer3_outputs(4554)) and not (layer3_outputs(5020));
    layer4_outputs(2006) <= not(layer3_outputs(4936));
    layer4_outputs(2007) <= not(layer3_outputs(2702));
    layer4_outputs(2008) <= (layer3_outputs(1237)) or (layer3_outputs(1713));
    layer4_outputs(2009) <= (layer3_outputs(2877)) or (layer3_outputs(1531));
    layer4_outputs(2010) <= '1';
    layer4_outputs(2011) <= '0';
    layer4_outputs(2012) <= layer3_outputs(3150);
    layer4_outputs(2013) <= not(layer3_outputs(1052));
    layer4_outputs(2014) <= (layer3_outputs(417)) and not (layer3_outputs(2031));
    layer4_outputs(2015) <= '0';
    layer4_outputs(2016) <= (layer3_outputs(62)) or (layer3_outputs(474));
    layer4_outputs(2017) <= layer3_outputs(4972);
    layer4_outputs(2018) <= not(layer3_outputs(2007)) or (layer3_outputs(4339));
    layer4_outputs(2019) <= not(layer3_outputs(2165));
    layer4_outputs(2020) <= not((layer3_outputs(2324)) and (layer3_outputs(2389)));
    layer4_outputs(2021) <= '0';
    layer4_outputs(2022) <= not(layer3_outputs(3887));
    layer4_outputs(2023) <= not((layer3_outputs(699)) or (layer3_outputs(1464)));
    layer4_outputs(2024) <= layer3_outputs(5014);
    layer4_outputs(2025) <= (layer3_outputs(1765)) or (layer3_outputs(3411));
    layer4_outputs(2026) <= (layer3_outputs(4412)) and not (layer3_outputs(262));
    layer4_outputs(2027) <= (layer3_outputs(583)) and (layer3_outputs(4893));
    layer4_outputs(2028) <= not(layer3_outputs(3780)) or (layer3_outputs(1336));
    layer4_outputs(2029) <= not((layer3_outputs(3334)) or (layer3_outputs(1390)));
    layer4_outputs(2030) <= not((layer3_outputs(4717)) and (layer3_outputs(157)));
    layer4_outputs(2031) <= not(layer3_outputs(2412));
    layer4_outputs(2032) <= not(layer3_outputs(4935));
    layer4_outputs(2033) <= layer3_outputs(4793);
    layer4_outputs(2034) <= not((layer3_outputs(1609)) or (layer3_outputs(2505)));
    layer4_outputs(2035) <= not((layer3_outputs(3601)) and (layer3_outputs(4181)));
    layer4_outputs(2036) <= not(layer3_outputs(3204)) or (layer3_outputs(4467));
    layer4_outputs(2037) <= not(layer3_outputs(4166)) or (layer3_outputs(226));
    layer4_outputs(2038) <= layer3_outputs(4563);
    layer4_outputs(2039) <= layer3_outputs(3195);
    layer4_outputs(2040) <= layer3_outputs(2796);
    layer4_outputs(2041) <= layer3_outputs(1077);
    layer4_outputs(2042) <= (layer3_outputs(4636)) and not (layer3_outputs(1240));
    layer4_outputs(2043) <= layer3_outputs(712);
    layer4_outputs(2044) <= not(layer3_outputs(3717)) or (layer3_outputs(3631));
    layer4_outputs(2045) <= '1';
    layer4_outputs(2046) <= (layer3_outputs(4597)) or (layer3_outputs(320));
    layer4_outputs(2047) <= (layer3_outputs(927)) and (layer3_outputs(3418));
    layer4_outputs(2048) <= not(layer3_outputs(64)) or (layer3_outputs(3985));
    layer4_outputs(2049) <= not(layer3_outputs(3717)) or (layer3_outputs(987));
    layer4_outputs(2050) <= not(layer3_outputs(3219)) or (layer3_outputs(1718));
    layer4_outputs(2051) <= not((layer3_outputs(1129)) and (layer3_outputs(3832)));
    layer4_outputs(2052) <= not(layer3_outputs(1407));
    layer4_outputs(2053) <= layer3_outputs(12);
    layer4_outputs(2054) <= not(layer3_outputs(4267));
    layer4_outputs(2055) <= not((layer3_outputs(287)) and (layer3_outputs(714)));
    layer4_outputs(2056) <= (layer3_outputs(4693)) and not (layer3_outputs(937));
    layer4_outputs(2057) <= not(layer3_outputs(1050));
    layer4_outputs(2058) <= layer3_outputs(1161);
    layer4_outputs(2059) <= not(layer3_outputs(3914));
    layer4_outputs(2060) <= (layer3_outputs(3560)) or (layer3_outputs(4698));
    layer4_outputs(2061) <= not(layer3_outputs(4224));
    layer4_outputs(2062) <= (layer3_outputs(3989)) or (layer3_outputs(1532));
    layer4_outputs(2063) <= (layer3_outputs(972)) and not (layer3_outputs(3705));
    layer4_outputs(2064) <= layer3_outputs(869);
    layer4_outputs(2065) <= not(layer3_outputs(3565));
    layer4_outputs(2066) <= layer3_outputs(4129);
    layer4_outputs(2067) <= (layer3_outputs(1853)) and (layer3_outputs(4826));
    layer4_outputs(2068) <= not(layer3_outputs(1740));
    layer4_outputs(2069) <= layer3_outputs(2474);
    layer4_outputs(2070) <= '1';
    layer4_outputs(2071) <= not(layer3_outputs(1880));
    layer4_outputs(2072) <= not((layer3_outputs(1025)) and (layer3_outputs(744)));
    layer4_outputs(2073) <= (layer3_outputs(422)) and not (layer3_outputs(900));
    layer4_outputs(2074) <= (layer3_outputs(292)) and not (layer3_outputs(4535));
    layer4_outputs(2075) <= not((layer3_outputs(137)) xor (layer3_outputs(1802)));
    layer4_outputs(2076) <= not(layer3_outputs(4656)) or (layer3_outputs(423));
    layer4_outputs(2077) <= not(layer3_outputs(3176)) or (layer3_outputs(1222));
    layer4_outputs(2078) <= (layer3_outputs(456)) xor (layer3_outputs(2425));
    layer4_outputs(2079) <= (layer3_outputs(3299)) and not (layer3_outputs(3211));
    layer4_outputs(2080) <= not(layer3_outputs(4284));
    layer4_outputs(2081) <= layer3_outputs(2282);
    layer4_outputs(2082) <= (layer3_outputs(4842)) and not (layer3_outputs(1036));
    layer4_outputs(2083) <= not(layer3_outputs(4156));
    layer4_outputs(2084) <= layer3_outputs(308);
    layer4_outputs(2085) <= (layer3_outputs(3706)) and not (layer3_outputs(2564));
    layer4_outputs(2086) <= not(layer3_outputs(4759));
    layer4_outputs(2087) <= layer3_outputs(88);
    layer4_outputs(2088) <= layer3_outputs(521);
    layer4_outputs(2089) <= not(layer3_outputs(2191)) or (layer3_outputs(1872));
    layer4_outputs(2090) <= layer3_outputs(4485);
    layer4_outputs(2091) <= (layer3_outputs(5051)) or (layer3_outputs(519));
    layer4_outputs(2092) <= not(layer3_outputs(4259)) or (layer3_outputs(3286));
    layer4_outputs(2093) <= layer3_outputs(3899);
    layer4_outputs(2094) <= not(layer3_outputs(1418)) or (layer3_outputs(4068));
    layer4_outputs(2095) <= layer3_outputs(4750);
    layer4_outputs(2096) <= '1';
    layer4_outputs(2097) <= layer3_outputs(1805);
    layer4_outputs(2098) <= (layer3_outputs(1489)) or (layer3_outputs(3489));
    layer4_outputs(2099) <= not(layer3_outputs(2099)) or (layer3_outputs(3049));
    layer4_outputs(2100) <= not(layer3_outputs(3310));
    layer4_outputs(2101) <= not(layer3_outputs(4561)) or (layer3_outputs(2085));
    layer4_outputs(2102) <= layer3_outputs(5038);
    layer4_outputs(2103) <= layer3_outputs(3621);
    layer4_outputs(2104) <= layer3_outputs(150);
    layer4_outputs(2105) <= (layer3_outputs(4021)) and not (layer3_outputs(4234));
    layer4_outputs(2106) <= not(layer3_outputs(4285)) or (layer3_outputs(1870));
    layer4_outputs(2107) <= (layer3_outputs(3016)) xor (layer3_outputs(1584));
    layer4_outputs(2108) <= (layer3_outputs(1428)) and (layer3_outputs(4078));
    layer4_outputs(2109) <= (layer3_outputs(762)) and not (layer3_outputs(276));
    layer4_outputs(2110) <= (layer3_outputs(1971)) and not (layer3_outputs(1551));
    layer4_outputs(2111) <= not(layer3_outputs(1136));
    layer4_outputs(2112) <= not((layer3_outputs(254)) and (layer3_outputs(2012)));
    layer4_outputs(2113) <= not((layer3_outputs(5015)) or (layer3_outputs(2594)));
    layer4_outputs(2114) <= not(layer3_outputs(3844)) or (layer3_outputs(3711));
    layer4_outputs(2115) <= not((layer3_outputs(3366)) or (layer3_outputs(1350)));
    layer4_outputs(2116) <= not(layer3_outputs(3772));
    layer4_outputs(2117) <= not(layer3_outputs(4748));
    layer4_outputs(2118) <= layer3_outputs(1492);
    layer4_outputs(2119) <= not(layer3_outputs(3734));
    layer4_outputs(2120) <= not(layer3_outputs(499));
    layer4_outputs(2121) <= (layer3_outputs(4005)) and not (layer3_outputs(218));
    layer4_outputs(2122) <= layer3_outputs(3909);
    layer4_outputs(2123) <= not(layer3_outputs(167)) or (layer3_outputs(4161));
    layer4_outputs(2124) <= not((layer3_outputs(2385)) or (layer3_outputs(2280)));
    layer4_outputs(2125) <= not(layer3_outputs(1233)) or (layer3_outputs(4467));
    layer4_outputs(2126) <= (layer3_outputs(411)) and not (layer3_outputs(4851));
    layer4_outputs(2127) <= '0';
    layer4_outputs(2128) <= (layer3_outputs(1163)) or (layer3_outputs(2993));
    layer4_outputs(2129) <= '0';
    layer4_outputs(2130) <= (layer3_outputs(4426)) or (layer3_outputs(1243));
    layer4_outputs(2131) <= not((layer3_outputs(1493)) and (layer3_outputs(3435)));
    layer4_outputs(2132) <= not(layer3_outputs(2866));
    layer4_outputs(2133) <= '1';
    layer4_outputs(2134) <= '1';
    layer4_outputs(2135) <= layer3_outputs(3380);
    layer4_outputs(2136) <= (layer3_outputs(4817)) and (layer3_outputs(2473));
    layer4_outputs(2137) <= not(layer3_outputs(1538)) or (layer3_outputs(4216));
    layer4_outputs(2138) <= not(layer3_outputs(4061)) or (layer3_outputs(227));
    layer4_outputs(2139) <= not((layer3_outputs(3302)) or (layer3_outputs(1890)));
    layer4_outputs(2140) <= '0';
    layer4_outputs(2141) <= not(layer3_outputs(1526));
    layer4_outputs(2142) <= (layer3_outputs(2017)) and not (layer3_outputs(3122));
    layer4_outputs(2143) <= not(layer3_outputs(2446));
    layer4_outputs(2144) <= '0';
    layer4_outputs(2145) <= not(layer3_outputs(3546));
    layer4_outputs(2146) <= (layer3_outputs(3500)) and (layer3_outputs(4859));
    layer4_outputs(2147) <= layer3_outputs(3106);
    layer4_outputs(2148) <= layer3_outputs(610);
    layer4_outputs(2149) <= not((layer3_outputs(5107)) or (layer3_outputs(4472)));
    layer4_outputs(2150) <= '1';
    layer4_outputs(2151) <= not((layer3_outputs(1494)) and (layer3_outputs(2736)));
    layer4_outputs(2152) <= layer3_outputs(2956);
    layer4_outputs(2153) <= not((layer3_outputs(3359)) or (layer3_outputs(3148)));
    layer4_outputs(2154) <= layer3_outputs(3945);
    layer4_outputs(2155) <= (layer3_outputs(1649)) and not (layer3_outputs(2129));
    layer4_outputs(2156) <= (layer3_outputs(3280)) and not (layer3_outputs(713));
    layer4_outputs(2157) <= (layer3_outputs(3994)) or (layer3_outputs(2141));
    layer4_outputs(2158) <= not(layer3_outputs(3018)) or (layer3_outputs(3266));
    layer4_outputs(2159) <= not(layer3_outputs(1372)) or (layer3_outputs(3746));
    layer4_outputs(2160) <= not(layer3_outputs(1918));
    layer4_outputs(2161) <= (layer3_outputs(187)) and not (layer3_outputs(1540));
    layer4_outputs(2162) <= '0';
    layer4_outputs(2163) <= (layer3_outputs(4831)) and (layer3_outputs(2372));
    layer4_outputs(2164) <= layer3_outputs(4715);
    layer4_outputs(2165) <= not(layer3_outputs(2166)) or (layer3_outputs(4074));
    layer4_outputs(2166) <= layer3_outputs(1744);
    layer4_outputs(2167) <= not(layer3_outputs(2252));
    layer4_outputs(2168) <= not(layer3_outputs(4488));
    layer4_outputs(2169) <= (layer3_outputs(2131)) and (layer3_outputs(1911));
    layer4_outputs(2170) <= not(layer3_outputs(222));
    layer4_outputs(2171) <= not(layer3_outputs(4206)) or (layer3_outputs(2654));
    layer4_outputs(2172) <= '0';
    layer4_outputs(2173) <= layer3_outputs(2643);
    layer4_outputs(2174) <= not((layer3_outputs(905)) or (layer3_outputs(4247)));
    layer4_outputs(2175) <= (layer3_outputs(3234)) and not (layer3_outputs(276));
    layer4_outputs(2176) <= not(layer3_outputs(3596)) or (layer3_outputs(715));
    layer4_outputs(2177) <= not(layer3_outputs(2133));
    layer4_outputs(2178) <= '0';
    layer4_outputs(2179) <= layer3_outputs(369);
    layer4_outputs(2180) <= (layer3_outputs(3156)) and (layer3_outputs(1958));
    layer4_outputs(2181) <= not((layer3_outputs(2778)) or (layer3_outputs(3666)));
    layer4_outputs(2182) <= not(layer3_outputs(3058));
    layer4_outputs(2183) <= not((layer3_outputs(2644)) and (layer3_outputs(3555)));
    layer4_outputs(2184) <= not(layer3_outputs(840)) or (layer3_outputs(3165));
    layer4_outputs(2185) <= not((layer3_outputs(3970)) and (layer3_outputs(849)));
    layer4_outputs(2186) <= (layer3_outputs(2009)) or (layer3_outputs(2862));
    layer4_outputs(2187) <= '1';
    layer4_outputs(2188) <= not(layer3_outputs(1341)) or (layer3_outputs(4229));
    layer4_outputs(2189) <= not(layer3_outputs(1329));
    layer4_outputs(2190) <= not((layer3_outputs(3828)) or (layer3_outputs(1348)));
    layer4_outputs(2191) <= (layer3_outputs(5112)) xor (layer3_outputs(4253));
    layer4_outputs(2192) <= not(layer3_outputs(230));
    layer4_outputs(2193) <= not(layer3_outputs(1963));
    layer4_outputs(2194) <= (layer3_outputs(4768)) or (layer3_outputs(2647));
    layer4_outputs(2195) <= not((layer3_outputs(3473)) or (layer3_outputs(3416)));
    layer4_outputs(2196) <= (layer3_outputs(1767)) or (layer3_outputs(265));
    layer4_outputs(2197) <= not(layer3_outputs(310));
    layer4_outputs(2198) <= '0';
    layer4_outputs(2199) <= not((layer3_outputs(2978)) and (layer3_outputs(2525)));
    layer4_outputs(2200) <= not(layer3_outputs(855));
    layer4_outputs(2201) <= not(layer3_outputs(933)) or (layer3_outputs(3604));
    layer4_outputs(2202) <= not(layer3_outputs(3733));
    layer4_outputs(2203) <= not(layer3_outputs(2997)) or (layer3_outputs(2140));
    layer4_outputs(2204) <= (layer3_outputs(4541)) and not (layer3_outputs(4436));
    layer4_outputs(2205) <= not((layer3_outputs(825)) and (layer3_outputs(3953)));
    layer4_outputs(2206) <= '0';
    layer4_outputs(2207) <= not((layer3_outputs(2573)) and (layer3_outputs(4242)));
    layer4_outputs(2208) <= not(layer3_outputs(4311)) or (layer3_outputs(2183));
    layer4_outputs(2209) <= layer3_outputs(3155);
    layer4_outputs(2210) <= not(layer3_outputs(1601)) or (layer3_outputs(3509));
    layer4_outputs(2211) <= '1';
    layer4_outputs(2212) <= not(layer3_outputs(4980));
    layer4_outputs(2213) <= not(layer3_outputs(4410));
    layer4_outputs(2214) <= not(layer3_outputs(1314)) or (layer3_outputs(36));
    layer4_outputs(2215) <= not((layer3_outputs(5064)) xor (layer3_outputs(878)));
    layer4_outputs(2216) <= not(layer3_outputs(2358));
    layer4_outputs(2217) <= not(layer3_outputs(3856));
    layer4_outputs(2218) <= layer3_outputs(3922);
    layer4_outputs(2219) <= (layer3_outputs(4808)) or (layer3_outputs(4848));
    layer4_outputs(2220) <= '1';
    layer4_outputs(2221) <= '0';
    layer4_outputs(2222) <= (layer3_outputs(2881)) and (layer3_outputs(1083));
    layer4_outputs(2223) <= not((layer3_outputs(450)) and (layer3_outputs(1910)));
    layer4_outputs(2224) <= (layer3_outputs(2002)) or (layer3_outputs(1906));
    layer4_outputs(2225) <= not(layer3_outputs(2837)) or (layer3_outputs(3228));
    layer4_outputs(2226) <= (layer3_outputs(2098)) xor (layer3_outputs(4497));
    layer4_outputs(2227) <= (layer3_outputs(607)) and (layer3_outputs(2448));
    layer4_outputs(2228) <= layer3_outputs(5087);
    layer4_outputs(2229) <= not((layer3_outputs(464)) or (layer3_outputs(4689)));
    layer4_outputs(2230) <= not(layer3_outputs(2672));
    layer4_outputs(2231) <= not(layer3_outputs(4908)) or (layer3_outputs(259));
    layer4_outputs(2232) <= '1';
    layer4_outputs(2233) <= layer3_outputs(1510);
    layer4_outputs(2234) <= not(layer3_outputs(534)) or (layer3_outputs(888));
    layer4_outputs(2235) <= not(layer3_outputs(2260));
    layer4_outputs(2236) <= (layer3_outputs(2281)) and not (layer3_outputs(84));
    layer4_outputs(2237) <= (layer3_outputs(1184)) and not (layer3_outputs(3868));
    layer4_outputs(2238) <= (layer3_outputs(3998)) and not (layer3_outputs(3065));
    layer4_outputs(2239) <= (layer3_outputs(4286)) and not (layer3_outputs(3955));
    layer4_outputs(2240) <= not(layer3_outputs(1704)) or (layer3_outputs(267));
    layer4_outputs(2241) <= layer3_outputs(1192);
    layer4_outputs(2242) <= layer3_outputs(427);
    layer4_outputs(2243) <= not(layer3_outputs(2631));
    layer4_outputs(2244) <= not((layer3_outputs(4742)) or (layer3_outputs(2917)));
    layer4_outputs(2245) <= (layer3_outputs(2781)) and not (layer3_outputs(618));
    layer4_outputs(2246) <= layer3_outputs(735);
    layer4_outputs(2247) <= '1';
    layer4_outputs(2248) <= (layer3_outputs(4803)) and not (layer3_outputs(1109));
    layer4_outputs(2249) <= not((layer3_outputs(3657)) or (layer3_outputs(3548)));
    layer4_outputs(2250) <= '1';
    layer4_outputs(2251) <= '1';
    layer4_outputs(2252) <= '1';
    layer4_outputs(2253) <= layer3_outputs(313);
    layer4_outputs(2254) <= layer3_outputs(3173);
    layer4_outputs(2255) <= (layer3_outputs(4968)) or (layer3_outputs(786));
    layer4_outputs(2256) <= (layer3_outputs(4630)) and (layer3_outputs(3307));
    layer4_outputs(2257) <= not(layer3_outputs(477));
    layer4_outputs(2258) <= (layer3_outputs(3027)) and not (layer3_outputs(533));
    layer4_outputs(2259) <= not(layer3_outputs(4131)) or (layer3_outputs(2040));
    layer4_outputs(2260) <= not(layer3_outputs(1404)) or (layer3_outputs(4775));
    layer4_outputs(2261) <= not((layer3_outputs(2090)) xor (layer3_outputs(835)));
    layer4_outputs(2262) <= not(layer3_outputs(2914));
    layer4_outputs(2263) <= (layer3_outputs(1536)) and not (layer3_outputs(2410));
    layer4_outputs(2264) <= (layer3_outputs(4096)) or (layer3_outputs(3278));
    layer4_outputs(2265) <= (layer3_outputs(2874)) and (layer3_outputs(4219));
    layer4_outputs(2266) <= (layer3_outputs(4389)) and (layer3_outputs(3912));
    layer4_outputs(2267) <= (layer3_outputs(603)) or (layer3_outputs(446));
    layer4_outputs(2268) <= (layer3_outputs(4910)) or (layer3_outputs(297));
    layer4_outputs(2269) <= '1';
    layer4_outputs(2270) <= layer3_outputs(3603);
    layer4_outputs(2271) <= (layer3_outputs(1162)) and not (layer3_outputs(4567));
    layer4_outputs(2272) <= not(layer3_outputs(105));
    layer4_outputs(2273) <= '1';
    layer4_outputs(2274) <= not(layer3_outputs(1557));
    layer4_outputs(2275) <= (layer3_outputs(1102)) and not (layer3_outputs(4906));
    layer4_outputs(2276) <= layer3_outputs(286);
    layer4_outputs(2277) <= not((layer3_outputs(4998)) and (layer3_outputs(918)));
    layer4_outputs(2278) <= not(layer3_outputs(4982));
    layer4_outputs(2279) <= not((layer3_outputs(3312)) and (layer3_outputs(1808)));
    layer4_outputs(2280) <= not((layer3_outputs(1486)) and (layer3_outputs(5017)));
    layer4_outputs(2281) <= '1';
    layer4_outputs(2282) <= (layer3_outputs(4048)) and not (layer3_outputs(2546));
    layer4_outputs(2283) <= '0';
    layer4_outputs(2284) <= not((layer3_outputs(1599)) or (layer3_outputs(3255)));
    layer4_outputs(2285) <= layer3_outputs(2468);
    layer4_outputs(2286) <= layer3_outputs(3602);
    layer4_outputs(2287) <= not((layer3_outputs(703)) or (layer3_outputs(2604)));
    layer4_outputs(2288) <= not(layer3_outputs(3558));
    layer4_outputs(2289) <= layer3_outputs(2532);
    layer4_outputs(2290) <= not(layer3_outputs(4682)) or (layer3_outputs(3686));
    layer4_outputs(2291) <= not(layer3_outputs(488)) or (layer3_outputs(1835));
    layer4_outputs(2292) <= not(layer3_outputs(955));
    layer4_outputs(2293) <= (layer3_outputs(1300)) and not (layer3_outputs(4004));
    layer4_outputs(2294) <= (layer3_outputs(1871)) or (layer3_outputs(1254));
    layer4_outputs(2295) <= (layer3_outputs(310)) and (layer3_outputs(1831));
    layer4_outputs(2296) <= (layer3_outputs(38)) and (layer3_outputs(3749));
    layer4_outputs(2297) <= not(layer3_outputs(4196)) or (layer3_outputs(4644));
    layer4_outputs(2298) <= not(layer3_outputs(944)) or (layer3_outputs(4089));
    layer4_outputs(2299) <= not(layer3_outputs(1428)) or (layer3_outputs(405));
    layer4_outputs(2300) <= not(layer3_outputs(1244));
    layer4_outputs(2301) <= (layer3_outputs(886)) or (layer3_outputs(4800));
    layer4_outputs(2302) <= not((layer3_outputs(4385)) or (layer3_outputs(2062)));
    layer4_outputs(2303) <= '1';
    layer4_outputs(2304) <= (layer3_outputs(1442)) and (layer3_outputs(4719));
    layer4_outputs(2305) <= layer3_outputs(1420);
    layer4_outputs(2306) <= (layer3_outputs(4534)) and (layer3_outputs(1936));
    layer4_outputs(2307) <= '1';
    layer4_outputs(2308) <= (layer3_outputs(2313)) and not (layer3_outputs(4662));
    layer4_outputs(2309) <= (layer3_outputs(3563)) or (layer3_outputs(1605));
    layer4_outputs(2310) <= not((layer3_outputs(144)) and (layer3_outputs(4357)));
    layer4_outputs(2311) <= not((layer3_outputs(2321)) and (layer3_outputs(5012)));
    layer4_outputs(2312) <= not((layer3_outputs(4423)) and (layer3_outputs(3128)));
    layer4_outputs(2313) <= not(layer3_outputs(1258)) or (layer3_outputs(3892));
    layer4_outputs(2314) <= (layer3_outputs(1280)) and not (layer3_outputs(3613));
    layer4_outputs(2315) <= layer3_outputs(2102);
    layer4_outputs(2316) <= '1';
    layer4_outputs(2317) <= not(layer3_outputs(3860)) or (layer3_outputs(3572));
    layer4_outputs(2318) <= '1';
    layer4_outputs(2319) <= layer3_outputs(2075);
    layer4_outputs(2320) <= not((layer3_outputs(5119)) and (layer3_outputs(403)));
    layer4_outputs(2321) <= (layer3_outputs(3219)) and not (layer3_outputs(1115));
    layer4_outputs(2322) <= (layer3_outputs(2152)) and (layer3_outputs(2823));
    layer4_outputs(2323) <= not(layer3_outputs(1100));
    layer4_outputs(2324) <= not((layer3_outputs(3486)) and (layer3_outputs(4743)));
    layer4_outputs(2325) <= (layer3_outputs(2277)) and (layer3_outputs(671));
    layer4_outputs(2326) <= layer3_outputs(820);
    layer4_outputs(2327) <= layer3_outputs(3989);
    layer4_outputs(2328) <= (layer3_outputs(4916)) and not (layer3_outputs(2154));
    layer4_outputs(2329) <= '0';
    layer4_outputs(2330) <= layer3_outputs(4747);
    layer4_outputs(2331) <= not((layer3_outputs(899)) or (layer3_outputs(4786)));
    layer4_outputs(2332) <= '1';
    layer4_outputs(2333) <= not((layer3_outputs(658)) or (layer3_outputs(4907)));
    layer4_outputs(2334) <= not(layer3_outputs(438)) or (layer3_outputs(2932));
    layer4_outputs(2335) <= layer3_outputs(4009);
    layer4_outputs(2336) <= not(layer3_outputs(3788)) or (layer3_outputs(2023));
    layer4_outputs(2337) <= (layer3_outputs(3302)) and not (layer3_outputs(2501));
    layer4_outputs(2338) <= not(layer3_outputs(2227)) or (layer3_outputs(3283));
    layer4_outputs(2339) <= not(layer3_outputs(733)) or (layer3_outputs(4448));
    layer4_outputs(2340) <= (layer3_outputs(946)) xor (layer3_outputs(1762));
    layer4_outputs(2341) <= '1';
    layer4_outputs(2342) <= '1';
    layer4_outputs(2343) <= not(layer3_outputs(3789));
    layer4_outputs(2344) <= not(layer3_outputs(1085));
    layer4_outputs(2345) <= '1';
    layer4_outputs(2346) <= (layer3_outputs(4573)) and (layer3_outputs(797));
    layer4_outputs(2347) <= layer3_outputs(2231);
    layer4_outputs(2348) <= (layer3_outputs(1550)) and not (layer3_outputs(737));
    layer4_outputs(2349) <= not((layer3_outputs(4301)) and (layer3_outputs(1838)));
    layer4_outputs(2350) <= '0';
    layer4_outputs(2351) <= (layer3_outputs(4959)) and not (layer3_outputs(1898));
    layer4_outputs(2352) <= layer3_outputs(2064);
    layer4_outputs(2353) <= (layer3_outputs(2800)) and not (layer3_outputs(4069));
    layer4_outputs(2354) <= (layer3_outputs(5113)) and not (layer3_outputs(3564));
    layer4_outputs(2355) <= '1';
    layer4_outputs(2356) <= not((layer3_outputs(496)) and (layer3_outputs(4331)));
    layer4_outputs(2357) <= '0';
    layer4_outputs(2358) <= (layer3_outputs(1750)) and (layer3_outputs(2629));
    layer4_outputs(2359) <= (layer3_outputs(1121)) or (layer3_outputs(224));
    layer4_outputs(2360) <= layer3_outputs(5089);
    layer4_outputs(2361) <= '1';
    layer4_outputs(2362) <= (layer3_outputs(2410)) and (layer3_outputs(803));
    layer4_outputs(2363) <= not((layer3_outputs(751)) and (layer3_outputs(997)));
    layer4_outputs(2364) <= (layer3_outputs(4695)) and not (layer3_outputs(628));
    layer4_outputs(2365) <= not(layer3_outputs(3528)) or (layer3_outputs(3058));
    layer4_outputs(2366) <= layer3_outputs(2582);
    layer4_outputs(2367) <= (layer3_outputs(4226)) or (layer3_outputs(2873));
    layer4_outputs(2368) <= not(layer3_outputs(4077)) or (layer3_outputs(958));
    layer4_outputs(2369) <= (layer3_outputs(2037)) or (layer3_outputs(594));
    layer4_outputs(2370) <= not((layer3_outputs(1288)) and (layer3_outputs(370)));
    layer4_outputs(2371) <= not((layer3_outputs(2704)) and (layer3_outputs(4393)));
    layer4_outputs(2372) <= not(layer3_outputs(508));
    layer4_outputs(2373) <= not(layer3_outputs(3827));
    layer4_outputs(2374) <= '0';
    layer4_outputs(2375) <= (layer3_outputs(4587)) and (layer3_outputs(1086));
    layer4_outputs(2376) <= (layer3_outputs(85)) and not (layer3_outputs(2244));
    layer4_outputs(2377) <= not(layer3_outputs(1514)) or (layer3_outputs(4002));
    layer4_outputs(2378) <= (layer3_outputs(2625)) or (layer3_outputs(4478));
    layer4_outputs(2379) <= '1';
    layer4_outputs(2380) <= (layer3_outputs(3871)) and not (layer3_outputs(4135));
    layer4_outputs(2381) <= not((layer3_outputs(4894)) or (layer3_outputs(2285)));
    layer4_outputs(2382) <= layer3_outputs(1774);
    layer4_outputs(2383) <= layer3_outputs(4484);
    layer4_outputs(2384) <= (layer3_outputs(2374)) and (layer3_outputs(3884));
    layer4_outputs(2385) <= (layer3_outputs(2630)) xor (layer3_outputs(2444));
    layer4_outputs(2386) <= not(layer3_outputs(4925)) or (layer3_outputs(171));
    layer4_outputs(2387) <= not(layer3_outputs(3205)) or (layer3_outputs(1073));
    layer4_outputs(2388) <= not(layer3_outputs(1193)) or (layer3_outputs(1622));
    layer4_outputs(2389) <= (layer3_outputs(868)) and not (layer3_outputs(147));
    layer4_outputs(2390) <= (layer3_outputs(5075)) and not (layer3_outputs(2148));
    layer4_outputs(2391) <= not(layer3_outputs(252));
    layer4_outputs(2392) <= layer3_outputs(2483);
    layer4_outputs(2393) <= '1';
    layer4_outputs(2394) <= not(layer3_outputs(4341)) or (layer3_outputs(1973));
    layer4_outputs(2395) <= (layer3_outputs(2355)) and (layer3_outputs(1525));
    layer4_outputs(2396) <= layer3_outputs(4569);
    layer4_outputs(2397) <= not(layer3_outputs(5067)) or (layer3_outputs(4934));
    layer4_outputs(2398) <= not(layer3_outputs(3100));
    layer4_outputs(2399) <= '1';
    layer4_outputs(2400) <= layer3_outputs(3751);
    layer4_outputs(2401) <= layer3_outputs(2035);
    layer4_outputs(2402) <= not(layer3_outputs(890));
    layer4_outputs(2403) <= layer3_outputs(554);
    layer4_outputs(2404) <= layer3_outputs(377);
    layer4_outputs(2405) <= layer3_outputs(264);
    layer4_outputs(2406) <= layer3_outputs(4092);
    layer4_outputs(2407) <= (layer3_outputs(762)) and (layer3_outputs(3422));
    layer4_outputs(2408) <= not(layer3_outputs(4271)) or (layer3_outputs(470));
    layer4_outputs(2409) <= not((layer3_outputs(916)) or (layer3_outputs(3254)));
    layer4_outputs(2410) <= not(layer3_outputs(173));
    layer4_outputs(2411) <= not(layer3_outputs(4663)) or (layer3_outputs(846));
    layer4_outputs(2412) <= not(layer3_outputs(92));
    layer4_outputs(2413) <= '1';
    layer4_outputs(2414) <= not(layer3_outputs(2560));
    layer4_outputs(2415) <= '1';
    layer4_outputs(2416) <= layer3_outputs(4798);
    layer4_outputs(2417) <= (layer3_outputs(4980)) and (layer3_outputs(5010));
    layer4_outputs(2418) <= (layer3_outputs(1858)) or (layer3_outputs(1657));
    layer4_outputs(2419) <= not(layer3_outputs(1504));
    layer4_outputs(2420) <= (layer3_outputs(51)) and (layer3_outputs(3913));
    layer4_outputs(2421) <= (layer3_outputs(1678)) xor (layer3_outputs(3492));
    layer4_outputs(2422) <= not(layer3_outputs(819));
    layer4_outputs(2423) <= layer3_outputs(3603);
    layer4_outputs(2424) <= not(layer3_outputs(581));
    layer4_outputs(2425) <= layer3_outputs(2899);
    layer4_outputs(2426) <= not((layer3_outputs(677)) and (layer3_outputs(3490)));
    layer4_outputs(2427) <= '0';
    layer4_outputs(2428) <= layer3_outputs(3385);
    layer4_outputs(2429) <= layer3_outputs(77);
    layer4_outputs(2430) <= '1';
    layer4_outputs(2431) <= not(layer3_outputs(374)) or (layer3_outputs(46));
    layer4_outputs(2432) <= not((layer3_outputs(1159)) or (layer3_outputs(3941)));
    layer4_outputs(2433) <= (layer3_outputs(1219)) and (layer3_outputs(4571));
    layer4_outputs(2434) <= (layer3_outputs(551)) and not (layer3_outputs(1596));
    layer4_outputs(2435) <= '1';
    layer4_outputs(2436) <= layer3_outputs(676);
    layer4_outputs(2437) <= layer3_outputs(1779);
    layer4_outputs(2438) <= '1';
    layer4_outputs(2439) <= not((layer3_outputs(928)) or (layer3_outputs(4420)));
    layer4_outputs(2440) <= (layer3_outputs(630)) xor (layer3_outputs(2384));
    layer4_outputs(2441) <= not(layer3_outputs(4269));
    layer4_outputs(2442) <= not(layer3_outputs(366));
    layer4_outputs(2443) <= (layer3_outputs(1000)) and (layer3_outputs(2965));
    layer4_outputs(2444) <= layer3_outputs(848);
    layer4_outputs(2445) <= (layer3_outputs(4324)) or (layer3_outputs(3269));
    layer4_outputs(2446) <= not((layer3_outputs(2360)) and (layer3_outputs(2406)));
    layer4_outputs(2447) <= (layer3_outputs(2310)) and (layer3_outputs(1299));
    layer4_outputs(2448) <= not(layer3_outputs(5046));
    layer4_outputs(2449) <= (layer3_outputs(2039)) or (layer3_outputs(1552));
    layer4_outputs(2450) <= not(layer3_outputs(3797));
    layer4_outputs(2451) <= (layer3_outputs(4695)) and not (layer3_outputs(726));
    layer4_outputs(2452) <= '1';
    layer4_outputs(2453) <= not((layer3_outputs(4345)) or (layer3_outputs(5086)));
    layer4_outputs(2454) <= not(layer3_outputs(4528)) or (layer3_outputs(4326));
    layer4_outputs(2455) <= '0';
    layer4_outputs(2456) <= not(layer3_outputs(1821));
    layer4_outputs(2457) <= not((layer3_outputs(2759)) xor (layer3_outputs(1639)));
    layer4_outputs(2458) <= (layer3_outputs(2332)) or (layer3_outputs(3049));
    layer4_outputs(2459) <= layer3_outputs(1981);
    layer4_outputs(2460) <= not(layer3_outputs(968));
    layer4_outputs(2461) <= not((layer3_outputs(2931)) xor (layer3_outputs(4472)));
    layer4_outputs(2462) <= not((layer3_outputs(3060)) and (layer3_outputs(4139)));
    layer4_outputs(2463) <= not((layer3_outputs(2534)) or (layer3_outputs(3619)));
    layer4_outputs(2464) <= not(layer3_outputs(1572));
    layer4_outputs(2465) <= not(layer3_outputs(4444));
    layer4_outputs(2466) <= (layer3_outputs(1844)) or (layer3_outputs(1097));
    layer4_outputs(2467) <= (layer3_outputs(1490)) and (layer3_outputs(110));
    layer4_outputs(2468) <= (layer3_outputs(243)) xor (layer3_outputs(643));
    layer4_outputs(2469) <= (layer3_outputs(4041)) and (layer3_outputs(23));
    layer4_outputs(2470) <= not(layer3_outputs(940));
    layer4_outputs(2471) <= '0';
    layer4_outputs(2472) <= '0';
    layer4_outputs(2473) <= (layer3_outputs(2162)) and (layer3_outputs(2239));
    layer4_outputs(2474) <= not((layer3_outputs(3966)) and (layer3_outputs(985)));
    layer4_outputs(2475) <= (layer3_outputs(1062)) and not (layer3_outputs(3221));
    layer4_outputs(2476) <= (layer3_outputs(3317)) and not (layer3_outputs(3589));
    layer4_outputs(2477) <= (layer3_outputs(2349)) xor (layer3_outputs(3205));
    layer4_outputs(2478) <= (layer3_outputs(3210)) and not (layer3_outputs(4866));
    layer4_outputs(2479) <= not(layer3_outputs(4031)) or (layer3_outputs(3700));
    layer4_outputs(2480) <= (layer3_outputs(3892)) and not (layer3_outputs(1464));
    layer4_outputs(2481) <= '0';
    layer4_outputs(2482) <= layer3_outputs(138);
    layer4_outputs(2483) <= (layer3_outputs(1955)) and not (layer3_outputs(3189));
    layer4_outputs(2484) <= (layer3_outputs(4665)) and not (layer3_outputs(2230));
    layer4_outputs(2485) <= '1';
    layer4_outputs(2486) <= '0';
    layer4_outputs(2487) <= not(layer3_outputs(2632));
    layer4_outputs(2488) <= not(layer3_outputs(4615)) or (layer3_outputs(4541));
    layer4_outputs(2489) <= (layer3_outputs(2965)) and (layer3_outputs(2910));
    layer4_outputs(2490) <= not(layer3_outputs(3642));
    layer4_outputs(2491) <= (layer3_outputs(1835)) and not (layer3_outputs(3162));
    layer4_outputs(2492) <= (layer3_outputs(1922)) and not (layer3_outputs(1737));
    layer4_outputs(2493) <= '1';
    layer4_outputs(2494) <= (layer3_outputs(775)) and not (layer3_outputs(2163));
    layer4_outputs(2495) <= not((layer3_outputs(740)) and (layer3_outputs(674)));
    layer4_outputs(2496) <= not((layer3_outputs(4348)) and (layer3_outputs(1187)));
    layer4_outputs(2497) <= layer3_outputs(1847);
    layer4_outputs(2498) <= layer3_outputs(1084);
    layer4_outputs(2499) <= layer3_outputs(376);
    layer4_outputs(2500) <= (layer3_outputs(4639)) and not (layer3_outputs(2793));
    layer4_outputs(2501) <= not(layer3_outputs(4633));
    layer4_outputs(2502) <= not(layer3_outputs(2066));
    layer4_outputs(2503) <= layer3_outputs(732);
    layer4_outputs(2504) <= not((layer3_outputs(3278)) or (layer3_outputs(1660)));
    layer4_outputs(2505) <= not(layer3_outputs(5007));
    layer4_outputs(2506) <= (layer3_outputs(4582)) and not (layer3_outputs(4600));
    layer4_outputs(2507) <= not(layer3_outputs(1655)) or (layer3_outputs(172));
    layer4_outputs(2508) <= layer3_outputs(3808);
    layer4_outputs(2509) <= not((layer3_outputs(2711)) xor (layer3_outputs(1789)));
    layer4_outputs(2510) <= '1';
    layer4_outputs(2511) <= layer3_outputs(3965);
    layer4_outputs(2512) <= (layer3_outputs(48)) and not (layer3_outputs(3912));
    layer4_outputs(2513) <= not(layer3_outputs(3308)) or (layer3_outputs(1516));
    layer4_outputs(2514) <= '0';
    layer4_outputs(2515) <= not(layer3_outputs(2521));
    layer4_outputs(2516) <= not((layer3_outputs(1516)) and (layer3_outputs(1827)));
    layer4_outputs(2517) <= layer3_outputs(3644);
    layer4_outputs(2518) <= not(layer3_outputs(1928)) or (layer3_outputs(5068));
    layer4_outputs(2519) <= not(layer3_outputs(3042));
    layer4_outputs(2520) <= '1';
    layer4_outputs(2521) <= (layer3_outputs(3559)) or (layer3_outputs(4704));
    layer4_outputs(2522) <= (layer3_outputs(521)) and not (layer3_outputs(2320));
    layer4_outputs(2523) <= not(layer3_outputs(3285));
    layer4_outputs(2524) <= not(layer3_outputs(4761));
    layer4_outputs(2525) <= not(layer3_outputs(3825));
    layer4_outputs(2526) <= (layer3_outputs(1996)) or (layer3_outputs(2189));
    layer4_outputs(2527) <= '1';
    layer4_outputs(2528) <= not(layer3_outputs(2903));
    layer4_outputs(2529) <= layer3_outputs(887);
    layer4_outputs(2530) <= not(layer3_outputs(4668));
    layer4_outputs(2531) <= not((layer3_outputs(960)) and (layer3_outputs(3763)));
    layer4_outputs(2532) <= not((layer3_outputs(3137)) or (layer3_outputs(3957)));
    layer4_outputs(2533) <= '1';
    layer4_outputs(2534) <= not((layer3_outputs(999)) or (layer3_outputs(4966)));
    layer4_outputs(2535) <= not(layer3_outputs(1948));
    layer4_outputs(2536) <= not(layer3_outputs(2957));
    layer4_outputs(2537) <= '1';
    layer4_outputs(2538) <= (layer3_outputs(2357)) and not (layer3_outputs(893));
    layer4_outputs(2539) <= not(layer3_outputs(1662)) or (layer3_outputs(1128));
    layer4_outputs(2540) <= (layer3_outputs(1268)) or (layer3_outputs(1904));
    layer4_outputs(2541) <= not(layer3_outputs(2551)) or (layer3_outputs(2705));
    layer4_outputs(2542) <= not(layer3_outputs(3575));
    layer4_outputs(2543) <= layer3_outputs(2915);
    layer4_outputs(2544) <= layer3_outputs(2344);
    layer4_outputs(2545) <= not(layer3_outputs(4918));
    layer4_outputs(2546) <= '0';
    layer4_outputs(2547) <= (layer3_outputs(2301)) and (layer3_outputs(3094));
    layer4_outputs(2548) <= not((layer3_outputs(4473)) and (layer3_outputs(4552)));
    layer4_outputs(2549) <= not((layer3_outputs(1154)) xor (layer3_outputs(2517)));
    layer4_outputs(2550) <= not((layer3_outputs(588)) or (layer3_outputs(1886)));
    layer4_outputs(2551) <= (layer3_outputs(2450)) or (layer3_outputs(2354));
    layer4_outputs(2552) <= not(layer3_outputs(1372));
    layer4_outputs(2553) <= layer3_outputs(568);
    layer4_outputs(2554) <= not(layer3_outputs(2813));
    layer4_outputs(2555) <= '1';
    layer4_outputs(2556) <= not((layer3_outputs(1477)) and (layer3_outputs(917)));
    layer4_outputs(2557) <= '0';
    layer4_outputs(2558) <= not(layer3_outputs(3981)) or (layer3_outputs(2934));
    layer4_outputs(2559) <= layer3_outputs(1803);
    layer4_outputs(2560) <= not(layer3_outputs(4681));
    layer4_outputs(2561) <= not(layer3_outputs(898)) or (layer3_outputs(167));
    layer4_outputs(2562) <= not(layer3_outputs(2819));
    layer4_outputs(2563) <= not((layer3_outputs(3883)) and (layer3_outputs(4870)));
    layer4_outputs(2564) <= not(layer3_outputs(678));
    layer4_outputs(2565) <= not(layer3_outputs(3799)) or (layer3_outputs(43));
    layer4_outputs(2566) <= not(layer3_outputs(1620));
    layer4_outputs(2567) <= not((layer3_outputs(3108)) or (layer3_outputs(2186)));
    layer4_outputs(2568) <= (layer3_outputs(1202)) and not (layer3_outputs(4543));
    layer4_outputs(2569) <= layer3_outputs(148);
    layer4_outputs(2570) <= not(layer3_outputs(2913));
    layer4_outputs(2571) <= not(layer3_outputs(4648)) or (layer3_outputs(299));
    layer4_outputs(2572) <= '0';
    layer4_outputs(2573) <= '1';
    layer4_outputs(2574) <= (layer3_outputs(4599)) and (layer3_outputs(5031));
    layer4_outputs(2575) <= '1';
    layer4_outputs(2576) <= (layer3_outputs(1555)) and not (layer3_outputs(2190));
    layer4_outputs(2577) <= (layer3_outputs(1186)) or (layer3_outputs(3084));
    layer4_outputs(2578) <= not((layer3_outputs(5018)) and (layer3_outputs(3614)));
    layer4_outputs(2579) <= not((layer3_outputs(1116)) or (layer3_outputs(4762)));
    layer4_outputs(2580) <= not((layer3_outputs(4640)) and (layer3_outputs(4277)));
    layer4_outputs(2581) <= (layer3_outputs(3257)) and not (layer3_outputs(2154));
    layer4_outputs(2582) <= (layer3_outputs(2848)) and not (layer3_outputs(3586));
    layer4_outputs(2583) <= not(layer3_outputs(1909)) or (layer3_outputs(34));
    layer4_outputs(2584) <= not((layer3_outputs(2556)) and (layer3_outputs(1502)));
    layer4_outputs(2585) <= layer3_outputs(1775);
    layer4_outputs(2586) <= (layer3_outputs(3783)) and not (layer3_outputs(3419));
    layer4_outputs(2587) <= not(layer3_outputs(1307));
    layer4_outputs(2588) <= not((layer3_outputs(138)) and (layer3_outputs(3988)));
    layer4_outputs(2589) <= (layer3_outputs(1112)) and (layer3_outputs(1590));
    layer4_outputs(2590) <= not((layer3_outputs(1798)) or (layer3_outputs(2820)));
    layer4_outputs(2591) <= not((layer3_outputs(1983)) or (layer3_outputs(1053)));
    layer4_outputs(2592) <= not((layer3_outputs(4408)) or (layer3_outputs(2228)));
    layer4_outputs(2593) <= (layer3_outputs(3982)) and (layer3_outputs(136));
    layer4_outputs(2594) <= (layer3_outputs(936)) and not (layer3_outputs(1089));
    layer4_outputs(2595) <= not(layer3_outputs(1203));
    layer4_outputs(2596) <= (layer3_outputs(1347)) and not (layer3_outputs(4077));
    layer4_outputs(2597) <= (layer3_outputs(2533)) and not (layer3_outputs(1479));
    layer4_outputs(2598) <= (layer3_outputs(807)) and (layer3_outputs(1437));
    layer4_outputs(2599) <= (layer3_outputs(1840)) and not (layer3_outputs(2078));
    layer4_outputs(2600) <= not(layer3_outputs(2891)) or (layer3_outputs(448));
    layer4_outputs(2601) <= '0';
    layer4_outputs(2602) <= not((layer3_outputs(3946)) and (layer3_outputs(1415)));
    layer4_outputs(2603) <= (layer3_outputs(1980)) xor (layer3_outputs(2682));
    layer4_outputs(2604) <= '1';
    layer4_outputs(2605) <= '0';
    layer4_outputs(2606) <= not(layer3_outputs(4653));
    layer4_outputs(2607) <= not((layer3_outputs(1911)) or (layer3_outputs(1182)));
    layer4_outputs(2608) <= not(layer3_outputs(2952));
    layer4_outputs(2609) <= not(layer3_outputs(1172)) or (layer3_outputs(2231));
    layer4_outputs(2610) <= (layer3_outputs(4489)) and not (layer3_outputs(2061));
    layer4_outputs(2611) <= (layer3_outputs(3331)) xor (layer3_outputs(4225));
    layer4_outputs(2612) <= '0';
    layer4_outputs(2613) <= layer3_outputs(3759);
    layer4_outputs(2614) <= (layer3_outputs(152)) and not (layer3_outputs(3230));
    layer4_outputs(2615) <= (layer3_outputs(33)) or (layer3_outputs(1379));
    layer4_outputs(2616) <= layer3_outputs(678);
    layer4_outputs(2617) <= layer3_outputs(288);
    layer4_outputs(2618) <= (layer3_outputs(1105)) and not (layer3_outputs(510));
    layer4_outputs(2619) <= not(layer3_outputs(770));
    layer4_outputs(2620) <= layer3_outputs(1794);
    layer4_outputs(2621) <= (layer3_outputs(1693)) or (layer3_outputs(1658));
    layer4_outputs(2622) <= '1';
    layer4_outputs(2623) <= '1';
    layer4_outputs(2624) <= not((layer3_outputs(2793)) or (layer3_outputs(4267)));
    layer4_outputs(2625) <= (layer3_outputs(217)) and (layer3_outputs(1512));
    layer4_outputs(2626) <= not(layer3_outputs(1746));
    layer4_outputs(2627) <= (layer3_outputs(4977)) or (layer3_outputs(3927));
    layer4_outputs(2628) <= layer3_outputs(2941);
    layer4_outputs(2629) <= '1';
    layer4_outputs(2630) <= not(layer3_outputs(3033)) or (layer3_outputs(2715));
    layer4_outputs(2631) <= '1';
    layer4_outputs(2632) <= not((layer3_outputs(2731)) xor (layer3_outputs(1191)));
    layer4_outputs(2633) <= (layer3_outputs(3337)) and (layer3_outputs(1096));
    layer4_outputs(2634) <= not(layer3_outputs(2562)) or (layer3_outputs(2932));
    layer4_outputs(2635) <= not(layer3_outputs(1174)) or (layer3_outputs(1920));
    layer4_outputs(2636) <= not(layer3_outputs(4121)) or (layer3_outputs(5002));
    layer4_outputs(2637) <= '0';
    layer4_outputs(2638) <= layer3_outputs(1925);
    layer4_outputs(2639) <= (layer3_outputs(1228)) and not (layer3_outputs(3710));
    layer4_outputs(2640) <= '0';
    layer4_outputs(2641) <= (layer3_outputs(2210)) or (layer3_outputs(416));
    layer4_outputs(2642) <= (layer3_outputs(3787)) and (layer3_outputs(4392));
    layer4_outputs(2643) <= not(layer3_outputs(3139)) or (layer3_outputs(1977));
    layer4_outputs(2644) <= not(layer3_outputs(3761)) or (layer3_outputs(1060));
    layer4_outputs(2645) <= (layer3_outputs(3945)) and (layer3_outputs(5036));
    layer4_outputs(2646) <= (layer3_outputs(375)) and not (layer3_outputs(4683));
    layer4_outputs(2647) <= not((layer3_outputs(3046)) or (layer3_outputs(2502)));
    layer4_outputs(2648) <= (layer3_outputs(4188)) and not (layer3_outputs(4125));
    layer4_outputs(2649) <= layer3_outputs(1541);
    layer4_outputs(2650) <= '0';
    layer4_outputs(2651) <= layer3_outputs(3672);
    layer4_outputs(2652) <= (layer3_outputs(1424)) and not (layer3_outputs(1506));
    layer4_outputs(2653) <= '1';
    layer4_outputs(2654) <= not(layer3_outputs(480));
    layer4_outputs(2655) <= layer3_outputs(163);
    layer4_outputs(2656) <= layer3_outputs(4054);
    layer4_outputs(2657) <= not((layer3_outputs(2520)) and (layer3_outputs(572)));
    layer4_outputs(2658) <= layer3_outputs(646);
    layer4_outputs(2659) <= not(layer3_outputs(1398));
    layer4_outputs(2660) <= layer3_outputs(2875);
    layer4_outputs(2661) <= layer3_outputs(3483);
    layer4_outputs(2662) <= '0';
    layer4_outputs(2663) <= not(layer3_outputs(1180)) or (layer3_outputs(2471));
    layer4_outputs(2664) <= layer3_outputs(4809);
    layer4_outputs(2665) <= (layer3_outputs(856)) or (layer3_outputs(1292));
    layer4_outputs(2666) <= '0';
    layer4_outputs(2667) <= not((layer3_outputs(618)) and (layer3_outputs(889)));
    layer4_outputs(2668) <= not(layer3_outputs(625)) or (layer3_outputs(2431));
    layer4_outputs(2669) <= '0';
    layer4_outputs(2670) <= layer3_outputs(563);
    layer4_outputs(2671) <= not((layer3_outputs(1604)) or (layer3_outputs(69)));
    layer4_outputs(2672) <= (layer3_outputs(2034)) and not (layer3_outputs(4029));
    layer4_outputs(2673) <= not(layer3_outputs(453)) or (layer3_outputs(908));
    layer4_outputs(2674) <= layer3_outputs(3005);
    layer4_outputs(2675) <= layer3_outputs(4594);
    layer4_outputs(2676) <= not((layer3_outputs(836)) or (layer3_outputs(1018)));
    layer4_outputs(2677) <= '1';
    layer4_outputs(2678) <= (layer3_outputs(2897)) and not (layer3_outputs(4408));
    layer4_outputs(2679) <= not(layer3_outputs(3788)) or (layer3_outputs(4355));
    layer4_outputs(2680) <= layer3_outputs(3779);
    layer4_outputs(2681) <= not(layer3_outputs(4136));
    layer4_outputs(2682) <= not(layer3_outputs(420));
    layer4_outputs(2683) <= '1';
    layer4_outputs(2684) <= '0';
    layer4_outputs(2685) <= (layer3_outputs(978)) and not (layer3_outputs(1978));
    layer4_outputs(2686) <= not(layer3_outputs(4070));
    layer4_outputs(2687) <= '0';
    layer4_outputs(2688) <= not((layer3_outputs(1731)) or (layer3_outputs(4879)));
    layer4_outputs(2689) <= '0';
    layer4_outputs(2690) <= '0';
    layer4_outputs(2691) <= layer3_outputs(2186);
    layer4_outputs(2692) <= layer3_outputs(2570);
    layer4_outputs(2693) <= not(layer3_outputs(1048));
    layer4_outputs(2694) <= not(layer3_outputs(4046));
    layer4_outputs(2695) <= not(layer3_outputs(3392)) or (layer3_outputs(1110));
    layer4_outputs(2696) <= layer3_outputs(2803);
    layer4_outputs(2697) <= layer3_outputs(2626);
    layer4_outputs(2698) <= not(layer3_outputs(1343));
    layer4_outputs(2699) <= not(layer3_outputs(3214));
    layer4_outputs(2700) <= not(layer3_outputs(909)) or (layer3_outputs(1279));
    layer4_outputs(2701) <= layer3_outputs(1631);
    layer4_outputs(2702) <= '1';
    layer4_outputs(2703) <= not(layer3_outputs(4307));
    layer4_outputs(2704) <= not(layer3_outputs(1014)) or (layer3_outputs(4463));
    layer4_outputs(2705) <= not(layer3_outputs(1990));
    layer4_outputs(2706) <= '0';
    layer4_outputs(2707) <= not((layer3_outputs(4265)) or (layer3_outputs(4000)));
    layer4_outputs(2708) <= layer3_outputs(998);
    layer4_outputs(2709) <= not((layer3_outputs(2307)) and (layer3_outputs(3252)));
    layer4_outputs(2710) <= not(layer3_outputs(852)) or (layer3_outputs(1017));
    layer4_outputs(2711) <= not((layer3_outputs(4864)) and (layer3_outputs(1002)));
    layer4_outputs(2712) <= layer3_outputs(3527);
    layer4_outputs(2713) <= (layer3_outputs(2318)) and (layer3_outputs(586));
    layer4_outputs(2714) <= (layer3_outputs(2219)) and not (layer3_outputs(1313));
    layer4_outputs(2715) <= layer3_outputs(938);
    layer4_outputs(2716) <= layer3_outputs(1382);
    layer4_outputs(2717) <= not(layer3_outputs(501)) or (layer3_outputs(606));
    layer4_outputs(2718) <= layer3_outputs(28);
    layer4_outputs(2719) <= not(layer3_outputs(3822)) or (layer3_outputs(4191));
    layer4_outputs(2720) <= not(layer3_outputs(3425)) or (layer3_outputs(4836));
    layer4_outputs(2721) <= layer3_outputs(1397);
    layer4_outputs(2722) <= '1';
    layer4_outputs(2723) <= layer3_outputs(599);
    layer4_outputs(2724) <= (layer3_outputs(462)) and not (layer3_outputs(632));
    layer4_outputs(2725) <= layer3_outputs(4094);
    layer4_outputs(2726) <= (layer3_outputs(2868)) and not (layer3_outputs(778));
    layer4_outputs(2727) <= (layer3_outputs(4862)) and (layer3_outputs(1438));
    layer4_outputs(2728) <= '0';
    layer4_outputs(2729) <= (layer3_outputs(3911)) or (layer3_outputs(965));
    layer4_outputs(2730) <= '1';
    layer4_outputs(2731) <= (layer3_outputs(4567)) and (layer3_outputs(5119));
    layer4_outputs(2732) <= layer3_outputs(3503);
    layer4_outputs(2733) <= (layer3_outputs(4360)) and (layer3_outputs(4570));
    layer4_outputs(2734) <= (layer3_outputs(1446)) or (layer3_outputs(2240));
    layer4_outputs(2735) <= (layer3_outputs(1623)) and not (layer3_outputs(2890));
    layer4_outputs(2736) <= not((layer3_outputs(2536)) and (layer3_outputs(35)));
    layer4_outputs(2737) <= not((layer3_outputs(4862)) and (layer3_outputs(2707)));
    layer4_outputs(2738) <= (layer3_outputs(1404)) or (layer3_outputs(1217));
    layer4_outputs(2739) <= layer3_outputs(1128);
    layer4_outputs(2740) <= layer3_outputs(5024);
    layer4_outputs(2741) <= not(layer3_outputs(3129));
    layer4_outputs(2742) <= (layer3_outputs(709)) or (layer3_outputs(1776));
    layer4_outputs(2743) <= '0';
    layer4_outputs(2744) <= not((layer3_outputs(814)) and (layer3_outputs(75)));
    layer4_outputs(2745) <= not(layer3_outputs(3645));
    layer4_outputs(2746) <= '0';
    layer4_outputs(2747) <= not(layer3_outputs(2825));
    layer4_outputs(2748) <= (layer3_outputs(1172)) and (layer3_outputs(1335));
    layer4_outputs(2749) <= not(layer3_outputs(3354)) or (layer3_outputs(3112));
    layer4_outputs(2750) <= (layer3_outputs(3652)) or (layer3_outputs(2568));
    layer4_outputs(2751) <= (layer3_outputs(4863)) xor (layer3_outputs(2079));
    layer4_outputs(2752) <= layer3_outputs(3980);
    layer4_outputs(2753) <= not(layer3_outputs(4684));
    layer4_outputs(2754) <= not(layer3_outputs(1363)) or (layer3_outputs(1032));
    layer4_outputs(2755) <= not(layer3_outputs(5071));
    layer4_outputs(2756) <= not((layer3_outputs(2328)) and (layer3_outputs(3748)));
    layer4_outputs(2757) <= not(layer3_outputs(1218));
    layer4_outputs(2758) <= not(layer3_outputs(5082));
    layer4_outputs(2759) <= '1';
    layer4_outputs(2760) <= (layer3_outputs(1693)) and not (layer3_outputs(1959));
    layer4_outputs(2761) <= '0';
    layer4_outputs(2762) <= '1';
    layer4_outputs(2763) <= '1';
    layer4_outputs(2764) <= not(layer3_outputs(4284));
    layer4_outputs(2765) <= not(layer3_outputs(2481)) or (layer3_outputs(458));
    layer4_outputs(2766) <= not(layer3_outputs(3423));
    layer4_outputs(2767) <= '1';
    layer4_outputs(2768) <= (layer3_outputs(4251)) and not (layer3_outputs(271));
    layer4_outputs(2769) <= not((layer3_outputs(1385)) and (layer3_outputs(2914)));
    layer4_outputs(2770) <= layer3_outputs(3664);
    layer4_outputs(2771) <= layer3_outputs(2525);
    layer4_outputs(2772) <= (layer3_outputs(1408)) and not (layer3_outputs(3660));
    layer4_outputs(2773) <= (layer3_outputs(2680)) or (layer3_outputs(1048));
    layer4_outputs(2774) <= (layer3_outputs(4036)) and (layer3_outputs(991));
    layer4_outputs(2775) <= not((layer3_outputs(180)) and (layer3_outputs(4781)));
    layer4_outputs(2776) <= layer3_outputs(2212);
    layer4_outputs(2777) <= not(layer3_outputs(2269));
    layer4_outputs(2778) <= '0';
    layer4_outputs(2779) <= not(layer3_outputs(2665)) or (layer3_outputs(2597));
    layer4_outputs(2780) <= layer3_outputs(3332);
    layer4_outputs(2781) <= not((layer3_outputs(3817)) or (layer3_outputs(2019)));
    layer4_outputs(2782) <= '0';
    layer4_outputs(2783) <= (layer3_outputs(2337)) or (layer3_outputs(470));
    layer4_outputs(2784) <= (layer3_outputs(674)) and not (layer3_outputs(2121));
    layer4_outputs(2785) <= layer3_outputs(1714);
    layer4_outputs(2786) <= not((layer3_outputs(1657)) or (layer3_outputs(1283)));
    layer4_outputs(2787) <= (layer3_outputs(3584)) and not (layer3_outputs(3256));
    layer4_outputs(2788) <= layer3_outputs(3704);
    layer4_outputs(2789) <= layer3_outputs(2592);
    layer4_outputs(2790) <= (layer3_outputs(3806)) or (layer3_outputs(1384));
    layer4_outputs(2791) <= '0';
    layer4_outputs(2792) <= layer3_outputs(3142);
    layer4_outputs(2793) <= not(layer3_outputs(4713)) or (layer3_outputs(1506));
    layer4_outputs(2794) <= not(layer3_outputs(4712)) or (layer3_outputs(802));
    layer4_outputs(2795) <= layer3_outputs(3844);
    layer4_outputs(2796) <= not(layer3_outputs(98));
    layer4_outputs(2797) <= '1';
    layer4_outputs(2798) <= '1';
    layer4_outputs(2799) <= not((layer3_outputs(2725)) or (layer3_outputs(2277)));
    layer4_outputs(2800) <= (layer3_outputs(53)) and not (layer3_outputs(3480));
    layer4_outputs(2801) <= (layer3_outputs(1646)) and not (layer3_outputs(1862));
    layer4_outputs(2802) <= not(layer3_outputs(322));
    layer4_outputs(2803) <= not((layer3_outputs(3548)) xor (layer3_outputs(1393)));
    layer4_outputs(2804) <= (layer3_outputs(3062)) or (layer3_outputs(1096));
    layer4_outputs(2805) <= not(layer3_outputs(2476)) or (layer3_outputs(4049));
    layer4_outputs(2806) <= '0';
    layer4_outputs(2807) <= '1';
    layer4_outputs(2808) <= '1';
    layer4_outputs(2809) <= '1';
    layer4_outputs(2810) <= (layer3_outputs(3578)) and not (layer3_outputs(5063));
    layer4_outputs(2811) <= layer3_outputs(4896);
    layer4_outputs(2812) <= not((layer3_outputs(3527)) and (layer3_outputs(1292)));
    layer4_outputs(2813) <= not((layer3_outputs(2967)) or (layer3_outputs(918)));
    layer4_outputs(2814) <= (layer3_outputs(4494)) and not (layer3_outputs(1129));
    layer4_outputs(2815) <= not((layer3_outputs(845)) and (layer3_outputs(4737)));
    layer4_outputs(2816) <= not((layer3_outputs(4539)) or (layer3_outputs(3636)));
    layer4_outputs(2817) <= not((layer3_outputs(3605)) or (layer3_outputs(3438)));
    layer4_outputs(2818) <= not(layer3_outputs(2755));
    layer4_outputs(2819) <= (layer3_outputs(5006)) and (layer3_outputs(1264));
    layer4_outputs(2820) <= not(layer3_outputs(16)) or (layer3_outputs(636));
    layer4_outputs(2821) <= '0';
    layer4_outputs(2822) <= not((layer3_outputs(437)) or (layer3_outputs(1185)));
    layer4_outputs(2823) <= (layer3_outputs(3606)) and not (layer3_outputs(312));
    layer4_outputs(2824) <= layer3_outputs(4079);
    layer4_outputs(2825) <= layer3_outputs(4024);
    layer4_outputs(2826) <= not((layer3_outputs(3314)) and (layer3_outputs(1391)));
    layer4_outputs(2827) <= not(layer3_outputs(754));
    layer4_outputs(2828) <= (layer3_outputs(3879)) and (layer3_outputs(1600));
    layer4_outputs(2829) <= not(layer3_outputs(1378)) or (layer3_outputs(745));
    layer4_outputs(2830) <= (layer3_outputs(1589)) and not (layer3_outputs(2498));
    layer4_outputs(2831) <= (layer3_outputs(3556)) and not (layer3_outputs(5051));
    layer4_outputs(2832) <= (layer3_outputs(4290)) and not (layer3_outputs(126));
    layer4_outputs(2833) <= not(layer3_outputs(454));
    layer4_outputs(2834) <= not(layer3_outputs(3726)) or (layer3_outputs(3993));
    layer4_outputs(2835) <= '0';
    layer4_outputs(2836) <= not(layer3_outputs(4260));
    layer4_outputs(2837) <= layer3_outputs(4883);
    layer4_outputs(2838) <= not(layer3_outputs(3739));
    layer4_outputs(2839) <= (layer3_outputs(3495)) xor (layer3_outputs(591));
    layer4_outputs(2840) <= (layer3_outputs(2737)) and not (layer3_outputs(4646));
    layer4_outputs(2841) <= not(layer3_outputs(2980));
    layer4_outputs(2842) <= (layer3_outputs(736)) or (layer3_outputs(2093));
    layer4_outputs(2843) <= layer3_outputs(3109);
    layer4_outputs(2844) <= not((layer3_outputs(1227)) or (layer3_outputs(2748)));
    layer4_outputs(2845) <= layer3_outputs(1039);
    layer4_outputs(2846) <= (layer3_outputs(3536)) and not (layer3_outputs(782));
    layer4_outputs(2847) <= not(layer3_outputs(3067));
    layer4_outputs(2848) <= not(layer3_outputs(4574));
    layer4_outputs(2849) <= '0';
    layer4_outputs(2850) <= not((layer3_outputs(1793)) and (layer3_outputs(4418)));
    layer4_outputs(2851) <= '1';
    layer4_outputs(2852) <= '1';
    layer4_outputs(2853) <= not(layer3_outputs(932));
    layer4_outputs(2854) <= not(layer3_outputs(3747));
    layer4_outputs(2855) <= '1';
    layer4_outputs(2856) <= (layer3_outputs(2481)) xor (layer3_outputs(4114));
    layer4_outputs(2857) <= not(layer3_outputs(2187)) or (layer3_outputs(3235));
    layer4_outputs(2858) <= layer3_outputs(2988);
    layer4_outputs(2859) <= layer3_outputs(4852);
    layer4_outputs(2860) <= layer3_outputs(2577);
    layer4_outputs(2861) <= layer3_outputs(1049);
    layer4_outputs(2862) <= layer3_outputs(2000);
    layer4_outputs(2863) <= not((layer3_outputs(621)) and (layer3_outputs(912)));
    layer4_outputs(2864) <= not((layer3_outputs(826)) and (layer3_outputs(182)));
    layer4_outputs(2865) <= not((layer3_outputs(1595)) and (layer3_outputs(2516)));
    layer4_outputs(2866) <= layer3_outputs(385);
    layer4_outputs(2867) <= not(layer3_outputs(3973));
    layer4_outputs(2868) <= not(layer3_outputs(3820));
    layer4_outputs(2869) <= (layer3_outputs(4525)) or (layer3_outputs(4644));
    layer4_outputs(2870) <= layer3_outputs(2105);
    layer4_outputs(2871) <= not(layer3_outputs(2668)) or (layer3_outputs(2586));
    layer4_outputs(2872) <= not(layer3_outputs(4899));
    layer4_outputs(2873) <= not((layer3_outputs(5008)) or (layer3_outputs(1908)));
    layer4_outputs(2874) <= not(layer3_outputs(1736)) or (layer3_outputs(3563));
    layer4_outputs(2875) <= not((layer3_outputs(2576)) or (layer3_outputs(2938)));
    layer4_outputs(2876) <= (layer3_outputs(3171)) or (layer3_outputs(4235));
    layer4_outputs(2877) <= (layer3_outputs(4658)) or (layer3_outputs(4203));
    layer4_outputs(2878) <= not(layer3_outputs(1274)) or (layer3_outputs(2361));
    layer4_outputs(2879) <= (layer3_outputs(2103)) or (layer3_outputs(2476));
    layer4_outputs(2880) <= (layer3_outputs(3068)) or (layer3_outputs(2453));
    layer4_outputs(2881) <= (layer3_outputs(723)) or (layer3_outputs(2046));
    layer4_outputs(2882) <= (layer3_outputs(1175)) and not (layer3_outputs(5002));
    layer4_outputs(2883) <= (layer3_outputs(4816)) xor (layer3_outputs(3323));
    layer4_outputs(2884) <= (layer3_outputs(179)) and not (layer3_outputs(2392));
    layer4_outputs(2885) <= '1';
    layer4_outputs(2886) <= not(layer3_outputs(4690));
    layer4_outputs(2887) <= not(layer3_outputs(2692));
    layer4_outputs(2888) <= (layer3_outputs(4405)) and (layer3_outputs(2209));
    layer4_outputs(2889) <= (layer3_outputs(3659)) and not (layer3_outputs(1210));
    layer4_outputs(2890) <= not(layer3_outputs(2217)) or (layer3_outputs(2068));
    layer4_outputs(2891) <= not(layer3_outputs(4347));
    layer4_outputs(2892) <= not(layer3_outputs(4454));
    layer4_outputs(2893) <= layer3_outputs(2202);
    layer4_outputs(2894) <= not(layer3_outputs(1453));
    layer4_outputs(2895) <= layer3_outputs(1636);
    layer4_outputs(2896) <= not((layer3_outputs(388)) xor (layer3_outputs(2513)));
    layer4_outputs(2897) <= not(layer3_outputs(3690));
    layer4_outputs(2898) <= layer3_outputs(3247);
    layer4_outputs(2899) <= not((layer3_outputs(2895)) or (layer3_outputs(1557)));
    layer4_outputs(2900) <= '0';
    layer4_outputs(2901) <= (layer3_outputs(1874)) and (layer3_outputs(1520));
    layer4_outputs(2902) <= '0';
    layer4_outputs(2903) <= (layer3_outputs(2383)) and not (layer3_outputs(4397));
    layer4_outputs(2904) <= not((layer3_outputs(3352)) or (layer3_outputs(5009)));
    layer4_outputs(2905) <= not(layer3_outputs(5014));
    layer4_outputs(2906) <= (layer3_outputs(690)) and not (layer3_outputs(2160));
    layer4_outputs(2907) <= not(layer3_outputs(1680));
    layer4_outputs(2908) <= layer3_outputs(765);
    layer4_outputs(2909) <= not(layer3_outputs(990));
    layer4_outputs(2910) <= '1';
    layer4_outputs(2911) <= layer3_outputs(3852);
    layer4_outputs(2912) <= not((layer3_outputs(2349)) or (layer3_outputs(3818)));
    layer4_outputs(2913) <= (layer3_outputs(1685)) and not (layer3_outputs(37));
    layer4_outputs(2914) <= (layer3_outputs(481)) and not (layer3_outputs(4672));
    layer4_outputs(2915) <= not((layer3_outputs(1173)) and (layer3_outputs(4337)));
    layer4_outputs(2916) <= not((layer3_outputs(2157)) and (layer3_outputs(4433)));
    layer4_outputs(2917) <= not(layer3_outputs(2041)) or (layer3_outputs(3522));
    layer4_outputs(2918) <= not(layer3_outputs(1792)) or (layer3_outputs(2962));
    layer4_outputs(2919) <= (layer3_outputs(265)) and not (layer3_outputs(2693));
    layer4_outputs(2920) <= layer3_outputs(4814);
    layer4_outputs(2921) <= not(layer3_outputs(4195));
    layer4_outputs(2922) <= layer3_outputs(4642);
    layer4_outputs(2923) <= not((layer3_outputs(3387)) or (layer3_outputs(80)));
    layer4_outputs(2924) <= layer3_outputs(1800);
    layer4_outputs(2925) <= layer3_outputs(2463);
    layer4_outputs(2926) <= '1';
    layer4_outputs(2927) <= not(layer3_outputs(519)) or (layer3_outputs(349));
    layer4_outputs(2928) <= layer3_outputs(3867);
    layer4_outputs(2929) <= layer3_outputs(4212);
    layer4_outputs(2930) <= (layer3_outputs(366)) and not (layer3_outputs(4725));
    layer4_outputs(2931) <= not((layer3_outputs(1228)) or (layer3_outputs(2661)));
    layer4_outputs(2932) <= (layer3_outputs(1779)) and not (layer3_outputs(323));
    layer4_outputs(2933) <= layer3_outputs(4897);
    layer4_outputs(2934) <= not(layer3_outputs(3516)) or (layer3_outputs(828));
    layer4_outputs(2935) <= not(layer3_outputs(2508)) or (layer3_outputs(4387));
    layer4_outputs(2936) <= not(layer3_outputs(4986));
    layer4_outputs(2937) <= not((layer3_outputs(3962)) and (layer3_outputs(2335)));
    layer4_outputs(2938) <= '1';
    layer4_outputs(2939) <= not(layer3_outputs(4117)) or (layer3_outputs(6));
    layer4_outputs(2940) <= (layer3_outputs(3133)) and not (layer3_outputs(2273));
    layer4_outputs(2941) <= (layer3_outputs(4361)) and (layer3_outputs(1766));
    layer4_outputs(2942) <= not(layer3_outputs(2723));
    layer4_outputs(2943) <= '0';
    layer4_outputs(2944) <= (layer3_outputs(4684)) and not (layer3_outputs(116));
    layer4_outputs(2945) <= (layer3_outputs(2065)) and not (layer3_outputs(4740));
    layer4_outputs(2946) <= not(layer3_outputs(4528));
    layer4_outputs(2947) <= not(layer3_outputs(4299));
    layer4_outputs(2948) <= not(layer3_outputs(472));
    layer4_outputs(2949) <= (layer3_outputs(4109)) or (layer3_outputs(4060));
    layer4_outputs(2950) <= '1';
    layer4_outputs(2951) <= not(layer3_outputs(4196)) or (layer3_outputs(311));
    layer4_outputs(2952) <= not(layer3_outputs(908));
    layer4_outputs(2953) <= (layer3_outputs(3479)) and not (layer3_outputs(720));
    layer4_outputs(2954) <= (layer3_outputs(5065)) and (layer3_outputs(1324));
    layer4_outputs(2955) <= not((layer3_outputs(1075)) and (layer3_outputs(1926)));
    layer4_outputs(2956) <= not(layer3_outputs(3996)) or (layer3_outputs(4411));
    layer4_outputs(2957) <= (layer3_outputs(1156)) and not (layer3_outputs(1852));
    layer4_outputs(2958) <= (layer3_outputs(1092)) xor (layer3_outputs(409));
    layer4_outputs(2959) <= not(layer3_outputs(2241));
    layer4_outputs(2960) <= not(layer3_outputs(2279)) or (layer3_outputs(4733));
    layer4_outputs(2961) <= '0';
    layer4_outputs(2962) <= (layer3_outputs(4442)) or (layer3_outputs(4504));
    layer4_outputs(2963) <= (layer3_outputs(2833)) or (layer3_outputs(337));
    layer4_outputs(2964) <= (layer3_outputs(2774)) and not (layer3_outputs(2828));
    layer4_outputs(2965) <= not(layer3_outputs(2968)) or (layer3_outputs(4418));
    layer4_outputs(2966) <= not(layer3_outputs(4514));
    layer4_outputs(2967) <= not(layer3_outputs(1872));
    layer4_outputs(2968) <= not((layer3_outputs(1787)) or (layer3_outputs(4133)));
    layer4_outputs(2969) <= not((layer3_outputs(1230)) or (layer3_outputs(3135)));
    layer4_outputs(2970) <= not(layer3_outputs(4356)) or (layer3_outputs(1608));
    layer4_outputs(2971) <= (layer3_outputs(4758)) xor (layer3_outputs(394));
    layer4_outputs(2972) <= not(layer3_outputs(1547));
    layer4_outputs(2973) <= '1';
    layer4_outputs(2974) <= layer3_outputs(1794);
    layer4_outputs(2975) <= not((layer3_outputs(1519)) or (layer3_outputs(1688)));
    layer4_outputs(2976) <= (layer3_outputs(4435)) and (layer3_outputs(897));
    layer4_outputs(2977) <= not(layer3_outputs(360));
    layer4_outputs(2978) <= layer3_outputs(2867);
    layer4_outputs(2979) <= (layer3_outputs(4911)) and not (layer3_outputs(3202));
    layer4_outputs(2980) <= '0';
    layer4_outputs(2981) <= layer3_outputs(1861);
    layer4_outputs(2982) <= not((layer3_outputs(442)) or (layer3_outputs(4430)));
    layer4_outputs(2983) <= not((layer3_outputs(100)) and (layer3_outputs(1674)));
    layer4_outputs(2984) <= layer3_outputs(473);
    layer4_outputs(2985) <= layer3_outputs(1884);
    layer4_outputs(2986) <= (layer3_outputs(1941)) and not (layer3_outputs(250));
    layer4_outputs(2987) <= '0';
    layer4_outputs(2988) <= not(layer3_outputs(1621));
    layer4_outputs(2989) <= (layer3_outputs(4333)) or (layer3_outputs(1262));
    layer4_outputs(2990) <= layer3_outputs(4362);
    layer4_outputs(2991) <= (layer3_outputs(5093)) and not (layer3_outputs(4698));
    layer4_outputs(2992) <= layer3_outputs(3322);
    layer4_outputs(2993) <= (layer3_outputs(3074)) and not (layer3_outputs(2409));
    layer4_outputs(2994) <= (layer3_outputs(1763)) xor (layer3_outputs(3979));
    layer4_outputs(2995) <= layer3_outputs(4116);
    layer4_outputs(2996) <= not(layer3_outputs(5103));
    layer4_outputs(2997) <= not(layer3_outputs(4974)) or (layer3_outputs(3037));
    layer4_outputs(2998) <= '0';
    layer4_outputs(2999) <= layer3_outputs(1131);
    layer4_outputs(3000) <= (layer3_outputs(3532)) and not (layer3_outputs(1931));
    layer4_outputs(3001) <= (layer3_outputs(2532)) or (layer3_outputs(2854));
    layer4_outputs(3002) <= not(layer3_outputs(2689));
    layer4_outputs(3003) <= '0';
    layer4_outputs(3004) <= (layer3_outputs(760)) and (layer3_outputs(3918));
    layer4_outputs(3005) <= not(layer3_outputs(3944));
    layer4_outputs(3006) <= (layer3_outputs(1176)) and (layer3_outputs(439));
    layer4_outputs(3007) <= not(layer3_outputs(2005));
    layer4_outputs(3008) <= '1';
    layer4_outputs(3009) <= not(layer3_outputs(743)) or (layer3_outputs(2453));
    layer4_outputs(3010) <= (layer3_outputs(1134)) and not (layer3_outputs(2415));
    layer4_outputs(3011) <= '1';
    layer4_outputs(3012) <= (layer3_outputs(2044)) or (layer3_outputs(4570));
    layer4_outputs(3013) <= (layer3_outputs(4549)) and not (layer3_outputs(4629));
    layer4_outputs(3014) <= '0';
    layer4_outputs(3015) <= '0';
    layer4_outputs(3016) <= not(layer3_outputs(193));
    layer4_outputs(3017) <= layer3_outputs(92);
    layer4_outputs(3018) <= not(layer3_outputs(2857));
    layer4_outputs(3019) <= not((layer3_outputs(2657)) and (layer3_outputs(3668)));
    layer4_outputs(3020) <= (layer3_outputs(3010)) and not (layer3_outputs(4051));
    layer4_outputs(3021) <= layer3_outputs(3741);
    layer4_outputs(3022) <= not((layer3_outputs(3083)) or (layer3_outputs(185)));
    layer4_outputs(3023) <= (layer3_outputs(2384)) and not (layer3_outputs(1235));
    layer4_outputs(3024) <= not(layer3_outputs(3050));
    layer4_outputs(3025) <= not(layer3_outputs(907));
    layer4_outputs(3026) <= layer3_outputs(2933);
    layer4_outputs(3027) <= not((layer3_outputs(455)) and (layer3_outputs(3543)));
    layer4_outputs(3028) <= (layer3_outputs(552)) and not (layer3_outputs(727));
    layer4_outputs(3029) <= '1';
    layer4_outputs(3030) <= (layer3_outputs(4212)) or (layer3_outputs(1694));
    layer4_outputs(3031) <= (layer3_outputs(2500)) or (layer3_outputs(2111));
    layer4_outputs(3032) <= (layer3_outputs(3627)) and not (layer3_outputs(3947));
    layer4_outputs(3033) <= (layer3_outputs(3829)) or (layer3_outputs(1150));
    layer4_outputs(3034) <= (layer3_outputs(2449)) and (layer3_outputs(4065));
    layer4_outputs(3035) <= not(layer3_outputs(3414));
    layer4_outputs(3036) <= '1';
    layer4_outputs(3037) <= not(layer3_outputs(3079));
    layer4_outputs(3038) <= not(layer3_outputs(2756)) or (layer3_outputs(4651));
    layer4_outputs(3039) <= not(layer3_outputs(3736));
    layer4_outputs(3040) <= layer3_outputs(2747);
    layer4_outputs(3041) <= not(layer3_outputs(1376)) or (layer3_outputs(1091));
    layer4_outputs(3042) <= (layer3_outputs(1214)) xor (layer3_outputs(957));
    layer4_outputs(3043) <= not(layer3_outputs(148));
    layer4_outputs(3044) <= '1';
    layer4_outputs(3045) <= not(layer3_outputs(4136));
    layer4_outputs(3046) <= not(layer3_outputs(4176));
    layer4_outputs(3047) <= (layer3_outputs(4363)) and not (layer3_outputs(3092));
    layer4_outputs(3048) <= not(layer3_outputs(1581)) or (layer3_outputs(178));
    layer4_outputs(3049) <= not(layer3_outputs(4611)) or (layer3_outputs(3950));
    layer4_outputs(3050) <= not(layer3_outputs(1555));
    layer4_outputs(3051) <= '0';
    layer4_outputs(3052) <= not((layer3_outputs(4983)) and (layer3_outputs(2555)));
    layer4_outputs(3053) <= not((layer3_outputs(3273)) xor (layer3_outputs(2831)));
    layer4_outputs(3054) <= not(layer3_outputs(263));
    layer4_outputs(3055) <= '0';
    layer4_outputs(3056) <= not(layer3_outputs(3356));
    layer4_outputs(3057) <= not(layer3_outputs(2050)) or (layer3_outputs(1280));
    layer4_outputs(3058) <= not((layer3_outputs(3544)) and (layer3_outputs(3305)));
    layer4_outputs(3059) <= (layer3_outputs(592)) xor (layer3_outputs(467));
    layer4_outputs(3060) <= not((layer3_outputs(2746)) and (layer3_outputs(2375)));
    layer4_outputs(3061) <= not(layer3_outputs(1326));
    layer4_outputs(3062) <= not((layer3_outputs(1432)) or (layer3_outputs(3241)));
    layer4_outputs(3063) <= (layer3_outputs(5096)) and not (layer3_outputs(4617));
    layer4_outputs(3064) <= '0';
    layer4_outputs(3065) <= layer3_outputs(5027);
    layer4_outputs(3066) <= (layer3_outputs(2911)) and (layer3_outputs(4093));
    layer4_outputs(3067) <= not(layer3_outputs(4113));
    layer4_outputs(3068) <= not(layer3_outputs(2030)) or (layer3_outputs(2055));
    layer4_outputs(3069) <= '1';
    layer4_outputs(3070) <= layer3_outputs(1186);
    layer4_outputs(3071) <= not(layer3_outputs(536));
    layer4_outputs(3072) <= layer3_outputs(1363);
    layer4_outputs(3073) <= not(layer3_outputs(1522));
    layer4_outputs(3074) <= not(layer3_outputs(4224)) or (layer3_outputs(1482));
    layer4_outputs(3075) <= layer3_outputs(1187);
    layer4_outputs(3076) <= not((layer3_outputs(1982)) and (layer3_outputs(1714)));
    layer4_outputs(3077) <= '1';
    layer4_outputs(3078) <= not(layer3_outputs(1603)) or (layer3_outputs(5059));
    layer4_outputs(3079) <= not((layer3_outputs(3599)) or (layer3_outputs(543)));
    layer4_outputs(3080) <= layer3_outputs(2873);
    layer4_outputs(3081) <= (layer3_outputs(251)) and not (layer3_outputs(549));
    layer4_outputs(3082) <= (layer3_outputs(2819)) and (layer3_outputs(2907));
    layer4_outputs(3083) <= '0';
    layer4_outputs(3084) <= (layer3_outputs(1249)) and (layer3_outputs(3350));
    layer4_outputs(3085) <= '1';
    layer4_outputs(3086) <= not(layer3_outputs(4438)) or (layer3_outputs(2675));
    layer4_outputs(3087) <= not((layer3_outputs(2494)) or (layer3_outputs(1888)));
    layer4_outputs(3088) <= not(layer3_outputs(4060));
    layer4_outputs(3089) <= not(layer3_outputs(4533));
    layer4_outputs(3090) <= '1';
    layer4_outputs(3091) <= not((layer3_outputs(4334)) and (layer3_outputs(2607)));
    layer4_outputs(3092) <= not((layer3_outputs(3187)) and (layer3_outputs(4824)));
    layer4_outputs(3093) <= not((layer3_outputs(637)) and (layer3_outputs(859)));
    layer4_outputs(3094) <= not(layer3_outputs(2679)) or (layer3_outputs(1143));
    layer4_outputs(3095) <= (layer3_outputs(3767)) and (layer3_outputs(1005));
    layer4_outputs(3096) <= not(layer3_outputs(1481)) or (layer3_outputs(3866));
    layer4_outputs(3097) <= layer3_outputs(477);
    layer4_outputs(3098) <= not(layer3_outputs(4456));
    layer4_outputs(3099) <= not(layer3_outputs(3073)) or (layer3_outputs(3500));
    layer4_outputs(3100) <= (layer3_outputs(289)) and not (layer3_outputs(4507));
    layer4_outputs(3101) <= (layer3_outputs(2537)) and not (layer3_outputs(2897));
    layer4_outputs(3102) <= not(layer3_outputs(1973));
    layer4_outputs(3103) <= not((layer3_outputs(4557)) and (layer3_outputs(1768)));
    layer4_outputs(3104) <= not((layer3_outputs(3073)) and (layer3_outputs(1823)));
    layer4_outputs(3105) <= not((layer3_outputs(3265)) or (layer3_outputs(4664)));
    layer4_outputs(3106) <= (layer3_outputs(2115)) or (layer3_outputs(4815));
    layer4_outputs(3107) <= '0';
    layer4_outputs(3108) <= not(layer3_outputs(1200));
    layer4_outputs(3109) <= not((layer3_outputs(4333)) or (layer3_outputs(2855)));
    layer4_outputs(3110) <= (layer3_outputs(1232)) and (layer3_outputs(4300));
    layer4_outputs(3111) <= not(layer3_outputs(270));
    layer4_outputs(3112) <= (layer3_outputs(3339)) or (layer3_outputs(3795));
    layer4_outputs(3113) <= not(layer3_outputs(78));
    layer4_outputs(3114) <= (layer3_outputs(2214)) xor (layer3_outputs(4340));
    layer4_outputs(3115) <= layer3_outputs(750);
    layer4_outputs(3116) <= (layer3_outputs(4400)) or (layer3_outputs(1029));
    layer4_outputs(3117) <= not(layer3_outputs(1733));
    layer4_outputs(3118) <= not((layer3_outputs(2944)) or (layer3_outputs(4431)));
    layer4_outputs(3119) <= not(layer3_outputs(589)) or (layer3_outputs(1749));
    layer4_outputs(3120) <= (layer3_outputs(2042)) or (layer3_outputs(1583));
    layer4_outputs(3121) <= not(layer3_outputs(4486)) or (layer3_outputs(969));
    layer4_outputs(3122) <= layer3_outputs(1056);
    layer4_outputs(3123) <= (layer3_outputs(3885)) or (layer3_outputs(1161));
    layer4_outputs(3124) <= '1';
    layer4_outputs(3125) <= not(layer3_outputs(1364)) or (layer3_outputs(3351));
    layer4_outputs(3126) <= not(layer3_outputs(2635)) or (layer3_outputs(239));
    layer4_outputs(3127) <= layer3_outputs(2445);
    layer4_outputs(3128) <= '0';
    layer4_outputs(3129) <= not((layer3_outputs(97)) and (layer3_outputs(3046)));
    layer4_outputs(3130) <= not((layer3_outputs(3134)) and (layer3_outputs(3132)));
    layer4_outputs(3131) <= not((layer3_outputs(4109)) or (layer3_outputs(951)));
    layer4_outputs(3132) <= not((layer3_outputs(1214)) or (layer3_outputs(3117)));
    layer4_outputs(3133) <= not(layer3_outputs(2684)) or (layer3_outputs(4122));
    layer4_outputs(3134) <= not(layer3_outputs(1954)) or (layer3_outputs(3726));
    layer4_outputs(3135) <= (layer3_outputs(917)) and not (layer3_outputs(3443));
    layer4_outputs(3136) <= not(layer3_outputs(415));
    layer4_outputs(3137) <= '1';
    layer4_outputs(3138) <= layer3_outputs(4922);
    layer4_outputs(3139) <= '0';
    layer4_outputs(3140) <= not(layer3_outputs(1979)) or (layer3_outputs(4236));
    layer4_outputs(3141) <= not(layer3_outputs(644)) or (layer3_outputs(892));
    layer4_outputs(3142) <= (layer3_outputs(3687)) xor (layer3_outputs(4882));
    layer4_outputs(3143) <= (layer3_outputs(4783)) and not (layer3_outputs(2764));
    layer4_outputs(3144) <= not(layer3_outputs(2887)) or (layer3_outputs(2972));
    layer4_outputs(3145) <= not(layer3_outputs(1358)) or (layer3_outputs(1880));
    layer4_outputs(3146) <= not((layer3_outputs(1902)) and (layer3_outputs(2563)));
    layer4_outputs(3147) <= not((layer3_outputs(4220)) or (layer3_outputs(2886)));
    layer4_outputs(3148) <= not(layer3_outputs(4111)) or (layer3_outputs(4524));
    layer4_outputs(3149) <= not((layer3_outputs(1011)) or (layer3_outputs(2367)));
    layer4_outputs(3150) <= '1';
    layer4_outputs(3151) <= '1';
    layer4_outputs(3152) <= not(layer3_outputs(399));
    layer4_outputs(3153) <= layer3_outputs(4758);
    layer4_outputs(3154) <= not((layer3_outputs(3836)) and (layer3_outputs(3292)));
    layer4_outputs(3155) <= layer3_outputs(4015);
    layer4_outputs(3156) <= (layer3_outputs(4818)) and not (layer3_outputs(2396));
    layer4_outputs(3157) <= layer3_outputs(1995);
    layer4_outputs(3158) <= (layer3_outputs(434)) or (layer3_outputs(3));
    layer4_outputs(3159) <= not(layer3_outputs(1848));
    layer4_outputs(3160) <= (layer3_outputs(1323)) xor (layer3_outputs(4623));
    layer4_outputs(3161) <= not((layer3_outputs(700)) and (layer3_outputs(3112)));
    layer4_outputs(3162) <= '1';
    layer4_outputs(3163) <= (layer3_outputs(4606)) and not (layer3_outputs(177));
    layer4_outputs(3164) <= layer3_outputs(3390);
    layer4_outputs(3165) <= (layer3_outputs(3624)) and not (layer3_outputs(2821));
    layer4_outputs(3166) <= layer3_outputs(1190);
    layer4_outputs(3167) <= (layer3_outputs(3051)) or (layer3_outputs(1120));
    layer4_outputs(3168) <= layer3_outputs(931);
    layer4_outputs(3169) <= not((layer3_outputs(4985)) or (layer3_outputs(2595)));
    layer4_outputs(3170) <= '0';
    layer4_outputs(3171) <= (layer3_outputs(4009)) or (layer3_outputs(4840));
    layer4_outputs(3172) <= not((layer3_outputs(3837)) or (layer3_outputs(676)));
    layer4_outputs(3173) <= (layer3_outputs(1960)) xor (layer3_outputs(728));
    layer4_outputs(3174) <= '1';
    layer4_outputs(3175) <= layer3_outputs(4760);
    layer4_outputs(3176) <= not(layer3_outputs(3347));
    layer4_outputs(3177) <= '1';
    layer4_outputs(3178) <= (layer3_outputs(1613)) or (layer3_outputs(2325));
    layer4_outputs(3179) <= (layer3_outputs(1646)) and not (layer3_outputs(4909));
    layer4_outputs(3180) <= not(layer3_outputs(2317));
    layer4_outputs(3181) <= not((layer3_outputs(4413)) or (layer3_outputs(1946)));
    layer4_outputs(3182) <= '0';
    layer4_outputs(3183) <= not(layer3_outputs(3568)) or (layer3_outputs(246));
    layer4_outputs(3184) <= (layer3_outputs(3985)) or (layer3_outputs(2412));
    layer4_outputs(3185) <= (layer3_outputs(4182)) and not (layer3_outputs(2578));
    layer4_outputs(3186) <= not(layer3_outputs(795)) or (layer3_outputs(2357));
    layer4_outputs(3187) <= '1';
    layer4_outputs(3188) <= not(layer3_outputs(64)) or (layer3_outputs(2606));
    layer4_outputs(3189) <= (layer3_outputs(3176)) and not (layer3_outputs(4446));
    layer4_outputs(3190) <= not((layer3_outputs(1224)) or (layer3_outputs(2241)));
    layer4_outputs(3191) <= (layer3_outputs(4953)) and (layer3_outputs(4965));
    layer4_outputs(3192) <= (layer3_outputs(4742)) xor (layer3_outputs(2045));
    layer4_outputs(3193) <= not(layer3_outputs(3061)) or (layer3_outputs(3076));
    layer4_outputs(3194) <= '0';
    layer4_outputs(3195) <= not(layer3_outputs(4249)) or (layer3_outputs(4280));
    layer4_outputs(3196) <= '1';
    layer4_outputs(3197) <= layer3_outputs(2280);
    layer4_outputs(3198) <= not((layer3_outputs(301)) or (layer3_outputs(2973)));
    layer4_outputs(3199) <= (layer3_outputs(70)) and not (layer3_outputs(4297));
    layer4_outputs(3200) <= layer3_outputs(2148);
    layer4_outputs(3201) <= (layer3_outputs(794)) or (layer3_outputs(4678));
    layer4_outputs(3202) <= not(layer3_outputs(4839));
    layer4_outputs(3203) <= '0';
    layer4_outputs(3204) <= (layer3_outputs(3493)) and (layer3_outputs(3948));
    layer4_outputs(3205) <= layer3_outputs(1993);
    layer4_outputs(3206) <= not(layer3_outputs(355));
    layer4_outputs(3207) <= not((layer3_outputs(635)) and (layer3_outputs(1679)));
    layer4_outputs(3208) <= not(layer3_outputs(1245));
    layer4_outputs(3209) <= '1';
    layer4_outputs(3210) <= (layer3_outputs(4296)) and not (layer3_outputs(5053));
    layer4_outputs(3211) <= not(layer3_outputs(2710));
    layer4_outputs(3212) <= not((layer3_outputs(680)) or (layer3_outputs(861)));
    layer4_outputs(3213) <= not(layer3_outputs(936));
    layer4_outputs(3214) <= '1';
    layer4_outputs(3215) <= (layer3_outputs(317)) xor (layer3_outputs(4750));
    layer4_outputs(3216) <= (layer3_outputs(5041)) xor (layer3_outputs(2138));
    layer4_outputs(3217) <= layer3_outputs(1424);
    layer4_outputs(3218) <= not(layer3_outputs(1468)) or (layer3_outputs(4763));
    layer4_outputs(3219) <= not((layer3_outputs(3966)) or (layer3_outputs(4380)));
    layer4_outputs(3220) <= '0';
    layer4_outputs(3221) <= not(layer3_outputs(2685));
    layer4_outputs(3222) <= not((layer3_outputs(986)) or (layer3_outputs(4493)));
    layer4_outputs(3223) <= not((layer3_outputs(2984)) and (layer3_outputs(2181)));
    layer4_outputs(3224) <= not((layer3_outputs(3345)) and (layer3_outputs(1182)));
    layer4_outputs(3225) <= not((layer3_outputs(4066)) xor (layer3_outputs(2126)));
    layer4_outputs(3226) <= (layer3_outputs(1670)) and (layer3_outputs(2899));
    layer4_outputs(3227) <= '1';
    layer4_outputs(3228) <= (layer3_outputs(593)) and (layer3_outputs(2572));
    layer4_outputs(3229) <= not((layer3_outputs(1884)) and (layer3_outputs(803)));
    layer4_outputs(3230) <= '0';
    layer4_outputs(3231) <= (layer3_outputs(881)) xor (layer3_outputs(255));
    layer4_outputs(3232) <= (layer3_outputs(601)) and (layer3_outputs(4247));
    layer4_outputs(3233) <= layer3_outputs(3175);
    layer4_outputs(3234) <= (layer3_outputs(776)) and not (layer3_outputs(2445));
    layer4_outputs(3235) <= (layer3_outputs(342)) and (layer3_outputs(840));
    layer4_outputs(3236) <= layer3_outputs(4716);
    layer4_outputs(3237) <= not(layer3_outputs(1202));
    layer4_outputs(3238) <= (layer3_outputs(963)) and (layer3_outputs(3353));
    layer4_outputs(3239) <= not(layer3_outputs(5012));
    layer4_outputs(3240) <= not((layer3_outputs(3001)) and (layer3_outputs(2396)));
    layer4_outputs(3241) <= (layer3_outputs(2060)) and not (layer3_outputs(83));
    layer4_outputs(3242) <= layer3_outputs(1707);
    layer4_outputs(3243) <= (layer3_outputs(1566)) and (layer3_outputs(4038));
    layer4_outputs(3244) <= (layer3_outputs(3003)) xor (layer3_outputs(1830));
    layer4_outputs(3245) <= not(layer3_outputs(1342)) or (layer3_outputs(1104));
    layer4_outputs(3246) <= (layer3_outputs(668)) and not (layer3_outputs(2226));
    layer4_outputs(3247) <= not(layer3_outputs(3570)) or (layer3_outputs(1265));
    layer4_outputs(3248) <= (layer3_outputs(2405)) and not (layer3_outputs(4132));
    layer4_outputs(3249) <= layer3_outputs(4784);
    layer4_outputs(3250) <= (layer3_outputs(604)) and not (layer3_outputs(307));
    layer4_outputs(3251) <= (layer3_outputs(4337)) and not (layer3_outputs(3704));
    layer4_outputs(3252) <= not(layer3_outputs(1034)) or (layer3_outputs(3600));
    layer4_outputs(3253) <= (layer3_outputs(2683)) or (layer3_outputs(1431));
    layer4_outputs(3254) <= not((layer3_outputs(1399)) and (layer3_outputs(3346)));
    layer4_outputs(3255) <= not(layer3_outputs(3776));
    layer4_outputs(3256) <= not((layer3_outputs(824)) or (layer3_outputs(52)));
    layer4_outputs(3257) <= not(layer3_outputs(4578)) or (layer3_outputs(2271));
    layer4_outputs(3258) <= not((layer3_outputs(179)) or (layer3_outputs(3222)));
    layer4_outputs(3259) <= layer3_outputs(256);
    layer4_outputs(3260) <= layer3_outputs(701);
    layer4_outputs(3261) <= layer3_outputs(3706);
    layer4_outputs(3262) <= not((layer3_outputs(1039)) and (layer3_outputs(3002)));
    layer4_outputs(3263) <= not(layer3_outputs(1819)) or (layer3_outputs(1626));
    layer4_outputs(3264) <= layer3_outputs(3404);
    layer4_outputs(3265) <= (layer3_outputs(3161)) and not (layer3_outputs(5099));
    layer4_outputs(3266) <= not((layer3_outputs(3071)) or (layer3_outputs(2292)));
    layer4_outputs(3267) <= not(layer3_outputs(2117)) or (layer3_outputs(4536));
    layer4_outputs(3268) <= not(layer3_outputs(687)) or (layer3_outputs(4912));
    layer4_outputs(3269) <= '0';
    layer4_outputs(3270) <= '1';
    layer4_outputs(3271) <= layer3_outputs(698);
    layer4_outputs(3272) <= (layer3_outputs(2860)) xor (layer3_outputs(348));
    layer4_outputs(3273) <= '0';
    layer4_outputs(3274) <= layer3_outputs(1803);
    layer4_outputs(3275) <= '1';
    layer4_outputs(3276) <= '0';
    layer4_outputs(3277) <= (layer3_outputs(4111)) and not (layer3_outputs(426));
    layer4_outputs(3278) <= '0';
    layer4_outputs(3279) <= not(layer3_outputs(3411));
    layer4_outputs(3280) <= '1';
    layer4_outputs(3281) <= (layer3_outputs(1139)) and not (layer3_outputs(170));
    layer4_outputs(3282) <= (layer3_outputs(3896)) and (layer3_outputs(2871));
    layer4_outputs(3283) <= (layer3_outputs(1583)) xor (layer3_outputs(3549));
    layer4_outputs(3284) <= '1';
    layer4_outputs(3285) <= '1';
    layer4_outputs(3286) <= not((layer3_outputs(219)) or (layer3_outputs(870)));
    layer4_outputs(3287) <= not((layer3_outputs(4101)) or (layer3_outputs(1345)));
    layer4_outputs(3288) <= not(layer3_outputs(560));
    layer4_outputs(3289) <= '0';
    layer4_outputs(3290) <= not(layer3_outputs(3429)) or (layer3_outputs(4614));
    layer4_outputs(3291) <= not(layer3_outputs(2553)) or (layer3_outputs(2200));
    layer4_outputs(3292) <= (layer3_outputs(3327)) and (layer3_outputs(2807));
    layer4_outputs(3293) <= '0';
    layer4_outputs(3294) <= not(layer3_outputs(1770)) or (layer3_outputs(3095));
    layer4_outputs(3295) <= not(layer3_outputs(4072));
    layer4_outputs(3296) <= not(layer3_outputs(781));
    layer4_outputs(3297) <= (layer3_outputs(4010)) and not (layer3_outputs(2125));
    layer4_outputs(3298) <= layer3_outputs(4686);
    layer4_outputs(3299) <= layer3_outputs(4329);
    layer4_outputs(3300) <= not((layer3_outputs(1650)) and (layer3_outputs(3028)));
    layer4_outputs(3301) <= (layer3_outputs(1593)) xor (layer3_outputs(3539));
    layer4_outputs(3302) <= not((layer3_outputs(2258)) or (layer3_outputs(3197)));
    layer4_outputs(3303) <= layer3_outputs(1291);
    layer4_outputs(3304) <= layer3_outputs(2503);
    layer4_outputs(3305) <= not(layer3_outputs(4547)) or (layer3_outputs(2430));
    layer4_outputs(3306) <= not(layer3_outputs(2358));
    layer4_outputs(3307) <= not(layer3_outputs(1242)) or (layer3_outputs(3935));
    layer4_outputs(3308) <= '0';
    layer4_outputs(3309) <= layer3_outputs(1511);
    layer4_outputs(3310) <= not((layer3_outputs(613)) and (layer3_outputs(4244)));
    layer4_outputs(3311) <= not((layer3_outputs(4253)) and (layer3_outputs(4592)));
    layer4_outputs(3312) <= '0';
    layer4_outputs(3313) <= (layer3_outputs(2334)) and not (layer3_outputs(815));
    layer4_outputs(3314) <= not((layer3_outputs(1718)) or (layer3_outputs(4255)));
    layer4_outputs(3315) <= not(layer3_outputs(125));
    layer4_outputs(3316) <= (layer3_outputs(3048)) and (layer3_outputs(3320));
    layer4_outputs(3317) <= layer3_outputs(1537);
    layer4_outputs(3318) <= '1';
    layer4_outputs(3319) <= '1';
    layer4_outputs(3320) <= '0';
    layer4_outputs(3321) <= (layer3_outputs(203)) and not (layer3_outputs(4798));
    layer4_outputs(3322) <= (layer3_outputs(5006)) and not (layer3_outputs(1700));
    layer4_outputs(3323) <= layer3_outputs(3047);
    layer4_outputs(3324) <= (layer3_outputs(4126)) and (layer3_outputs(4984));
    layer4_outputs(3325) <= (layer3_outputs(775)) and not (layer3_outputs(4513));
    layer4_outputs(3326) <= '1';
    layer4_outputs(3327) <= not(layer3_outputs(1634));
    layer4_outputs(3328) <= not(layer3_outputs(1786)) or (layer3_outputs(4934));
    layer4_outputs(3329) <= (layer3_outputs(3125)) and (layer3_outputs(4992));
    layer4_outputs(3330) <= (layer3_outputs(4316)) and (layer3_outputs(3716));
    layer4_outputs(3331) <= '0';
    layer4_outputs(3332) <= not(layer3_outputs(1750));
    layer4_outputs(3333) <= not(layer3_outputs(4966));
    layer4_outputs(3334) <= '0';
    layer4_outputs(3335) <= '0';
    layer4_outputs(3336) <= not((layer3_outputs(518)) or (layer3_outputs(204)));
    layer4_outputs(3337) <= not((layer3_outputs(3381)) and (layer3_outputs(182)));
    layer4_outputs(3338) <= '0';
    layer4_outputs(3339) <= layer3_outputs(430);
    layer4_outputs(3340) <= (layer3_outputs(4629)) or (layer3_outputs(2656));
    layer4_outputs(3341) <= (layer3_outputs(403)) and not (layer3_outputs(4503));
    layer4_outputs(3342) <= not(layer3_outputs(2908));
    layer4_outputs(3343) <= layer3_outputs(686);
    layer4_outputs(3344) <= '1';
    layer4_outputs(3345) <= not(layer3_outputs(2460));
    layer4_outputs(3346) <= (layer3_outputs(3228)) and not (layer3_outputs(2875));
    layer4_outputs(3347) <= (layer3_outputs(3873)) and not (layer3_outputs(1704));
    layer4_outputs(3348) <= not(layer3_outputs(5095)) or (layer3_outputs(4098));
    layer4_outputs(3349) <= (layer3_outputs(5074)) and not (layer3_outputs(2860));
    layer4_outputs(3350) <= not(layer3_outputs(2053));
    layer4_outputs(3351) <= not((layer3_outputs(2385)) and (layer3_outputs(1686)));
    layer4_outputs(3352) <= layer3_outputs(3230);
    layer4_outputs(3353) <= (layer3_outputs(3668)) or (layer3_outputs(4354));
    layer4_outputs(3354) <= (layer3_outputs(1999)) and not (layer3_outputs(2434));
    layer4_outputs(3355) <= '1';
    layer4_outputs(3356) <= not(layer3_outputs(2178)) or (layer3_outputs(1321));
    layer4_outputs(3357) <= (layer3_outputs(3281)) and not (layer3_outputs(444));
    layer4_outputs(3358) <= not((layer3_outputs(5106)) and (layer3_outputs(3814)));
    layer4_outputs(3359) <= layer3_outputs(4031);
    layer4_outputs(3360) <= not(layer3_outputs(3360)) or (layer3_outputs(4873));
    layer4_outputs(3361) <= (layer3_outputs(334)) and not (layer3_outputs(3877));
    layer4_outputs(3362) <= (layer3_outputs(3826)) and not (layer3_outputs(4609));
    layer4_outputs(3363) <= not(layer3_outputs(3498)) or (layer3_outputs(3591));
    layer4_outputs(3364) <= '0';
    layer4_outputs(3365) <= layer3_outputs(2420);
    layer4_outputs(3366) <= not(layer3_outputs(2074)) or (layer3_outputs(1703));
    layer4_outputs(3367) <= not((layer3_outputs(540)) or (layer3_outputs(1676)));
    layer4_outputs(3368) <= not(layer3_outputs(1993)) or (layer3_outputs(4107));
    layer4_outputs(3369) <= not(layer3_outputs(234));
    layer4_outputs(3370) <= not(layer3_outputs(283));
    layer4_outputs(3371) <= '0';
    layer4_outputs(3372) <= not((layer3_outputs(4079)) or (layer3_outputs(4628)));
    layer4_outputs(3373) <= layer3_outputs(4168);
    layer4_outputs(3374) <= not(layer3_outputs(2617));
    layer4_outputs(3375) <= not((layer3_outputs(3437)) and (layer3_outputs(801)));
    layer4_outputs(3376) <= not(layer3_outputs(2815));
    layer4_outputs(3377) <= not((layer3_outputs(3882)) xor (layer3_outputs(2140)));
    layer4_outputs(3378) <= (layer3_outputs(3262)) and not (layer3_outputs(1436));
    layer4_outputs(3379) <= (layer3_outputs(4501)) or (layer3_outputs(4641));
    layer4_outputs(3380) <= not((layer3_outputs(1782)) or (layer3_outputs(4550)));
    layer4_outputs(3381) <= layer3_outputs(3338);
    layer4_outputs(3382) <= (layer3_outputs(2544)) and (layer3_outputs(4823));
    layer4_outputs(3383) <= not(layer3_outputs(4430)) or (layer3_outputs(947));
    layer4_outputs(3384) <= not(layer3_outputs(1971)) or (layer3_outputs(3035));
    layer4_outputs(3385) <= layer3_outputs(1501);
    layer4_outputs(3386) <= (layer3_outputs(1909)) and not (layer3_outputs(3615));
    layer4_outputs(3387) <= (layer3_outputs(3075)) and not (layer3_outputs(3561));
    layer4_outputs(3388) <= layer3_outputs(2363);
    layer4_outputs(3389) <= not(layer3_outputs(4124));
    layer4_outputs(3390) <= layer3_outputs(3866);
    layer4_outputs(3391) <= not(layer3_outputs(549));
    layer4_outputs(3392) <= layer3_outputs(2757);
    layer4_outputs(3393) <= not(layer3_outputs(1726));
    layer4_outputs(3394) <= (layer3_outputs(3183)) or (layer3_outputs(3026));
    layer4_outputs(3395) <= (layer3_outputs(528)) and not (layer3_outputs(299));
    layer4_outputs(3396) <= (layer3_outputs(1244)) and not (layer3_outputs(1956));
    layer4_outputs(3397) <= not(layer3_outputs(3048)) or (layer3_outputs(1153));
    layer4_outputs(3398) <= '1';
    layer4_outputs(3399) <= '0';
    layer4_outputs(3400) <= layer3_outputs(1373);
    layer4_outputs(3401) <= not((layer3_outputs(4207)) or (layer3_outputs(1729)));
    layer4_outputs(3402) <= (layer3_outputs(4011)) and (layer3_outputs(3714));
    layer4_outputs(3403) <= (layer3_outputs(533)) and (layer3_outputs(550));
    layer4_outputs(3404) <= (layer3_outputs(4889)) and not (layer3_outputs(3853));
    layer4_outputs(3405) <= '1';
    layer4_outputs(3406) <= not((layer3_outputs(3361)) and (layer3_outputs(4669)));
    layer4_outputs(3407) <= (layer3_outputs(3903)) and (layer3_outputs(2167));
    layer4_outputs(3408) <= not((layer3_outputs(2386)) and (layer3_outputs(2077)));
    layer4_outputs(3409) <= not((layer3_outputs(3719)) and (layer3_outputs(2297)));
    layer4_outputs(3410) <= not((layer3_outputs(4916)) or (layer3_outputs(2382)));
    layer4_outputs(3411) <= not(layer3_outputs(810));
    layer4_outputs(3412) <= (layer3_outputs(1589)) and not (layer3_outputs(4796));
    layer4_outputs(3413) <= layer3_outputs(4514);
    layer4_outputs(3414) <= '0';
    layer4_outputs(3415) <= not(layer3_outputs(2062)) or (layer3_outputs(2615));
    layer4_outputs(3416) <= not(layer3_outputs(3273)) or (layer3_outputs(193));
    layer4_outputs(3417) <= not(layer3_outputs(3436)) or (layer3_outputs(66));
    layer4_outputs(3418) <= (layer3_outputs(2049)) and not (layer3_outputs(4859));
    layer4_outputs(3419) <= '0';
    layer4_outputs(3420) <= not((layer3_outputs(2193)) and (layer3_outputs(2144)));
    layer4_outputs(3421) <= layer3_outputs(2221);
    layer4_outputs(3422) <= not(layer3_outputs(702)) or (layer3_outputs(4744));
    layer4_outputs(3423) <= not(layer3_outputs(949));
    layer4_outputs(3424) <= not((layer3_outputs(3956)) and (layer3_outputs(2754)));
    layer4_outputs(3425) <= '0';
    layer4_outputs(3426) <= (layer3_outputs(1274)) and not (layer3_outputs(4661));
    layer4_outputs(3427) <= layer3_outputs(1212);
    layer4_outputs(3428) <= not(layer3_outputs(1342)) or (layer3_outputs(5095));
    layer4_outputs(3429) <= layer3_outputs(1239);
    layer4_outputs(3430) <= not((layer3_outputs(4890)) or (layer3_outputs(1116)));
    layer4_outputs(3431) <= '0';
    layer4_outputs(3432) <= not(layer3_outputs(1044));
    layer4_outputs(3433) <= (layer3_outputs(4115)) and (layer3_outputs(1063));
    layer4_outputs(3434) <= (layer3_outputs(3721)) and not (layer3_outputs(4650));
    layer4_outputs(3435) <= not(layer3_outputs(3867)) or (layer3_outputs(1666));
    layer4_outputs(3436) <= layer3_outputs(3420);
    layer4_outputs(3437) <= '1';
    layer4_outputs(3438) <= (layer3_outputs(236)) and (layer3_outputs(785));
    layer4_outputs(3439) <= not(layer3_outputs(3684)) or (layer3_outputs(4561));
    layer4_outputs(3440) <= '0';
    layer4_outputs(3441) <= not(layer3_outputs(3598));
    layer4_outputs(3442) <= (layer3_outputs(4732)) and (layer3_outputs(1932));
    layer4_outputs(3443) <= layer3_outputs(1298);
    layer4_outputs(3444) <= layer3_outputs(4040);
    layer4_outputs(3445) <= not(layer3_outputs(3778));
    layer4_outputs(3446) <= not(layer3_outputs(152)) or (layer3_outputs(4463));
    layer4_outputs(3447) <= (layer3_outputs(644)) and (layer3_outputs(794));
    layer4_outputs(3448) <= not(layer3_outputs(1306));
    layer4_outputs(3449) <= '0';
    layer4_outputs(3450) <= not(layer3_outputs(2738)) or (layer3_outputs(4942));
    layer4_outputs(3451) <= layer3_outputs(689);
    layer4_outputs(3452) <= '0';
    layer4_outputs(3453) <= (layer3_outputs(112)) and (layer3_outputs(4490));
    layer4_outputs(3454) <= not((layer3_outputs(4764)) and (layer3_outputs(1324)));
    layer4_outputs(3455) <= not(layer3_outputs(3362)) or (layer3_outputs(34));
    layer4_outputs(3456) <= not(layer3_outputs(2070));
    layer4_outputs(3457) <= not((layer3_outputs(4612)) or (layer3_outputs(2159)));
    layer4_outputs(3458) <= (layer3_outputs(2842)) and not (layer3_outputs(4833));
    layer4_outputs(3459) <= not((layer3_outputs(72)) and (layer3_outputs(2430)));
    layer4_outputs(3460) <= not(layer3_outputs(3225));
    layer4_outputs(3461) <= not(layer3_outputs(3244));
    layer4_outputs(3462) <= '1';
    layer4_outputs(3463) <= not(layer3_outputs(1903)) or (layer3_outputs(3384));
    layer4_outputs(3464) <= not(layer3_outputs(30));
    layer4_outputs(3465) <= layer3_outputs(3771);
    layer4_outputs(3466) <= (layer3_outputs(2380)) or (layer3_outputs(2642));
    layer4_outputs(3467) <= layer3_outputs(4290);
    layer4_outputs(3468) <= (layer3_outputs(3929)) xor (layer3_outputs(3834));
    layer4_outputs(3469) <= not(layer3_outputs(8)) or (layer3_outputs(4708));
    layer4_outputs(3470) <= (layer3_outputs(4868)) and not (layer3_outputs(1031));
    layer4_outputs(3471) <= not(layer3_outputs(615));
    layer4_outputs(3472) <= not(layer3_outputs(685)) or (layer3_outputs(2128));
    layer4_outputs(3473) <= not(layer3_outputs(1006));
    layer4_outputs(3474) <= layer3_outputs(4974);
    layer4_outputs(3475) <= (layer3_outputs(4328)) and not (layer3_outputs(5059));
    layer4_outputs(3476) <= (layer3_outputs(4351)) and not (layer3_outputs(209));
    layer4_outputs(3477) <= layer3_outputs(2200);
    layer4_outputs(3478) <= (layer3_outputs(1415)) and not (layer3_outputs(3146));
    layer4_outputs(3479) <= not((layer3_outputs(1943)) xor (layer3_outputs(281)));
    layer4_outputs(3480) <= not(layer3_outputs(1944));
    layer4_outputs(3481) <= not((layer3_outputs(4396)) and (layer3_outputs(4135)));
    layer4_outputs(3482) <= '1';
    layer4_outputs(3483) <= '1';
    layer4_outputs(3484) <= not(layer3_outputs(2150)) or (layer3_outputs(3953));
    layer4_outputs(3485) <= (layer3_outputs(2634)) xor (layer3_outputs(4972));
    layer4_outputs(3486) <= (layer3_outputs(2164)) and not (layer3_outputs(17));
    layer4_outputs(3487) <= (layer3_outputs(2057)) and not (layer3_outputs(2596));
    layer4_outputs(3488) <= (layer3_outputs(4479)) and not (layer3_outputs(1151));
    layer4_outputs(3489) <= not(layer3_outputs(2077));
    layer4_outputs(3490) <= not((layer3_outputs(4892)) and (layer3_outputs(3940)));
    layer4_outputs(3491) <= (layer3_outputs(2815)) or (layer3_outputs(3823));
    layer4_outputs(3492) <= not((layer3_outputs(482)) or (layer3_outputs(2493)));
    layer4_outputs(3493) <= not(layer3_outputs(4325));
    layer4_outputs(3494) <= layer3_outputs(2663);
    layer4_outputs(3495) <= not(layer3_outputs(2781));
    layer4_outputs(3496) <= (layer3_outputs(5097)) and not (layer3_outputs(4902));
    layer4_outputs(3497) <= (layer3_outputs(239)) and (layer3_outputs(2324));
    layer4_outputs(3498) <= (layer3_outputs(3712)) and (layer3_outputs(2421));
    layer4_outputs(3499) <= not((layer3_outputs(576)) or (layer3_outputs(987)));
    layer4_outputs(3500) <= '1';
    layer4_outputs(3501) <= layer3_outputs(2250);
    layer4_outputs(3502) <= not(layer3_outputs(4734));
    layer4_outputs(3503) <= not(layer3_outputs(4325)) or (layer3_outputs(4174));
    layer4_outputs(3504) <= layer3_outputs(1112);
    layer4_outputs(3505) <= (layer3_outputs(2059)) xor (layer3_outputs(1199));
    layer4_outputs(3506) <= not(layer3_outputs(2176));
    layer4_outputs(3507) <= layer3_outputs(3714);
    layer4_outputs(3508) <= (layer3_outputs(1510)) or (layer3_outputs(4002));
    layer4_outputs(3509) <= not((layer3_outputs(4119)) or (layer3_outputs(1276)));
    layer4_outputs(3510) <= (layer3_outputs(3902)) and not (layer3_outputs(4806));
    layer4_outputs(3511) <= '1';
    layer4_outputs(3512) <= layer3_outputs(2347);
    layer4_outputs(3513) <= layer3_outputs(94);
    layer4_outputs(3514) <= not((layer3_outputs(638)) and (layer3_outputs(1793)));
    layer4_outputs(3515) <= (layer3_outputs(433)) and not (layer3_outputs(1410));
    layer4_outputs(3516) <= not(layer3_outputs(2004));
    layer4_outputs(3517) <= (layer3_outputs(3560)) and not (layer3_outputs(1709));
    layer4_outputs(3518) <= not((layer3_outputs(5049)) or (layer3_outputs(3466)));
    layer4_outputs(3519) <= '0';
    layer4_outputs(3520) <= not(layer3_outputs(895));
    layer4_outputs(3521) <= '0';
    layer4_outputs(3522) <= layer3_outputs(3191);
    layer4_outputs(3523) <= (layer3_outputs(4963)) and not (layer3_outputs(4028));
    layer4_outputs(3524) <= (layer3_outputs(4230)) and (layer3_outputs(716));
    layer4_outputs(3525) <= not(layer3_outputs(701)) or (layer3_outputs(109));
    layer4_outputs(3526) <= layer3_outputs(1752);
    layer4_outputs(3527) <= '0';
    layer4_outputs(3528) <= not((layer3_outputs(2479)) or (layer3_outputs(1159)));
    layer4_outputs(3529) <= not(layer3_outputs(760));
    layer4_outputs(3530) <= layer3_outputs(2182);
    layer4_outputs(3531) <= not((layer3_outputs(4221)) or (layer3_outputs(915)));
    layer4_outputs(3532) <= (layer3_outputs(1912)) and not (layer3_outputs(2471));
    layer4_outputs(3533) <= (layer3_outputs(3999)) and not (layer3_outputs(1833));
    layer4_outputs(3534) <= '1';
    layer4_outputs(3535) <= '1';
    layer4_outputs(3536) <= not((layer3_outputs(1455)) and (layer3_outputs(3480)));
    layer4_outputs(3537) <= not(layer3_outputs(633)) or (layer3_outputs(4563));
    layer4_outputs(3538) <= '1';
    layer4_outputs(3539) <= not((layer3_outputs(4772)) or (layer3_outputs(3594)));
    layer4_outputs(3540) <= (layer3_outputs(1056)) and not (layer3_outputs(949));
    layer4_outputs(3541) <= (layer3_outputs(1420)) xor (layer3_outputs(466));
    layer4_outputs(3542) <= (layer3_outputs(469)) or (layer3_outputs(1915));
    layer4_outputs(3543) <= not((layer3_outputs(3764)) or (layer3_outputs(2237)));
    layer4_outputs(3544) <= (layer3_outputs(696)) and (layer3_outputs(2203));
    layer4_outputs(3545) <= '1';
    layer4_outputs(3546) <= (layer3_outputs(2403)) or (layer3_outputs(2487));
    layer4_outputs(3547) <= '1';
    layer4_outputs(3548) <= (layer3_outputs(3728)) and not (layer3_outputs(4232));
    layer4_outputs(3549) <= (layer3_outputs(1951)) xor (layer3_outputs(4728));
    layer4_outputs(3550) <= layer3_outputs(2928);
    layer4_outputs(3551) <= not(layer3_outputs(2716)) or (layer3_outputs(2289));
    layer4_outputs(3552) <= not(layer3_outputs(982)) or (layer3_outputs(1094));
    layer4_outputs(3553) <= layer3_outputs(4992);
    layer4_outputs(3554) <= layer3_outputs(1730);
    layer4_outputs(3555) <= (layer3_outputs(4593)) and not (layer3_outputs(60));
    layer4_outputs(3556) <= (layer3_outputs(1469)) and not (layer3_outputs(3828));
    layer4_outputs(3557) <= not(layer3_outputs(362));
    layer4_outputs(3558) <= layer3_outputs(4749);
    layer4_outputs(3559) <= (layer3_outputs(201)) or (layer3_outputs(842));
    layer4_outputs(3560) <= layer3_outputs(673);
    layer4_outputs(3561) <= not((layer3_outputs(3855)) and (layer3_outputs(1876)));
    layer4_outputs(3562) <= not(layer3_outputs(916));
    layer4_outputs(3563) <= not((layer3_outputs(1629)) or (layer3_outputs(3957)));
    layer4_outputs(3564) <= not((layer3_outputs(4404)) and (layer3_outputs(1297)));
    layer4_outputs(3565) <= not(layer3_outputs(4432));
    layer4_outputs(3566) <= not((layer3_outputs(361)) or (layer3_outputs(4264)));
    layer4_outputs(3567) <= (layer3_outputs(1257)) and (layer3_outputs(4157));
    layer4_outputs(3568) <= (layer3_outputs(3899)) and (layer3_outputs(3086));
    layer4_outputs(3569) <= (layer3_outputs(4505)) and not (layer3_outputs(4821));
    layer4_outputs(3570) <= not(layer3_outputs(3859)) or (layer3_outputs(2135));
    layer4_outputs(3571) <= (layer3_outputs(2235)) and not (layer3_outputs(3349));
    layer4_outputs(3572) <= not(layer3_outputs(2226));
    layer4_outputs(3573) <= not(layer3_outputs(4584)) or (layer3_outputs(4676));
    layer4_outputs(3574) <= '1';
    layer4_outputs(3575) <= not(layer3_outputs(4828)) or (layer3_outputs(3906));
    layer4_outputs(3576) <= (layer3_outputs(2964)) or (layer3_outputs(779));
    layer4_outputs(3577) <= (layer3_outputs(2943)) or (layer3_outputs(4988));
    layer4_outputs(3578) <= '0';
    layer4_outputs(3579) <= not(layer3_outputs(1080));
    layer4_outputs(3580) <= layer3_outputs(4263);
    layer4_outputs(3581) <= not(layer3_outputs(2119)) or (layer3_outputs(3068));
    layer4_outputs(3582) <= not(layer3_outputs(206));
    layer4_outputs(3583) <= not(layer3_outputs(1013));
    layer4_outputs(3584) <= not(layer3_outputs(1563)) or (layer3_outputs(3169));
    layer4_outputs(3585) <= not(layer3_outputs(742));
    layer4_outputs(3586) <= (layer3_outputs(257)) xor (layer3_outputs(97));
    layer4_outputs(3587) <= layer3_outputs(2379);
    layer4_outputs(3588) <= not(layer3_outputs(114));
    layer4_outputs(3589) <= layer3_outputs(2774);
    layer4_outputs(3590) <= (layer3_outputs(114)) and not (layer3_outputs(3451));
    layer4_outputs(3591) <= '1';
    layer4_outputs(3592) <= '0';
    layer4_outputs(3593) <= (layer3_outputs(1231)) or (layer3_outputs(1068));
    layer4_outputs(3594) <= not(layer3_outputs(2007)) or (layer3_outputs(3738));
    layer4_outputs(3595) <= layer3_outputs(1078);
    layer4_outputs(3596) <= layer3_outputs(3942);
    layer4_outputs(3597) <= not(layer3_outputs(4905)) or (layer3_outputs(4289));
    layer4_outputs(3598) <= not((layer3_outputs(4174)) xor (layer3_outputs(1681)));
    layer4_outputs(3599) <= not(layer3_outputs(4692));
    layer4_outputs(3600) <= '1';
    layer4_outputs(3601) <= '0';
    layer4_outputs(3602) <= layer3_outputs(4660);
    layer4_outputs(3603) <= '0';
    layer4_outputs(3604) <= (layer3_outputs(2353)) and not (layer3_outputs(1303));
    layer4_outputs(3605) <= layer3_outputs(1358);
    layer4_outputs(3606) <= not(layer3_outputs(4270));
    layer4_outputs(3607) <= '0';
    layer4_outputs(3608) <= '0';
    layer4_outputs(3609) <= not(layer3_outputs(2344));
    layer4_outputs(3610) <= (layer3_outputs(1085)) and not (layer3_outputs(2877));
    layer4_outputs(3611) <= (layer3_outputs(1037)) and not (layer3_outputs(3906));
    layer4_outputs(3612) <= layer3_outputs(955);
    layer4_outputs(3613) <= not((layer3_outputs(4550)) or (layer3_outputs(4735)));
    layer4_outputs(3614) <= (layer3_outputs(3220)) and (layer3_outputs(4616));
    layer4_outputs(3615) <= not(layer3_outputs(3348));
    layer4_outputs(3616) <= '0';
    layer4_outputs(3617) <= layer3_outputs(3510);
    layer4_outputs(3618) <= (layer3_outputs(691)) or (layer3_outputs(1177));
    layer4_outputs(3619) <= '0';
    layer4_outputs(3620) <= (layer3_outputs(553)) and (layer3_outputs(3343));
    layer4_outputs(3621) <= (layer3_outputs(893)) and not (layer3_outputs(1340));
    layer4_outputs(3622) <= not(layer3_outputs(2089));
    layer4_outputs(3623) <= (layer3_outputs(2204)) and (layer3_outputs(3364));
    layer4_outputs(3624) <= '1';
    layer4_outputs(3625) <= '0';
    layer4_outputs(3626) <= not((layer3_outputs(2177)) xor (layer3_outputs(3994)));
    layer4_outputs(3627) <= not(layer3_outputs(263)) or (layer3_outputs(4617));
    layer4_outputs(3628) <= '1';
    layer4_outputs(3629) <= (layer3_outputs(4723)) and not (layer3_outputs(4303));
    layer4_outputs(3630) <= not((layer3_outputs(4578)) and (layer3_outputs(2426)));
    layer4_outputs(3631) <= not(layer3_outputs(1071));
    layer4_outputs(3632) <= '1';
    layer4_outputs(3633) <= layer3_outputs(2461);
    layer4_outputs(3634) <= '0';
    layer4_outputs(3635) <= '1';
    layer4_outputs(3636) <= not(layer3_outputs(4991)) or (layer3_outputs(3937));
    layer4_outputs(3637) <= not(layer3_outputs(5045)) or (layer3_outputs(4099));
    layer4_outputs(3638) <= (layer3_outputs(3798)) or (layer3_outputs(1217));
    layer4_outputs(3639) <= layer3_outputs(211);
    layer4_outputs(3640) <= '1';
    layer4_outputs(3641) <= (layer3_outputs(3950)) and not (layer3_outputs(3535));
    layer4_outputs(3642) <= not((layer3_outputs(4396)) and (layer3_outputs(1167)));
    layer4_outputs(3643) <= (layer3_outputs(341)) or (layer3_outputs(739));
    layer4_outputs(3644) <= not((layer3_outputs(773)) or (layer3_outputs(2869)));
    layer4_outputs(3645) <= layer3_outputs(2464);
    layer4_outputs(3646) <= '0';
    layer4_outputs(3647) <= not((layer3_outputs(2740)) xor (layer3_outputs(4727)));
    layer4_outputs(3648) <= not(layer3_outputs(1701));
    layer4_outputs(3649) <= not(layer3_outputs(1297)) or (layer3_outputs(3138));
    layer4_outputs(3650) <= (layer3_outputs(1)) and (layer3_outputs(3633));
    layer4_outputs(3651) <= layer3_outputs(2766);
    layer4_outputs(3652) <= layer3_outputs(4465);
    layer4_outputs(3653) <= '0';
    layer4_outputs(3654) <= '1';
    layer4_outputs(3655) <= '0';
    layer4_outputs(3656) <= (layer3_outputs(4182)) and not (layer3_outputs(1825));
    layer4_outputs(3657) <= (layer3_outputs(3151)) xor (layer3_outputs(3522));
    layer4_outputs(3658) <= layer3_outputs(5023);
    layer4_outputs(3659) <= not(layer3_outputs(128));
    layer4_outputs(3660) <= not(layer3_outputs(4082)) or (layer3_outputs(2294));
    layer4_outputs(3661) <= (layer3_outputs(5004)) and (layer3_outputs(884));
    layer4_outputs(3662) <= not(layer3_outputs(2368));
    layer4_outputs(3663) <= not(layer3_outputs(1038)) or (layer3_outputs(709));
    layer4_outputs(3664) <= not(layer3_outputs(4422)) or (layer3_outputs(4920));
    layer4_outputs(3665) <= '0';
    layer4_outputs(3666) <= (layer3_outputs(2427)) and not (layer3_outputs(3386));
    layer4_outputs(3667) <= not((layer3_outputs(808)) and (layer3_outputs(569)));
    layer4_outputs(3668) <= '1';
    layer4_outputs(3669) <= '0';
    layer4_outputs(3670) <= not((layer3_outputs(3762)) and (layer3_outputs(2885)));
    layer4_outputs(3671) <= not(layer3_outputs(3556)) or (layer3_outputs(1578));
    layer4_outputs(3672) <= not(layer3_outputs(4987));
    layer4_outputs(3673) <= not((layer3_outputs(1965)) and (layer3_outputs(2744)));
    layer4_outputs(3674) <= (layer3_outputs(4864)) or (layer3_outputs(679));
    layer4_outputs(3675) <= (layer3_outputs(3392)) and (layer3_outputs(4564));
    layer4_outputs(3676) <= not((layer3_outputs(3919)) and (layer3_outputs(2010)));
    layer4_outputs(3677) <= not(layer3_outputs(3441));
    layer4_outputs(3678) <= '1';
    layer4_outputs(3679) <= (layer3_outputs(4470)) xor (layer3_outputs(395));
    layer4_outputs(3680) <= not((layer3_outputs(1006)) or (layer3_outputs(4309)));
    layer4_outputs(3681) <= not(layer3_outputs(4679));
    layer4_outputs(3682) <= '1';
    layer4_outputs(3683) <= not(layer3_outputs(622));
    layer4_outputs(3684) <= (layer3_outputs(2698)) xor (layer3_outputs(4803));
    layer4_outputs(3685) <= '0';
    layer4_outputs(3686) <= layer3_outputs(543);
    layer4_outputs(3687) <= not(layer3_outputs(3857));
    layer4_outputs(3688) <= not((layer3_outputs(1107)) or (layer3_outputs(388)));
    layer4_outputs(3689) <= '0';
    layer4_outputs(3690) <= (layer3_outputs(4965)) and not (layer3_outputs(3451));
    layer4_outputs(3691) <= not(layer3_outputs(4159)) or (layer3_outputs(238));
    layer4_outputs(3692) <= layer3_outputs(3671);
    layer4_outputs(3693) <= not(layer3_outputs(2796)) or (layer3_outputs(1568));
    layer4_outputs(3694) <= not((layer3_outputs(4046)) and (layer3_outputs(4565)));
    layer4_outputs(3695) <= (layer3_outputs(2523)) and not (layer3_outputs(567));
    layer4_outputs(3696) <= not(layer3_outputs(3301)) or (layer3_outputs(2323));
    layer4_outputs(3697) <= layer3_outputs(3926);
    layer4_outputs(3698) <= layer3_outputs(737);
    layer4_outputs(3699) <= layer3_outputs(5028);
    layer4_outputs(3700) <= (layer3_outputs(2534)) or (layer3_outputs(4025));
    layer4_outputs(3701) <= (layer3_outputs(2345)) and (layer3_outputs(183));
    layer4_outputs(3702) <= layer3_outputs(836);
    layer4_outputs(3703) <= not(layer3_outputs(5041));
    layer4_outputs(3704) <= '1';
    layer4_outputs(3705) <= not(layer3_outputs(258)) or (layer3_outputs(1507));
    layer4_outputs(3706) <= (layer3_outputs(826)) and (layer3_outputs(2533));
    layer4_outputs(3707) <= layer3_outputs(1015);
    layer4_outputs(3708) <= not((layer3_outputs(902)) or (layer3_outputs(2988)));
    layer4_outputs(3709) <= not((layer3_outputs(641)) and (layer3_outputs(1903)));
    layer4_outputs(3710) <= (layer3_outputs(3530)) and not (layer3_outputs(4912));
    layer4_outputs(3711) <= not(layer3_outputs(531)) or (layer3_outputs(4140));
    layer4_outputs(3712) <= not((layer3_outputs(3891)) or (layer3_outputs(4881)));
    layer4_outputs(3713) <= not((layer3_outputs(3709)) and (layer3_outputs(4731)));
    layer4_outputs(3714) <= not((layer3_outputs(2867)) and (layer3_outputs(4632)));
    layer4_outputs(3715) <= (layer3_outputs(4944)) and (layer3_outputs(4588));
    layer4_outputs(3716) <= (layer3_outputs(50)) and (layer3_outputs(3390));
    layer4_outputs(3717) <= not((layer3_outputs(2414)) xor (layer3_outputs(2613)));
    layer4_outputs(3718) <= not(layer3_outputs(4826)) or (layer3_outputs(707));
    layer4_outputs(3719) <= not((layer3_outputs(4181)) or (layer3_outputs(1564)));
    layer4_outputs(3720) <= (layer3_outputs(2194)) and not (layer3_outputs(2645));
    layer4_outputs(3721) <= not(layer3_outputs(2330));
    layer4_outputs(3722) <= (layer3_outputs(4995)) and not (layer3_outputs(1877));
    layer4_outputs(3723) <= layer3_outputs(729);
    layer4_outputs(3724) <= not((layer3_outputs(2170)) or (layer3_outputs(962)));
    layer4_outputs(3725) <= (layer3_outputs(3757)) and not (layer3_outputs(3641));
    layer4_outputs(3726) <= layer3_outputs(4835);
    layer4_outputs(3727) <= layer3_outputs(2609);
    layer4_outputs(3728) <= layer3_outputs(2332);
    layer4_outputs(3729) <= not(layer3_outputs(688));
    layer4_outputs(3730) <= not(layer3_outputs(724)) or (layer3_outputs(471));
    layer4_outputs(3731) <= '0';
    layer4_outputs(3732) <= (layer3_outputs(1140)) or (layer3_outputs(1423));
    layer4_outputs(3733) <= not(layer3_outputs(1469));
    layer4_outputs(3734) <= layer3_outputs(2261);
    layer4_outputs(3735) <= not(layer3_outputs(4316)) or (layer3_outputs(345));
    layer4_outputs(3736) <= not(layer3_outputs(4407));
    layer4_outputs(3737) <= not(layer3_outputs(1571)) or (layer3_outputs(31));
    layer4_outputs(3738) <= (layer3_outputs(3692)) and not (layer3_outputs(1580));
    layer4_outputs(3739) <= '0';
    layer4_outputs(3740) <= '0';
    layer4_outputs(3741) <= layer3_outputs(1125);
    layer4_outputs(3742) <= layer3_outputs(3165);
    layer4_outputs(3743) <= not(layer3_outputs(3961)) or (layer3_outputs(1698));
    layer4_outputs(3744) <= layer3_outputs(921);
    layer4_outputs(3745) <= not(layer3_outputs(3217));
    layer4_outputs(3746) <= not((layer3_outputs(4633)) and (layer3_outputs(4871)));
    layer4_outputs(3747) <= not(layer3_outputs(2098)) or (layer3_outputs(746));
    layer4_outputs(3748) <= (layer3_outputs(3037)) and (layer3_outputs(168));
    layer4_outputs(3749) <= (layer3_outputs(3054)) and not (layer3_outputs(2225));
    layer4_outputs(3750) <= (layer3_outputs(4634)) or (layer3_outputs(1734));
    layer4_outputs(3751) <= (layer3_outputs(1281)) and not (layer3_outputs(3252));
    layer4_outputs(3752) <= (layer3_outputs(1523)) and (layer3_outputs(1508));
    layer4_outputs(3753) <= (layer3_outputs(1867)) or (layer3_outputs(5115));
    layer4_outputs(3754) <= not((layer3_outputs(2067)) and (layer3_outputs(2561)));
    layer4_outputs(3755) <= '1';
    layer4_outputs(3756) <= '1';
    layer4_outputs(3757) <= not((layer3_outputs(4646)) or (layer3_outputs(1565)));
    layer4_outputs(3758) <= not(layer3_outputs(3513));
    layer4_outputs(3759) <= (layer3_outputs(1528)) and (layer3_outputs(3195));
    layer4_outputs(3760) <= not(layer3_outputs(1145)) or (layer3_outputs(3142));
    layer4_outputs(3761) <= '1';
    layer4_outputs(3762) <= (layer3_outputs(858)) or (layer3_outputs(4545));
    layer4_outputs(3763) <= not(layer3_outputs(819));
    layer4_outputs(3764) <= not(layer3_outputs(1727)) or (layer3_outputs(4994));
    layer4_outputs(3765) <= '0';
    layer4_outputs(3766) <= not((layer3_outputs(2696)) and (layer3_outputs(3683)));
    layer4_outputs(3767) <= not((layer3_outputs(3358)) xor (layer3_outputs(2614)));
    layer4_outputs(3768) <= '1';
    layer4_outputs(3769) <= not(layer3_outputs(4209)) or (layer3_outputs(2517));
    layer4_outputs(3770) <= not((layer3_outputs(4970)) xor (layer3_outputs(1929)));
    layer4_outputs(3771) <= not(layer3_outputs(1963)) or (layer3_outputs(2347));
    layer4_outputs(3772) <= not(layer3_outputs(2451)) or (layer3_outputs(2202));
    layer4_outputs(3773) <= (layer3_outputs(3645)) and not (layer3_outputs(1976));
    layer4_outputs(3774) <= (layer3_outputs(2250)) and not (layer3_outputs(3881));
    layer4_outputs(3775) <= '0';
    layer4_outputs(3776) <= (layer3_outputs(866)) and (layer3_outputs(4421));
    layer4_outputs(3777) <= (layer3_outputs(4766)) or (layer3_outputs(2879));
    layer4_outputs(3778) <= not((layer3_outputs(2136)) or (layer3_outputs(233)));
    layer4_outputs(3779) <= not(layer3_outputs(970));
    layer4_outputs(3780) <= not((layer3_outputs(2443)) and (layer3_outputs(1008)));
    layer4_outputs(3781) <= (layer3_outputs(4282)) and not (layer3_outputs(1893));
    layer4_outputs(3782) <= (layer3_outputs(546)) and not (layer3_outputs(1147));
    layer4_outputs(3783) <= '0';
    layer4_outputs(3784) <= layer3_outputs(1548);
    layer4_outputs(3785) <= layer3_outputs(240);
    layer4_outputs(3786) <= not((layer3_outputs(3955)) or (layer3_outputs(2798)));
    layer4_outputs(3787) <= layer3_outputs(1177);
    layer4_outputs(3788) <= layer3_outputs(2519);
    layer4_outputs(3789) <= not(layer3_outputs(2835)) or (layer3_outputs(855));
    layer4_outputs(3790) <= '1';
    layer4_outputs(3791) <= not((layer3_outputs(1047)) and (layer3_outputs(2594)));
    layer4_outputs(3792) <= not(layer3_outputs(1760)) or (layer3_outputs(847));
    layer4_outputs(3793) <= '0';
    layer4_outputs(3794) <= '1';
    layer4_outputs(3795) <= not(layer3_outputs(4680));
    layer4_outputs(3796) <= (layer3_outputs(3321)) and (layer3_outputs(2330));
    layer4_outputs(3797) <= '0';
    layer4_outputs(3798) <= (layer3_outputs(3900)) and not (layer3_outputs(4));
    layer4_outputs(3799) <= layer3_outputs(1797);
    layer4_outputs(3800) <= '1';
    layer4_outputs(3801) <= not(layer3_outputs(2719)) or (layer3_outputs(1485));
    layer4_outputs(3802) <= (layer3_outputs(4846)) and not (layer3_outputs(3819));
    layer4_outputs(3803) <= (layer3_outputs(4685)) and not (layer3_outputs(539));
    layer4_outputs(3804) <= (layer3_outputs(1003)) and (layer3_outputs(4377));
    layer4_outputs(3805) <= (layer3_outputs(1556)) xor (layer3_outputs(2282));
    layer4_outputs(3806) <= (layer3_outputs(4310)) and not (layer3_outputs(389));
    layer4_outputs(3807) <= not(layer3_outputs(2266)) or (layer3_outputs(3250));
    layer4_outputs(3808) <= '1';
    layer4_outputs(3809) <= layer3_outputs(715);
    layer4_outputs(3810) <= '1';
    layer4_outputs(3811) <= not((layer3_outputs(979)) and (layer3_outputs(2130)));
    layer4_outputs(3812) <= not(layer3_outputs(2434)) or (layer3_outputs(4891));
    layer4_outputs(3813) <= (layer3_outputs(3400)) and not (layer3_outputs(4759));
    layer4_outputs(3814) <= not(layer3_outputs(2340));
    layer4_outputs(3815) <= not(layer3_outputs(3898));
    layer4_outputs(3816) <= not(layer3_outputs(4223)) or (layer3_outputs(1968));
    layer4_outputs(3817) <= layer3_outputs(844);
    layer4_outputs(3818) <= '1';
    layer4_outputs(3819) <= not(layer3_outputs(2728));
    layer4_outputs(3820) <= (layer3_outputs(1388)) and not (layer3_outputs(1320));
    layer4_outputs(3821) <= '1';
    layer4_outputs(3822) <= layer3_outputs(2489);
    layer4_outputs(3823) <= not((layer3_outputs(1885)) or (layer3_outputs(2180)));
    layer4_outputs(3824) <= layer3_outputs(2073);
    layer4_outputs(3825) <= not((layer3_outputs(4143)) xor (layer3_outputs(4020)));
    layer4_outputs(3826) <= not((layer3_outputs(3928)) and (layer3_outputs(402)));
    layer4_outputs(3827) <= layer3_outputs(2566);
    layer4_outputs(3828) <= (layer3_outputs(2040)) and not (layer3_outputs(1057));
    layer4_outputs(3829) <= not((layer3_outputs(4674)) and (layer3_outputs(4470)));
    layer4_outputs(3830) <= not((layer3_outputs(929)) and (layer3_outputs(213)));
    layer4_outputs(3831) <= '1';
    layer4_outputs(3832) <= not((layer3_outputs(4532)) and (layer3_outputs(5022)));
    layer4_outputs(3833) <= (layer3_outputs(4003)) and not (layer3_outputs(973));
    layer4_outputs(3834) <= not((layer3_outputs(1269)) or (layer3_outputs(774)));
    layer4_outputs(3835) <= not((layer3_outputs(3168)) and (layer3_outputs(525)));
    layer4_outputs(3836) <= (layer3_outputs(1544)) and (layer3_outputs(13));
    layer4_outputs(3837) <= '1';
    layer4_outputs(3838) <= layer3_outputs(4283);
    layer4_outputs(3839) <= not(layer3_outputs(3839)) or (layer3_outputs(2531));
    layer4_outputs(3840) <= not(layer3_outputs(1484));
    layer4_outputs(3841) <= (layer3_outputs(2068)) and not (layer3_outputs(2407));
    layer4_outputs(3842) <= (layer3_outputs(2853)) and not (layer3_outputs(1992));
    layer4_outputs(3843) <= not(layer3_outputs(1519)) or (layer3_outputs(396));
    layer4_outputs(3844) <= (layer3_outputs(981)) and not (layer3_outputs(1875));
    layer4_outputs(3845) <= layer3_outputs(2085);
    layer4_outputs(3846) <= (layer3_outputs(4733)) and (layer3_outputs(2630));
    layer4_outputs(3847) <= (layer3_outputs(4947)) and not (layer3_outputs(2479));
    layer4_outputs(3848) <= (layer3_outputs(1410)) and (layer3_outputs(4481));
    layer4_outputs(3849) <= not(layer3_outputs(4437)) or (layer3_outputs(1434));
    layer4_outputs(3850) <= not(layer3_outputs(4865));
    layer4_outputs(3851) <= (layer3_outputs(2352)) and not (layer3_outputs(317));
    layer4_outputs(3852) <= (layer3_outputs(698)) and not (layer3_outputs(890));
    layer4_outputs(3853) <= layer3_outputs(1058);
    layer4_outputs(3854) <= not((layer3_outputs(3314)) or (layer3_outputs(756)));
    layer4_outputs(3855) <= not(layer3_outputs(1705)) or (layer3_outputs(3732));
    layer4_outputs(3856) <= not(layer3_outputs(2192));
    layer4_outputs(3857) <= not(layer3_outputs(3248));
    layer4_outputs(3858) <= (layer3_outputs(661)) xor (layer3_outputs(86));
    layer4_outputs(3859) <= not((layer3_outputs(3484)) xor (layer3_outputs(1338)));
    layer4_outputs(3860) <= (layer3_outputs(3775)) and (layer3_outputs(1592));
    layer4_outputs(3861) <= (layer3_outputs(535)) and not (layer3_outputs(1259));
    layer4_outputs(3862) <= (layer3_outputs(3583)) and not (layer3_outputs(1822));
    layer4_outputs(3863) <= not(layer3_outputs(4217));
    layer4_outputs(3864) <= '1';
    layer4_outputs(3865) <= not((layer3_outputs(3279)) and (layer3_outputs(2518)));
    layer4_outputs(3866) <= (layer3_outputs(1549)) and not (layer3_outputs(3821));
    layer4_outputs(3867) <= not((layer3_outputs(2192)) and (layer3_outputs(3193)));
    layer4_outputs(3868) <= (layer3_outputs(2851)) and not (layer3_outputs(2647));
    layer4_outputs(3869) <= not(layer3_outputs(3703));
    layer4_outputs(3870) <= not(layer3_outputs(2538));
    layer4_outputs(3871) <= layer3_outputs(3951);
    layer4_outputs(3872) <= not(layer3_outputs(1357));
    layer4_outputs(3873) <= '1';
    layer4_outputs(3874) <= (layer3_outputs(1074)) xor (layer3_outputs(2641));
    layer4_outputs(3875) <= not(layer3_outputs(3103)) or (layer3_outputs(363));
    layer4_outputs(3876) <= (layer3_outputs(3846)) and not (layer3_outputs(1211));
    layer4_outputs(3877) <= layer3_outputs(4142);
    layer4_outputs(3878) <= '0';
    layer4_outputs(3879) <= (layer3_outputs(3333)) and not (layer3_outputs(1025));
    layer4_outputs(3880) <= (layer3_outputs(1846)) xor (layer3_outputs(1255));
    layer4_outputs(3881) <= (layer3_outputs(4849)) or (layer3_outputs(3834));
    layer4_outputs(3882) <= not(layer3_outputs(1741));
    layer4_outputs(3883) <= not(layer3_outputs(568)) or (layer3_outputs(5098));
    layer4_outputs(3884) <= not((layer3_outputs(2028)) xor (layer3_outputs(672)));
    layer4_outputs(3885) <= not(layer3_outputs(372));
    layer4_outputs(3886) <= not((layer3_outputs(3939)) and (layer3_outputs(2690)));
    layer4_outputs(3887) <= not(layer3_outputs(391));
    layer4_outputs(3888) <= '1';
    layer4_outputs(3889) <= (layer3_outputs(4231)) and (layer3_outputs(2272));
    layer4_outputs(3890) <= (layer3_outputs(1444)) and not (layer3_outputs(2783));
    layer4_outputs(3891) <= (layer3_outputs(26)) and not (layer3_outputs(1677));
    layer4_outputs(3892) <= '0';
    layer4_outputs(3893) <= layer3_outputs(2554);
    layer4_outputs(3894) <= not((layer3_outputs(1924)) or (layer3_outputs(3456)));
    layer4_outputs(3895) <= layer3_outputs(3702);
    layer4_outputs(3896) <= not(layer3_outputs(922));
    layer4_outputs(3897) <= (layer3_outputs(1550)) or (layer3_outputs(475));
    layer4_outputs(3898) <= not(layer3_outputs(1597));
    layer4_outputs(3899) <= '1';
    layer4_outputs(3900) <= (layer3_outputs(4330)) or (layer3_outputs(46));
    layer4_outputs(3901) <= layer3_outputs(957);
    layer4_outputs(3902) <= (layer3_outputs(3587)) xor (layer3_outputs(446));
    layer4_outputs(3903) <= (layer3_outputs(1894)) and not (layer3_outputs(4515));
    layer4_outputs(3904) <= not(layer3_outputs(3320)) or (layer3_outputs(360));
    layer4_outputs(3905) <= not(layer3_outputs(143));
    layer4_outputs(3906) <= not((layer3_outputs(1136)) and (layer3_outputs(3447)));
    layer4_outputs(3907) <= layer3_outputs(2930);
    layer4_outputs(3908) <= (layer3_outputs(3649)) and not (layer3_outputs(3901));
    layer4_outputs(3909) <= not((layer3_outputs(2104)) or (layer3_outputs(4845)));
    layer4_outputs(3910) <= not(layer3_outputs(879));
    layer4_outputs(3911) <= not((layer3_outputs(520)) or (layer3_outputs(4133)));
    layer4_outputs(3912) <= not(layer3_outputs(4036)) or (layer3_outputs(4596));
    layer4_outputs(3913) <= not((layer3_outputs(1817)) or (layer3_outputs(3185)));
    layer4_outputs(3914) <= layer3_outputs(155);
    layer4_outputs(3915) <= layer3_outputs(4156);
    layer4_outputs(3916) <= not((layer3_outputs(2694)) or (layer3_outputs(1170)));
    layer4_outputs(3917) <= not((layer3_outputs(699)) or (layer3_outputs(4529)));
    layer4_outputs(3918) <= '1';
    layer4_outputs(3919) <= (layer3_outputs(4292)) and (layer3_outputs(63));
    layer4_outputs(3920) <= not((layer3_outputs(3586)) or (layer3_outputs(4854)));
    layer4_outputs(3921) <= (layer3_outputs(2989)) and not (layer3_outputs(4655));
    layer4_outputs(3922) <= '0';
    layer4_outputs(3923) <= not(layer3_outputs(4838));
    layer4_outputs(3924) <= not((layer3_outputs(3588)) or (layer3_outputs(2730)));
    layer4_outputs(3925) <= '1';
    layer4_outputs(3926) <= (layer3_outputs(1459)) and not (layer3_outputs(4453));
    layer4_outputs(3927) <= not(layer3_outputs(693));
    layer4_outputs(3928) <= (layer3_outputs(982)) and not (layer3_outputs(2526));
    layer4_outputs(3929) <= layer3_outputs(134);
    layer4_outputs(3930) <= not((layer3_outputs(3395)) or (layer3_outputs(4517)));
    layer4_outputs(3931) <= (layer3_outputs(2733)) or (layer3_outputs(2810));
    layer4_outputs(3932) <= (layer3_outputs(4732)) and not (layer3_outputs(2397));
    layer4_outputs(3933) <= layer3_outputs(1565);
    layer4_outputs(3934) <= (layer3_outputs(4773)) and (layer3_outputs(2008));
    layer4_outputs(3935) <= '0';
    layer4_outputs(3936) <= '0';
    layer4_outputs(3937) <= layer3_outputs(4302);
    layer4_outputs(3938) <= not(layer3_outputs(818)) or (layer3_outputs(4610));
    layer4_outputs(3939) <= not(layer3_outputs(4812)) or (layer3_outputs(2395));
    layer4_outputs(3940) <= '0';
    layer4_outputs(3941) <= (layer3_outputs(2870)) and not (layer3_outputs(547));
    layer4_outputs(3942) <= (layer3_outputs(141)) or (layer3_outputs(1571));
    layer4_outputs(3943) <= layer3_outputs(4384);
    layer4_outputs(3944) <= not(layer3_outputs(665));
    layer4_outputs(3945) <= layer3_outputs(2311);
    layer4_outputs(3946) <= not(layer3_outputs(9)) or (layer3_outputs(1566));
    layer4_outputs(3947) <= (layer3_outputs(4614)) and not (layer3_outputs(5089));
    layer4_outputs(3948) <= (layer3_outputs(4091)) and not (layer3_outputs(1367));
    layer4_outputs(3949) <= not(layer3_outputs(3809)) or (layer3_outputs(4932));
    layer4_outputs(3950) <= '0';
    layer4_outputs(3951) <= not(layer3_outputs(5093)) or (layer3_outputs(1619));
    layer4_outputs(3952) <= not(layer3_outputs(697));
    layer4_outputs(3953) <= not(layer3_outputs(3111)) or (layer3_outputs(2748));
    layer4_outputs(3954) <= (layer3_outputs(1503)) or (layer3_outputs(5092));
    layer4_outputs(3955) <= (layer3_outputs(1409)) or (layer3_outputs(2850));
    layer4_outputs(3956) <= not((layer3_outputs(2168)) or (layer3_outputs(5109)));
    layer4_outputs(3957) <= not(layer3_outputs(3297));
    layer4_outputs(3958) <= not((layer3_outputs(3127)) xor (layer3_outputs(1692)));
    layer4_outputs(3959) <= not(layer3_outputs(2386)) or (layer3_outputs(4105));
    layer4_outputs(3960) <= not(layer3_outputs(4287));
    layer4_outputs(3961) <= layer3_outputs(4175);
    layer4_outputs(3962) <= not(layer3_outputs(2295));
    layer4_outputs(3963) <= (layer3_outputs(2036)) xor (layer3_outputs(73));
    layer4_outputs(3964) <= not((layer3_outputs(4233)) or (layer3_outputs(724)));
    layer4_outputs(3965) <= not((layer3_outputs(2579)) or (layer3_outputs(956)));
    layer4_outputs(3966) <= not(layer3_outputs(4322));
    layer4_outputs(3967) <= not(layer3_outputs(854));
    layer4_outputs(3968) <= (layer3_outputs(4026)) and not (layer3_outputs(2197));
    layer4_outputs(3969) <= (layer3_outputs(531)) and not (layer3_outputs(4211));
    layer4_outputs(3970) <= not(layer3_outputs(1773));
    layer4_outputs(3971) <= '1';
    layer4_outputs(3972) <= layer3_outputs(4384);
    layer4_outputs(3973) <= '1';
    layer4_outputs(3974) <= (layer3_outputs(3787)) or (layer3_outputs(1275));
    layer4_outputs(3975) <= '1';
    layer4_outputs(3976) <= not(layer3_outputs(4590));
    layer4_outputs(3977) <= (layer3_outputs(4103)) and (layer3_outputs(3070));
    layer4_outputs(3978) <= not((layer3_outputs(2705)) and (layer3_outputs(1653)));
    layer4_outputs(3979) <= '0';
    layer4_outputs(3980) <= not((layer3_outputs(1969)) or (layer3_outputs(4779)));
    layer4_outputs(3981) <= layer3_outputs(2076);
    layer4_outputs(3982) <= not(layer3_outputs(765));
    layer4_outputs(3983) <= layer3_outputs(532);
    layer4_outputs(3984) <= (layer3_outputs(49)) and (layer3_outputs(2417));
    layer4_outputs(3985) <= (layer3_outputs(2363)) or (layer3_outputs(2843));
    layer4_outputs(3986) <= (layer3_outputs(639)) or (layer3_outputs(2298));
    layer4_outputs(3987) <= '0';
    layer4_outputs(3988) <= not((layer3_outputs(4526)) or (layer3_outputs(4496)));
    layer4_outputs(3989) <= not(layer3_outputs(5008));
    layer4_outputs(3990) <= (layer3_outputs(146)) or (layer3_outputs(3721));
    layer4_outputs(3991) <= not(layer3_outputs(3963));
    layer4_outputs(3992) <= not(layer3_outputs(1457)) or (layer3_outputs(4042));
    layer4_outputs(3993) <= layer3_outputs(1649);
    layer4_outputs(3994) <= not(layer3_outputs(1667)) or (layer3_outputs(3893));
    layer4_outputs(3995) <= layer3_outputs(3954);
    layer4_outputs(3996) <= not(layer3_outputs(4959));
    layer4_outputs(3997) <= layer3_outputs(2082);
    layer4_outputs(3998) <= (layer3_outputs(1239)) and not (layer3_outputs(2979));
    layer4_outputs(3999) <= '1';
    layer4_outputs(4000) <= not(layer3_outputs(105)) or (layer3_outputs(1430));
    layer4_outputs(4001) <= layer3_outputs(3811);
    layer4_outputs(4002) <= (layer3_outputs(3034)) and (layer3_outputs(5114));
    layer4_outputs(4003) <= layer3_outputs(3489);
    layer4_outputs(4004) <= not(layer3_outputs(1070)) or (layer3_outputs(3638));
    layer4_outputs(4005) <= (layer3_outputs(504)) and not (layer3_outputs(4044));
    layer4_outputs(4006) <= layer3_outputs(590);
    layer4_outputs(4007) <= '0';
    layer4_outputs(4008) <= not(layer3_outputs(2016));
    layer4_outputs(4009) <= '1';
    layer4_outputs(4010) <= layer3_outputs(4607);
    layer4_outputs(4011) <= not(layer3_outputs(104)) or (layer3_outputs(2549));
    layer4_outputs(4012) <= layer3_outputs(3244);
    layer4_outputs(4013) <= not((layer3_outputs(3447)) and (layer3_outputs(2173)));
    layer4_outputs(4014) <= not(layer3_outputs(2878));
    layer4_outputs(4015) <= not(layer3_outputs(2066)) or (layer3_outputs(2727));
    layer4_outputs(4016) <= not(layer3_outputs(4569)) or (layer3_outputs(2986));
    layer4_outputs(4017) <= layer3_outputs(754);
    layer4_outputs(4018) <= not(layer3_outputs(3936));
    layer4_outputs(4019) <= layer3_outputs(1003);
    layer4_outputs(4020) <= '1';
    layer4_outputs(4021) <= '0';
    layer4_outputs(4022) <= layer3_outputs(2446);
    layer4_outputs(4023) <= (layer3_outputs(4414)) and (layer3_outputs(3402));
    layer4_outputs(4024) <= not((layer3_outputs(168)) xor (layer3_outputs(3813)));
    layer4_outputs(4025) <= layer3_outputs(435);
    layer4_outputs(4026) <= not(layer3_outputs(3530));
    layer4_outputs(4027) <= (layer3_outputs(408)) and not (layer3_outputs(4480));
    layer4_outputs(4028) <= layer3_outputs(579);
    layer4_outputs(4029) <= layer3_outputs(3539);
    layer4_outputs(4030) <= not(layer3_outputs(1427)) or (layer3_outputs(3712));
    layer4_outputs(4031) <= (layer3_outputs(3108)) and (layer3_outputs(570));
    layer4_outputs(4032) <= not(layer3_outputs(4415));
    layer4_outputs(4033) <= not(layer3_outputs(2770)) or (layer3_outputs(20));
    layer4_outputs(4034) <= not(layer3_outputs(2579));
    layer4_outputs(4035) <= not((layer3_outputs(2952)) xor (layer3_outputs(4837)));
    layer4_outputs(4036) <= '1';
    layer4_outputs(4037) <= not(layer3_outputs(3478)) or (layer3_outputs(1069));
    layer4_outputs(4038) <= layer3_outputs(1075);
    layer4_outputs(4039) <= (layer3_outputs(2859)) and not (layer3_outputs(1259));
    layer4_outputs(4040) <= (layer3_outputs(5098)) or (layer3_outputs(5088));
    layer4_outputs(4041) <= not((layer3_outputs(2601)) and (layer3_outputs(4232)));
    layer4_outputs(4042) <= not(layer3_outputs(1578));
    layer4_outputs(4043) <= '1';
    layer4_outputs(4044) <= not(layer3_outputs(18)) or (layer3_outputs(1809));
    layer4_outputs(4045) <= not(layer3_outputs(853));
    layer4_outputs(4046) <= not(layer3_outputs(1664));
    layer4_outputs(4047) <= (layer3_outputs(6)) and not (layer3_outputs(913));
    layer4_outputs(4048) <= not(layer3_outputs(984)) or (layer3_outputs(3580));
    layer4_outputs(4049) <= not((layer3_outputs(4795)) or (layer3_outputs(536)));
    layer4_outputs(4050) <= (layer3_outputs(1784)) and (layer3_outputs(1144));
    layer4_outputs(4051) <= (layer3_outputs(1221)) and not (layer3_outputs(3737));
    layer4_outputs(4052) <= not((layer3_outputs(5067)) and (layer3_outputs(2338)));
    layer4_outputs(4053) <= layer3_outputs(2926);
    layer4_outputs(4054) <= layer3_outputs(1184);
    layer4_outputs(4055) <= not(layer3_outputs(1199)) or (layer3_outputs(4721));
    layer4_outputs(4056) <= not(layer3_outputs(4252)) or (layer3_outputs(295));
    layer4_outputs(4057) <= (layer3_outputs(22)) and (layer3_outputs(368));
    layer4_outputs(4058) <= (layer3_outputs(593)) and not (layer3_outputs(1403));
    layer4_outputs(4059) <= not((layer3_outputs(2556)) xor (layer3_outputs(104)));
    layer4_outputs(4060) <= not(layer3_outputs(3802)) or (layer3_outputs(2802));
    layer4_outputs(4061) <= layer3_outputs(1028);
    layer4_outputs(4062) <= layer3_outputs(1706);
    layer4_outputs(4063) <= '0';
    layer4_outputs(4064) <= not((layer3_outputs(4301)) and (layer3_outputs(4666)));
    layer4_outputs(4065) <= not(layer3_outputs(1375)) or (layer3_outputs(3352));
    layer4_outputs(4066) <= not(layer3_outputs(4317));
    layer4_outputs(4067) <= (layer3_outputs(4245)) or (layer3_outputs(4477));
    layer4_outputs(4068) <= '0';
    layer4_outputs(4069) <= (layer3_outputs(2571)) and not (layer3_outputs(2359));
    layer4_outputs(4070) <= layer3_outputs(3597);
    layer4_outputs(4071) <= (layer3_outputs(4461)) and not (layer3_outputs(5044));
    layer4_outputs(4072) <= (layer3_outputs(1603)) and not (layer3_outputs(4315));
    layer4_outputs(4073) <= (layer3_outputs(3040)) and not (layer3_outputs(4668));
    layer4_outputs(4074) <= layer3_outputs(194);
    layer4_outputs(4075) <= (layer3_outputs(3383)) and not (layer3_outputs(3143));
    layer4_outputs(4076) <= (layer3_outputs(4719)) and (layer3_outputs(4318));
    layer4_outputs(4077) <= not((layer3_outputs(4832)) or (layer3_outputs(5113)));
    layer4_outputs(4078) <= '0';
    layer4_outputs(4079) <= '1';
    layer4_outputs(4080) <= '0';
    layer4_outputs(4081) <= not(layer3_outputs(4080));
    layer4_outputs(4082) <= not(layer3_outputs(4445)) or (layer3_outputs(2436));
    layer4_outputs(4083) <= '1';
    layer4_outputs(4084) <= not(layer3_outputs(3524));
    layer4_outputs(4085) <= (layer3_outputs(2884)) and not (layer3_outputs(2591));
    layer4_outputs(4086) <= '1';
    layer4_outputs(4087) <= not(layer3_outputs(4853));
    layer4_outputs(4088) <= layer3_outputs(3240);
    layer4_outputs(4089) <= not(layer3_outputs(1303)) or (layer3_outputs(3101));
    layer4_outputs(4090) <= layer3_outputs(4322);
    layer4_outputs(4091) <= not(layer3_outputs(3931)) or (layer3_outputs(942));
    layer4_outputs(4092) <= layer3_outputs(4537);
    layer4_outputs(4093) <= not(layer3_outputs(2365)) or (layer3_outputs(805));
    layer4_outputs(4094) <= not(layer3_outputs(2263));
    layer4_outputs(4095) <= not(layer3_outputs(1397));
    layer4_outputs(4096) <= (layer3_outputs(3053)) and (layer3_outputs(1346));
    layer4_outputs(4097) <= (layer3_outputs(1842)) and (layer3_outputs(2201));
    layer4_outputs(4098) <= layer3_outputs(4040);
    layer4_outputs(4099) <= not(layer3_outputs(3208)) or (layer3_outputs(2472));
    layer4_outputs(4100) <= not((layer3_outputs(784)) or (layer3_outputs(5056)));
    layer4_outputs(4101) <= layer3_outputs(714);
    layer4_outputs(4102) <= not(layer3_outputs(1686));
    layer4_outputs(4103) <= (layer3_outputs(1156)) and (layer3_outputs(3173));
    layer4_outputs(4104) <= not(layer3_outputs(930));
    layer4_outputs(4105) <= not(layer3_outputs(4283)) or (layer3_outputs(336));
    layer4_outputs(4106) <= not((layer3_outputs(2294)) xor (layer3_outputs(633)));
    layer4_outputs(4107) <= layer3_outputs(3274);
    layer4_outputs(4108) <= (layer3_outputs(4782)) and (layer3_outputs(476));
    layer4_outputs(4109) <= layer3_outputs(757);
    layer4_outputs(4110) <= (layer3_outputs(1336)) and not (layer3_outputs(288));
    layer4_outputs(4111) <= (layer3_outputs(2794)) or (layer3_outputs(2962));
    layer4_outputs(4112) <= (layer3_outputs(4722)) or (layer3_outputs(4279));
    layer4_outputs(4113) <= not((layer3_outputs(589)) and (layer3_outputs(1553)));
    layer4_outputs(4114) <= '0';
    layer4_outputs(4115) <= (layer3_outputs(1592)) or (layer3_outputs(171));
    layer4_outputs(4116) <= not((layer3_outputs(2012)) and (layer3_outputs(2397)));
    layer4_outputs(4117) <= not(layer3_outputs(369)) or (layer3_outputs(2298));
    layer4_outputs(4118) <= not((layer3_outputs(4905)) xor (layer3_outputs(880)));
    layer4_outputs(4119) <= '1';
    layer4_outputs(4120) <= not(layer3_outputs(2905));
    layer4_outputs(4121) <= layer3_outputs(4625);
    layer4_outputs(4122) <= (layer3_outputs(4703)) and not (layer3_outputs(2270));
    layer4_outputs(4123) <= (layer3_outputs(4649)) and (layer3_outputs(429));
    layer4_outputs(4124) <= not(layer3_outputs(3399));
    layer4_outputs(4125) <= '1';
    layer4_outputs(4126) <= (layer3_outputs(3519)) and (layer3_outputs(614));
    layer4_outputs(4127) <= (layer3_outputs(1643)) and not (layer3_outputs(4696));
    layer4_outputs(4128) <= (layer3_outputs(4149)) and not (layer3_outputs(201));
    layer4_outputs(4129) <= (layer3_outputs(1773)) and not (layer3_outputs(3134));
    layer4_outputs(4130) <= (layer3_outputs(685)) and (layer3_outputs(4595));
    layer4_outputs(4131) <= '0';
    layer4_outputs(4132) <= (layer3_outputs(4175)) and not (layer3_outputs(684));
    layer4_outputs(4133) <= not(layer3_outputs(2317));
    layer4_outputs(4134) <= not((layer3_outputs(2401)) xor (layer3_outputs(3295)));
    layer4_outputs(4135) <= not(layer3_outputs(373));
    layer4_outputs(4136) <= not(layer3_outputs(2994));
    layer4_outputs(4137) <= not(layer3_outputs(2655)) or (layer3_outputs(3168));
    layer4_outputs(4138) <= not((layer3_outputs(123)) xor (layer3_outputs(4250)));
    layer4_outputs(4139) <= (layer3_outputs(5079)) and not (layer3_outputs(2360));
    layer4_outputs(4140) <= (layer3_outputs(2254)) and not (layer3_outputs(3772));
    layer4_outputs(4141) <= not(layer3_outputs(3607));
    layer4_outputs(4142) <= '1';
    layer4_outputs(4143) <= not((layer3_outputs(2485)) and (layer3_outputs(4022)));
    layer4_outputs(4144) <= layer3_outputs(67);
    layer4_outputs(4145) <= (layer3_outputs(1672)) and (layer3_outputs(1289));
    layer4_outputs(4146) <= '1';
    layer4_outputs(4147) <= (layer3_outputs(3919)) and not (layer3_outputs(2912));
    layer4_outputs(4148) <= layer3_outputs(2097);
    layer4_outputs(4149) <= not(layer3_outputs(3592));
    layer4_outputs(4150) <= (layer3_outputs(292)) xor (layer3_outputs(399));
    layer4_outputs(4151) <= (layer3_outputs(3817)) and not (layer3_outputs(4089));
    layer4_outputs(4152) <= '1';
    layer4_outputs(4153) <= layer3_outputs(1254);
    layer4_outputs(4154) <= not((layer3_outputs(3398)) xor (layer3_outputs(3404)));
    layer4_outputs(4155) <= not(layer3_outputs(214)) or (layer3_outputs(4548));
    layer4_outputs(4156) <= '0';
    layer4_outputs(4157) <= layer3_outputs(1758);
    layer4_outputs(4158) <= not(layer3_outputs(2541)) or (layer3_outputs(2485));
    layer4_outputs(4159) <= (layer3_outputs(18)) and not (layer3_outputs(4875));
    layer4_outputs(4160) <= layer3_outputs(2773);
    layer4_outputs(4161) <= layer3_outputs(4815);
    layer4_outputs(4162) <= not((layer3_outputs(4259)) or (layer3_outputs(3926)));
    layer4_outputs(4163) <= not((layer3_outputs(2663)) and (layer3_outputs(1133)));
    layer4_outputs(4164) <= not((layer3_outputs(4954)) and (layer3_outputs(3421)));
    layer4_outputs(4165) <= '0';
    layer4_outputs(4166) <= '1';
    layer4_outputs(4167) <= (layer3_outputs(2769)) and (layer3_outputs(1669));
    layer4_outputs(4168) <= '0';
    layer4_outputs(4169) <= (layer3_outputs(1539)) and not (layer3_outputs(2640));
    layer4_outputs(4170) <= not((layer3_outputs(463)) or (layer3_outputs(834)));
    layer4_outputs(4171) <= not(layer3_outputs(1322));
    layer4_outputs(4172) <= (layer3_outputs(3960)) and not (layer3_outputs(3190));
    layer4_outputs(4173) <= layer3_outputs(93);
    layer4_outputs(4174) <= not(layer3_outputs(617));
    layer4_outputs(4175) <= (layer3_outputs(1726)) and not (layer3_outputs(2505));
    layer4_outputs(4176) <= '0';
    layer4_outputs(4177) <= not(layer3_outputs(75));
    layer4_outputs(4178) <= (layer3_outputs(2662)) or (layer3_outputs(4510));
    layer4_outputs(4179) <= (layer3_outputs(1717)) or (layer3_outputs(3573));
    layer4_outputs(4180) <= not(layer3_outputs(2858));
    layer4_outputs(4181) <= not(layer3_outputs(113)) or (layer3_outputs(2665));
    layer4_outputs(4182) <= not(layer3_outputs(1999));
    layer4_outputs(4183) <= not(layer3_outputs(3567));
    layer4_outputs(4184) <= '0';
    layer4_outputs(4185) <= not((layer3_outputs(3071)) and (layer3_outputs(1775)));
    layer4_outputs(4186) <= layer3_outputs(681);
    layer4_outputs(4187) <= '1';
    layer4_outputs(4188) <= not(layer3_outputs(3893)) or (layer3_outputs(2708));
    layer4_outputs(4189) <= (layer3_outputs(2552)) and (layer3_outputs(2961));
    layer4_outputs(4190) <= not((layer3_outputs(1723)) and (layer3_outputs(2504)));
    layer4_outputs(4191) <= layer3_outputs(1018);
    layer4_outputs(4192) <= layer3_outputs(1596);
    layer4_outputs(4193) <= (layer3_outputs(423)) xor (layer3_outputs(2466));
    layer4_outputs(4194) <= (layer3_outputs(1233)) and not (layer3_outputs(4163));
    layer4_outputs(4195) <= (layer3_outputs(237)) or (layer3_outputs(4888));
    layer4_outputs(4196) <= not((layer3_outputs(1859)) and (layer3_outputs(623)));
    layer4_outputs(4197) <= '0';
    layer4_outputs(4198) <= not(layer3_outputs(3111));
    layer4_outputs(4199) <= (layer3_outputs(2828)) and not (layer3_outputs(3409));
    layer4_outputs(4200) <= layer3_outputs(4262);
    layer4_outputs(4201) <= not(layer3_outputs(68)) or (layer3_outputs(623));
    layer4_outputs(4202) <= '1';
    layer4_outputs(4203) <= (layer3_outputs(2440)) and not (layer3_outputs(656));
    layer4_outputs(4204) <= not(layer3_outputs(1665)) or (layer3_outputs(847));
    layer4_outputs(4205) <= (layer3_outputs(848)) or (layer3_outputs(1183));
    layer4_outputs(4206) <= '1';
    layer4_outputs(4207) <= layer3_outputs(1291);
    layer4_outputs(4208) <= layer3_outputs(410);
    layer4_outputs(4209) <= (layer3_outputs(2754)) and not (layer3_outputs(3845));
    layer4_outputs(4210) <= '1';
    layer4_outputs(4211) <= not(layer3_outputs(1642));
    layer4_outputs(4212) <= '1';
    layer4_outputs(4213) <= layer3_outputs(4886);
    layer4_outputs(4214) <= '0';
    layer4_outputs(4215) <= not((layer3_outputs(161)) or (layer3_outputs(4064)));
    layer4_outputs(4216) <= (layer3_outputs(1622)) or (layer3_outputs(334));
    layer4_outputs(4217) <= not(layer3_outputs(1517));
    layer4_outputs(4218) <= (layer3_outputs(759)) or (layer3_outputs(1302));
    layer4_outputs(4219) <= '0';
    layer4_outputs(4220) <= not((layer3_outputs(3610)) or (layer3_outputs(2539)));
    layer4_outputs(4221) <= layer3_outputs(3676);
    layer4_outputs(4222) <= not(layer3_outputs(894)) or (layer3_outputs(2415));
    layer4_outputs(4223) <= (layer3_outputs(1683)) and not (layer3_outputs(5078));
    layer4_outputs(4224) <= not(layer3_outputs(1370)) or (layer3_outputs(4195));
    layer4_outputs(4225) <= '1';
    layer4_outputs(4226) <= not((layer3_outputs(4705)) and (layer3_outputs(940)));
    layer4_outputs(4227) <= (layer3_outputs(2680)) or (layer3_outputs(332));
    layer4_outputs(4228) <= layer3_outputs(4540);
    layer4_outputs(4229) <= (layer3_outputs(4437)) and not (layer3_outputs(3694));
    layer4_outputs(4230) <= '1';
    layer4_outputs(4231) <= (layer3_outputs(854)) and not (layer3_outputs(4776));
    layer4_outputs(4232) <= not(layer3_outputs(1755)) or (layer3_outputs(2272));
    layer4_outputs(4233) <= not(layer3_outputs(2198)) or (layer3_outputs(649));
    layer4_outputs(4234) <= (layer3_outputs(928)) and not (layer3_outputs(1369));
    layer4_outputs(4235) <= not((layer3_outputs(3517)) and (layer3_outputs(562)));
    layer4_outputs(4236) <= (layer3_outputs(3105)) xor (layer3_outputs(3218));
    layer4_outputs(4237) <= (layer3_outputs(1401)) and (layer3_outputs(2380));
    layer4_outputs(4238) <= not((layer3_outputs(101)) and (layer3_outputs(572)));
    layer4_outputs(4239) <= not((layer3_outputs(1845)) or (layer3_outputs(3920)));
    layer4_outputs(4240) <= layer3_outputs(194);
    layer4_outputs(4241) <= not(layer3_outputs(1426));
    layer4_outputs(4242) <= not(layer3_outputs(2365)) or (layer3_outputs(3238));
    layer4_outputs(4243) <= not(layer3_outputs(585));
    layer4_outputs(4244) <= (layer3_outputs(1508)) and not (layer3_outputs(1402));
    layer4_outputs(4245) <= not(layer3_outputs(5090)) or (layer3_outputs(420));
    layer4_outputs(4246) <= not((layer3_outputs(391)) or (layer3_outputs(5117)));
    layer4_outputs(4247) <= not(layer3_outputs(2215)) or (layer3_outputs(1854));
    layer4_outputs(4248) <= layer3_outputs(1520);
    layer4_outputs(4249) <= layer3_outputs(4626);
    layer4_outputs(4250) <= (layer3_outputs(1016)) and (layer3_outputs(1944));
    layer4_outputs(4251) <= '1';
    layer4_outputs(4252) <= not((layer3_outputs(3339)) and (layer3_outputs(4553)));
    layer4_outputs(4253) <= (layer3_outputs(2927)) and (layer3_outputs(1473));
    layer4_outputs(4254) <= (layer3_outputs(35)) and not (layer3_outputs(2058));
    layer4_outputs(4255) <= not(layer3_outputs(3959)) or (layer3_outputs(33));
    layer4_outputs(4256) <= not(layer3_outputs(2702));
    layer4_outputs(4257) <= (layer3_outputs(1530)) and not (layer3_outputs(4975));
    layer4_outputs(4258) <= layer3_outputs(3285);
    layer4_outputs(4259) <= (layer3_outputs(2786)) or (layer3_outputs(3986));
    layer4_outputs(4260) <= (layer3_outputs(4153)) or (layer3_outputs(1721));
    layer4_outputs(4261) <= '1';
    layer4_outputs(4262) <= '1';
    layer4_outputs(4263) <= layer3_outputs(2506);
    layer4_outputs(4264) <= layer3_outputs(1840);
    layer4_outputs(4265) <= '0';
    layer4_outputs(4266) <= not((layer3_outputs(3703)) and (layer3_outputs(1575)));
    layer4_outputs(4267) <= not(layer3_outputs(2138)) or (layer3_outputs(500));
    layer4_outputs(4268) <= not(layer3_outputs(2643)) or (layer3_outputs(435));
    layer4_outputs(4269) <= not(layer3_outputs(3752)) or (layer3_outputs(3876));
    layer4_outputs(4270) <= (layer3_outputs(1360)) and not (layer3_outputs(331));
    layer4_outputs(4271) <= not(layer3_outputs(4124)) or (layer3_outputs(3154));
    layer4_outputs(4272) <= '1';
    layer4_outputs(4273) <= (layer3_outputs(67)) xor (layer3_outputs(2092));
    layer4_outputs(4274) <= layer3_outputs(1066);
    layer4_outputs(4275) <= not((layer3_outputs(2547)) or (layer3_outputs(1598)));
    layer4_outputs(4276) <= not(layer3_outputs(321));
    layer4_outputs(4277) <= layer3_outputs(2439);
    layer4_outputs(4278) <= layer3_outputs(789);
    layer4_outputs(4279) <= '1';
    layer4_outputs(4280) <= not(layer3_outputs(3572));
    layer4_outputs(4281) <= (layer3_outputs(210)) and not (layer3_outputs(1470));
    layer4_outputs(4282) <= layer3_outputs(1247);
    layer4_outputs(4283) <= not(layer3_outputs(4028));
    layer4_outputs(4284) <= '0';
    layer4_outputs(4285) <= (layer3_outputs(229)) or (layer3_outputs(333));
    layer4_outputs(4286) <= '0';
    layer4_outputs(4287) <= (layer3_outputs(3943)) and not (layer3_outputs(612));
    layer4_outputs(4288) <= (layer3_outputs(857)) and not (layer3_outputs(1488));
    layer4_outputs(4289) <= not((layer3_outputs(5114)) xor (layer3_outputs(57)));
    layer4_outputs(4290) <= not((layer3_outputs(414)) or (layer3_outputs(2590)));
    layer4_outputs(4291) <= not((layer3_outputs(785)) and (layer3_outputs(2043)));
    layer4_outputs(4292) <= (layer3_outputs(1947)) and not (layer3_outputs(3482));
    layer4_outputs(4293) <= not(layer3_outputs(2633));
    layer4_outputs(4294) <= not((layer3_outputs(3213)) or (layer3_outputs(1073)));
    layer4_outputs(4295) <= (layer3_outputs(1477)) and (layer3_outputs(1702));
    layer4_outputs(4296) <= (layer3_outputs(4447)) or (layer3_outputs(4157));
    layer4_outputs(4297) <= (layer3_outputs(4033)) and not (layer3_outputs(1337));
    layer4_outputs(4298) <= layer3_outputs(2119);
    layer4_outputs(4299) <= not((layer3_outputs(5071)) or (layer3_outputs(4766)));
    layer4_outputs(4300) <= not(layer3_outputs(599));
    layer4_outputs(4301) <= layer3_outputs(4693);
    layer4_outputs(4302) <= layer3_outputs(286);
    layer4_outputs(4303) <= not(layer3_outputs(4210));
    layer4_outputs(4304) <= not(layer3_outputs(948)) or (layer3_outputs(687));
    layer4_outputs(4305) <= (layer3_outputs(235)) and not (layer3_outputs(1403));
    layer4_outputs(4306) <= not((layer3_outputs(2809)) and (layer3_outputs(4378)));
    layer4_outputs(4307) <= (layer3_outputs(659)) and (layer3_outputs(671));
    layer4_outputs(4308) <= not(layer3_outputs(151));
    layer4_outputs(4309) <= not(layer3_outputs(2571)) or (layer3_outputs(3427));
    layer4_outputs(4310) <= not(layer3_outputs(1314)) or (layer3_outputs(257));
    layer4_outputs(4311) <= not((layer3_outputs(770)) or (layer3_outputs(3981)));
    layer4_outputs(4312) <= not((layer3_outputs(2206)) and (layer3_outputs(562)));
    layer4_outputs(4313) <= '1';
    layer4_outputs(4314) <= not(layer3_outputs(1395)) or (layer3_outputs(873));
    layer4_outputs(4315) <= not(layer3_outputs(4519));
    layer4_outputs(4316) <= (layer3_outputs(3196)) and not (layer3_outputs(2983));
    layer4_outputs(4317) <= layer3_outputs(4017);
    layer4_outputs(4318) <= '1';
    layer4_outputs(4319) <= layer3_outputs(4884);
    layer4_outputs(4320) <= (layer3_outputs(2381)) and not (layer3_outputs(1027));
    layer4_outputs(4321) <= '1';
    layer4_outputs(4322) <= not((layer3_outputs(2544)) or (layer3_outputs(429)));
    layer4_outputs(4323) <= (layer3_outputs(1703)) and not (layer3_outputs(4952));
    layer4_outputs(4324) <= not(layer3_outputs(2419)) or (layer3_outputs(5057));
    layer4_outputs(4325) <= not((layer3_outputs(1866)) and (layer3_outputs(1827)));
    layer4_outputs(4326) <= not(layer3_outputs(1777));
    layer4_outputs(4327) <= layer3_outputs(4052);
    layer4_outputs(4328) <= '0';
    layer4_outputs(4329) <= not(layer3_outputs(3055)) or (layer3_outputs(1057));
    layer4_outputs(4330) <= '1';
    layer4_outputs(4331) <= layer3_outputs(2743);
    layer4_outputs(4332) <= (layer3_outputs(1020)) and not (layer3_outputs(3887));
    layer4_outputs(4333) <= not((layer3_outputs(3471)) or (layer3_outputs(4294)));
    layer4_outputs(4334) <= not(layer3_outputs(2633));
    layer4_outputs(4335) <= layer3_outputs(4014);
    layer4_outputs(4336) <= not(layer3_outputs(4776));
    layer4_outputs(4337) <= (layer3_outputs(427)) and (layer3_outputs(3816));
    layer4_outputs(4338) <= layer3_outputs(3693);
    layer4_outputs(4339) <= not((layer3_outputs(3420)) or (layer3_outputs(499)));
    layer4_outputs(4340) <= not(layer3_outputs(3841)) or (layer3_outputs(4024));
    layer4_outputs(4341) <= (layer3_outputs(103)) or (layer3_outputs(4172));
    layer4_outputs(4342) <= layer3_outputs(2354);
    layer4_outputs(4343) <= not(layer3_outputs(3689)) or (layer3_outputs(298));
    layer4_outputs(4344) <= not(layer3_outputs(153)) or (layer3_outputs(659));
    layer4_outputs(4345) <= not(layer3_outputs(2893)) or (layer3_outputs(1458));
    layer4_outputs(4346) <= (layer3_outputs(4648)) or (layer3_outputs(4741));
    layer4_outputs(4347) <= not((layer3_outputs(843)) or (layer3_outputs(885)));
    layer4_outputs(4348) <= layer3_outputs(1082);
    layer4_outputs(4349) <= not(layer3_outputs(1330)) or (layer3_outputs(1141));
    layer4_outputs(4350) <= not(layer3_outputs(3294));
    layer4_outputs(4351) <= not(layer3_outputs(483));
    layer4_outputs(4352) <= not(layer3_outputs(4576));
    layer4_outputs(4353) <= not((layer3_outputs(4984)) and (layer3_outputs(2492)));
    layer4_outputs(4354) <= not((layer3_outputs(5032)) and (layer3_outputs(4836)));
    layer4_outputs(4355) <= not((layer3_outputs(3258)) xor (layer3_outputs(3757)));
    layer4_outputs(4356) <= layer3_outputs(2024);
    layer4_outputs(4357) <= not((layer3_outputs(3813)) or (layer3_outputs(4979)));
    layer4_outputs(4358) <= layer3_outputs(4414);
    layer4_outputs(4359) <= layer3_outputs(2728);
    layer4_outputs(4360) <= '1';
    layer4_outputs(4361) <= not(layer3_outputs(2837)) or (layer3_outputs(1253));
    layer4_outputs(4362) <= layer3_outputs(2322);
    layer4_outputs(4363) <= (layer3_outputs(2311)) and not (layer3_outputs(1130));
    layer4_outputs(4364) <= not(layer3_outputs(4336));
    layer4_outputs(4365) <= not(layer3_outputs(1383)) or (layer3_outputs(2864));
    layer4_outputs(4366) <= not(layer3_outputs(1905)) or (layer3_outputs(694));
    layer4_outputs(4367) <= (layer3_outputs(2717)) and not (layer3_outputs(1052));
    layer4_outputs(4368) <= layer3_outputs(4014);
    layer4_outputs(4369) <= (layer3_outputs(2659)) and not (layer3_outputs(4394));
    layer4_outputs(4370) <= not(layer3_outputs(2444));
    layer4_outputs(4371) <= layer3_outputs(41);
    layer4_outputs(4372) <= '0';
    layer4_outputs(4373) <= '1';
    layer4_outputs(4374) <= layer3_outputs(3082);
    layer4_outputs(4375) <= not((layer3_outputs(4022)) xor (layer3_outputs(186)));
    layer4_outputs(4376) <= layer3_outputs(837);
    layer4_outputs(4377) <= not(layer3_outputs(3384)) or (layer3_outputs(1609));
    layer4_outputs(4378) <= (layer3_outputs(2876)) and not (layer3_outputs(2494));
    layer4_outputs(4379) <= not(layer3_outputs(482)) or (layer3_outputs(628));
    layer4_outputs(4380) <= (layer3_outputs(1849)) and not (layer3_outputs(584));
    layer4_outputs(4381) <= layer3_outputs(971);
    layer4_outputs(4382) <= not((layer3_outputs(3651)) and (layer3_outputs(1089)));
    layer4_outputs(4383) <= (layer3_outputs(4556)) and (layer3_outputs(4607));
    layer4_outputs(4384) <= not((layer3_outputs(1249)) and (layer3_outputs(3127)));
    layer4_outputs(4385) <= '1';
    layer4_outputs(4386) <= (layer3_outputs(4973)) and not (layer3_outputs(3028));
    layer4_outputs(4387) <= (layer3_outputs(4432)) and not (layer3_outputs(2708));
    layer4_outputs(4388) <= '1';
    layer4_outputs(4389) <= '0';
    layer4_outputs(4390) <= (layer3_outputs(1621)) and (layer3_outputs(4238));
    layer4_outputs(4391) <= '0';
    layer4_outputs(4392) <= (layer3_outputs(503)) and not (layer3_outputs(2827));
    layer4_outputs(4393) <= not(layer3_outputs(2587));
    layer4_outputs(4394) <= (layer3_outputs(192)) or (layer3_outputs(4920));
    layer4_outputs(4395) <= not((layer3_outputs(4908)) and (layer3_outputs(1783)));
    layer4_outputs(4396) <= '1';
    layer4_outputs(4397) <= not((layer3_outputs(707)) or (layer3_outputs(3677)));
    layer4_outputs(4398) <= not((layer3_outputs(2882)) and (layer3_outputs(1853)));
    layer4_outputs(4399) <= layer3_outputs(2059);
    layer4_outputs(4400) <= '0';
    layer4_outputs(4401) <= (layer3_outputs(3816)) or (layer3_outputs(4073));
    layer4_outputs(4402) <= not((layer3_outputs(3995)) and (layer3_outputs(2977)));
    layer4_outputs(4403) <= layer3_outputs(3861);
    layer4_outputs(4404) <= (layer3_outputs(2457)) or (layer3_outputs(711));
    layer4_outputs(4405) <= layer3_outputs(241);
    layer4_outputs(4406) <= (layer3_outputs(229)) or (layer3_outputs(4678));
    layer4_outputs(4407) <= (layer3_outputs(1770)) and not (layer3_outputs(4346));
    layer4_outputs(4408) <= (layer3_outputs(4268)) and not (layer3_outputs(1421));
    layer4_outputs(4409) <= not(layer3_outputs(280)) or (layer3_outputs(3934));
    layer4_outputs(4410) <= not((layer3_outputs(4642)) and (layer3_outputs(285)));
    layer4_outputs(4411) <= (layer3_outputs(4881)) or (layer3_outputs(1665));
    layer4_outputs(4412) <= (layer3_outputs(2789)) and not (layer3_outputs(4673));
    layer4_outputs(4413) <= not(layer3_outputs(1994)) or (layer3_outputs(3524));
    layer4_outputs(4414) <= not(layer3_outputs(3555));
    layer4_outputs(4415) <= layer3_outputs(4727);
    layer4_outputs(4416) <= (layer3_outputs(1058)) and not (layer3_outputs(3847));
    layer4_outputs(4417) <= '0';
    layer4_outputs(4418) <= not(layer3_outputs(864));
    layer4_outputs(4419) <= layer3_outputs(688);
    layer4_outputs(4420) <= (layer3_outputs(1807)) and (layer3_outputs(3180));
    layer4_outputs(4421) <= not(layer3_outputs(1339)) or (layer3_outputs(3944));
    layer4_outputs(4422) <= (layer3_outputs(4583)) xor (layer3_outputs(1191));
    layer4_outputs(4423) <= not((layer3_outputs(1376)) and (layer3_outputs(4165)));
    layer4_outputs(4424) <= (layer3_outputs(2844)) and not (layer3_outputs(749));
    layer4_outputs(4425) <= not(layer3_outputs(1540)) or (layer3_outputs(1558));
    layer4_outputs(4426) <= not((layer3_outputs(4890)) or (layer3_outputs(2898)));
    layer4_outputs(4427) <= layer3_outputs(4107);
    layer4_outputs(4428) <= not(layer3_outputs(4443)) or (layer3_outputs(1623));
    layer4_outputs(4429) <= '1';
    layer4_outputs(4430) <= (layer3_outputs(4187)) and (layer3_outputs(4382));
    layer4_outputs(4431) <= not(layer3_outputs(2368)) or (layer3_outputs(4956));
    layer4_outputs(4432) <= (layer3_outputs(3646)) or (layer3_outputs(839));
    layer4_outputs(4433) <= '0';
    layer4_outputs(4434) <= not((layer3_outputs(939)) and (layer3_outputs(4293)));
    layer4_outputs(4435) <= layer3_outputs(3905);
    layer4_outputs(4436) <= (layer3_outputs(2712)) and (layer3_outputs(2020));
    layer4_outputs(4437) <= not(layer3_outputs(12));
    layer4_outputs(4438) <= not((layer3_outputs(964)) and (layer3_outputs(2911)));
    layer4_outputs(4439) <= not((layer3_outputs(3958)) and (layer3_outputs(2871)));
    layer4_outputs(4440) <= not((layer3_outputs(4170)) or (layer3_outputs(481)));
    layer4_outputs(4441) <= not(layer3_outputs(2300));
    layer4_outputs(4442) <= not(layer3_outputs(1062));
    layer4_outputs(4443) <= (layer3_outputs(3635)) and (layer3_outputs(1394));
    layer4_outputs(4444) <= not(layer3_outputs(867));
    layer4_outputs(4445) <= (layer3_outputs(166)) and not (layer3_outputs(1648));
    layer4_outputs(4446) <= not(layer3_outputs(287));
    layer4_outputs(4447) <= not(layer3_outputs(4838));
    layer4_outputs(4448) <= not(layer3_outputs(2108));
    layer4_outputs(4449) <= not(layer3_outputs(3502));
    layer4_outputs(4450) <= '1';
    layer4_outputs(4451) <= not((layer3_outputs(4676)) or (layer3_outputs(474)));
    layer4_outputs(4452) <= (layer3_outputs(1627)) and not (layer3_outputs(828));
    layer4_outputs(4453) <= not((layer3_outputs(3800)) or (layer3_outputs(2149)));
    layer4_outputs(4454) <= layer3_outputs(4260);
    layer4_outputs(4455) <= (layer3_outputs(3740)) and not (layer3_outputs(430));
    layer4_outputs(4456) <= layer3_outputs(4939);
    layer4_outputs(4457) <= (layer3_outputs(19)) or (layer3_outputs(2726));
    layer4_outputs(4458) <= not(layer3_outputs(1881));
    layer4_outputs(4459) <= not(layer3_outputs(125)) or (layer3_outputs(1027));
    layer4_outputs(4460) <= '1';
    layer4_outputs(4461) <= not((layer3_outputs(65)) xor (layer3_outputs(1277)));
    layer4_outputs(4462) <= not(layer3_outputs(1602)) or (layer3_outputs(4222));
    layer4_outputs(4463) <= (layer3_outputs(767)) and not (layer3_outputs(503));
    layer4_outputs(4464) <= layer3_outputs(4624);
    layer4_outputs(4465) <= (layer3_outputs(1864)) or (layer3_outputs(4606));
    layer4_outputs(4466) <= (layer3_outputs(3643)) and (layer3_outputs(3381));
    layer4_outputs(4467) <= not(layer3_outputs(2036)) or (layer3_outputs(2979));
    layer4_outputs(4468) <= not((layer3_outputs(4930)) or (layer3_outputs(3863)));
    layer4_outputs(4469) <= (layer3_outputs(1178)) and (layer3_outputs(472));
    layer4_outputs(4470) <= not((layer3_outputs(1366)) or (layer3_outputs(1717)));
    layer4_outputs(4471) <= not(layer3_outputs(660)) or (layer3_outputs(3116));
    layer4_outputs(4472) <= not((layer3_outputs(3212)) and (layer3_outputs(140)));
    layer4_outputs(4473) <= (layer3_outputs(3485)) and not (layer3_outputs(1712));
    layer4_outputs(4474) <= (layer3_outputs(2111)) and not (layer3_outputs(3025));
    layer4_outputs(4475) <= '1';
    layer4_outputs(4476) <= layer3_outputs(2383);
    layer4_outputs(4477) <= not(layer3_outputs(1988)) or (layer3_outputs(4619));
    layer4_outputs(4478) <= not((layer3_outputs(5029)) or (layer3_outputs(4500)));
    layer4_outputs(4479) <= not(layer3_outputs(117)) or (layer3_outputs(634));
    layer4_outputs(4480) <= '1';
    layer4_outputs(4481) <= not(layer3_outputs(915));
    layer4_outputs(4482) <= layer3_outputs(3444);
    layer4_outputs(4483) <= (layer3_outputs(3171)) and (layer3_outputs(2732));
    layer4_outputs(4484) <= not(layer3_outputs(3730)) or (layer3_outputs(2834));
    layer4_outputs(4485) <= (layer3_outputs(3571)) and (layer3_outputs(1276));
    layer4_outputs(4486) <= (layer3_outputs(2496)) and not (layer3_outputs(1380));
    layer4_outputs(4487) <= not((layer3_outputs(2259)) and (layer3_outputs(450)));
    layer4_outputs(4488) <= '1';
    layer4_outputs(4489) <= not((layer3_outputs(756)) or (layer3_outputs(1765)));
    layer4_outputs(4490) <= (layer3_outputs(4586)) and (layer3_outputs(603));
    layer4_outputs(4491) <= not(layer3_outputs(2175)) or (layer3_outputs(2374));
    layer4_outputs(4492) <= '1';
    layer4_outputs(4493) <= '1';
    layer4_outputs(4494) <= layer3_outputs(3975);
    layer4_outputs(4495) <= (layer3_outputs(1976)) and not (layer3_outputs(3549));
    layer4_outputs(4496) <= (layer3_outputs(1616)) and not (layer3_outputs(4341));
    layer4_outputs(4497) <= not((layer3_outputs(3329)) or (layer3_outputs(4554)));
    layer4_outputs(4498) <= layer3_outputs(4198);
    layer4_outputs(4499) <= layer3_outputs(2431);
    layer4_outputs(4500) <= not(layer3_outputs(3641));
    layer4_outputs(4501) <= not(layer3_outputs(1354)) or (layer3_outputs(4717));
    layer4_outputs(4502) <= not(layer3_outputs(3426));
    layer4_outputs(4503) <= (layer3_outputs(2039)) and not (layer3_outputs(142));
    layer4_outputs(4504) <= '0';
    layer4_outputs(4505) <= '0';
    layer4_outputs(4506) <= '0';
    layer4_outputs(4507) <= '1';
    layer4_outputs(4508) <= layer3_outputs(3076);
    layer4_outputs(4509) <= not((layer3_outputs(4927)) and (layer3_outputs(1306)));
    layer4_outputs(4510) <= layer3_outputs(791);
    layer4_outputs(4511) <= not(layer3_outputs(1639));
    layer4_outputs(4512) <= (layer3_outputs(2457)) or (layer3_outputs(3433));
    layer4_outputs(4513) <= not(layer3_outputs(1162));
    layer4_outputs(4514) <= layer3_outputs(4218);
    layer4_outputs(4515) <= (layer3_outputs(2084)) and not (layer3_outputs(1743));
    layer4_outputs(4516) <= '0';
    layer4_outputs(4517) <= not(layer3_outputs(4858));
    layer4_outputs(4518) <= (layer3_outputs(3006)) and not (layer3_outputs(2477));
    layer4_outputs(4519) <= not(layer3_outputs(1007)) or (layer3_outputs(78));
    layer4_outputs(4520) <= (layer3_outputs(5055)) and not (layer3_outputs(4686));
    layer4_outputs(4521) <= '1';
    layer4_outputs(4522) <= not(layer3_outputs(1167));
    layer4_outputs(4523) <= (layer3_outputs(2480)) or (layer3_outputs(4498));
    layer4_outputs(4524) <= '1';
    layer4_outputs(4525) <= layer3_outputs(5094);
    layer4_outputs(4526) <= (layer3_outputs(2782)) and not (layer3_outputs(4011));
    layer4_outputs(4527) <= (layer3_outputs(866)) and not (layer3_outputs(1008));
    layer4_outputs(4528) <= not(layer3_outputs(786)) or (layer3_outputs(3542));
    layer4_outputs(4529) <= (layer3_outputs(4947)) or (layer3_outputs(994));
    layer4_outputs(4530) <= not(layer3_outputs(2761));
    layer4_outputs(4531) <= not((layer3_outputs(1489)) and (layer3_outputs(4379)));
    layer4_outputs(4532) <= '1';
    layer4_outputs(4533) <= not(layer3_outputs(3253));
    layer4_outputs(4534) <= (layer3_outputs(629)) or (layer3_outputs(422));
    layer4_outputs(4535) <= not((layer3_outputs(1858)) and (layer3_outputs(1413)));
    layer4_outputs(4536) <= (layer3_outputs(2993)) and (layer3_outputs(4855));
    layer4_outputs(4537) <= layer3_outputs(4946);
    layer4_outputs(4538) <= not(layer3_outputs(3079)) or (layer3_outputs(1284));
    layer4_outputs(4539) <= not(layer3_outputs(570));
    layer4_outputs(4540) <= layer3_outputs(3322);
    layer4_outputs(4541) <= not(layer3_outputs(3414));
    layer4_outputs(4542) <= not(layer3_outputs(624));
    layer4_outputs(4543) <= '0';
    layer4_outputs(4544) <= (layer3_outputs(4070)) or (layer3_outputs(553));
    layer4_outputs(4545) <= not(layer3_outputs(2139)) or (layer3_outputs(540));
    layer4_outputs(4546) <= '0';
    layer4_outputs(4547) <= (layer3_outputs(3850)) or (layer3_outputs(4724));
    layer4_outputs(4548) <= (layer3_outputs(4145)) or (layer3_outputs(2713));
    layer4_outputs(4549) <= not(layer3_outputs(4704));
    layer4_outputs(4550) <= not((layer3_outputs(3792)) and (layer3_outputs(3097)));
    layer4_outputs(4551) <= not(layer3_outputs(1651));
    layer4_outputs(4552) <= not(layer3_outputs(3072));
    layer4_outputs(4553) <= (layer3_outputs(2371)) or (layer3_outputs(4164));
    layer4_outputs(4554) <= not(layer3_outputs(1744));
    layer4_outputs(4555) <= layer3_outputs(729);
    layer4_outputs(4556) <= not((layer3_outputs(4439)) or (layer3_outputs(4478)));
    layer4_outputs(4557) <= '0';
    layer4_outputs(4558) <= (layer3_outputs(2852)) or (layer3_outputs(3676));
    layer4_outputs(4559) <= not(layer3_outputs(1095));
    layer4_outputs(4560) <= not((layer3_outputs(3263)) and (layer3_outputs(3140)));
    layer4_outputs(4561) <= '1';
    layer4_outputs(4562) <= not((layer3_outputs(2199)) xor (layer3_outputs(1308)));
    layer4_outputs(4563) <= not((layer3_outputs(1823)) or (layer3_outputs(3377)));
    layer4_outputs(4564) <= '0';
    layer4_outputs(4565) <= (layer3_outputs(547)) or (layer3_outputs(5073));
    layer4_outputs(4566) <= not((layer3_outputs(1614)) or (layer3_outputs(2763)));
    layer4_outputs(4567) <= not(layer3_outputs(4023)) or (layer3_outputs(3290));
    layer4_outputs(4568) <= layer3_outputs(3394);
    layer4_outputs(4569) <= (layer3_outputs(824)) and not (layer3_outputs(2245));
    layer4_outputs(4570) <= not(layer3_outputs(1984)) or (layer3_outputs(4254));
    layer4_outputs(4571) <= not(layer3_outputs(445)) or (layer3_outputs(3223));
    layer4_outputs(4572) <= not(layer3_outputs(3909)) or (layer3_outputs(2495));
    layer4_outputs(4573) <= not((layer3_outputs(1123)) and (layer3_outputs(1939)));
    layer4_outputs(4574) <= (layer3_outputs(439)) and not (layer3_outputs(2146));
    layer4_outputs(4575) <= not((layer3_outputs(4948)) and (layer3_outputs(3476)));
    layer4_outputs(4576) <= '1';
    layer4_outputs(4577) <= layer3_outputs(4808);
    layer4_outputs(4578) <= (layer3_outputs(3765)) and not (layer3_outputs(4735));
    layer4_outputs(4579) <= not(layer3_outputs(3472)) or (layer3_outputs(1379));
    layer4_outputs(4580) <= layer3_outputs(2535);
    layer4_outputs(4581) <= not(layer3_outputs(2878));
    layer4_outputs(4582) <= layer3_outputs(1321);
    layer4_outputs(4583) <= not((layer3_outputs(3670)) and (layer3_outputs(2413)));
    layer4_outputs(4584) <= (layer3_outputs(3241)) and (layer3_outputs(2426));
    layer4_outputs(4585) <= not(layer3_outputs(3946)) or (layer3_outputs(3251));
    layer4_outputs(4586) <= (layer3_outputs(1978)) and (layer3_outputs(2134));
    layer4_outputs(4587) <= (layer3_outputs(282)) and not (layer3_outputs(1505));
    layer4_outputs(4588) <= not(layer3_outputs(961)) or (layer3_outputs(1248));
    layer4_outputs(4589) <= not(layer3_outputs(976));
    layer4_outputs(4590) <= '0';
    layer4_outputs(4591) <= layer3_outputs(5039);
    layer4_outputs(4592) <= not(layer3_outputs(651));
    layer4_outputs(4593) <= (layer3_outputs(2892)) or (layer3_outputs(1678));
    layer4_outputs(4594) <= '0';
    layer4_outputs(4595) <= (layer3_outputs(2685)) and not (layer3_outputs(4683));
    layer4_outputs(4596) <= not(layer3_outputs(4791)) or (layer3_outputs(3745));
    layer4_outputs(4597) <= (layer3_outputs(3890)) and not (layer3_outputs(3459));
    layer4_outputs(4598) <= (layer3_outputs(2766)) and (layer3_outputs(4512));
    layer4_outputs(4599) <= not((layer3_outputs(4007)) and (layer3_outputs(4071)));
    layer4_outputs(4600) <= layer3_outputs(258);
    layer4_outputs(4601) <= layer3_outputs(3272);
    layer4_outputs(4602) <= not((layer3_outputs(279)) or (layer3_outputs(4302)));
    layer4_outputs(4603) <= not(layer3_outputs(205));
    layer4_outputs(4604) <= '1';
    layer4_outputs(4605) <= '0';
    layer4_outputs(4606) <= not(layer3_outputs(3550)) or (layer3_outputs(1364));
    layer4_outputs(4607) <= layer3_outputs(3138);
    layer4_outputs(4608) <= not(layer3_outputs(1740)) or (layer3_outputs(3008));
    layer4_outputs(4609) <= (layer3_outputs(3786)) or (layer3_outputs(3602));
    layer4_outputs(4610) <= not(layer3_outputs(71));
    layer4_outputs(4611) <= (layer3_outputs(108)) and not (layer3_outputs(2578));
    layer4_outputs(4612) <= '1';
    layer4_outputs(4613) <= not(layer3_outputs(3082));
    layer4_outputs(4614) <= (layer3_outputs(1785)) and not (layer3_outputs(4588));
    layer4_outputs(4615) <= layer3_outputs(3115);
    layer4_outputs(4616) <= not(layer3_outputs(4183)) or (layer3_outputs(2391));
    layer4_outputs(4617) <= '0';
    layer4_outputs(4618) <= (layer3_outputs(1922)) and not (layer3_outputs(3090));
    layer4_outputs(4619) <= '0';
    layer4_outputs(4620) <= layer3_outputs(900);
    layer4_outputs(4621) <= layer3_outputs(5055);
    layer4_outputs(4622) <= (layer3_outputs(2388)) and not (layer3_outputs(1648));
    layer4_outputs(4623) <= layer3_outputs(413);
    layer4_outputs(4624) <= not(layer3_outputs(4359)) or (layer3_outputs(956));
    layer4_outputs(4625) <= '0';
    layer4_outputs(4626) <= layer3_outputs(2032);
    layer4_outputs(4627) <= (layer3_outputs(475)) or (layer3_outputs(2083));
    layer4_outputs(4628) <= layer3_outputs(243);
    layer4_outputs(4629) <= layer3_outputs(2288);
    layer4_outputs(4630) <= '0';
    layer4_outputs(4631) <= '1';
    layer4_outputs(4632) <= not((layer3_outputs(2343)) or (layer3_outputs(1382)));
    layer4_outputs(4633) <= not(layer3_outputs(4370)) or (layer3_outputs(953));
    layer4_outputs(4634) <= '1';
    layer4_outputs(4635) <= (layer3_outputs(1034)) or (layer3_outputs(4462));
    layer4_outputs(4636) <= '0';
    layer4_outputs(4637) <= (layer3_outputs(1814)) or (layer3_outputs(975));
    layer4_outputs(4638) <= (layer3_outputs(2688)) and not (layer3_outputs(1513));
    layer4_outputs(4639) <= not(layer3_outputs(2676)) or (layer3_outputs(1201));
    layer4_outputs(4640) <= layer3_outputs(447);
    layer4_outputs(4641) <= (layer3_outputs(382)) and not (layer3_outputs(4843));
    layer4_outputs(4642) <= (layer3_outputs(3145)) and (layer3_outputs(376));
    layer4_outputs(4643) <= not(layer3_outputs(3067));
    layer4_outputs(4644) <= '1';
    layer4_outputs(4645) <= not((layer3_outputs(4652)) and (layer3_outputs(2823)));
    layer4_outputs(4646) <= not((layer3_outputs(872)) and (layer3_outputs(4406)));
    layer4_outputs(4647) <= (layer3_outputs(3442)) and (layer3_outputs(787));
    layer4_outputs(4648) <= not(layer3_outputs(2492)) or (layer3_outputs(4471));
    layer4_outputs(4649) <= not(layer3_outputs(3001));
    layer4_outputs(4650) <= not((layer3_outputs(4640)) or (layer3_outputs(1885)));
    layer4_outputs(4651) <= not(layer3_outputs(1757)) or (layer3_outputs(4213));
    layer4_outputs(4652) <= '0';
    layer4_outputs(4653) <= (layer3_outputs(3691)) and (layer3_outputs(4486));
    layer4_outputs(4654) <= not((layer3_outputs(4730)) or (layer3_outputs(5091)));
    layer4_outputs(4655) <= (layer3_outputs(2428)) and (layer3_outputs(1130));
    layer4_outputs(4656) <= not(layer3_outputs(2799)) or (layer3_outputs(643));
    layer4_outputs(4657) <= (layer3_outputs(582)) and not (layer3_outputs(304));
    layer4_outputs(4658) <= not(layer3_outputs(4597));
    layer4_outputs(4659) <= '1';
    layer4_outputs(4660) <= '1';
    layer4_outputs(4661) <= not((layer3_outputs(3009)) or (layer3_outputs(3238)));
    layer4_outputs(4662) <= not(layer3_outputs(2267));
    layer4_outputs(4663) <= not(layer3_outputs(4097));
    layer4_outputs(4664) <= layer3_outputs(280);
    layer4_outputs(4665) <= (layer3_outputs(4964)) or (layer3_outputs(1189));
    layer4_outputs(4666) <= not(layer3_outputs(2698));
    layer4_outputs(4667) <= not((layer3_outputs(2536)) and (layer3_outputs(1613)));
    layer4_outputs(4668) <= not((layer3_outputs(1850)) and (layer3_outputs(3674)));
    layer4_outputs(4669) <= not(layer3_outputs(1091));
    layer4_outputs(4670) <= '0';
    layer4_outputs(4671) <= not(layer3_outputs(2925)) or (layer3_outputs(1147));
    layer4_outputs(4672) <= not((layer3_outputs(5019)) xor (layer3_outputs(3399)));
    layer4_outputs(4673) <= layer3_outputs(153);
    layer4_outputs(4674) <= (layer3_outputs(2848)) and (layer3_outputs(863));
    layer4_outputs(4675) <= not(layer3_outputs(4577)) or (layer3_outputs(1991));
    layer4_outputs(4676) <= '1';
    layer4_outputs(4677) <= (layer3_outputs(2256)) and not (layer3_outputs(4297));
    layer4_outputs(4678) <= (layer3_outputs(672)) and not (layer3_outputs(1169));
    layer4_outputs(4679) <= layer3_outputs(544);
    layer4_outputs(4680) <= not(layer3_outputs(871));
    layer4_outputs(4681) <= not((layer3_outputs(637)) and (layer3_outputs(4266)));
    layer4_outputs(4682) <= '0';
    layer4_outputs(4683) <= not(layer3_outputs(2714)) or (layer3_outputs(160));
    layer4_outputs(4684) <= layer3_outputs(1329);
    layer4_outputs(4685) <= not((layer3_outputs(4850)) and (layer3_outputs(2827)));
    layer4_outputs(4686) <= not(layer3_outputs(4272)) or (layer3_outputs(3905));
    layer4_outputs(4687) <= not((layer3_outputs(5084)) and (layer3_outputs(1673)));
    layer4_outputs(4688) <= '1';
    layer4_outputs(4689) <= '1';
    layer4_outputs(4690) <= '0';
    layer4_outputs(4691) <= not((layer3_outputs(808)) and (layer3_outputs(1194)));
    layer4_outputs(4692) <= not(layer3_outputs(734)) or (layer3_outputs(1810));
    layer4_outputs(4693) <= layer3_outputs(1617);
    layer4_outputs(4694) <= (layer3_outputs(454)) and (layer3_outputs(3976));
    layer4_outputs(4695) <= (layer3_outputs(2580)) and (layer3_outputs(2217));
    layer4_outputs(4696) <= layer3_outputs(2655);
    layer4_outputs(4697) <= layer3_outputs(2764);
    layer4_outputs(4698) <= not((layer3_outputs(3220)) and (layer3_outputs(758)));
    layer4_outputs(4699) <= (layer3_outputs(3628)) or (layer3_outputs(4853));
    layer4_outputs(4700) <= '1';
    layer4_outputs(4701) <= (layer3_outputs(1236)) and (layer3_outputs(3013));
    layer4_outputs(4702) <= layer3_outputs(3481);
    layer4_outputs(4703) <= layer3_outputs(3897);
    layer4_outputs(4704) <= (layer3_outputs(4149)) and not (layer3_outputs(2288));
    layer4_outputs(4705) <= not(layer3_outputs(4697));
    layer4_outputs(4706) <= not(layer3_outputs(4118)) or (layer3_outputs(225));
    layer4_outputs(4707) <= not(layer3_outputs(4165));
    layer4_outputs(4708) <= not((layer3_outputs(4770)) and (layer3_outputs(4587)));
    layer4_outputs(4709) <= not(layer3_outputs(1958)) or (layer3_outputs(2719));
    layer4_outputs(4710) <= not(layer3_outputs(3359)) or (layer3_outputs(3043));
    layer4_outputs(4711) <= not((layer3_outputs(1812)) or (layer3_outputs(3573)));
    layer4_outputs(4712) <= layer3_outputs(598);
    layer4_outputs(4713) <= (layer3_outputs(3382)) and not (layer3_outputs(2465));
    layer4_outputs(4714) <= (layer3_outputs(2166)) and not (layer3_outputs(1989));
    layer4_outputs(4715) <= (layer3_outputs(3525)) and (layer3_outputs(3088));
    layer4_outputs(4716) <= (layer3_outputs(2557)) and not (layer3_outputs(4940));
    layer4_outputs(4717) <= not(layer3_outputs(3829)) or (layer3_outputs(4875));
    layer4_outputs(4718) <= (layer3_outputs(4371)) and (layer3_outputs(4964));
    layer4_outputs(4719) <= layer3_outputs(378);
    layer4_outputs(4720) <= layer3_outputs(3424);
    layer4_outputs(4721) <= not(layer3_outputs(3502)) or (layer3_outputs(1074));
    layer4_outputs(4722) <= (layer3_outputs(1689)) and (layer3_outputs(5052));
    layer4_outputs(4723) <= (layer3_outputs(145)) or (layer3_outputs(3756));
    layer4_outputs(4724) <= '0';
    layer4_outputs(4725) <= (layer3_outputs(2768)) and not (layer3_outputs(326));
    layer4_outputs(4726) <= not((layer3_outputs(4510)) and (layer3_outputs(834)));
    layer4_outputs(4727) <= (layer3_outputs(2264)) or (layer3_outputs(1308));
    layer4_outputs(4728) <= (layer3_outputs(1465)) and not (layer3_outputs(910));
    layer4_outputs(4729) <= (layer3_outputs(1935)) or (layer3_outputs(4151));
    layer4_outputs(4730) <= not(layer3_outputs(3496));
    layer4_outputs(4731) <= layer3_outputs(2580);
    layer4_outputs(4732) <= not((layer3_outputs(4866)) and (layer3_outputs(3354)));
    layer4_outputs(4733) <= (layer3_outputs(3445)) xor (layer3_outputs(1710));
    layer4_outputs(4734) <= layer3_outputs(2026);
    layer4_outputs(4735) <= (layer3_outputs(319)) and not (layer3_outputs(4178));
    layer4_outputs(4736) <= not((layer3_outputs(2027)) and (layer3_outputs(4976)));
    layer4_outputs(4737) <= not(layer3_outputs(4081)) or (layer3_outputs(3764));
    layer4_outputs(4738) <= '1';
    layer4_outputs(4739) <= (layer3_outputs(798)) and not (layer3_outputs(1809));
    layer4_outputs(4740) <= not(layer3_outputs(2824));
    layer4_outputs(4741) <= (layer3_outputs(2669)) and (layer3_outputs(4841));
    layer4_outputs(4742) <= not(layer3_outputs(309));
    layer4_outputs(4743) <= not(layer3_outputs(2618));
    layer4_outputs(4744) <= (layer3_outputs(2496)) and (layer3_outputs(1985));
    layer4_outputs(4745) <= layer3_outputs(3995);
    layer4_outputs(4746) <= not((layer3_outputs(2666)) or (layer3_outputs(3842)));
    layer4_outputs(4747) <= not((layer3_outputs(3147)) and (layer3_outputs(3900)));
    layer4_outputs(4748) <= (layer3_outputs(5022)) or (layer3_outputs(1644));
    layer4_outputs(4749) <= (layer3_outputs(4517)) or (layer3_outputs(2504));
    layer4_outputs(4750) <= (layer3_outputs(1577)) or (layer3_outputs(1412));
    layer4_outputs(4751) <= layer3_outputs(1289);
    layer4_outputs(4752) <= '0';
    layer4_outputs(4753) <= (layer3_outputs(3518)) and (layer3_outputs(1335));
    layer4_outputs(4754) <= not(layer3_outputs(3090));
    layer4_outputs(4755) <= '1';
    layer4_outputs(4756) <= (layer3_outputs(2032)) or (layer3_outputs(3002));
    layer4_outputs(4757) <= '1';
    layer4_outputs(4758) <= not((layer3_outputs(4375)) xor (layer3_outputs(5116)));
    layer4_outputs(4759) <= not(layer3_outputs(922));
    layer4_outputs(4760) <= (layer3_outputs(4981)) and not (layer3_outputs(4197));
    layer4_outputs(4761) <= (layer3_outputs(4988)) and (layer3_outputs(4340));
    layer4_outputs(4762) <= not(layer3_outputs(25));
    layer4_outputs(4763) <= not((layer3_outputs(4352)) xor (layer3_outputs(1298)));
    layer4_outputs(4764) <= not((layer3_outputs(1658)) or (layer3_outputs(567)));
    layer4_outputs(4765) <= not(layer3_outputs(3478)) or (layer3_outputs(1188));
    layer4_outputs(4766) <= '0';
    layer4_outputs(4767) <= (layer3_outputs(3122)) or (layer3_outputs(1828));
    layer4_outputs(4768) <= layer3_outputs(309);
    layer4_outputs(4769) <= not(layer3_outputs(4637));
    layer4_outputs(4770) <= layer3_outputs(532);
    layer4_outputs(4771) <= not(layer3_outputs(692));
    layer4_outputs(4772) <= (layer3_outputs(2198)) or (layer3_outputs(2455));
    layer4_outputs(4773) <= (layer3_outputs(3937)) or (layer3_outputs(2961));
    layer4_outputs(4774) <= (layer3_outputs(453)) and not (layer3_outputs(3907));
    layer4_outputs(4775) <= not(layer3_outputs(1627));
    layer4_outputs(4776) <= not(layer3_outputs(3822)) or (layer3_outputs(3282));
    layer4_outputs(4777) <= '1';
    layer4_outputs(4778) <= not((layer3_outputs(486)) or (layer3_outputs(2958)));
    layer4_outputs(4779) <= not(layer3_outputs(2303)) or (layer3_outputs(816));
    layer4_outputs(4780) <= (layer3_outputs(4152)) and (layer3_outputs(5003));
    layer4_outputs(4781) <= not(layer3_outputs(529));
    layer4_outputs(4782) <= '1';
    layer4_outputs(4783) <= not(layer3_outputs(4962));
    layer4_outputs(4784) <= (layer3_outputs(2652)) or (layer3_outputs(1425));
    layer4_outputs(4785) <= '0';
    layer4_outputs(4786) <= not((layer3_outputs(492)) and (layer3_outputs(364)));
    layer4_outputs(4787) <= not(layer3_outputs(657)) or (layer3_outputs(959));
    layer4_outputs(4788) <= not((layer3_outputs(2895)) and (layer3_outputs(1207)));
    layer4_outputs(4789) <= (layer3_outputs(4177)) and (layer3_outputs(4529));
    layer4_outputs(4790) <= layer3_outputs(1579);
    layer4_outputs(4791) <= (layer3_outputs(1630)) or (layer3_outputs(1769));
    layer4_outputs(4792) <= (layer3_outputs(3640)) or (layer3_outputs(2900));
    layer4_outputs(4793) <= not(layer3_outputs(863)) or (layer3_outputs(896));
    layer4_outputs(4794) <= layer3_outputs(3439);
    layer4_outputs(4795) <= not(layer3_outputs(812));
    layer4_outputs(4796) <= layer3_outputs(2801);
    layer4_outputs(4797) <= '1';
    layer4_outputs(4798) <= not((layer3_outputs(563)) and (layer3_outputs(85)));
    layer4_outputs(4799) <= layer3_outputs(2744);
    layer4_outputs(4800) <= not(layer3_outputs(1680)) or (layer3_outputs(4446));
    layer4_outputs(4801) <= (layer3_outputs(1822)) or (layer3_outputs(1165));
    layer4_outputs(4802) <= not(layer3_outputs(648));
    layer4_outputs(4803) <= not(layer3_outputs(1166)) or (layer3_outputs(4870));
    layer4_outputs(4804) <= (layer3_outputs(731)) and not (layer3_outputs(2387));
    layer4_outputs(4805) <= not(layer3_outputs(2093)) or (layer3_outputs(4680));
    layer4_outputs(4806) <= (layer3_outputs(3592)) and not (layer3_outputs(4610));
    layer4_outputs(4807) <= (layer3_outputs(3674)) and not (layer3_outputs(4099));
    layer4_outputs(4808) <= '1';
    layer4_outputs(4809) <= (layer3_outputs(1046)) and not (layer3_outputs(675));
    layer4_outputs(4810) <= not(layer3_outputs(2408)) or (layer3_outputs(684));
    layer4_outputs(4811) <= (layer3_outputs(813)) and not (layer3_outputs(1908));
    layer4_outputs(4812) <= (layer3_outputs(1151)) or (layer3_outputs(689));
    layer4_outputs(4813) <= (layer3_outputs(4313)) and not (layer3_outputs(3126));
    layer4_outputs(4814) <= not((layer3_outputs(362)) or (layer3_outputs(1563)));
    layer4_outputs(4815) <= (layer3_outputs(4685)) and not (layer3_outputs(3291));
    layer4_outputs(4816) <= layer3_outputs(1174);
    layer4_outputs(4817) <= (layer3_outputs(1467)) and not (layer3_outputs(3428));
    layer4_outputs(4818) <= layer3_outputs(4585);
    layer4_outputs(4819) <= not((layer3_outputs(825)) and (layer3_outputs(879)));
    layer4_outputs(4820) <= not(layer3_outputs(2779)) or (layer3_outputs(3004));
    layer4_outputs(4821) <= not(layer3_outputs(4689));
    layer4_outputs(4822) <= '1';
    layer4_outputs(4823) <= (layer3_outputs(1493)) and not (layer3_outputs(4303));
    layer4_outputs(4824) <= (layer3_outputs(1422)) and not (layer3_outputs(4507));
    layer4_outputs(4825) <= not((layer3_outputs(2888)) and (layer3_outputs(4032)));
    layer4_outputs(4826) <= '1';
    layer4_outputs(4827) <= not(layer3_outputs(3261));
    layer4_outputs(4828) <= (layer3_outputs(38)) and not (layer3_outputs(3719));
    layer4_outputs(4829) <= (layer3_outputs(3938)) or (layer3_outputs(4707));
    layer4_outputs(4830) <= layer3_outputs(4045);
    layer4_outputs(4831) <= not(layer3_outputs(1356)) or (layer3_outputs(3130));
    layer4_outputs(4832) <= layer3_outputs(3629);
    layer4_outputs(4833) <= (layer3_outputs(39)) and not (layer3_outputs(370));
    layer4_outputs(4834) <= (layer3_outputs(530)) and not (layer3_outputs(2981));
    layer4_outputs(4835) <= (layer3_outputs(4782)) and (layer3_outputs(2718));
    layer4_outputs(4836) <= layer3_outputs(3546);
    layer4_outputs(4837) <= layer3_outputs(1081);
    layer4_outputs(4838) <= (layer3_outputs(4455)) and not (layer3_outputs(1671));
    layer4_outputs(4839) <= '1';
    layer4_outputs(4840) <= not(layer3_outputs(3488)) or (layer3_outputs(443));
    layer4_outputs(4841) <= '0';
    layer4_outputs(4842) <= layer3_outputs(1695);
    layer4_outputs(4843) <= (layer3_outputs(2970)) and not (layer3_outputs(4477));
    layer4_outputs(4844) <= not((layer3_outputs(991)) and (layer3_outputs(1849)));
    layer4_outputs(4845) <= (layer3_outputs(1981)) and (layer3_outputs(476));
    layer4_outputs(4846) <= layer3_outputs(1486);
    layer4_outputs(4847) <= layer3_outputs(2656);
    layer4_outputs(4848) <= '0';
    layer4_outputs(4849) <= (layer3_outputs(1294)) or (layer3_outputs(4228));
    layer4_outputs(4850) <= (layer3_outputs(3930)) and not (layer3_outputs(2964));
    layer4_outputs(4851) <= not(layer3_outputs(4825));
    layer4_outputs(4852) <= (layer3_outputs(4398)) and not (layer3_outputs(4367));
    layer4_outputs(4853) <= '0';
    layer4_outputs(4854) <= (layer3_outputs(3988)) and not (layer3_outputs(3454));
    layer4_outputs(4855) <= (layer3_outputs(3971)) and not (layer3_outputs(1672));
    layer4_outputs(4856) <= not(layer3_outputs(3748));
    layer4_outputs(4857) <= not((layer3_outputs(4821)) or (layer3_outputs(2509)));
    layer4_outputs(4858) <= not(layer3_outputs(2839));
    layer4_outputs(4859) <= layer3_outputs(1054);
    layer4_outputs(4860) <= (layer3_outputs(2916)) and (layer3_outputs(248));
    layer4_outputs(4861) <= not(layer3_outputs(2812)) or (layer3_outputs(1305));
    layer4_outputs(4862) <= not((layer3_outputs(3286)) xor (layer3_outputs(3179)));
    layer4_outputs(4863) <= '0';
    layer4_outputs(4864) <= layer3_outputs(274);
    layer4_outputs(4865) <= not((layer3_outputs(1115)) or (layer3_outputs(2687)));
    layer4_outputs(4866) <= not((layer3_outputs(2441)) and (layer3_outputs(2281)));
    layer4_outputs(4867) <= not(layer3_outputs(4455));
    layer4_outputs(4868) <= (layer3_outputs(4928)) and (layer3_outputs(882));
    layer4_outputs(4869) <= layer3_outputs(4496);
    layer4_outputs(4870) <= layer3_outputs(2435);
    layer4_outputs(4871) <= not(layer3_outputs(3686)) or (layer3_outputs(3041));
    layer4_outputs(4872) <= not(layer3_outputs(2404));
    layer4_outputs(4873) <= layer3_outputs(130);
    layer4_outputs(4874) <= not(layer3_outputs(1733));
    layer4_outputs(4875) <= not(layer3_outputs(3233)) or (layer3_outputs(870));
    layer4_outputs(4876) <= '1';
    layer4_outputs(4877) <= (layer3_outputs(3577)) and not (layer3_outputs(4800));
    layer4_outputs(4878) <= not(layer3_outputs(2341));
    layer4_outputs(4879) <= layer3_outputs(594);
    layer4_outputs(4880) <= (layer3_outputs(269)) and (layer3_outputs(5083));
    layer4_outputs(4881) <= not(layer3_outputs(3253)) or (layer3_outputs(3249));
    layer4_outputs(4882) <= layer3_outputs(505);
    layer4_outputs(4883) <= not(layer3_outputs(3427)) or (layer3_outputs(27));
    layer4_outputs(4884) <= not(layer3_outputs(2088));
    layer4_outputs(4885) <= not(layer3_outputs(3374));
    layer4_outputs(4886) <= layer3_outputs(493);
    layer4_outputs(4887) <= layer3_outputs(4202);
    layer4_outputs(4888) <= not(layer3_outputs(3141));
    layer4_outputs(4889) <= not((layer3_outputs(4452)) or (layer3_outputs(4120)));
    layer4_outputs(4890) <= (layer3_outputs(1097)) and not (layer3_outputs(1114));
    layer4_outputs(4891) <= not(layer3_outputs(146)) or (layer3_outputs(255));
    layer4_outputs(4892) <= not((layer3_outputs(4580)) and (layer3_outputs(15)));
    layer4_outputs(4893) <= not(layer3_outputs(407)) or (layer3_outputs(3083));
    layer4_outputs(4894) <= (layer3_outputs(3695)) and not (layer3_outputs(1226));
    layer4_outputs(4895) <= not(layer3_outputs(3514));
    layer4_outputs(4896) <= (layer3_outputs(2334)) and not (layer3_outputs(1079));
    layer4_outputs(4897) <= not(layer3_outputs(4296));
    layer4_outputs(4898) <= not((layer3_outputs(1487)) or (layer3_outputs(1451)));
    layer4_outputs(4899) <= (layer3_outputs(691)) and not (layer3_outputs(1607));
    layer4_outputs(4900) <= not((layer3_outputs(3157)) and (layer3_outputs(1836)));
    layer4_outputs(4901) <= (layer3_outputs(580)) xor (layer3_outputs(755));
    layer4_outputs(4902) <= (layer3_outputs(5077)) and not (layer3_outputs(5042));
    layer4_outputs(4903) <= layer3_outputs(3713);
    layer4_outputs(4904) <= layer3_outputs(22);
    layer4_outputs(4905) <= '0';
    layer4_outputs(4906) <= (layer3_outputs(4391)) or (layer3_outputs(159));
    layer4_outputs(4907) <= layer3_outputs(91);
    layer4_outputs(4908) <= '1';
    layer4_outputs(4909) <= '0';
    layer4_outputs(4910) <= (layer3_outputs(2697)) and not (layer3_outputs(3729));
    layer4_outputs(4911) <= not((layer3_outputs(2398)) and (layer3_outputs(1234)));
    layer4_outputs(4912) <= not((layer3_outputs(4458)) and (layer3_outputs(3262)));
    layer4_outputs(4913) <= layer3_outputs(2120);
    layer4_outputs(4914) <= (layer3_outputs(2581)) xor (layer3_outputs(4710));
    layer4_outputs(4915) <= not((layer3_outputs(1675)) and (layer3_outputs(3814)));
    layer4_outputs(4916) <= not(layer3_outputs(4475)) or (layer3_outputs(3488));
    layer4_outputs(4917) <= not((layer3_outputs(923)) or (layer3_outputs(1959)));
    layer4_outputs(4918) <= (layer3_outputs(690)) or (layer3_outputs(2963));
    layer4_outputs(4919) <= layer3_outputs(483);
    layer4_outputs(4920) <= (layer3_outputs(2254)) xor (layer3_outputs(3186));
    layer4_outputs(4921) <= (layer3_outputs(811)) and not (layer3_outputs(1632));
    layer4_outputs(4922) <= layer3_outputs(2738);
    layer4_outputs(4923) <= layer3_outputs(3978);
    layer4_outputs(4924) <= layer3_outputs(3345);
    layer4_outputs(4925) <= (layer3_outputs(2584)) and not (layer3_outputs(2213));
    layer4_outputs(4926) <= '1';
    layer4_outputs(4927) <= not(layer3_outputs(872)) or (layer3_outputs(2470));
    layer4_outputs(4928) <= (layer3_outputs(4035)) and not (layer3_outputs(4110));
    layer4_outputs(4929) <= (layer3_outputs(1042)) and (layer3_outputs(2370));
    layer4_outputs(4930) <= not(layer3_outputs(45)) or (layer3_outputs(1492));
    layer4_outputs(4931) <= layer3_outputs(4225);
    layer4_outputs(4932) <= not(layer3_outputs(4855)) or (layer3_outputs(3374));
    layer4_outputs(4933) <= layer3_outputs(3170);
    layer4_outputs(4934) <= '0';
    layer4_outputs(4935) <= (layer3_outputs(1099)) and not (layer3_outputs(2307));
    layer4_outputs(4936) <= not(layer3_outputs(451));
    layer4_outputs(4937) <= (layer3_outputs(66)) and (layer3_outputs(3687));
    layer4_outputs(4938) <= not(layer3_outputs(4320)) or (layer3_outputs(3481));
    layer4_outputs(4939) <= layer3_outputs(3609);
    layer4_outputs(4940) <= layer3_outputs(200);
    layer4_outputs(4941) <= (layer3_outputs(2739)) and (layer3_outputs(4090));
    layer4_outputs(4942) <= not(layer3_outputs(2648));
    layer4_outputs(4943) <= (layer3_outputs(3880)) or (layer3_outputs(1137));
    layer4_outputs(4944) <= '0';
    layer4_outputs(4945) <= layer3_outputs(1406);
    layer4_outputs(4946) <= not(layer3_outputs(4922)) or (layer3_outputs(5118));
    layer4_outputs(4947) <= not(layer3_outputs(460)) or (layer3_outputs(4873));
    layer4_outputs(4948) <= (layer3_outputs(967)) or (layer3_outputs(4688));
    layer4_outputs(4949) <= (layer3_outputs(1471)) and (layer3_outputs(2807));
    layer4_outputs(4950) <= (layer3_outputs(2094)) and not (layer3_outputs(480));
    layer4_outputs(4951) <= (layer3_outputs(2420)) or (layer3_outputs(1069));
    layer4_outputs(4952) <= layer3_outputs(3183);
    layer4_outputs(4953) <= not(layer3_outputs(1330));
    layer4_outputs(4954) <= (layer3_outputs(2775)) and not (layer3_outputs(3699));
    layer4_outputs(4955) <= not((layer3_outputs(3330)) and (layer3_outputs(3033)));
    layer4_outputs(4956) <= layer3_outputs(3315);
    layer4_outputs(4957) <= not(layer3_outputs(4797));
    layer4_outputs(4958) <= not(layer3_outputs(1762));
    layer4_outputs(4959) <= layer3_outputs(4033);
    layer4_outputs(4960) <= not(layer3_outputs(2623));
    layer4_outputs(4961) <= layer3_outputs(1377);
    layer4_outputs(4962) <= not((layer3_outputs(4479)) and (layer3_outputs(2253)));
    layer4_outputs(4963) <= not(layer3_outputs(2394));
    layer4_outputs(4964) <= not(layer3_outputs(156));
    layer4_outputs(4965) <= layer3_outputs(2267);
    layer4_outputs(4966) <= (layer3_outputs(69)) and not (layer3_outputs(608));
    layer4_outputs(4967) <= (layer3_outputs(2359)) xor (layer3_outputs(885));
    layer4_outputs(4968) <= not(layer3_outputs(1282));
    layer4_outputs(4969) <= layer3_outputs(3815);
    layer4_outputs(4970) <= not(layer3_outputs(5034));
    layer4_outputs(4971) <= '0';
    layer4_outputs(4972) <= '0';
    layer4_outputs(4973) <= layer3_outputs(2615);
    layer4_outputs(4974) <= (layer3_outputs(3462)) and (layer3_outputs(941));
    layer4_outputs(4975) <= '0';
    layer4_outputs(4976) <= (layer3_outputs(3408)) or (layer3_outputs(2044));
    layer4_outputs(4977) <= not(layer3_outputs(4598)) or (layer3_outputs(1121));
    layer4_outputs(4978) <= (layer3_outputs(2418)) and not (layer3_outputs(4411));
    layer4_outputs(4979) <= (layer3_outputs(130)) and not (layer3_outputs(4096));
    layer4_outputs(4980) <= not(layer3_outputs(1474)) or (layer3_outputs(1497));
    layer4_outputs(4981) <= not(layer3_outputs(2240)) or (layer3_outputs(293));
    layer4_outputs(4982) <= '0';
    layer4_outputs(4983) <= '1';
    layer4_outputs(4984) <= '0';
    layer4_outputs(4985) <= (layer3_outputs(1322)) and not (layer3_outputs(4448));
    layer4_outputs(4986) <= not((layer3_outputs(4499)) and (layer3_outputs(3442)));
    layer4_outputs(4987) <= not((layer3_outputs(3791)) or (layer3_outputs(1334)));
    layer4_outputs(4988) <= layer3_outputs(2152);
    layer4_outputs(4989) <= '1';
    layer4_outputs(4990) <= (layer3_outputs(2990)) and not (layer3_outputs(4537));
    layer4_outputs(4991) <= '1';
    layer4_outputs(4992) <= layer3_outputs(2853);
    layer4_outputs(4993) <= (layer3_outputs(99)) and not (layer3_outputs(1743));
    layer4_outputs(4994) <= not(layer3_outputs(3365));
    layer4_outputs(4995) <= not((layer3_outputs(1295)) and (layer3_outputs(3019)));
    layer4_outputs(4996) <= (layer3_outputs(2468)) and not (layer3_outputs(457));
    layer4_outputs(4997) <= not(layer3_outputs(4626));
    layer4_outputs(4998) <= (layer3_outputs(3662)) or (layer3_outputs(1594));
    layer4_outputs(4999) <= not(layer3_outputs(4773));
    layer4_outputs(5000) <= not(layer3_outputs(1065)) or (layer3_outputs(1278));
    layer4_outputs(5001) <= not((layer3_outputs(3260)) or (layer3_outputs(1043)));
    layer4_outputs(5002) <= '0';
    layer4_outputs(5003) <= (layer3_outputs(2512)) or (layer3_outputs(2478));
    layer4_outputs(5004) <= layer3_outputs(822);
    layer4_outputs(5005) <= not((layer3_outputs(2590)) or (layer3_outputs(392)));
    layer4_outputs(5006) <= (layer3_outputs(4736)) and (layer3_outputs(2257));
    layer4_outputs(5007) <= not((layer3_outputs(4790)) or (layer3_outputs(1862)));
    layer4_outputs(5008) <= (layer3_outputs(3770)) and not (layer3_outputs(600));
    layer4_outputs(5009) <= (layer3_outputs(4525)) and not (layer3_outputs(4064));
    layer4_outputs(5010) <= not(layer3_outputs(3648));
    layer4_outputs(5011) <= not(layer3_outputs(2109)) or (layer3_outputs(3616));
    layer4_outputs(5012) <= (layer3_outputs(1319)) and not (layer3_outputs(3923));
    layer4_outputs(5013) <= layer3_outputs(4013);
    layer4_outputs(5014) <= '0';
    layer4_outputs(5015) <= layer3_outputs(4416);
    layer4_outputs(5016) <= (layer3_outputs(3770)) and (layer3_outputs(1789));
    layer4_outputs(5017) <= layer3_outputs(1730);
    layer4_outputs(5018) <= layer3_outputs(223);
    layer4_outputs(5019) <= '1';
    layer4_outputs(5020) <= not(layer3_outputs(1881));
    layer4_outputs(5021) <= (layer3_outputs(4215)) and not (layer3_outputs(4346));
    layer4_outputs(5022) <= '0';
    layer4_outputs(5023) <= (layer3_outputs(2336)) or (layer3_outputs(4402));
    layer4_outputs(5024) <= (layer3_outputs(390)) or (layer3_outputs(2097));
    layer4_outputs(5025) <= '1';
    layer4_outputs(5026) <= layer3_outputs(3849);
    layer4_outputs(5027) <= (layer3_outputs(4102)) xor (layer3_outputs(4848));
    layer4_outputs(5028) <= '1';
    layer4_outputs(5029) <= not(layer3_outputs(3969));
    layer4_outputs(5030) <= layer3_outputs(5000);
    layer4_outputs(5031) <= '0';
    layer4_outputs(5032) <= (layer3_outputs(4941)) and (layer3_outputs(3907));
    layer4_outputs(5033) <= not((layer3_outputs(2287)) and (layer3_outputs(2830)));
    layer4_outputs(5034) <= not((layer3_outputs(3450)) and (layer3_outputs(1090)));
    layer4_outputs(5035) <= not((layer3_outputs(3369)) and (layer3_outputs(4493)));
    layer4_outputs(5036) <= layer3_outputs(4943);
    layer4_outputs(5037) <= '0';
    layer4_outputs(5038) <= not(layer3_outputs(5070)) or (layer3_outputs(2149));
    layer4_outputs(5039) <= not((layer3_outputs(4527)) and (layer3_outputs(1904)));
    layer4_outputs(5040) <= '0';
    layer4_outputs(5041) <= (layer3_outputs(392)) and (layer3_outputs(3484));
    layer4_outputs(5042) <= not((layer3_outputs(2443)) xor (layer3_outputs(5086)));
    layer4_outputs(5043) <= '1';
    layer4_outputs(5044) <= (layer3_outputs(4499)) and (layer3_outputs(270));
    layer4_outputs(5045) <= not((layer3_outputs(504)) and (layer3_outputs(3101)));
    layer4_outputs(5046) <= layer3_outputs(4080);
    layer4_outputs(5047) <= not(layer3_outputs(2378)) or (layer3_outputs(2390));
    layer4_outputs(5048) <= not(layer3_outputs(195)) or (layer3_outputs(660));
    layer4_outputs(5049) <= layer3_outputs(3309);
    layer4_outputs(5050) <= not(layer3_outputs(4865));
    layer4_outputs(5051) <= '1';
    layer4_outputs(5052) <= (layer3_outputs(1834)) or (layer3_outputs(3229));
    layer4_outputs(5053) <= not((layer3_outputs(2745)) or (layer3_outputs(4777)));
    layer4_outputs(5054) <= '0';
    layer4_outputs(5055) <= (layer3_outputs(1708)) and (layer3_outputs(3718));
    layer4_outputs(5056) <= not(layer3_outputs(302)) or (layer3_outputs(4995));
    layer4_outputs(5057) <= not(layer3_outputs(1687));
    layer4_outputs(5058) <= not((layer3_outputs(3335)) and (layer3_outputs(3201)));
    layer4_outputs(5059) <= (layer3_outputs(4041)) and (layer3_outputs(467));
    layer4_outputs(5060) <= not((layer3_outputs(639)) or (layer3_outputs(465)));
    layer4_outputs(5061) <= not(layer3_outputs(379)) or (layer3_outputs(642));
    layer4_outputs(5062) <= (layer3_outputs(1094)) and not (layer3_outputs(4482));
    layer4_outputs(5063) <= not(layer3_outputs(4882)) or (layer3_outputs(1001));
    layer4_outputs(5064) <= not(layer3_outputs(198)) or (layer3_outputs(4381));
    layer4_outputs(5065) <= layer3_outputs(2243);
    layer4_outputs(5066) <= (layer3_outputs(1777)) xor (layer3_outputs(20));
    layer4_outputs(5067) <= layer3_outputs(3098);
    layer4_outputs(5068) <= '0';
    layer4_outputs(5069) <= not(layer3_outputs(1836));
    layer4_outputs(5070) <= not((layer3_outputs(2799)) and (layer3_outputs(3380)));
    layer4_outputs(5071) <= '0';
    layer4_outputs(5072) <= '1';
    layer4_outputs(5073) <= (layer3_outputs(1185)) and not (layer3_outputs(2742));
    layer4_outputs(5074) <= '0';
    layer4_outputs(5075) <= (layer3_outputs(1707)) xor (layer3_outputs(4560));
    layer4_outputs(5076) <= not((layer3_outputs(1400)) or (layer3_outputs(1198)));
    layer4_outputs(5077) <= not(layer3_outputs(4093));
    layer4_outputs(5078) <= layer3_outputs(2935);
    layer4_outputs(5079) <= not(layer3_outputs(4208));
    layer4_outputs(5080) <= layer3_outputs(3736);
    layer4_outputs(5081) <= (layer3_outputs(5047)) and not (layer3_outputs(1810));
    layer4_outputs(5082) <= layer3_outputs(296);
    layer4_outputs(5083) <= (layer3_outputs(1180)) and (layer3_outputs(1618));
    layer4_outputs(5084) <= '0';
    layer4_outputs(5085) <= not((layer3_outputs(3858)) or (layer3_outputs(517)));
    layer4_outputs(5086) <= not(layer3_outputs(3865)) or (layer3_outputs(1534));
    layer4_outputs(5087) <= layer3_outputs(9);
    layer4_outputs(5088) <= (layer3_outputs(3888)) and not (layer3_outputs(1991));
    layer4_outputs(5089) <= not((layer3_outputs(2901)) and (layer3_outputs(4178)));
    layer4_outputs(5090) <= (layer3_outputs(2110)) or (layer3_outputs(1669));
    layer4_outputs(5091) <= (layer3_outputs(4148)) or (layer3_outputs(352));
    layer4_outputs(5092) <= (layer3_outputs(1900)) or (layer3_outputs(783));
    layer4_outputs(5093) <= layer3_outputs(960);
    layer4_outputs(5094) <= layer3_outputs(3326);
    layer4_outputs(5095) <= layer3_outputs(127);
    layer4_outputs(5096) <= (layer3_outputs(2283)) and not (layer3_outputs(3833));
    layer4_outputs(5097) <= not(layer3_outputs(3487));
    layer4_outputs(5098) <= (layer3_outputs(812)) and not (layer3_outputs(1119));
    layer4_outputs(5099) <= '1';
    layer4_outputs(5100) <= not(layer3_outputs(419));
    layer4_outputs(5101) <= '1';
    layer4_outputs(5102) <= not((layer3_outputs(3317)) and (layer3_outputs(2784)));
    layer4_outputs(5103) <= not((layer3_outputs(3551)) and (layer3_outputs(1719)));
    layer4_outputs(5104) <= (layer3_outputs(3340)) and not (layer3_outputs(3344));
    layer4_outputs(5105) <= (layer3_outputs(3533)) and not (layer3_outputs(3465));
    layer4_outputs(5106) <= not((layer3_outputs(1001)) or (layer3_outputs(875)));
    layer4_outputs(5107) <= layer3_outputs(1729);
    layer4_outputs(5108) <= not((layer3_outputs(877)) or (layer3_outputs(1441)));
    layer4_outputs(5109) <= '1';
    layer4_outputs(5110) <= not((layer3_outputs(4419)) or (layer3_outputs(973)));
    layer4_outputs(5111) <= layer3_outputs(1209);
    layer4_outputs(5112) <= '0';
    layer4_outputs(5113) <= layer3_outputs(139);
    layer4_outputs(5114) <= layer3_outputs(2769);
    layer4_outputs(5115) <= '1';
    layer4_outputs(5116) <= not(layer3_outputs(4961));
    layer4_outputs(5117) <= not(layer3_outputs(268));
    layer4_outputs(5118) <= not(layer3_outputs(2467)) or (layer3_outputs(3700));
    layer4_outputs(5119) <= (layer3_outputs(620)) xor (layer3_outputs(3078));
    layer5_outputs(0) <= '1';
    layer5_outputs(1) <= layer4_outputs(4132);
    layer5_outputs(2) <= not((layer4_outputs(2623)) or (layer4_outputs(651)));
    layer5_outputs(3) <= not(layer4_outputs(3572)) or (layer4_outputs(4932));
    layer5_outputs(4) <= (layer4_outputs(2924)) and (layer4_outputs(3725));
    layer5_outputs(5) <= (layer4_outputs(1065)) and not (layer4_outputs(1387));
    layer5_outputs(6) <= (layer4_outputs(3580)) and (layer4_outputs(3403));
    layer5_outputs(7) <= layer4_outputs(1279);
    layer5_outputs(8) <= not(layer4_outputs(145));
    layer5_outputs(9) <= (layer4_outputs(1260)) xor (layer4_outputs(1186));
    layer5_outputs(10) <= layer4_outputs(3242);
    layer5_outputs(11) <= not(layer4_outputs(1166));
    layer5_outputs(12) <= (layer4_outputs(1152)) or (layer4_outputs(665));
    layer5_outputs(13) <= not(layer4_outputs(1253));
    layer5_outputs(14) <= (layer4_outputs(1984)) or (layer4_outputs(3428));
    layer5_outputs(15) <= layer4_outputs(3763);
    layer5_outputs(16) <= layer4_outputs(1558);
    layer5_outputs(17) <= '0';
    layer5_outputs(18) <= not(layer4_outputs(3522));
    layer5_outputs(19) <= (layer4_outputs(4340)) and not (layer4_outputs(4136));
    layer5_outputs(20) <= (layer4_outputs(1085)) and not (layer4_outputs(2210));
    layer5_outputs(21) <= '0';
    layer5_outputs(22) <= layer4_outputs(1379);
    layer5_outputs(23) <= layer4_outputs(965);
    layer5_outputs(24) <= not((layer4_outputs(1939)) and (layer4_outputs(953)));
    layer5_outputs(25) <= layer4_outputs(2024);
    layer5_outputs(26) <= layer4_outputs(1462);
    layer5_outputs(27) <= layer4_outputs(3695);
    layer5_outputs(28) <= layer4_outputs(4500);
    layer5_outputs(29) <= layer4_outputs(2959);
    layer5_outputs(30) <= not((layer4_outputs(2433)) or (layer4_outputs(1162)));
    layer5_outputs(31) <= not((layer4_outputs(318)) and (layer4_outputs(3313)));
    layer5_outputs(32) <= not(layer4_outputs(4446));
    layer5_outputs(33) <= layer4_outputs(74);
    layer5_outputs(34) <= not(layer4_outputs(319)) or (layer4_outputs(4543));
    layer5_outputs(35) <= not(layer4_outputs(4397));
    layer5_outputs(36) <= layer4_outputs(4412);
    layer5_outputs(37) <= (layer4_outputs(159)) and not (layer4_outputs(3515));
    layer5_outputs(38) <= not((layer4_outputs(1392)) or (layer4_outputs(389)));
    layer5_outputs(39) <= layer4_outputs(3621);
    layer5_outputs(40) <= (layer4_outputs(3014)) xor (layer4_outputs(4953));
    layer5_outputs(41) <= not(layer4_outputs(2273));
    layer5_outputs(42) <= (layer4_outputs(3551)) and (layer4_outputs(492));
    layer5_outputs(43) <= (layer4_outputs(4151)) or (layer4_outputs(3772));
    layer5_outputs(44) <= not((layer4_outputs(75)) and (layer4_outputs(1866)));
    layer5_outputs(45) <= layer4_outputs(2405);
    layer5_outputs(46) <= '1';
    layer5_outputs(47) <= not((layer4_outputs(784)) and (layer4_outputs(3768)));
    layer5_outputs(48) <= not(layer4_outputs(2212)) or (layer4_outputs(5072));
    layer5_outputs(49) <= layer4_outputs(2977);
    layer5_outputs(50) <= not(layer4_outputs(3175)) or (layer4_outputs(3546));
    layer5_outputs(51) <= not(layer4_outputs(3425)) or (layer4_outputs(1760));
    layer5_outputs(52) <= (layer4_outputs(2825)) or (layer4_outputs(5057));
    layer5_outputs(53) <= layer4_outputs(2542);
    layer5_outputs(54) <= not(layer4_outputs(1736));
    layer5_outputs(55) <= not(layer4_outputs(2105)) or (layer4_outputs(180));
    layer5_outputs(56) <= not(layer4_outputs(4240));
    layer5_outputs(57) <= not(layer4_outputs(1412));
    layer5_outputs(58) <= not(layer4_outputs(2369));
    layer5_outputs(59) <= not(layer4_outputs(875)) or (layer4_outputs(1652));
    layer5_outputs(60) <= '1';
    layer5_outputs(61) <= '0';
    layer5_outputs(62) <= not(layer4_outputs(3026));
    layer5_outputs(63) <= not(layer4_outputs(4476));
    layer5_outputs(64) <= not(layer4_outputs(5081)) or (layer4_outputs(4544));
    layer5_outputs(65) <= layer4_outputs(283);
    layer5_outputs(66) <= layer4_outputs(1322);
    layer5_outputs(67) <= layer4_outputs(1430);
    layer5_outputs(68) <= (layer4_outputs(4629)) or (layer4_outputs(3588));
    layer5_outputs(69) <= not(layer4_outputs(4113));
    layer5_outputs(70) <= layer4_outputs(692);
    layer5_outputs(71) <= not(layer4_outputs(2168)) or (layer4_outputs(1466));
    layer5_outputs(72) <= layer4_outputs(769);
    layer5_outputs(73) <= not((layer4_outputs(916)) xor (layer4_outputs(1543)));
    layer5_outputs(74) <= (layer4_outputs(5007)) and (layer4_outputs(3891));
    layer5_outputs(75) <= (layer4_outputs(294)) and not (layer4_outputs(1183));
    layer5_outputs(76) <= not(layer4_outputs(1448));
    layer5_outputs(77) <= (layer4_outputs(4476)) and not (layer4_outputs(3768));
    layer5_outputs(78) <= not(layer4_outputs(3412));
    layer5_outputs(79) <= not(layer4_outputs(1783)) or (layer4_outputs(2598));
    layer5_outputs(80) <= not(layer4_outputs(3923)) or (layer4_outputs(4051));
    layer5_outputs(81) <= (layer4_outputs(4416)) and not (layer4_outputs(146));
    layer5_outputs(82) <= (layer4_outputs(2400)) xor (layer4_outputs(1796));
    layer5_outputs(83) <= (layer4_outputs(3399)) and not (layer4_outputs(3121));
    layer5_outputs(84) <= layer4_outputs(912);
    layer5_outputs(85) <= layer4_outputs(3780);
    layer5_outputs(86) <= not(layer4_outputs(3648));
    layer5_outputs(87) <= not(layer4_outputs(4845));
    layer5_outputs(88) <= (layer4_outputs(633)) and not (layer4_outputs(1287));
    layer5_outputs(89) <= not((layer4_outputs(4846)) and (layer4_outputs(4362)));
    layer5_outputs(90) <= '0';
    layer5_outputs(91) <= layer4_outputs(4472);
    layer5_outputs(92) <= layer4_outputs(3984);
    layer5_outputs(93) <= '1';
    layer5_outputs(94) <= layer4_outputs(397);
    layer5_outputs(95) <= not(layer4_outputs(4145));
    layer5_outputs(96) <= (layer4_outputs(660)) or (layer4_outputs(3935));
    layer5_outputs(97) <= layer4_outputs(4267);
    layer5_outputs(98) <= not(layer4_outputs(2644));
    layer5_outputs(99) <= (layer4_outputs(2333)) and (layer4_outputs(4713));
    layer5_outputs(100) <= not((layer4_outputs(2016)) or (layer4_outputs(4676)));
    layer5_outputs(101) <= (layer4_outputs(2118)) and not (layer4_outputs(5074));
    layer5_outputs(102) <= not(layer4_outputs(1051)) or (layer4_outputs(657));
    layer5_outputs(103) <= not((layer4_outputs(1286)) or (layer4_outputs(1033)));
    layer5_outputs(104) <= not(layer4_outputs(3715)) or (layer4_outputs(2412));
    layer5_outputs(105) <= not((layer4_outputs(2972)) or (layer4_outputs(106)));
    layer5_outputs(106) <= (layer4_outputs(4758)) and not (layer4_outputs(2463));
    layer5_outputs(107) <= (layer4_outputs(1058)) and (layer4_outputs(3555));
    layer5_outputs(108) <= '1';
    layer5_outputs(109) <= layer4_outputs(4904);
    layer5_outputs(110) <= (layer4_outputs(2155)) and not (layer4_outputs(3801));
    layer5_outputs(111) <= not((layer4_outputs(911)) and (layer4_outputs(794)));
    layer5_outputs(112) <= layer4_outputs(3876);
    layer5_outputs(113) <= (layer4_outputs(1122)) and not (layer4_outputs(3811));
    layer5_outputs(114) <= not((layer4_outputs(487)) or (layer4_outputs(4141)));
    layer5_outputs(115) <= not((layer4_outputs(3881)) or (layer4_outputs(1767)));
    layer5_outputs(116) <= '0';
    layer5_outputs(117) <= (layer4_outputs(1840)) and (layer4_outputs(1987));
    layer5_outputs(118) <= not(layer4_outputs(1783));
    layer5_outputs(119) <= not(layer4_outputs(738));
    layer5_outputs(120) <= layer4_outputs(4819);
    layer5_outputs(121) <= (layer4_outputs(3060)) and not (layer4_outputs(652));
    layer5_outputs(122) <= '1';
    layer5_outputs(123) <= (layer4_outputs(4017)) and (layer4_outputs(4462));
    layer5_outputs(124) <= (layer4_outputs(1363)) xor (layer4_outputs(2721));
    layer5_outputs(125) <= not(layer4_outputs(2896));
    layer5_outputs(126) <= '0';
    layer5_outputs(127) <= (layer4_outputs(2096)) and not (layer4_outputs(4996));
    layer5_outputs(128) <= layer4_outputs(1860);
    layer5_outputs(129) <= not((layer4_outputs(2868)) and (layer4_outputs(2465)));
    layer5_outputs(130) <= (layer4_outputs(4565)) and not (layer4_outputs(228));
    layer5_outputs(131) <= layer4_outputs(3782);
    layer5_outputs(132) <= not((layer4_outputs(2921)) and (layer4_outputs(4317)));
    layer5_outputs(133) <= not(layer4_outputs(987));
    layer5_outputs(134) <= not(layer4_outputs(3502)) or (layer4_outputs(705));
    layer5_outputs(135) <= '1';
    layer5_outputs(136) <= not(layer4_outputs(4223));
    layer5_outputs(137) <= not(layer4_outputs(1069)) or (layer4_outputs(2362));
    layer5_outputs(138) <= (layer4_outputs(3138)) and not (layer4_outputs(4272));
    layer5_outputs(139) <= '1';
    layer5_outputs(140) <= '1';
    layer5_outputs(141) <= layer4_outputs(4810);
    layer5_outputs(142) <= layer4_outputs(1262);
    layer5_outputs(143) <= (layer4_outputs(980)) or (layer4_outputs(670));
    layer5_outputs(144) <= layer4_outputs(130);
    layer5_outputs(145) <= (layer4_outputs(3560)) and not (layer4_outputs(2112));
    layer5_outputs(146) <= not(layer4_outputs(3701)) or (layer4_outputs(4104));
    layer5_outputs(147) <= (layer4_outputs(3072)) or (layer4_outputs(401));
    layer5_outputs(148) <= not((layer4_outputs(4557)) and (layer4_outputs(205)));
    layer5_outputs(149) <= not(layer4_outputs(3243)) or (layer4_outputs(2898));
    layer5_outputs(150) <= not(layer4_outputs(2728));
    layer5_outputs(151) <= layer4_outputs(2341);
    layer5_outputs(152) <= not((layer4_outputs(1057)) or (layer4_outputs(1148)));
    layer5_outputs(153) <= layer4_outputs(3655);
    layer5_outputs(154) <= not((layer4_outputs(1356)) xor (layer4_outputs(2062)));
    layer5_outputs(155) <= not(layer4_outputs(2198)) or (layer4_outputs(5063));
    layer5_outputs(156) <= layer4_outputs(151);
    layer5_outputs(157) <= layer4_outputs(5002);
    layer5_outputs(158) <= not(layer4_outputs(4859)) or (layer4_outputs(3746));
    layer5_outputs(159) <= not(layer4_outputs(4275)) or (layer4_outputs(2273));
    layer5_outputs(160) <= (layer4_outputs(4798)) or (layer4_outputs(3384));
    layer5_outputs(161) <= not(layer4_outputs(78));
    layer5_outputs(162) <= not(layer4_outputs(1770)) or (layer4_outputs(1541));
    layer5_outputs(163) <= (layer4_outputs(679)) and not (layer4_outputs(4303));
    layer5_outputs(164) <= layer4_outputs(758);
    layer5_outputs(165) <= (layer4_outputs(3535)) or (layer4_outputs(3311));
    layer5_outputs(166) <= (layer4_outputs(2659)) and not (layer4_outputs(1916));
    layer5_outputs(167) <= layer4_outputs(3716);
    layer5_outputs(168) <= layer4_outputs(4287);
    layer5_outputs(169) <= (layer4_outputs(3001)) xor (layer4_outputs(4762));
    layer5_outputs(170) <= (layer4_outputs(3776)) xor (layer4_outputs(3931));
    layer5_outputs(171) <= '0';
    layer5_outputs(172) <= layer4_outputs(1480);
    layer5_outputs(173) <= (layer4_outputs(364)) or (layer4_outputs(3927));
    layer5_outputs(174) <= not((layer4_outputs(2004)) or (layer4_outputs(3799)));
    layer5_outputs(175) <= not(layer4_outputs(2858));
    layer5_outputs(176) <= not(layer4_outputs(1878));
    layer5_outputs(177) <= not(layer4_outputs(4430)) or (layer4_outputs(5031));
    layer5_outputs(178) <= (layer4_outputs(1199)) and not (layer4_outputs(1747));
    layer5_outputs(179) <= '1';
    layer5_outputs(180) <= (layer4_outputs(4685)) or (layer4_outputs(1523));
    layer5_outputs(181) <= not(layer4_outputs(2966));
    layer5_outputs(182) <= not((layer4_outputs(2429)) or (layer4_outputs(4421)));
    layer5_outputs(183) <= not(layer4_outputs(134));
    layer5_outputs(184) <= not(layer4_outputs(1960));
    layer5_outputs(185) <= layer4_outputs(2487);
    layer5_outputs(186) <= layer4_outputs(3760);
    layer5_outputs(187) <= (layer4_outputs(354)) or (layer4_outputs(1284));
    layer5_outputs(188) <= '0';
    layer5_outputs(189) <= (layer4_outputs(3751)) and not (layer4_outputs(3669));
    layer5_outputs(190) <= not(layer4_outputs(2257)) or (layer4_outputs(2328));
    layer5_outputs(191) <= not(layer4_outputs(752));
    layer5_outputs(192) <= (layer4_outputs(1683)) or (layer4_outputs(357));
    layer5_outputs(193) <= (layer4_outputs(2694)) and not (layer4_outputs(828));
    layer5_outputs(194) <= not(layer4_outputs(3680));
    layer5_outputs(195) <= not(layer4_outputs(4056));
    layer5_outputs(196) <= (layer4_outputs(1578)) and not (layer4_outputs(1516));
    layer5_outputs(197) <= not(layer4_outputs(2725));
    layer5_outputs(198) <= (layer4_outputs(87)) and not (layer4_outputs(4896));
    layer5_outputs(199) <= (layer4_outputs(4630)) and not (layer4_outputs(864));
    layer5_outputs(200) <= not(layer4_outputs(252));
    layer5_outputs(201) <= not((layer4_outputs(4244)) and (layer4_outputs(1496)));
    layer5_outputs(202) <= layer4_outputs(3909);
    layer5_outputs(203) <= not((layer4_outputs(3339)) and (layer4_outputs(1203)));
    layer5_outputs(204) <= not((layer4_outputs(132)) and (layer4_outputs(1289)));
    layer5_outputs(205) <= not(layer4_outputs(4996));
    layer5_outputs(206) <= not((layer4_outputs(517)) and (layer4_outputs(31)));
    layer5_outputs(207) <= (layer4_outputs(3903)) and not (layer4_outputs(1998));
    layer5_outputs(208) <= not(layer4_outputs(571));
    layer5_outputs(209) <= '1';
    layer5_outputs(210) <= not((layer4_outputs(510)) xor (layer4_outputs(3884)));
    layer5_outputs(211) <= (layer4_outputs(72)) and not (layer4_outputs(4965));
    layer5_outputs(212) <= (layer4_outputs(1862)) and (layer4_outputs(1594));
    layer5_outputs(213) <= not(layer4_outputs(3625));
    layer5_outputs(214) <= not(layer4_outputs(4131));
    layer5_outputs(215) <= (layer4_outputs(1517)) xor (layer4_outputs(4888));
    layer5_outputs(216) <= (layer4_outputs(2363)) or (layer4_outputs(5052));
    layer5_outputs(217) <= not(layer4_outputs(3249));
    layer5_outputs(218) <= '0';
    layer5_outputs(219) <= not(layer4_outputs(1479));
    layer5_outputs(220) <= layer4_outputs(2472);
    layer5_outputs(221) <= not(layer4_outputs(5031));
    layer5_outputs(222) <= '1';
    layer5_outputs(223) <= not((layer4_outputs(3926)) xor (layer4_outputs(4658)));
    layer5_outputs(224) <= not(layer4_outputs(12));
    layer5_outputs(225) <= layer4_outputs(1511);
    layer5_outputs(226) <= not(layer4_outputs(3056));
    layer5_outputs(227) <= (layer4_outputs(4998)) or (layer4_outputs(1518));
    layer5_outputs(228) <= not(layer4_outputs(126));
    layer5_outputs(229) <= '1';
    layer5_outputs(230) <= not(layer4_outputs(1872));
    layer5_outputs(231) <= (layer4_outputs(2689)) and not (layer4_outputs(1942));
    layer5_outputs(232) <= not(layer4_outputs(4008)) or (layer4_outputs(932));
    layer5_outputs(233) <= '0';
    layer5_outputs(234) <= (layer4_outputs(1476)) or (layer4_outputs(4861));
    layer5_outputs(235) <= (layer4_outputs(1226)) and (layer4_outputs(3321));
    layer5_outputs(236) <= (layer4_outputs(595)) and not (layer4_outputs(3736));
    layer5_outputs(237) <= layer4_outputs(1765);
    layer5_outputs(238) <= not(layer4_outputs(1472));
    layer5_outputs(239) <= layer4_outputs(1479);
    layer5_outputs(240) <= not(layer4_outputs(3478));
    layer5_outputs(241) <= not(layer4_outputs(5082));
    layer5_outputs(242) <= '0';
    layer5_outputs(243) <= not(layer4_outputs(730)) or (layer4_outputs(1212));
    layer5_outputs(244) <= not(layer4_outputs(1325));
    layer5_outputs(245) <= layer4_outputs(5045);
    layer5_outputs(246) <= layer4_outputs(1216);
    layer5_outputs(247) <= not((layer4_outputs(4347)) and (layer4_outputs(3045)));
    layer5_outputs(248) <= '0';
    layer5_outputs(249) <= (layer4_outputs(4591)) and not (layer4_outputs(891));
    layer5_outputs(250) <= not(layer4_outputs(2254));
    layer5_outputs(251) <= layer4_outputs(598);
    layer5_outputs(252) <= layer4_outputs(2670);
    layer5_outputs(253) <= '0';
    layer5_outputs(254) <= not(layer4_outputs(2211));
    layer5_outputs(255) <= not(layer4_outputs(3118)) or (layer4_outputs(4550));
    layer5_outputs(256) <= layer4_outputs(3216);
    layer5_outputs(257) <= not(layer4_outputs(4659));
    layer5_outputs(258) <= not(layer4_outputs(1958)) or (layer4_outputs(2381));
    layer5_outputs(259) <= not(layer4_outputs(4846));
    layer5_outputs(260) <= not((layer4_outputs(2778)) xor (layer4_outputs(4919)));
    layer5_outputs(261) <= (layer4_outputs(1179)) and not (layer4_outputs(3160));
    layer5_outputs(262) <= not((layer4_outputs(604)) or (layer4_outputs(2604)));
    layer5_outputs(263) <= layer4_outputs(2895);
    layer5_outputs(264) <= (layer4_outputs(694)) and not (layer4_outputs(3961));
    layer5_outputs(265) <= (layer4_outputs(1912)) and (layer4_outputs(1005));
    layer5_outputs(266) <= '0';
    layer5_outputs(267) <= (layer4_outputs(2060)) and (layer4_outputs(3124));
    layer5_outputs(268) <= not(layer4_outputs(718));
    layer5_outputs(269) <= not(layer4_outputs(2864)) or (layer4_outputs(4150));
    layer5_outputs(270) <= (layer4_outputs(1666)) and (layer4_outputs(1138));
    layer5_outputs(271) <= layer4_outputs(3067);
    layer5_outputs(272) <= not(layer4_outputs(676));
    layer5_outputs(273) <= not((layer4_outputs(4962)) or (layer4_outputs(4787)));
    layer5_outputs(274) <= not(layer4_outputs(1879));
    layer5_outputs(275) <= layer4_outputs(3413);
    layer5_outputs(276) <= not(layer4_outputs(4367));
    layer5_outputs(277) <= not((layer4_outputs(4911)) or (layer4_outputs(2420)));
    layer5_outputs(278) <= (layer4_outputs(1919)) and (layer4_outputs(934));
    layer5_outputs(279) <= (layer4_outputs(1422)) and not (layer4_outputs(2285));
    layer5_outputs(280) <= not(layer4_outputs(1006));
    layer5_outputs(281) <= not((layer4_outputs(3364)) and (layer4_outputs(993)));
    layer5_outputs(282) <= (layer4_outputs(2579)) and not (layer4_outputs(605));
    layer5_outputs(283) <= layer4_outputs(1847);
    layer5_outputs(284) <= '0';
    layer5_outputs(285) <= (layer4_outputs(946)) and (layer4_outputs(528));
    layer5_outputs(286) <= layer4_outputs(1156);
    layer5_outputs(287) <= (layer4_outputs(108)) or (layer4_outputs(3214));
    layer5_outputs(288) <= layer4_outputs(4994);
    layer5_outputs(289) <= not((layer4_outputs(1624)) xor (layer4_outputs(4669)));
    layer5_outputs(290) <= (layer4_outputs(2162)) and not (layer4_outputs(978));
    layer5_outputs(291) <= (layer4_outputs(1153)) and (layer4_outputs(4244));
    layer5_outputs(292) <= layer4_outputs(1996);
    layer5_outputs(293) <= layer4_outputs(3026);
    layer5_outputs(294) <= (layer4_outputs(273)) and not (layer4_outputs(3356));
    layer5_outputs(295) <= (layer4_outputs(1533)) and not (layer4_outputs(650));
    layer5_outputs(296) <= '0';
    layer5_outputs(297) <= not(layer4_outputs(815));
    layer5_outputs(298) <= not((layer4_outputs(850)) xor (layer4_outputs(567)));
    layer5_outputs(299) <= (layer4_outputs(4857)) and not (layer4_outputs(3910));
    layer5_outputs(300) <= layer4_outputs(1541);
    layer5_outputs(301) <= not(layer4_outputs(3484));
    layer5_outputs(302) <= layer4_outputs(2461);
    layer5_outputs(303) <= not(layer4_outputs(1771)) or (layer4_outputs(4266));
    layer5_outputs(304) <= layer4_outputs(2698);
    layer5_outputs(305) <= (layer4_outputs(3506)) and not (layer4_outputs(4036));
    layer5_outputs(306) <= not((layer4_outputs(2123)) and (layer4_outputs(3445)));
    layer5_outputs(307) <= (layer4_outputs(2265)) xor (layer4_outputs(829));
    layer5_outputs(308) <= not(layer4_outputs(5001)) or (layer4_outputs(874));
    layer5_outputs(309) <= (layer4_outputs(3142)) and not (layer4_outputs(4001));
    layer5_outputs(310) <= layer4_outputs(1856);
    layer5_outputs(311) <= (layer4_outputs(2093)) and not (layer4_outputs(2826));
    layer5_outputs(312) <= (layer4_outputs(4223)) xor (layer4_outputs(1992));
    layer5_outputs(313) <= (layer4_outputs(3418)) and not (layer4_outputs(1973));
    layer5_outputs(314) <= not(layer4_outputs(2987)) or (layer4_outputs(2775));
    layer5_outputs(315) <= layer4_outputs(544);
    layer5_outputs(316) <= not(layer4_outputs(3157)) or (layer4_outputs(2349));
    layer5_outputs(317) <= (layer4_outputs(4848)) and not (layer4_outputs(1426));
    layer5_outputs(318) <= (layer4_outputs(3925)) or (layer4_outputs(997));
    layer5_outputs(319) <= not((layer4_outputs(558)) or (layer4_outputs(1782)));
    layer5_outputs(320) <= not((layer4_outputs(1786)) or (layer4_outputs(3702)));
    layer5_outputs(321) <= '1';
    layer5_outputs(322) <= not(layer4_outputs(4246)) or (layer4_outputs(1249));
    layer5_outputs(323) <= not(layer4_outputs(2082)) or (layer4_outputs(868));
    layer5_outputs(324) <= not(layer4_outputs(710)) or (layer4_outputs(4854));
    layer5_outputs(325) <= not(layer4_outputs(3215));
    layer5_outputs(326) <= not(layer4_outputs(236)) or (layer4_outputs(1204));
    layer5_outputs(327) <= not(layer4_outputs(4767));
    layer5_outputs(328) <= not(layer4_outputs(3803));
    layer5_outputs(329) <= not(layer4_outputs(1670));
    layer5_outputs(330) <= (layer4_outputs(2753)) and not (layer4_outputs(4170));
    layer5_outputs(331) <= not(layer4_outputs(4070)) or (layer4_outputs(2351));
    layer5_outputs(332) <= not(layer4_outputs(2126));
    layer5_outputs(333) <= not((layer4_outputs(384)) xor (layer4_outputs(4920)));
    layer5_outputs(334) <= (layer4_outputs(4545)) or (layer4_outputs(4757));
    layer5_outputs(335) <= not((layer4_outputs(602)) and (layer4_outputs(4047)));
    layer5_outputs(336) <= layer4_outputs(2465);
    layer5_outputs(337) <= layer4_outputs(672);
    layer5_outputs(338) <= not((layer4_outputs(4755)) or (layer4_outputs(2251)));
    layer5_outputs(339) <= (layer4_outputs(3701)) and (layer4_outputs(5014));
    layer5_outputs(340) <= (layer4_outputs(3179)) and not (layer4_outputs(2761));
    layer5_outputs(341) <= '1';
    layer5_outputs(342) <= (layer4_outputs(691)) and not (layer4_outputs(3398));
    layer5_outputs(343) <= layer4_outputs(3752);
    layer5_outputs(344) <= not(layer4_outputs(3383));
    layer5_outputs(345) <= not(layer4_outputs(1310));
    layer5_outputs(346) <= (layer4_outputs(578)) and (layer4_outputs(4727));
    layer5_outputs(347) <= not((layer4_outputs(395)) or (layer4_outputs(4053)));
    layer5_outputs(348) <= (layer4_outputs(3570)) xor (layer4_outputs(3150));
    layer5_outputs(349) <= (layer4_outputs(4701)) and not (layer4_outputs(208));
    layer5_outputs(350) <= not(layer4_outputs(675));
    layer5_outputs(351) <= (layer4_outputs(3979)) and not (layer4_outputs(2536));
    layer5_outputs(352) <= not(layer4_outputs(1031));
    layer5_outputs(353) <= layer4_outputs(4458);
    layer5_outputs(354) <= not((layer4_outputs(2372)) xor (layer4_outputs(1788)));
    layer5_outputs(355) <= not(layer4_outputs(1294));
    layer5_outputs(356) <= layer4_outputs(4416);
    layer5_outputs(357) <= not((layer4_outputs(3775)) and (layer4_outputs(3205)));
    layer5_outputs(358) <= layer4_outputs(2035);
    layer5_outputs(359) <= '0';
    layer5_outputs(360) <= layer4_outputs(2469);
    layer5_outputs(361) <= not(layer4_outputs(1956));
    layer5_outputs(362) <= (layer4_outputs(3206)) and not (layer4_outputs(3571));
    layer5_outputs(363) <= not(layer4_outputs(3130)) or (layer4_outputs(28));
    layer5_outputs(364) <= (layer4_outputs(2732)) and not (layer4_outputs(4011));
    layer5_outputs(365) <= layer4_outputs(4843);
    layer5_outputs(366) <= not(layer4_outputs(439));
    layer5_outputs(367) <= '0';
    layer5_outputs(368) <= (layer4_outputs(1081)) xor (layer4_outputs(4990));
    layer5_outputs(369) <= not((layer4_outputs(4437)) xor (layer4_outputs(531)));
    layer5_outputs(370) <= '0';
    layer5_outputs(371) <= layer4_outputs(4447);
    layer5_outputs(372) <= (layer4_outputs(4149)) or (layer4_outputs(3703));
    layer5_outputs(373) <= not(layer4_outputs(2821)) or (layer4_outputs(5034));
    layer5_outputs(374) <= (layer4_outputs(1125)) and not (layer4_outputs(1028));
    layer5_outputs(375) <= layer4_outputs(3104);
    layer5_outputs(376) <= '1';
    layer5_outputs(377) <= (layer4_outputs(1819)) and (layer4_outputs(3194));
    layer5_outputs(378) <= not((layer4_outputs(1423)) or (layer4_outputs(3115)));
    layer5_outputs(379) <= not((layer4_outputs(968)) and (layer4_outputs(4677)));
    layer5_outputs(380) <= not((layer4_outputs(3151)) and (layer4_outputs(3859)));
    layer5_outputs(381) <= layer4_outputs(3882);
    layer5_outputs(382) <= layer4_outputs(1433);
    layer5_outputs(383) <= layer4_outputs(3696);
    layer5_outputs(384) <= not((layer4_outputs(2235)) and (layer4_outputs(2489)));
    layer5_outputs(385) <= layer4_outputs(5008);
    layer5_outputs(386) <= not(layer4_outputs(377));
    layer5_outputs(387) <= '1';
    layer5_outputs(388) <= (layer4_outputs(4959)) and not (layer4_outputs(3420));
    layer5_outputs(389) <= not((layer4_outputs(1036)) or (layer4_outputs(2114)));
    layer5_outputs(390) <= '1';
    layer5_outputs(391) <= layer4_outputs(3954);
    layer5_outputs(392) <= '1';
    layer5_outputs(393) <= not(layer4_outputs(2117));
    layer5_outputs(394) <= (layer4_outputs(4235)) xor (layer4_outputs(1092));
    layer5_outputs(395) <= not((layer4_outputs(545)) or (layer4_outputs(3240)));
    layer5_outputs(396) <= layer4_outputs(3017);
    layer5_outputs(397) <= not(layer4_outputs(4103)) or (layer4_outputs(410));
    layer5_outputs(398) <= not(layer4_outputs(1314));
    layer5_outputs(399) <= not(layer4_outputs(4389)) or (layer4_outputs(3343));
    layer5_outputs(400) <= (layer4_outputs(1689)) and not (layer4_outputs(4412));
    layer5_outputs(401) <= '1';
    layer5_outputs(402) <= not((layer4_outputs(2348)) and (layer4_outputs(3204)));
    layer5_outputs(403) <= '0';
    layer5_outputs(404) <= not(layer4_outputs(4306));
    layer5_outputs(405) <= not(layer4_outputs(3916)) or (layer4_outputs(3195));
    layer5_outputs(406) <= not(layer4_outputs(4160));
    layer5_outputs(407) <= not(layer4_outputs(2392)) or (layer4_outputs(975));
    layer5_outputs(408) <= not((layer4_outputs(3552)) and (layer4_outputs(4117)));
    layer5_outputs(409) <= (layer4_outputs(9)) and (layer4_outputs(4964));
    layer5_outputs(410) <= layer4_outputs(2054);
    layer5_outputs(411) <= (layer4_outputs(1588)) xor (layer4_outputs(4674));
    layer5_outputs(412) <= not(layer4_outputs(2662)) or (layer4_outputs(3730));
    layer5_outputs(413) <= (layer4_outputs(3980)) and (layer4_outputs(3911));
    layer5_outputs(414) <= (layer4_outputs(1333)) and not (layer4_outputs(3330));
    layer5_outputs(415) <= not((layer4_outputs(4735)) and (layer4_outputs(4869)));
    layer5_outputs(416) <= not((layer4_outputs(3879)) and (layer4_outputs(2822)));
    layer5_outputs(417) <= layer4_outputs(3997);
    layer5_outputs(418) <= layer4_outputs(3997);
    layer5_outputs(419) <= not(layer4_outputs(13));
    layer5_outputs(420) <= not(layer4_outputs(1556));
    layer5_outputs(421) <= (layer4_outputs(433)) xor (layer4_outputs(1456));
    layer5_outputs(422) <= (layer4_outputs(3146)) and not (layer4_outputs(181));
    layer5_outputs(423) <= not(layer4_outputs(2014)) or (layer4_outputs(2477));
    layer5_outputs(424) <= (layer4_outputs(1762)) or (layer4_outputs(5033));
    layer5_outputs(425) <= (layer4_outputs(3786)) xor (layer4_outputs(441));
    layer5_outputs(426) <= not((layer4_outputs(2050)) or (layer4_outputs(230)));
    layer5_outputs(427) <= not((layer4_outputs(2843)) or (layer4_outputs(3681)));
    layer5_outputs(428) <= (layer4_outputs(298)) and (layer4_outputs(3296));
    layer5_outputs(429) <= (layer4_outputs(3851)) and not (layer4_outputs(2556));
    layer5_outputs(430) <= not(layer4_outputs(814));
    layer5_outputs(431) <= (layer4_outputs(2980)) and not (layer4_outputs(3036));
    layer5_outputs(432) <= not(layer4_outputs(2691));
    layer5_outputs(433) <= (layer4_outputs(2077)) and not (layer4_outputs(3638));
    layer5_outputs(434) <= (layer4_outputs(3614)) and (layer4_outputs(2530));
    layer5_outputs(435) <= (layer4_outputs(80)) and (layer4_outputs(1211));
    layer5_outputs(436) <= not(layer4_outputs(1558));
    layer5_outputs(437) <= layer4_outputs(2571);
    layer5_outputs(438) <= not(layer4_outputs(974)) or (layer4_outputs(4692));
    layer5_outputs(439) <= layer4_outputs(2362);
    layer5_outputs(440) <= not((layer4_outputs(4736)) or (layer4_outputs(2292)));
    layer5_outputs(441) <= not(layer4_outputs(3602)) or (layer4_outputs(805));
    layer5_outputs(442) <= (layer4_outputs(1487)) or (layer4_outputs(194));
    layer5_outputs(443) <= layer4_outputs(4036);
    layer5_outputs(444) <= layer4_outputs(5083);
    layer5_outputs(445) <= layer4_outputs(3335);
    layer5_outputs(446) <= (layer4_outputs(4197)) and (layer4_outputs(2754));
    layer5_outputs(447) <= '1';
    layer5_outputs(448) <= not(layer4_outputs(2139)) or (layer4_outputs(2517));
    layer5_outputs(449) <= (layer4_outputs(4077)) and not (layer4_outputs(2935));
    layer5_outputs(450) <= not((layer4_outputs(2677)) and (layer4_outputs(4813)));
    layer5_outputs(451) <= '1';
    layer5_outputs(452) <= not(layer4_outputs(1167));
    layer5_outputs(453) <= not(layer4_outputs(3517)) or (layer4_outputs(2330));
    layer5_outputs(454) <= '0';
    layer5_outputs(455) <= not((layer4_outputs(52)) and (layer4_outputs(1949)));
    layer5_outputs(456) <= not(layer4_outputs(2130)) or (layer4_outputs(282));
    layer5_outputs(457) <= not(layer4_outputs(687)) or (layer4_outputs(2603));
    layer5_outputs(458) <= (layer4_outputs(3966)) or (layer4_outputs(5102));
    layer5_outputs(459) <= (layer4_outputs(242)) xor (layer4_outputs(733));
    layer5_outputs(460) <= not(layer4_outputs(1833));
    layer5_outputs(461) <= not(layer4_outputs(4648));
    layer5_outputs(462) <= not(layer4_outputs(834));
    layer5_outputs(463) <= not(layer4_outputs(253));
    layer5_outputs(464) <= (layer4_outputs(4694)) and (layer4_outputs(1207));
    layer5_outputs(465) <= (layer4_outputs(3221)) or (layer4_outputs(3713));
    layer5_outputs(466) <= layer4_outputs(2847);
    layer5_outputs(467) <= (layer4_outputs(2984)) and (layer4_outputs(4418));
    layer5_outputs(468) <= (layer4_outputs(2870)) and (layer4_outputs(290));
    layer5_outputs(469) <= (layer4_outputs(3193)) xor (layer4_outputs(1716));
    layer5_outputs(470) <= layer4_outputs(475);
    layer5_outputs(471) <= not(layer4_outputs(934));
    layer5_outputs(472) <= (layer4_outputs(2882)) xor (layer4_outputs(128));
    layer5_outputs(473) <= (layer4_outputs(1586)) and not (layer4_outputs(902));
    layer5_outputs(474) <= '1';
    layer5_outputs(475) <= not(layer4_outputs(231));
    layer5_outputs(476) <= (layer4_outputs(204)) or (layer4_outputs(1299));
    layer5_outputs(477) <= not(layer4_outputs(5044));
    layer5_outputs(478) <= '1';
    layer5_outputs(479) <= (layer4_outputs(1937)) and (layer4_outputs(3742));
    layer5_outputs(480) <= not(layer4_outputs(882));
    layer5_outputs(481) <= layer4_outputs(2859);
    layer5_outputs(482) <= layer4_outputs(2974);
    layer5_outputs(483) <= not((layer4_outputs(2084)) and (layer4_outputs(3898)));
    layer5_outputs(484) <= not(layer4_outputs(4502));
    layer5_outputs(485) <= not((layer4_outputs(4426)) or (layer4_outputs(668)));
    layer5_outputs(486) <= not((layer4_outputs(4064)) or (layer4_outputs(3500)));
    layer5_outputs(487) <= not(layer4_outputs(3223));
    layer5_outputs(488) <= not(layer4_outputs(1821));
    layer5_outputs(489) <= layer4_outputs(1011);
    layer5_outputs(490) <= (layer4_outputs(240)) and not (layer4_outputs(4703));
    layer5_outputs(491) <= '0';
    layer5_outputs(492) <= not(layer4_outputs(296));
    layer5_outputs(493) <= (layer4_outputs(4278)) and (layer4_outputs(4563));
    layer5_outputs(494) <= '0';
    layer5_outputs(495) <= not(layer4_outputs(2286));
    layer5_outputs(496) <= not((layer4_outputs(255)) and (layer4_outputs(1206)));
    layer5_outputs(497) <= (layer4_outputs(2564)) or (layer4_outputs(2951));
    layer5_outputs(498) <= (layer4_outputs(4572)) and not (layer4_outputs(4731));
    layer5_outputs(499) <= (layer4_outputs(1228)) and (layer4_outputs(2442));
    layer5_outputs(500) <= not(layer4_outputs(3062));
    layer5_outputs(501) <= (layer4_outputs(263)) and (layer4_outputs(1418));
    layer5_outputs(502) <= layer4_outputs(2168);
    layer5_outputs(503) <= not(layer4_outputs(614));
    layer5_outputs(504) <= (layer4_outputs(3292)) and (layer4_outputs(683));
    layer5_outputs(505) <= not(layer4_outputs(3578)) or (layer4_outputs(1915));
    layer5_outputs(506) <= not(layer4_outputs(3767));
    layer5_outputs(507) <= layer4_outputs(704);
    layer5_outputs(508) <= not(layer4_outputs(3070));
    layer5_outputs(509) <= not(layer4_outputs(2915)) or (layer4_outputs(4365));
    layer5_outputs(510) <= not(layer4_outputs(4685));
    layer5_outputs(511) <= (layer4_outputs(2998)) and (layer4_outputs(2436));
    layer5_outputs(512) <= (layer4_outputs(2148)) and not (layer4_outputs(97));
    layer5_outputs(513) <= layer4_outputs(2283);
    layer5_outputs(514) <= not((layer4_outputs(3101)) and (layer4_outputs(5017)));
    layer5_outputs(515) <= (layer4_outputs(2221)) or (layer4_outputs(3459));
    layer5_outputs(516) <= (layer4_outputs(4320)) and not (layer4_outputs(2532));
    layer5_outputs(517) <= not((layer4_outputs(5119)) xor (layer4_outputs(3609)));
    layer5_outputs(518) <= not(layer4_outputs(594));
    layer5_outputs(519) <= (layer4_outputs(725)) xor (layer4_outputs(3983));
    layer5_outputs(520) <= layer4_outputs(144);
    layer5_outputs(521) <= not(layer4_outputs(2454));
    layer5_outputs(522) <= (layer4_outputs(3659)) xor (layer4_outputs(582));
    layer5_outputs(523) <= (layer4_outputs(3414)) and (layer4_outputs(543));
    layer5_outputs(524) <= not(layer4_outputs(1313)) or (layer4_outputs(1290));
    layer5_outputs(525) <= (layer4_outputs(3273)) and not (layer4_outputs(3781));
    layer5_outputs(526) <= layer4_outputs(376);
    layer5_outputs(527) <= layer4_outputs(2629);
    layer5_outputs(528) <= layer4_outputs(1580);
    layer5_outputs(529) <= not(layer4_outputs(2098)) or (layer4_outputs(3640));
    layer5_outputs(530) <= not(layer4_outputs(3661));
    layer5_outputs(531) <= '1';
    layer5_outputs(532) <= layer4_outputs(1233);
    layer5_outputs(533) <= not((layer4_outputs(3990)) or (layer4_outputs(1784)));
    layer5_outputs(534) <= not(layer4_outputs(4005));
    layer5_outputs(535) <= (layer4_outputs(434)) or (layer4_outputs(4438));
    layer5_outputs(536) <= layer4_outputs(4864);
    layer5_outputs(537) <= not((layer4_outputs(3601)) and (layer4_outputs(1880)));
    layer5_outputs(538) <= (layer4_outputs(2063)) and not (layer4_outputs(3668));
    layer5_outputs(539) <= not(layer4_outputs(954));
    layer5_outputs(540) <= (layer4_outputs(2498)) and not (layer4_outputs(3188));
    layer5_outputs(541) <= not((layer4_outputs(987)) or (layer4_outputs(4584)));
    layer5_outputs(542) <= not((layer4_outputs(34)) xor (layer4_outputs(3788)));
    layer5_outputs(543) <= not(layer4_outputs(1525));
    layer5_outputs(544) <= '1';
    layer5_outputs(545) <= not((layer4_outputs(1169)) xor (layer4_outputs(4963)));
    layer5_outputs(546) <= layer4_outputs(831);
    layer5_outputs(547) <= layer4_outputs(1424);
    layer5_outputs(548) <= not(layer4_outputs(4564)) or (layer4_outputs(3721));
    layer5_outputs(549) <= not(layer4_outputs(1397));
    layer5_outputs(550) <= '0';
    layer5_outputs(551) <= (layer4_outputs(3566)) and (layer4_outputs(3589));
    layer5_outputs(552) <= not((layer4_outputs(1832)) or (layer4_outputs(3735)));
    layer5_outputs(553) <= not(layer4_outputs(2627)) or (layer4_outputs(1732));
    layer5_outputs(554) <= not(layer4_outputs(4930)) or (layer4_outputs(3363));
    layer5_outputs(555) <= layer4_outputs(4014);
    layer5_outputs(556) <= not((layer4_outputs(3890)) and (layer4_outputs(4850)));
    layer5_outputs(557) <= not(layer4_outputs(1983)) or (layer4_outputs(292));
    layer5_outputs(558) <= layer4_outputs(371);
    layer5_outputs(559) <= '1';
    layer5_outputs(560) <= not(layer4_outputs(2705)) or (layer4_outputs(1644));
    layer5_outputs(561) <= not(layer4_outputs(852));
    layer5_outputs(562) <= '1';
    layer5_outputs(563) <= not((layer4_outputs(513)) or (layer4_outputs(2647)));
    layer5_outputs(564) <= (layer4_outputs(2270)) or (layer4_outputs(2946));
    layer5_outputs(565) <= not(layer4_outputs(3146)) or (layer4_outputs(3981));
    layer5_outputs(566) <= not(layer4_outputs(2120));
    layer5_outputs(567) <= '1';
    layer5_outputs(568) <= (layer4_outputs(3185)) or (layer4_outputs(910));
    layer5_outputs(569) <= not(layer4_outputs(849));
    layer5_outputs(570) <= layer4_outputs(2069);
    layer5_outputs(571) <= layer4_outputs(3651);
    layer5_outputs(572) <= layer4_outputs(4157);
    layer5_outputs(573) <= (layer4_outputs(1719)) and (layer4_outputs(2720));
    layer5_outputs(574) <= (layer4_outputs(3539)) and (layer4_outputs(2296));
    layer5_outputs(575) <= layer4_outputs(2022);
    layer5_outputs(576) <= not(layer4_outputs(2374)) or (layer4_outputs(331));
    layer5_outputs(577) <= (layer4_outputs(762)) or (layer4_outputs(3930));
    layer5_outputs(578) <= not((layer4_outputs(2071)) and (layer4_outputs(967)));
    layer5_outputs(579) <= not(layer4_outputs(1617));
    layer5_outputs(580) <= not(layer4_outputs(360));
    layer5_outputs(581) <= (layer4_outputs(2826)) or (layer4_outputs(1219));
    layer5_outputs(582) <= not(layer4_outputs(3634));
    layer5_outputs(583) <= (layer4_outputs(1388)) or (layer4_outputs(59));
    layer5_outputs(584) <= '0';
    layer5_outputs(585) <= not((layer4_outputs(2395)) and (layer4_outputs(4811)));
    layer5_outputs(586) <= (layer4_outputs(2182)) and not (layer4_outputs(4296));
    layer5_outputs(587) <= (layer4_outputs(1157)) and not (layer4_outputs(3354));
    layer5_outputs(588) <= not(layer4_outputs(2491)) or (layer4_outputs(2862));
    layer5_outputs(589) <= not((layer4_outputs(1761)) or (layer4_outputs(2230)));
    layer5_outputs(590) <= (layer4_outputs(3724)) and (layer4_outputs(2784));
    layer5_outputs(591) <= (layer4_outputs(957)) or (layer4_outputs(1870));
    layer5_outputs(592) <= not(layer4_outputs(2243));
    layer5_outputs(593) <= '1';
    layer5_outputs(594) <= (layer4_outputs(1595)) and (layer4_outputs(2765));
    layer5_outputs(595) <= layer4_outputs(3436);
    layer5_outputs(596) <= (layer4_outputs(1350)) or (layer4_outputs(2151));
    layer5_outputs(597) <= not(layer4_outputs(1579)) or (layer4_outputs(3611));
    layer5_outputs(598) <= (layer4_outputs(4046)) and not (layer4_outputs(356));
    layer5_outputs(599) <= not(layer4_outputs(4949)) or (layer4_outputs(1823));
    layer5_outputs(600) <= (layer4_outputs(877)) and not (layer4_outputs(4056));
    layer5_outputs(601) <= layer4_outputs(3953);
    layer5_outputs(602) <= not(layer4_outputs(1825)) or (layer4_outputs(1736));
    layer5_outputs(603) <= (layer4_outputs(1943)) and (layer4_outputs(824));
    layer5_outputs(604) <= not((layer4_outputs(2750)) and (layer4_outputs(3579)));
    layer5_outputs(605) <= (layer4_outputs(3401)) and not (layer4_outputs(3165));
    layer5_outputs(606) <= not(layer4_outputs(4891));
    layer5_outputs(607) <= '1';
    layer5_outputs(608) <= not(layer4_outputs(588)) or (layer4_outputs(2979));
    layer5_outputs(609) <= (layer4_outputs(5015)) and (layer4_outputs(4662));
    layer5_outputs(610) <= '1';
    layer5_outputs(611) <= not(layer4_outputs(1281)) or (layer4_outputs(4444));
    layer5_outputs(612) <= layer4_outputs(3206);
    layer5_outputs(613) <= not(layer4_outputs(3491)) or (layer4_outputs(3231));
    layer5_outputs(614) <= not((layer4_outputs(2551)) or (layer4_outputs(1475)));
    layer5_outputs(615) <= '0';
    layer5_outputs(616) <= (layer4_outputs(396)) and not (layer4_outputs(33));
    layer5_outputs(617) <= layer4_outputs(2147);
    layer5_outputs(618) <= layer4_outputs(715);
    layer5_outputs(619) <= layer4_outputs(2592);
    layer5_outputs(620) <= not(layer4_outputs(992)) or (layer4_outputs(4710));
    layer5_outputs(621) <= not(layer4_outputs(2568));
    layer5_outputs(622) <= not((layer4_outputs(4841)) and (layer4_outputs(2687)));
    layer5_outputs(623) <= layer4_outputs(4066);
    layer5_outputs(624) <= layer4_outputs(4567);
    layer5_outputs(625) <= not(layer4_outputs(1235));
    layer5_outputs(626) <= not((layer4_outputs(956)) and (layer4_outputs(1770)));
    layer5_outputs(627) <= (layer4_outputs(1173)) and (layer4_outputs(4679));
    layer5_outputs(628) <= not(layer4_outputs(342));
    layer5_outputs(629) <= (layer4_outputs(4511)) and not (layer4_outputs(4388));
    layer5_outputs(630) <= not((layer4_outputs(2635)) and (layer4_outputs(4300)));
    layer5_outputs(631) <= layer4_outputs(3814);
    layer5_outputs(632) <= (layer4_outputs(3469)) xor (layer4_outputs(2446));
    layer5_outputs(633) <= layer4_outputs(3753);
    layer5_outputs(634) <= (layer4_outputs(5007)) or (layer4_outputs(1243));
    layer5_outputs(635) <= (layer4_outputs(15)) and (layer4_outputs(653));
    layer5_outputs(636) <= layer4_outputs(3023);
    layer5_outputs(637) <= not(layer4_outputs(3687));
    layer5_outputs(638) <= layer4_outputs(754);
    layer5_outputs(639) <= not(layer4_outputs(4162)) or (layer4_outputs(4212));
    layer5_outputs(640) <= layer4_outputs(4933);
    layer5_outputs(641) <= layer4_outputs(689);
    layer5_outputs(642) <= layer4_outputs(640);
    layer5_outputs(643) <= not(layer4_outputs(1245));
    layer5_outputs(644) <= not((layer4_outputs(4084)) and (layer4_outputs(4696)));
    layer5_outputs(645) <= (layer4_outputs(856)) and not (layer4_outputs(3210));
    layer5_outputs(646) <= not((layer4_outputs(1640)) or (layer4_outputs(4336)));
    layer5_outputs(647) <= not(layer4_outputs(2813));
    layer5_outputs(648) <= layer4_outputs(2057);
    layer5_outputs(649) <= '0';
    layer5_outputs(650) <= not(layer4_outputs(1125)) or (layer4_outputs(4255));
    layer5_outputs(651) <= layer4_outputs(3476);
    layer5_outputs(652) <= not(layer4_outputs(3077));
    layer5_outputs(653) <= (layer4_outputs(2611)) xor (layer4_outputs(5115));
    layer5_outputs(654) <= (layer4_outputs(4584)) xor (layer4_outputs(1650));
    layer5_outputs(655) <= not((layer4_outputs(3220)) xor (layer4_outputs(8)));
    layer5_outputs(656) <= not(layer4_outputs(3604));
    layer5_outputs(657) <= not(layer4_outputs(3826)) or (layer4_outputs(4196));
    layer5_outputs(658) <= layer4_outputs(3693);
    layer5_outputs(659) <= (layer4_outputs(1344)) xor (layer4_outputs(4473));
    layer5_outputs(660) <= not(layer4_outputs(4828)) or (layer4_outputs(1349));
    layer5_outputs(661) <= (layer4_outputs(241)) or (layer4_outputs(4762));
    layer5_outputs(662) <= not((layer4_outputs(3800)) or (layer4_outputs(2879)));
    layer5_outputs(663) <= not(layer4_outputs(4893));
    layer5_outputs(664) <= '1';
    layer5_outputs(665) <= not(layer4_outputs(3365));
    layer5_outputs(666) <= layer4_outputs(4792);
    layer5_outputs(667) <= (layer4_outputs(1137)) and not (layer4_outputs(3407));
    layer5_outputs(668) <= not((layer4_outputs(1325)) and (layer4_outputs(2945)));
    layer5_outputs(669) <= not(layer4_outputs(2279));
    layer5_outputs(670) <= '1';
    layer5_outputs(671) <= layer4_outputs(1357);
    layer5_outputs(672) <= layer4_outputs(612);
    layer5_outputs(673) <= not(layer4_outputs(1721)) or (layer4_outputs(986));
    layer5_outputs(674) <= not(layer4_outputs(806));
    layer5_outputs(675) <= (layer4_outputs(3367)) or (layer4_outputs(2053));
    layer5_outputs(676) <= not(layer4_outputs(1384));
    layer5_outputs(677) <= not(layer4_outputs(3451));
    layer5_outputs(678) <= not(layer4_outputs(2523));
    layer5_outputs(679) <= (layer4_outputs(229)) xor (layer4_outputs(3685));
    layer5_outputs(680) <= (layer4_outputs(2713)) or (layer4_outputs(1687));
    layer5_outputs(681) <= not(layer4_outputs(4877));
    layer5_outputs(682) <= not(layer4_outputs(3153));
    layer5_outputs(683) <= layer4_outputs(3902);
    layer5_outputs(684) <= (layer4_outputs(2837)) or (layer4_outputs(1082));
    layer5_outputs(685) <= not((layer4_outputs(2594)) or (layer4_outputs(3190)));
    layer5_outputs(686) <= not(layer4_outputs(698));
    layer5_outputs(687) <= not(layer4_outputs(1089));
    layer5_outputs(688) <= not(layer4_outputs(1540)) or (layer4_outputs(4644));
    layer5_outputs(689) <= not(layer4_outputs(3462));
    layer5_outputs(690) <= '1';
    layer5_outputs(691) <= not((layer4_outputs(1514)) and (layer4_outputs(2954)));
    layer5_outputs(692) <= not(layer4_outputs(1486));
    layer5_outputs(693) <= (layer4_outputs(688)) or (layer4_outputs(1530));
    layer5_outputs(694) <= not(layer4_outputs(3995)) or (layer4_outputs(4791));
    layer5_outputs(695) <= (layer4_outputs(1501)) and (layer4_outputs(900));
    layer5_outputs(696) <= not(layer4_outputs(214)) or (layer4_outputs(207));
    layer5_outputs(697) <= (layer4_outputs(4637)) and not (layer4_outputs(5));
    layer5_outputs(698) <= (layer4_outputs(2577)) xor (layer4_outputs(3221));
    layer5_outputs(699) <= (layer4_outputs(4969)) or (layer4_outputs(2698));
    layer5_outputs(700) <= layer4_outputs(297);
    layer5_outputs(701) <= not((layer4_outputs(4406)) xor (layer4_outputs(3228)));
    layer5_outputs(702) <= not(layer4_outputs(2736));
    layer5_outputs(703) <= layer4_outputs(216);
    layer5_outputs(704) <= not(layer4_outputs(2666));
    layer5_outputs(705) <= layer4_outputs(3714);
    layer5_outputs(706) <= layer4_outputs(4907);
    layer5_outputs(707) <= '0';
    layer5_outputs(708) <= (layer4_outputs(2762)) xor (layer4_outputs(529));
    layer5_outputs(709) <= (layer4_outputs(1003)) and not (layer4_outputs(2502));
    layer5_outputs(710) <= not(layer4_outputs(4585));
    layer5_outputs(711) <= layer4_outputs(3041);
    layer5_outputs(712) <= (layer4_outputs(2593)) and (layer4_outputs(1155));
    layer5_outputs(713) <= (layer4_outputs(3448)) xor (layer4_outputs(3601));
    layer5_outputs(714) <= (layer4_outputs(3977)) and not (layer4_outputs(4864));
    layer5_outputs(715) <= layer4_outputs(4066);
    layer5_outputs(716) <= (layer4_outputs(1866)) and not (layer4_outputs(1196));
    layer5_outputs(717) <= (layer4_outputs(4023)) and not (layer4_outputs(4484));
    layer5_outputs(718) <= (layer4_outputs(3685)) and not (layer4_outputs(3483));
    layer5_outputs(719) <= (layer4_outputs(1710)) or (layer4_outputs(3865));
    layer5_outputs(720) <= '1';
    layer5_outputs(721) <= (layer4_outputs(3474)) and not (layer4_outputs(3678));
    layer5_outputs(722) <= layer4_outputs(2181);
    layer5_outputs(723) <= not(layer4_outputs(1446));
    layer5_outputs(724) <= (layer4_outputs(5030)) and not (layer4_outputs(5004));
    layer5_outputs(725) <= not(layer4_outputs(2306)) or (layer4_outputs(1895));
    layer5_outputs(726) <= layer4_outputs(2735);
    layer5_outputs(727) <= layer4_outputs(1545);
    layer5_outputs(728) <= not((layer4_outputs(3946)) xor (layer4_outputs(4124)));
    layer5_outputs(729) <= layer4_outputs(220);
    layer5_outputs(730) <= '0';
    layer5_outputs(731) <= (layer4_outputs(1192)) or (layer4_outputs(4616));
    layer5_outputs(732) <= not(layer4_outputs(4322)) or (layer4_outputs(2937));
    layer5_outputs(733) <= not(layer4_outputs(2681));
    layer5_outputs(734) <= not((layer4_outputs(3523)) and (layer4_outputs(2928)));
    layer5_outputs(735) <= not(layer4_outputs(1083));
    layer5_outputs(736) <= (layer4_outputs(4558)) or (layer4_outputs(3812));
    layer5_outputs(737) <= not(layer4_outputs(3852));
    layer5_outputs(738) <= (layer4_outputs(4400)) and not (layer4_outputs(1095));
    layer5_outputs(739) <= not(layer4_outputs(2337));
    layer5_outputs(740) <= (layer4_outputs(1997)) and not (layer4_outputs(2424));
    layer5_outputs(741) <= not(layer4_outputs(4161)) or (layer4_outputs(38));
    layer5_outputs(742) <= not(layer4_outputs(3058)) or (layer4_outputs(4796));
    layer5_outputs(743) <= (layer4_outputs(3509)) or (layer4_outputs(1801));
    layer5_outputs(744) <= not(layer4_outputs(4843));
    layer5_outputs(745) <= not(layer4_outputs(5096)) or (layer4_outputs(389));
    layer5_outputs(746) <= not(layer4_outputs(409));
    layer5_outputs(747) <= layer4_outputs(3351);
    layer5_outputs(748) <= '1';
    layer5_outputs(749) <= layer4_outputs(1915);
    layer5_outputs(750) <= not(layer4_outputs(348));
    layer5_outputs(751) <= layer4_outputs(1643);
    layer5_outputs(752) <= not(layer4_outputs(4488));
    layer5_outputs(753) <= (layer4_outputs(3847)) xor (layer4_outputs(4726));
    layer5_outputs(754) <= not(layer4_outputs(3224));
    layer5_outputs(755) <= '0';
    layer5_outputs(756) <= not(layer4_outputs(3124));
    layer5_outputs(757) <= '1';
    layer5_outputs(758) <= not(layer4_outputs(4019));
    layer5_outputs(759) <= '0';
    layer5_outputs(760) <= (layer4_outputs(4701)) and not (layer4_outputs(4116));
    layer5_outputs(761) <= not((layer4_outputs(472)) and (layer4_outputs(4508)));
    layer5_outputs(762) <= layer4_outputs(2028);
    layer5_outputs(763) <= (layer4_outputs(2619)) and not (layer4_outputs(1888));
    layer5_outputs(764) <= '1';
    layer5_outputs(765) <= not((layer4_outputs(2042)) and (layer4_outputs(1875)));
    layer5_outputs(766) <= not(layer4_outputs(3289)) or (layer4_outputs(1671));
    layer5_outputs(767) <= not(layer4_outputs(1054));
    layer5_outputs(768) <= layer4_outputs(3694);
    layer5_outputs(769) <= (layer4_outputs(4926)) and (layer4_outputs(2534));
    layer5_outputs(770) <= layer4_outputs(1559);
    layer5_outputs(771) <= '1';
    layer5_outputs(772) <= layer4_outputs(77);
    layer5_outputs(773) <= not(layer4_outputs(731));
    layer5_outputs(774) <= layer4_outputs(741);
    layer5_outputs(775) <= not((layer4_outputs(4199)) xor (layer4_outputs(3449)));
    layer5_outputs(776) <= (layer4_outputs(703)) and (layer4_outputs(3279));
    layer5_outputs(777) <= not((layer4_outputs(915)) or (layer4_outputs(4509)));
    layer5_outputs(778) <= not((layer4_outputs(1339)) and (layer4_outputs(3677)));
    layer5_outputs(779) <= layer4_outputs(4759);
    layer5_outputs(780) <= not((layer4_outputs(225)) or (layer4_outputs(3035)));
    layer5_outputs(781) <= not(layer4_outputs(549)) or (layer4_outputs(2520));
    layer5_outputs(782) <= layer4_outputs(4628);
    layer5_outputs(783) <= not(layer4_outputs(3781));
    layer5_outputs(784) <= '1';
    layer5_outputs(785) <= (layer4_outputs(3686)) and not (layer4_outputs(817));
    layer5_outputs(786) <= (layer4_outputs(2085)) xor (layer4_outputs(1359));
    layer5_outputs(787) <= layer4_outputs(4018);
    layer5_outputs(788) <= (layer4_outputs(1370)) and not (layer4_outputs(4166));
    layer5_outputs(789) <= not(layer4_outputs(3369));
    layer5_outputs(790) <= not(layer4_outputs(519)) or (layer4_outputs(544));
    layer5_outputs(791) <= layer4_outputs(2803);
    layer5_outputs(792) <= (layer4_outputs(1571)) and (layer4_outputs(1827));
    layer5_outputs(793) <= layer4_outputs(4487);
    layer5_outputs(794) <= (layer4_outputs(827)) or (layer4_outputs(434));
    layer5_outputs(795) <= (layer4_outputs(999)) and (layer4_outputs(2263));
    layer5_outputs(796) <= not((layer4_outputs(3463)) xor (layer4_outputs(601)));
    layer5_outputs(797) <= not(layer4_outputs(2424));
    layer5_outputs(798) <= not(layer4_outputs(3407));
    layer5_outputs(799) <= not((layer4_outputs(1318)) xor (layer4_outputs(2892)));
    layer5_outputs(800) <= '0';
    layer5_outputs(801) <= (layer4_outputs(1366)) xor (layer4_outputs(4512));
    layer5_outputs(802) <= not((layer4_outputs(1920)) and (layer4_outputs(1760)));
    layer5_outputs(803) <= (layer4_outputs(2945)) and not (layer4_outputs(4754));
    layer5_outputs(804) <= (layer4_outputs(2630)) and not (layer4_outputs(609));
    layer5_outputs(805) <= layer4_outputs(3627);
    layer5_outputs(806) <= not(layer4_outputs(3915));
    layer5_outputs(807) <= not((layer4_outputs(1086)) and (layer4_outputs(4834)));
    layer5_outputs(808) <= layer4_outputs(1651);
    layer5_outputs(809) <= layer4_outputs(2719);
    layer5_outputs(810) <= not((layer4_outputs(2544)) and (layer4_outputs(936)));
    layer5_outputs(811) <= not(layer4_outputs(4780)) or (layer4_outputs(844));
    layer5_outputs(812) <= not(layer4_outputs(4676)) or (layer4_outputs(2271));
    layer5_outputs(813) <= not(layer4_outputs(985)) or (layer4_outputs(743));
    layer5_outputs(814) <= not((layer4_outputs(4405)) xor (layer4_outputs(2600)));
    layer5_outputs(815) <= not(layer4_outputs(4110));
    layer5_outputs(816) <= not(layer4_outputs(3604)) or (layer4_outputs(4498));
    layer5_outputs(817) <= not(layer4_outputs(16));
    layer5_outputs(818) <= layer4_outputs(1793);
    layer5_outputs(819) <= not(layer4_outputs(1698));
    layer5_outputs(820) <= not((layer4_outputs(1094)) or (layer4_outputs(2656)));
    layer5_outputs(821) <= not(layer4_outputs(3121));
    layer5_outputs(822) <= not(layer4_outputs(2721));
    layer5_outputs(823) <= (layer4_outputs(4806)) and not (layer4_outputs(1256));
    layer5_outputs(824) <= not(layer4_outputs(1176)) or (layer4_outputs(4033));
    layer5_outputs(825) <= (layer4_outputs(154)) or (layer4_outputs(2641));
    layer5_outputs(826) <= layer4_outputs(388);
    layer5_outputs(827) <= not(layer4_outputs(1824));
    layer5_outputs(828) <= not((layer4_outputs(3760)) or (layer4_outputs(1000)));
    layer5_outputs(829) <= not(layer4_outputs(4169)) or (layer4_outputs(4112));
    layer5_outputs(830) <= not((layer4_outputs(2567)) and (layer4_outputs(73)));
    layer5_outputs(831) <= not((layer4_outputs(486)) or (layer4_outputs(2479)));
    layer5_outputs(832) <= (layer4_outputs(2906)) and not (layer4_outputs(421));
    layer5_outputs(833) <= not((layer4_outputs(2305)) and (layer4_outputs(1130)));
    layer5_outputs(834) <= '0';
    layer5_outputs(835) <= '1';
    layer5_outputs(836) <= layer4_outputs(4614);
    layer5_outputs(837) <= (layer4_outputs(1925)) and (layer4_outputs(1257));
    layer5_outputs(838) <= (layer4_outputs(4304)) or (layer4_outputs(3894));
    layer5_outputs(839) <= layer4_outputs(1234);
    layer5_outputs(840) <= (layer4_outputs(937)) and not (layer4_outputs(2872));
    layer5_outputs(841) <= (layer4_outputs(5041)) and not (layer4_outputs(3178));
    layer5_outputs(842) <= not(layer4_outputs(1700)) or (layer4_outputs(2327));
    layer5_outputs(843) <= layer4_outputs(4466);
    layer5_outputs(844) <= not((layer4_outputs(1669)) and (layer4_outputs(3247)));
    layer5_outputs(845) <= (layer4_outputs(1963)) and not (layer4_outputs(5055));
    layer5_outputs(846) <= (layer4_outputs(3030)) and not (layer4_outputs(2434));
    layer5_outputs(847) <= layer4_outputs(2311);
    layer5_outputs(848) <= (layer4_outputs(5046)) or (layer4_outputs(3387));
    layer5_outputs(849) <= layer4_outputs(2302);
    layer5_outputs(850) <= (layer4_outputs(4080)) and not (layer4_outputs(4034));
    layer5_outputs(851) <= not(layer4_outputs(3125));
    layer5_outputs(852) <= not((layer4_outputs(3008)) or (layer4_outputs(27)));
    layer5_outputs(853) <= (layer4_outputs(4747)) or (layer4_outputs(3022));
    layer5_outputs(854) <= layer4_outputs(117);
    layer5_outputs(855) <= not(layer4_outputs(1739));
    layer5_outputs(856) <= layer4_outputs(1467);
    layer5_outputs(857) <= layer4_outputs(4179);
    layer5_outputs(858) <= not((layer4_outputs(2652)) xor (layer4_outputs(4910)));
    layer5_outputs(859) <= not(layer4_outputs(2585));
    layer5_outputs(860) <= not(layer4_outputs(5070)) or (layer4_outputs(4079));
    layer5_outputs(861) <= not((layer4_outputs(4801)) and (layer4_outputs(2277)));
    layer5_outputs(862) <= layer4_outputs(519);
    layer5_outputs(863) <= not(layer4_outputs(1841));
    layer5_outputs(864) <= (layer4_outputs(401)) and (layer4_outputs(4307));
    layer5_outputs(865) <= layer4_outputs(370);
    layer5_outputs(866) <= '1';
    layer5_outputs(867) <= not(layer4_outputs(364)) or (layer4_outputs(2894));
    layer5_outputs(868) <= not(layer4_outputs(4195));
    layer5_outputs(869) <= not(layer4_outputs(3644)) or (layer4_outputs(336));
    layer5_outputs(870) <= '0';
    layer5_outputs(871) <= (layer4_outputs(1794)) and not (layer4_outputs(3955));
    layer5_outputs(872) <= layer4_outputs(2214);
    layer5_outputs(873) <= '1';
    layer5_outputs(874) <= not((layer4_outputs(4551)) xor (layer4_outputs(4817)));
    layer5_outputs(875) <= layer4_outputs(4183);
    layer5_outputs(876) <= not(layer4_outputs(4328)) or (layer4_outputs(2804));
    layer5_outputs(877) <= layer4_outputs(4889);
    layer5_outputs(878) <= (layer4_outputs(313)) xor (layer4_outputs(696));
    layer5_outputs(879) <= (layer4_outputs(23)) and not (layer4_outputs(259));
    layer5_outputs(880) <= '1';
    layer5_outputs(881) <= not(layer4_outputs(618)) or (layer4_outputs(1436));
    layer5_outputs(882) <= layer4_outputs(1163);
    layer5_outputs(883) <= (layer4_outputs(4057)) xor (layer4_outputs(1914));
    layer5_outputs(884) <= not(layer4_outputs(2088));
    layer5_outputs(885) <= layer4_outputs(4966);
    layer5_outputs(886) <= (layer4_outputs(2343)) or (layer4_outputs(1304));
    layer5_outputs(887) <= not(layer4_outputs(893)) or (layer4_outputs(552));
    layer5_outputs(888) <= layer4_outputs(194);
    layer5_outputs(889) <= not((layer4_outputs(4226)) or (layer4_outputs(2983)));
    layer5_outputs(890) <= (layer4_outputs(3442)) and not (layer4_outputs(4217));
    layer5_outputs(891) <= layer4_outputs(1966);
    layer5_outputs(892) <= not(layer4_outputs(3679)) or (layer4_outputs(232));
    layer5_outputs(893) <= not((layer4_outputs(1156)) and (layer4_outputs(4007)));
    layer5_outputs(894) <= (layer4_outputs(3334)) and (layer4_outputs(4941));
    layer5_outputs(895) <= not((layer4_outputs(2219)) or (layer4_outputs(3597)));
    layer5_outputs(896) <= not(layer4_outputs(1075));
    layer5_outputs(897) <= (layer4_outputs(3802)) and not (layer4_outputs(4067));
    layer5_outputs(898) <= '0';
    layer5_outputs(899) <= (layer4_outputs(4622)) and not (layer4_outputs(3670));
    layer5_outputs(900) <= (layer4_outputs(4941)) and not (layer4_outputs(3214));
    layer5_outputs(901) <= '0';
    layer5_outputs(902) <= (layer4_outputs(2492)) and not (layer4_outputs(1554));
    layer5_outputs(903) <= (layer4_outputs(2116)) or (layer4_outputs(4444));
    layer5_outputs(904) <= layer4_outputs(2384);
    layer5_outputs(905) <= layer4_outputs(297);
    layer5_outputs(906) <= (layer4_outputs(2624)) and (layer4_outputs(2799));
    layer5_outputs(907) <= layer4_outputs(5112);
    layer5_outputs(908) <= not((layer4_outputs(4522)) and (layer4_outputs(2710)));
    layer5_outputs(909) <= (layer4_outputs(2414)) and not (layer4_outputs(2296));
    layer5_outputs(910) <= not(layer4_outputs(1481));
    layer5_outputs(911) <= layer4_outputs(4318);
    layer5_outputs(912) <= '0';
    layer5_outputs(913) <= not(layer4_outputs(502));
    layer5_outputs(914) <= (layer4_outputs(484)) and (layer4_outputs(606));
    layer5_outputs(915) <= layer4_outputs(3283);
    layer5_outputs(916) <= layer4_outputs(5061);
    layer5_outputs(917) <= not(layer4_outputs(881));
    layer5_outputs(918) <= not(layer4_outputs(4836));
    layer5_outputs(919) <= (layer4_outputs(973)) and (layer4_outputs(4582));
    layer5_outputs(920) <= (layer4_outputs(2960)) or (layer4_outputs(4326));
    layer5_outputs(921) <= not(layer4_outputs(4312)) or (layer4_outputs(5018));
    layer5_outputs(922) <= not((layer4_outputs(3542)) or (layer4_outputs(1455)));
    layer5_outputs(923) <= not(layer4_outputs(1015)) or (layer4_outputs(1721));
    layer5_outputs(924) <= not(layer4_outputs(1870));
    layer5_outputs(925) <= not((layer4_outputs(1102)) or (layer4_outputs(4261)));
    layer5_outputs(926) <= not(layer4_outputs(1641)) or (layer4_outputs(3663));
    layer5_outputs(927) <= not(layer4_outputs(4075)) or (layer4_outputs(4548));
    layer5_outputs(928) <= not(layer4_outputs(4363));
    layer5_outputs(929) <= not(layer4_outputs(2690)) or (layer4_outputs(2320));
    layer5_outputs(930) <= layer4_outputs(1926);
    layer5_outputs(931) <= not(layer4_outputs(3763));
    layer5_outputs(932) <= not(layer4_outputs(3117)) or (layer4_outputs(3737));
    layer5_outputs(933) <= (layer4_outputs(482)) and not (layer4_outputs(584));
    layer5_outputs(934) <= layer4_outputs(2765);
    layer5_outputs(935) <= not((layer4_outputs(2658)) and (layer4_outputs(2624)));
    layer5_outputs(936) <= (layer4_outputs(3404)) xor (layer4_outputs(4025));
    layer5_outputs(937) <= (layer4_outputs(3423)) xor (layer4_outputs(4773));
    layer5_outputs(938) <= not((layer4_outputs(593)) and (layer4_outputs(3289)));
    layer5_outputs(939) <= '1';
    layer5_outputs(940) <= '1';
    layer5_outputs(941) <= '1';
    layer5_outputs(942) <= (layer4_outputs(4935)) xor (layer4_outputs(3959));
    layer5_outputs(943) <= not(layer4_outputs(3111));
    layer5_outputs(944) <= layer4_outputs(1822);
    layer5_outputs(945) <= (layer4_outputs(5006)) or (layer4_outputs(93));
    layer5_outputs(946) <= (layer4_outputs(649)) or (layer4_outputs(4868));
    layer5_outputs(947) <= (layer4_outputs(121)) and not (layer4_outputs(392));
    layer5_outputs(948) <= not(layer4_outputs(2755));
    layer5_outputs(949) <= (layer4_outputs(693)) xor (layer4_outputs(2015));
    layer5_outputs(950) <= not(layer4_outputs(3943));
    layer5_outputs(951) <= layer4_outputs(3216);
    layer5_outputs(952) <= not(layer4_outputs(2414));
    layer5_outputs(953) <= (layer4_outputs(1116)) and (layer4_outputs(2760));
    layer5_outputs(954) <= (layer4_outputs(1798)) and (layer4_outputs(435));
    layer5_outputs(955) <= (layer4_outputs(3066)) and (layer4_outputs(4374));
    layer5_outputs(956) <= not(layer4_outputs(1812)) or (layer4_outputs(4380));
    layer5_outputs(957) <= not(layer4_outputs(3083));
    layer5_outputs(958) <= layer4_outputs(1189);
    layer5_outputs(959) <= layer4_outputs(4113);
    layer5_outputs(960) <= (layer4_outputs(3297)) and (layer4_outputs(3536));
    layer5_outputs(961) <= (layer4_outputs(4621)) and not (layer4_outputs(4503));
    layer5_outputs(962) <= layer4_outputs(334);
    layer5_outputs(963) <= not(layer4_outputs(5014)) or (layer4_outputs(2537));
    layer5_outputs(964) <= not(layer4_outputs(783)) or (layer4_outputs(2617));
    layer5_outputs(965) <= (layer4_outputs(3553)) or (layer4_outputs(1685));
    layer5_outputs(966) <= not(layer4_outputs(343)) or (layer4_outputs(414));
    layer5_outputs(967) <= not(layer4_outputs(2508));
    layer5_outputs(968) <= not((layer4_outputs(4234)) or (layer4_outputs(1060)));
    layer5_outputs(969) <= layer4_outputs(4379);
    layer5_outputs(970) <= not(layer4_outputs(2702));
    layer5_outputs(971) <= (layer4_outputs(1153)) and not (layer4_outputs(1183));
    layer5_outputs(972) <= layer4_outputs(4293);
    layer5_outputs(973) <= (layer4_outputs(4951)) and not (layer4_outputs(886));
    layer5_outputs(974) <= not(layer4_outputs(1936));
    layer5_outputs(975) <= not((layer4_outputs(4986)) xor (layer4_outputs(549)));
    layer5_outputs(976) <= (layer4_outputs(1774)) or (layer4_outputs(3719));
    layer5_outputs(977) <= not(layer4_outputs(3921)) or (layer4_outputs(1132));
    layer5_outputs(978) <= (layer4_outputs(3610)) xor (layer4_outputs(2715));
    layer5_outputs(979) <= (layer4_outputs(788)) and not (layer4_outputs(2650));
    layer5_outputs(980) <= not((layer4_outputs(1878)) or (layer4_outputs(3468)));
    layer5_outputs(981) <= not(layer4_outputs(1779));
    layer5_outputs(982) <= not((layer4_outputs(971)) xor (layer4_outputs(4898)));
    layer5_outputs(983) <= not(layer4_outputs(3920)) or (layer4_outputs(5038));
    layer5_outputs(984) <= (layer4_outputs(1894)) and not (layer4_outputs(818));
    layer5_outputs(985) <= not(layer4_outputs(3499));
    layer5_outputs(986) <= not(layer4_outputs(3459)) or (layer4_outputs(2008));
    layer5_outputs(987) <= (layer4_outputs(2817)) and (layer4_outputs(2800));
    layer5_outputs(988) <= not(layer4_outputs(1093));
    layer5_outputs(989) <= layer4_outputs(2217);
    layer5_outputs(990) <= (layer4_outputs(2893)) and not (layer4_outputs(2047));
    layer5_outputs(991) <= layer4_outputs(2852);
    layer5_outputs(992) <= (layer4_outputs(723)) and (layer4_outputs(4940));
    layer5_outputs(993) <= not(layer4_outputs(3831));
    layer5_outputs(994) <= not(layer4_outputs(4805));
    layer5_outputs(995) <= layer4_outputs(349);
    layer5_outputs(996) <= (layer4_outputs(3357)) and not (layer4_outputs(3462));
    layer5_outputs(997) <= (layer4_outputs(2639)) xor (layer4_outputs(2828));
    layer5_outputs(998) <= not((layer4_outputs(3393)) xor (layer4_outputs(302)));
    layer5_outputs(999) <= '1';
    layer5_outputs(1000) <= not((layer4_outputs(2776)) xor (layer4_outputs(3667)));
    layer5_outputs(1001) <= (layer4_outputs(2910)) or (layer4_outputs(4033));
    layer5_outputs(1002) <= (layer4_outputs(1120)) xor (layer4_outputs(652));
    layer5_outputs(1003) <= layer4_outputs(1425);
    layer5_outputs(1004) <= not((layer4_outputs(3929)) and (layer4_outputs(2835)));
    layer5_outputs(1005) <= layer4_outputs(2061);
    layer5_outputs(1006) <= not((layer4_outputs(3273)) or (layer4_outputs(1809)));
    layer5_outputs(1007) <= '0';
    layer5_outputs(1008) <= not((layer4_outputs(4392)) or (layer4_outputs(2132)));
    layer5_outputs(1009) <= not(layer4_outputs(380)) or (layer4_outputs(2309));
    layer5_outputs(1010) <= not((layer4_outputs(4164)) or (layer4_outputs(1232)));
    layer5_outputs(1011) <= not(layer4_outputs(2970));
    layer5_outputs(1012) <= layer4_outputs(2518);
    layer5_outputs(1013) <= (layer4_outputs(1657)) or (layer4_outputs(667));
    layer5_outputs(1014) <= '1';
    layer5_outputs(1015) <= layer4_outputs(2164);
    layer5_outputs(1016) <= layer4_outputs(3875);
    layer5_outputs(1017) <= not(layer4_outputs(4796)) or (layer4_outputs(4216));
    layer5_outputs(1018) <= not(layer4_outputs(2612)) or (layer4_outputs(4779));
    layer5_outputs(1019) <= (layer4_outputs(3647)) and (layer4_outputs(969));
    layer5_outputs(1020) <= not(layer4_outputs(3844)) or (layer4_outputs(592));
    layer5_outputs(1021) <= '1';
    layer5_outputs(1022) <= not(layer4_outputs(3003));
    layer5_outputs(1023) <= not(layer4_outputs(3990)) or (layer4_outputs(889));
    layer5_outputs(1024) <= not((layer4_outputs(3393)) and (layer4_outputs(304)));
    layer5_outputs(1025) <= not(layer4_outputs(2166));
    layer5_outputs(1026) <= layer4_outputs(4031);
    layer5_outputs(1027) <= not(layer4_outputs(1359));
    layer5_outputs(1028) <= not(layer4_outputs(4858));
    layer5_outputs(1029) <= not(layer4_outputs(3106)) or (layer4_outputs(3869));
    layer5_outputs(1030) <= (layer4_outputs(4878)) and (layer4_outputs(460));
    layer5_outputs(1031) <= (layer4_outputs(1336)) and (layer4_outputs(2779));
    layer5_outputs(1032) <= not(layer4_outputs(3382));
    layer5_outputs(1033) <= (layer4_outputs(4740)) and not (layer4_outputs(387));
    layer5_outputs(1034) <= '0';
    layer5_outputs(1035) <= not((layer4_outputs(2960)) and (layer4_outputs(4229)));
    layer5_outputs(1036) <= not(layer4_outputs(4270));
    layer5_outputs(1037) <= (layer4_outputs(1108)) or (layer4_outputs(1618));
    layer5_outputs(1038) <= not((layer4_outputs(4610)) xor (layer4_outputs(3272)));
    layer5_outputs(1039) <= (layer4_outputs(3790)) and not (layer4_outputs(3004));
    layer5_outputs(1040) <= layer4_outputs(3176);
    layer5_outputs(1041) <= (layer4_outputs(2300)) and not (layer4_outputs(121));
    layer5_outputs(1042) <= (layer4_outputs(3281)) and (layer4_outputs(785));
    layer5_outputs(1043) <= (layer4_outputs(3182)) or (layer4_outputs(4671));
    layer5_outputs(1044) <= (layer4_outputs(4979)) and not (layer4_outputs(2926));
    layer5_outputs(1045) <= '1';
    layer5_outputs(1046) <= not((layer4_outputs(875)) or (layer4_outputs(3208)));
    layer5_outputs(1047) <= layer4_outputs(4981);
    layer5_outputs(1048) <= not((layer4_outputs(3418)) or (layer4_outputs(1600)));
    layer5_outputs(1049) <= '0';
    layer5_outputs(1050) <= layer4_outputs(865);
    layer5_outputs(1051) <= not((layer4_outputs(3260)) or (layer4_outputs(1298)));
    layer5_outputs(1052) <= not((layer4_outputs(2468)) and (layer4_outputs(3908)));
    layer5_outputs(1053) <= not((layer4_outputs(950)) or (layer4_outputs(3068)));
    layer5_outputs(1054) <= (layer4_outputs(842)) and (layer4_outputs(886));
    layer5_outputs(1055) <= not(layer4_outputs(1324));
    layer5_outputs(1056) <= (layer4_outputs(4402)) and not (layer4_outputs(4829));
    layer5_outputs(1057) <= layer4_outputs(1113);
    layer5_outputs(1058) <= layer4_outputs(3919);
    layer5_outputs(1059) <= (layer4_outputs(2446)) xor (layer4_outputs(1626));
    layer5_outputs(1060) <= not(layer4_outputs(4635));
    layer5_outputs(1061) <= '1';
    layer5_outputs(1062) <= layer4_outputs(3852);
    layer5_outputs(1063) <= not(layer4_outputs(3518));
    layer5_outputs(1064) <= (layer4_outputs(506)) or (layer4_outputs(3467));
    layer5_outputs(1065) <= not(layer4_outputs(1037));
    layer5_outputs(1066) <= (layer4_outputs(2098)) and not (layer4_outputs(3882));
    layer5_outputs(1067) <= not((layer4_outputs(2146)) and (layer4_outputs(4984)));
    layer5_outputs(1068) <= '0';
    layer5_outputs(1069) <= layer4_outputs(2632);
    layer5_outputs(1070) <= '0';
    layer5_outputs(1071) <= not(layer4_outputs(1892));
    layer5_outputs(1072) <= layer4_outputs(755);
    layer5_outputs(1073) <= not(layer4_outputs(3854));
    layer5_outputs(1074) <= not((layer4_outputs(3315)) or (layer4_outputs(1410)));
    layer5_outputs(1075) <= not(layer4_outputs(1375));
    layer5_outputs(1076) <= not(layer4_outputs(1252)) or (layer4_outputs(3500));
    layer5_outputs(1077) <= not((layer4_outputs(530)) or (layer4_outputs(1803)));
    layer5_outputs(1078) <= (layer4_outputs(2845)) or (layer4_outputs(2272));
    layer5_outputs(1079) <= not(layer4_outputs(1172)) or (layer4_outputs(958));
    layer5_outputs(1080) <= not(layer4_outputs(2028)) or (layer4_outputs(1991));
    layer5_outputs(1081) <= not(layer4_outputs(2390));
    layer5_outputs(1082) <= not(layer4_outputs(5052));
    layer5_outputs(1083) <= layer4_outputs(3109);
    layer5_outputs(1084) <= (layer4_outputs(1172)) xor (layer4_outputs(1751));
    layer5_outputs(1085) <= '1';
    layer5_outputs(1086) <= not(layer4_outputs(2633));
    layer5_outputs(1087) <= not(layer4_outputs(4135)) or (layer4_outputs(1198));
    layer5_outputs(1088) <= (layer4_outputs(1385)) and not (layer4_outputs(2981));
    layer5_outputs(1089) <= '0';
    layer5_outputs(1090) <= not(layer4_outputs(5095));
    layer5_outputs(1091) <= not(layer4_outputs(1381));
    layer5_outputs(1092) <= not((layer4_outputs(2918)) or (layer4_outputs(2680)));
    layer5_outputs(1093) <= layer4_outputs(4141);
    layer5_outputs(1094) <= not(layer4_outputs(615));
    layer5_outputs(1095) <= not(layer4_outputs(1831)) or (layer4_outputs(3135));
    layer5_outputs(1096) <= layer4_outputs(2291);
    layer5_outputs(1097) <= layer4_outputs(3317);
    layer5_outputs(1098) <= not(layer4_outputs(2390));
    layer5_outputs(1099) <= (layer4_outputs(4470)) or (layer4_outputs(1572));
    layer5_outputs(1100) <= not(layer4_outputs(235));
    layer5_outputs(1101) <= (layer4_outputs(1371)) and not (layer4_outputs(4243));
    layer5_outputs(1102) <= not((layer4_outputs(1120)) and (layer4_outputs(3355)));
    layer5_outputs(1103) <= (layer4_outputs(4824)) and (layer4_outputs(3880));
    layer5_outputs(1104) <= not(layer4_outputs(1941));
    layer5_outputs(1105) <= layer4_outputs(4424);
    layer5_outputs(1106) <= (layer4_outputs(2466)) and not (layer4_outputs(2202));
    layer5_outputs(1107) <= '0';
    layer5_outputs(1108) <= not(layer4_outputs(3047));
    layer5_outputs(1109) <= not(layer4_outputs(4974));
    layer5_outputs(1110) <= not((layer4_outputs(680)) or (layer4_outputs(518)));
    layer5_outputs(1111) <= layer4_outputs(2716);
    layer5_outputs(1112) <= (layer4_outputs(4097)) and not (layer4_outputs(866));
    layer5_outputs(1113) <= not(layer4_outputs(2668));
    layer5_outputs(1114) <= layer4_outputs(1123);
    layer5_outputs(1115) <= '0';
    layer5_outputs(1116) <= layer4_outputs(2216);
    layer5_outputs(1117) <= not((layer4_outputs(4248)) xor (layer4_outputs(4039)));
    layer5_outputs(1118) <= layer4_outputs(4481);
    layer5_outputs(1119) <= not(layer4_outputs(2238));
    layer5_outputs(1120) <= not((layer4_outputs(3832)) and (layer4_outputs(2001)));
    layer5_outputs(1121) <= layer4_outputs(51);
    layer5_outputs(1122) <= layer4_outputs(3843);
    layer5_outputs(1123) <= not(layer4_outputs(272));
    layer5_outputs(1124) <= not(layer4_outputs(2093));
    layer5_outputs(1125) <= not(layer4_outputs(3567));
    layer5_outputs(1126) <= not(layer4_outputs(2641));
    layer5_outputs(1127) <= (layer4_outputs(547)) or (layer4_outputs(268));
    layer5_outputs(1128) <= not(layer4_outputs(3741));
    layer5_outputs(1129) <= not(layer4_outputs(812));
    layer5_outputs(1130) <= not(layer4_outputs(5089)) or (layer4_outputs(683));
    layer5_outputs(1131) <= (layer4_outputs(3967)) xor (layer4_outputs(796));
    layer5_outputs(1132) <= not(layer4_outputs(570));
    layer5_outputs(1133) <= not(layer4_outputs(3924));
    layer5_outputs(1134) <= not((layer4_outputs(3290)) and (layer4_outputs(2655)));
    layer5_outputs(1135) <= layer4_outputs(1055);
    layer5_outputs(1136) <= layer4_outputs(4899);
    layer5_outputs(1137) <= layer4_outputs(172);
    layer5_outputs(1138) <= not(layer4_outputs(870));
    layer5_outputs(1139) <= '0';
    layer5_outputs(1140) <= layer4_outputs(1200);
    layer5_outputs(1141) <= layer4_outputs(4133);
    layer5_outputs(1142) <= (layer4_outputs(329)) and (layer4_outputs(4665));
    layer5_outputs(1143) <= not((layer4_outputs(2419)) or (layer4_outputs(1527)));
    layer5_outputs(1144) <= not(layer4_outputs(4313));
    layer5_outputs(1145) <= not((layer4_outputs(2646)) and (layer4_outputs(1591)));
    layer5_outputs(1146) <= (layer4_outputs(3323)) and (layer4_outputs(1087));
    layer5_outputs(1147) <= not((layer4_outputs(1181)) and (layer4_outputs(184)));
    layer5_outputs(1148) <= (layer4_outputs(587)) and (layer4_outputs(3110));
    layer5_outputs(1149) <= layer4_outputs(3173);
    layer5_outputs(1150) <= not(layer4_outputs(1247));
    layer5_outputs(1151) <= layer4_outputs(4672);
    layer5_outputs(1152) <= (layer4_outputs(62)) or (layer4_outputs(3542));
    layer5_outputs(1153) <= layer4_outputs(2912);
    layer5_outputs(1154) <= (layer4_outputs(112)) and not (layer4_outputs(1088));
    layer5_outputs(1155) <= (layer4_outputs(237)) or (layer4_outputs(363));
    layer5_outputs(1156) <= not(layer4_outputs(2943));
    layer5_outputs(1157) <= '0';
    layer5_outputs(1158) <= not(layer4_outputs(2884)) or (layer4_outputs(4800));
    layer5_outputs(1159) <= (layer4_outputs(4228)) and (layer4_outputs(4168));
    layer5_outputs(1160) <= not((layer4_outputs(1542)) xor (layer4_outputs(4569)));
    layer5_outputs(1161) <= (layer4_outputs(2260)) or (layer4_outputs(4666));
    layer5_outputs(1162) <= layer4_outputs(4560);
    layer5_outputs(1163) <= not((layer4_outputs(4698)) or (layer4_outputs(362)));
    layer5_outputs(1164) <= '0';
    layer5_outputs(1165) <= not(layer4_outputs(858));
    layer5_outputs(1166) <= (layer4_outputs(2481)) and not (layer4_outputs(3477));
    layer5_outputs(1167) <= '1';
    layer5_outputs(1168) <= '0';
    layer5_outputs(1169) <= not((layer4_outputs(2425)) xor (layer4_outputs(3743)));
    layer5_outputs(1170) <= (layer4_outputs(359)) and not (layer4_outputs(787));
    layer5_outputs(1171) <= (layer4_outputs(1450)) and not (layer4_outputs(2192));
    layer5_outputs(1172) <= not(layer4_outputs(4608)) or (layer4_outputs(2313));
    layer5_outputs(1173) <= not((layer4_outputs(4716)) and (layer4_outputs(5113)));
    layer5_outputs(1174) <= not(layer4_outputs(4896));
    layer5_outputs(1175) <= not((layer4_outputs(690)) and (layer4_outputs(1132)));
    layer5_outputs(1176) <= (layer4_outputs(2516)) and not (layer4_outputs(3550));
    layer5_outputs(1177) <= not(layer4_outputs(3930)) or (layer4_outputs(2756));
    layer5_outputs(1178) <= (layer4_outputs(861)) or (layer4_outputs(1334));
    layer5_outputs(1179) <= not(layer4_outputs(1609));
    layer5_outputs(1180) <= not(layer4_outputs(3910));
    layer5_outputs(1181) <= not(layer4_outputs(2007)) or (layer4_outputs(857));
    layer5_outputs(1182) <= not(layer4_outputs(3626)) or (layer4_outputs(3252));
    layer5_outputs(1183) <= (layer4_outputs(4528)) or (layer4_outputs(3611));
    layer5_outputs(1184) <= (layer4_outputs(4710)) or (layer4_outputs(3809));
    layer5_outputs(1185) <= not(layer4_outputs(4153));
    layer5_outputs(1186) <= not(layer4_outputs(311));
    layer5_outputs(1187) <= not((layer4_outputs(4229)) xor (layer4_outputs(4900)));
    layer5_outputs(1188) <= not((layer4_outputs(2291)) or (layer4_outputs(322)));
    layer5_outputs(1189) <= '1';
    layer5_outputs(1190) <= not(layer4_outputs(2274));
    layer5_outputs(1191) <= (layer4_outputs(2428)) and (layer4_outputs(4464));
    layer5_outputs(1192) <= not((layer4_outputs(114)) xor (layer4_outputs(3643)));
    layer5_outputs(1193) <= not(layer4_outputs(222)) or (layer4_outputs(2157));
    layer5_outputs(1194) <= not((layer4_outputs(2587)) or (layer4_outputs(245)));
    layer5_outputs(1195) <= layer4_outputs(345);
    layer5_outputs(1196) <= (layer4_outputs(2448)) and not (layer4_outputs(2391));
    layer5_outputs(1197) <= layer4_outputs(677);
    layer5_outputs(1198) <= not(layer4_outputs(3796));
    layer5_outputs(1199) <= not(layer4_outputs(1416));
    layer5_outputs(1200) <= not(layer4_outputs(1780)) or (layer4_outputs(2195));
    layer5_outputs(1201) <= not((layer4_outputs(3120)) or (layer4_outputs(1886)));
    layer5_outputs(1202) <= layer4_outputs(992);
    layer5_outputs(1203) <= (layer4_outputs(3117)) and not (layer4_outputs(2331));
    layer5_outputs(1204) <= '1';
    layer5_outputs(1205) <= not((layer4_outputs(1116)) xor (layer4_outputs(1198)));
    layer5_outputs(1206) <= not(layer4_outputs(1944));
    layer5_outputs(1207) <= (layer4_outputs(3815)) or (layer4_outputs(885));
    layer5_outputs(1208) <= (layer4_outputs(4905)) and not (layer4_outputs(3368));
    layer5_outputs(1209) <= not(layer4_outputs(1440));
    layer5_outputs(1210) <= not((layer4_outputs(3710)) xor (layer4_outputs(41)));
    layer5_outputs(1211) <= not((layer4_outputs(3673)) and (layer4_outputs(2661)));
    layer5_outputs(1212) <= (layer4_outputs(873)) or (layer4_outputs(2151));
    layer5_outputs(1213) <= not((layer4_outputs(2131)) or (layer4_outputs(2)));
    layer5_outputs(1214) <= '0';
    layer5_outputs(1215) <= (layer4_outputs(2244)) and not (layer4_outputs(5063));
    layer5_outputs(1216) <= not((layer4_outputs(563)) and (layer4_outputs(3266)));
    layer5_outputs(1217) <= not(layer4_outputs(2965));
    layer5_outputs(1218) <= '0';
    layer5_outputs(1219) <= not((layer4_outputs(209)) and (layer4_outputs(4526)));
    layer5_outputs(1220) <= layer4_outputs(1578);
    layer5_outputs(1221) <= layer4_outputs(3156);
    layer5_outputs(1222) <= not(layer4_outputs(3823)) or (layer4_outputs(3046));
    layer5_outputs(1223) <= not((layer4_outputs(1839)) and (layer4_outputs(831)));
    layer5_outputs(1224) <= (layer4_outputs(812)) or (layer4_outputs(290));
    layer5_outputs(1225) <= not(layer4_outputs(2833));
    layer5_outputs(1226) <= '1';
    layer5_outputs(1227) <= layer4_outputs(1726);
    layer5_outputs(1228) <= not(layer4_outputs(4613));
    layer5_outputs(1229) <= not(layer4_outputs(4975)) or (layer4_outputs(438));
    layer5_outputs(1230) <= layer4_outputs(1179);
    layer5_outputs(1231) <= not(layer4_outputs(2323)) or (layer4_outputs(1376));
    layer5_outputs(1232) <= not(layer4_outputs(2596));
    layer5_outputs(1233) <= (layer4_outputs(4867)) or (layer4_outputs(2408));
    layer5_outputs(1234) <= layer4_outputs(4572);
    layer5_outputs(1235) <= layer4_outputs(4002);
    layer5_outputs(1236) <= layer4_outputs(5049);
    layer5_outputs(1237) <= not((layer4_outputs(2472)) or (layer4_outputs(1393)));
    layer5_outputs(1238) <= (layer4_outputs(3158)) and (layer4_outputs(1258));
    layer5_outputs(1239) <= '1';
    layer5_outputs(1240) <= not((layer4_outputs(1036)) or (layer4_outputs(3388)));
    layer5_outputs(1241) <= (layer4_outputs(4091)) and not (layer4_outputs(3767));
    layer5_outputs(1242) <= layer4_outputs(2812);
    layer5_outputs(1243) <= (layer4_outputs(358)) and not (layer4_outputs(2533));
    layer5_outputs(1244) <= '0';
    layer5_outputs(1245) <= layer4_outputs(2003);
    layer5_outputs(1246) <= not(layer4_outputs(3585)) or (layer4_outputs(2271));
    layer5_outputs(1247) <= '1';
    layer5_outputs(1248) <= (layer4_outputs(2216)) or (layer4_outputs(4403));
    layer5_outputs(1249) <= not(layer4_outputs(3010));
    layer5_outputs(1250) <= not(layer4_outputs(4825));
    layer5_outputs(1251) <= not(layer4_outputs(2593));
    layer5_outputs(1252) <= layer4_outputs(419);
    layer5_outputs(1253) <= layer4_outputs(2196);
    layer5_outputs(1254) <= '1';
    layer5_outputs(1255) <= not(layer4_outputs(918));
    layer5_outputs(1256) <= '1';
    layer5_outputs(1257) <= not(layer4_outputs(2546)) or (layer4_outputs(468));
    layer5_outputs(1258) <= not(layer4_outputs(1848));
    layer5_outputs(1259) <= not(layer4_outputs(2530));
    layer5_outputs(1260) <= not(layer4_outputs(1415));
    layer5_outputs(1261) <= not(layer4_outputs(1115));
    layer5_outputs(1262) <= (layer4_outputs(1805)) and (layer4_outputs(3386));
    layer5_outputs(1263) <= (layer4_outputs(430)) and not (layer4_outputs(2437));
    layer5_outputs(1264) <= not(layer4_outputs(3972));
    layer5_outputs(1265) <= not(layer4_outputs(3504)) or (layer4_outputs(5086));
    layer5_outputs(1266) <= layer4_outputs(2275);
    layer5_outputs(1267) <= not(layer4_outputs(2027)) or (layer4_outputs(913));
    layer5_outputs(1268) <= (layer4_outputs(3322)) and not (layer4_outputs(317));
    layer5_outputs(1269) <= not(layer4_outputs(3029));
    layer5_outputs(1270) <= not((layer4_outputs(694)) and (layer4_outputs(4715)));
    layer5_outputs(1271) <= (layer4_outputs(1363)) and not (layer4_outputs(3696));
    layer5_outputs(1272) <= (layer4_outputs(3174)) and not (layer4_outputs(3862));
    layer5_outputs(1273) <= not((layer4_outputs(3277)) xor (layer4_outputs(1230)));
    layer5_outputs(1274) <= not(layer4_outputs(3533)) or (layer4_outputs(516));
    layer5_outputs(1275) <= '1';
    layer5_outputs(1276) <= layer4_outputs(4699);
    layer5_outputs(1277) <= (layer4_outputs(4815)) and (layer4_outputs(583));
    layer5_outputs(1278) <= (layer4_outputs(2121)) or (layer4_outputs(2205));
    layer5_outputs(1279) <= not(layer4_outputs(999)) or (layer4_outputs(374));
    layer5_outputs(1280) <= not(layer4_outputs(4116)) or (layer4_outputs(4425));
    layer5_outputs(1281) <= not((layer4_outputs(3718)) or (layer4_outputs(429)));
    layer5_outputs(1282) <= '0';
    layer5_outputs(1283) <= not(layer4_outputs(1306)) or (layer4_outputs(4743));
    layer5_outputs(1284) <= not(layer4_outputs(1458)) or (layer4_outputs(702));
    layer5_outputs(1285) <= not(layer4_outputs(4535));
    layer5_outputs(1286) <= '1';
    layer5_outputs(1287) <= not(layer4_outputs(3178));
    layer5_outputs(1288) <= (layer4_outputs(3280)) and not (layer4_outputs(2317));
    layer5_outputs(1289) <= (layer4_outputs(2222)) and not (layer4_outputs(1858));
    layer5_outputs(1290) <= (layer4_outputs(969)) and (layer4_outputs(2957));
    layer5_outputs(1291) <= not((layer4_outputs(540)) and (layer4_outputs(1948)));
    layer5_outputs(1292) <= not((layer4_outputs(1146)) xor (layer4_outputs(3623)));
    layer5_outputs(1293) <= '0';
    layer5_outputs(1294) <= not(layer4_outputs(2421)) or (layer4_outputs(2160));
    layer5_outputs(1295) <= (layer4_outputs(554)) xor (layer4_outputs(4175));
    layer5_outputs(1296) <= not(layer4_outputs(460));
    layer5_outputs(1297) <= (layer4_outputs(2963)) and not (layer4_outputs(4104));
    layer5_outputs(1298) <= not(layer4_outputs(1702)) or (layer4_outputs(3756));
    layer5_outputs(1299) <= (layer4_outputs(4874)) or (layer4_outputs(3098));
    layer5_outputs(1300) <= not(layer4_outputs(2068)) or (layer4_outputs(610));
    layer5_outputs(1301) <= (layer4_outputs(2247)) and not (layer4_outputs(710));
    layer5_outputs(1302) <= (layer4_outputs(3011)) and not (layer4_outputs(921));
    layer5_outputs(1303) <= not(layer4_outputs(1776)) or (layer4_outputs(2069));
    layer5_outputs(1304) <= not(layer4_outputs(3856));
    layer5_outputs(1305) <= not((layer4_outputs(1700)) or (layer4_outputs(1775)));
    layer5_outputs(1306) <= (layer4_outputs(2812)) or (layer4_outputs(821));
    layer5_outputs(1307) <= not(layer4_outputs(2409));
    layer5_outputs(1308) <= (layer4_outputs(2193)) xor (layer4_outputs(3776));
    layer5_outputs(1309) <= (layer4_outputs(3629)) xor (layer4_outputs(1208));
    layer5_outputs(1310) <= (layer4_outputs(1174)) and (layer4_outputs(497));
    layer5_outputs(1311) <= not(layer4_outputs(1646)) or (layer4_outputs(3433));
    layer5_outputs(1312) <= layer4_outputs(4722);
    layer5_outputs(1313) <= not(layer4_outputs(271)) or (layer4_outputs(448));
    layer5_outputs(1314) <= layer4_outputs(2753);
    layer5_outputs(1315) <= layer4_outputs(26);
    layer5_outputs(1316) <= not((layer4_outputs(1709)) or (layer4_outputs(1629)));
    layer5_outputs(1317) <= layer4_outputs(4170);
    layer5_outputs(1318) <= (layer4_outputs(2964)) or (layer4_outputs(1843));
    layer5_outputs(1319) <= not(layer4_outputs(4859)) or (layer4_outputs(2303));
    layer5_outputs(1320) <= not(layer4_outputs(654)) or (layer4_outputs(1602));
    layer5_outputs(1321) <= '1';
    layer5_outputs(1322) <= (layer4_outputs(3757)) and not (layer4_outputs(3952));
    layer5_outputs(1323) <= '0';
    layer5_outputs(1324) <= '0';
    layer5_outputs(1325) <= not((layer4_outputs(1850)) xor (layer4_outputs(1619)));
    layer5_outputs(1326) <= not(layer4_outputs(1196));
    layer5_outputs(1327) <= (layer4_outputs(1900)) xor (layer4_outputs(2043));
    layer5_outputs(1328) <= (layer4_outputs(100)) and not (layer4_outputs(4549));
    layer5_outputs(1329) <= layer4_outputs(1779);
    layer5_outputs(1330) <= not(layer4_outputs(3568)) or (layer4_outputs(2997));
    layer5_outputs(1331) <= (layer4_outputs(2061)) and not (layer4_outputs(1048));
    layer5_outputs(1332) <= layer4_outputs(4769);
    layer5_outputs(1333) <= not((layer4_outputs(2288)) and (layer4_outputs(2018)));
    layer5_outputs(1334) <= layer4_outputs(2508);
    layer5_outputs(1335) <= not((layer4_outputs(3921)) and (layer4_outputs(4485)));
    layer5_outputs(1336) <= not((layer4_outputs(2255)) or (layer4_outputs(2393)));
    layer5_outputs(1337) <= (layer4_outputs(2854)) and not (layer4_outputs(1955));
    layer5_outputs(1338) <= not(layer4_outputs(1513)) or (layer4_outputs(1255));
    layer5_outputs(1339) <= layer4_outputs(3747);
    layer5_outputs(1340) <= not(layer4_outputs(5113));
    layer5_outputs(1341) <= '0';
    layer5_outputs(1342) <= layer4_outputs(3808);
    layer5_outputs(1343) <= not(layer4_outputs(1828));
    layer5_outputs(1344) <= '0';
    layer5_outputs(1345) <= not((layer4_outputs(4277)) xor (layer4_outputs(372)));
    layer5_outputs(1346) <= (layer4_outputs(3082)) xor (layer4_outputs(4087));
    layer5_outputs(1347) <= layer4_outputs(1324);
    layer5_outputs(1348) <= '1';
    layer5_outputs(1349) <= not((layer4_outputs(455)) and (layer4_outputs(1217)));
    layer5_outputs(1350) <= not(layer4_outputs(339));
    layer5_outputs(1351) <= layer4_outputs(2664);
    layer5_outputs(1352) <= layer4_outputs(287);
    layer5_outputs(1353) <= not((layer4_outputs(3171)) or (layer4_outputs(780)));
    layer5_outputs(1354) <= (layer4_outputs(4693)) and not (layer4_outputs(1807));
    layer5_outputs(1355) <= not(layer4_outputs(3632)) or (layer4_outputs(4997));
    layer5_outputs(1356) <= layer4_outputs(2127);
    layer5_outputs(1357) <= layer4_outputs(3424);
    layer5_outputs(1358) <= layer4_outputs(1986);
    layer5_outputs(1359) <= (layer4_outputs(92)) or (layer4_outputs(2074));
    layer5_outputs(1360) <= (layer4_outputs(1041)) and not (layer4_outputs(2621));
    layer5_outputs(1361) <= '1';
    layer5_outputs(1362) <= (layer4_outputs(4074)) and not (layer4_outputs(2166));
    layer5_outputs(1363) <= (layer4_outputs(2825)) and not (layer4_outputs(5051));
    layer5_outputs(1364) <= layer4_outputs(1863);
    layer5_outputs(1365) <= '0';
    layer5_outputs(1366) <= not(layer4_outputs(95));
    layer5_outputs(1367) <= (layer4_outputs(3229)) and (layer4_outputs(2911));
    layer5_outputs(1368) <= (layer4_outputs(3898)) or (layer4_outputs(722));
    layer5_outputs(1369) <= (layer4_outputs(2581)) xor (layer4_outputs(263));
    layer5_outputs(1370) <= (layer4_outputs(1999)) or (layer4_outputs(836));
    layer5_outputs(1371) <= not(layer4_outputs(1520));
    layer5_outputs(1372) <= not((layer4_outputs(101)) and (layer4_outputs(256)));
    layer5_outputs(1373) <= not(layer4_outputs(2231)) or (layer4_outputs(3580));
    layer5_outputs(1374) <= not(layer4_outputs(4718)) or (layer4_outputs(2588));
    layer5_outputs(1375) <= not(layer4_outputs(1733));
    layer5_outputs(1376) <= (layer4_outputs(968)) and (layer4_outputs(2511));
    layer5_outputs(1377) <= (layer4_outputs(1536)) and (layer4_outputs(1498));
    layer5_outputs(1378) <= not(layer4_outputs(2054));
    layer5_outputs(1379) <= layer4_outputs(4895);
    layer5_outputs(1380) <= not((layer4_outputs(2404)) and (layer4_outputs(4609)));
    layer5_outputs(1381) <= not(layer4_outputs(4684));
    layer5_outputs(1382) <= not(layer4_outputs(3009));
    layer5_outputs(1383) <= not(layer4_outputs(4004)) or (layer4_outputs(1666));
    layer5_outputs(1384) <= layer4_outputs(1974);
    layer5_outputs(1385) <= (layer4_outputs(4208)) or (layer4_outputs(641));
    layer5_outputs(1386) <= (layer4_outputs(3797)) and not (layer4_outputs(4775));
    layer5_outputs(1387) <= not(layer4_outputs(3877));
    layer5_outputs(1388) <= layer4_outputs(1014);
    layer5_outputs(1389) <= (layer4_outputs(4997)) xor (layer4_outputs(514));
    layer5_outputs(1390) <= not((layer4_outputs(4395)) xor (layer4_outputs(4472)));
    layer5_outputs(1391) <= layer4_outputs(3000);
    layer5_outputs(1392) <= layer4_outputs(3554);
    layer5_outputs(1393) <= not(layer4_outputs(3870));
    layer5_outputs(1394) <= not(layer4_outputs(4189));
    layer5_outputs(1395) <= not((layer4_outputs(2642)) and (layer4_outputs(1662)));
    layer5_outputs(1396) <= not(layer4_outputs(2748));
    layer5_outputs(1397) <= layer4_outputs(4643);
    layer5_outputs(1398) <= not(layer4_outputs(2173));
    layer5_outputs(1399) <= not((layer4_outputs(4020)) xor (layer4_outputs(1199)));
    layer5_outputs(1400) <= not(layer4_outputs(3942));
    layer5_outputs(1401) <= (layer4_outputs(823)) and not (layer4_outputs(3830));
    layer5_outputs(1402) <= layer4_outputs(23);
    layer5_outputs(1403) <= (layer4_outputs(938)) and not (layer4_outputs(4872));
    layer5_outputs(1404) <= '1';
    layer5_outputs(1405) <= layer4_outputs(1929);
    layer5_outputs(1406) <= not(layer4_outputs(739));
    layer5_outputs(1407) <= (layer4_outputs(1757)) and not (layer4_outputs(4337));
    layer5_outputs(1408) <= layer4_outputs(4871);
    layer5_outputs(1409) <= layer4_outputs(3451);
    layer5_outputs(1410) <= (layer4_outputs(2052)) and not (layer4_outputs(249));
    layer5_outputs(1411) <= not(layer4_outputs(4759));
    layer5_outputs(1412) <= not(layer4_outputs(5042));
    layer5_outputs(1413) <= (layer4_outputs(3822)) and not (layer4_outputs(3471));
    layer5_outputs(1414) <= (layer4_outputs(3480)) and (layer4_outputs(228));
    layer5_outputs(1415) <= layer4_outputs(4586);
    layer5_outputs(1416) <= (layer4_outputs(906)) and not (layer4_outputs(4937));
    layer5_outputs(1417) <= (layer4_outputs(553)) or (layer4_outputs(2997));
    layer5_outputs(1418) <= layer4_outputs(3199);
    layer5_outputs(1419) <= not((layer4_outputs(2267)) and (layer4_outputs(542)));
    layer5_outputs(1420) <= not(layer4_outputs(2383)) or (layer4_outputs(896));
    layer5_outputs(1421) <= layer4_outputs(1815);
    layer5_outputs(1422) <= not(layer4_outputs(3985));
    layer5_outputs(1423) <= not(layer4_outputs(2994)) or (layer4_outputs(1553));
    layer5_outputs(1424) <= '1';
    layer5_outputs(1425) <= (layer4_outputs(4861)) and not (layer4_outputs(3541));
    layer5_outputs(1426) <= not(layer4_outputs(3998));
    layer5_outputs(1427) <= (layer4_outputs(2726)) and not (layer4_outputs(915));
    layer5_outputs(1428) <= layer4_outputs(295);
    layer5_outputs(1429) <= not(layer4_outputs(2610));
    layer5_outputs(1430) <= layer4_outputs(477);
    layer5_outputs(1431) <= not(layer4_outputs(4084));
    layer5_outputs(1432) <= (layer4_outputs(3650)) and not (layer4_outputs(547));
    layer5_outputs(1433) <= (layer4_outputs(4633)) xor (layer4_outputs(3128));
    layer5_outputs(1434) <= (layer4_outputs(3659)) xor (layer4_outputs(2914));
    layer5_outputs(1435) <= not(layer4_outputs(3814)) or (layer4_outputs(1581));
    layer5_outputs(1436) <= not(layer4_outputs(2497));
    layer5_outputs(1437) <= layer4_outputs(1340);
    layer5_outputs(1438) <= (layer4_outputs(2108)) and not (layer4_outputs(4062));
    layer5_outputs(1439) <= not(layer4_outputs(1654)) or (layer4_outputs(2497));
    layer5_outputs(1440) <= (layer4_outputs(4637)) and (layer4_outputs(5084));
    layer5_outputs(1441) <= not(layer4_outputs(2848)) or (layer4_outputs(4772));
    layer5_outputs(1442) <= not(layer4_outputs(4993)) or (layer4_outputs(4414));
    layer5_outputs(1443) <= not(layer4_outputs(1932));
    layer5_outputs(1444) <= not(layer4_outputs(3332)) or (layer4_outputs(3854));
    layer5_outputs(1445) <= not(layer4_outputs(2547));
    layer5_outputs(1446) <= not((layer4_outputs(3728)) or (layer4_outputs(4451)));
    layer5_outputs(1447) <= (layer4_outputs(689)) and not (layer4_outputs(5106));
    layer5_outputs(1448) <= (layer4_outputs(506)) and not (layer4_outputs(5080));
    layer5_outputs(1449) <= (layer4_outputs(2392)) and (layer4_outputs(4135));
    layer5_outputs(1450) <= not(layer4_outputs(2620)) or (layer4_outputs(4086));
    layer5_outputs(1451) <= not((layer4_outputs(2931)) and (layer4_outputs(385)));
    layer5_outputs(1452) <= layer4_outputs(2615);
    layer5_outputs(1453) <= not(layer4_outputs(2890)) or (layer4_outputs(4115));
    layer5_outputs(1454) <= '0';
    layer5_outputs(1455) <= (layer4_outputs(3342)) or (layer4_outputs(4385));
    layer5_outputs(1456) <= (layer4_outputs(1003)) and not (layer4_outputs(4227));
    layer5_outputs(1457) <= not((layer4_outputs(3888)) or (layer4_outputs(4260)));
    layer5_outputs(1458) <= not(layer4_outputs(4161));
    layer5_outputs(1459) <= (layer4_outputs(2578)) and not (layer4_outputs(2316));
    layer5_outputs(1460) <= not((layer4_outputs(1079)) and (layer4_outputs(857)));
    layer5_outputs(1461) <= not(layer4_outputs(916));
    layer5_outputs(1462) <= '1';
    layer5_outputs(1463) <= '1';
    layer5_outputs(1464) <= (layer4_outputs(169)) and not (layer4_outputs(3191));
    layer5_outputs(1465) <= not(layer4_outputs(3415));
    layer5_outputs(1466) <= (layer4_outputs(4652)) and not (layer4_outputs(4329));
    layer5_outputs(1467) <= not((layer4_outputs(4936)) or (layer4_outputs(2899)));
    layer5_outputs(1468) <= not(layer4_outputs(2823));
    layer5_outputs(1469) <= not(layer4_outputs(734));
    layer5_outputs(1470) <= (layer4_outputs(2696)) and not (layer4_outputs(935));
    layer5_outputs(1471) <= not(layer4_outputs(1537)) or (layer4_outputs(4893));
    layer5_outputs(1472) <= not(layer4_outputs(786));
    layer5_outputs(1473) <= not((layer4_outputs(2315)) and (layer4_outputs(336)));
    layer5_outputs(1474) <= not(layer4_outputs(466));
    layer5_outputs(1475) <= not((layer4_outputs(4901)) xor (layer4_outputs(734)));
    layer5_outputs(1476) <= (layer4_outputs(408)) xor (layer4_outputs(2888));
    layer5_outputs(1477) <= (layer4_outputs(4785)) and (layer4_outputs(2540));
    layer5_outputs(1478) <= '0';
    layer5_outputs(1479) <= not(layer4_outputs(3720));
    layer5_outputs(1480) <= layer4_outputs(4217);
    layer5_outputs(1481) <= '1';
    layer5_outputs(1482) <= not((layer4_outputs(4892)) or (layer4_outputs(2347)));
    layer5_outputs(1483) <= (layer4_outputs(224)) and not (layer4_outputs(4309));
    layer5_outputs(1484) <= not(layer4_outputs(3249)) or (layer4_outputs(1577));
    layer5_outputs(1485) <= (layer4_outputs(4907)) or (layer4_outputs(3932));
    layer5_outputs(1486) <= not(layer4_outputs(2936));
    layer5_outputs(1487) <= '0';
    layer5_outputs(1488) <= (layer4_outputs(2241)) xor (layer4_outputs(13));
    layer5_outputs(1489) <= (layer4_outputs(2747)) and not (layer4_outputs(2890));
    layer5_outputs(1490) <= (layer4_outputs(3292)) xor (layer4_outputs(2885));
    layer5_outputs(1491) <= layer4_outputs(1096);
    layer5_outputs(1492) <= not((layer4_outputs(4118)) xor (layer4_outputs(4486)));
    layer5_outputs(1493) <= not((layer4_outputs(4102)) and (layer4_outputs(1032)));
    layer5_outputs(1494) <= not(layer4_outputs(3481));
    layer5_outputs(1495) <= (layer4_outputs(4544)) or (layer4_outputs(1524));
    layer5_outputs(1496) <= '0';
    layer5_outputs(1497) <= (layer4_outputs(2281)) or (layer4_outputs(2863));
    layer5_outputs(1498) <= not(layer4_outputs(3606));
    layer5_outputs(1499) <= not((layer4_outputs(418)) and (layer4_outputs(4546)));
    layer5_outputs(1500) <= not(layer4_outputs(2452));
    layer5_outputs(1501) <= not(layer4_outputs(2878)) or (layer4_outputs(834));
    layer5_outputs(1502) <= not((layer4_outputs(2778)) or (layer4_outputs(1893)));
    layer5_outputs(1503) <= not((layer4_outputs(3621)) and (layer4_outputs(120)));
    layer5_outputs(1504) <= not(layer4_outputs(4664));
    layer5_outputs(1505) <= (layer4_outputs(3302)) and (layer4_outputs(2212));
    layer5_outputs(1506) <= not((layer4_outputs(4650)) and (layer4_outputs(2625)));
    layer5_outputs(1507) <= layer4_outputs(92);
    layer5_outputs(1508) <= (layer4_outputs(2340)) and not (layer4_outputs(4368));
    layer5_outputs(1509) <= not(layer4_outputs(4722));
    layer5_outputs(1510) <= layer4_outputs(2982);
    layer5_outputs(1511) <= layer4_outputs(413);
    layer5_outputs(1512) <= layer4_outputs(1521);
    layer5_outputs(1513) <= not(layer4_outputs(4961));
    layer5_outputs(1514) <= not((layer4_outputs(978)) xor (layer4_outputs(170)));
    layer5_outputs(1515) <= (layer4_outputs(933)) xor (layer4_outputs(134));
    layer5_outputs(1516) <= layer4_outputs(4570);
    layer5_outputs(1517) <= (layer4_outputs(3005)) and (layer4_outputs(3951));
    layer5_outputs(1518) <= layer4_outputs(4638);
    layer5_outputs(1519) <= not(layer4_outputs(4805));
    layer5_outputs(1520) <= not(layer4_outputs(1391));
    layer5_outputs(1521) <= not((layer4_outputs(3514)) or (layer4_outputs(98)));
    layer5_outputs(1522) <= (layer4_outputs(2891)) and not (layer4_outputs(1160));
    layer5_outputs(1523) <= (layer4_outputs(3066)) or (layer4_outputs(3427));
    layer5_outputs(1524) <= not((layer4_outputs(4958)) and (layer4_outputs(1186)));
    layer5_outputs(1525) <= (layer4_outputs(4933)) and not (layer4_outputs(3532));
    layer5_outputs(1526) <= (layer4_outputs(70)) and (layer4_outputs(551));
    layer5_outputs(1527) <= (layer4_outputs(4614)) or (layer4_outputs(4776));
    layer5_outputs(1528) <= not(layer4_outputs(1638));
    layer5_outputs(1529) <= not(layer4_outputs(2810));
    layer5_outputs(1530) <= layer4_outputs(5109);
    layer5_outputs(1531) <= not(layer4_outputs(3052));
    layer5_outputs(1532) <= not(layer4_outputs(4132));
    layer5_outputs(1533) <= layer4_outputs(2832);
    layer5_outputs(1534) <= layer4_outputs(239);
    layer5_outputs(1535) <= (layer4_outputs(2391)) or (layer4_outputs(1701));
    layer5_outputs(1536) <= layer4_outputs(4678);
    layer5_outputs(1537) <= not((layer4_outputs(3774)) xor (layer4_outputs(564)));
    layer5_outputs(1538) <= layer4_outputs(1046);
    layer5_outputs(1539) <= '0';
    layer5_outputs(1540) <= not(layer4_outputs(2176));
    layer5_outputs(1541) <= layer4_outputs(4443);
    layer5_outputs(1542) <= layer4_outputs(3225);
    layer5_outputs(1543) <= (layer4_outputs(4177)) xor (layer4_outputs(4184));
    layer5_outputs(1544) <= (layer4_outputs(1846)) or (layer4_outputs(1477));
    layer5_outputs(1545) <= not(layer4_outputs(1301)) or (layer4_outputs(3829));
    layer5_outputs(1546) <= '0';
    layer5_outputs(1547) <= (layer4_outputs(1362)) and (layer4_outputs(2344));
    layer5_outputs(1548) <= (layer4_outputs(4315)) and (layer4_outputs(162));
    layer5_outputs(1549) <= not(layer4_outputs(4680));
    layer5_outputs(1550) <= layer4_outputs(3827);
    layer5_outputs(1551) <= '0';
    layer5_outputs(1552) <= layer4_outputs(4335);
    layer5_outputs(1553) <= layer4_outputs(2896);
    layer5_outputs(1554) <= not(layer4_outputs(4158));
    layer5_outputs(1555) <= not(layer4_outputs(706));
    layer5_outputs(1556) <= not(layer4_outputs(3588)) or (layer4_outputs(3464));
    layer5_outputs(1557) <= (layer4_outputs(1980)) or (layer4_outputs(3270));
    layer5_outputs(1558) <= (layer4_outputs(1270)) and not (layer4_outputs(2729));
    layer5_outputs(1559) <= '0';
    layer5_outputs(1560) <= not(layer4_outputs(1084));
    layer5_outputs(1561) <= '1';
    layer5_outputs(1562) <= not(layer4_outputs(448)) or (layer4_outputs(425));
    layer5_outputs(1563) <= (layer4_outputs(1376)) or (layer4_outputs(3529));
    layer5_outputs(1564) <= layer4_outputs(2811);
    layer5_outputs(1565) <= not(layer4_outputs(929)) or (layer4_outputs(2220));
    layer5_outputs(1566) <= not((layer4_outputs(1613)) or (layer4_outputs(3512)));
    layer5_outputs(1567) <= layer4_outputs(2954);
    layer5_outputs(1568) <= not((layer4_outputs(4079)) or (layer4_outputs(663)));
    layer5_outputs(1569) <= layer4_outputs(132);
    layer5_outputs(1570) <= not((layer4_outputs(5082)) xor (layer4_outputs(4968)));
    layer5_outputs(1571) <= not(layer4_outputs(4236));
    layer5_outputs(1572) <= not(layer4_outputs(5092));
    layer5_outputs(1573) <= not(layer4_outputs(2507));
    layer5_outputs(1574) <= (layer4_outputs(1890)) and not (layer4_outputs(3424));
    layer5_outputs(1575) <= layer4_outputs(4918);
    layer5_outputs(1576) <= not((layer4_outputs(1778)) or (layer4_outputs(4880)));
    layer5_outputs(1577) <= not((layer4_outputs(2284)) and (layer4_outputs(162)));
    layer5_outputs(1578) <= (layer4_outputs(2801)) and not (layer4_outputs(3461));
    layer5_outputs(1579) <= not((layer4_outputs(4823)) xor (layer4_outputs(3813)));
    layer5_outputs(1580) <= (layer4_outputs(3576)) and not (layer4_outputs(2224));
    layer5_outputs(1581) <= layer4_outputs(4729);
    layer5_outputs(1582) <= not(layer4_outputs(3294));
    layer5_outputs(1583) <= layer4_outputs(4727);
    layer5_outputs(1584) <= not(layer4_outputs(2704));
    layer5_outputs(1585) <= not(layer4_outputs(4310));
    layer5_outputs(1586) <= not(layer4_outputs(2304)) or (layer4_outputs(3085));
    layer5_outputs(1587) <= (layer4_outputs(928)) or (layer4_outputs(3860));
    layer5_outputs(1588) <= not(layer4_outputs(4999)) or (layer4_outputs(511));
    layer5_outputs(1589) <= layer4_outputs(1906);
    layer5_outputs(1590) <= '1';
    layer5_outputs(1591) <= not((layer4_outputs(3504)) or (layer4_outputs(3860)));
    layer5_outputs(1592) <= not(layer4_outputs(2619)) or (layer4_outputs(4970));
    layer5_outputs(1593) <= (layer4_outputs(1457)) xor (layer4_outputs(202));
    layer5_outputs(1594) <= layer4_outputs(4193);
    layer5_outputs(1595) <= (layer4_outputs(174)) and not (layer4_outputs(1077));
    layer5_outputs(1596) <= (layer4_outputs(2639)) and not (layer4_outputs(601));
    layer5_outputs(1597) <= '1';
    layer5_outputs(1598) <= layer4_outputs(1420);
    layer5_outputs(1599) <= layer4_outputs(4702);
    layer5_outputs(1600) <= not((layer4_outputs(155)) and (layer4_outputs(2810)));
    layer5_outputs(1601) <= (layer4_outputs(3874)) and not (layer4_outputs(3453));
    layer5_outputs(1602) <= not(layer4_outputs(2649));
    layer5_outputs(1603) <= '1';
    layer5_outputs(1604) <= not((layer4_outputs(84)) and (layer4_outputs(1981)));
    layer5_outputs(1605) <= not(layer4_outputs(431)) or (layer4_outputs(2111));
    layer5_outputs(1606) <= not(layer4_outputs(1748));
    layer5_outputs(1607) <= not(layer4_outputs(4489)) or (layer4_outputs(3514));
    layer5_outputs(1608) <= (layer4_outputs(3562)) and not (layer4_outputs(1072));
    layer5_outputs(1609) <= not(layer4_outputs(2662));
    layer5_outputs(1610) <= not(layer4_outputs(3080));
    layer5_outputs(1611) <= not(layer4_outputs(1488)) or (layer4_outputs(1600));
    layer5_outputs(1612) <= layer4_outputs(4497);
    layer5_outputs(1613) <= layer4_outputs(1264);
    layer5_outputs(1614) <= layer4_outputs(3520);
    layer5_outputs(1615) <= not(layer4_outputs(1679));
    layer5_outputs(1616) <= '0';
    layer5_outputs(1617) <= (layer4_outputs(1925)) and not (layer4_outputs(2967));
    layer5_outputs(1618) <= (layer4_outputs(913)) or (layer4_outputs(5039));
    layer5_outputs(1619) <= not(layer4_outputs(930)) or (layer4_outputs(2969));
    layer5_outputs(1620) <= (layer4_outputs(2413)) and not (layer4_outputs(701));
    layer5_outputs(1621) <= layer4_outputs(690);
    layer5_outputs(1622) <= not(layer4_outputs(3482));
    layer5_outputs(1623) <= (layer4_outputs(3246)) and (layer4_outputs(4174));
    layer5_outputs(1624) <= '0';
    layer5_outputs(1625) <= (layer4_outputs(4897)) or (layer4_outputs(3691));
    layer5_outputs(1626) <= (layer4_outputs(2525)) or (layer4_outputs(127));
    layer5_outputs(1627) <= not((layer4_outputs(4556)) and (layer4_outputs(4780)));
    layer5_outputs(1628) <= layer4_outputs(4353);
    layer5_outputs(1629) <= (layer4_outputs(2692)) and not (layer4_outputs(1738));
    layer5_outputs(1630) <= (layer4_outputs(11)) xor (layer4_outputs(5066));
    layer5_outputs(1631) <= not(layer4_outputs(1618));
    layer5_outputs(1632) <= (layer4_outputs(2692)) and not (layer4_outputs(3458));
    layer5_outputs(1633) <= not((layer4_outputs(399)) or (layer4_outputs(3383)));
    layer5_outputs(1634) <= not(layer4_outputs(825));
    layer5_outputs(1635) <= not(layer4_outputs(3055));
    layer5_outputs(1636) <= layer4_outputs(2020);
    layer5_outputs(1637) <= not(layer4_outputs(2993));
    layer5_outputs(1638) <= (layer4_outputs(4885)) xor (layer4_outputs(1416));
    layer5_outputs(1639) <= layer4_outputs(1053);
    layer5_outputs(1640) <= not(layer4_outputs(226));
    layer5_outputs(1641) <= '0';
    layer5_outputs(1642) <= (layer4_outputs(3724)) and not (layer4_outputs(229));
    layer5_outputs(1643) <= layer4_outputs(2366);
    layer5_outputs(1644) <= layer4_outputs(3006);
    layer5_outputs(1645) <= not(layer4_outputs(2170));
    layer5_outputs(1646) <= not(layer4_outputs(2766)) or (layer4_outputs(4254));
    layer5_outputs(1647) <= not(layer4_outputs(4737));
    layer5_outputs(1648) <= layer4_outputs(3841);
    layer5_outputs(1649) <= (layer4_outputs(3523)) and not (layer4_outputs(3231));
    layer5_outputs(1650) <= (layer4_outputs(2916)) and not (layer4_outputs(87));
    layer5_outputs(1651) <= not(layer4_outputs(427));
    layer5_outputs(1652) <= not((layer4_outputs(3598)) xor (layer4_outputs(4543)));
    layer5_outputs(1653) <= (layer4_outputs(1301)) and not (layer4_outputs(131));
    layer5_outputs(1654) <= not(layer4_outputs(3446));
    layer5_outputs(1655) <= not((layer4_outputs(4374)) and (layer4_outputs(2972)));
    layer5_outputs(1656) <= layer4_outputs(2455);
    layer5_outputs(1657) <= layer4_outputs(281);
    layer5_outputs(1658) <= not(layer4_outputs(3177));
    layer5_outputs(1659) <= (layer4_outputs(147)) xor (layer4_outputs(286));
    layer5_outputs(1660) <= layer4_outputs(4589);
    layer5_outputs(1661) <= layer4_outputs(3235);
    layer5_outputs(1662) <= (layer4_outputs(3100)) and not (layer4_outputs(665));
    layer5_outputs(1663) <= '0';
    layer5_outputs(1664) <= not(layer4_outputs(4838));
    layer5_outputs(1665) <= layer4_outputs(697);
    layer5_outputs(1666) <= layer4_outputs(2255);
    layer5_outputs(1667) <= not(layer4_outputs(4323)) or (layer4_outputs(4255));
    layer5_outputs(1668) <= not(layer4_outputs(1883)) or (layer4_outputs(3732));
    layer5_outputs(1669) <= (layer4_outputs(789)) or (layer4_outputs(3093));
    layer5_outputs(1670) <= not(layer4_outputs(2005)) or (layer4_outputs(250));
    layer5_outputs(1671) <= layer4_outputs(2428);
    layer5_outputs(1672) <= '0';
    layer5_outputs(1673) <= not((layer4_outputs(2012)) or (layer4_outputs(2906)));
    layer5_outputs(1674) <= not(layer4_outputs(2090));
    layer5_outputs(1675) <= '1';
    layer5_outputs(1676) <= layer4_outputs(1139);
    layer5_outputs(1677) <= layer4_outputs(2146);
    layer5_outputs(1678) <= layer4_outputs(22);
    layer5_outputs(1679) <= not(layer4_outputs(803));
    layer5_outputs(1680) <= layer4_outputs(550);
    layer5_outputs(1681) <= not(layer4_outputs(4273)) or (layer4_outputs(4391));
    layer5_outputs(1682) <= '0';
    layer5_outputs(1683) <= not(layer4_outputs(2012));
    layer5_outputs(1684) <= not(layer4_outputs(1412));
    layer5_outputs(1685) <= not(layer4_outputs(3015));
    layer5_outputs(1686) <= (layer4_outputs(4464)) and (layer4_outputs(2234));
    layer5_outputs(1687) <= (layer4_outputs(4361)) and not (layer4_outputs(105));
    layer5_outputs(1688) <= not((layer4_outputs(1411)) and (layer4_outputs(4408)));
    layer5_outputs(1689) <= not(layer4_outputs(3821)) or (layer4_outputs(36));
    layer5_outputs(1690) <= (layer4_outputs(4549)) xor (layer4_outputs(1382));
    layer5_outputs(1691) <= not(layer4_outputs(817)) or (layer4_outputs(4365));
    layer5_outputs(1692) <= (layer4_outputs(388)) or (layer4_outputs(2990));
    layer5_outputs(1693) <= (layer4_outputs(3002)) or (layer4_outputs(2809));
    layer5_outputs(1694) <= not(layer4_outputs(1298)) or (layer4_outputs(4528));
    layer5_outputs(1695) <= not(layer4_outputs(2676));
    layer5_outputs(1696) <= not(layer4_outputs(985)) or (layer4_outputs(1816));
    layer5_outputs(1697) <= '0';
    layer5_outputs(1698) <= (layer4_outputs(2035)) or (layer4_outputs(3700));
    layer5_outputs(1699) <= '0';
    layer5_outputs(1700) <= (layer4_outputs(4433)) and not (layer4_outputs(737));
    layer5_outputs(1701) <= (layer4_outputs(3001)) and not (layer4_outputs(3577));
    layer5_outputs(1702) <= not(layer4_outputs(1145));
    layer5_outputs(1703) <= not((layer4_outputs(2322)) and (layer4_outputs(781)));
    layer5_outputs(1704) <= '1';
    layer5_outputs(1705) <= not(layer4_outputs(4872));
    layer5_outputs(1706) <= (layer4_outputs(221)) and not (layer4_outputs(2798));
    layer5_outputs(1707) <= not(layer4_outputs(139));
    layer5_outputs(1708) <= not(layer4_outputs(1751));
    layer5_outputs(1709) <= '0';
    layer5_outputs(1710) <= layer4_outputs(320);
    layer5_outputs(1711) <= (layer4_outputs(655)) and (layer4_outputs(3950));
    layer5_outputs(1712) <= not(layer4_outputs(3711));
    layer5_outputs(1713) <= layer4_outputs(1741);
    layer5_outputs(1714) <= layer4_outputs(3465);
    layer5_outputs(1715) <= (layer4_outputs(481)) and (layer4_outputs(3616));
    layer5_outputs(1716) <= not(layer4_outputs(1672)) or (layer4_outputs(43));
    layer5_outputs(1717) <= not(layer4_outputs(3398));
    layer5_outputs(1718) <= layer4_outputs(3271);
    layer5_outputs(1719) <= not(layer4_outputs(3996));
    layer5_outputs(1720) <= not(layer4_outputs(4539)) or (layer4_outputs(4194));
    layer5_outputs(1721) <= layer4_outputs(4706);
    layer5_outputs(1722) <= not((layer4_outputs(4192)) or (layer4_outputs(340)));
    layer5_outputs(1723) <= not(layer4_outputs(2914)) or (layer4_outputs(4602));
    layer5_outputs(1724) <= (layer4_outputs(1178)) or (layer4_outputs(4159));
    layer5_outputs(1725) <= '0';
    layer5_outputs(1726) <= not(layer4_outputs(1792)) or (layer4_outputs(4016));
    layer5_outputs(1727) <= layer4_outputs(4035);
    layer5_outputs(1728) <= (layer4_outputs(3293)) and not (layer4_outputs(38));
    layer5_outputs(1729) <= '1';
    layer5_outputs(1730) <= (layer4_outputs(2801)) and not (layer4_outputs(1664));
    layer5_outputs(1731) <= (layer4_outputs(1897)) and (layer4_outputs(4904));
    layer5_outputs(1732) <= layer4_outputs(18);
    layer5_outputs(1733) <= not(layer4_outputs(2109));
    layer5_outputs(1734) <= '1';
    layer5_outputs(1735) <= not(layer4_outputs(4581));
    layer5_outputs(1736) <= not(layer4_outputs(4636)) or (layer4_outputs(2876));
    layer5_outputs(1737) <= layer4_outputs(4807);
    layer5_outputs(1738) <= not(layer4_outputs(1281));
    layer5_outputs(1739) <= (layer4_outputs(3726)) or (layer4_outputs(1257));
    layer5_outputs(1740) <= '1';
    layer5_outputs(1741) <= not(layer4_outputs(4918));
    layer5_outputs(1742) <= (layer4_outputs(2201)) or (layer4_outputs(3877));
    layer5_outputs(1743) <= not(layer4_outputs(963));
    layer5_outputs(1744) <= not((layer4_outputs(3544)) and (layer4_outputs(1431)));
    layer5_outputs(1745) <= not(layer4_outputs(3386)) or (layer4_outputs(4757));
    layer5_outputs(1746) <= not(layer4_outputs(1854)) or (layer4_outputs(3498));
    layer5_outputs(1747) <= not((layer4_outputs(935)) xor (layer4_outputs(4382)));
    layer5_outputs(1748) <= not(layer4_outputs(111));
    layer5_outputs(1749) <= not(layer4_outputs(4248));
    layer5_outputs(1750) <= layer4_outputs(559);
    layer5_outputs(1751) <= not((layer4_outputs(2116)) and (layer4_outputs(4357)));
    layer5_outputs(1752) <= (layer4_outputs(522)) and not (layer4_outputs(2441));
    layer5_outputs(1753) <= '0';
    layer5_outputs(1754) <= (layer4_outputs(960)) and not (layer4_outputs(2364));
    layer5_outputs(1755) <= (layer4_outputs(2851)) and not (layer4_outputs(1795));
    layer5_outputs(1756) <= not(layer4_outputs(3791));
    layer5_outputs(1757) <= layer4_outputs(2376);
    layer5_outputs(1758) <= '1';
    layer5_outputs(1759) <= not(layer4_outputs(4708));
    layer5_outputs(1760) <= not(layer4_outputs(3167));
    layer5_outputs(1761) <= not((layer4_outputs(5101)) or (layer4_outputs(2931)));
    layer5_outputs(1762) <= layer4_outputs(1371);
    layer5_outputs(1763) <= layer4_outputs(3820);
    layer5_outputs(1764) <= layer4_outputs(4737);
    layer5_outputs(1765) <= not((layer4_outputs(1034)) or (layer4_outputs(4325)));
    layer5_outputs(1766) <= '1';
    layer5_outputs(1767) <= not(layer4_outputs(2842));
    layer5_outputs(1768) <= not(layer4_outputs(2717)) or (layer4_outputs(764));
    layer5_outputs(1769) <= (layer4_outputs(2595)) and not (layer4_outputs(498));
    layer5_outputs(1770) <= not(layer4_outputs(1170));
    layer5_outputs(1771) <= not(layer4_outputs(3170));
    layer5_outputs(1772) <= not(layer4_outputs(1079));
    layer5_outputs(1773) <= layer4_outputs(4456);
    layer5_outputs(1774) <= layer4_outputs(1569);
    layer5_outputs(1775) <= '0';
    layer5_outputs(1776) <= layer4_outputs(5093);
    layer5_outputs(1777) <= layer4_outputs(2871);
    layer5_outputs(1778) <= (layer4_outputs(4250)) and not (layer4_outputs(3624));
    layer5_outputs(1779) <= (layer4_outputs(3147)) and (layer4_outputs(2488));
    layer5_outputs(1780) <= layer4_outputs(2486);
    layer5_outputs(1781) <= layer4_outputs(124);
    layer5_outputs(1782) <= (layer4_outputs(1164)) and (layer4_outputs(2164));
    layer5_outputs(1783) <= not(layer4_outputs(2921));
    layer5_outputs(1784) <= not(layer4_outputs(5020));
    layer5_outputs(1785) <= '0';
    layer5_outputs(1786) <= layer4_outputs(1025);
    layer5_outputs(1787) <= not(layer4_outputs(2674));
    layer5_outputs(1788) <= (layer4_outputs(3030)) and not (layer4_outputs(1984));
    layer5_outputs(1789) <= not(layer4_outputs(4168)) or (layer4_outputs(2502));
    layer5_outputs(1790) <= not(layer4_outputs(2396));
    layer5_outputs(1791) <= '1';
    layer5_outputs(1792) <= not((layer4_outputs(1389)) and (layer4_outputs(4039)));
    layer5_outputs(1793) <= layer4_outputs(2875);
    layer5_outputs(1794) <= layer4_outputs(4832);
    layer5_outputs(1795) <= (layer4_outputs(3885)) and not (layer4_outputs(4127));
    layer5_outputs(1796) <= not((layer4_outputs(3527)) xor (layer4_outputs(2021)));
    layer5_outputs(1797) <= not((layer4_outputs(724)) or (layer4_outputs(1062)));
    layer5_outputs(1798) <= layer4_outputs(4467);
    layer5_outputs(1799) <= '0';
    layer5_outputs(1800) <= layer4_outputs(128);
    layer5_outputs(1801) <= not(layer4_outputs(4457));
    layer5_outputs(1802) <= '0';
    layer5_outputs(1803) <= layer4_outputs(1854);
    layer5_outputs(1804) <= layer4_outputs(1927);
    layer5_outputs(1805) <= not((layer4_outputs(4873)) and (layer4_outputs(4988)));
    layer5_outputs(1806) <= layer4_outputs(5077);
    layer5_outputs(1807) <= not(layer4_outputs(5023));
    layer5_outputs(1808) <= layer4_outputs(2693);
    layer5_outputs(1809) <= (layer4_outputs(4520)) and not (layer4_outputs(4989));
    layer5_outputs(1810) <= (layer4_outputs(3890)) and not (layer4_outputs(907));
    layer5_outputs(1811) <= not(layer4_outputs(3016));
    layer5_outputs(1812) <= not(layer4_outputs(4595)) or (layer4_outputs(932));
    layer5_outputs(1813) <= '1';
    layer5_outputs(1814) <= '1';
    layer5_outputs(1815) <= not(layer4_outputs(3536)) or (layer4_outputs(711));
    layer5_outputs(1816) <= '1';
    layer5_outputs(1817) <= (layer4_outputs(2584)) and not (layer4_outputs(3726));
    layer5_outputs(1818) <= not(layer4_outputs(227));
    layer5_outputs(1819) <= (layer4_outputs(1725)) and (layer4_outputs(1970));
    layer5_outputs(1820) <= not(layer4_outputs(370));
    layer5_outputs(1821) <= '1';
    layer5_outputs(1822) <= '1';
    layer5_outputs(1823) <= layer4_outputs(1744);
    layer5_outputs(1824) <= not((layer4_outputs(2120)) and (layer4_outputs(2214)));
    layer5_outputs(1825) <= layer4_outputs(2158);
    layer5_outputs(1826) <= '1';
    layer5_outputs(1827) <= not(layer4_outputs(1004)) or (layer4_outputs(3453));
    layer5_outputs(1828) <= (layer4_outputs(4761)) and not (layer4_outputs(2415));
    layer5_outputs(1829) <= '0';
    layer5_outputs(1830) <= not(layer4_outputs(863)) or (layer4_outputs(3465));
    layer5_outputs(1831) <= (layer4_outputs(12)) and (layer4_outputs(4625));
    layer5_outputs(1832) <= (layer4_outputs(323)) and not (layer4_outputs(3772));
    layer5_outputs(1833) <= (layer4_outputs(3053)) and not (layer4_outputs(1990));
    layer5_outputs(1834) <= not((layer4_outputs(1218)) or (layer4_outputs(49)));
    layer5_outputs(1835) <= layer4_outputs(1570);
    layer5_outputs(1836) <= not(layer4_outputs(80));
    layer5_outputs(1837) <= not(layer4_outputs(1144));
    layer5_outputs(1838) <= '0';
    layer5_outputs(1839) <= not(layer4_outputs(2582)) or (layer4_outputs(898));
    layer5_outputs(1840) <= '0';
    layer5_outputs(1841) <= layer4_outputs(103);
    layer5_outputs(1842) <= not((layer4_outputs(2984)) and (layer4_outputs(3742)));
    layer5_outputs(1843) <= (layer4_outputs(4931)) and (layer4_outputs(1995));
    layer5_outputs(1844) <= (layer4_outputs(1340)) or (layer4_outputs(4080));
    layer5_outputs(1845) <= (layer4_outputs(824)) and (layer4_outputs(3198));
    layer5_outputs(1846) <= layer4_outputs(1873);
    layer5_outputs(1847) <= '1';
    layer5_outputs(1848) <= not(layer4_outputs(1012)) or (layer4_outputs(2439));
    layer5_outputs(1849) <= not((layer4_outputs(3661)) xor (layer4_outputs(2067)));
    layer5_outputs(1850) <= not(layer4_outputs(2781));
    layer5_outputs(1851) <= not(layer4_outputs(3960));
    layer5_outputs(1852) <= (layer4_outputs(4195)) or (layer4_outputs(1033));
    layer5_outputs(1853) <= '0';
    layer5_outputs(1854) <= (layer4_outputs(285)) or (layer4_outputs(1178));
    layer5_outputs(1855) <= layer4_outputs(3987);
    layer5_outputs(1856) <= (layer4_outputs(1585)) and (layer4_outputs(4219));
    layer5_outputs(1857) <= not(layer4_outputs(723));
    layer5_outputs(1858) <= layer4_outputs(2372);
    layer5_outputs(1859) <= (layer4_outputs(5100)) xor (layer4_outputs(3856));
    layer5_outputs(1860) <= (layer4_outputs(600)) and not (layer4_outputs(411));
    layer5_outputs(1861) <= not(layer4_outputs(1460));
    layer5_outputs(1862) <= layer4_outputs(2858);
    layer5_outputs(1863) <= '0';
    layer5_outputs(1864) <= (layer4_outputs(1746)) and (layer4_outputs(4695));
    layer5_outputs(1865) <= layer4_outputs(2747);
    layer5_outputs(1866) <= '0';
    layer5_outputs(1867) <= not(layer4_outputs(1367));
    layer5_outputs(1868) <= layer4_outputs(4316);
    layer5_outputs(1869) <= not((layer4_outputs(3496)) and (layer4_outputs(2031)));
    layer5_outputs(1870) <= (layer4_outputs(1615)) and not (layer4_outputs(1861));
    layer5_outputs(1871) <= (layer4_outputs(843)) or (layer4_outputs(2527));
    layer5_outputs(1872) <= not(layer4_outputs(190)) or (layer4_outputs(4292));
    layer5_outputs(1873) <= '1';
    layer5_outputs(1874) <= (layer4_outputs(2306)) or (layer4_outputs(4115));
    layer5_outputs(1875) <= not(layer4_outputs(4962));
    layer5_outputs(1876) <= layer4_outputs(1834);
    layer5_outputs(1877) <= not((layer4_outputs(2813)) xor (layer4_outputs(900)));
    layer5_outputs(1878) <= (layer4_outputs(3266)) and not (layer4_outputs(1143));
    layer5_outputs(1879) <= not(layer4_outputs(4366)) or (layer4_outputs(3417));
    layer5_outputs(1880) <= not(layer4_outputs(1826));
    layer5_outputs(1881) <= (layer4_outputs(896)) or (layer4_outputs(3319));
    layer5_outputs(1882) <= not(layer4_outputs(407));
    layer5_outputs(1883) <= not(layer4_outputs(2085)) or (layer4_outputs(2426));
    layer5_outputs(1884) <= not(layer4_outputs(2100)) or (layer4_outputs(340));
    layer5_outputs(1885) <= not(layer4_outputs(1685));
    layer5_outputs(1886) <= layer4_outputs(3561);
    layer5_outputs(1887) <= layer4_outputs(208);
    layer5_outputs(1888) <= (layer4_outputs(1705)) and not (layer4_outputs(4645));
    layer5_outputs(1889) <= not((layer4_outputs(193)) and (layer4_outputs(2660)));
    layer5_outputs(1890) <= '0';
    layer5_outputs(1891) <= not(layer4_outputs(1920));
    layer5_outputs(1892) <= not(layer4_outputs(3751));
    layer5_outputs(1893) <= (layer4_outputs(3498)) and (layer4_outputs(3139));
    layer5_outputs(1894) <= not((layer4_outputs(3012)) and (layer4_outputs(4986)));
    layer5_outputs(1895) <= not((layer4_outputs(2147)) xor (layer4_outputs(1701)));
    layer5_outputs(1896) <= not(layer4_outputs(989)) or (layer4_outputs(837));
    layer5_outputs(1897) <= '1';
    layer5_outputs(1898) <= not(layer4_outputs(595));
    layer5_outputs(1899) <= not(layer4_outputs(373)) or (layer4_outputs(3036));
    layer5_outputs(1900) <= (layer4_outputs(5022)) or (layer4_outputs(422));
    layer5_outputs(1901) <= not(layer4_outputs(1103)) or (layer4_outputs(324));
    layer5_outputs(1902) <= (layer4_outputs(2397)) and (layer4_outputs(1628));
    layer5_outputs(1903) <= not(layer4_outputs(3018)) or (layer4_outputs(1852));
    layer5_outputs(1904) <= '0';
    layer5_outputs(1905) <= not(layer4_outputs(1391));
    layer5_outputs(1906) <= not(layer4_outputs(2078));
    layer5_outputs(1907) <= (layer4_outputs(4554)) and not (layer4_outputs(2881));
    layer5_outputs(1908) <= '0';
    layer5_outputs(1909) <= (layer4_outputs(3914)) and (layer4_outputs(1781));
    layer5_outputs(1910) <= (layer4_outputs(3430)) and not (layer4_outputs(4673));
    layer5_outputs(1911) <= not(layer4_outputs(2435)) or (layer4_outputs(664));
    layer5_outputs(1912) <= not(layer4_outputs(3014));
    layer5_outputs(1913) <= (layer4_outputs(139)) and not (layer4_outputs(439));
    layer5_outputs(1914) <= layer4_outputs(1342);
    layer5_outputs(1915) <= not(layer4_outputs(4782));
    layer5_outputs(1916) <= layer4_outputs(2490);
    layer5_outputs(1917) <= '1';
    layer5_outputs(1918) <= not(layer4_outputs(4956));
    layer5_outputs(1919) <= layer4_outputs(4626);
    layer5_outputs(1920) <= not((layer4_outputs(1988)) and (layer4_outputs(3147)));
    layer5_outputs(1921) <= not(layer4_outputs(2026)) or (layer4_outputs(876));
    layer5_outputs(1922) <= not((layer4_outputs(1078)) and (layer4_outputs(4789)));
    layer5_outputs(1923) <= (layer4_outputs(4358)) and (layer4_outputs(3300));
    layer5_outputs(1924) <= (layer4_outputs(2673)) and not (layer4_outputs(2878));
    layer5_outputs(1925) <= not(layer4_outputs(2369));
    layer5_outputs(1926) <= layer4_outputs(3607);
    layer5_outputs(1927) <= not((layer4_outputs(1188)) or (layer4_outputs(2668)));
    layer5_outputs(1928) <= layer4_outputs(3392);
    layer5_outputs(1929) <= layer4_outputs(4975);
    layer5_outputs(1930) <= not(layer4_outputs(4853)) or (layer4_outputs(210));
    layer5_outputs(1931) <= not(layer4_outputs(1058)) or (layer4_outputs(2336));
    layer5_outputs(1932) <= '0';
    layer5_outputs(1933) <= layer4_outputs(4337);
    layer5_outputs(1934) <= (layer4_outputs(1429)) and not (layer4_outputs(1519));
    layer5_outputs(1935) <= (layer4_outputs(2552)) and (layer4_outputs(3347));
    layer5_outputs(1936) <= (layer4_outputs(113)) and not (layer4_outputs(1893));
    layer5_outputs(1937) <= not(layer4_outputs(2933)) or (layer4_outputs(1818));
    layer5_outputs(1938) <= not(layer4_outputs(1619));
    layer5_outputs(1939) <= '0';
    layer5_outputs(1940) <= '0';
    layer5_outputs(1941) <= (layer4_outputs(2498)) and (layer4_outputs(1601));
    layer5_outputs(1942) <= (layer4_outputs(2938)) and not (layer4_outputs(3138));
    layer5_outputs(1943) <= layer4_outputs(3609);
    layer5_outputs(1944) <= not(layer4_outputs(1295)) or (layer4_outputs(2679));
    layer5_outputs(1945) <= (layer4_outputs(4862)) and (layer4_outputs(1424));
    layer5_outputs(1946) <= not(layer4_outputs(4661));
    layer5_outputs(1947) <= not(layer4_outputs(2861)) or (layer4_outputs(4376));
    layer5_outputs(1948) <= not(layer4_outputs(1262));
    layer5_outputs(1949) <= (layer4_outputs(471)) and not (layer4_outputs(981));
    layer5_outputs(1950) <= layer4_outputs(4525);
    layer5_outputs(1951) <= layer4_outputs(1061);
    layer5_outputs(1952) <= not(layer4_outputs(2693));
    layer5_outputs(1953) <= not((layer4_outputs(1761)) or (layer4_outputs(2208)));
    layer5_outputs(1954) <= not(layer4_outputs(533));
    layer5_outputs(1955) <= layer4_outputs(1648);
    layer5_outputs(1956) <= layer4_outputs(2777);
    layer5_outputs(1957) <= (layer4_outputs(3281)) and (layer4_outputs(2089));
    layer5_outputs(1958) <= not(layer4_outputs(1718)) or (layer4_outputs(409));
    layer5_outputs(1959) <= not(layer4_outputs(2686));
    layer5_outputs(1960) <= not((layer4_outputs(4333)) and (layer4_outputs(2840)));
    layer5_outputs(1961) <= not(layer4_outputs(3599)) or (layer4_outputs(34));
    layer5_outputs(1962) <= not((layer4_outputs(218)) and (layer4_outputs(4332)));
    layer5_outputs(1963) <= not(layer4_outputs(2763));
    layer5_outputs(1964) <= (layer4_outputs(5078)) and not (layer4_outputs(3830));
    layer5_outputs(1965) <= not(layer4_outputs(4849)) or (layer4_outputs(196));
    layer5_outputs(1966) <= not(layer4_outputs(277)) or (layer4_outputs(4106));
    layer5_outputs(1967) <= not(layer4_outputs(1439)) or (layer4_outputs(2493));
    layer5_outputs(1968) <= (layer4_outputs(1290)) or (layer4_outputs(4553));
    layer5_outputs(1969) <= layer4_outputs(3094);
    layer5_outputs(1970) <= not(layer4_outputs(3897));
    layer5_outputs(1971) <= layer4_outputs(1556);
    layer5_outputs(1972) <= not(layer4_outputs(1022));
    layer5_outputs(1973) <= '1';
    layer5_outputs(1974) <= (layer4_outputs(4600)) and not (layer4_outputs(1885));
    layer5_outputs(1975) <= layer4_outputs(4943);
    layer5_outputs(1976) <= not(layer4_outputs(5029));
    layer5_outputs(1977) <= not(layer4_outputs(1154)) or (layer4_outputs(4879));
    layer5_outputs(1978) <= not(layer4_outputs(2807));
    layer5_outputs(1979) <= layer4_outputs(3092);
    layer5_outputs(1980) <= not(layer4_outputs(1655)) or (layer4_outputs(2555));
    layer5_outputs(1981) <= layer4_outputs(415);
    layer5_outputs(1982) <= '0';
    layer5_outputs(1983) <= (layer4_outputs(3478)) and (layer4_outputs(3179));
    layer5_outputs(1984) <= layer4_outputs(2353);
    layer5_outputs(1985) <= (layer4_outputs(4274)) xor (layer4_outputs(1840));
    layer5_outputs(1986) <= not(layer4_outputs(3878)) or (layer4_outputs(3055));
    layer5_outputs(1987) <= (layer4_outputs(2819)) and not (layer4_outputs(2051));
    layer5_outputs(1988) <= not(layer4_outputs(2975));
    layer5_outputs(1989) <= layer4_outputs(350);
    layer5_outputs(1990) <= not((layer4_outputs(2329)) or (layer4_outputs(1090)));
    layer5_outputs(1991) <= (layer4_outputs(3805)) and not (layer4_outputs(4581));
    layer5_outputs(1992) <= layer4_outputs(3945);
    layer5_outputs(1993) <= layer4_outputs(2429);
    layer5_outputs(1994) <= not(layer4_outputs(3164));
    layer5_outputs(1995) <= layer4_outputs(5064);
    layer5_outputs(1996) <= not(layer4_outputs(4575));
    layer5_outputs(1997) <= (layer4_outputs(4763)) and not (layer4_outputs(3025));
    layer5_outputs(1998) <= not(layer4_outputs(1555));
    layer5_outputs(1999) <= (layer4_outputs(1707)) xor (layer4_outputs(1663));
    layer5_outputs(2000) <= (layer4_outputs(2102)) and not (layer4_outputs(3722));
    layer5_outputs(2001) <= (layer4_outputs(643)) and not (layer4_outputs(3490));
    layer5_outputs(2002) <= not(layer4_outputs(3277));
    layer5_outputs(2003) <= not(layer4_outputs(4045)) or (layer4_outputs(2783));
    layer5_outputs(2004) <= not((layer4_outputs(403)) or (layer4_outputs(2087)));
    layer5_outputs(2005) <= not(layer4_outputs(3098));
    layer5_outputs(2006) <= '1';
    layer5_outputs(2007) <= (layer4_outputs(4162)) and not (layer4_outputs(3821));
    layer5_outputs(2008) <= not((layer4_outputs(2932)) and (layer4_outputs(772)));
    layer5_outputs(2009) <= not(layer4_outputs(4249));
    layer5_outputs(2010) <= (layer4_outputs(984)) and not (layer4_outputs(1310));
    layer5_outputs(2011) <= not(layer4_outputs(2013)) or (layer4_outputs(2634));
    layer5_outputs(2012) <= (layer4_outputs(3679)) and (layer4_outputs(3755));
    layer5_outputs(2013) <= not(layer4_outputs(1354)) or (layer4_outputs(1139));
    layer5_outputs(2014) <= layer4_outputs(1194);
    layer5_outputs(2015) <= not(layer4_outputs(2455)) or (layer4_outputs(1307));
    layer5_outputs(2016) <= layer4_outputs(2345);
    layer5_outputs(2017) <= (layer4_outputs(1074)) and not (layer4_outputs(4037));
    layer5_outputs(2018) <= layer4_outputs(4154);
    layer5_outputs(2019) <= (layer4_outputs(507)) and (layer4_outputs(3899));
    layer5_outputs(2020) <= (layer4_outputs(2499)) and not (layer4_outputs(3064));
    layer5_outputs(2021) <= '0';
    layer5_outputs(2022) <= not(layer4_outputs(5022)) or (layer4_outputs(3538));
    layer5_outputs(2023) <= layer4_outputs(363);
    layer5_outputs(2024) <= layer4_outputs(1131);
    layer5_outputs(2025) <= not(layer4_outputs(1352)) or (layer4_outputs(2398));
    layer5_outputs(2026) <= not((layer4_outputs(3749)) and (layer4_outputs(4901)));
    layer5_outputs(2027) <= layer4_outputs(664);
    layer5_outputs(2028) <= (layer4_outputs(832)) and (layer4_outputs(3040));
    layer5_outputs(2029) <= not((layer4_outputs(3681)) or (layer4_outputs(2558)));
    layer5_outputs(2030) <= not(layer4_outputs(2126));
    layer5_outputs(2031) <= not(layer4_outputs(1917));
    layer5_outputs(2032) <= not(layer4_outputs(3443));
    layer5_outputs(2033) <= '1';
    layer5_outputs(2034) <= not(layer4_outputs(240));
    layer5_outputs(2035) <= layer4_outputs(3405);
    layer5_outputs(2036) <= not(layer4_outputs(4518));
    layer5_outputs(2037) <= not(layer4_outputs(3851)) or (layer4_outputs(1867));
    layer5_outputs(2038) <= '0';
    layer5_outputs(2039) <= (layer4_outputs(1978)) and not (layer4_outputs(4995));
    layer5_outputs(2040) <= (layer4_outputs(4680)) and not (layer4_outputs(2136));
    layer5_outputs(2041) <= not(layer4_outputs(1800)) or (layer4_outputs(640));
    layer5_outputs(2042) <= not(layer4_outputs(4072)) or (layer4_outputs(1445));
    layer5_outputs(2043) <= not(layer4_outputs(1401));
    layer5_outputs(2044) <= (layer4_outputs(1758)) or (layer4_outputs(1189));
    layer5_outputs(2045) <= (layer4_outputs(192)) and not (layer4_outputs(1755));
    layer5_outputs(2046) <= not(layer4_outputs(4087)) or (layer4_outputs(2295));
    layer5_outputs(2047) <= not(layer4_outputs(3125)) or (layer4_outputs(3792));
    layer5_outputs(2048) <= layer4_outputs(2576);
    layer5_outputs(2049) <= not(layer4_outputs(1931)) or (layer4_outputs(800));
    layer5_outputs(2050) <= not(layer4_outputs(675)) or (layer4_outputs(4013));
    layer5_outputs(2051) <= (layer4_outputs(2490)) xor (layer4_outputs(1355));
    layer5_outputs(2052) <= not(layer4_outputs(3733));
    layer5_outputs(2053) <= layer4_outputs(2267);
    layer5_outputs(2054) <= layer4_outputs(5037);
    layer5_outputs(2055) <= layer4_outputs(2294);
    layer5_outputs(2056) <= not(layer4_outputs(2966));
    layer5_outputs(2057) <= not((layer4_outputs(1563)) and (layer4_outputs(3422)));
    layer5_outputs(2058) <= not(layer4_outputs(3212)) or (layer4_outputs(269));
    layer5_outputs(2059) <= '0';
    layer5_outputs(2060) <= '1';
    layer5_outputs(2061) <= not(layer4_outputs(341));
    layer5_outputs(2062) <= not(layer4_outputs(4262)) or (layer4_outputs(3883));
    layer5_outputs(2063) <= '0';
    layer5_outputs(2064) <= not(layer4_outputs(5071)) or (layer4_outputs(3594));
    layer5_outputs(2065) <= (layer4_outputs(1517)) xor (layer4_outputs(3142));
    layer5_outputs(2066) <= not((layer4_outputs(4479)) xor (layer4_outputs(4501)));
    layer5_outputs(2067) <= (layer4_outputs(4191)) and (layer4_outputs(4069));
    layer5_outputs(2068) <= not(layer4_outputs(2887));
    layer5_outputs(2069) <= (layer4_outputs(2533)) or (layer4_outputs(2903));
    layer5_outputs(2070) <= not(layer4_outputs(1803));
    layer5_outputs(2071) <= (layer4_outputs(768)) and (layer4_outputs(4107));
    layer5_outputs(2072) <= not((layer4_outputs(3084)) and (layer4_outputs(2460)));
    layer5_outputs(2073) <= layer4_outputs(2365);
    layer5_outputs(2074) <= not(layer4_outputs(766));
    layer5_outputs(2075) <= (layer4_outputs(26)) xor (layer4_outputs(4394));
    layer5_outputs(2076) <= layer4_outputs(4485);
    layer5_outputs(2077) <= (layer4_outputs(3896)) or (layer4_outputs(1264));
    layer5_outputs(2078) <= layer4_outputs(2566);
    layer5_outputs(2079) <= '1';
    layer5_outputs(2080) <= '0';
    layer5_outputs(2081) <= (layer4_outputs(4421)) xor (layer4_outputs(457));
    layer5_outputs(2082) <= not(layer4_outputs(703));
    layer5_outputs(2083) <= layer4_outputs(3399);
    layer5_outputs(2084) <= not(layer4_outputs(1830));
    layer5_outputs(2085) <= not((layer4_outputs(2180)) xor (layer4_outputs(2004)));
    layer5_outputs(2086) <= not((layer4_outputs(1791)) and (layer4_outputs(739)));
    layer5_outputs(2087) <= (layer4_outputs(1720)) xor (layer4_outputs(2115));
    layer5_outputs(2088) <= (layer4_outputs(2526)) xor (layer4_outputs(410));
    layer5_outputs(2089) <= (layer4_outputs(928)) and (layer4_outputs(761));
    layer5_outputs(2090) <= not((layer4_outputs(4208)) or (layer4_outputs(682)));
    layer5_outputs(2091) <= layer4_outputs(3867);
    layer5_outputs(2092) <= layer4_outputs(1811);
    layer5_outputs(2093) <= not(layer4_outputs(35)) or (layer4_outputs(3819));
    layer5_outputs(2094) <= layer4_outputs(3103);
    layer5_outputs(2095) <= layer4_outputs(282);
    layer5_outputs(2096) <= (layer4_outputs(1656)) and (layer4_outputs(4021));
    layer5_outputs(2097) <= not((layer4_outputs(4647)) and (layer4_outputs(771)));
    layer5_outputs(2098) <= layer4_outputs(709);
    layer5_outputs(2099) <= (layer4_outputs(3889)) and not (layer4_outputs(4623));
    layer5_outputs(2100) <= layer4_outputs(2626);
    layer5_outputs(2101) <= not((layer4_outputs(1164)) or (layer4_outputs(2503)));
    layer5_outputs(2102) <= not(layer4_outputs(3300));
    layer5_outputs(2103) <= (layer4_outputs(1582)) and (layer4_outputs(454));
    layer5_outputs(2104) <= not((layer4_outputs(4478)) and (layer4_outputs(1384)));
    layer5_outputs(2105) <= (layer4_outputs(2442)) and not (layer4_outputs(143));
    layer5_outputs(2106) <= not(layer4_outputs(4948));
    layer5_outputs(2107) <= (layer4_outputs(4093)) and not (layer4_outputs(1756));
    layer5_outputs(2108) <= (layer4_outputs(839)) xor (layer4_outputs(3977));
    layer5_outputs(2109) <= not((layer4_outputs(4649)) and (layer4_outputs(914)));
    layer5_outputs(2110) <= not((layer4_outputs(3316)) xor (layer4_outputs(1185)));
    layer5_outputs(2111) <= (layer4_outputs(3812)) and not (layer4_outputs(1154));
    layer5_outputs(2112) <= (layer4_outputs(4921)) or (layer4_outputs(2244));
    layer5_outputs(2113) <= layer4_outputs(2134);
    layer5_outputs(2114) <= not(layer4_outputs(1993)) or (layer4_outputs(3169));
    layer5_outputs(2115) <= layer4_outputs(613);
    layer5_outputs(2116) <= layer4_outputs(1971);
    layer5_outputs(2117) <= (layer4_outputs(4636)) and (layer4_outputs(1692));
    layer5_outputs(2118) <= not(layer4_outputs(3279));
    layer5_outputs(2119) <= layer4_outputs(1565);
    layer5_outputs(2120) <= not((layer4_outputs(3520)) xor (layer4_outputs(4375)));
    layer5_outputs(2121) <= not(layer4_outputs(1590)) or (layer4_outputs(3169));
    layer5_outputs(2122) <= not(layer4_outputs(4271));
    layer5_outputs(2123) <= (layer4_outputs(3093)) or (layer4_outputs(4738));
    layer5_outputs(2124) <= not(layer4_outputs(4599));
    layer5_outputs(2125) <= not(layer4_outputs(2229));
    layer5_outputs(2126) <= not((layer4_outputs(4622)) xor (layer4_outputs(3421)));
    layer5_outputs(2127) <= (layer4_outputs(2849)) and not (layer4_outputs(1919));
    layer5_outputs(2128) <= not(layer4_outputs(4887)) or (layer4_outputs(2664));
    layer5_outputs(2129) <= layer4_outputs(3853);
    layer5_outputs(2130) <= (layer4_outputs(2630)) and (layer4_outputs(967));
    layer5_outputs(2131) <= (layer4_outputs(2197)) and (layer4_outputs(4215));
    layer5_outputs(2132) <= not((layer4_outputs(1628)) and (layer4_outputs(186)));
    layer5_outputs(2133) <= not((layer4_outputs(801)) or (layer4_outputs(432)));
    layer5_outputs(2134) <= not(layer4_outputs(3620)) or (layer4_outputs(4966));
    layer5_outputs(2135) <= not((layer4_outputs(3108)) xor (layer4_outputs(4647)));
    layer5_outputs(2136) <= (layer4_outputs(3780)) and (layer4_outputs(3797));
    layer5_outputs(2137) <= (layer4_outputs(1335)) or (layer4_outputs(3203));
    layer5_outputs(2138) <= (layer4_outputs(1549)) or (layer4_outputs(4341));
    layer5_outputs(2139) <= (layer4_outputs(1574)) and not (layer4_outputs(3974));
    layer5_outputs(2140) <= not((layer4_outputs(3019)) or (layer4_outputs(4587)));
    layer5_outputs(2141) <= layer4_outputs(2986);
    layer5_outputs(2142) <= '0';
    layer5_outputs(2143) <= (layer4_outputs(507)) xor (layer4_outputs(2749));
    layer5_outputs(2144) <= not(layer4_outputs(3647)) or (layer4_outputs(4592));
    layer5_outputs(2145) <= not(layer4_outputs(1964));
    layer5_outputs(2146) <= layer4_outputs(157);
    layer5_outputs(2147) <= (layer4_outputs(2963)) or (layer4_outputs(4512));
    layer5_outputs(2148) <= not((layer4_outputs(3894)) or (layer4_outputs(1467)));
    layer5_outputs(2149) <= '0';
    layer5_outputs(2150) <= (layer4_outputs(2017)) and (layer4_outputs(3395));
    layer5_outputs(2151) <= not((layer4_outputs(4475)) or (layer4_outputs(239)));
    layer5_outputs(2152) <= '0';
    layer5_outputs(2153) <= (layer4_outputs(790)) and not (layer4_outputs(3477));
    layer5_outputs(2154) <= layer4_outputs(5118);
    layer5_outputs(2155) <= (layer4_outputs(4681)) and not (layer4_outputs(1268));
    layer5_outputs(2156) <= not((layer4_outputs(3074)) and (layer4_outputs(1073)));
    layer5_outputs(2157) <= not(layer4_outputs(2179));
    layer5_outputs(2158) <= (layer4_outputs(5102)) and not (layer4_outputs(4448));
    layer5_outputs(2159) <= not(layer4_outputs(2181)) or (layer4_outputs(1491));
    layer5_outputs(2160) <= layer4_outputs(2800);
    layer5_outputs(2161) <= layer4_outputs(4073);
    layer5_outputs(2162) <= (layer4_outputs(4373)) or (layer4_outputs(2080));
    layer5_outputs(2163) <= not((layer4_outputs(4688)) or (layer4_outputs(596)));
    layer5_outputs(2164) <= not((layer4_outputs(3723)) or (layer4_outputs(3807)));
    layer5_outputs(2165) <= not(layer4_outputs(2223));
    layer5_outputs(2166) <= not(layer4_outputs(1966));
    layer5_outputs(2167) <= not(layer4_outputs(1398));
    layer5_outputs(2168) <= not(layer4_outputs(3495));
    layer5_outputs(2169) <= (layer4_outputs(2575)) or (layer4_outputs(5036));
    layer5_outputs(2170) <= not(layer4_outputs(763));
    layer5_outputs(2171) <= not((layer4_outputs(2500)) and (layer4_outputs(2144)));
    layer5_outputs(2172) <= layer4_outputs(4632);
    layer5_outputs(2173) <= not((layer4_outputs(5062)) xor (layer4_outputs(4045)));
    layer5_outputs(2174) <= not((layer4_outputs(924)) or (layer4_outputs(2743)));
    layer5_outputs(2175) <= not((layer4_outputs(2612)) and (layer4_outputs(4180)));
    layer5_outputs(2176) <= not((layer4_outputs(4455)) and (layer4_outputs(322)));
    layer5_outputs(2177) <= not((layer4_outputs(816)) or (layer4_outputs(2764)));
    layer5_outputs(2178) <= layer4_outputs(4842);
    layer5_outputs(2179) <= not(layer4_outputs(988));
    layer5_outputs(2180) <= (layer4_outputs(3937)) and not (layer4_outputs(5064));
    layer5_outputs(2181) <= (layer4_outputs(2875)) and (layer4_outputs(4954));
    layer5_outputs(2182) <= not(layer4_outputs(1111));
    layer5_outputs(2183) <= not((layer4_outputs(3162)) and (layer4_outputs(4840)));
    layer5_outputs(2184) <= not(layer4_outputs(4028));
    layer5_outputs(2185) <= not(layer4_outputs(4787)) or (layer4_outputs(3741));
    layer5_outputs(2186) <= (layer4_outputs(1637)) or (layer4_outputs(4283));
    layer5_outputs(2187) <= not(layer4_outputs(4958)) or (layer4_outputs(2525));
    layer5_outputs(2188) <= not(layer4_outputs(3091));
    layer5_outputs(2189) <= not(layer4_outputs(2110));
    layer5_outputs(2190) <= not(layer4_outputs(2528)) or (layer4_outputs(4237));
    layer5_outputs(2191) <= not(layer4_outputs(3699)) or (layer4_outputs(1297));
    layer5_outputs(2192) <= '1';
    layer5_outputs(2193) <= not((layer4_outputs(2537)) or (layer4_outputs(1682)));
    layer5_outputs(2194) <= (layer4_outputs(988)) and not (layer4_outputs(342));
    layer5_outputs(2195) <= layer4_outputs(557);
    layer5_outputs(2196) <= '0';
    layer5_outputs(2197) <= not(layer4_outputs(1197));
    layer5_outputs(2198) <= not(layer4_outputs(2585));
    layer5_outputs(2199) <= not(layer4_outputs(77)) or (layer4_outputs(3377));
    layer5_outputs(2200) <= '1';
    layer5_outputs(2201) <= not(layer4_outputs(4746)) or (layer4_outputs(4423));
    layer5_outputs(2202) <= not(layer4_outputs(2995));
    layer5_outputs(2203) <= '0';
    layer5_outputs(2204) <= not((layer4_outputs(673)) or (layer4_outputs(3409)));
    layer5_outputs(2205) <= (layer4_outputs(4521)) and not (layer4_outputs(4753));
    layer5_outputs(2206) <= not((layer4_outputs(3756)) or (layer4_outputs(904)));
    layer5_outputs(2207) <= '1';
    layer5_outputs(2208) <= (layer4_outputs(499)) xor (layer4_outputs(1463));
    layer5_outputs(2209) <= (layer4_outputs(5117)) and not (layer4_outputs(4273));
    layer5_outputs(2210) <= not(layer4_outputs(2245)) or (layer4_outputs(4363));
    layer5_outputs(2211) <= layer4_outputs(465);
    layer5_outputs(2212) <= not(layer4_outputs(41));
    layer5_outputs(2213) <= layer4_outputs(3506);
    layer5_outputs(2214) <= not(layer4_outputs(3263));
    layer5_outputs(2215) <= not(layer4_outputs(1503)) or (layer4_outputs(3628));
    layer5_outputs(2216) <= (layer4_outputs(1749)) or (layer4_outputs(2360));
    layer5_outputs(2217) <= layer4_outputs(576);
    layer5_outputs(2218) <= layer4_outputs(909);
    layer5_outputs(2219) <= '1';
    layer5_outputs(2220) <= '1';
    layer5_outputs(2221) <= not(layer4_outputs(1056));
    layer5_outputs(2222) <= layer4_outputs(1273);
    layer5_outputs(2223) <= layer4_outputs(3677);
    layer5_outputs(2224) <= (layer4_outputs(4298)) or (layer4_outputs(1191));
    layer5_outputs(2225) <= (layer4_outputs(4563)) xor (layer4_outputs(422));
    layer5_outputs(2226) <= not((layer4_outputs(729)) and (layer4_outputs(3329)));
    layer5_outputs(2227) <= not(layer4_outputs(2816)) or (layer4_outputs(215));
    layer5_outputs(2228) <= (layer4_outputs(4173)) and not (layer4_outputs(3932));
    layer5_outputs(2229) <= '1';
    layer5_outputs(2230) <= (layer4_outputs(2743)) and not (layer4_outputs(4654));
    layer5_outputs(2231) <= layer4_outputs(4677);
    layer5_outputs(2232) <= layer4_outputs(1967);
    layer5_outputs(2233) <= not((layer4_outputs(1643)) or (layer4_outputs(2050)));
    layer5_outputs(2234) <= (layer4_outputs(3924)) and not (layer4_outputs(1008));
    layer5_outputs(2235) <= not(layer4_outputs(591));
    layer5_outputs(2236) <= not(layer4_outputs(1818));
    layer5_outputs(2237) <= (layer4_outputs(474)) xor (layer4_outputs(2509));
    layer5_outputs(2238) <= not(layer4_outputs(5076));
    layer5_outputs(2239) <= not((layer4_outputs(4779)) xor (layer4_outputs(3444)));
    layer5_outputs(2240) <= not((layer4_outputs(4767)) or (layer4_outputs(2729)));
    layer5_outputs(2241) <= layer4_outputs(579);
    layer5_outputs(2242) <= not(layer4_outputs(4445));
    layer5_outputs(2243) <= not(layer4_outputs(2062)) or (layer4_outputs(5097));
    layer5_outputs(2244) <= not(layer4_outputs(4205));
    layer5_outputs(2245) <= not((layer4_outputs(465)) xor (layer4_outputs(2850)));
    layer5_outputs(2246) <= not(layer4_outputs(4439));
    layer5_outputs(2247) <= layer4_outputs(1763);
    layer5_outputs(2248) <= (layer4_outputs(3130)) and (layer4_outputs(2996));
    layer5_outputs(2249) <= not(layer4_outputs(2247));
    layer5_outputs(2250) <= not(layer4_outputs(3455));
    layer5_outputs(2251) <= not(layer4_outputs(1050)) or (layer4_outputs(1097));
    layer5_outputs(2252) <= not(layer4_outputs(3304)) or (layer4_outputs(2219));
    layer5_outputs(2253) <= (layer4_outputs(3031)) and not (layer4_outputs(2353));
    layer5_outputs(2254) <= layer4_outputs(3239);
    layer5_outputs(2255) <= not(layer4_outputs(1737));
    layer5_outputs(2256) <= (layer4_outputs(1465)) and not (layer4_outputs(423));
    layer5_outputs(2257) <= (layer4_outputs(2706)) and not (layer4_outputs(2402));
    layer5_outputs(2258) <= (layer4_outputs(1559)) or (layer4_outputs(4784));
    layer5_outputs(2259) <= (layer4_outputs(4114)) and (layer4_outputs(3341));
    layer5_outputs(2260) <= (layer4_outputs(3306)) and (layer4_outputs(1059));
    layer5_outputs(2261) <= not((layer4_outputs(1067)) xor (layer4_outputs(3762)));
    layer5_outputs(2262) <= (layer4_outputs(4732)) and not (layer4_outputs(3881));
    layer5_outputs(2263) <= not((layer4_outputs(619)) and (layer4_outputs(2803)));
    layer5_outputs(2264) <= (layer4_outputs(452)) and not (layer4_outputs(3771));
    layer5_outputs(2265) <= layer4_outputs(1885);
    layer5_outputs(2266) <= layer4_outputs(1627);
    layer5_outputs(2267) <= not(layer4_outputs(3560)) or (layer4_outputs(2404));
    layer5_outputs(2268) <= (layer4_outputs(180)) and not (layer4_outputs(2580));
    layer5_outputs(2269) <= not((layer4_outputs(4272)) or (layer4_outputs(2927)));
    layer5_outputs(2270) <= (layer4_outputs(3434)) and not (layer4_outputs(2696));
    layer5_outputs(2271) <= layer4_outputs(1750);
    layer5_outputs(2272) <= not((layer4_outputs(1138)) or (layer4_outputs(1955)));
    layer5_outputs(2273) <= layer4_outputs(3202);
    layer5_outputs(2274) <= (layer4_outputs(5103)) or (layer4_outputs(3564));
    layer5_outputs(2275) <= not(layer4_outputs(1099));
    layer5_outputs(2276) <= not((layer4_outputs(1291)) and (layer4_outputs(1626)));
    layer5_outputs(2277) <= (layer4_outputs(4332)) and not (layer4_outputs(1968));
    layer5_outputs(2278) <= not(layer4_outputs(1714));
    layer5_outputs(2279) <= (layer4_outputs(3444)) and not (layer4_outputs(2501));
    layer5_outputs(2280) <= not(layer4_outputs(2233)) or (layer4_outputs(343));
    layer5_outputs(2281) <= layer4_outputs(1648);
    layer5_outputs(2282) <= layer4_outputs(528);
    layer5_outputs(2283) <= not(layer4_outputs(3056));
    layer5_outputs(2284) <= not((layer4_outputs(2036)) and (layer4_outputs(3312)));
    layer5_outputs(2285) <= not(layer4_outputs(2140));
    layer5_outputs(2286) <= not(layer4_outputs(860)) or (layer4_outputs(1909));
    layer5_outputs(2287) <= (layer4_outputs(2313)) xor (layer4_outputs(2002));
    layer5_outputs(2288) <= not(layer4_outputs(2334)) or (layer4_outputs(4393));
    layer5_outputs(2289) <= layer4_outputs(1300);
    layer5_outputs(2290) <= not(layer4_outputs(1490)) or (layer4_outputs(3038));
    layer5_outputs(2291) <= layer4_outputs(2091);
    layer5_outputs(2292) <= not(layer4_outputs(1835)) or (layer4_outputs(3534));
    layer5_outputs(2293) <= not(layer4_outputs(3964));
    layer5_outputs(2294) <= not((layer4_outputs(1217)) and (layer4_outputs(4348)));
    layer5_outputs(2295) <= not((layer4_outputs(3698)) or (layer4_outputs(2808)));
    layer5_outputs(2296) <= not(layer4_outputs(3643));
    layer5_outputs(2297) <= not(layer4_outputs(807));
    layer5_outputs(2298) <= (layer4_outputs(3656)) xor (layer4_outputs(4429));
    layer5_outputs(2299) <= not(layer4_outputs(398)) or (layer4_outputs(1529));
    layer5_outputs(2300) <= (layer4_outputs(2976)) and not (layer4_outputs(458));
    layer5_outputs(2301) <= '0';
    layer5_outputs(2302) <= layer4_outputs(2911);
    layer5_outputs(2303) <= (layer4_outputs(4089)) and not (layer4_outputs(1908));
    layer5_outputs(2304) <= not(layer4_outputs(3721));
    layer5_outputs(2305) <= (layer4_outputs(4794)) and not (layer4_outputs(2242));
    layer5_outputs(2306) <= not(layer4_outputs(559));
    layer5_outputs(2307) <= not(layer4_outputs(4605));
    layer5_outputs(2308) <= not(layer4_outputs(3302));
    layer5_outputs(2309) <= not(layer4_outputs(2535));
    layer5_outputs(2310) <= not(layer4_outputs(1766));
    layer5_outputs(2311) <= not(layer4_outputs(797)) or (layer4_outputs(1134));
    layer5_outputs(2312) <= not((layer4_outputs(3986)) and (layer4_outputs(1091)));
    layer5_outputs(2313) <= layer4_outputs(4632);
    layer5_outputs(2314) <= not(layer4_outputs(1508));
    layer5_outputs(2315) <= not(layer4_outputs(4027)) or (layer4_outputs(513));
    layer5_outputs(2316) <= not(layer4_outputs(2355));
    layer5_outputs(2317) <= '1';
    layer5_outputs(2318) <= (layer4_outputs(1593)) and not (layer4_outputs(4289));
    layer5_outputs(2319) <= layer4_outputs(1845);
    layer5_outputs(2320) <= not(layer4_outputs(1284)) or (layer4_outputs(1839));
    layer5_outputs(2321) <= not(layer4_outputs(2195)) or (layer4_outputs(3423));
    layer5_outputs(2322) <= '0';
    layer5_outputs(2323) <= not(layer4_outputs(3159));
    layer5_outputs(2324) <= layer4_outputs(3028);
    layer5_outputs(2325) <= '1';
    layer5_outputs(2326) <= (layer4_outputs(3409)) and (layer4_outputs(3346));
    layer5_outputs(2327) <= not(layer4_outputs(2947)) or (layer4_outputs(1965));
    layer5_outputs(2328) <= not(layer4_outputs(191));
    layer5_outputs(2329) <= not((layer4_outputs(4119)) xor (layer4_outputs(1941)));
    layer5_outputs(2330) <= (layer4_outputs(970)) and (layer4_outputs(3475));
    layer5_outputs(2331) <= not(layer4_outputs(4190)) or (layer4_outputs(839));
    layer5_outputs(2332) <= (layer4_outputs(362)) and not (layer4_outputs(2430));
    layer5_outputs(2333) <= (layer4_outputs(2059)) and (layer4_outputs(421));
    layer5_outputs(2334) <= not((layer4_outputs(3965)) and (layer4_outputs(4979)));
    layer5_outputs(2335) <= (layer4_outputs(1308)) and not (layer4_outputs(4130));
    layer5_outputs(2336) <= not((layer4_outputs(279)) or (layer4_outputs(442)));
    layer5_outputs(2337) <= (layer4_outputs(502)) and (layer4_outputs(2385));
    layer5_outputs(2338) <= layer4_outputs(681);
    layer5_outputs(2339) <= '0';
    layer5_outputs(2340) <= not((layer4_outputs(3865)) or (layer4_outputs(4221)));
    layer5_outputs(2341) <= not(layer4_outputs(2884)) or (layer4_outputs(889));
    layer5_outputs(2342) <= not(layer4_outputs(1111));
    layer5_outputs(2343) <= '0';
    layer5_outputs(2344) <= not(layer4_outputs(2534));
    layer5_outputs(2345) <= layer4_outputs(2191);
    layer5_outputs(2346) <= not((layer4_outputs(2416)) and (layer4_outputs(843)));
    layer5_outputs(2347) <= layer4_outputs(4848);
    layer5_outputs(2348) <= (layer4_outputs(4815)) xor (layer4_outputs(3645));
    layer5_outputs(2349) <= layer4_outputs(1483);
    layer5_outputs(2350) <= (layer4_outputs(198)) and (layer4_outputs(3631));
    layer5_outputs(2351) <= layer4_outputs(523);
    layer5_outputs(2352) <= not(layer4_outputs(1738)) or (layer4_outputs(4059));
    layer5_outputs(2353) <= not(layer4_outputs(2471)) or (layer4_outputs(2075));
    layer5_outputs(2354) <= not(layer4_outputs(3622));
    layer5_outputs(2355) <= not(layer4_outputs(1880)) or (layer4_outputs(892));
    layer5_outputs(2356) <= (layer4_outputs(3434)) and not (layer4_outputs(990));
    layer5_outputs(2357) <= not(layer4_outputs(213));
    layer5_outputs(2358) <= not((layer4_outputs(2319)) and (layer4_outputs(1000)));
    layer5_outputs(2359) <= (layer4_outputs(2425)) and (layer4_outputs(2651));
    layer5_outputs(2360) <= (layer4_outputs(2250)) or (layer4_outputs(2780));
    layer5_outputs(2361) <= '1';
    layer5_outputs(2362) <= not(layer4_outputs(3165)) or (layer4_outputs(2663));
    layer5_outputs(2363) <= not(layer4_outputs(5027));
    layer5_outputs(2364) <= (layer4_outputs(3144)) and not (layer4_outputs(178));
    layer5_outputs(2365) <= not(layer4_outputs(3524));
    layer5_outputs(2366) <= not(layer4_outputs(1828));
    layer5_outputs(2367) <= layer4_outputs(4641);
    layer5_outputs(2368) <= not(layer4_outputs(3976));
    layer5_outputs(2369) <= not((layer4_outputs(3983)) xor (layer4_outputs(2653)));
    layer5_outputs(2370) <= not(layer4_outputs(3832));
    layer5_outputs(2371) <= layer4_outputs(4914);
    layer5_outputs(2372) <= layer4_outputs(2737);
    layer5_outputs(2373) <= (layer4_outputs(1539)) and (layer4_outputs(4369));
    layer5_outputs(2374) <= '0';
    layer5_outputs(2375) <= layer4_outputs(3887);
    layer5_outputs(2376) <= layer4_outputs(2174);
    layer5_outputs(2377) <= not((layer4_outputs(3439)) xor (layer4_outputs(3145)));
    layer5_outputs(2378) <= not(layer4_outputs(393)) or (layer4_outputs(840));
    layer5_outputs(2379) <= (layer4_outputs(3519)) and (layer4_outputs(1698));
    layer5_outputs(2380) <= layer4_outputs(266);
    layer5_outputs(2381) <= (layer4_outputs(3585)) and not (layer4_outputs(1795));
    layer5_outputs(2382) <= not(layer4_outputs(2849)) or (layer4_outputs(807));
    layer5_outputs(2383) <= (layer4_outputs(761)) or (layer4_outputs(4474));
    layer5_outputs(2384) <= not((layer4_outputs(458)) or (layer4_outputs(3872)));
    layer5_outputs(2385) <= '1';
    layer5_outputs(2386) <= not((layer4_outputs(2685)) or (layer4_outputs(4978)));
    layer5_outputs(2387) <= not((layer4_outputs(2666)) and (layer4_outputs(5084)));
    layer5_outputs(2388) <= '0';
    layer5_outputs(2389) <= layer4_outputs(4094);
    layer5_outputs(2390) <= not(layer4_outputs(4085)) or (layer4_outputs(3189));
    layer5_outputs(2391) <= not(layer4_outputs(3455));
    layer5_outputs(2392) <= not(layer4_outputs(1867)) or (layer4_outputs(2560));
    layer5_outputs(2393) <= (layer4_outputs(4507)) and (layer4_outputs(3060));
    layer5_outputs(2394) <= layer4_outputs(1443);
    layer5_outputs(2395) <= not(layer4_outputs(2197));
    layer5_outputs(2396) <= (layer4_outputs(530)) and (layer4_outputs(535));
    layer5_outputs(2397) <= layer4_outputs(3102);
    layer5_outputs(2398) <= layer4_outputs(2726);
    layer5_outputs(2399) <= layer4_outputs(3998);
    layer5_outputs(2400) <= not(layer4_outputs(1379));
    layer5_outputs(2401) <= not(layer4_outputs(2907));
    layer5_outputs(2402) <= not(layer4_outputs(2745));
    layer5_outputs(2403) <= not((layer4_outputs(3298)) or (layer4_outputs(2345)));
    layer5_outputs(2404) <= not(layer4_outputs(4386));
    layer5_outputs(2405) <= layer4_outputs(2509);
    layer5_outputs(2406) <= not((layer4_outputs(3372)) and (layer4_outputs(493)));
    layer5_outputs(2407) <= layer4_outputs(286);
    layer5_outputs(2408) <= (layer4_outputs(1166)) or (layer4_outputs(3631));
    layer5_outputs(2409) <= not(layer4_outputs(5112)) or (layer4_outputs(830));
    layer5_outputs(2410) <= (layer4_outputs(4108)) xor (layer4_outputs(3435));
    layer5_outputs(2411) <= (layer4_outputs(4668)) and not (layer4_outputs(4683));
    layer5_outputs(2412) <= '1';
    layer5_outputs(2413) <= not(layer4_outputs(4586));
    layer5_outputs(2414) <= '1';
    layer5_outputs(2415) <= (layer4_outputs(4289)) or (layer4_outputs(4049));
    layer5_outputs(2416) <= not(layer4_outputs(1749));
    layer5_outputs(2417) <= not((layer4_outputs(2051)) or (layer4_outputs(3291)));
    layer5_outputs(2418) <= not(layer4_outputs(3864));
    layer5_outputs(2419) <= '1';
    layer5_outputs(2420) <= layer4_outputs(3891);
    layer5_outputs(2421) <= not(layer4_outputs(1045));
    layer5_outputs(2422) <= (layer4_outputs(3808)) or (layer4_outputs(1806));
    layer5_outputs(2423) <= '0';
    layer5_outputs(2424) <= not(layer4_outputs(1047)) or (layer4_outputs(2703));
    layer5_outputs(2425) <= layer4_outputs(4293);
    layer5_outputs(2426) <= layer4_outputs(1428);
    layer5_outputs(2427) <= (layer4_outputs(674)) and not (layer4_outputs(3936));
    layer5_outputs(2428) <= '1';
    layer5_outputs(2429) <= layer4_outputs(1639);
    layer5_outputs(2430) <= '0';
    layer5_outputs(2431) <= not((layer4_outputs(1190)) and (layer4_outputs(1943)));
    layer5_outputs(2432) <= (layer4_outputs(1485)) or (layer4_outputs(3469));
    layer5_outputs(2433) <= (layer4_outputs(4797)) and not (layer4_outputs(4013));
    layer5_outputs(2434) <= (layer4_outputs(400)) and (layer4_outputs(1552));
    layer5_outputs(2435) <= not(layer4_outputs(1048));
    layer5_outputs(2436) <= not(layer4_outputs(2204));
    layer5_outputs(2437) <= layer4_outputs(2135);
    layer5_outputs(2438) <= layer4_outputs(3176);
    layer5_outputs(2439) <= (layer4_outputs(4378)) xor (layer4_outputs(1500));
    layer5_outputs(2440) <= not(layer4_outputs(3879));
    layer5_outputs(2441) <= not((layer4_outputs(3562)) and (layer4_outputs(3917)));
    layer5_outputs(2442) <= not(layer4_outputs(1016));
    layer5_outputs(2443) <= (layer4_outputs(3057)) and (layer4_outputs(2266));
    layer5_outputs(2444) <= (layer4_outputs(3021)) or (layer4_outputs(1684));
    layer5_outputs(2445) <= (layer4_outputs(572)) xor (layer4_outputs(3440));
    layer5_outputs(2446) <= (layer4_outputs(2594)) and not (layer4_outputs(3035));
    layer5_outputs(2447) <= (layer4_outputs(3044)) or (layer4_outputs(2937));
    layer5_outputs(2448) <= '1';
    layer5_outputs(2449) <= not(layer4_outputs(1436));
    layer5_outputs(2450) <= (layer4_outputs(124)) and not (layer4_outputs(2278));
    layer5_outputs(2451) <= '0';
    layer5_outputs(2452) <= (layer4_outputs(383)) or (layer4_outputs(3600));
    layer5_outputs(2453) <= layer4_outputs(1507);
    layer5_outputs(2454) <= not(layer4_outputs(4359));
    layer5_outputs(2455) <= (layer4_outputs(2628)) or (layer4_outputs(168));
    layer5_outputs(2456) <= not((layer4_outputs(4555)) and (layer4_outputs(1267)));
    layer5_outputs(2457) <= not((layer4_outputs(810)) and (layer4_outputs(3708)));
    layer5_outputs(2458) <= (layer4_outputs(781)) and not (layer4_outputs(4644));
    layer5_outputs(2459) <= layer4_outputs(4055);
    layer5_outputs(2460) <= (layer4_outputs(2034)) and (layer4_outputs(2784));
    layer5_outputs(2461) <= layer4_outputs(271);
    layer5_outputs(2462) <= layer4_outputs(3473);
    layer5_outputs(2463) <= not((layer4_outputs(1304)) or (layer4_outputs(3951)));
    layer5_outputs(2464) <= not((layer4_outputs(4171)) or (layer4_outputs(5013)));
    layer5_outputs(2465) <= layer4_outputs(772);
    layer5_outputs(2466) <= not((layer4_outputs(3825)) xor (layer4_outputs(5091)));
    layer5_outputs(2467) <= not(layer4_outputs(1484));
    layer5_outputs(2468) <= not(layer4_outputs(496));
    layer5_outputs(2469) <= (layer4_outputs(4764)) and not (layer4_outputs(1234));
    layer5_outputs(2470) <= not(layer4_outputs(2124));
    layer5_outputs(2471) <= '0';
    layer5_outputs(2472) <= not(layer4_outputs(2175));
    layer5_outputs(2473) <= (layer4_outputs(2178)) and not (layer4_outputs(1283));
    layer5_outputs(2474) <= (layer4_outputs(1876)) and not (layer4_outputs(1229));
    layer5_outputs(2475) <= '1';
    layer5_outputs(2476) <= layer4_outputs(819);
    layer5_outputs(2477) <= (layer4_outputs(4379)) and not (layer4_outputs(3127));
    layer5_outputs(2478) <= not(layer4_outputs(3470)) or (layer4_outputs(998));
    layer5_outputs(2479) <= (layer4_outputs(2501)) or (layer4_outputs(4777));
    layer5_outputs(2480) <= not(layer4_outputs(4948));
    layer5_outputs(2481) <= '0';
    layer5_outputs(2482) <= not((layer4_outputs(3168)) or (layer4_outputs(4276)));
    layer5_outputs(2483) <= '0';
    layer5_outputs(2484) <= not(layer4_outputs(691));
    layer5_outputs(2485) <= not((layer4_outputs(3268)) or (layer4_outputs(3085)));
    layer5_outputs(2486) <= '0';
    layer5_outputs(2487) <= (layer4_outputs(4474)) and (layer4_outputs(4719));
    layer5_outputs(2488) <= not(layer4_outputs(3245));
    layer5_outputs(2489) <= not((layer4_outputs(3204)) and (layer4_outputs(4139)));
    layer5_outputs(2490) <= not(layer4_outputs(3321));
    layer5_outputs(2491) <= layer4_outputs(2685);
    layer5_outputs(2492) <= not(layer4_outputs(2779));
    layer5_outputs(2493) <= (layer4_outputs(4611)) and not (layer4_outputs(3447));
    layer5_outputs(2494) <= layer4_outputs(20);
    layer5_outputs(2495) <= not(layer4_outputs(4917)) or (layer4_outputs(1086));
    layer5_outputs(2496) <= '0';
    layer5_outputs(2497) <= (layer4_outputs(2678)) and not (layer4_outputs(979));
    layer5_outputs(2498) <= (layer4_outputs(2788)) and not (layer4_outputs(3719));
    layer5_outputs(2499) <= not(layer4_outputs(1274)) or (layer4_outputs(1435));
    layer5_outputs(2500) <= not((layer4_outputs(293)) and (layer4_outputs(4473)));
    layer5_outputs(2501) <= '0';
    layer5_outputs(2502) <= (layer4_outputs(4232)) xor (layer4_outputs(1158));
    layer5_outputs(2503) <= '1';
    layer5_outputs(2504) <= not(layer4_outputs(2366));
    layer5_outputs(2505) <= not((layer4_outputs(4463)) or (layer4_outputs(3511)));
    layer5_outputs(2506) <= (layer4_outputs(404)) and not (layer4_outputs(3252));
    layer5_outputs(2507) <= (layer4_outputs(667)) and (layer4_outputs(3859));
    layer5_outputs(2508) <= layer4_outputs(4821);
    layer5_outputs(2509) <= (layer4_outputs(472)) and not (layer4_outputs(1095));
    layer5_outputs(2510) <= layer4_outputs(4689);
    layer5_outputs(2511) <= (layer4_outputs(4292)) and not (layer4_outputs(897));
    layer5_outputs(2512) <= not(layer4_outputs(4234)) or (layer4_outputs(4353));
    layer5_outputs(2513) <= not(layer4_outputs(1580));
    layer5_outputs(2514) <= (layer4_outputs(1372)) or (layer4_outputs(946));
    layer5_outputs(2515) <= (layer4_outputs(264)) and not (layer4_outputs(4324));
    layer5_outputs(2516) <= not(layer4_outputs(1319));
    layer5_outputs(2517) <= (layer4_outputs(1431)) or (layer4_outputs(1728));
    layer5_outputs(2518) <= not((layer4_outputs(5095)) and (layer4_outputs(3988)));
    layer5_outputs(2519) <= (layer4_outputs(4576)) or (layer4_outputs(4881));
    layer5_outputs(2520) <= not(layer4_outputs(938)) or (layer4_outputs(3714));
    layer5_outputs(2521) <= (layer4_outputs(1595)) and not (layer4_outputs(488));
    layer5_outputs(2522) <= (layer4_outputs(878)) xor (layer4_outputs(2237));
    layer5_outputs(2523) <= not(layer4_outputs(979));
    layer5_outputs(2524) <= layer4_outputs(1244);
    layer5_outputs(2525) <= '1';
    layer5_outputs(2526) <= layer4_outputs(2559);
    layer5_outputs(2527) <= layer4_outputs(2741);
    layer5_outputs(2528) <= layer4_outputs(1687);
    layer5_outputs(2529) <= not((layer4_outputs(1706)) or (layer4_outputs(3676)));
    layer5_outputs(2530) <= (layer4_outputs(2202)) or (layer4_outputs(4983));
    layer5_outputs(2531) <= not((layer4_outputs(3048)) and (layer4_outputs(543)));
    layer5_outputs(2532) <= layer4_outputs(1406);
    layer5_outputs(2533) <= not(layer4_outputs(4233)) or (layer4_outputs(3426));
    layer5_outputs(2534) <= not(layer4_outputs(780)) or (layer4_outputs(2928));
    layer5_outputs(2535) <= not((layer4_outputs(4969)) and (layer4_outputs(2688)));
    layer5_outputs(2536) <= not(layer4_outputs(2175));
    layer5_outputs(2537) <= not(layer4_outputs(1557)) or (layer4_outputs(3282));
    layer5_outputs(2538) <= not(layer4_outputs(3271));
    layer5_outputs(2539) <= not((layer4_outputs(1109)) and (layer4_outputs(3798)));
    layer5_outputs(2540) <= not(layer4_outputs(2855));
    layer5_outputs(2541) <= '0';
    layer5_outputs(2542) <= (layer4_outputs(3517)) and (layer4_outputs(2016));
    layer5_outputs(2543) <= layer4_outputs(3945);
    layer5_outputs(2544) <= (layer4_outputs(1706)) xor (layer4_outputs(4917));
    layer5_outputs(2545) <= not((layer4_outputs(4152)) or (layer4_outputs(845)));
    layer5_outputs(2546) <= not(layer4_outputs(476));
    layer5_outputs(2547) <= not(layer4_outputs(459)) or (layer4_outputs(2418));
    layer5_outputs(2548) <= layer4_outputs(1018);
    layer5_outputs(2549) <= not(layer4_outputs(1782)) or (layer4_outputs(4009));
    layer5_outputs(2550) <= (layer4_outputs(4817)) and not (layer4_outputs(4011));
    layer5_outputs(2551) <= not((layer4_outputs(186)) and (layer4_outputs(4972)));
    layer5_outputs(2552) <= not((layer4_outputs(2048)) or (layer4_outputs(4425)));
    layer5_outputs(2553) <= not(layer4_outputs(3605));
    layer5_outputs(2554) <= not(layer4_outputs(3025));
    layer5_outputs(2555) <= not((layer4_outputs(1772)) or (layer4_outputs(525)));
    layer5_outputs(2556) <= not(layer4_outputs(1327)) or (layer4_outputs(1891));
    layer5_outputs(2557) <= not((layer4_outputs(1505)) and (layer4_outputs(2932)));
    layer5_outputs(2558) <= not((layer4_outputs(3425)) or (layer4_outputs(588)));
    layer5_outputs(2559) <= not(layer4_outputs(4947)) or (layer4_outputs(1954));
    layer5_outputs(2560) <= not(layer4_outputs(2550));
    layer5_outputs(2561) <= not(layer4_outputs(2682));
    layer5_outputs(2562) <= not(layer4_outputs(3073)) or (layer4_outputs(2694));
    layer5_outputs(2563) <= not(layer4_outputs(1932));
    layer5_outputs(2564) <= not(layer4_outputs(4007)) or (layer4_outputs(1023));
    layer5_outputs(2565) <= not((layer4_outputs(3748)) and (layer4_outputs(2293)));
    layer5_outputs(2566) <= (layer4_outputs(52)) and (layer4_outputs(1203));
    layer5_outputs(2567) <= not((layer4_outputs(443)) and (layer4_outputs(3485)));
    layer5_outputs(2568) <= (layer4_outputs(1240)) and not (layer4_outputs(2572));
    layer5_outputs(2569) <= layer4_outputs(2613);
    layer5_outputs(2570) <= not((layer4_outputs(3114)) and (layer4_outputs(4041)));
    layer5_outputs(2571) <= not((layer4_outputs(2889)) xor (layer4_outputs(676)));
    layer5_outputs(2572) <= (layer4_outputs(4921)) or (layer4_outputs(351));
    layer5_outputs(2573) <= layer4_outputs(3);
    layer5_outputs(2574) <= (layer4_outputs(3710)) and (layer4_outputs(58));
    layer5_outputs(2575) <= (layer4_outputs(3987)) and not (layer4_outputs(2082));
    layer5_outputs(2576) <= not((layer4_outputs(4783)) and (layer4_outputs(4734)));
    layer5_outputs(2577) <= not((layer4_outputs(5118)) or (layer4_outputs(2836)));
    layer5_outputs(2578) <= layer4_outputs(4129);
    layer5_outputs(2579) <= (layer4_outputs(1632)) or (layer4_outputs(1830));
    layer5_outputs(2580) <= layer4_outputs(1603);
    layer5_outputs(2581) <= not(layer4_outputs(4334));
    layer5_outputs(2582) <= not(layer4_outputs(589)) or (layer4_outputs(3849));
    layer5_outputs(2583) <= not(layer4_outputs(3706)) or (layer4_outputs(3527));
    layer5_outputs(2584) <= not((layer4_outputs(262)) or (layer4_outputs(3154)));
    layer5_outputs(2585) <= not(layer4_outputs(4536));
    layer5_outputs(2586) <= not(layer4_outputs(1241)) or (layer4_outputs(4603));
    layer5_outputs(2587) <= '1';
    layer5_outputs(2588) <= '1';
    layer5_outputs(2589) <= not(layer4_outputs(1791)) or (layer4_outputs(4302));
    layer5_outputs(2590) <= (layer4_outputs(1380)) and (layer4_outputs(641));
    layer5_outputs(2591) <= not(layer4_outputs(4606)) or (layer4_outputs(3259));
    layer5_outputs(2592) <= not(layer4_outputs(42)) or (layer4_outputs(2860));
    layer5_outputs(2593) <= (layer4_outputs(1532)) and (layer4_outputs(2200));
    layer5_outputs(2594) <= not(layer4_outputs(4065));
    layer5_outputs(2595) <= not(layer4_outputs(3497)) or (layer4_outputs(4593));
    layer5_outputs(2596) <= not(layer4_outputs(1133)) or (layer4_outputs(3986));
    layer5_outputs(2597) <= not(layer4_outputs(5033));
    layer5_outputs(2598) <= layer4_outputs(3603);
    layer5_outputs(2599) <= not(layer4_outputs(1360)) or (layer4_outputs(4610));
    layer5_outputs(2600) <= not(layer4_outputs(352));
    layer5_outputs(2601) <= (layer4_outputs(771)) xor (layer4_outputs(560));
    layer5_outputs(2602) <= (layer4_outputs(1952)) and (layer4_outputs(1175));
    layer5_outputs(2603) <= (layer4_outputs(1005)) and not (layer4_outputs(3209));
    layer5_outputs(2604) <= not(layer4_outputs(1631)) or (layer4_outputs(884));
    layer5_outputs(2605) <= (layer4_outputs(1900)) and not (layer4_outputs(2859));
    layer5_outputs(2606) <= not(layer4_outputs(199)) or (layer4_outputs(1778));
    layer5_outputs(2607) <= '0';
    layer5_outputs(2608) <= not(layer4_outputs(4156)) or (layer4_outputs(4052));
    layer5_outputs(2609) <= not(layer4_outputs(1369));
    layer5_outputs(2610) <= not(layer4_outputs(3598)) or (layer4_outputs(2738));
    layer5_outputs(2611) <= not(layer4_outputs(418)) or (layer4_outputs(2125));
    layer5_outputs(2612) <= not((layer4_outputs(3785)) xor (layer4_outputs(2378)));
    layer5_outputs(2613) <= not(layer4_outputs(604));
    layer5_outputs(2614) <= not(layer4_outputs(2328));
    layer5_outputs(2615) <= layer4_outputs(2610);
    layer5_outputs(2616) <= not((layer4_outputs(4742)) and (layer4_outputs(4328)));
    layer5_outputs(2617) <= (layer4_outputs(2532)) and not (layer4_outputs(2307));
    layer5_outputs(2618) <= layer4_outputs(3237);
    layer5_outputs(2619) <= not(layer4_outputs(4791));
    layer5_outputs(2620) <= layer4_outputs(686);
    layer5_outputs(2621) <= (layer4_outputs(4111)) and not (layer4_outputs(4258));
    layer5_outputs(2622) <= not(layer4_outputs(98));
    layer5_outputs(2623) <= (layer4_outputs(1926)) and not (layer4_outputs(4029));
    layer5_outputs(2624) <= (layer4_outputs(4751)) and not (layer4_outputs(4106));
    layer5_outputs(2625) <= not(layer4_outputs(711));
    layer5_outputs(2626) <= (layer4_outputs(888)) or (layer4_outputs(85));
    layer5_outputs(2627) <= layer4_outputs(2621);
    layer5_outputs(2628) <= not(layer4_outputs(3089));
    layer5_outputs(2629) <= not(layer4_outputs(4187));
    layer5_outputs(2630) <= layer4_outputs(1462);
    layer5_outputs(2631) <= (layer4_outputs(4054)) or (layer4_outputs(2897));
    layer5_outputs(2632) <= layer4_outputs(2352);
    layer5_outputs(2633) <= not(layer4_outputs(2867));
    layer5_outputs(2634) <= not((layer4_outputs(4688)) xor (layer4_outputs(2041)));
    layer5_outputs(2635) <= '1';
    layer5_outputs(2636) <= not(layer4_outputs(2246));
    layer5_outputs(2637) <= not(layer4_outputs(1239)) or (layer4_outputs(2543));
    layer5_outputs(2638) <= '1';
    layer5_outputs(2639) <= layer4_outputs(2992);
    layer5_outputs(2640) <= (layer4_outputs(4771)) and not (layer4_outputs(1775));
    layer5_outputs(2641) <= not(layer4_outputs(3807));
    layer5_outputs(2642) <= (layer4_outputs(3803)) and (layer4_outputs(4652));
    layer5_outputs(2643) <= not(layer4_outputs(4937)) or (layer4_outputs(4631));
    layer5_outputs(2644) <= (layer4_outputs(2792)) and (layer4_outputs(3000));
    layer5_outputs(2645) <= not(layer4_outputs(3799));
    layer5_outputs(2646) <= (layer4_outputs(1566)) and not (layer4_outputs(4266));
    layer5_outputs(2647) <= layer4_outputs(757);
    layer5_outputs(2648) <= layer4_outputs(1066);
    layer5_outputs(2649) <= not((layer4_outputs(4825)) or (layer4_outputs(800)));
    layer5_outputs(2650) <= not(layer4_outputs(2162));
    layer5_outputs(2651) <= not(layer4_outputs(3039));
    layer5_outputs(2652) <= not(layer4_outputs(1417)) or (layer4_outputs(2948));
    layer5_outputs(2653) <= not((layer4_outputs(3683)) and (layer4_outputs(3749)));
    layer5_outputs(2654) <= (layer4_outputs(2652)) and not (layer4_outputs(2935));
    layer5_outputs(2655) <= not((layer4_outputs(1450)) and (layer4_outputs(3115)));
    layer5_outputs(2656) <= not(layer4_outputs(220));
    layer5_outputs(2657) <= layer4_outputs(2606);
    layer5_outputs(2658) <= not((layer4_outputs(4834)) xor (layer4_outputs(2920)));
    layer5_outputs(2659) <= (layer4_outputs(2640)) and (layer4_outputs(2514));
    layer5_outputs(2660) <= not((layer4_outputs(3614)) and (layer4_outputs(4851)));
    layer5_outputs(2661) <= layer4_outputs(4671);
    layer5_outputs(2662) <= '0';
    layer5_outputs(2663) <= layer4_outputs(1908);
    layer5_outputs(2664) <= layer4_outputs(2322);
    layer5_outputs(2665) <= (layer4_outputs(161)) xor (layer4_outputs(1490));
    layer5_outputs(2666) <= layer4_outputs(1910);
    layer5_outputs(2667) <= not(layer4_outputs(3876));
    layer5_outputs(2668) <= not((layer4_outputs(2467)) and (layer4_outputs(3984)));
    layer5_outputs(2669) <= (layer4_outputs(4894)) and not (layer4_outputs(4538));
    layer5_outputs(2670) <= '0';
    layer5_outputs(2671) <= not(layer4_outputs(4944)) or (layer4_outputs(2789));
    layer5_outputs(2672) <= not(layer4_outputs(5029)) or (layer4_outputs(4133));
    layer5_outputs(2673) <= not(layer4_outputs(1193));
    layer5_outputs(2674) <= not(layer4_outputs(1756));
    layer5_outputs(2675) <= not(layer4_outputs(2189)) or (layer4_outputs(1954));
    layer5_outputs(2676) <= '0';
    layer5_outputs(2677) <= layer4_outputs(3381);
    layer5_outputs(2678) <= '0';
    layer5_outputs(2679) <= (layer4_outputs(2930)) and not (layer4_outputs(104));
    layer5_outputs(2680) <= not(layer4_outputs(2688));
    layer5_outputs(2681) <= not(layer4_outputs(3608));
    layer5_outputs(2682) <= '1';
    layer5_outputs(2683) <= not((layer4_outputs(4616)) xor (layer4_outputs(3106)));
    layer5_outputs(2684) <= (layer4_outputs(1141)) and (layer4_outputs(1029));
    layer5_outputs(2685) <= not(layer4_outputs(315));
    layer5_outputs(2686) <= layer4_outputs(4591);
    layer5_outputs(2687) <= (layer4_outputs(611)) xor (layer4_outputs(1512));
    layer5_outputs(2688) <= not((layer4_outputs(1505)) or (layer4_outputs(2456)));
    layer5_outputs(2689) <= (layer4_outputs(743)) and not (layer4_outputs(4296));
    layer5_outputs(2690) <= not(layer4_outputs(4513));
    layer5_outputs(2691) <= not(layer4_outputs(390)) or (layer4_outputs(5010));
    layer5_outputs(2692) <= not(layer4_outputs(2149));
    layer5_outputs(2693) <= (layer4_outputs(3674)) or (layer4_outputs(2423));
    layer5_outputs(2694) <= (layer4_outputs(2918)) and not (layer4_outputs(942));
    layer5_outputs(2695) <= (layer4_outputs(2258)) and not (layer4_outputs(3978));
    layer5_outputs(2696) <= not(layer4_outputs(1934)) or (layer4_outputs(4351));
    layer5_outputs(2697) <= layer4_outputs(152);
    layer5_outputs(2698) <= (layer4_outputs(4228)) and not (layer4_outputs(4912));
    layer5_outputs(2699) <= layer4_outputs(1088);
    layer5_outputs(2700) <= '0';
    layer5_outputs(2701) <= not(layer4_outputs(1444));
    layer5_outputs(2702) <= (layer4_outputs(698)) or (layer4_outputs(4874));
    layer5_outputs(2703) <= (layer4_outputs(4020)) xor (layer4_outputs(3132));
    layer5_outputs(2704) <= '1';
    layer5_outputs(2705) <= layer4_outputs(5083);
    layer5_outputs(2706) <= layer4_outputs(1123);
    layer5_outputs(2707) <= not((layer4_outputs(4462)) and (layer4_outputs(2444)));
    layer5_outputs(2708) <= '0';
    layer5_outputs(2709) <= not(layer4_outputs(584));
    layer5_outputs(2710) <= not(layer4_outputs(3255));
    layer5_outputs(2711) <= not(layer4_outputs(746));
    layer5_outputs(2712) <= layer4_outputs(570);
    layer5_outputs(2713) <= (layer4_outputs(4233)) and not (layer4_outputs(82));
    layer5_outputs(2714) <= layer4_outputs(2172);
    layer5_outputs(2715) <= layer4_outputs(2504);
    layer5_outputs(2716) <= '0';
    layer5_outputs(2717) <= '1';
    layer5_outputs(2718) <= not(layer4_outputs(4158)) or (layer4_outputs(4577));
    layer5_outputs(2719) <= (layer4_outputs(493)) and not (layer4_outputs(1246));
    layer5_outputs(2720) <= not((layer4_outputs(2620)) and (layer4_outputs(4428)));
    layer5_outputs(2721) <= (layer4_outputs(3081)) and not (layer4_outputs(2759));
    layer5_outputs(2722) <= not(layer4_outputs(4297)) or (layer4_outputs(1904));
    layer5_outputs(2723) <= not(layer4_outputs(3840)) or (layer4_outputs(2315));
    layer5_outputs(2724) <= (layer4_outputs(3370)) and not (layer4_outputs(3624));
    layer5_outputs(2725) <= not((layer4_outputs(1495)) and (layer4_outputs(172)));
    layer5_outputs(2726) <= layer4_outputs(2052);
    layer5_outputs(2727) <= not(layer4_outputs(1368)) or (layer4_outputs(1882));
    layer5_outputs(2728) <= (layer4_outputs(599)) xor (layer4_outputs(4740));
    layer5_outputs(2729) <= (layer4_outputs(5089)) and not (layer4_outputs(356));
    layer5_outputs(2730) <= (layer4_outputs(238)) and not (layer4_outputs(4186));
    layer5_outputs(2731) <= '1';
    layer5_outputs(2732) <= not(layer4_outputs(2443));
    layer5_outputs(2733) <= (layer4_outputs(4415)) and not (layer4_outputs(2924));
    layer5_outputs(2734) <= (layer4_outputs(2840)) and not (layer4_outputs(4809));
    layer5_outputs(2735) <= not(layer4_outputs(3076));
    layer5_outputs(2736) <= not(layer4_outputs(1898)) or (layer4_outputs(1793));
    layer5_outputs(2737) <= not(layer4_outputs(2143)) or (layer4_outputs(1465));
    layer5_outputs(2738) <= '0';
    layer5_outputs(2739) <= not(layer4_outputs(647));
    layer5_outputs(2740) <= not(layer4_outputs(10)) or (layer4_outputs(4758));
    layer5_outputs(2741) <= (layer4_outputs(3654)) and (layer4_outputs(706));
    layer5_outputs(2742) <= not(layer4_outputs(3864));
    layer5_outputs(2743) <= not(layer4_outputs(3267)) or (layer4_outputs(4418));
    layer5_outputs(2744) <= layer4_outputs(1013);
    layer5_outputs(2745) <= layer4_outputs(5093);
    layer5_outputs(2746) <= (layer4_outputs(4654)) or (layer4_outputs(3376));
    layer5_outputs(2747) <= not(layer4_outputs(2961));
    layer5_outputs(2748) <= not((layer4_outputs(3240)) and (layer4_outputs(688)));
    layer5_outputs(2749) <= not(layer4_outputs(2445));
    layer5_outputs(2750) <= not((layer4_outputs(2134)) or (layer4_outputs(2493)));
    layer5_outputs(2751) <= not(layer4_outputs(3065));
    layer5_outputs(2752) <= not(layer4_outputs(2303));
    layer5_outputs(2753) <= '1';
    layer5_outputs(2754) <= '1';
    layer5_outputs(2755) <= not((layer4_outputs(4645)) or (layer4_outputs(4862)));
    layer5_outputs(2756) <= (layer4_outputs(104)) or (layer4_outputs(1772));
    layer5_outputs(2757) <= layer4_outputs(835);
    layer5_outputs(2758) <= not(layer4_outputs(1740)) or (layer4_outputs(635));
    layer5_outputs(2759) <= not(layer4_outputs(2709));
    layer5_outputs(2760) <= not(layer4_outputs(1825));
    layer5_outputs(2761) <= layer4_outputs(1055);
    layer5_outputs(2762) <= not(layer4_outputs(377));
    layer5_outputs(2763) <= (layer4_outputs(1670)) and not (layer4_outputs(4040));
    layer5_outputs(2764) <= not(layer4_outputs(3618));
    layer5_outputs(2765) <= not(layer4_outputs(627));
    layer5_outputs(2766) <= layer4_outputs(3794);
    layer5_outputs(2767) <= not(layer4_outputs(4624));
    layer5_outputs(2768) <= layer4_outputs(169);
    layer5_outputs(2769) <= layer4_outputs(17);
    layer5_outputs(2770) <= '1';
    layer5_outputs(2771) <= not(layer4_outputs(3752)) or (layer4_outputs(3825));
    layer5_outputs(2772) <= (layer4_outputs(3341)) and not (layer4_outputs(4612));
    layer5_outputs(2773) <= not(layer4_outputs(1810)) or (layer4_outputs(3052));
    layer5_outputs(2774) <= (layer4_outputs(2125)) and (layer4_outputs(4038));
    layer5_outputs(2775) <= (layer4_outputs(1533)) and not (layer4_outputs(1838));
    layer5_outputs(2776) <= not((layer4_outputs(810)) and (layer4_outputs(1549)));
    layer5_outputs(2777) <= not(layer4_outputs(3617));
    layer5_outputs(2778) <= '0';
    layer5_outputs(2779) <= not((layer4_outputs(1868)) or (layer4_outputs(2865)));
    layer5_outputs(2780) <= (layer4_outputs(2235)) and (layer4_outputs(74));
    layer5_outputs(2781) <= (layer4_outputs(2700)) or (layer4_outputs(1260));
    layer5_outputs(2782) <= (layer4_outputs(3411)) and (layer4_outputs(5055));
    layer5_outputs(2783) <= not(layer4_outputs(4401));
    layer5_outputs(2784) <= not((layer4_outputs(66)) xor (layer4_outputs(5108)));
    layer5_outputs(2785) <= (layer4_outputs(1269)) or (layer4_outputs(4245));
    layer5_outputs(2786) <= not(layer4_outputs(2338));
    layer5_outputs(2787) <= (layer4_outputs(3828)) and not (layer4_outputs(2527));
    layer5_outputs(2788) <= (layer4_outputs(414)) and not (layer4_outputs(1724));
    layer5_outputs(2789) <= layer4_outputs(2218);
    layer5_outputs(2790) <= not(layer4_outputs(2547));
    layer5_outputs(2791) <= (layer4_outputs(4940)) and not (layer4_outputs(852));
    layer5_outputs(2792) <= layer4_outputs(3595);
    layer5_outputs(2793) <= layer4_outputs(2883);
    layer5_outputs(2794) <= (layer4_outputs(945)) and not (layer4_outputs(2451));
    layer5_outputs(2795) <= '1';
    layer5_outputs(2796) <= '0';
    layer5_outputs(2797) <= not(layer4_outputs(1649));
    layer5_outputs(2798) <= not((layer4_outputs(1409)) and (layer4_outputs(3636)));
    layer5_outputs(2799) <= not(layer4_outputs(4540));
    layer5_outputs(2800) <= (layer4_outputs(3061)) and not (layer4_outputs(4268));
    layer5_outputs(2801) <= layer4_outputs(4992);
    layer5_outputs(2802) <= not(layer4_outputs(1191)) or (layer4_outputs(4844));
    layer5_outputs(2803) <= not(layer4_outputs(1180));
    layer5_outputs(2804) <= '0';
    layer5_outputs(2805) <= not((layer4_outputs(3810)) or (layer4_outputs(4247)));
    layer5_outputs(2806) <= (layer4_outputs(5053)) or (layer4_outputs(2037));
    layer5_outputs(2807) <= layer4_outputs(2274);
    layer5_outputs(2808) <= (layer4_outputs(4714)) and (layer4_outputs(4201));
    layer5_outputs(2809) <= '0';
    layer5_outputs(2810) <= not(layer4_outputs(4952));
    layer5_outputs(2811) <= not((layer4_outputs(3177)) xor (layer4_outputs(1427)));
    layer5_outputs(2812) <= not((layer4_outputs(2558)) or (layer4_outputs(4903)));
    layer5_outputs(2813) <= not(layer4_outputs(4777)) or (layer4_outputs(1892));
    layer5_outputs(2814) <= not(layer4_outputs(942));
    layer5_outputs(2815) <= not(layer4_outputs(535));
    layer5_outputs(2816) <= not(layer4_outputs(3051));
    layer5_outputs(2817) <= (layer4_outputs(4532)) or (layer4_outputs(1101));
    layer5_outputs(2818) <= layer4_outputs(4882);
    layer5_outputs(2819) <= layer4_outputs(4344);
    layer5_outputs(2820) <= not(layer4_outputs(4018)) or (layer4_outputs(3558));
    layer5_outputs(2821) <= not(layer4_outputs(2477));
    layer5_outputs(2822) <= not(layer4_outputs(4865)) or (layer4_outputs(4726));
    layer5_outputs(2823) <= layer4_outputs(1540);
    layer5_outputs(2824) <= not((layer4_outputs(4793)) and (layer4_outputs(2824)));
    layer5_outputs(2825) <= layer4_outputs(171);
    layer5_outputs(2826) <= (layer4_outputs(2133)) and not (layer4_outputs(1584));
    layer5_outputs(2827) <= not(layer4_outputs(300)) or (layer4_outputs(4750));
    layer5_outputs(2828) <= not((layer4_outputs(3972)) xor (layer4_outputs(100)));
    layer5_outputs(2829) <= not((layer4_outputs(2364)) and (layer4_outputs(1809)));
    layer5_outputs(2830) <= '0';
    layer5_outputs(2831) <= (layer4_outputs(2774)) and (layer4_outputs(4202));
    layer5_outputs(2832) <= not(layer4_outputs(2583)) or (layer4_outputs(4356));
    layer5_outputs(2833) <= not((layer4_outputs(204)) or (layer4_outputs(1407)));
    layer5_outputs(2834) <= '1';
    layer5_outputs(2835) <= (layer4_outputs(4856)) and (layer4_outputs(3114));
    layer5_outputs(2836) <= '0';
    layer5_outputs(2837) <= '1';
    layer5_outputs(2838) <= layer4_outputs(1836);
    layer5_outputs(2839) <= not(layer4_outputs(2625)) or (layer4_outputs(4465));
    layer5_outputs(2840) <= not(layer4_outputs(3236));
    layer5_outputs(2841) <= not(layer4_outputs(2993)) or (layer4_outputs(3140));
    layer5_outputs(2842) <= not(layer4_outputs(3432)) or (layer4_outputs(2276));
    layer5_outputs(2843) <= not(layer4_outputs(17));
    layer5_outputs(2844) <= not(layer4_outputs(1351)) or (layer4_outputs(4607));
    layer5_outputs(2845) <= (layer4_outputs(3786)) and not (layer4_outputs(4090));
    layer5_outputs(2846) <= layer4_outputs(1414);
    layer5_outputs(2847) <= layer4_outputs(2996);
    layer5_outputs(2848) <= not(layer4_outputs(3717));
    layer5_outputs(2849) <= layer4_outputs(3447);
    layer5_outputs(2850) <= not(layer4_outputs(3766));
    layer5_outputs(2851) <= not((layer4_outputs(2071)) or (layer4_outputs(2264)));
    layer5_outputs(2852) <= not(layer4_outputs(5097));
    layer5_outputs(2853) <= (layer4_outputs(1887)) or (layer4_outputs(3989));
    layer5_outputs(2854) <= '1';
    layer5_outputs(2855) <= not((layer4_outputs(3154)) or (layer4_outputs(2550)));
    layer5_outputs(2856) <= '0';
    layer5_outputs(2857) <= '0';
    layer5_outputs(2858) <= '0';
    layer5_outputs(2859) <= layer4_outputs(2311);
    layer5_outputs(2860) <= not((layer4_outputs(1080)) xor (layer4_outputs(1347)));
    layer5_outputs(2861) <= (layer4_outputs(3933)) and (layer4_outputs(1289));
    layer5_outputs(2862) <= not(layer4_outputs(4513));
    layer5_outputs(2863) <= (layer4_outputs(4364)) and (layer4_outputs(1674));
    layer5_outputs(2864) <= (layer4_outputs(2796)) and not (layer4_outputs(841));
    layer5_outputs(2865) <= (layer4_outputs(1587)) and not (layer4_outputs(2560));
    layer5_outputs(2866) <= (layer4_outputs(4895)) or (layer4_outputs(3889));
    layer5_outputs(2867) <= (layer4_outputs(296)) and (layer4_outputs(4371));
    layer5_outputs(2868) <= not((layer4_outputs(1712)) or (layer4_outputs(4022)));
    layer5_outputs(2869) <= not(layer4_outputs(1342)) or (layer4_outputs(3037));
    layer5_outputs(2870) <= not(layer4_outputs(4873));
    layer5_outputs(2871) <= not((layer4_outputs(4338)) xor (layer4_outputs(1591)));
    layer5_outputs(2872) <= not(layer4_outputs(243));
    layer5_outputs(2873) <= '0';
    layer5_outputs(2874) <= not(layer4_outputs(3869));
    layer5_outputs(2875) <= layer4_outputs(2657);
    layer5_outputs(2876) <= not((layer4_outputs(2524)) and (layer4_outputs(1420)));
    layer5_outputs(2877) <= '0';
    layer5_outputs(2878) <= not(layer4_outputs(2339)) or (layer4_outputs(2145));
    layer5_outputs(2879) <= (layer4_outputs(1368)) or (layer4_outputs(2119));
    layer5_outputs(2880) <= not(layer4_outputs(533));
    layer5_outputs(2881) <= not(layer4_outputs(1953));
    layer5_outputs(2882) <= not(layer4_outputs(2577));
    layer5_outputs(2883) <= layer4_outputs(4294);
    layer5_outputs(2884) <= layer4_outputs(3550);
    layer5_outputs(2885) <= not(layer4_outputs(1398));
    layer5_outputs(2886) <= (layer4_outputs(50)) xor (layer4_outputs(2388));
    layer5_outputs(2887) <= (layer4_outputs(1373)) xor (layer4_outputs(3613));
    layer5_outputs(2888) <= (layer4_outputs(751)) and (layer4_outputs(3188));
    layer5_outputs(2889) <= (layer4_outputs(3251)) or (layer4_outputs(1449));
    layer5_outputs(2890) <= layer4_outputs(603);
    layer5_outputs(2891) <= not((layer4_outputs(2752)) xor (layer4_outputs(1201)));
    layer5_outputs(2892) <= (layer4_outputs(2282)) and not (layer4_outputs(705));
    layer5_outputs(2893) <= not((layer4_outputs(995)) or (layer4_outputs(5050)));
    layer5_outputs(2894) <= layer4_outputs(2457);
    layer5_outputs(2895) <= '0';
    layer5_outputs(2896) <= '1';
    layer5_outputs(2897) <= not(layer4_outputs(4539)) or (layer4_outputs(1308));
    layer5_outputs(2898) <= '0';
    layer5_outputs(2899) <= layer4_outputs(2749);
    layer5_outputs(2900) <= not((layer4_outputs(2873)) and (layer4_outputs(314)));
    layer5_outputs(2901) <= not((layer4_outputs(1989)) and (layer4_outputs(3332)));
    layer5_outputs(2902) <= not(layer4_outputs(3622));
    layer5_outputs(2903) <= layer4_outputs(4960);
    layer5_outputs(2904) <= not((layer4_outputs(3454)) or (layer4_outputs(3722)));
    layer5_outputs(2905) <= layer4_outputs(4542);
    layer5_outputs(2906) <= layer4_outputs(2478);
    layer5_outputs(2907) <= layer4_outputs(3087);
    layer5_outputs(2908) <= not((layer4_outputs(1017)) and (layer4_outputs(602)));
    layer5_outputs(2909) <= layer4_outputs(485);
    layer5_outputs(2910) <= (layer4_outputs(435)) and not (layer4_outputs(1040));
    layer5_outputs(2911) <= not(layer4_outputs(2521));
    layer5_outputs(2912) <= (layer4_outputs(4897)) and not (layer4_outputs(338));
    layer5_outputs(2913) <= '0';
    layer5_outputs(2914) <= layer4_outputs(3417);
    layer5_outputs(2915) <= not(layer4_outputs(2916));
    layer5_outputs(2916) <= (layer4_outputs(3606)) and (layer4_outputs(4305));
    layer5_outputs(2917) <= (layer4_outputs(2196)) xor (layer4_outputs(4742));
    layer5_outputs(2918) <= (layer4_outputs(189)) and not (layer4_outputs(3662));
    layer5_outputs(2919) <= not(layer4_outputs(2063)) or (layer4_outputs(1581));
    layer5_outputs(2920) <= not((layer4_outputs(1589)) and (layer4_outputs(2757)));
    layer5_outputs(2921) <= layer4_outputs(159);
    layer5_outputs(2922) <= not(layer4_outputs(291));
    layer5_outputs(2923) <= not(layer4_outputs(4945));
    layer5_outputs(2924) <= not(layer4_outputs(3164));
    layer5_outputs(2925) <= (layer4_outputs(4971)) and not (layer4_outputs(2909));
    layer5_outputs(2926) <= not(layer4_outputs(1551)) or (layer4_outputs(4252));
    layer5_outputs(2927) <= not(layer4_outputs(1250));
    layer5_outputs(2928) <= not((layer4_outputs(1461)) and (layer4_outputs(3385)));
    layer5_outputs(2929) <= not((layer4_outputs(4821)) or (layer4_outputs(3770)));
    layer5_outputs(2930) <= not(layer4_outputs(4354));
    layer5_outputs(2931) <= not((layer4_outputs(1592)) and (layer4_outputs(2034)));
    layer5_outputs(2932) <= '1';
    layer5_outputs(2933) <= (layer4_outputs(2432)) and not (layer4_outputs(4068));
    layer5_outputs(2934) <= not(layer4_outputs(1474));
    layer5_outputs(2935) <= (layer4_outputs(4813)) and (layer4_outputs(5105));
    layer5_outputs(2936) <= not((layer4_outputs(464)) and (layer4_outputs(3023)));
    layer5_outputs(2937) <= not(layer4_outputs(1743));
    layer5_outputs(2938) <= not((layer4_outputs(3954)) xor (layer4_outputs(1395)));
    layer5_outputs(2939) <= layer4_outputs(1985);
    layer5_outputs(2940) <= not(layer4_outputs(2177)) or (layer4_outputs(4955));
    layer5_outputs(2941) <= not(layer4_outputs(4124));
    layer5_outputs(2942) <= not((layer4_outputs(1254)) xor (layer4_outputs(444)));
    layer5_outputs(2943) <= not(layer4_outputs(4192)) or (layer4_outputs(1129));
    layer5_outputs(2944) <= not(layer4_outputs(1535));
    layer5_outputs(2945) <= not(layer4_outputs(3996));
    layer5_outputs(2946) <= layer4_outputs(4242);
    layer5_outputs(2947) <= not(layer4_outputs(4088));
    layer5_outputs(2948) <= not((layer4_outputs(605)) or (layer4_outputs(750)));
    layer5_outputs(2949) <= not(layer4_outputs(5015)) or (layer4_outputs(1852));
    layer5_outputs(2950) <= (layer4_outputs(1334)) or (layer4_outputs(1858));
    layer5_outputs(2951) <= layer4_outputs(5041);
    layer5_outputs(2952) <= not(layer4_outputs(2857));
    layer5_outputs(2953) <= not(layer4_outputs(4790));
    layer5_outputs(2954) <= layer4_outputs(5111);
    layer5_outputs(2955) <= (layer4_outputs(4381)) xor (layer4_outputs(2708));
    layer5_outputs(2956) <= '1';
    layer5_outputs(2957) <= not((layer4_outputs(3276)) xor (layer4_outputs(3224)));
    layer5_outputs(2958) <= not(layer4_outputs(3507));
    layer5_outputs(2959) <= (layer4_outputs(1719)) and (layer4_outputs(3764));
    layer5_outputs(2960) <= not(layer4_outputs(3350)) or (layer4_outputs(3344));
    layer5_outputs(2961) <= not((layer4_outputs(4301)) or (layer4_outputs(4749)));
    layer5_outputs(2962) <= not(layer4_outputs(2897));
    layer5_outputs(2963) <= (layer4_outputs(2824)) or (layer4_outputs(3143));
    layer5_outputs(2964) <= not(layer4_outputs(567));
    layer5_outputs(2965) <= not(layer4_outputs(3738)) or (layer4_outputs(4995));
    layer5_outputs(2966) <= '0';
    layer5_outputs(2967) <= not((layer4_outputs(4517)) xor (layer4_outputs(3805)));
    layer5_outputs(2968) <= (layer4_outputs(302)) and not (layer4_outputs(1644));
    layer5_outputs(2969) <= not(layer4_outputs(450));
    layer5_outputs(2970) <= not(layer4_outputs(3846));
    layer5_outputs(2971) <= not(layer4_outputs(4653)) or (layer4_outputs(5030));
    layer5_outputs(2972) <= (layer4_outputs(3103)) and not (layer4_outputs(669));
    layer5_outputs(2973) <= not((layer4_outputs(2714)) and (layer4_outputs(3660)));
    layer5_outputs(2974) <= not((layer4_outputs(1294)) and (layer4_outputs(684)));
    layer5_outputs(2975) <= layer4_outputs(4554);
    layer5_outputs(2976) <= not(layer4_outputs(2669));
    layer5_outputs(2977) <= (layer4_outputs(1413)) and not (layer4_outputs(2379));
    layer5_outputs(2978) <= (layer4_outputs(3949)) and not (layer4_outputs(306));
    layer5_outputs(2979) <= not((layer4_outputs(1400)) or (layer4_outputs(2111)));
    layer5_outputs(2980) <= not(layer4_outputs(1898)) or (layer4_outputs(2278));
    layer5_outputs(2981) <= (layer4_outputs(3853)) and (layer4_outputs(2941));
    layer5_outputs(2982) <= layer4_outputs(2008);
    layer5_outputs(2983) <= '0';
    layer5_outputs(2984) <= layer4_outputs(4435);
    layer5_outputs(2985) <= (layer4_outputs(3031)) and not (layer4_outputs(304));
    layer5_outputs(2986) <= (layer4_outputs(1128)) xor (layer4_outputs(4383));
    layer5_outputs(2987) <= layer4_outputs(4592);
    layer5_outputs(2988) <= (layer4_outputs(1002)) or (layer4_outputs(3171));
    layer5_outputs(2989) <= not(layer4_outputs(395));
    layer5_outputs(2990) <= not((layer4_outputs(4806)) or (layer4_outputs(1529)));
    layer5_outputs(2991) <= layer4_outputs(4350);
    layer5_outputs(2992) <= not(layer4_outputs(4973)) or (layer4_outputs(2995));
    layer5_outputs(2993) <= layer4_outputs(4058);
    layer5_outputs(2994) <= not(layer4_outputs(1458)) or (layer4_outputs(4081));
    layer5_outputs(2995) <= not(layer4_outputs(825));
    layer5_outputs(2996) <= (layer4_outputs(4743)) and not (layer4_outputs(94));
    layer5_outputs(2997) <= (layer4_outputs(2838)) or (layer4_outputs(4291));
    layer5_outputs(2998) <= (layer4_outputs(3918)) and not (layer4_outputs(4026));
    layer5_outputs(2999) <= (layer4_outputs(4078)) and not (layer4_outputs(2711));
    layer5_outputs(3000) <= '1';
    layer5_outputs(3001) <= (layer4_outputs(1610)) and (layer4_outputs(4605));
    layer5_outputs(3002) <= not(layer4_outputs(1679));
    layer5_outputs(3003) <= layer4_outputs(2780);
    layer5_outputs(3004) <= not((layer4_outputs(3617)) or (layer4_outputs(1349)));
    layer5_outputs(3005) <= not((layer4_outputs(1594)) and (layer4_outputs(2903)));
    layer5_outputs(3006) <= not((layer4_outputs(4373)) and (layer4_outputs(3548)));
    layer5_outputs(3007) <= (layer4_outputs(1182)) and not (layer4_outputs(2150));
    layer5_outputs(3008) <= (layer4_outputs(671)) and (layer4_outputs(659));
    layer5_outputs(3009) <= not(layer4_outputs(4707)) or (layer4_outputs(2257));
    layer5_outputs(3010) <= layer4_outputs(4801);
    layer5_outputs(3011) <= not((layer4_outputs(3516)) or (layer4_outputs(3158)));
    layer5_outputs(3012) <= layer4_outputs(2346);
    layer5_outputs(3013) <= layer4_outputs(2412);
    layer5_outputs(3014) <= not((layer4_outputs(1710)) xor (layer4_outputs(4615)));
    layer5_outputs(3015) <= not(layer4_outputs(2683));
    layer5_outputs(3016) <= not(layer4_outputs(28));
    layer5_outputs(3017) <= '1';
    layer5_outputs(3018) <= '1';
    layer5_outputs(3019) <= layer4_outputs(1833);
    layer5_outputs(3020) <= not(layer4_outputs(2083));
    layer5_outputs(3021) <= (layer4_outputs(3509)) or (layer4_outputs(1265));
    layer5_outputs(3022) <= not(layer4_outputs(1857)) or (layer4_outputs(4057));
    layer5_outputs(3023) <= not(layer4_outputs(4301)) or (layer4_outputs(3883));
    layer5_outputs(3024) <= layer4_outputs(631);
    layer5_outputs(3025) <= not(layer4_outputs(495)) or (layer4_outputs(2290));
    layer5_outputs(3026) <= not(layer4_outputs(2380));
    layer5_outputs(3027) <= (layer4_outputs(1928)) and not (layer4_outputs(826));
    layer5_outputs(3028) <= layer4_outputs(1764);
    layer5_outputs(3029) <= layer4_outputs(491);
    layer5_outputs(3030) <= not(layer4_outputs(4227));
    layer5_outputs(3031) <= not(layer4_outputs(1280)) or (layer4_outputs(964));
    layer5_outputs(3032) <= (layer4_outputs(1126)) and not (layer4_outputs(2287));
    layer5_outputs(3033) <= not((layer4_outputs(2237)) or (layer4_outputs(3783)));
    layer5_outputs(3034) <= not(layer4_outputs(4323)) or (layer4_outputs(2204));
    layer5_outputs(3035) <= '1';
    layer5_outputs(3036) <= (layer4_outputs(3306)) and (layer4_outputs(1934));
    layer5_outputs(3037) <= not((layer4_outputs(4593)) or (layer4_outputs(4276)));
    layer5_outputs(3038) <= (layer4_outputs(1668)) and not (layer4_outputs(4802));
    layer5_outputs(3039) <= not((layer4_outputs(2272)) and (layer4_outputs(3590)));
    layer5_outputs(3040) <= (layer4_outputs(569)) xor (layer4_outputs(2917));
    layer5_outputs(3041) <= (layer4_outputs(365)) and not (layer4_outputs(486));
    layer5_outputs(3042) <= layer4_outputs(3419);
    layer5_outputs(3043) <= not(layer4_outputs(2154)) or (layer4_outputs(3913));
    layer5_outputs(3044) <= not(layer4_outputs(3246));
    layer5_outputs(3045) <= layer4_outputs(4649);
    layer5_outputs(3046) <= '1';
    layer5_outputs(3047) <= not(layer4_outputs(195));
    layer5_outputs(3048) <= (layer4_outputs(917)) and not (layer4_outputs(1254));
    layer5_outputs(3049) <= (layer4_outputs(1798)) and (layer4_outputs(473));
    layer5_outputs(3050) <= not((layer4_outputs(707)) and (layer4_outputs(3765)));
    layer5_outputs(3051) <= not(layer4_outputs(4359));
    layer5_outputs(3052) <= layer4_outputs(5000);
    layer5_outputs(3053) <= not((layer4_outputs(390)) or (layer4_outputs(4911)));
    layer5_outputs(3054) <= not(layer4_outputs(4409));
    layer5_outputs(3055) <= not(layer4_outputs(4594)) or (layer4_outputs(2565));
    layer5_outputs(3056) <= (layer4_outputs(5099)) and (layer4_outputs(2359));
    layer5_outputs(3057) <= not((layer4_outputs(4338)) and (layer4_outputs(3392)));
    layer5_outputs(3058) <= (layer4_outputs(1889)) or (layer4_outputs(2531));
    layer5_outputs(3059) <= layer4_outputs(3265);
    layer5_outputs(3060) <= (layer4_outputs(1752)) and (layer4_outputs(2249));
    layer5_outputs(3061) <= not((layer4_outputs(2365)) or (layer4_outputs(4000)));
    layer5_outputs(3062) <= layer4_outputs(71);
    layer5_outputs(3063) <= not((layer4_outputs(4440)) and (layer4_outputs(2951)));
    layer5_outputs(3064) <= (layer4_outputs(1266)) xor (layer4_outputs(4440));
    layer5_outputs(3065) <= layer4_outputs(2242);
    layer5_outputs(3066) <= not(layer4_outputs(268)) or (layer4_outputs(2374));
    layer5_outputs(3067) <= (layer4_outputs(3596)) and not (layer4_outputs(3351));
    layer5_outputs(3068) <= layer4_outputs(156);
    layer5_outputs(3069) <= not(layer4_outputs(4611)) or (layer4_outputs(4835));
    layer5_outputs(3070) <= not(layer4_outputs(294)) or (layer4_outputs(1645));
    layer5_outputs(3071) <= not(layer4_outputs(4308));
    layer5_outputs(3072) <= not(layer4_outputs(2227)) or (layer4_outputs(1837));
    layer5_outputs(3073) <= (layer4_outputs(3707)) or (layer4_outputs(4949));
    layer5_outputs(3074) <= not(layer4_outputs(193)) or (layer4_outputs(2211));
    layer5_outputs(3075) <= (layer4_outputs(4553)) or (layer4_outputs(2677));
    layer5_outputs(3076) <= not(layer4_outputs(1040)) or (layer4_outputs(3769));
    layer5_outputs(3077) <= not(layer4_outputs(2213));
    layer5_outputs(3078) <= not(layer4_outputs(1609));
    layer5_outputs(3079) <= not((layer4_outputs(2622)) xor (layer4_outputs(2568)));
    layer5_outputs(3080) <= not((layer4_outputs(1658)) and (layer4_outputs(2902)));
    layer5_outputs(3081) <= layer4_outputs(906);
    layer5_outputs(3082) <= (layer4_outputs(2744)) and not (layer4_outputs(2697));
    layer5_outputs(3083) <= not(layer4_outputs(3784));
    layer5_outputs(3084) <= layer4_outputs(4097);
    layer5_outputs(3085) <= not(layer4_outputs(5079)) or (layer4_outputs(962));
    layer5_outputs(3086) <= not(layer4_outputs(1));
    layer5_outputs(3087) <= layer4_outputs(2456);
    layer5_outputs(3088) <= layer4_outputs(4035);
    layer5_outputs(3089) <= (layer4_outputs(2218)) or (layer4_outputs(2757));
    layer5_outputs(3090) <= '0';
    layer5_outputs(3091) <= not(layer4_outputs(2952));
    layer5_outputs(3092) <= not(layer4_outputs(4415)) or (layer4_outputs(1029));
    layer5_outputs(3093) <= '0';
    layer5_outputs(3094) <= not(layer4_outputs(4723));
    layer5_outputs(3095) <= not((layer4_outputs(4388)) or (layer4_outputs(4240)));
    layer5_outputs(3096) <= (layer4_outputs(4085)) or (layer4_outputs(4325));
    layer5_outputs(3097) <= not(layer4_outputs(2607));
    layer5_outputs(3098) <= layer4_outputs(4042);
    layer5_outputs(3099) <= not(layer4_outputs(71));
    layer5_outputs(3100) <= not(layer4_outputs(576));
    layer5_outputs(3101) <= not(layer4_outputs(3371));
    layer5_outputs(3102) <= not((layer4_outputs(3789)) or (layer4_outputs(4449)));
    layer5_outputs(3103) <= not((layer4_outputs(2516)) or (layer4_outputs(718)));
    layer5_outputs(3104) <= layer4_outputs(1014);
    layer5_outputs(3105) <= not(layer4_outputs(4249));
    layer5_outputs(3106) <= (layer4_outputs(2223)) or (layer4_outputs(116));
    layer5_outputs(3107) <= layer4_outputs(2030);
    layer5_outputs(3108) <= '1';
    layer5_outputs(3109) <= not((layer4_outputs(2681)) or (layer4_outputs(213)));
    layer5_outputs(3110) <= layer4_outputs(2159);
    layer5_outputs(3111) <= not((layer4_outputs(801)) and (layer4_outputs(1855)));
    layer5_outputs(3112) <= not(layer4_outputs(440));
    layer5_outputs(3113) <= not((layer4_outputs(4679)) or (layer4_outputs(991)));
    layer5_outputs(3114) <= '1';
    layer5_outputs(3115) <= not(layer4_outputs(4457)) or (layer4_outputs(1443));
    layer5_outputs(3116) <= (layer4_outputs(4342)) or (layer4_outputs(4998));
    layer5_outputs(3117) <= (layer4_outputs(4065)) and (layer4_outputs(4144));
    layer5_outputs(3118) <= not(layer4_outputs(2441)) or (layer4_outputs(141));
    layer5_outputs(3119) <= not((layer4_outputs(1691)) or (layer4_outputs(2399)));
    layer5_outputs(3120) <= not(layer4_outputs(8));
    layer5_outputs(3121) <= layer4_outputs(509);
    layer5_outputs(3122) <= (layer4_outputs(4295)) and not (layer4_outputs(1611));
    layer5_outputs(3123) <= not((layer4_outputs(2118)) or (layer4_outputs(2209)));
    layer5_outputs(3124) <= not(layer4_outputs(2781)) or (layer4_outputs(569));
    layer5_outputs(3125) <= not(layer4_outputs(4047)) or (layer4_outputs(3905));
    layer5_outputs(3126) <= not((layer4_outputs(4355)) or (layer4_outputs(1092)));
    layer5_outputs(3127) <= not(layer4_outputs(4827)) or (layer4_outputs(632));
    layer5_outputs(3128) <= (layer4_outputs(3479)) or (layer4_outputs(2361));
    layer5_outputs(3129) <= '1';
    layer5_outputs(3130) <= '0';
    layer5_outputs(3131) <= not(layer4_outputs(1425));
    layer5_outputs(3132) <= (layer4_outputs(515)) xor (layer4_outputs(4697));
    layer5_outputs(3133) <= (layer4_outputs(1080)) xor (layer4_outputs(2521));
    layer5_outputs(3134) <= '0';
    layer5_outputs(3135) <= '1';
    layer5_outputs(3136) <= (layer4_outputs(4960)) and not (layer4_outputs(5005));
    layer5_outputs(3137) <= not((layer4_outputs(1712)) and (layer4_outputs(1689)));
    layer5_outputs(3138) <= not(layer4_outputs(4929)) or (layer4_outputs(770));
    layer5_outputs(3139) <= layer4_outputs(2043);
    layer5_outputs(3140) <= layer4_outputs(2109);
    layer5_outputs(3141) <= not(layer4_outputs(4844)) or (layer4_outputs(1471));
    layer5_outputs(3142) <= '1';
    layer5_outputs(3143) <= '0';
    layer5_outputs(3144) <= layer4_outputs(2777);
    layer5_outputs(3145) <= not(layer4_outputs(1419));
    layer5_outputs(3146) <= layer4_outputs(2398);
    layer5_outputs(3147) <= not(layer4_outputs(1711)) or (layer4_outputs(2317));
    layer5_outputs(3148) <= (layer4_outputs(2697)) and (layer4_outputs(4447));
    layer5_outputs(3149) <= layer4_outputs(4840);
    layer5_outputs(3150) <= '1';
    layer5_outputs(3151) <= not(layer4_outputs(3993));
    layer5_outputs(3152) <= not((layer4_outputs(527)) and (layer4_outputs(1481)));
    layer5_outputs(3153) <= not((layer4_outputs(2344)) or (layer4_outputs(3416)));
    layer5_outputs(3154) <= not((layer4_outputs(3118)) xor (layer4_outputs(3032)));
    layer5_outputs(3155) <= (layer4_outputs(3925)) xor (layer4_outputs(745));
    layer5_outputs(3156) <= '0';
    layer5_outputs(3157) <= (layer4_outputs(628)) or (layer4_outputs(2018));
    layer5_outputs(3158) <= '0';
    layer5_outputs(3159) <= not((layer4_outputs(931)) or (layer4_outputs(4797)));
    layer5_outputs(3160) <= not(layer4_outputs(3820));
    layer5_outputs(3161) <= not(layer4_outputs(1006)) or (layer4_outputs(4524));
    layer5_outputs(3162) <= layer4_outputs(1826);
    layer5_outputs(3163) <= not(layer4_outputs(4690)) or (layer4_outputs(4322));
    layer5_outputs(3164) <= not((layer4_outputs(984)) or (layer4_outputs(1303)));
    layer5_outputs(3165) <= not(layer4_outputs(4108));
    layer5_outputs(3166) <= layer4_outputs(1667);
    layer5_outputs(3167) <= (layer4_outputs(3546)) or (layer4_outputs(4788));
    layer5_outputs(3168) <= not(layer4_outputs(1488)) or (layer4_outputs(3197));
    layer5_outputs(3169) <= not(layer4_outputs(2614)) or (layer4_outputs(3101));
    layer5_outputs(3170) <= not((layer4_outputs(3666)) and (layer4_outputs(3338)));
    layer5_outputs(3171) <= (layer4_outputs(3457)) and not (layer4_outputs(4604));
    layer5_outputs(3172) <= not((layer4_outputs(3904)) or (layer4_outputs(1365)));
    layer5_outputs(3173) <= layer4_outputs(3053);
    layer5_outputs(3174) <= (layer4_outputs(1135)) and not (layer4_outputs(4965));
    layer5_outputs(3175) <= layer4_outputs(2774);
    layer5_outputs(3176) <= '1';
    layer5_outputs(3177) <= (layer4_outputs(1305)) and not (layer4_outputs(959));
    layer5_outputs(3178) <= not(layer4_outputs(2738));
    layer5_outputs(3179) <= not(layer4_outputs(3274));
    layer5_outputs(3180) <= not(layer4_outputs(4349)) or (layer4_outputs(1042));
    layer5_outputs(3181) <= not((layer4_outputs(265)) and (layer4_outputs(4488)));
    layer5_outputs(3182) <= layer4_outputs(2822);
    layer5_outputs(3183) <= not(layer4_outputs(3886));
    layer5_outputs(3184) <= (layer4_outputs(4167)) and (layer4_outputs(4143));
    layer5_outputs(3185) <= '1';
    layer5_outputs(3186) <= not((layer4_outputs(4245)) or (layer4_outputs(3861)));
    layer5_outputs(3187) <= not(layer4_outputs(3230)) or (layer4_outputs(610));
    layer5_outputs(3188) <= not(layer4_outputs(4491));
    layer5_outputs(3189) <= not((layer4_outputs(3201)) and (layer4_outputs(4858)));
    layer5_outputs(3190) <= not(layer4_outputs(1872)) or (layer4_outputs(2943));
    layer5_outputs(3191) <= layer4_outputs(2080);
    layer5_outputs(3192) <= not((layer4_outputs(4601)) or (layer4_outputs(5051)));
    layer5_outputs(3193) <= not((layer4_outputs(1410)) and (layer4_outputs(2336)));
    layer5_outputs(3194) <= not((layer4_outputs(1608)) or (layer4_outputs(66)));
    layer5_outputs(3195) <= not((layer4_outputs(3422)) or (layer4_outputs(303)));
    layer5_outputs(3196) <= not(layer4_outputs(259)) or (layer4_outputs(2339));
    layer5_outputs(3197) <= layer4_outputs(428);
    layer5_outputs(3198) <= not(layer4_outputs(225)) or (layer4_outputs(1344));
    layer5_outputs(3199) <= '0';
    layer5_outputs(3200) <= not((layer4_outputs(2096)) or (layer4_outputs(3573)));
    layer5_outputs(3201) <= (layer4_outputs(1248)) xor (layer4_outputs(4903));
    layer5_outputs(3202) <= layer4_outputs(2);
    layer5_outputs(3203) <= (layer4_outputs(278)) and (layer4_outputs(912));
    layer5_outputs(3204) <= not(layer4_outputs(4091));
    layer5_outputs(3205) <= not((layer4_outputs(1149)) and (layer4_outputs(5059)));
    layer5_outputs(3206) <= (layer4_outputs(3441)) or (layer4_outputs(3072));
    layer5_outputs(3207) <= (layer4_outputs(1216)) and (layer4_outputs(1986));
    layer5_outputs(3208) <= not(layer4_outputs(3819));
    layer5_outputs(3209) <= (layer4_outputs(4648)) and not (layer4_outputs(3162));
    layer5_outputs(3210) <= (layer4_outputs(733)) and (layer4_outputs(1242));
    layer5_outputs(3211) <= not((layer4_outputs(3773)) or (layer4_outputs(2019)));
    layer5_outputs(3212) <= not((layer4_outputs(4667)) xor (layer4_outputs(4674)));
    layer5_outputs(3213) <= (layer4_outputs(5020)) or (layer4_outputs(2474));
    layer5_outputs(3214) <= (layer4_outputs(4241)) and not (layer4_outputs(93));
    layer5_outputs(3215) <= not(layer4_outputs(4368));
    layer5_outputs(3216) <= layer4_outputs(796);
    layer5_outputs(3217) <= layer4_outputs(285);
    layer5_outputs(3218) <= not(layer4_outputs(2640)) or (layer4_outputs(3522));
    layer5_outputs(3219) <= '1';
    layer5_outputs(3220) <= not(layer4_outputs(4515)) or (layer4_outputs(3319));
    layer5_outputs(3221) <= not(layer4_outputs(291)) or (layer4_outputs(2410));
    layer5_outputs(3222) <= layer4_outputs(1696);
    layer5_outputs(3223) <= not(layer4_outputs(4519)) or (layer4_outputs(1821));
    layer5_outputs(3224) <= layer4_outputs(2866);
    layer5_outputs(3225) <= (layer4_outputs(3773)) or (layer4_outputs(3172));
    layer5_outputs(3226) <= not(layer4_outputs(461));
    layer5_outputs(3227) <= layer4_outputs(4401);
    layer5_outputs(3228) <= (layer4_outputs(2059)) and not (layer4_outputs(4409));
    layer5_outputs(3229) <= (layer4_outputs(3007)) xor (layer4_outputs(1194));
    layer5_outputs(3230) <= (layer4_outputs(1402)) or (layer4_outputs(2265));
    layer5_outputs(3231) <= layer4_outputs(1667);
    layer5_outputs(3232) <= not(layer4_outputs(1930)) or (layer4_outputs(4165));
    layer5_outputs(3233) <= not(layer4_outputs(14));
    layer5_outputs(3234) <= not((layer4_outputs(283)) and (layer4_outputs(4583)));
    layer5_outputs(3235) <= (layer4_outputs(1068)) or (layer4_outputs(2024));
    layer5_outputs(3236) <= not(layer4_outputs(1148)) or (layer4_outputs(1453));
    layer5_outputs(3237) <= layer4_outputs(4712);
    layer5_outputs(3238) <= (layer4_outputs(3649)) or (layer4_outputs(2269));
    layer5_outputs(3239) <= not(layer4_outputs(3720)) or (layer4_outputs(4344));
    layer5_outputs(3240) <= layer4_outputs(1259);
    layer5_outputs(3241) <= layer4_outputs(2902);
    layer5_outputs(3242) <= layer4_outputs(3473);
    layer5_outputs(3243) <= '0';
    layer5_outputs(3244) <= '1';
    layer5_outputs(3245) <= '0';
    layer5_outputs(3246) <= not((layer4_outputs(4026)) or (layer4_outputs(2201)));
    layer5_outputs(3247) <= not(layer4_outputs(895)) or (layer4_outputs(245));
    layer5_outputs(3248) <= (layer4_outputs(624)) or (layer4_outputs(4926));
    layer5_outputs(3249) <= not((layer4_outputs(1393)) and (layer4_outputs(3087)));
    layer5_outputs(3250) <= not(layer4_outputs(1329)) or (layer4_outputs(4609));
    layer5_outputs(3251) <= '1';
    layer5_outputs(3252) <= (layer4_outputs(2913)) and not (layer4_outputs(1509));
    layer5_outputs(3253) <= not((layer4_outputs(4461)) and (layer4_outputs(4176)));
    layer5_outputs(3254) <= '0';
    layer5_outputs(3255) <= not(layer4_outputs(1072));
    layer5_outputs(3256) <= not((layer4_outputs(3937)) or (layer4_outputs(119)));
    layer5_outputs(3257) <= not(layer4_outputs(2676));
    layer5_outputs(3258) <= layer4_outputs(3380);
    layer5_outputs(3259) <= layer4_outputs(115);
    layer5_outputs(3260) <= (layer4_outputs(562)) and (layer4_outputs(4150));
    layer5_outputs(3261) <= (layer4_outputs(174)) and (layer4_outputs(3727));
    layer5_outputs(3262) <= not(layer4_outputs(3497));
    layer5_outputs(3263) <= (layer4_outputs(1377)) and (layer4_outputs(3313));
    layer5_outputs(3264) <= layer4_outputs(963);
    layer5_outputs(3265) <= (layer4_outputs(135)) or (layer4_outputs(925));
    layer5_outputs(3266) <= (layer4_outputs(2506)) and (layer4_outputs(2675));
    layer5_outputs(3267) <= not(layer4_outputs(4422));
    layer5_outputs(3268) <= '0';
    layer5_outputs(3269) <= not(layer4_outputs(3795));
    layer5_outputs(3270) <= not(layer4_outputs(173)) or (layer4_outputs(1451));
    layer5_outputs(3271) <= not(layer4_outputs(3510));
    layer5_outputs(3272) <= layer4_outputs(3953);
    layer5_outputs(3273) <= (layer4_outputs(4566)) and (layer4_outputs(1261));
    layer5_outputs(3274) <= not((layer4_outputs(3186)) or (layer4_outputs(1314)));
    layer5_outputs(3275) <= (layer4_outputs(1903)) and not (layer4_outputs(349));
    layer5_outputs(3276) <= not(layer4_outputs(1439)) or (layer4_outputs(3705));
    layer5_outputs(3277) <= (layer4_outputs(2333)) and (layer4_outputs(323));
    layer5_outputs(3278) <= layer4_outputs(2519);
    layer5_outputs(3279) <= not(layer4_outputs(4191));
    layer5_outputs(3280) <= (layer4_outputs(851)) and not (layer4_outputs(3050));
    layer5_outputs(3281) <= layer4_outputs(1081);
    layer5_outputs(3282) <= not(layer4_outputs(1317));
    layer5_outputs(3283) <= layer4_outputs(1338);
    layer5_outputs(3284) <= not(layer4_outputs(1137));
    layer5_outputs(3285) <= not(layer4_outputs(4939));
    layer5_outputs(3286) <= (layer4_outputs(2049)) xor (layer4_outputs(3783));
    layer5_outputs(3287) <= layer4_outputs(1620);
    layer5_outputs(3288) <= (layer4_outputs(687)) and not (layer4_outputs(1720));
    layer5_outputs(3289) <= not((layer4_outputs(2601)) and (layer4_outputs(1052)));
    layer5_outputs(3290) <= (layer4_outputs(2863)) xor (layer4_outputs(3479));
    layer5_outputs(3291) <= not(layer4_outputs(3414)) or (layer4_outputs(150));
    layer5_outputs(3292) <= not((layer4_outputs(2789)) and (layer4_outputs(2895)));
    layer5_outputs(3293) <= layer4_outputs(4775);
    layer5_outputs(3294) <= not((layer4_outputs(1653)) or (layer4_outputs(2386)));
    layer5_outputs(3295) <= layer4_outputs(3345);
    layer5_outputs(3296) <= (layer4_outputs(2207)) and not (layer4_outputs(2978));
    layer5_outputs(3297) <= not(layer4_outputs(3834)) or (layer4_outputs(2967));
    layer5_outputs(3298) <= not(layer4_outputs(4198)) or (layer4_outputs(1444));
    layer5_outputs(3299) <= layer4_outputs(3225);
    layer5_outputs(3300) <= not(layer4_outputs(904));
    layer5_outputs(3301) <= not((layer4_outputs(3901)) or (layer4_outputs(2321)));
    layer5_outputs(3302) <= not(layer4_outputs(3991));
    layer5_outputs(3303) <= not((layer4_outputs(2332)) or (layer4_outputs(4812)));
    layer5_outputs(3304) <= not(layer4_outputs(355));
    layer5_outputs(3305) <= not((layer4_outputs(1611)) xor (layer4_outputs(1070)));
    layer5_outputs(3306) <= layer4_outputs(2396);
    layer5_outputs(3307) <= not(layer4_outputs(18));
    layer5_outputs(3308) <= '1';
    layer5_outputs(3309) <= (layer4_outputs(353)) or (layer4_outputs(1346));
    layer5_outputs(3310) <= (layer4_outputs(280)) or (layer4_outputs(335));
    layer5_outputs(3311) <= not((layer4_outputs(211)) and (layer4_outputs(2144)));
    layer5_outputs(3312) <= not(layer4_outputs(4712)) or (layer4_outputs(2590));
    layer5_outputs(3313) <= not((layer4_outputs(242)) or (layer4_outputs(5003)));
    layer5_outputs(3314) <= (layer4_outputs(1274)) xor (layer4_outputs(3058));
    layer5_outputs(3315) <= (layer4_outputs(1386)) and (layer4_outputs(307));
    layer5_outputs(3316) <= '0';
    layer5_outputs(3317) <= '0';
    layer5_outputs(3318) <= layer4_outputs(464);
    layer5_outputs(3319) <= (layer4_outputs(590)) and (layer4_outputs(3235));
    layer5_outputs(3320) <= (layer4_outputs(3378)) xor (layer4_outputs(90));
    layer5_outputs(3321) <= layer4_outputs(1408);
    layer5_outputs(3322) <= layer4_outputs(4534);
    layer5_outputs(3323) <= (layer4_outputs(3104)) and (layer4_outputs(3112));
    layer5_outputs(3324) <= (layer4_outputs(2874)) and not (layer4_outputs(5044));
    layer5_outputs(3325) <= not((layer4_outputs(2762)) and (layer4_outputs(332)));
    layer5_outputs(3326) <= layer4_outputs(776);
    layer5_outputs(3327) <= not(layer4_outputs(4527)) or (layer4_outputs(4530));
    layer5_outputs(3328) <= not(layer4_outputs(2021));
    layer5_outputs(3329) <= layer4_outputs(4319);
    layer5_outputs(3330) <= not(layer4_outputs(1568));
    layer5_outputs(3331) <= not(layer4_outputs(4756)) or (layer4_outputs(3508));
    layer5_outputs(3332) <= layer4_outputs(2337);
    layer5_outputs(3333) <= not(layer4_outputs(962));
    layer5_outputs(3334) <= not(layer4_outputs(3113));
    layer5_outputs(3335) <= layer4_outputs(500);
    layer5_outputs(3336) <= not(layer4_outputs(385)) or (layer4_outputs(3137));
    layer5_outputs(3337) <= (layer4_outputs(512)) and (layer4_outputs(3922));
    layer5_outputs(3338) <= (layer4_outputs(548)) and (layer4_outputs(182));
    layer5_outputs(3339) <= (layer4_outputs(1622)) and not (layer4_outputs(3495));
    layer5_outputs(3340) <= (layer4_outputs(3367)) and not (layer4_outputs(1543));
    layer5_outputs(3341) <= not(layer4_outputs(3787));
    layer5_outputs(3342) <= layer4_outputs(1140);
    layer5_outputs(3343) <= not(layer4_outputs(620));
    layer5_outputs(3344) <= (layer4_outputs(1511)) or (layer4_outputs(3390));
    layer5_outputs(3345) <= layer4_outputs(982);
    layer5_outputs(3346) <= layer4_outputs(2124);
    layer5_outputs(3347) <= not(layer4_outputs(372)) or (layer4_outputs(1177));
    layer5_outputs(3348) <= '1';
    layer5_outputs(3349) <= not(layer4_outputs(1861)) or (layer4_outputs(106));
    layer5_outputs(3350) <= (layer4_outputs(3549)) and (layer4_outputs(4700));
    layer5_outputs(3351) <= not(layer4_outputs(2988));
    layer5_outputs(3352) <= '0';
    layer5_outputs(3353) <= not((layer4_outputs(1232)) and (layer4_outputs(538)));
    layer5_outputs(3354) <= layer4_outputs(4299);
    layer5_outputs(3355) <= not((layer4_outputs(5018)) and (layer4_outputs(3596)));
    layer5_outputs(3356) <= layer4_outputs(247);
    layer5_outputs(3357) <= not(layer4_outputs(4750));
    layer5_outputs(3358) <= (layer4_outputs(1583)) and not (layer4_outputs(2007));
    layer5_outputs(3359) <= not(layer4_outputs(4309)) or (layer4_outputs(5010));
    layer5_outputs(3360) <= not(layer4_outputs(1790));
    layer5_outputs(3361) <= (layer4_outputs(4279)) or (layer4_outputs(4698));
    layer5_outputs(3362) <= not(layer4_outputs(267));
    layer5_outputs(3363) <= '1';
    layer5_outputs(3364) <= not((layer4_outputs(2535)) and (layer4_outputs(3731)));
    layer5_outputs(3365) <= (layer4_outputs(656)) and not (layer4_outputs(872));
    layer5_outputs(3366) <= '1';
    layer5_outputs(3367) <= (layer4_outputs(3128)) and (layer4_outputs(1959));
    layer5_outputs(3368) <= (layer4_outputs(1526)) or (layer4_outputs(1647));
    layer5_outputs(3369) <= (layer4_outputs(5088)) and not (layer4_outputs(4852));
    layer5_outputs(3370) <= (layer4_outputs(4847)) and not (layer4_outputs(168));
    layer5_outputs(3371) <= (layer4_outputs(965)) and not (layer4_outputs(2998));
    layer5_outputs(3372) <= not(layer4_outputs(2557)) or (layer4_outputs(1733));
    layer5_outputs(3373) <= layer4_outputs(4134);
    layer5_outputs(3374) <= '0';
    layer5_outputs(3375) <= (layer4_outputs(3110)) and not (layer4_outputs(1979));
    layer5_outputs(3376) <= layer4_outputs(1753);
    layer5_outputs(3377) <= (layer4_outputs(1951)) and not (layer4_outputs(1142));
    layer5_outputs(3378) <= (layer4_outputs(110)) and not (layer4_outputs(2161));
    layer5_outputs(3379) <= not(layer4_outputs(2148)) or (layer4_outputs(4517));
    layer5_outputs(3380) <= (layer4_outputs(779)) and (layer4_outputs(4327));
    layer5_outputs(3381) <= not(layer4_outputs(3345));
    layer5_outputs(3382) <= (layer4_outputs(1453)) or (layer4_outputs(3668));
    layer5_outputs(3383) <= layer4_outputs(592);
    layer5_outputs(3384) <= not(layer4_outputs(1660));
    layer5_outputs(3385) <= layer4_outputs(3708);
    layer5_outputs(3386) <= not(layer4_outputs(2879));
    layer5_outputs(3387) <= (layer4_outputs(379)) xor (layer4_outputs(4453));
    layer5_outputs(3388) <= '1';
    layer5_outputs(3389) <= (layer4_outputs(1489)) and not (layer4_outputs(1754));
    layer5_outputs(3390) <= not(layer4_outputs(3817)) or (layer4_outputs(3715));
    layer5_outputs(3391) <= layer4_outputs(99);
    layer5_outputs(3392) <= (layer4_outputs(4265)) and (layer4_outputs(4495));
    layer5_outputs(3393) <= (layer4_outputs(1451)) xor (layer4_outputs(483));
    layer5_outputs(3394) <= not(layer4_outputs(3847)) or (layer4_outputs(3912));
    layer5_outputs(3395) <= layer4_outputs(1550);
    layer5_outputs(3396) <= (layer4_outputs(2473)) and (layer4_outputs(1311));
    layer5_outputs(3397) <= (layer4_outputs(1526)) and not (layer4_outputs(2797));
    layer5_outputs(3398) <= not(layer4_outputs(4736));
    layer5_outputs(3399) <= not(layer4_outputs(3944));
    layer5_outputs(3400) <= layer4_outputs(2802);
    layer5_outputs(3401) <= '1';
    layer5_outputs(3402) <= not(layer4_outputs(2040)) or (layer4_outputs(731));
    layer5_outputs(3403) <= not(layer4_outputs(668));
    layer5_outputs(3404) <= not(layer4_outputs(4004));
    layer5_outputs(3405) <= not(layer4_outputs(4880)) or (layer4_outputs(483));
    layer5_outputs(3406) <= not((layer4_outputs(2163)) or (layer4_outputs(3537)));
    layer5_outputs(3407) <= not(layer4_outputs(4833)) or (layer4_outputs(276));
    layer5_outputs(3408) <= (layer4_outputs(5059)) and not (layer4_outputs(2458));
    layer5_outputs(3409) <= not(layer4_outputs(1804));
    layer5_outputs(3410) <= not(layer4_outputs(1686)) or (layer4_outputs(541));
    layer5_outputs(3411) <= (layer4_outputs(4694)) and not (layer4_outputs(185));
    layer5_outputs(3412) <= (layer4_outputs(2727)) or (layer4_outputs(1277));
    layer5_outputs(3413) <= not(layer4_outputs(2468));
    layer5_outputs(3414) <= (layer4_outputs(3481)) and not (layer4_outputs(565));
    layer5_outputs(3415) <= layer4_outputs(4978);
    layer5_outputs(3416) <= not((layer4_outputs(867)) or (layer4_outputs(1935)));
    layer5_outputs(3417) <= not(layer4_outputs(5090));
    layer5_outputs(3418) <= (layer4_outputs(1606)) and not (layer4_outputs(4450));
    layer5_outputs(3419) <= (layer4_outputs(1126)) and (layer4_outputs(1403));
    layer5_outputs(3420) <= (layer4_outputs(4100)) and not (layer4_outputs(3466));
    layer5_outputs(3421) <= not(layer4_outputs(3460));
    layer5_outputs(3422) <= layer4_outputs(3886);
    layer5_outputs(3423) <= layer4_outputs(2444);
    layer5_outputs(3424) <= (layer4_outputs(480)) and (layer4_outputs(1151));
    layer5_outputs(3425) <= layer4_outputs(3097);
    layer5_outputs(3426) <= layer4_outputs(4720);
    layer5_outputs(3427) <= not((layer4_outputs(728)) and (layer4_outputs(2032)));
    layer5_outputs(3428) <= not(layer4_outputs(4669)) or (layer4_outputs(5058));
    layer5_outputs(3429) <= (layer4_outputs(4781)) and not (layer4_outputs(662));
    layer5_outputs(3430) <= not(layer4_outputs(3529)) or (layer4_outputs(2172));
    layer5_outputs(3431) <= not((layer4_outputs(3513)) or (layer4_outputs(1525)));
    layer5_outputs(3432) <= (layer4_outputs(1231)) and not (layer4_outputs(3728));
    layer5_outputs(3433) <= '0';
    layer5_outputs(3434) <= layer4_outputs(1038);
    layer5_outputs(3435) <= '0';
    layer5_outputs(3436) <= layer4_outputs(4936);
    layer5_outputs(3437) <= layer4_outputs(4856);
    layer5_outputs(3438) <= not((layer4_outputs(1219)) and (layer4_outputs(2492)));
    layer5_outputs(3439) <= '0';
    layer5_outputs(3440) <= not((layer4_outputs(4596)) or (layer4_outputs(2252)));
    layer5_outputs(3441) <= (layer4_outputs(4559)) or (layer4_outputs(81));
    layer5_outputs(3442) <= not(layer4_outputs(3131));
    layer5_outputs(3443) <= (layer4_outputs(574)) and (layer4_outputs(4789));
    layer5_outputs(3444) <= layer4_outputs(2206);
    layer5_outputs(3445) <= not(layer4_outputs(309));
    layer5_outputs(3446) <= layer4_outputs(2892);
    layer5_outputs(3447) <= (layer4_outputs(4270)) xor (layer4_outputs(4606));
    layer5_outputs(3448) <= not((layer4_outputs(1587)) and (layer4_outputs(1530)));
    layer5_outputs(3449) <= layer4_outputs(661);
    layer5_outputs(3450) <= layer4_outputs(4826);
    layer5_outputs(3451) <= (layer4_outputs(3901)) and not (layer4_outputs(1787));
    layer5_outputs(3452) <= not(layer4_outputs(4798)) or (layer4_outputs(3356));
    layer5_outputs(3453) <= not((layer4_outputs(4038)) and (layer4_outputs(455)));
    layer5_outputs(3454) <= not(layer4_outputs(1409));
    layer5_outputs(3455) <= not((layer4_outputs(224)) or (layer4_outputs(3182)));
    layer5_outputs(3456) <= (layer4_outputs(2771)) and not (layer4_outputs(950));
    layer5_outputs(3457) <= (layer4_outputs(2844)) xor (layer4_outputs(620));
    layer5_outputs(3458) <= not(layer4_outputs(3284)) or (layer4_outputs(1168));
    layer5_outputs(3459) <= not((layer4_outputs(2203)) or (layer4_outputs(4163)));
    layer5_outputs(3460) <= not(layer4_outputs(4691)) or (layer4_outputs(3366));
    layer5_outputs(3461) <= not(layer4_outputs(4453)) or (layer4_outputs(2794));
    layer5_outputs(3462) <= not((layer4_outputs(1158)) and (layer4_outputs(1482)));
    layer5_outputs(3463) <= not(layer4_outputs(2261));
    layer5_outputs(3464) <= (layer4_outputs(4099)) or (layer4_outputs(1343));
    layer5_outputs(3465) <= not(layer4_outputs(4417));
    layer5_outputs(3466) <= not(layer4_outputs(3833));
    layer5_outputs(3467) <= not(layer4_outputs(467)) or (layer4_outputs(629));
    layer5_outputs(3468) <= '1';
    layer5_outputs(3469) <= layer4_outputs(4348);
    layer5_outputs(3470) <= not((layer4_outputs(4909)) or (layer4_outputs(960)));
    layer5_outputs(3471) <= (layer4_outputs(1843)) and not (layer4_outputs(1470));
    layer5_outputs(3472) <= '1';
    layer5_outputs(3473) <= (layer4_outputs(891)) and not (layer4_outputs(2113));
    layer5_outputs(3474) <= layer4_outputs(3241);
    layer5_outputs(3475) <= not(layer4_outputs(3));
    layer5_outputs(3476) <= not((layer4_outputs(3015)) and (layer4_outputs(365)));
    layer5_outputs(3477) <= '1';
    layer5_outputs(3478) <= '0';
    layer5_outputs(3479) <= not(layer4_outputs(1713));
    layer5_outputs(3480) <= (layer4_outputs(5098)) and not (layer4_outputs(4693));
    layer5_outputs(3481) <= not((layer4_outputs(3395)) and (layer4_outputs(3403)));
    layer5_outputs(3482) <= '0';
    layer5_outputs(3483) <= (layer4_outputs(4346)) and (layer4_outputs(899));
    layer5_outputs(3484) <= not((layer4_outputs(972)) or (layer4_outputs(1614)));
    layer5_outputs(3485) <= (layer4_outputs(4839)) and not (layer4_outputs(2847));
    layer5_outputs(3486) <= (layer4_outputs(1319)) and not (layer4_outputs(1404));
    layer5_outputs(3487) <= (layer4_outputs(44)) and (layer4_outputs(732));
    layer5_outputs(3488) <= (layer4_outputs(2048)) or (layer4_outputs(2518));
    layer5_outputs(3489) <= not((layer4_outputs(5011)) and (layer4_outputs(197)));
    layer5_outputs(3490) <= not((layer4_outputs(790)) and (layer4_outputs(2883)));
    layer5_outputs(3491) <= not((layer4_outputs(2684)) and (layer4_outputs(2329)));
    layer5_outputs(3492) <= '1';
    layer5_outputs(3493) <= '0';
    layer5_outputs(3494) <= not(layer4_outputs(4752)) or (layer4_outputs(2722));
    layer5_outputs(3495) <= (layer4_outputs(1432)) or (layer4_outputs(514));
    layer5_outputs(3496) <= layer4_outputs(2169);
    layer5_outputs(3497) <= not(layer4_outputs(4749)) or (layer4_outputs(129));
    layer5_outputs(3498) <= not(layer4_outputs(236));
    layer5_outputs(3499) <= not((layer4_outputs(3893)) xor (layer4_outputs(1209)));
    layer5_outputs(3500) <= '1';
    layer5_outputs(3501) <= not(layer4_outputs(2905)) or (layer4_outputs(3818));
    layer5_outputs(3502) <= not(layer4_outputs(1419)) or (layer4_outputs(4717));
    layer5_outputs(3503) <= '1';
    layer5_outputs(3504) <= (layer4_outputs(975)) and not (layer4_outputs(1115));
    layer5_outputs(3505) <= (layer4_outputs(3004)) and not (layer4_outputs(1034));
    layer5_outputs(3506) <= not(layer4_outputs(4627));
    layer5_outputs(3507) <= not(layer4_outputs(2213));
    layer5_outputs(3508) <= not(layer4_outputs(2948));
    layer5_outputs(3509) <= (layer4_outputs(3335)) or (layer4_outputs(2982));
    layer5_outputs(3510) <= not(layer4_outputs(1842));
    layer5_outputs(3511) <= layer4_outputs(2557);
    layer5_outputs(3512) <= not(layer4_outputs(787));
    layer5_outputs(3513) <= (layer4_outputs(597)) and (layer4_outputs(4589));
    layer5_outputs(3514) <= not(layer4_outputs(3626));
    layer5_outputs(3515) <= layer4_outputs(3845);
    layer5_outputs(3516) <= not(layer4_outputs(3234));
    layer5_outputs(3517) <= layer4_outputs(4560);
    layer5_outputs(3518) <= layer4_outputs(1039);
    layer5_outputs(3519) <= layer4_outputs(4306);
    layer5_outputs(3520) <= layer4_outputs(2732);
    layer5_outputs(3521) <= (layer4_outputs(2095)) and not (layer4_outputs(1108));
    layer5_outputs(3522) <= layer4_outputs(207);
    layer5_outputs(3523) <= not(layer4_outputs(4070)) or (layer4_outputs(3665));
    layer5_outputs(3524) <= not((layer4_outputs(1350)) or (layer4_outputs(417)));
    layer5_outputs(3525) <= layer4_outputs(1917);
    layer5_outputs(3526) <= not(layer4_outputs(476));
    layer5_outputs(3527) <= not(layer4_outputs(760)) or (layer4_outputs(947));
    layer5_outputs(3528) <= not((layer4_outputs(1121)) and (layer4_outputs(222)));
    layer5_outputs(3529) <= (layer4_outputs(1638)) and (layer4_outputs(1032));
    layer5_outputs(3530) <= '1';
    layer5_outputs(3531) <= layer4_outputs(822);
    layer5_outputs(3532) <= '0';
    layer5_outputs(3533) <= layer4_outputs(645);
    layer5_outputs(3534) <= (layer4_outputs(2283)) and (layer4_outputs(2806));
    layer5_outputs(3535) <= not((layer4_outputs(2631)) and (layer4_outputs(4357)));
    layer5_outputs(3536) <= (layer4_outputs(307)) or (layer4_outputs(3791));
    layer5_outputs(3537) <= not((layer4_outputs(4619)) and (layer4_outputs(1747)));
    layer5_outputs(3538) <= (layer4_outputs(2893)) and not (layer4_outputs(937));
    layer5_outputs(3539) <= not((layer4_outputs(5048)) and (layer4_outputs(1307)));
    layer5_outputs(3540) <= layer4_outputs(2326);
    layer5_outputs(3541) <= layer4_outputs(1422);
    layer5_outputs(3542) <= (layer4_outputs(40)) xor (layer4_outputs(2453));
    layer5_outputs(3543) <= layer4_outputs(1022);
    layer5_outputs(3544) <= not((layer4_outputs(4278)) or (layer4_outputs(524)));
    layer5_outputs(3545) <= layer4_outputs(621);
    layer5_outputs(3546) <= not(layer4_outputs(3557));
    layer5_outputs(3547) <= not(layer4_outputs(221));
    layer5_outputs(3548) <= not((layer4_outputs(4540)) and (layer4_outputs(4518)));
    layer5_outputs(3549) <= not(layer4_outputs(1649)) or (layer4_outputs(2370));
    layer5_outputs(3550) <= not((layer4_outputs(1427)) and (layer4_outputs(3857)));
    layer5_outputs(3551) <= not(layer4_outputs(3431));
    layer5_outputs(3552) <= not(layer4_outputs(3893));
    layer5_outputs(3553) <= (layer4_outputs(3627)) and not (layer4_outputs(4076));
    layer5_outputs(3554) <= layer4_outputs(3850);
    layer5_outputs(3555) <= not((layer4_outputs(447)) xor (layer4_outputs(4445)));
    layer5_outputs(3556) <= not(layer4_outputs(2661));
    layer5_outputs(3557) <= (layer4_outputs(2599)) and not (layer4_outputs(2908));
    layer5_outputs(3558) <= not(layer4_outputs(2773));
    layer5_outputs(3559) <= (layer4_outputs(4568)) and not (layer4_outputs(918));
    layer5_outputs(3560) <= not(layer4_outputs(4386));
    layer5_outputs(3561) <= not(layer4_outputs(4550));
    layer5_outputs(3562) <= (layer4_outputs(4403)) xor (layer4_outputs(3253));
    layer5_outputs(3563) <= (layer4_outputs(2177)) and (layer4_outputs(2552));
    layer5_outputs(3564) <= not(layer4_outputs(4974));
    layer5_outputs(3565) <= not((layer4_outputs(250)) and (layer4_outputs(469)));
    layer5_outputs(3566) <= not(layer4_outputs(334));
    layer5_outputs(3567) <= layer4_outputs(1496);
    layer5_outputs(3568) <= (layer4_outputs(2746)) and not (layer4_outputs(740));
    layer5_outputs(3569) <= not((layer4_outputs(3123)) xor (layer4_outputs(4639)));
    layer5_outputs(3570) <= not(layer4_outputs(1546)) or (layer4_outputs(3437));
    layer5_outputs(3571) <= not((layer4_outputs(36)) and (layer4_outputs(4842)));
    layer5_outputs(3572) <= not(layer4_outputs(3250));
    layer5_outputs(3573) <= '0';
    layer5_outputs(3574) <= (layer4_outputs(4230)) or (layer4_outputs(2699));
    layer5_outputs(3575) <= (layer4_outputs(73)) and (layer4_outputs(2987));
    layer5_outputs(3576) <= not(layer4_outputs(3080));
    layer5_outputs(3577) <= not(layer4_outputs(3660));
    layer5_outputs(3578) <= layer4_outputs(4659);
    layer5_outputs(3579) <= layer4_outputs(753);
    layer5_outputs(3580) <= not(layer4_outputs(416));
    layer5_outputs(3581) <= not(layer4_outputs(2340));
    layer5_outputs(3582) <= not(layer4_outputs(2079));
    layer5_outputs(3583) <= (layer4_outputs(167)) and not (layer4_outputs(4310));
    layer5_outputs(3584) <= layer4_outputs(3508);
    layer5_outputs(3585) <= not(layer4_outputs(3232)) or (layer4_outputs(144));
    layer5_outputs(3586) <= '0';
    layer5_outputs(3587) <= (layer4_outputs(4215)) and (layer4_outputs(4987));
    layer5_outputs(3588) <= (layer4_outputs(4953)) and (layer4_outputs(1602));
    layer5_outputs(3589) <= '0';
    layer5_outputs(3590) <= not((layer4_outputs(4816)) and (layer4_outputs(40)));
    layer5_outputs(3591) <= '1';
    layer5_outputs(3592) <= layer4_outputs(4551);
    layer5_outputs(3593) <= (layer4_outputs(3836)) and (layer4_outputs(3793));
    layer5_outputs(3594) <= (layer4_outputs(394)) and not (layer4_outputs(4243));
    layer5_outputs(3595) <= not(layer4_outputs(480));
    layer5_outputs(3596) <= not(layer4_outputs(2264));
    layer5_outputs(3597) <= not(layer4_outputs(1276));
    layer5_outputs(3598) <= layer4_outputs(2350);
    layer5_outputs(3599) <= layer4_outputs(3835);
    layer5_outputs(3600) <= not(layer4_outputs(518));
    layer5_outputs(3601) <= (layer4_outputs(4657)) and (layer4_outputs(33));
    layer5_outputs(3602) <= (layer4_outputs(3652)) and not (layer4_outputs(3586));
    layer5_outputs(3603) <= not(layer4_outputs(503));
    layer5_outputs(3604) <= layer4_outputs(838);
    layer5_outputs(3605) <= layer4_outputs(3296);
    layer5_outputs(3606) <= not((layer4_outputs(3796)) or (layer4_outputs(1545)));
    layer5_outputs(3607) <= not((layer4_outputs(2735)) and (layer4_outputs(3868)));
    layer5_outputs(3608) <= not(layer4_outputs(3287)) or (layer4_outputs(3472));
    layer5_outputs(3609) <= not(layer4_outputs(3184));
    layer5_outputs(3610) <= '0';
    layer5_outputs(3611) <= not((layer4_outputs(3049)) xor (layer4_outputs(1221)));
    layer5_outputs(3612) <= (layer4_outputs(3532)) and not (layer4_outputs(3559));
    layer5_outputs(3613) <= layer4_outputs(2830);
    layer5_outputs(3614) <= layer4_outputs(714);
    layer5_outputs(3615) <= (layer4_outputs(212)) and not (layer4_outputs(6));
    layer5_outputs(3616) <= not((layer4_outputs(2733)) and (layer4_outputs(3934)));
    layer5_outputs(3617) <= layer4_outputs(532);
    layer5_outputs(3618) <= not((layer4_outputs(2485)) or (layer4_outputs(2829)));
    layer5_outputs(3619) <= (layer4_outputs(4241)) and (layer4_outputs(4220));
    layer5_outputs(3620) <= (layer4_outputs(1440)) or (layer4_outputs(2815));
    layer5_outputs(3621) <= '1';
    layer5_outputs(3622) <= layer4_outputs(1097);
    layer5_outputs(3623) <= not((layer4_outputs(2173)) or (layer4_outputs(2976)));
    layer5_outputs(3624) <= (layer4_outputs(3295)) xor (layer4_outputs(3167));
    layer5_outputs(3625) <= (layer4_outputs(58)) and (layer4_outputs(2152));
    layer5_outputs(3626) <= (layer4_outputs(1177)) and (layer4_outputs(1265));
    layer5_outputs(3627) <= not((layer4_outputs(4060)) and (layer4_outputs(4256)));
    layer5_outputs(3628) <= '1';
    layer5_outputs(3629) <= (layer4_outputs(3297)) and (layer4_outputs(3175));
    layer5_outputs(3630) <= not(layer4_outputs(1155));
    layer5_outputs(3631) <= (layer4_outputs(3744)) xor (layer4_outputs(585));
    layer5_outputs(3632) <= not(layer4_outputs(3396));
    layer5_outputs(3633) <= not(layer4_outputs(4103));
    layer5_outputs(3634) <= not(layer4_outputs(1456)) or (layer4_outputs(2541));
    layer5_outputs(3635) <= not(layer4_outputs(3521));
    layer5_outputs(3636) <= (layer4_outputs(462)) xor (layer4_outputs(3016));
    layer5_outputs(3637) <= (layer4_outputs(4012)) and (layer4_outputs(4331));
    layer5_outputs(3638) <= layer4_outputs(1312);
    layer5_outputs(3639) <= (layer4_outputs(3324)) and not (layer4_outputs(1143));
    layer5_outputs(3640) <= not((layer4_outputs(5106)) and (layer4_outputs(2968)));
    layer5_outputs(3641) <= (layer4_outputs(4298)) and not (layer4_outputs(5047));
    layer5_outputs(3642) <= layer4_outputs(2769);
    layer5_outputs(3643) <= not(layer4_outputs(4165)) or (layer4_outputs(219));
    layer5_outputs(3644) <= layer4_outputs(920);
    layer5_outputs(3645) <= layer4_outputs(1275);
    layer5_outputs(3646) <= not(layer4_outputs(4521));
    layer5_outputs(3647) <= (layer4_outputs(2581)) and not (layer4_outputs(4382));
    layer5_outputs(3648) <= not(layer4_outputs(3699));
    layer5_outputs(3649) <= layer4_outputs(2540);
    layer5_outputs(3650) <= not(layer4_outputs(4924));
    layer5_outputs(3651) <= (layer4_outputs(774)) and not (layer4_outputs(2623));
    layer5_outputs(3652) <= '1';
    layer5_outputs(3653) <= not((layer4_outputs(4442)) and (layer4_outputs(4689)));
    layer5_outputs(3654) <= not(layer4_outputs(2695));
    layer5_outputs(3655) <= not((layer4_outputs(3350)) and (layer4_outputs(318)));
    layer5_outputs(3656) <= '1';
    layer5_outputs(3657) <= layer4_outputs(4968);
    layer5_outputs(3658) <= layer4_outputs(4950);
    layer5_outputs(3659) <= (layer4_outputs(4526)) and (layer4_outputs(4925));
    layer5_outputs(3660) <= layer4_outputs(642);
    layer5_outputs(3661) <= not((layer4_outputs(109)) and (layer4_outputs(1351)));
    layer5_outputs(3662) <= (layer4_outputs(2586)) and not (layer4_outputs(4803));
    layer5_outputs(3663) <= not(layer4_outputs(3437)) or (layer4_outputs(22));
    layer5_outputs(3664) <= not((layer4_outputs(3493)) or (layer4_outputs(4571)));
    layer5_outputs(3665) <= (layer4_outputs(1731)) or (layer4_outputs(716));
    layer5_outputs(3666) <= not(layer4_outputs(4724)) or (layer4_outputs(4354));
    layer5_outputs(3667) <= not(layer4_outputs(4718)) or (layer4_outputs(2097));
    layer5_outputs(3668) <= not(layer4_outputs(791));
    layer5_outputs(3669) <= not(layer4_outputs(25));
    layer5_outputs(3670) <= not(layer4_outputs(3268));
    layer5_outputs(3671) <= layer4_outputs(426);
    layer5_outputs(3672) <= (layer4_outputs(1592)) and not (layer4_outputs(660));
    layer5_outputs(3673) <= layer4_outputs(4667);
    layer5_outputs(3674) <= not((layer4_outputs(1758)) xor (layer4_outputs(3287)));
    layer5_outputs(3675) <= layer4_outputs(983);
    layer5_outputs(3676) <= layer4_outputs(1315);
    layer5_outputs(3677) <= layer4_outputs(1433);
    layer5_outputs(3678) <= not(layer4_outputs(2249));
    layer5_outputs(3679) <= layer4_outputs(3672);
    layer5_outputs(3680) <= (layer4_outputs(48)) and not (layer4_outputs(662));
    layer5_outputs(3681) <= layer4_outputs(855);
    layer5_outputs(3682) <= (layer4_outputs(59)) and (layer4_outputs(3042));
    layer5_outputs(3683) <= not((layer4_outputs(1009)) or (layer4_outputs(3991)));
    layer5_outputs(3684) <= '0';
    layer5_outputs(3685) <= layer4_outputs(4263);
    layer5_outputs(3686) <= not((layer4_outputs(2019)) or (layer4_outputs(1950)));
    layer5_outputs(3687) <= not(layer4_outputs(1007));
    layer5_outputs(3688) <= (layer4_outputs(1992)) and (layer4_outputs(1740));
    layer5_outputs(3689) <= layer4_outputs(3969);
    layer5_outputs(3690) <= not(layer4_outputs(3839)) or (layer4_outputs(2236));
    layer5_outputs(3691) <= (layer4_outputs(989)) xor (layer4_outputs(539));
    layer5_outputs(3692) <= layer4_outputs(3075);
    layer5_outputs(3693) <= (layer4_outputs(2427)) and (layer4_outputs(760));
    layer5_outputs(3694) <= '0';
    layer5_outputs(3695) <= '1';
    layer5_outputs(3696) <= '1';
    layer5_outputs(3697) <= not(layer4_outputs(4571));
    layer5_outputs(3698) <= (layer4_outputs(3578)) and (layer4_outputs(3833));
    layer5_outputs(3699) <= '0';
    layer5_outputs(3700) <= (layer4_outputs(4882)) and (layer4_outputs(1117));
    layer5_outputs(3701) <= not(layer4_outputs(997));
    layer5_outputs(3702) <= not((layer4_outputs(205)) xor (layer4_outputs(4590)));
    layer5_outputs(3703) <= layer4_outputs(1624);
    layer5_outputs(3704) <= layer4_outputs(4556);
    layer5_outputs(3705) <= not((layer4_outputs(517)) and (layer4_outputs(1085)));
    layer5_outputs(3706) <= '1';
    layer5_outputs(3707) <= not((layer4_outputs(4280)) or (layer4_outputs(5066)));
    layer5_outputs(3708) <= '1';
    layer5_outputs(3709) <= not(layer4_outputs(2888));
    layer5_outputs(3710) <= (layer4_outputs(487)) and (layer4_outputs(3982));
    layer5_outputs(3711) <= not(layer4_outputs(1589)) or (layer4_outputs(46));
    layer5_outputs(3712) <= (layer4_outputs(3357)) or (layer4_outputs(55));
    layer5_outputs(3713) <= (layer4_outputs(643)) and not (layer4_outputs(4242));
    layer5_outputs(3714) <= (layer4_outputs(1727)) and not (layer4_outputs(1220));
    layer5_outputs(3715) <= layer4_outputs(3494);
    layer5_outputs(3716) <= not(layer4_outputs(5042)) or (layer4_outputs(2850));
    layer5_outputs(3717) <= not(layer4_outputs(2222)) or (layer4_outputs(1015));
    layer5_outputs(3718) <= layer4_outputs(2719);
    layer5_outputs(3719) <= (layer4_outputs(102)) and (layer4_outputs(3065));
    layer5_outputs(3720) <= not((layer4_outputs(3108)) or (layer4_outputs(3191)));
    layer5_outputs(3721) <= (layer4_outputs(4260)) xor (layer4_outputs(5034));
    layer5_outputs(3722) <= not((layer4_outputs(4006)) and (layer4_outputs(1752)));
    layer5_outputs(3723) <= (layer4_outputs(4312)) or (layer4_outputs(4410));
    layer5_outputs(3724) <= (layer4_outputs(2138)) and not (layer4_outputs(1734));
    layer5_outputs(3725) <= layer4_outputs(5067);
    layer5_outputs(3726) <= not(layer4_outputs(2574)) or (layer4_outputs(3938));
    layer5_outputs(3727) <= (layer4_outputs(2880)) and not (layer4_outputs(392));
    layer5_outputs(3728) <= (layer4_outputs(2232)) and (layer4_outputs(3298));
    layer5_outputs(3729) <= not(layer4_outputs(2725));
    layer5_outputs(3730) <= layer4_outputs(4906);
    layer5_outputs(3731) <= layer4_outputs(3402);
    layer5_outputs(3732) <= not(layer4_outputs(1171));
    layer5_outputs(3733) <= layer4_outputs(2793);
    layer5_outputs(3734) <= not(layer4_outputs(2286)) or (layer4_outputs(267));
    layer5_outputs(3735) <= not(layer4_outputs(3569));
    layer5_outputs(3736) <= (layer4_outputs(140)) xor (layer4_outputs(1956));
    layer5_outputs(3737) <= '0';
    layer5_outputs(3738) <= '1';
    layer5_outputs(3739) <= not((layer4_outputs(2709)) and (layer4_outputs(1817)));
    layer5_outputs(3740) <= (layer4_outputs(692)) and (layer4_outputs(1597));
    layer5_outputs(3741) <= '1';
    layer5_outputs(3742) <= not((layer4_outputs(2422)) and (layer4_outputs(83)));
    layer5_outputs(3743) <= layer4_outputs(1441);
    layer5_outputs(3744) <= (layer4_outputs(5025)) and not (layer4_outputs(2958));
    layer5_outputs(3745) <= not(layer4_outputs(1332)) or (layer4_outputs(2187));
    layer5_outputs(3746) <= layer4_outputs(1374);
    layer5_outputs(3747) <= not(layer4_outputs(3126)) or (layer4_outputs(609));
    layer5_outputs(3748) <= (layer4_outputs(4705)) and not (layer4_outputs(4733));
    layer5_outputs(3749) <= layer4_outputs(2670);
    layer5_outputs(3750) <= (layer4_outputs(4394)) and not (layer4_outputs(295));
    layer5_outputs(3751) <= (layer4_outputs(3476)) xor (layer4_outputs(1845));
    layer5_outputs(3752) <= not(layer4_outputs(3071)) or (layer4_outputs(2926));
    layer5_outputs(3753) <= not(layer4_outputs(3838));
    layer5_outputs(3754) <= '1';
    layer5_outputs(3755) <= not((layer4_outputs(3435)) and (layer4_outputs(1273)));
    layer5_outputs(3756) <= not(layer4_outputs(2554));
    layer5_outputs(3757) <= not(layer4_outputs(1651)) or (layer4_outputs(2443));
    layer5_outputs(3758) <= not(layer4_outputs(3361)) or (layer4_outputs(4030));
    layer5_outputs(3759) <= (layer4_outputs(4411)) or (layer4_outputs(4785));
    layer5_outputs(3760) <= (layer4_outputs(1711)) and not (layer4_outputs(2643));
    layer5_outputs(3761) <= '0';
    layer5_outputs(3762) <= (layer4_outputs(2225)) and (layer4_outputs(2382));
    layer5_outputs(3763) <= (layer4_outputs(2100)) and not (layer4_outputs(2380));
    layer5_outputs(3764) <= not(layer4_outputs(644));
    layer5_outputs(3765) <= not(layer4_outputs(2899)) or (layer4_outputs(1518));
    layer5_outputs(3766) <= not(layer4_outputs(368));
    layer5_outputs(3767) <= not(layer4_outputs(5078));
    layer5_outputs(3768) <= not((layer4_outputs(2866)) or (layer4_outputs(4884)));
    layer5_outputs(3769) <= not(layer4_outputs(2484)) or (layer4_outputs(357));
    layer5_outputs(3770) <= layer4_outputs(4930);
    layer5_outputs(3771) <= not(layer4_outputs(4755)) or (layer4_outputs(4660));
    layer5_outputs(3772) <= (layer4_outputs(4420)) and not (layer4_outputs(2717));
    layer5_outputs(3773) <= (layer4_outputs(1522)) and (layer4_outputs(3406));
    layer5_outputs(3774) <= layer4_outputs(151);
    layer5_outputs(3775) <= not((layer4_outputs(3211)) or (layer4_outputs(618)));
    layer5_outputs(3776) <= (layer4_outputs(2609)) or (layer4_outputs(1336));
    layer5_outputs(3777) <= (layer4_outputs(1106)) and (layer4_outputs(76));
    layer5_outputs(3778) <= not((layer4_outputs(3919)) and (layer4_outputs(2703)));
    layer5_outputs(3779) <= not(layer4_outputs(2680)) or (layer4_outputs(3848));
    layer5_outputs(3780) <= (layer4_outputs(3426)) and not (layer4_outputs(2290));
    layer5_outputs(3781) <= not((layer4_outputs(5004)) or (layer4_outputs(3261)));
    layer5_outputs(3782) <= not(layer4_outputs(490));
    layer5_outputs(3783) <= layer4_outputs(1690);
    layer5_outputs(3784) <= '0';
    layer5_outputs(3785) <= (layer4_outputs(4906)) and not (layer4_outputs(1103));
    layer5_outputs(3786) <= not(layer4_outputs(2471));
    layer5_outputs(3787) <= not(layer4_outputs(1868));
    layer5_outputs(3788) <= not(layer4_outputs(2901));
    layer5_outputs(3789) <= (layer4_outputs(3338)) and not (layer4_outputs(1165));
    layer5_outputs(3790) <= not(layer4_outputs(740));
    layer5_outputs(3791) <= not((layer4_outputs(4167)) and (layer4_outputs(890)));
    layer5_outputs(3792) <= not((layer4_outputs(3573)) and (layer4_outputs(2655)));
    layer5_outputs(3793) <= '1';
    layer5_outputs(3794) <= (layer4_outputs(1432)) and not (layer4_outputs(680));
    layer5_outputs(3795) <= (layer4_outputs(2121)) and not (layer4_outputs(2191));
    layer5_outputs(3796) <= layer4_outputs(3608);
    layer5_outputs(3797) <= (layer4_outputs(809)) and (layer4_outputs(1853));
    layer5_outputs(3798) <= layer4_outputs(4193);
    layer5_outputs(3799) <= not(layer4_outputs(1206));
    layer5_outputs(3800) <= not(layer4_outputs(778)) or (layer4_outputs(1339));
    layer5_outputs(3801) <= not(layer4_outputs(2691)) or (layer4_outputs(931));
    layer5_outputs(3802) <= (layer4_outputs(1377)) and not (layer4_outputs(4678));
    layer5_outputs(3803) <= layer4_outputs(3102);
    layer5_outputs(3804) <= not((layer4_outputs(1098)) or (layer4_outputs(2495)));
    layer5_outputs(3805) <= layer4_outputs(2107);
    layer5_outputs(3806) <= layer4_outputs(3530);
    layer5_outputs(3807) <= layer4_outputs(4419);
    layer5_outputs(3808) <= not(layer4_outputs(2939)) or (layer4_outputs(2736));
    layer5_outputs(3809) <= not((layer4_outputs(384)) xor (layer4_outputs(1675)));
    layer5_outputs(3810) <= (layer4_outputs(1150)) and not (layer4_outputs(2590));
    layer5_outputs(3811) <= not((layer4_outputs(68)) xor (layer4_outputs(717)));
    layer5_outputs(3812) <= layer4_outputs(4770);
    layer5_outputs(3813) <= (layer4_outputs(3547)) and (layer4_outputs(846));
    layer5_outputs(3814) <= layer4_outputs(64);
    layer5_outputs(3815) <= not((layer4_outputs(495)) and (layer4_outputs(278)));
    layer5_outputs(3816) <= '0';
    layer5_outputs(3817) <= layer4_outputs(1946);
    layer5_outputs(3818) <= (layer4_outputs(4934)) and not (layer4_outputs(2805));
    layer5_outputs(3819) <= not(layer4_outputs(2814)) or (layer4_outputs(4121));
    layer5_outputs(3820) <= not(layer4_outputs(3233));
    layer5_outputs(3821) <= layer4_outputs(1411);
    layer5_outputs(3822) <= not(layer4_outputs(2944)) or (layer4_outputs(3337));
    layer5_outputs(3823) <= (layer4_outputs(127)) xor (layer4_outputs(4032));
    layer5_outputs(3824) <= (layer4_outputs(3155)) or (layer4_outputs(2741));
    layer5_outputs(3825) <= layer4_outputs(3112);
    layer5_outputs(3826) <= not(layer4_outputs(4349)) or (layer4_outputs(2183));
    layer5_outputs(3827) <= layer4_outputs(607);
    layer5_outputs(3828) <= '0';
    layer5_outputs(3829) <= layer4_outputs(2432);
    layer5_outputs(3830) <= (layer4_outputs(1928)) and not (layer4_outputs(2371));
    layer5_outputs(3831) <= not(layer4_outputs(2480)) or (layer4_outputs(1717));
    layer5_outputs(3832) <= not(layer4_outputs(3213));
    layer5_outputs(3833) <= layer4_outputs(1110);
    layer5_outputs(3834) <= not((layer4_outputs(4017)) and (layer4_outputs(2383)));
    layer5_outputs(3835) <= not(layer4_outputs(1971));
    layer5_outputs(3836) <= '1';
    layer5_outputs(3837) <= not(layer4_outputs(3275)) or (layer4_outputs(4508));
    layer5_outputs(3838) <= not((layer4_outputs(1802)) xor (layer4_outputs(4450)));
    layer5_outputs(3839) <= layer4_outputs(909);
    layer5_outputs(3840) <= not((layer4_outputs(3094)) or (layer4_outputs(1245)));
    layer5_outputs(3841) <= (layer4_outputs(742)) xor (layer4_outputs(1469));
    layer5_outputs(3842) <= layer4_outputs(3009);
    layer5_outputs(3843) <= not(layer4_outputs(3895)) or (layer4_outputs(1168));
    layer5_outputs(3844) <= layer4_outputs(4383);
    layer5_outputs(3845) <= not(layer4_outputs(2730)) or (layer4_outputs(4028));
    layer5_outputs(3846) <= not((layer4_outputs(3576)) and (layer4_outputs(4442)));
    layer5_outputs(3847) <= (layer4_outputs(2971)) or (layer4_outputs(3376));
    layer5_outputs(3848) <= not(layer4_outputs(3620));
    layer5_outputs(3849) <= not(layer4_outputs(907));
    layer5_outputs(3850) <= layer4_outputs(1329);
    layer5_outputs(3851) <= (layer4_outputs(1214)) or (layer4_outputs(3645));
    layer5_outputs(3852) <= not(layer4_outputs(2467));
    layer5_outputs(3853) <= (layer4_outputs(3442)) and (layer4_outputs(1544));
    layer5_outputs(3854) <= not((layer4_outputs(2605)) and (layer4_outputs(1187)));
    layer5_outputs(3855) <= not(layer4_outputs(802));
    layer5_outputs(3856) <= (layer4_outputs(3340)) or (layer4_outputs(1683));
    layer5_outputs(3857) <= not(layer4_outputs(3349));
    layer5_outputs(3858) <= not((layer4_outputs(1046)) xor (layer4_outputs(714)));
    layer5_outputs(3859) <= not((layer4_outputs(1855)) and (layer4_outputs(35)));
    layer5_outputs(3860) <= (layer4_outputs(2210)) or (layer4_outputs(1021));
    layer5_outputs(3861) <= layer4_outputs(3400);
    layer5_outputs(3862) <= not((layer4_outputs(1460)) and (layer4_outputs(4922)));
    layer5_outputs(3863) <= (layer4_outputs(3159)) and (layer4_outputs(4925));
    layer5_outputs(3864) <= not(layer4_outputs(3501));
    layer5_outputs(3865) <= (layer4_outputs(1276)) and (layer4_outputs(1073));
    layer5_outputs(3866) <= not(layer4_outputs(1099));
    layer5_outputs(3867) <= (layer4_outputs(1007)) xor (layer4_outputs(4752));
    layer5_outputs(3868) <= not(layer4_outputs(14));
    layer5_outputs(3869) <= not((layer4_outputs(3342)) xor (layer4_outputs(1709)));
    layer5_outputs(3870) <= (layer4_outputs(3615)) and (layer4_outputs(2695));
    layer5_outputs(3871) <= (layer4_outputs(4120)) xor (layer4_outputs(48));
    layer5_outputs(3872) <= not(layer4_outputs(4497)) or (layer4_outputs(4814));
    layer5_outputs(3873) <= (layer4_outputs(1317)) and not (layer4_outputs(305));
    layer5_outputs(3874) <= layer4_outputs(3571);
    layer5_outputs(3875) <= layer4_outputs(1856);
    layer5_outputs(3876) <= not(layer4_outputs(3548));
    layer5_outputs(3877) <= not(layer4_outputs(4818)) or (layer4_outputs(4656));
    layer5_outputs(3878) <= not(layer4_outputs(2450));
    layer5_outputs(3879) <= not((layer4_outputs(4110)) and (layer4_outputs(3152)));
    layer5_outputs(3880) <= not(layer4_outputs(4024));
    layer5_outputs(3881) <= not((layer4_outputs(2209)) or (layer4_outputs(1051)));
    layer5_outputs(3882) <= (layer4_outputs(3689)) and not (layer4_outputs(4369));
    layer5_outputs(3883) <= not(layer4_outputs(3717));
    layer5_outputs(3884) <= (layer4_outputs(2117)) and not (layer4_outputs(3233));
    layer5_outputs(3885) <= not(layer4_outputs(319));
    layer5_outputs(3886) <= (layer4_outputs(959)) and (layer4_outputs(2355));
    layer5_outputs(3887) <= not(layer4_outputs(4566)) or (layer4_outputs(4920));
    layer5_outputs(3888) <= layer4_outputs(3474);
    layer5_outputs(3889) <= not(layer4_outputs(2770));
    layer5_outputs(3890) <= layer4_outputs(5067);
    layer5_outputs(3891) <= not((layer4_outputs(2643)) or (layer4_outputs(730)));
    layer5_outputs(3892) <= layer4_outputs(4063);
    layer5_outputs(3893) <= (layer4_outputs(1653)) and (layer4_outputs(2647));
    layer5_outputs(3894) <= not(layer4_outputs(1293)) or (layer4_outputs(3638));
    layer5_outputs(3895) <= (layer4_outputs(2919)) and not (layer4_outputs(32));
    layer5_outputs(3896) <= (layer4_outputs(666)) or (layer4_outputs(862));
    layer5_outputs(3897) <= '0';
    layer5_outputs(3898) <= (layer4_outputs(3220)) and (layer4_outputs(1827));
    layer5_outputs(3899) <= not(layer4_outputs(1170)) or (layer4_outputs(1341));
    layer5_outputs(3900) <= layer4_outputs(4003);
    layer5_outputs(3901) <= (layer4_outputs(2304)) and (layer4_outputs(4945));
    layer5_outputs(3902) <= not((layer4_outputs(3734)) xor (layer4_outputs(4064)));
    layer5_outputs(3903) <= not(layer4_outputs(1715));
    layer5_outputs(3904) <= not(layer4_outputs(1374)) or (layer4_outputs(3095));
    layer5_outputs(3905) <= not(layer4_outputs(4314));
    layer5_outputs(3906) <= not((layer4_outputs(768)) xor (layer4_outputs(1428)));
    layer5_outputs(3907) <= layer4_outputs(1016);
    layer5_outputs(3908) <= not(layer4_outputs(2407));
    layer5_outputs(3909) <= not((layer4_outputs(252)) or (layer4_outputs(1201)));
    layer5_outputs(3910) <= not(layer4_outputs(1576));
    layer5_outputs(3911) <= not(layer4_outputs(4098));
    layer5_outputs(3912) <= layer4_outputs(1037);
    layer5_outputs(3913) <= not(layer4_outputs(1497));
    layer5_outputs(3914) <= not(layer4_outputs(1341)) or (layer4_outputs(558));
    layer5_outputs(3915) <= not(layer4_outputs(924));
    layer5_outputs(3916) <= (layer4_outputs(1874)) or (layer4_outputs(3561));
    layer5_outputs(3917) <= (layer4_outputs(2944)) and not (layer4_outputs(830));
    layer5_outputs(3918) <= '1';
    layer5_outputs(3919) <= (layer4_outputs(3593)) and not (layer4_outputs(2602));
    layer5_outputs(3920) <= layer4_outputs(3295);
    layer5_outputs(3921) <= '1';
    layer5_outputs(3922) <= not((layer4_outputs(2029)) and (layer4_outputs(4392)));
    layer5_outputs(3923) <= '1';
    layer5_outputs(3924) <= (layer4_outputs(550)) and (layer4_outputs(1174));
    layer5_outputs(3925) <= not(layer4_outputs(4516));
    layer5_outputs(3926) <= not(layer4_outputs(5081));
    layer5_outputs(3927) <= not((layer4_outputs(2485)) xor (layer4_outputs(264)));
    layer5_outputs(3928) <= layer4_outputs(3480);
    layer5_outputs(3929) <= (layer4_outputs(1399)) and not (layer4_outputs(4330));
    layer5_outputs(3930) <= layer4_outputs(3683);
    layer5_outputs(3931) <= not(layer4_outputs(1606));
    layer5_outputs(3932) <= not(layer4_outputs(3843));
    layer5_outputs(3933) <= '1';
    layer5_outputs(3934) <= not(layer4_outputs(3061));
    layer5_outputs(3935) <= (layer4_outputs(623)) and not (layer4_outputs(3779));
    layer5_outputs(3936) <= layer4_outputs(4657);
    layer5_outputs(3937) <= not(layer4_outputs(4504)) or (layer4_outputs(4414));
    layer5_outputs(3938) <= (layer4_outputs(2980)) and (layer4_outputs(2637));
    layer5_outputs(3939) <= (layer4_outputs(1922)) and (layer4_outputs(3650));
    layer5_outputs(3940) <= not((layer4_outputs(2512)) and (layer4_outputs(1474)));
    layer5_outputs(3941) <= not(layer4_outputs(2405)) or (layer4_outputs(303));
    layer5_outputs(3942) <= not((layer4_outputs(964)) or (layer4_outputs(2864)));
    layer5_outputs(3943) <= not((layer4_outputs(4486)) and (layer4_outputs(1321)));
    layer5_outputs(3944) <= not(layer4_outputs(2259)) or (layer4_outputs(2469));
    layer5_outputs(3945) <= not((layer4_outputs(2834)) and (layer4_outputs(1754)));
    layer5_outputs(3946) <= not((layer4_outputs(2243)) and (layer4_outputs(2104)));
    layer5_outputs(3947) <= not(layer4_outputs(2284));
    layer5_outputs(3948) <= not((layer4_outputs(4837)) xor (layer4_outputs(1094)));
    layer5_outputs(3949) <= (layer4_outputs(1813)) and (layer4_outputs(1846));
    layer5_outputs(3950) <= not(layer4_outputs(678));
    layer5_outputs(3951) <= '1';
    layer5_outputs(3952) <= layer4_outputs(4764);
    layer5_outputs(3953) <= not((layer4_outputs(3695)) and (layer4_outputs(3488)));
    layer5_outputs(3954) <= not((layer4_outputs(3217)) or (layer4_outputs(1136)));
    layer5_outputs(3955) <= '1';
    layer5_outputs(3956) <= layer4_outputs(2352);
    layer5_outputs(3957) <= layer4_outputs(185);
    layer5_outputs(3958) <= '1';
    layer5_outputs(3959) <= layer4_outputs(3981);
    layer5_outputs(3960) <= '0';
    layer5_outputs(3961) <= not((layer4_outputs(265)) and (layer4_outputs(5110)));
    layer5_outputs(3962) <= not(layer4_outputs(1996)) or (layer4_outputs(738));
    layer5_outputs(3963) <= (layer4_outputs(4804)) and not (layer4_outputs(945));
    layer5_outputs(3964) <= not(layer4_outputs(777)) or (layer4_outputs(2076));
    layer5_outputs(3965) <= layer4_outputs(200);
    layer5_outputs(3966) <= not(layer4_outputs(112));
    layer5_outputs(3967) <= layer4_outputs(4510);
    layer5_outputs(3968) <= not(layer4_outputs(5046));
    layer5_outputs(3969) <= layer4_outputs(627);
    layer5_outputs(3970) <= (layer4_outputs(3530)) xor (layer4_outputs(1744));
    layer5_outputs(3971) <= not(layer4_outputs(2298));
    layer5_outputs(3972) <= layer4_outputs(4398);
    layer5_outputs(3973) <= (layer4_outputs(3711)) or (layer4_outputs(4456));
    layer5_outputs(3974) <= layer4_outputs(3264);
    layer5_outputs(3975) <= (layer4_outputs(4760)) and not (layer4_outputs(3096));
    layer5_outputs(3976) <= not(layer4_outputs(1768)) or (layer4_outputs(4269));
    layer5_outputs(3977) <= (layer4_outputs(3913)) xor (layer4_outputs(2595));
    layer5_outputs(3978) <= layer4_outputs(4083);
    layer5_outputs(3979) <= (layer4_outputs(209)) or (layer4_outputs(4576));
    layer5_outputs(3980) <= not(layer4_outputs(4765));
    layer5_outputs(3981) <= (layer4_outputs(3173)) and not (layer4_outputs(1972));
    layer5_outputs(3982) <= '0';
    layer5_outputs(3983) <= not(layer4_outputs(3587));
    layer5_outputs(3984) <= '0';
    layer5_outputs(3985) <= not(layer4_outputs(1159));
    layer5_outputs(3986) <= (layer4_outputs(2758)) or (layer4_outputs(2262));
    layer5_outputs(3987) <= layer4_outputs(3045);
    layer5_outputs(3988) <= not(layer4_outputs(3885));
    layer5_outputs(3989) <= not((layer4_outputs(4615)) or (layer4_outputs(2782)));
    layer5_outputs(3990) <= not(layer4_outputs(4302)) or (layer4_outputs(1921));
    layer5_outputs(3991) <= layer4_outputs(2000);
    layer5_outputs(3992) <= '1';
    layer5_outputs(3993) <= layer4_outputs(3750);
    layer5_outputs(3994) <= layer4_outputs(2226);
    layer5_outputs(3995) <= (layer4_outputs(3180)) and not (layer4_outputs(3599));
    layer5_outputs(3996) <= not((layer4_outputs(148)) or (layer4_outputs(4384)));
    layer5_outputs(3997) <= (layer4_outputs(301)) and not (layer4_outputs(2385));
    layer5_outputs(3998) <= (layer4_outputs(798)) and not (layer4_outputs(947));
    layer5_outputs(3999) <= not(layer4_outputs(4703));
    layer5_outputs(4000) <= layer4_outputs(3141);
    layer5_outputs(4001) <= not((layer4_outputs(2030)) or (layer4_outputs(3734)));
    layer5_outputs(4002) <= not((layer4_outputs(4774)) and (layer4_outputs(138)));
    layer5_outputs(4003) <= layer4_outputs(3547);
    layer5_outputs(4004) <= (layer4_outputs(2869)) or (layer4_outputs(371));
    layer5_outputs(4005) <= (layer4_outputs(612)) and not (layer4_outputs(716));
    layer5_outputs(4006) <= layer4_outputs(2400);
    layer5_outputs(4007) <= (layer4_outputs(2476)) and (layer4_outputs(1309));
    layer5_outputs(4008) <= layer4_outputs(4014);
    layer5_outputs(4009) <= (layer4_outputs(1223)) and (layer4_outputs(2005));
    layer5_outputs(4010) <= not(layer4_outputs(2829));
    layer5_outputs(4011) <= layer4_outputs(249);
    layer5_outputs(4012) <= '1';
    layer5_outputs(4013) <= '1';
    layer5_outputs(4014) <= layer4_outputs(2248);
    layer5_outputs(4015) <= (layer4_outputs(3553)) and not (layer4_outputs(288));
    layer5_outputs(4016) <= (layer4_outputs(3428)) and (layer4_outputs(1785));
    layer5_outputs(4017) <= not((layer4_outputs(767)) or (layer4_outputs(438)));
    layer5_outputs(4018) <= '1';
    layer5_outputs(4019) <= (layer4_outputs(966)) and not (layer4_outputs(1386));
    layer5_outputs(4020) <= '0';
    layer5_outputs(4021) <= not((layer4_outputs(1090)) or (layer4_outputs(4269)));
    layer5_outputs(4022) <= (layer4_outputs(4417)) xor (layer4_outputs(4928));
    layer5_outputs(4023) <= not((layer4_outputs(1476)) or (layer4_outputs(3099)));
    layer5_outputs(4024) <= not(layer4_outputs(3789));
    layer5_outputs(4025) <= layer4_outputs(4870);
    layer5_outputs(4026) <= (layer4_outputs(5075)) and (layer4_outputs(44));
    layer5_outputs(4027) <= not(layer4_outputs(3563));
    layer5_outputs(4028) <= not(layer4_outputs(1662));
    layer5_outputs(4029) <= not((layer4_outputs(2165)) xor (layer4_outputs(1849)));
    layer5_outputs(4030) <= (layer4_outputs(4577)) or (layer4_outputs(685));
    layer5_outputs(4031) <= not((layer4_outputs(3068)) or (layer4_outputs(4427)));
    layer5_outputs(4032) <= not(layer4_outputs(4957));
    layer5_outputs(4033) <= not(layer4_outputs(3091));
    layer5_outputs(4034) <= not(layer4_outputs(243));
    layer5_outputs(4035) <= not((layer4_outputs(1933)) and (layer4_outputs(1266)));
    layer5_outputs(4036) <= '0';
    layer5_outputs(4037) <= (layer4_outputs(437)) and (layer4_outputs(4890));
    layer5_outputs(4038) <= not((layer4_outputs(3927)) or (layer4_outputs(4730)));
    layer5_outputs(4039) <= layer4_outputs(5021);
    layer5_outputs(4040) <= (layer4_outputs(2321)) and not (layer4_outputs(2312));
    layer5_outputs(4041) <= '0';
    layer5_outputs(4042) <= (layer4_outputs(4503)) and not (layer4_outputs(713));
    layer5_outputs(4043) <= layer4_outputs(2277);
    layer5_outputs(4044) <= (layer4_outputs(4929)) and (layer4_outputs(2597));
    layer5_outputs(4045) <= layer4_outputs(489);
    layer5_outputs(4046) <= not(layer4_outputs(2506)) or (layer4_outputs(3207));
    layer5_outputs(4047) <= (layer4_outputs(1110)) and (layer4_outputs(4126));
    layer5_outputs(4048) <= layer4_outputs(5090);
    layer5_outputs(4049) <= (layer4_outputs(2806)) and (layer4_outputs(3149));
    layer5_outputs(4050) <= (layer4_outputs(2545)) and not (layer4_outputs(4196));
    layer5_outputs(4051) <= layer4_outputs(4469);
    layer5_outputs(4052) <= not(layer4_outputs(4441));
    layer5_outputs(4053) <= not(layer4_outputs(4468));
    layer5_outputs(4054) <= (layer4_outputs(2217)) and not (layer4_outputs(1101));
    layer5_outputs(4055) <= not(layer4_outputs(4213));
    layer5_outputs(4056) <= not(layer4_outputs(5002)) or (layer4_outputs(177));
    layer5_outputs(4057) <= layer4_outputs(2373);
    layer5_outputs(4058) <= not((layer4_outputs(4831)) and (layer4_outputs(3330)));
    layer5_outputs(4059) <= layer4_outputs(3534);
    layer5_outputs(4060) <= not(layer4_outputs(1676));
    layer5_outputs(4061) <= not(layer4_outputs(2102));
    layer5_outputs(4062) <= not((layer4_outputs(65)) or (layer4_outputs(4509)));
    layer5_outputs(4063) <= not(layer4_outputs(443));
    layer5_outputs(4064) <= (layer4_outputs(556)) and (layer4_outputs(2480));
    layer5_outputs(4065) <= '0';
    layer5_outputs(4066) <= not(layer4_outputs(3961));
    layer5_outputs(4067) <= (layer4_outputs(4188)) or (layer4_outputs(2199));
    layer5_outputs(4068) <= (layer4_outputs(630)) and not (layer4_outputs(333));
    layer5_outputs(4069) <= (layer4_outputs(5011)) and not (layer4_outputs(2436));
    layer5_outputs(4070) <= (layer4_outputs(3545)) and not (layer4_outputs(1035));
    layer5_outputs(4071) <= (layer4_outputs(1562)) and not (layer4_outputs(933));
    layer5_outputs(4072) <= not(layer4_outputs(3968)) or (layer4_outputs(1499));
    layer5_outputs(4073) <= not(layer4_outputs(4189));
    layer5_outputs(4074) <= not(layer4_outputs(4504)) or (layer4_outputs(3999));
    layer5_outputs(4075) <= not(layer4_outputs(2020));
    layer5_outputs(4076) <= not(layer4_outputs(4839));
    layer5_outputs(4077) <= not(layer4_outputs(2427)) or (layer4_outputs(2072));
    layer5_outputs(4078) <= (layer4_outputs(203)) or (layer4_outputs(496));
    layer5_outputs(4079) <= not((layer4_outputs(2831)) or (layer4_outputs(2614)));
    layer5_outputs(4080) <= not(layer4_outputs(4642));
    layer5_outputs(4081) <= not(layer4_outputs(3973));
    layer5_outputs(4082) <= layer4_outputs(4259);
    layer5_outputs(4083) <= not(layer4_outputs(217));
    layer5_outputs(4084) <= layer4_outputs(1948);
    layer5_outputs(4085) <= (layer4_outputs(1850)) and not (layer4_outputs(4263));
    layer5_outputs(4086) <= (layer4_outputs(1454)) and not (layer4_outputs(699));
    layer5_outputs(4087) <= not(layer4_outputs(3388));
    layer5_outputs(4088) <= layer4_outputs(1550);
    layer5_outputs(4089) <= not((layer4_outputs(1454)) and (layer4_outputs(2793)));
    layer5_outputs(4090) <= '0';
    layer5_outputs(4091) <= layer4_outputs(366);
    layer5_outputs(4092) <= layer4_outputs(3602);
    layer5_outputs(4093) <= '1';
    layer5_outputs(4094) <= (layer4_outputs(600)) and not (layer4_outputs(1372));
    layer5_outputs(4095) <= not(layer4_outputs(84));
    layer5_outputs(4096) <= not(layer4_outputs(632)) or (layer4_outputs(420));
    layer5_outputs(4097) <= not((layer4_outputs(2128)) or (layer4_outputs(720)));
    layer5_outputs(4098) <= (layer4_outputs(4432)) or (layer4_outputs(1492));
    layer5_outputs(4099) <= layer4_outputs(4396);
    layer5_outputs(4100) <= layer4_outputs(2137);
    layer5_outputs(4101) <= layer4_outputs(822);
    layer5_outputs(4102) <= (layer4_outputs(4883)) and not (layer4_outputs(3811));
    layer5_outputs(4103) <= not((layer4_outputs(2791)) and (layer4_outputs(3325)));
    layer5_outputs(4104) <= layer4_outputs(3049);
    layer5_outputs(4105) <= not(layer4_outputs(1730));
    layer5_outputs(4106) <= not((layer4_outputs(1012)) and (layer4_outputs(1891)));
    layer5_outputs(4107) <= layer4_outputs(4498);
    layer5_outputs(4108) <= not(layer4_outputs(699));
    layer5_outputs(4109) <= not(layer4_outputs(4408));
    layer5_outputs(4110) <= (layer4_outputs(1330)) and not (layer4_outputs(2281));
    layer5_outputs(4111) <= not((layer4_outputs(4994)) or (layer4_outputs(3603)));
    layer5_outputs(4112) <= not((layer4_outputs(1131)) and (layer4_outputs(1692)));
    layer5_outputs(4113) <= not((layer4_outputs(2724)) xor (layer4_outputs(4720)));
    layer5_outputs(4114) <= layer4_outputs(1279);
    layer5_outputs(4115) <= '1';
    layer5_outputs(4116) <= not(layer4_outputs(616));
    layer5_outputs(4117) <= layer4_outputs(366);
    layer5_outputs(4118) <= (layer4_outputs(4339)) and not (layer4_outputs(2807));
    layer5_outputs(4119) <= not((layer4_outputs(4220)) and (layer4_outputs(4863)));
    layer5_outputs(4120) <= not((layer4_outputs(3095)) and (layer4_outputs(1659)));
    layer5_outputs(4121) <= not((layer4_outputs(2748)) and (layer4_outputs(3401)));
    layer5_outputs(4122) <= not((layer4_outputs(1469)) and (layer4_outputs(2239)));
    layer5_outputs(4123) <= not(layer4_outputs(1502));
    layer5_outputs(4124) <= not(layer4_outputs(721));
    layer5_outputs(4125) <= not(layer4_outputs(2609));
    layer5_outputs(4126) <= (layer4_outputs(56)) and (layer4_outputs(4136));
    layer5_outputs(4127) <= not(layer4_outputs(3445)) or (layer4_outputs(248));
    layer5_outputs(4128) <= (layer4_outputs(1657)) and (layer4_outputs(3579));
    layer5_outputs(4129) <= '1';
    layer5_outputs(4130) <= layer4_outputs(1776);
    layer5_outputs(4131) <= (layer4_outputs(2232)) or (layer4_outputs(354));
    layer5_outputs(4132) <= not(layer4_outputs(1446));
    layer5_outputs(4133) <= layer4_outputs(3076);
    layer5_outputs(4134) <= layer4_outputs(1516);
    layer5_outputs(4135) <= not((layer4_outputs(4236)) and (layer4_outputs(3782)));
    layer5_outputs(4136) <= (layer4_outputs(3320)) and not (layer4_outputs(897));
    layer5_outputs(4137) <= not(layer4_outputs(86));
    layer5_outputs(4138) <= not(layer4_outputs(2814)) or (layer4_outputs(3353));
    layer5_outputs(4139) <= (layer4_outputs(633)) or (layer4_outputs(4747));
    layer5_outputs(4140) <= layer4_outputs(1044);
    layer5_outputs(4141) <= not((layer4_outputs(3940)) and (layer4_outputs(2712)));
    layer5_outputs(4142) <= (layer4_outputs(170)) and not (layer4_outputs(1882));
    layer5_outputs(4143) <= not(layer4_outputs(4499));
    layer5_outputs(4144) <= not(layer4_outputs(3612)) or (layer4_outputs(226));
    layer5_outputs(4145) <= (layer4_outputs(4326)) and not (layer4_outputs(2797));
    layer5_outputs(4146) <= '1';
    layer5_outputs(4147) <= (layer4_outputs(61)) and not (layer4_outputs(973));
    layer5_outputs(4148) <= (layer4_outputs(4520)) and not (layer4_outputs(1918));
    layer5_outputs(4149) <= not(layer4_outputs(347));
    layer5_outputs(4150) <= (layer4_outputs(2387)) and (layer4_outputs(1282));
    layer5_outputs(4151) <= not(layer4_outputs(4598));
    layer5_outputs(4152) <= (layer4_outputs(4999)) and not (layer4_outputs(1573));
    layer5_outputs(4153) <= (layer4_outputs(3183)) or (layer4_outputs(2077));
    layer5_outputs(4154) <= not(layer4_outputs(1001)) or (layer4_outputs(4148));
    layer5_outputs(4155) <= not(layer4_outputs(2269));
    layer5_outputs(4156) <= (layer4_outputs(2755)) xor (layer4_outputs(1901));
    layer5_outputs(4157) <= (layer4_outputs(2845)) or (layer4_outputs(1493));
    layer5_outputs(4158) <= (layer4_outputs(4604)) xor (layer4_outputs(90));
    layer5_outputs(4159) <= not((layer4_outputs(2602)) or (layer4_outputs(1408)));
    layer5_outputs(4160) <= not(layer4_outputs(3122));
    layer5_outputs(4161) <= '0';
    layer5_outputs(4162) <= layer4_outputs(3936);
    layer5_outputs(4163) <= not(layer4_outputs(4643));
    layer5_outputs(4164) <= not(layer4_outputs(1575));
    layer5_outputs(4165) <= (layer4_outputs(4860)) and (layer4_outputs(1905));
    layer5_outputs(4166) <= (layer4_outputs(4711)) and (layer4_outputs(20));
    layer5_outputs(4167) <= not(layer4_outputs(686));
    layer5_outputs(4168) <= not(layer4_outputs(3892)) or (layer4_outputs(1911));
    layer5_outputs(4169) <= (layer4_outputs(4274)) and not (layer4_outputs(4947));
    layer5_outputs(4170) <= not((layer4_outputs(1510)) and (layer4_outputs(589)));
    layer5_outputs(4171) <= (layer4_outputs(3873)) or (layer4_outputs(2349));
    layer5_outputs(4172) <= not(layer4_outputs(4499)) or (layer4_outputs(3288));
    layer5_outputs(4173) <= layer4_outputs(3238);
    layer5_outputs(4174) <= not(layer4_outputs(4188));
    layer5_outputs(4175) <= not(layer4_outputs(4579));
    layer5_outputs(4176) <= (layer4_outputs(1789)) and not (layer4_outputs(3008));
    layer5_outputs(4177) <= not(layer4_outputs(2114));
    layer5_outputs(4178) <= (layer4_outputs(4391)) and not (layer4_outputs(4575));
    layer5_outputs(4179) <= (layer4_outputs(459)) and not (layer4_outputs(3086));
    layer5_outputs(4180) <= '1';
    layer5_outputs(4181) <= layer4_outputs(4052);
    layer5_outputs(4182) <= (layer4_outputs(2042)) and (layer4_outputs(345));
    layer5_outputs(4183) <= (layer4_outputs(2796)) and not (layer4_outputs(4502));
    layer5_outputs(4184) <= layer4_outputs(2876);
    layer5_outputs(4185) <= (layer4_outputs(2325)) and not (layer4_outputs(4356));
    layer5_outputs(4186) <= not((layer4_outputs(391)) xor (layer4_outputs(3556)));
    layer5_outputs(4187) <= '1';
    layer5_outputs(4188) <= (layer4_outputs(3294)) and not (layer4_outputs(2843));
    layer5_outputs(4189) <= layer4_outputs(2582);
    layer5_outputs(4190) <= layer4_outputs(5006);
    layer5_outputs(4191) <= not(layer4_outputs(2559)) or (layer4_outputs(2308));
    layer5_outputs(4192) <= layer4_outputs(1215);
    layer5_outputs(4193) <= not(layer4_outputs(1863));
    layer5_outputs(4194) <= not(layer4_outputs(2462));
    layer5_outputs(4195) <= not(layer4_outputs(2312));
    layer5_outputs(4196) <= layer4_outputs(3236);
    layer5_outputs(4197) <= (layer4_outputs(2474)) xor (layer4_outputs(2299));
    layer5_outputs(4198) <= not((layer4_outputs(841)) or (layer4_outputs(2049)));
    layer5_outputs(4199) <= layer4_outputs(4891);
    layer5_outputs(4200) <= (layer4_outputs(2671)) or (layer4_outputs(1625));
    layer5_outputs(4201) <= '1';
    layer5_outputs(4202) <= (layer4_outputs(1715)) or (layer4_outputs(735));
    layer5_outputs(4203) <= not((layer4_outputs(4666)) or (layer4_outputs(4071)));
    layer5_outputs(4204) <= (layer4_outputs(116)) and (layer4_outputs(1508));
    layer5_outputs(4205) <= (layer4_outputs(4751)) and (layer4_outputs(11));
    layer5_outputs(4206) <= (layer4_outputs(1560)) and not (layer4_outputs(1361));
    layer5_outputs(4207) <= layer4_outputs(4588);
    layer5_outputs(4208) <= (layer4_outputs(1817)) and not (layer4_outputs(3378));
    layer5_outputs(4209) <= (layer4_outputs(4072)) and not (layer4_outputs(3754));
    layer5_outputs(4210) <= not(layer4_outputs(4814)) or (layer4_outputs(1338));
    layer5_outputs(4211) <= not((layer4_outputs(4537)) xor (layer4_outputs(5074)));
    layer5_outputs(4212) <= not(layer4_outputs(3317));
    layer5_outputs(4213) <= (layer4_outputs(1664)) or (layer4_outputs(3955));
    layer5_outputs(4214) <= not(layer4_outputs(57));
    layer5_outputs(4215) <= (layer4_outputs(4431)) xor (layer4_outputs(2599));
    layer5_outputs(4216) <= (layer4_outputs(3275)) or (layer4_outputs(678));
    layer5_outputs(4217) <= not(layer4_outputs(2632));
    layer5_outputs(4218) <= not((layer4_outputs(926)) xor (layer4_outputs(955)));
    layer5_outputs(4219) <= layer4_outputs(2123);
    layer5_outputs(4220) <= not((layer4_outputs(451)) and (layer4_outputs(4318)));
    layer5_outputs(4221) <= not(layer4_outputs(1330));
    layer5_outputs(4222) <= layer4_outputs(1936);
    layer5_outputs(4223) <= not((layer4_outputs(2086)) and (layer4_outputs(3625)));
    layer5_outputs(4224) <= not(layer4_outputs(647));
    layer5_outputs(4225) <= '0';
    layer5_outputs(4226) <= (layer4_outputs(3795)) and not (layer4_outputs(2522));
    layer5_outputs(4227) <= not(layer4_outputs(4832));
    layer5_outputs(4228) <= not(layer4_outputs(3862));
    layer5_outputs(4229) <= not((layer4_outputs(4137)) and (layer4_outputs(4866)));
    layer5_outputs(4230) <= not(layer4_outputs(4954));
    layer5_outputs(4231) <= layer4_outputs(5104);
    layer5_outputs(4232) <= layer4_outputs(578);
    layer5_outputs(4233) <= layer4_outputs(1509);
    layer5_outputs(4234) <= (layer4_outputs(3248)) and (layer4_outputs(3308));
    layer5_outputs(4235) <= (layer4_outputs(4630)) and not (layer4_outputs(1635));
    layer5_outputs(4236) <= not(layer4_outputs(4105));
    layer5_outputs(4237) <= not(layer4_outputs(1707));
    layer5_outputs(4238) <= layer4_outputs(56);
    layer5_outputs(4239) <= not(layer4_outputs(2094)) or (layer4_outputs(4506));
    layer5_outputs(4240) <= not((layer4_outputs(953)) and (layer4_outputs(3359)));
    layer5_outputs(4241) <= layer4_outputs(3654);
    layer5_outputs(4242) <= layer4_outputs(1729);
    layer5_outputs(4243) <= layer4_outputs(337);
    layer5_outputs(4244) <= layer4_outputs(5009);
    layer5_outputs(4245) <= not(layer4_outputs(1331));
    layer5_outputs(4246) <= not(layer4_outputs(3450));
    layer5_outputs(4247) <= not(layer4_outputs(4185));
    layer5_outputs(4248) <= layer4_outputs(1691);
    layer5_outputs(4249) <= layer4_outputs(4109);
    layer5_outputs(4250) <= layer4_outputs(951);
    layer5_outputs(4251) <= not(layer4_outputs(4003));
    layer5_outputs(4252) <= not(layer4_outputs(4222));
    layer5_outputs(4253) <= (layer4_outputs(3778)) and not (layer4_outputs(2194));
    layer5_outputs(4254) <= not((layer4_outputs(4214)) and (layer4_outputs(198)));
    layer5_outputs(4255) <= not((layer4_outputs(4946)) or (layer4_outputs(1421)));
    layer5_outputs(4256) <= not((layer4_outputs(823)) xor (layer4_outputs(1182)));
    layer5_outputs(4257) <= (layer4_outputs(284)) and not (layer4_outputs(2569));
    layer5_outputs(4258) <= not((layer4_outputs(2122)) or (layer4_outputs(4040)));
    layer5_outputs(4259) <= not(layer4_outputs(274));
    layer5_outputs(4260) <= (layer4_outputs(4258)) and not (layer4_outputs(3903));
    layer5_outputs(4261) <= not(layer4_outputs(4847));
    layer5_outputs(4262) <= (layer4_outputs(2289)) or (layer4_outputs(1933));
    layer5_outputs(4263) <= (layer4_outputs(894)) xor (layer4_outputs(4465));
    layer5_outputs(4264) <= not((layer4_outputs(4865)) and (layer4_outputs(1916)));
    layer5_outputs(4265) <= not((layer4_outputs(339)) xor (layer4_outputs(1348)));
    layer5_outputs(4266) <= (layer4_outputs(1399)) xor (layer4_outputs(400));
    layer5_outputs(4267) <= not(layer4_outputs(2464)) or (layer4_outputs(3666));
    layer5_outputs(4268) <= (layer4_outputs(1473)) and not (layer4_outputs(331));
    layer5_outputs(4269) <= (layer4_outputs(4546)) and (layer4_outputs(1133));
    layer5_outputs(4270) <= (layer4_outputs(3083)) and not (layer4_outputs(4224));
    layer5_outputs(4271) <= (layer4_outputs(2183)) and (layer4_outputs(4733));
    layer5_outputs(4272) <= not(layer4_outputs(1769)) or (layer4_outputs(1021));
    layer5_outputs(4273) <= not((layer4_outputs(4327)) and (layer4_outputs(2584)));
    layer5_outputs(4274) <= not((layer4_outputs(2759)) and (layer4_outputs(4744)));
    layer5_outputs(4275) <= not(layer4_outputs(3690)) or (layer4_outputs(470));
    layer5_outputs(4276) <= not(layer4_outputs(1167));
    layer5_outputs(4277) <= not(layer4_outputs(2862));
    layer5_outputs(4278) <= not(layer4_outputs(2785));
    layer5_outputs(4279) <= layer4_outputs(4745);
    layer5_outputs(4280) <= layer4_outputs(2874);
    layer5_outputs(4281) <= (layer4_outputs(335)) or (layer4_outputs(417));
    layer5_outputs(4282) <= not(layer4_outputs(5040)) or (layer4_outputs(3484));
    layer5_outputs(4283) <= not(layer4_outputs(2039));
    layer5_outputs(4284) <= not(layer4_outputs(3092));
    layer5_outputs(4285) <= not(layer4_outputs(3074));
    layer5_outputs(4286) <= layer4_outputs(79);
    layer5_outputs(4287) <= not(layer4_outputs(2041));
    layer5_outputs(4288) <= layer4_outputs(3040);
    layer5_outputs(4289) <= layer4_outputs(2245);
    layer5_outputs(4290) <= not((layer4_outputs(4883)) and (layer4_outputs(468)));
    layer5_outputs(4291) <= layer4_outputs(2953);
    layer5_outputs(4292) <= not(layer4_outputs(260)) or (layer4_outputs(270));
    layer5_outputs(4293) <= not(layer4_outputs(3267)) or (layer4_outputs(2139));
    layer5_outputs(4294) <= '0';
    layer5_outputs(4295) <= not(layer4_outputs(957)) or (layer4_outputs(3254));
    layer5_outputs(4296) <= not(layer4_outputs(880));
    layer5_outputs(4297) <= '1';
    layer5_outputs(4298) <= '1';
    layer5_outputs(4299) <= layer4_outputs(762);
    layer5_outputs(4300) <= (layer4_outputs(70)) or (layer4_outputs(234));
    layer5_outputs(4301) <= (layer4_outputs(4955)) xor (layer4_outputs(3686));
    layer5_outputs(4302) <= layer4_outputs(1655);
    layer5_outputs(4303) <= (layer4_outputs(2669)) and (layer4_outputs(4739));
    layer5_outputs(4304) <= (layer4_outputs(4307)) and (layer4_outputs(1773));
    layer5_outputs(4305) <= (layer4_outputs(5072)) and not (layer4_outputs(232));
    layer5_outputs(4306) <= layer4_outputs(2663);
    layer5_outputs(4307) <= '1';
    layer5_outputs(4308) <= not((layer4_outputs(3994)) and (layer4_outputs(754)));
    layer5_outputs(4309) <= not(layer4_outputs(3928));
    layer5_outputs(4310) <= layer4_outputs(4709);
    layer5_outputs(4311) <= not(layer4_outputs(2316)) or (layer4_outputs(1897));
    layer5_outputs(4312) <= layer4_outputs(4496);
    layer5_outputs(4313) <= '1';
    layer5_outputs(4314) <= not((layer4_outputs(3637)) or (layer4_outputs(2644)));
    layer5_outputs(4315) <= not((layer4_outputs(2651)) and (layer4_outputs(598)));
    layer5_outputs(4316) <= layer4_outputs(1128);
    layer5_outputs(4317) <= (layer4_outputs(3149)) or (layer4_outputs(1623));
    layer5_outputs(4318) <= not(layer4_outputs(2841));
    layer5_outputs(4319) <= '1';
    layer5_outputs(4320) <= not((layer4_outputs(3969)) and (layer4_outputs(4420)));
    layer5_outputs(4321) <= not(layer4_outputs(3299));
    layer5_outputs(4322) <= layer4_outputs(65);
    layer5_outputs(4323) <= not(layer4_outputs(835));
    layer5_outputs(4324) <= (layer4_outputs(2289)) and not (layer4_outputs(650));
    layer5_outputs(4325) <= '0';
    layer5_outputs(4326) <= not((layer4_outputs(2792)) or (layer4_outputs(2115)));
    layer5_outputs(4327) <= layer4_outputs(1633);
    layer5_outputs(4328) <= not((layer4_outputs(645)) and (layer4_outputs(1447)));
    layer5_outputs(4329) <= (layer4_outputs(4773)) or (layer4_outputs(2707));
    layer5_outputs(4330) <= '1';
    layer5_outputs(4331) <= not(layer4_outputs(1729)) or (layer4_outputs(2103));
    layer5_outputs(4332) <= layer4_outputs(1247);
    layer5_outputs(4333) <= '0';
    layer5_outputs(4334) <= not((layer4_outputs(4130)) and (layer4_outputs(479)));
    layer5_outputs(4335) <= not((layer4_outputs(3861)) or (layer4_outputs(4350)));
    layer5_outputs(4336) <= (layer4_outputs(3940)) and not (layer4_outputs(2347));
    layer5_outputs(4337) <= (layer4_outputs(4625)) and (layer4_outputs(4982));
    layer5_outputs(4338) <= (layer4_outputs(3584)) and not (layer4_outputs(1842));
    layer5_outputs(4339) <= not((layer4_outputs(3043)) xor (layer4_outputs(1819)));
    layer5_outputs(4340) <= (layer4_outputs(4404)) or (layer4_outputs(3463));
    layer5_outputs(4341) <= not(layer4_outputs(2356));
    layer5_outputs(4342) <= not(layer4_outputs(2409)) or (layer4_outputs(157));
    layer5_outputs(4343) <= layer4_outputs(4155);
    layer5_outputs(4344) <= '0';
    layer5_outputs(4345) <= layer4_outputs(2047);
    layer5_outputs(4346) <= layer4_outputs(4640);
    layer5_outputs(4347) <= not((layer4_outputs(3702)) and (layer4_outputs(4765)));
    layer5_outputs(4348) <= not((layer4_outputs(481)) and (layer4_outputs(719)));
    layer5_outputs(4349) <= layer4_outputs(1471);
    layer5_outputs(4350) <= not(layer4_outputs(4264)) or (layer4_outputs(3215));
    layer5_outputs(4351) <= layer4_outputs(2060);
    layer5_outputs(4352) <= layer4_outputs(2519);
    layer5_outputs(4353) <= (layer4_outputs(1181)) or (layer4_outputs(4702));
    layer5_outputs(4354) <= not((layer4_outputs(3641)) and (layer4_outputs(2526)));
    layer5_outputs(4355) <= '1';
    layer5_outputs(4356) <= not(layer4_outputs(2104)) or (layer4_outputs(3443));
    layer5_outputs(4357) <= '0';
    layer5_outputs(4358) <= (layer4_outputs(3483)) or (layer4_outputs(3569));
    layer5_outputs(4359) <= not(layer4_outputs(2985));
    layer5_outputs(4360) <= (layer4_outputs(1918)) or (layer4_outputs(4620));
    layer5_outputs(4361) <= not((layer4_outputs(1382)) and (layer4_outputs(25)));
    layer5_outputs(4362) <= (layer4_outputs(2752)) or (layer4_outputs(585));
    layer5_outputs(4363) <= not(layer4_outputs(4177));
    layer5_outputs(4364) <= layer4_outputs(911);
    layer5_outputs(4365) <= not(layer4_outputs(1380)) or (layer4_outputs(2415));
    layer5_outputs(4366) <= not(layer4_outputs(4923));
    layer5_outputs(4367) <= layer4_outputs(3565);
    layer5_outputs(4368) <= not(layer4_outputs(4147));
    layer5_outputs(4369) <= not(layer4_outputs(1890)) or (layer4_outputs(4468));
    layer5_outputs(4370) <= layer4_outputs(2040);
    layer5_outputs(4371) <= layer4_outputs(4063);
    layer5_outputs(4372) <= (layer4_outputs(89)) and not (layer4_outputs(3029));
    layer5_outputs(4373) <= (layer4_outputs(2798)) or (layer4_outputs(2820));
    layer5_outputs(4374) <= (layer4_outputs(3043)) and not (layer4_outputs(1063));
    layer5_outputs(4375) <= layer4_outputs(2648);
    layer5_outputs(4376) <= not((layer4_outputs(2746)) and (layer4_outputs(160)));
    layer5_outputs(4377) <= not(layer4_outputs(96)) or (layer4_outputs(2022));
    layer5_outputs(4378) <= not(layer4_outputs(2886)) or (layer4_outputs(2074));
    layer5_outputs(4379) <= not(layer4_outputs(3871)) or (layer4_outputs(4235));
    layer5_outputs(4380) <= not(layer4_outputs(1225)) or (layer4_outputs(148));
    layer5_outputs(4381) <= (layer4_outputs(4054)) and (layer4_outputs(2133));
    layer5_outputs(4382) <= layer4_outputs(4828);
    layer5_outputs(4383) <= not((layer4_outputs(4541)) or (layer4_outputs(922)));
    layer5_outputs(4384) <= layer4_outputs(3372);
    layer5_outputs(4385) <= not((layer4_outputs(1415)) xor (layer4_outputs(3967)));
    layer5_outputs(4386) <= not(layer4_outputs(2650)) or (layer4_outputs(803));
    layer5_outputs(4387) <= (layer4_outputs(4448)) and (layer4_outputs(2808));
    layer5_outputs(4388) <= not((layer4_outputs(639)) xor (layer4_outputs(1367)));
    layer5_outputs(4389) <= (layer4_outputs(677)) or (layer4_outputs(5019));
    layer5_outputs(4390) <= layer4_outputs(770);
    layer5_outputs(4391) <= not(layer4_outputs(4932));
    layer5_outputs(4392) <= not((layer4_outputs(3787)) or (layer4_outputs(1348)));
    layer5_outputs(4393) <= (layer4_outputs(2513)) or (layer4_outputs(4596));
    layer5_outputs(4394) <= (layer4_outputs(2856)) and (layer4_outputs(2513));
    layer5_outputs(4395) <= not(layer4_outputs(3291));
    layer5_outputs(4396) <= layer4_outputs(1765);
    layer5_outputs(4397) <= (layer4_outputs(4172)) and not (layer4_outputs(2538));
    layer5_outputs(4398) <= (layer4_outputs(1263)) xor (layer4_outputs(2763));
    layer5_outputs(4399) <= not(layer4_outputs(3262));
    layer5_outputs(4400) <= not((layer4_outputs(3131)) and (layer4_outputs(1449)));
    layer5_outputs(4401) <= not((layer4_outputs(2157)) or (layer4_outputs(4786)));
    layer5_outputs(4402) <= layer4_outputs(2351);
    layer5_outputs(4403) <= layer4_outputs(1636);
    layer5_outputs(4404) <= not(layer4_outputs(3841)) or (layer4_outputs(4475));
    layer5_outputs(4405) <= (layer4_outputs(4527)) and not (layer4_outputs(403));
    layer5_outputs(4406) <= not(layer4_outputs(436));
    layer5_outputs(4407) <= (layer4_outputs(61)) and (layer4_outputs(1114));
    layer5_outputs(4408) <= layer4_outputs(2787);
    layer5_outputs(4409) <= layer4_outputs(1246);
    layer5_outputs(4410) <= not(layer4_outputs(4500));
    layer5_outputs(4411) <= layer4_outputs(2704);
    layer5_outputs(4412) <= (layer4_outputs(2438)) and not (layer4_outputs(3662));
    layer5_outputs(4413) <= layer4_outputs(4407);
    layer5_outputs(4414) <= (layer4_outputs(3590)) and not (layer4_outputs(4183));
    layer5_outputs(4415) <= not((layer4_outputs(275)) and (layer4_outputs(4899)));
    layer5_outputs(4416) <= layer4_outputs(2292);
    layer5_outputs(4417) <= '1';
    layer5_outputs(4418) <= (layer4_outputs(4095)) xor (layer4_outputs(394));
    layer5_outputs(4419) <= layer4_outputs(3333);
    layer5_outputs(4420) <= layer4_outputs(2186);
    layer5_outputs(4421) <= (layer4_outputs(3907)) and (layer4_outputs(53));
    layer5_outputs(4422) <= (layer4_outputs(4857)) and not (layer4_outputs(4876));
    layer5_outputs(4423) <= (layer4_outputs(3183)) and (layer4_outputs(2406));
    layer5_outputs(4424) <= not(layer4_outputs(3798)) or (layer4_outputs(4406));
    layer5_outputs(4425) <= layer4_outputs(1035);
    layer5_outputs(4426) <= layer4_outputs(4943);
    layer5_outputs(4427) <= not(layer4_outputs(4463)) or (layer4_outputs(4687));
    layer5_outputs(4428) <= (layer4_outputs(1607)) or (layer4_outputs(3957));
    layer5_outputs(4429) <= (layer4_outputs(31)) or (layer4_outputs(3020));
    layer5_outputs(4430) <= not(layer4_outputs(3003));
    layer5_outputs(4431) <= '1';
    layer5_outputs(4432) <= not(layer4_outputs(3971)) or (layer4_outputs(3116));
    layer5_outputs(4433) <= (layer4_outputs(1938)) or (layer4_outputs(1799));
    layer5_outputs(4434) <= not(layer4_outputs(1546));
    layer5_outputs(4435) <= not(layer4_outputs(3703));
    layer5_outputs(4436) <= '0';
    layer5_outputs(4437) <= '0';
    layer5_outputs(4438) <= (layer4_outputs(3655)) and not (layer4_outputs(3377));
    layer5_outputs(4439) <= not(layer4_outputs(3610));
    layer5_outputs(4440) <= (layer4_outputs(568)) or (layer4_outputs(2811));
    layer5_outputs(4441) <= (layer4_outputs(4311)) or (layer4_outputs(2718));
    layer5_outputs(4442) <= '0';
    layer5_outputs(4443) <= not(layer4_outputs(2841));
    layer5_outputs(4444) <= not(layer4_outputs(431)) or (layer4_outputs(2942));
    layer5_outputs(4445) <= (layer4_outputs(5056)) and not (layer4_outputs(4691));
    layer5_outputs(4446) <= not(layer4_outputs(515));
    layer5_outputs(4447) <= layer4_outputs(721);
    layer5_outputs(4448) <= '0';
    layer5_outputs(4449) <= not((layer4_outputs(908)) or (layer4_outputs(3636)));
    layer5_outputs(4450) <= (layer4_outputs(1352)) and (layer4_outputs(1959));
    layer5_outputs(4451) <= not(layer4_outputs(4012));
    layer5_outputs(4452) <= not((layer4_outputs(310)) and (layer4_outputs(2523)));
    layer5_outputs(4453) <= (layer4_outputs(1521)) and not (layer4_outputs(1610));
    layer5_outputs(4454) <= (layer4_outputs(136)) and not (layer4_outputs(4027));
    layer5_outputs(4455) <= '1';
    layer5_outputs(4456) <= not((layer4_outputs(621)) and (layer4_outputs(1554)));
    layer5_outputs(4457) <= not((layer4_outputs(178)) and (layer4_outputs(5119)));
    layer5_outputs(4458) <= (layer4_outputs(4915)) or (layer4_outputs(3461));
    layer5_outputs(4459) <= layer4_outputs(2672);
    layer5_outputs(4460) <= (layer4_outputs(4673)) and not (layer4_outputs(4915));
    layer5_outputs(4461) <= (layer4_outputs(4894)) xor (layer4_outputs(3468));
    layer5_outputs(4462) <= not(layer4_outputs(2253));
    layer5_outputs(4463) <= (layer4_outputs(3303)) and not (layer4_outputs(3042));
    layer5_outputs(4464) <= (layer4_outputs(2912)) and (layer4_outputs(1789));
    layer5_outputs(4465) <= not(layer4_outputs(4639)) or (layer4_outputs(3675));
    layer5_outputs(4466) <= not(layer4_outputs(2723));
    layer5_outputs(4467) <= not((layer4_outputs(4809)) xor (layer4_outputs(1472)));
    layer5_outputs(4468) <= not(layer4_outputs(37)) or (layer4_outputs(837));
    layer5_outputs(4469) <= not(layer4_outputs(308));
    layer5_outputs(4470) <= layer4_outputs(1019);
    layer5_outputs(4471) <= not(layer4_outputs(3197));
    layer5_outputs(4472) <= '1';
    layer5_outputs(4473) <= layer4_outputs(1287);
    layer5_outputs(4474) <= not(layer4_outputs(1970));
    layer5_outputs(4475) <= not(layer4_outputs(940));
    layer5_outputs(4476) <= (layer4_outputs(1923)) or (layer4_outputs(1278));
    layer5_outputs(4477) <= not((layer4_outputs(4175)) and (layer4_outputs(255)));
    layer5_outputs(4478) <= not(layer4_outputs(4029)) or (layer4_outputs(923));
    layer5_outputs(4479) <= not(layer4_outputs(54));
    layer5_outputs(4480) <= not(layer4_outputs(3427)) or (layer4_outputs(3829));
    layer5_outputs(4481) <= '1';
    layer5_outputs(4482) <= '1';
    layer5_outputs(4483) <= not(layer4_outputs(4077));
    layer5_outputs(4484) <= (layer4_outputs(4290)) and (layer4_outputs(606));
    layer5_outputs(4485) <= not(layer4_outputs(551)) or (layer4_outputs(3371));
    layer5_outputs(4486) <= not(layer4_outputs(4081));
    layer5_outputs(4487) <= not((layer4_outputs(1322)) and (layer4_outputs(4496)));
    layer5_outputs(4488) <= not((layer4_outputs(188)) and (layer4_outputs(3543)));
    layer5_outputs(4489) <= not((layer4_outputs(1732)) xor (layer4_outputs(2846)));
    layer5_outputs(4490) <= layer4_outputs(4613);
    layer5_outputs(4491) <= layer4_outputs(463);
    layer5_outputs(4492) <= (layer4_outputs(3420)) and (layer4_outputs(4098));
    layer5_outputs(4493) <= not(layer4_outputs(599)) or (layer4_outputs(4230));
    layer5_outputs(4494) <= not(layer4_outputs(4076)) or (layer4_outputs(697));
    layer5_outputs(4495) <= (layer4_outputs(2873)) and (layer4_outputs(201));
    layer5_outputs(4496) <= not(layer4_outputs(630)) or (layer4_outputs(2440));
    layer5_outputs(4497) <= '0';
    layer5_outputs(4498) <= layer4_outputs(2839);
    layer5_outputs(4499) <= not((layer4_outputs(3669)) xor (layer4_outputs(3229)));
    layer5_outputs(4500) <= (layer4_outputs(2846)) and not (layer4_outputs(4143));
    layer5_outputs(4501) <= layer4_outputs(3166);
    layer5_outputs(4502) <= (layer4_outputs(1076)) and not (layer4_outputs(3818));
    layer5_outputs(4503) <= not(layer4_outputs(3413));
    layer5_outputs(4504) <= '1';
    layer5_outputs(4505) <= '0';
    layer5_outputs(4506) <= not(layer4_outputs(777));
    layer5_outputs(4507) <= not(layer4_outputs(1876)) or (layer4_outputs(1096));
    layer5_outputs(4508) <= '0';
    layer5_outputs(4509) <= '0';
    layer5_outputs(4510) <= not(layer4_outputs(5032)) or (layer4_outputs(3835));
    layer5_outputs(4511) <= not(layer4_outputs(1357));
    layer5_outputs(4512) <= not(layer4_outputs(2305));
    layer5_outputs(4513) <= not(layer4_outputs(2318));
    layer5_outputs(4514) <= (layer4_outputs(1792)) and not (layer4_outputs(2310));
    layer5_outputs(4515) <= not((layer4_outputs(3928)) and (layer4_outputs(51)));
    layer5_outputs(4516) <= not((layer4_outputs(1553)) or (layer4_outputs(327)));
    layer5_outputs(4517) <= (layer4_outputs(1313)) or (layer4_outputs(149));
    layer5_outputs(4518) <= '1';
    layer5_outputs(4519) <= not((layer4_outputs(4991)) or (layer4_outputs(4812)));
    layer5_outputs(4520) <= (layer4_outputs(4093)) and not (layer4_outputs(773));
    layer5_outputs(4521) <= (layer4_outputs(1291)) and not (layer4_outputs(858));
    layer5_outputs(4522) <= (layer4_outputs(961)) and not (layer4_outputs(556));
    layer5_outputs(4523) <= not(layer4_outputs(866)) or (layer4_outputs(1999));
    layer5_outputs(4524) <= '0';
    layer5_outputs(4525) <= (layer4_outputs(2163)) and not (layer4_outputs(903));
    layer5_outputs(4526) <= (layer4_outputs(298)) and not (layer4_outputs(1209));
    layer5_outputs(4527) <= '0';
    layer5_outputs(4528) <= not(layer4_outputs(32));
    layer5_outputs(4529) <= layer4_outputs(3024);
    layer5_outputs(4530) <= layer4_outputs(917);
    layer5_outputs(4531) <= not(layer4_outputs(666));
    layer5_outputs(4532) <= layer4_outputs(3037);
    layer5_outputs(4533) <= layer4_outputs(2153);
    layer5_outputs(4534) <= layer4_outputs(1631);
    layer5_outputs(4535) <= (layer4_outputs(39)) and not (layer4_outputs(2068));
    layer5_outputs(4536) <= not(layer4_outputs(386));
    layer5_outputs(4537) <= not(layer4_outputs(1601));
    layer5_outputs(4538) <= layer4_outputs(3712);
    layer5_outputs(4539) <= (layer4_outputs(3257)) and not (layer4_outputs(2422));
    layer5_outputs(4540) <= (layer4_outputs(575)) and not (layer4_outputs(1604));
    layer5_outputs(4541) <= layer4_outputs(2470);
    layer5_outputs(4542) <= not((layer4_outputs(274)) or (layer4_outputs(316)));
    layer5_outputs(4543) <= not((layer4_outputs(1160)) xor (layer4_outputs(3639)));
    layer5_outputs(4544) <= not(layer4_outputs(3033));
    layer5_outputs(4545) <= not(layer4_outputs(792));
    layer5_outputs(4546) <= not(layer4_outputs(4320)) or (layer4_outputs(1052));
    layer5_outputs(4547) <= not(layer4_outputs(4122));
    layer5_outputs(4548) <= (layer4_outputs(2097)) xor (layer4_outputs(3316));
    layer5_outputs(4549) <= (layer4_outputs(3962)) and not (layer4_outputs(4331));
    layer5_outputs(4550) <= not(layer4_outputs(4529));
    layer5_outputs(4551) <= (layer4_outputs(1211)) and (layer4_outputs(2607));
    layer5_outputs(4552) <= layer4_outputs(3089);
    layer5_outputs(4553) <= not(layer4_outputs(2033));
    layer5_outputs(4554) <= (layer4_outputs(2129)) or (layer4_outputs(4282));
    layer5_outputs(4555) <= layer4_outputs(2450);
    layer5_outputs(4556) <= not(layer4_outputs(1762));
    layer5_outputs(4557) <= not((layer4_outputs(1994)) or (layer4_outputs(2367)));
    layer5_outputs(4558) <= layer4_outputs(3243);
    layer5_outputs(4559) <= not((layer4_outputs(534)) and (layer4_outputs(3758)));
    layer5_outputs(4560) <= (layer4_outputs(1347)) and not (layer4_outputs(1899));
    layer5_outputs(4561) <= not(layer4_outputs(4942)) or (layer4_outputs(2180));
    layer5_outputs(4562) <= not(layer4_outputs(442)) or (layer4_outputs(2360));
    layer5_outputs(4563) <= (layer4_outputs(1184)) and (layer4_outputs(2447));
    layer5_outputs(4564) <= not(layer4_outputs(3218)) or (layer4_outputs(3923));
    layer5_outputs(4565) <= not((layer4_outputs(2495)) or (layer4_outputs(2193)));
    layer5_outputs(4566) <= '1';
    layer5_outputs(4567) <= '1';
    layer5_outputs(4568) <= not((layer4_outputs(4778)) and (layer4_outputs(3452)));
    layer5_outputs(4569) <= not(layer4_outputs(2564)) or (layer4_outputs(2234));
    layer5_outputs(4570) <= layer4_outputs(3256);
    layer5_outputs(4571) <= not(layer4_outputs(2959)) or (layer4_outputs(3006));
    layer5_outputs(4572) <= '1';
    layer5_outputs(4573) <= not(layer4_outputs(2985)) or (layer4_outputs(4782));
    layer5_outputs(4574) <= (layer4_outputs(3804)) and not (layer4_outputs(2654));
    layer5_outputs(4575) <= not((layer4_outputs(1076)) xor (layer4_outputs(1394)));
    layer5_outputs(4576) <= (layer4_outputs(4501)) and not (layer4_outputs(4977));
    layer5_outputs(4577) <= '1';
    layer5_outputs(4578) <= layer4_outputs(3226);
    layer5_outputs(4579) <= not(layer4_outputs(2952));
    layer5_outputs(4580) <= '1';
    layer5_outputs(4581) <= not(layer4_outputs(1082));
    layer5_outputs(4582) <= (layer4_outputs(2969)) and not (layer4_outputs(430));
    layer5_outputs(4583) <= (layer4_outputs(1237)) and not (layer4_outputs(2949));
    layer5_outputs(4584) <= not(layer4_outputs(2108));
    layer5_outputs(4585) <= not(layer4_outputs(4048));
    layer5_outputs(4586) <= not((layer4_outputs(4294)) and (layer4_outputs(5098)));
    layer5_outputs(4587) <= not((layer4_outputs(1888)) or (layer4_outputs(1974)));
    layer5_outputs(4588) <= not(layer4_outputs(2772)) or (layer4_outputs(425));
    layer5_outputs(4589) <= (layer4_outputs(2101)) and not (layer4_outputs(1935));
    layer5_outputs(4590) <= layer4_outputs(46);
    layer5_outputs(4591) <= (layer4_outputs(4507)) and not (layer4_outputs(2140));
    layer5_outputs(4592) <= (layer4_outputs(2638)) or (layer4_outputs(4238));
    layer5_outputs(4593) <= (layer4_outputs(2645)) or (layer4_outputs(477));
    layer5_outputs(4594) <= not(layer4_outputs(2658)) or (layer4_outputs(4983));
    layer5_outputs(4595) <= not(layer4_outputs(4946));
    layer5_outputs(4596) <= not((layer4_outputs(2988)) and (layer4_outputs(1567)));
    layer5_outputs(4597) <= not(layer4_outputs(1390));
    layer5_outputs(4598) <= (layer4_outputs(1590)) and not (layer4_outputs(2531));
    layer5_outputs(4599) <= not((layer4_outputs(4317)) and (layer4_outputs(4176)));
    layer5_outputs(4600) <= not((layer4_outputs(4311)) xor (layer4_outputs(890)));
    layer5_outputs(4601) <= (layer4_outputs(3653)) and not (layer4_outputs(759));
    layer5_outputs(4602) <= not(layer4_outputs(1881)) or (layer4_outputs(1727));
    layer5_outputs(4603) <= not((layer4_outputs(4224)) or (layer4_outputs(1703)));
    layer5_outputs(4604) <= not(layer4_outputs(2189));
    layer5_outputs(4605) <= not(layer4_outputs(3570)) or (layer4_outputs(2964));
    layer5_outputs(4606) <= (layer4_outputs(2002)) and not (layer4_outputs(2989));
    layer5_outputs(4607) <= (layer4_outputs(2426)) and not (layer4_outputs(2745));
    layer5_outputs(4608) <= not(layer4_outputs(202)) or (layer4_outputs(3678));
    layer5_outputs(4609) <= layer4_outputs(3415);
    layer5_outputs(4610) <= not(layer4_outputs(3982));
    layer5_outputs(4611) <= '0';
    layer5_outputs(4612) <= not(layer4_outputs(494)) or (layer4_outputs(2334));
    layer5_outputs(4613) <= (layer4_outputs(3989)) and not (layer4_outputs(1047));
    layer5_outputs(4614) <= (layer4_outputs(2070)) and (layer4_outputs(571));
    layer5_outputs(4615) <= layer4_outputs(577);
    layer5_outputs(4616) <= layer4_outputs(1404);
    layer5_outputs(4617) <= layer4_outputs(2871);
    layer5_outputs(4618) <= layer4_outputs(4804);
    layer5_outputs(4619) <= not(layer4_outputs(3119)) or (layer4_outputs(510));
    layer5_outputs(4620) <= (layer4_outputs(3958)) and (layer4_outputs(1141));
    layer5_outputs(4621) <= not((layer4_outputs(3299)) and (layer4_outputs(927)));
    layer5_outputs(4622) <= not((layer4_outputs(4684)) xor (layer4_outputs(2368)));
    layer5_outputs(4623) <= layer4_outputs(4154);
    layer5_outputs(4624) <= (layer4_outputs(537)) and not (layer4_outputs(1697));
    layer5_outputs(4625) <= not(layer4_outputs(4030)) or (layer4_outputs(4992));
    layer5_outputs(4626) <= layer4_outputs(2894);
    layer5_outputs(4627) <= layer4_outputs(3328);
    layer5_outputs(4628) <= (layer4_outputs(3152)) and not (layer4_outputs(4601));
    layer5_outputs(4629) <= (layer4_outputs(1963)) and (layer4_outputs(3555));
    layer5_outputs(4630) <= (layer4_outputs(3539)) and (layer4_outputs(64));
    layer5_outputs(4631) <= not(layer4_outputs(3113));
    layer5_outputs(4632) <= (layer4_outputs(4083)) xor (layer4_outputs(1252));
    layer5_outputs(4633) <= layer4_outputs(135);
    layer5_outputs(4634) <= layer4_outputs(2107);
    layer5_outputs(4635) <= layer4_outputs(724);
    layer5_outputs(4636) <= layer4_outputs(2399);
    layer5_outputs(4637) <= (layer4_outputs(577)) and not (layer4_outputs(1551));
    layer5_outputs(4638) <= not((layer4_outputs(2653)) or (layer4_outputs(125)));
    layer5_outputs(4639) <= layer4_outputs(1231);
    layer5_outputs(4640) <= layer4_outputs(2723);
    layer5_outputs(4641) <= (layer4_outputs(2285)) and (layer4_outputs(3641));
    layer5_outputs(4642) <= (layer4_outputs(3100)) and (layer4_outputs(1140));
    layer5_outputs(4643) <= (layer4_outputs(4761)) and (layer4_outputs(2835));
    layer5_outputs(4644) <= layer4_outputs(1333);
    layer5_outputs(4645) <= (layer4_outputs(2017)) and not (layer4_outputs(3168));
    layer5_outputs(4646) <= '1';
    layer5_outputs(4647) <= not(layer4_outputs(3528)) or (layer4_outputs(3874));
    layer5_outputs(4648) <= not(layer4_outputs(3019)) or (layer4_outputs(3033));
    layer5_outputs(4649) <= not(layer4_outputs(566)) or (layer4_outputs(767));
    layer5_outputs(4650) <= not(layer4_outputs(3385));
    layer5_outputs(4651) <= layer4_outputs(3310);
    layer5_outputs(4652) <= layer4_outputs(2974);
    layer5_outputs(4653) <= (layer4_outputs(1805)) or (layer4_outputs(308));
    layer5_outputs(4654) <= not(layer4_outputs(3815));
    layer5_outputs(4655) <= not(layer4_outputs(1197));
    layer5_outputs(4656) <= not((layer4_outputs(1320)) and (layer4_outputs(466)));
    layer5_outputs(4657) <= (layer4_outputs(4424)) and not (layer4_outputs(4493));
    layer5_outputs(4658) <= layer4_outputs(3457);
    layer5_outputs(4659) <= layer4_outputs(919);
    layer5_outputs(4660) <= not((layer4_outputs(1565)) and (layer4_outputs(1064)));
    layer5_outputs(4661) <= not(layer4_outputs(3436));
    layer5_outputs(4662) <= layer4_outputs(2576);
    layer5_outputs(4663) <= not(layer4_outputs(842));
    layer5_outputs(4664) <= not(layer4_outputs(2908));
    layer5_outputs(4665) <= layer4_outputs(3172);
    layer5_outputs(4666) <= not(layer4_outputs(2011));
    layer5_outputs(4667) <= not(layer4_outputs(2591)) or (layer4_outputs(586));
    layer5_outputs(4668) <= '1';
    layer5_outputs(4669) <= (layer4_outputs(3210)) and not (layer4_outputs(3826));
    layer5_outputs(4670) <= not(layer4_outputs(5073));
    layer5_outputs(4671) <= layer4_outputs(1785);
    layer5_outputs(4672) <= (layer4_outputs(4041)) and not (layer4_outputs(1250));
    layer5_outputs(4673) <= (layer4_outputs(4237)) and not (layer4_outputs(4190));
    layer5_outputs(4674) <= '1';
    layer5_outputs(4675) <= layer4_outputs(3374);
    layer5_outputs(4676) <= not(layer4_outputs(568));
    layer5_outputs(4677) <= not((layer4_outputs(405)) or (layer4_outputs(1708)));
    layer5_outputs(4678) <= (layer4_outputs(2299)) or (layer4_outputs(1127));
    layer5_outputs(4679) <= not(layer4_outputs(4155));
    layer5_outputs(4680) <= '1';
    layer5_outputs(4681) <= '0';
    layer5_outputs(4682) <= (layer4_outputs(2965)) and not (layer4_outputs(3438));
    layer5_outputs(4683) <= not((layer4_outputs(1703)) or (layer4_outputs(4436)));
    layer5_outputs(4684) <= (layer4_outputs(2137)) and not (layer4_outputs(81));
    layer5_outputs(4685) <= (layer4_outputs(1207)) and not (layer4_outputs(2853));
    layer5_outputs(4686) <= layer4_outputs(179);
    layer5_outputs(4687) <= '0';
    layer5_outputs(4688) <= (layer4_outputs(1188)) and not (layer4_outputs(3274));
    layer5_outputs(4689) <= layer4_outputs(2711);
    layer5_outputs(4690) <= (layer4_outputs(1222)) or (layer4_outputs(4142));
    layer5_outputs(4691) <= layer4_outputs(3648);
    layer5_outputs(4692) <= not((layer4_outputs(4396)) or (layer4_outputs(4820)));
    layer5_outputs(4693) <= not(layer4_outputs(1599));
    layer5_outputs(4694) <= (layer4_outputs(1385)) and not (layer4_outputs(347));
    layer5_outputs(4695) <= (layer4_outputs(995)) and not (layer4_outputs(4768));
    layer5_outputs(4696) <= '1';
    layer5_outputs(4697) <= not((layer4_outputs(4297)) or (layer4_outputs(2319)));
    layer5_outputs(4698) <= (layer4_outputs(2857)) or (layer4_outputs(1990));
    layer5_outputs(4699) <= (layer4_outputs(1862)) xor (layer4_outputs(2923));
    layer5_outputs(4700) <= not((layer4_outputs(1345)) xor (layer4_outputs(463)));
    layer5_outputs(4701) <= layer4_outputs(3327);
    layer5_outputs(4702) <= not((layer4_outputs(1593)) xor (layer4_outputs(4580)));
    layer5_outputs(4703) <= (layer4_outputs(2634)) and not (layer4_outputs(2622));
    layer5_outputs(4704) <= (layer4_outputs(3948)) and not (layer4_outputs(1616));
    layer5_outputs(4705) <= not(layer4_outputs(413));
    layer5_outputs(4706) <= (layer4_outputs(111)) xor (layer4_outputs(1967));
    layer5_outputs(4707) <= not((layer4_outputs(3949)) and (layer4_outputs(3011)));
    layer5_outputs(4708) <= '0';
    layer5_outputs(4709) <= (layer4_outputs(815)) or (layer4_outputs(874));
    layer5_outputs(4710) <= not(layer4_outputs(55)) or (layer4_outputs(2950));
    layer5_outputs(4711) <= not(layer4_outputs(1699));
    layer5_outputs(4712) <= layer4_outputs(4025);
    layer5_outputs(4713) <= not((layer4_outputs(1452)) or (layer4_outputs(4395)));
    layer5_outputs(4714) <= (layer4_outputs(5050)) or (layer4_outputs(1902));
    layer5_outputs(4715) <= (layer4_outputs(1222)) or (layer4_outputs(3793));
    layer5_outputs(4716) <= '0';
    layer5_outputs(4717) <= not(layer4_outputs(1815));
    layer5_outputs(4718) <= (layer4_outputs(2314)) or (layer4_outputs(5075));
    layer5_outputs(4719) <= (layer4_outputs(478)) or (layer4_outputs(4185));
    layer5_outputs(4720) <= layer4_outputs(4492);
    layer5_outputs(4721) <= not(layer4_outputs(799));
    layer5_outputs(4722) <= (layer4_outputs(2323)) and (layer4_outputs(625));
    layer5_outputs(4723) <= not((layer4_outputs(1677)) and (layer4_outputs(142)));
    layer5_outputs(4724) <= not(layer4_outputs(949)) or (layer4_outputs(2037));
    layer5_outputs(4725) <= not(layer4_outputs(3157));
    layer5_outputs(4726) <= not(layer4_outputs(4967)) or (layer4_outputs(2280));
    layer5_outputs(4727) <= layer4_outputs(1930);
    layer5_outputs(4728) <= layer4_outputs(4531);
    layer5_outputs(4729) <= not((layer4_outputs(1534)) xor (layer4_outputs(1221)));
    layer5_outputs(4730) <= (layer4_outputs(646)) or (layer4_outputs(24));
    layer5_outputs(4731) <= not(layer4_outputs(2635));
    layer5_outputs(4732) <= not(layer4_outputs(1704)) or (layer4_outputs(4670));
    layer5_outputs(4733) <= not((layer4_outputs(3525)) and (layer4_outputs(2155)));
    layer5_outputs(4734) <= (layer4_outputs(2095)) and (layer4_outputs(4562));
    layer5_outputs(4735) <= not((layer4_outputs(4587)) xor (layer4_outputs(177)));
    layer5_outputs(4736) <= (layer4_outputs(3809)) xor (layer4_outputs(3739));
    layer5_outputs(4737) <= layer4_outputs(4300);
    layer5_outputs(4738) <= '1';
    layer5_outputs(4739) <= (layer4_outputs(3238)) and (layer4_outputs(1243));
    layer5_outputs(4740) <= '0';
    layer5_outputs(4741) <= layer4_outputs(4493);
    layer5_outputs(4742) <= (layer4_outputs(3680)) and (layer4_outputs(4877));
    layer5_outputs(4743) <= (layer4_outputs(613)) and not (layer4_outputs(4295));
    layer5_outputs(4744) <= not(layer4_outputs(2205)) or (layer4_outputs(2152));
    layer5_outputs(4745) <= not(layer4_outputs(3960)) or (layer4_outputs(1118));
    layer5_outputs(4746) <= layer4_outputs(4650);
    layer5_outputs(4747) <= (layer4_outputs(534)) and not (layer4_outputs(2737));
    layer5_outputs(4748) <= not((layer4_outputs(2785)) xor (layer4_outputs(3593)));
    layer5_outputs(4749) <= layer4_outputs(4308);
    layer5_outputs(4750) <= not((layer4_outputs(1019)) xor (layer4_outputs(4125)));
    layer5_outputs(4751) <= not((layer4_outputs(2417)) and (layer4_outputs(2149)));
    layer5_outputs(4752) <= (layer4_outputs(155)) and not (layer4_outputs(2860));
    layer5_outputs(4753) <= layer4_outputs(4547);
    layer5_outputs(4754) <= not((layer4_outputs(2992)) xor (layer4_outputs(2934)));
    layer5_outputs(4755) <= not(layer4_outputs(3211)) or (layer4_outputs(4105));
    layer5_outputs(4756) <= not((layer4_outputs(1822)) xor (layer4_outputs(3027)));
    layer5_outputs(4757) <= layer4_outputs(2072);
    layer5_outputs(4758) <= not((layer4_outputs(3978)) and (layer4_outputs(996)));
    layer5_outputs(4759) <= (layer4_outputs(2524)) xor (layer4_outputs(3737));
    layer5_outputs(4760) <= not((layer4_outputs(3369)) or (layer4_outputs(1569)));
    layer5_outputs(4761) <= layer4_outputs(580);
    layer5_outputs(4762) <= not(layer4_outputs(4988)) or (layer4_outputs(2962));
    layer5_outputs(4763) <= not((layer4_outputs(1309)) and (layer4_outputs(2645)));
    layer5_outputs(4764) <= not(layer4_outputs(1987));
    layer5_outputs(4765) <= not(layer4_outputs(3084)) or (layer4_outputs(1907));
    layer5_outputs(4766) <= not(layer4_outputs(1886));
    layer5_outputs(4767) <= (layer4_outputs(2187)) and not (layer4_outputs(2075));
    layer5_outputs(4768) <= '1';
    layer5_outputs(4769) <= layer4_outputs(5035);
    layer5_outputs(4770) <= layer4_outputs(488);
    layer5_outputs(4771) <= not(layer4_outputs(2094));
    layer5_outputs(4772) <= '1';
    layer5_outputs(4773) <= (layer4_outputs(4253)) and (layer4_outputs(2768));
    layer5_outputs(4774) <= (layer4_outputs(2827)) xor (layer4_outputs(4916));
    layer5_outputs(4775) <= not((layer4_outputs(3846)) and (layer4_outputs(473)));
    layer5_outputs(4776) <= layer4_outputs(4651);
    layer5_outputs(4777) <= layer4_outputs(238);
    layer5_outputs(4778) <= not(layer4_outputs(3303));
    layer5_outputs(4779) <= not(layer4_outputs(1043));
    layer5_outputs(4780) <= (layer4_outputs(3628)) or (layer4_outputs(161));
    layer5_outputs(4781) <= (layer4_outputs(3408)) and not (layer4_outputs(4174));
    layer5_outputs(4782) <= not(layer4_outputs(1786));
    layer5_outputs(4783) <= (layer4_outputs(1995)) and (layer4_outputs(919));
    layer5_outputs(4784) <= layer4_outputs(2279);
    layer5_outputs(4785) <= (layer4_outputs(4939)) and (layer4_outputs(299));
    layer5_outputs(4786) <= not(layer4_outputs(1884));
    layer5_outputs(4787) <= (layer4_outputs(4984)) xor (layer4_outputs(3762));
    layer5_outputs(4788) <= not((layer4_outputs(1567)) or (layer4_outputs(782)));
    layer5_outputs(4789) <= not(layer4_outputs(3709));
    layer5_outputs(4790) <= layer4_outputs(68);
    layer5_outputs(4791) <= (layer4_outputs(682)) or (layer4_outputs(784));
    layer5_outputs(4792) <= not(layer4_outputs(2816)) or (layer4_outputs(3352));
    layer5_outputs(4793) <= not(layer4_outputs(4211)) or (layer4_outputs(4545));
    layer5_outputs(4794) <= layer4_outputs(1157);
    layer5_outputs(4795) <= (layer4_outputs(2563)) or (layer4_outputs(3870));
    layer5_outputs(4796) <= (layer4_outputs(3494)) and not (layer4_outputs(5116));
    layer5_outputs(4797) <= layer4_outputs(3290);
    layer5_outputs(4798) <= '1';
    layer5_outputs(4799) <= (layer4_outputs(251)) or (layer4_outputs(2010));
    layer5_outputs(4800) <= (layer4_outputs(181)) or (layer4_outputs(3264));
    layer5_outputs(4801) <= layer4_outputs(3207);
    layer5_outputs(4802) <= (layer4_outputs(4402)) or (layer4_outputs(4120));
    layer5_outputs(4803) <= layer4_outputs(1621);
    layer5_outputs(4804) <= (layer4_outputs(1656)) or (layer4_outputs(4961));
    layer5_outputs(4805) <= not((layer4_outputs(1195)) and (layer4_outputs(1802)));
    layer5_outputs(4806) <= not(layer4_outputs(4059));
    layer5_outputs(4807) <= (layer4_outputs(1708)) and not (layer4_outputs(2962));
    layer5_outputs(4808) <= (layer4_outputs(3181)) and (layer4_outputs(4836));
    layer5_outputs(4809) <= layer4_outputs(412);
    layer5_outputs(4810) <= layer4_outputs(1937);
    layer5_outputs(4811) <= not((layer4_outputs(635)) and (layer4_outputs(3644)));
    layer5_outputs(4812) <= not((layer4_outputs(2705)) or (layer4_outputs(2026)));
    layer5_outputs(4813) <= (layer4_outputs(1831)) and not (layer4_outputs(2046));
    layer5_outputs(4814) <= '1';
    layer5_outputs(4815) <= layer4_outputs(3671);
    layer5_outputs(4816) <= layer4_outputs(3713);
    layer5_outputs(4817) <= layer4_outputs(1812);
    layer5_outputs(4818) <= not(layer4_outputs(3282));
    layer5_outputs(4819) <= (layer4_outputs(939)) xor (layer4_outputs(2791));
    layer5_outputs(4820) <= not(layer4_outputs(3007));
    layer5_outputs(4821) <= (layer4_outputs(4351)) and not (layer4_outputs(2818));
    layer5_outputs(4822) <= not(layer4_outputs(103));
    layer5_outputs(4823) <= (layer4_outputs(3430)) and (layer4_outputs(1370));
    layer5_outputs(4824) <= not((layer4_outputs(60)) or (layer4_outputs(3658)));
    layer5_outputs(4825) <= not(layer4_outputs(2308));
    layer5_outputs(4826) <= '1';
    layer5_outputs(4827) <= layer4_outputs(2608);
    layer5_outputs(4828) <= not((layer4_outputs(732)) or (layer4_outputs(4256)));
    layer5_outputs(4829) <= (layer4_outputs(2483)) and not (layer4_outputs(115));
    layer5_outputs(4830) <= '0';
    layer5_outputs(4831) <= not(layer4_outputs(1681)) or (layer4_outputs(3027));
    layer5_outputs(4832) <= not(layer4_outputs(1605)) or (layer4_outputs(3355));
    layer5_outputs(4833) <= (layer4_outputs(3806)) and (layer4_outputs(2499));
    layer5_outputs(4834) <= '1';
    layer5_outputs(4835) <= not(layer4_outputs(4147)) or (layer4_outputs(3326));
    layer5_outputs(4836) <= '0';
    layer5_outputs(4837) <= not(layer4_outputs(669));
    layer5_outputs(4838) <= layer4_outputs(4268);
    layer5_outputs(4839) <= not(layer4_outputs(2901));
    layer5_outputs(4840) <= not((layer4_outputs(757)) or (layer4_outputs(137)));
    layer5_outputs(4841) <= not(layer4_outputs(1742)) or (layer4_outputs(3254));
    layer5_outputs(4842) <= (layer4_outputs(3541)) and not (layer4_outputs(1045));
    layer5_outputs(4843) <= not((layer4_outputs(1869)) and (layer4_outputs(215)));
    layer5_outputs(4844) <= (layer4_outputs(4957)) and (layer4_outputs(1251));
    layer5_outputs(4845) <= not(layer4_outputs(4164));
    layer5_outputs(4846) <= (layer4_outputs(3020)) or (layer4_outputs(4459));
    layer5_outputs(4847) <= not(layer4_outputs(5054)) or (layer4_outputs(1774));
    layer5_outputs(4848) <= layer4_outputs(1991);
    layer5_outputs(4849) <= not((layer4_outputs(82)) and (layer4_outputs(3619)));
    layer5_outputs(4850) <= (layer4_outputs(3975)) or (layer4_outputs(4096));
    layer5_outputs(4851) <= '1';
    layer5_outputs(4852) <= (layer4_outputs(4153)) or (layer4_outputs(1566));
    layer5_outputs(4853) <= not(layer4_outputs(1435));
    layer5_outputs(4854) <= not(layer4_outputs(4205));
    layer5_outputs(4855) <= layer4_outputs(2654);
    layer5_outputs(4856) <= '1';
    layer5_outputs(4857) <= not((layer4_outputs(2185)) or (layer4_outputs(4330)));
    layer5_outputs(4858) <= (layer4_outputs(3394)) and not (layer4_outputs(1441));
    layer5_outputs(4859) <= (layer4_outputs(516)) and not (layer4_outputs(3373));
    layer5_outputs(4860) <= layer4_outputs(1982);
    layer5_outputs(4861) <= not(layer4_outputs(1661)) or (layer4_outputs(1303));
    layer5_outputs(4862) <= (layer4_outputs(3364)) and (layer4_outputs(848));
    layer5_outputs(4863) <= layer4_outputs(2297);
    layer5_outputs(4864) <= not(layer4_outputs(5008));
    layer5_outputs(4865) <= layer4_outputs(2905);
    layer5_outputs(4866) <= not((layer4_outputs(2190)) and (layer4_outputs(1923)));
    layer5_outputs(4867) <= not(layer4_outputs(1078));
    layer5_outputs(4868) <= not(layer4_outputs(4333)) or (layer4_outputs(4112));
    layer5_outputs(4869) <= (layer4_outputs(2009)) and not (layer4_outputs(1083));
    layer5_outputs(4870) <= layer4_outputs(2909);
    layer5_outputs(4871) <= '1';
    layer5_outputs(4872) <= '0';
    layer5_outputs(4873) <= not(layer4_outputs(1969));
    layer5_outputs(4874) <= layer4_outputs(149);
    layer5_outputs(4875) <= not(layer4_outputs(1896));
    layer5_outputs(4876) <= not(layer4_outputs(872));
    layer5_outputs(4877) <= not(layer4_outputs(774));
    layer5_outputs(4878) <= (layer4_outputs(4247)) or (layer4_outputs(1823));
    layer5_outputs(4879) <= not(layer4_outputs(4075));
    layer5_outputs(4880) <= not((layer4_outputs(4134)) or (layer4_outputs(3348)));
    layer5_outputs(4881) <= layer4_outputs(4370);
    layer5_outputs(4882) <= (layer4_outputs(2032)) and (layer4_outputs(4182));
    layer5_outputs(4883) <= not(layer4_outputs(4935)) or (layer4_outputs(158));
    layer5_outputs(4884) <= layer4_outputs(1061);
    layer5_outputs(4885) <= layer4_outputs(203);
    layer5_outputs(4886) <= not(layer4_outputs(4890)) or (layer4_outputs(827));
    layer5_outputs(4887) <= (layer4_outputs(9)) and not (layer4_outputs(3558));
    layer5_outputs(4888) <= not((layer4_outputs(3540)) and (layer4_outputs(1673)));
    layer5_outputs(4889) <= not(layer4_outputs(5017));
    layer5_outputs(4890) <= layer4_outputs(3528);
    layer5_outputs(4891) <= '0';
    layer5_outputs(4892) <= not(layer4_outputs(1084)) or (layer4_outputs(3902));
    layer5_outputs(4893) <= '0';
    layer5_outputs(4894) <= not(layer4_outputs(3410));
    layer5_outputs(4895) <= '1';
    layer5_outputs(4896) <= not(layer4_outputs(4140)) or (layer4_outputs(2529));
    layer5_outputs(4897) <= not(layer4_outputs(5056)) or (layer4_outputs(2130));
    layer5_outputs(4898) <= not(layer4_outputs(2950)) or (layer4_outputs(3429));
    layer5_outputs(4899) <= '1';
    layer5_outputs(4900) <= not(layer4_outputs(2473)) or (layer4_outputs(659));
    layer5_outputs(4901) <= (layer4_outputs(642)) and not (layer4_outputs(1161));
    layer5_outputs(4902) <= not(layer4_outputs(3228));
    layer5_outputs(4903) <= (layer4_outputs(1483)) and (layer4_outputs(4686));
    layer5_outputs(4904) <= not(layer4_outputs(1555));
    layer5_outputs(4905) <= (layer4_outputs(167)) and (layer4_outputs(850));
    layer5_outputs(4906) <= (layer4_outputs(1849)) and not (layer4_outputs(110));
    layer5_outputs(4907) <= layer4_outputs(5023);
    layer5_outputs(4908) <= not((layer4_outputs(5103)) and (layer4_outputs(3250)));
    layer5_outputs(4909) <= layer4_outputs(564);
    layer5_outputs(4910) <= layer4_outputs(2188);
    layer5_outputs(4911) <= not(layer4_outputs(3559)) or (layer4_outputs(2045));
    layer5_outputs(4912) <= (layer4_outputs(3195)) or (layer4_outputs(638));
    layer5_outputs(4913) <= not(layer4_outputs(4253)) or (layer4_outputs(845));
    layer5_outputs(4914) <= layer4_outputs(2156);
    layer5_outputs(4915) <= (layer4_outputs(1699)) and not (layer4_outputs(30));
    layer5_outputs(4916) <= not(layer4_outputs(3360)) or (layer4_outputs(2261));
    layer5_outputs(4917) <= not(layer4_outputs(4481));
    layer5_outputs(4918) <= (layer4_outputs(4641)) xor (layer4_outputs(3942));
    layer5_outputs(4919) <= not(layer4_outputs(3136));
    layer5_outputs(4920) <= layer4_outputs(1267);
    layer5_outputs(4921) <= not(layer4_outputs(3467));
    layer5_outputs(4922) <= not(layer4_outputs(3824));
    layer5_outputs(4923) <= (layer4_outputs(85)) and not (layer4_outputs(4634));
    layer5_outputs(4924) <= (layer4_outputs(2672)) and not (layer4_outputs(1759));
    layer5_outputs(4925) <= (layer4_outputs(3849)) and (layer4_outputs(29));
    layer5_outputs(4926) <= layer4_outputs(5026);
    layer5_outputs(4927) <= layer4_outputs(2588);
    layer5_outputs(4928) <= layer4_outputs(1205);
    layer5_outputs(4929) <= not(layer4_outputs(3301)) or (layer4_outputs(4160));
    layer5_outputs(4930) <= (layer4_outputs(3362)) and (layer4_outputs(3111));
    layer5_outputs(4931) <= not(layer4_outputs(2417));
    layer5_outputs(4932) <= not(layer4_outputs(211));
    layer5_outputs(4933) <= not(layer4_outputs(2767)) or (layer4_outputs(478));
    layer5_outputs(4934) <= not((layer4_outputs(1787)) or (layer4_outputs(4505)));
    layer5_outputs(4935) <= (layer4_outputs(1297)) or (layer4_outputs(4808));
    layer5_outputs(4936) <= (layer4_outputs(219)) or (layer4_outputs(4313));
    layer5_outputs(4937) <= layer4_outputs(2528);
    layer5_outputs(4938) <= not(layer4_outputs(1940)) or (layer4_outputs(5099));
    layer5_outputs(4939) <= not((layer4_outputs(804)) xor (layer4_outputs(4913)));
    layer5_outputs(4940) <= '1';
    layer5_outputs(4941) <= (layer4_outputs(2788)) and (layer4_outputs(2229));
    layer5_outputs(4942) <= layer4_outputs(2167);
    layer5_outputs(4943) <= layer4_outputs(4410);
    layer5_outputs(4944) <= not(layer4_outputs(525));
    layer5_outputs(4945) <= not(layer4_outputs(3071)) or (layer4_outputs(4291));
    layer5_outputs(4946) <= (layer4_outputs(4852)) or (layer4_outputs(2270));
    layer5_outputs(4947) <= (layer4_outputs(1731)) or (layer4_outputs(1678));
    layer5_outputs(4948) <= '0';
    layer5_outputs(4949) <= (layer4_outputs(695)) and (layer4_outputs(1913));
    layer5_outputs(4950) <= not((layer4_outputs(1434)) xor (layer4_outputs(1848)));
    layer5_outputs(4951) <= not((layer4_outputs(3554)) and (layer4_outputs(4031)));
    layer5_outputs(4952) <= not((layer4_outputs(1400)) and (layer4_outputs(1794)));
    layer5_outputs(4953) <= not(layer4_outputs(4345));
    layer5_outputs(4954) <= not(layer4_outputs(4125));
    layer5_outputs(4955) <= '0';
    layer5_outputs(4956) <= not(layer4_outputs(2275)) or (layer4_outputs(154));
    layer5_outputs(4957) <= layer4_outputs(1489);
    layer5_outputs(4958) <= not((layer4_outputs(3410)) xor (layer4_outputs(3899)));
    layer5_outputs(4959) <= layer4_outputs(522);
    layer5_outputs(4960) <= not(layer4_outputs(284)) or (layer4_outputs(2119));
    layer5_outputs(4961) <= layer4_outputs(3777);
    layer5_outputs(4962) <= not(layer4_outputs(1366)) or (layer4_outputs(2445));
    layer5_outputs(4963) <= not(layer4_outputs(2608)) or (layer4_outputs(4218));
    layer5_outputs(4964) <= (layer4_outputs(453)) and not (layer4_outputs(991));
    layer5_outputs(4965) <= (layer4_outputs(2023)) xor (layer4_outputs(2128));
    layer5_outputs(4966) <= (layer4_outputs(2294)) or (layer4_outputs(1889));
    layer5_outputs(4967) <= not(layer4_outputs(452)) or (layer4_outputs(3584));
    layer5_outputs(4968) <= layer4_outputs(1253);
    layer5_outputs(4969) <= (layer4_outputs(212)) and not (layer4_outputs(2851));
    layer5_outputs(4970) <= not(layer4_outputs(501)) or (layer4_outputs(1947));
    layer5_outputs(4971) <= not(layer4_outputs(3097));
    layer5_outputs(4972) <= (layer4_outputs(788)) and not (layer4_outputs(2136));
    layer5_outputs(4973) <= (layer4_outputs(2099)) and not (layer4_outputs(2440));
    layer5_outputs(4974) <= layer4_outputs(3327);
    layer5_outputs(4975) <= not((layer4_outputs(1557)) and (layer4_outputs(548)));
    layer5_outputs(4976) <= (layer4_outputs(261)) or (layer4_outputs(2541));
    layer5_outputs(4977) <= layer4_outputs(927);
    layer5_outputs(4978) <= layer4_outputs(3122);
    layer5_outputs(4979) <= (layer4_outputs(4870)) and not (layer4_outputs(4748));
    layer5_outputs(4980) <= not(layer4_outputs(2221));
    layer5_outputs(4981) <= (layer4_outputs(3966)) or (layer4_outputs(5086));
    layer5_outputs(4982) <= (layer4_outputs(1562)) and not (layer4_outputs(386));
    layer5_outputs(4983) <= layer4_outputs(397);
    layer5_outputs(4984) <= layer4_outputs(4071);
    layer5_outputs(4985) <= (layer4_outputs(1978)) and (layer4_outputs(355));
    layer5_outputs(4986) <= (layer4_outputs(1748)) or (layer4_outputs(4400));
    layer5_outputs(4987) <= (layer4_outputs(4990)) and not (layer4_outputs(5039));
    layer5_outputs(4988) <= not((layer4_outputs(616)) or (layer4_outputs(2001)));
    layer5_outputs(4989) <= (layer4_outputs(1238)) and not (layer4_outputs(565));
    layer5_outputs(4990) <= not(layer4_outputs(4728));
    layer5_outputs(4991) <= not((layer4_outputs(484)) or (layer4_outputs(3129)));
    layer5_outputs(4992) <= not(layer4_outputs(2904));
    layer5_outputs(4993) <= not((layer4_outputs(1299)) and (layer4_outputs(3594)));
    layer5_outputs(4994) <= layer4_outputs(4053);
    layer5_outputs(4995) <= layer4_outputs(1661);
    layer5_outputs(4996) <= not(layer4_outputs(3526));
    layer5_outputs(4997) <= not(layer4_outputs(1175));
    layer5_outputs(4998) <= not(layer4_outputs(4719)) or (layer4_outputs(5045));
    layer5_outputs(4999) <= not(layer4_outputs(1272));
    layer5_outputs(5000) <= '0';
    layer5_outputs(5001) <= not(layer4_outputs(1272));
    layer5_outputs(5002) <= (layer4_outputs(3566)) and not (layer4_outputs(2872));
    layer5_outputs(5003) <= (layer4_outputs(3667)) or (layer4_outputs(536));
    layer5_outputs(5004) <= layer4_outputs(608);
    layer5_outputs(5005) <= (layer4_outputs(5024)) xor (layer4_outputs(536));
    layer5_outputs(5006) <= (layer4_outputs(223)) and (layer4_outputs(996));
    layer5_outputs(5007) <= layer4_outputs(1176);
    layer5_outputs(5008) <= layer4_outputs(3872);
    layer5_outputs(5009) <= (layer4_outputs(540)) and (layer4_outputs(1764));
    layer5_outputs(5010) <= not((layer4_outputs(133)) and (layer4_outputs(4845)));
    layer5_outputs(5011) <= layer4_outputs(1790);
    layer5_outputs(5012) <= not((layer4_outputs(4723)) or (layer4_outputs(3792)));
    layer5_outputs(5013) <= layer4_outputs(1065);
    layer5_outputs(5014) <= '0';
    layer5_outputs(5015) <= (layer4_outputs(838)) and not (layer4_outputs(3174));
    layer5_outputs(5016) <= not((layer4_outputs(2258)) xor (layer4_outputs(2199)));
    layer5_outputs(5017) <= not((layer4_outputs(4889)) and (layer4_outputs(1233)));
    layer5_outputs(5018) <= (layer4_outputs(634)) and not (layer4_outputs(2989));
    layer5_outputs(5019) <= (layer4_outputs(4377)) and (layer4_outputs(1087));
    layer5_outputs(5020) <= layer4_outputs(1673);
    layer5_outputs(5021) <= (layer4_outputs(1278)) and not (layer4_outputs(3733));
    layer5_outputs(5022) <= layer4_outputs(324);
    layer5_outputs(5023) <= not(layer4_outputs(4772));
    layer5_outputs(5024) <= (layer4_outputs(1777)) and (layer4_outputs(3616));
    layer5_outputs(5025) <= (layer4_outputs(4390)) xor (layer4_outputs(3404));
    layer5_outputs(5026) <= layer4_outputs(580);
    layer5_outputs(5027) <= (layer4_outputs(4525)) and not (layer4_outputs(3380));
    layer5_outputs(5028) <= not(layer4_outputs(2489)) or (layer4_outputs(3375));
    layer5_outputs(5029) <= not(layer4_outputs(4138));
    layer5_outputs(5030) <= '1';
    layer5_outputs(5031) <= (layer4_outputs(1473)) and not (layer4_outputs(4745));
    layer5_outputs(5032) <= not((layer4_outputs(3222)) and (layer4_outputs(2156)));
    layer5_outputs(5033) <= layer4_outputs(2081);
    layer5_outputs(5034) <= (layer4_outputs(2545)) and (layer4_outputs(1623));
    layer5_outputs(5035) <= '1';
    layer5_outputs(5036) <= '1';
    layer5_outputs(5037) <= (layer4_outputs(681)) and not (layer4_outputs(2406));
    layer5_outputs(5038) <= '1';
    layer5_outputs(5039) <= (layer4_outputs(3041)) or (layer4_outputs(344));
    layer5_outputs(5040) <= not(layer4_outputs(5116)) or (layer4_outputs(3353));
    layer5_outputs(5041) <= (layer4_outputs(4078)) and not (layer4_outputs(4822));
    layer5_outputs(5042) <= not((layer4_outputs(3002)) and (layer4_outputs(1763)));
    layer5_outputs(5043) <= not((layer4_outputs(859)) and (layer4_outputs(3757)));
    layer5_outputs(5044) <= not((layer4_outputs(4008)) and (layer4_outputs(862)));
    layer5_outputs(5045) <= layer4_outputs(798);
    layer5_outputs(5046) <= (layer4_outputs(1859)) and not (layer4_outputs(10));
    layer5_outputs(5047) <= not(layer4_outputs(3866));
    layer5_outputs(5048) <= (layer4_outputs(1630)) and not (layer4_outputs(624));
    layer5_outputs(5049) <= not(layer4_outputs(4477));
    layer5_outputs(5050) <= not(layer4_outputs(4226));
    layer5_outputs(5051) <= not(layer4_outputs(2975)) or (layer4_outputs(2165));
    layer5_outputs(5052) <= (layer4_outputs(2006)) and (layer4_outputs(1598));
    layer5_outputs(5053) <= not((layer4_outputs(2929)) and (layer4_outputs(2138)));
    layer5_outputs(5054) <= not(layer4_outputs(4985)) or (layer4_outputs(382));
    layer5_outputs(5055) <= not((layer4_outputs(4800)) or (layer4_outputs(773)));
    layer5_outputs(5056) <= not(layer4_outputs(321));
    layer5_outputs(5057) <= '1';
    layer5_outputs(5058) <= layer4_outputs(3778);
    layer5_outputs(5059) <= not(layer4_outputs(4111));
    layer5_outputs(5060) <= (layer4_outputs(4833)) and (layer4_outputs(622));
    layer5_outputs(5061) <= (layer4_outputs(736)) and (layer4_outputs(7));
    layer5_outputs(5062) <= '0';
    layer5_outputs(5063) <= not(layer4_outputs(1829)) or (layer4_outputs(4470));
    layer5_outputs(5064) <= layer4_outputs(1109);
    layer5_outputs(5065) <= layer4_outputs(2877);
    layer5_outputs(5066) <= not(layer4_outputs(2795)) or (layer4_outputs(3581));
    layer5_outputs(5067) <= '1';
    layer5_outputs(5068) <= not(layer4_outputs(4734));
    layer5_outputs(5069) <= not((layer4_outputs(1734)) or (layer4_outputs(1255)));
    layer5_outputs(5070) <= not(layer4_outputs(2744));
    layer5_outputs(5071) <= not((layer4_outputs(2379)) or (layer4_outputs(759)));
    layer5_outputs(5072) <= not((layer4_outputs(3970)) xor (layer4_outputs(2542)));
    layer5_outputs(5073) <= (layer4_outputs(2066)) and (layer4_outputs(2690));
    layer5_outputs(5074) <= not((layer4_outputs(3460)) and (layer4_outputs(3613)));
    layer5_outputs(5075) <= not((layer4_outputs(4082)) xor (layer4_outputs(45)));
    layer5_outputs(5076) <= (layer4_outputs(183)) and not (layer4_outputs(753));
    layer5_outputs(5077) <= not(layer4_outputs(201)) or (layer4_outputs(2790));
    layer5_outputs(5078) <= (layer4_outputs(2592)) and not (layer4_outputs(2616));
    layer5_outputs(5079) <= not((layer4_outputs(1249)) and (layer4_outputs(2852)));
    layer5_outputs(5080) <= not(layer4_outputs(4704)) or (layer4_outputs(3247));
    layer5_outputs(5081) <= not(layer4_outputs(603));
    layer5_outputs(5082) <= (layer4_outputs(2724)) and not (layer4_outputs(2939));
    layer5_outputs(5083) <= (layer4_outputs(3884)) and not (layer4_outputs(1844));
    layer5_outputs(5084) <= layer4_outputs(332);
    layer5_outputs(5085) <= (layer4_outputs(4599)) and (layer4_outputs(1421));
    layer5_outputs(5086) <= not((layer4_outputs(4128)) or (layer4_outputs(1520)));
    layer5_outputs(5087) <= (layer4_outputs(4646)) and not (layer4_outputs(542));
    layer5_outputs(5088) <= not(layer4_outputs(4494)) or (layer4_outputs(183));
    layer5_outputs(5089) <= not(layer4_outputs(3394)) or (layer4_outputs(3842));
    layer5_outputs(5090) <= layer4_outputs(1912);
    layer5_outputs(5091) <= (layer4_outputs(3557)) and not (layer4_outputs(2268));
    layer5_outputs(5092) <= (layer4_outputs(2357)) and not (layer4_outputs(4533));
    layer5_outputs(5093) <= (layer4_outputs(885)) and not (layer4_outputs(1576));
    layer5_outputs(5094) <= layer4_outputs(1024);
    layer5_outputs(5095) <= (layer4_outputs(3633)) and (layer4_outputs(1977));
    layer5_outputs(5096) <= not(layer4_outputs(2459));
    layer5_outputs(5097) <= not(layer4_outputs(4257));
    layer5_outputs(5098) <= layer4_outputs(3526);
    layer5_outputs(5099) <= layer4_outputs(4006);
    layer5_outputs(5100) <= layer4_outputs(3050);
    layer5_outputs(5101) <= layer4_outputs(883);
    layer5_outputs(5102) <= not(layer4_outputs(4206)) or (layer4_outputs(658));
    layer5_outputs(5103) <= (layer4_outputs(4725)) and not (layer4_outputs(3217));
    layer5_outputs(5104) <= (layer4_outputs(1746)) and not (layer4_outputs(4562));
    layer5_outputs(5105) <= '1';
    layer5_outputs(5106) <= (layer4_outputs(4138)) or (layer4_outputs(727));
    layer5_outputs(5107) <= layer4_outputs(1331);
    layer5_outputs(5108) <= (layer4_outputs(359)) and (layer4_outputs(1515));
    layer5_outputs(5109) <= layer4_outputs(3069);
    layer5_outputs(5110) <= (layer4_outputs(974)) and (layer4_outputs(2817));
    layer5_outputs(5111) <= not(layer4_outputs(3933)) or (layer4_outputs(4044));
    layer5_outputs(5112) <= not(layer4_outputs(1755)) or (layer4_outputs(2208));
    layer5_outputs(5113) <= not(layer4_outputs(672)) or (layer4_outputs(2548));
    layer5_outputs(5114) <= not(layer4_outputs(583)) or (layer4_outputs(1204));
    layer5_outputs(5115) <= (layer4_outputs(320)) or (layer4_outputs(3831));
    layer5_outputs(5116) <= not((layer4_outputs(3788)) and (layer4_outputs(3619)));
    layer5_outputs(5117) <= (layer4_outputs(91)) and not (layer4_outputs(2160));
    layer5_outputs(5118) <= (layer4_outputs(4696)) and not (layer4_outputs(1375));
    layer5_outputs(5119) <= not(layer4_outputs(3946));
    layer6_outputs(0) <= not((layer5_outputs(4840)) and (layer5_outputs(1884)));
    layer6_outputs(1) <= '1';
    layer6_outputs(2) <= (layer5_outputs(5053)) xor (layer5_outputs(2966));
    layer6_outputs(3) <= '1';
    layer6_outputs(4) <= '1';
    layer6_outputs(5) <= layer5_outputs(1716);
    layer6_outputs(6) <= not(layer5_outputs(1021));
    layer6_outputs(7) <= (layer5_outputs(1842)) and not (layer5_outputs(2965));
    layer6_outputs(8) <= layer5_outputs(3592);
    layer6_outputs(9) <= layer5_outputs(3099);
    layer6_outputs(10) <= not(layer5_outputs(1945));
    layer6_outputs(11) <= (layer5_outputs(2866)) or (layer5_outputs(2076));
    layer6_outputs(12) <= not(layer5_outputs(3265));
    layer6_outputs(13) <= not(layer5_outputs(1722));
    layer6_outputs(14) <= (layer5_outputs(1507)) and (layer5_outputs(993));
    layer6_outputs(15) <= not(layer5_outputs(2945));
    layer6_outputs(16) <= '0';
    layer6_outputs(17) <= not(layer5_outputs(3092));
    layer6_outputs(18) <= (layer5_outputs(1561)) and not (layer5_outputs(2156));
    layer6_outputs(19) <= not(layer5_outputs(1871));
    layer6_outputs(20) <= not((layer5_outputs(172)) or (layer5_outputs(421)));
    layer6_outputs(21) <= not((layer5_outputs(1822)) or (layer5_outputs(4343)));
    layer6_outputs(22) <= '0';
    layer6_outputs(23) <= layer5_outputs(4475);
    layer6_outputs(24) <= not(layer5_outputs(4733));
    layer6_outputs(25) <= not(layer5_outputs(4349));
    layer6_outputs(26) <= not(layer5_outputs(5081));
    layer6_outputs(27) <= not(layer5_outputs(1670));
    layer6_outputs(28) <= not((layer5_outputs(2586)) and (layer5_outputs(2936)));
    layer6_outputs(29) <= not(layer5_outputs(1620));
    layer6_outputs(30) <= not(layer5_outputs(2822));
    layer6_outputs(31) <= layer5_outputs(577);
    layer6_outputs(32) <= layer5_outputs(965);
    layer6_outputs(33) <= (layer5_outputs(695)) or (layer5_outputs(4433));
    layer6_outputs(34) <= not(layer5_outputs(3393));
    layer6_outputs(35) <= layer5_outputs(3166);
    layer6_outputs(36) <= (layer5_outputs(1178)) and not (layer5_outputs(2639));
    layer6_outputs(37) <= (layer5_outputs(1773)) and (layer5_outputs(725));
    layer6_outputs(38) <= layer5_outputs(4094);
    layer6_outputs(39) <= (layer5_outputs(4697)) xor (layer5_outputs(3178));
    layer6_outputs(40) <= (layer5_outputs(3674)) and not (layer5_outputs(4748));
    layer6_outputs(41) <= layer5_outputs(4752);
    layer6_outputs(42) <= '1';
    layer6_outputs(43) <= (layer5_outputs(2812)) and not (layer5_outputs(1079));
    layer6_outputs(44) <= layer5_outputs(2878);
    layer6_outputs(45) <= not(layer5_outputs(3422));
    layer6_outputs(46) <= not(layer5_outputs(3116));
    layer6_outputs(47) <= layer5_outputs(73);
    layer6_outputs(48) <= not(layer5_outputs(251));
    layer6_outputs(49) <= not(layer5_outputs(2109)) or (layer5_outputs(3999));
    layer6_outputs(50) <= not(layer5_outputs(3535));
    layer6_outputs(51) <= not(layer5_outputs(510));
    layer6_outputs(52) <= not(layer5_outputs(3006));
    layer6_outputs(53) <= not((layer5_outputs(3427)) or (layer5_outputs(4600)));
    layer6_outputs(54) <= not((layer5_outputs(4736)) xor (layer5_outputs(3844)));
    layer6_outputs(55) <= (layer5_outputs(1322)) or (layer5_outputs(713));
    layer6_outputs(56) <= (layer5_outputs(3699)) and not (layer5_outputs(1635));
    layer6_outputs(57) <= not(layer5_outputs(2318));
    layer6_outputs(58) <= layer5_outputs(3353);
    layer6_outputs(59) <= not(layer5_outputs(1624)) or (layer5_outputs(4442));
    layer6_outputs(60) <= not(layer5_outputs(1144));
    layer6_outputs(61) <= not(layer5_outputs(782));
    layer6_outputs(62) <= not(layer5_outputs(1674));
    layer6_outputs(63) <= layer5_outputs(2271);
    layer6_outputs(64) <= (layer5_outputs(2123)) xor (layer5_outputs(4521));
    layer6_outputs(65) <= (layer5_outputs(452)) and not (layer5_outputs(216));
    layer6_outputs(66) <= not(layer5_outputs(4561));
    layer6_outputs(67) <= not((layer5_outputs(2800)) xor (layer5_outputs(1153)));
    layer6_outputs(68) <= not(layer5_outputs(4044));
    layer6_outputs(69) <= (layer5_outputs(4551)) or (layer5_outputs(2148));
    layer6_outputs(70) <= layer5_outputs(1380);
    layer6_outputs(71) <= (layer5_outputs(2556)) and (layer5_outputs(3929));
    layer6_outputs(72) <= not(layer5_outputs(3084)) or (layer5_outputs(530));
    layer6_outputs(73) <= '1';
    layer6_outputs(74) <= (layer5_outputs(3560)) and not (layer5_outputs(1140));
    layer6_outputs(75) <= (layer5_outputs(4823)) and not (layer5_outputs(3239));
    layer6_outputs(76) <= '1';
    layer6_outputs(77) <= not((layer5_outputs(2132)) or (layer5_outputs(1012)));
    layer6_outputs(78) <= not((layer5_outputs(2926)) or (layer5_outputs(2636)));
    layer6_outputs(79) <= (layer5_outputs(206)) and not (layer5_outputs(3759));
    layer6_outputs(80) <= not((layer5_outputs(1577)) or (layer5_outputs(1460)));
    layer6_outputs(81) <= not(layer5_outputs(4747)) or (layer5_outputs(1417));
    layer6_outputs(82) <= layer5_outputs(3309);
    layer6_outputs(83) <= not(layer5_outputs(4421)) or (layer5_outputs(2835));
    layer6_outputs(84) <= not((layer5_outputs(4159)) xor (layer5_outputs(3148)));
    layer6_outputs(85) <= not(layer5_outputs(3878));
    layer6_outputs(86) <= layer5_outputs(1299);
    layer6_outputs(87) <= (layer5_outputs(84)) or (layer5_outputs(4967));
    layer6_outputs(88) <= not((layer5_outputs(3224)) xor (layer5_outputs(2013)));
    layer6_outputs(89) <= (layer5_outputs(386)) and not (layer5_outputs(2389));
    layer6_outputs(90) <= not(layer5_outputs(2253));
    layer6_outputs(91) <= not(layer5_outputs(1195));
    layer6_outputs(92) <= not(layer5_outputs(2442)) or (layer5_outputs(4701));
    layer6_outputs(93) <= not(layer5_outputs(3179));
    layer6_outputs(94) <= layer5_outputs(4938);
    layer6_outputs(95) <= layer5_outputs(2469);
    layer6_outputs(96) <= (layer5_outputs(2279)) and (layer5_outputs(1225));
    layer6_outputs(97) <= not(layer5_outputs(981));
    layer6_outputs(98) <= not(layer5_outputs(469));
    layer6_outputs(99) <= not(layer5_outputs(1371));
    layer6_outputs(100) <= not((layer5_outputs(3653)) xor (layer5_outputs(4979)));
    layer6_outputs(101) <= not((layer5_outputs(2315)) and (layer5_outputs(1154)));
    layer6_outputs(102) <= (layer5_outputs(2252)) and not (layer5_outputs(190));
    layer6_outputs(103) <= '1';
    layer6_outputs(104) <= (layer5_outputs(149)) and (layer5_outputs(3004));
    layer6_outputs(105) <= (layer5_outputs(3213)) and not (layer5_outputs(4055));
    layer6_outputs(106) <= not(layer5_outputs(984)) or (layer5_outputs(3739));
    layer6_outputs(107) <= not(layer5_outputs(1459)) or (layer5_outputs(699));
    layer6_outputs(108) <= not((layer5_outputs(3523)) or (layer5_outputs(3143)));
    layer6_outputs(109) <= not(layer5_outputs(2418));
    layer6_outputs(110) <= layer5_outputs(3651);
    layer6_outputs(111) <= (layer5_outputs(161)) and not (layer5_outputs(1405));
    layer6_outputs(112) <= not(layer5_outputs(3331));
    layer6_outputs(113) <= not((layer5_outputs(633)) or (layer5_outputs(1453)));
    layer6_outputs(114) <= (layer5_outputs(1609)) or (layer5_outputs(2230));
    layer6_outputs(115) <= (layer5_outputs(1940)) and (layer5_outputs(2343));
    layer6_outputs(116) <= (layer5_outputs(2792)) and not (layer5_outputs(3458));
    layer6_outputs(117) <= (layer5_outputs(3004)) and not (layer5_outputs(372));
    layer6_outputs(118) <= (layer5_outputs(4429)) and not (layer5_outputs(4745));
    layer6_outputs(119) <= '0';
    layer6_outputs(120) <= (layer5_outputs(2887)) and not (layer5_outputs(3328));
    layer6_outputs(121) <= (layer5_outputs(4923)) or (layer5_outputs(3939));
    layer6_outputs(122) <= not((layer5_outputs(3310)) and (layer5_outputs(462)));
    layer6_outputs(123) <= (layer5_outputs(3635)) or (layer5_outputs(4101));
    layer6_outputs(124) <= (layer5_outputs(1566)) or (layer5_outputs(361));
    layer6_outputs(125) <= not((layer5_outputs(3016)) xor (layer5_outputs(4729)));
    layer6_outputs(126) <= not(layer5_outputs(1032));
    layer6_outputs(127) <= layer5_outputs(1303);
    layer6_outputs(128) <= not(layer5_outputs(4080));
    layer6_outputs(129) <= not(layer5_outputs(1801));
    layer6_outputs(130) <= not((layer5_outputs(1265)) or (layer5_outputs(1691)));
    layer6_outputs(131) <= (layer5_outputs(4833)) and not (layer5_outputs(2558));
    layer6_outputs(132) <= layer5_outputs(2177);
    layer6_outputs(133) <= (layer5_outputs(4628)) or (layer5_outputs(1408));
    layer6_outputs(134) <= layer5_outputs(700);
    layer6_outputs(135) <= not(layer5_outputs(836));
    layer6_outputs(136) <= not(layer5_outputs(2188)) or (layer5_outputs(5096));
    layer6_outputs(137) <= (layer5_outputs(574)) and (layer5_outputs(3082));
    layer6_outputs(138) <= not(layer5_outputs(2827));
    layer6_outputs(139) <= not(layer5_outputs(175));
    layer6_outputs(140) <= not(layer5_outputs(2282));
    layer6_outputs(141) <= layer5_outputs(94);
    layer6_outputs(142) <= not((layer5_outputs(3186)) xor (layer5_outputs(2431)));
    layer6_outputs(143) <= not((layer5_outputs(4117)) or (layer5_outputs(2988)));
    layer6_outputs(144) <= (layer5_outputs(3236)) and not (layer5_outputs(2084));
    layer6_outputs(145) <= (layer5_outputs(3942)) and not (layer5_outputs(4528));
    layer6_outputs(146) <= '1';
    layer6_outputs(147) <= not((layer5_outputs(2257)) and (layer5_outputs(2957)));
    layer6_outputs(148) <= layer5_outputs(714);
    layer6_outputs(149) <= layer5_outputs(2161);
    layer6_outputs(150) <= not(layer5_outputs(4582));
    layer6_outputs(151) <= layer5_outputs(2340);
    layer6_outputs(152) <= (layer5_outputs(1467)) and not (layer5_outputs(4275));
    layer6_outputs(153) <= layer5_outputs(2048);
    layer6_outputs(154) <= not(layer5_outputs(3032));
    layer6_outputs(155) <= layer5_outputs(557);
    layer6_outputs(156) <= not((layer5_outputs(2481)) xor (layer5_outputs(252)));
    layer6_outputs(157) <= layer5_outputs(2375);
    layer6_outputs(158) <= not(layer5_outputs(4347));
    layer6_outputs(159) <= (layer5_outputs(3816)) and not (layer5_outputs(1411));
    layer6_outputs(160) <= layer5_outputs(4119);
    layer6_outputs(161) <= not(layer5_outputs(876)) or (layer5_outputs(4061));
    layer6_outputs(162) <= (layer5_outputs(4471)) and not (layer5_outputs(2980));
    layer6_outputs(163) <= not(layer5_outputs(1663));
    layer6_outputs(164) <= '1';
    layer6_outputs(165) <= not(layer5_outputs(1252)) or (layer5_outputs(3757));
    layer6_outputs(166) <= not(layer5_outputs(4281));
    layer6_outputs(167) <= not(layer5_outputs(4160));
    layer6_outputs(168) <= not(layer5_outputs(2621));
    layer6_outputs(169) <= (layer5_outputs(2325)) and not (layer5_outputs(2898));
    layer6_outputs(170) <= not(layer5_outputs(2044));
    layer6_outputs(171) <= layer5_outputs(2498);
    layer6_outputs(172) <= not(layer5_outputs(1891)) or (layer5_outputs(446));
    layer6_outputs(173) <= not(layer5_outputs(2375));
    layer6_outputs(174) <= not(layer5_outputs(60));
    layer6_outputs(175) <= not(layer5_outputs(3974));
    layer6_outputs(176) <= not(layer5_outputs(3284));
    layer6_outputs(177) <= layer5_outputs(1568);
    layer6_outputs(178) <= not(layer5_outputs(3897));
    layer6_outputs(179) <= (layer5_outputs(3508)) and not (layer5_outputs(4520));
    layer6_outputs(180) <= not(layer5_outputs(3139)) or (layer5_outputs(2954));
    layer6_outputs(181) <= not((layer5_outputs(168)) xor (layer5_outputs(1158)));
    layer6_outputs(182) <= (layer5_outputs(2334)) or (layer5_outputs(2747));
    layer6_outputs(183) <= (layer5_outputs(679)) or (layer5_outputs(4952));
    layer6_outputs(184) <= (layer5_outputs(2967)) and not (layer5_outputs(1726));
    layer6_outputs(185) <= layer5_outputs(2446);
    layer6_outputs(186) <= not(layer5_outputs(793));
    layer6_outputs(187) <= '1';
    layer6_outputs(188) <= layer5_outputs(3095);
    layer6_outputs(189) <= not(layer5_outputs(1842));
    layer6_outputs(190) <= not(layer5_outputs(2303)) or (layer5_outputs(279));
    layer6_outputs(191) <= not((layer5_outputs(1838)) xor (layer5_outputs(2631)));
    layer6_outputs(192) <= not(layer5_outputs(3463));
    layer6_outputs(193) <= layer5_outputs(2183);
    layer6_outputs(194) <= not((layer5_outputs(3260)) and (layer5_outputs(3013)));
    layer6_outputs(195) <= (layer5_outputs(2461)) xor (layer5_outputs(1543));
    layer6_outputs(196) <= not(layer5_outputs(1181));
    layer6_outputs(197) <= not(layer5_outputs(2070));
    layer6_outputs(198) <= not(layer5_outputs(4836)) or (layer5_outputs(2616));
    layer6_outputs(199) <= (layer5_outputs(1348)) or (layer5_outputs(2756));
    layer6_outputs(200) <= (layer5_outputs(4329)) or (layer5_outputs(4866));
    layer6_outputs(201) <= layer5_outputs(1938);
    layer6_outputs(202) <= not(layer5_outputs(1275)) or (layer5_outputs(2784));
    layer6_outputs(203) <= layer5_outputs(1701);
    layer6_outputs(204) <= not(layer5_outputs(4455)) or (layer5_outputs(3992));
    layer6_outputs(205) <= layer5_outputs(3209);
    layer6_outputs(206) <= not(layer5_outputs(151));
    layer6_outputs(207) <= not((layer5_outputs(3144)) or (layer5_outputs(1887)));
    layer6_outputs(208) <= '0';
    layer6_outputs(209) <= (layer5_outputs(2760)) or (layer5_outputs(3012));
    layer6_outputs(210) <= not(layer5_outputs(290)) or (layer5_outputs(4273));
    layer6_outputs(211) <= not((layer5_outputs(2521)) or (layer5_outputs(239)));
    layer6_outputs(212) <= not(layer5_outputs(1991));
    layer6_outputs(213) <= (layer5_outputs(3357)) and not (layer5_outputs(4142));
    layer6_outputs(214) <= not(layer5_outputs(4752));
    layer6_outputs(215) <= (layer5_outputs(1321)) or (layer5_outputs(4630));
    layer6_outputs(216) <= not(layer5_outputs(3600));
    layer6_outputs(217) <= '1';
    layer6_outputs(218) <= layer5_outputs(1337);
    layer6_outputs(219) <= layer5_outputs(1872);
    layer6_outputs(220) <= not(layer5_outputs(4216));
    layer6_outputs(221) <= (layer5_outputs(2497)) xor (layer5_outputs(692));
    layer6_outputs(222) <= layer5_outputs(2075);
    layer6_outputs(223) <= layer5_outputs(440);
    layer6_outputs(224) <= not(layer5_outputs(1165));
    layer6_outputs(225) <= not((layer5_outputs(3110)) or (layer5_outputs(582)));
    layer6_outputs(226) <= layer5_outputs(632);
    layer6_outputs(227) <= layer5_outputs(927);
    layer6_outputs(228) <= not(layer5_outputs(4285));
    layer6_outputs(229) <= (layer5_outputs(1851)) and (layer5_outputs(2973));
    layer6_outputs(230) <= not(layer5_outputs(2045));
    layer6_outputs(231) <= not(layer5_outputs(372));
    layer6_outputs(232) <= layer5_outputs(1743);
    layer6_outputs(233) <= layer5_outputs(4411);
    layer6_outputs(234) <= layer5_outputs(3127);
    layer6_outputs(235) <= '1';
    layer6_outputs(236) <= (layer5_outputs(4432)) or (layer5_outputs(3501));
    layer6_outputs(237) <= layer5_outputs(1741);
    layer6_outputs(238) <= (layer5_outputs(3473)) or (layer5_outputs(768));
    layer6_outputs(239) <= (layer5_outputs(1876)) and not (layer5_outputs(3475));
    layer6_outputs(240) <= not((layer5_outputs(4394)) xor (layer5_outputs(4990)));
    layer6_outputs(241) <= not(layer5_outputs(4235)) or (layer5_outputs(957));
    layer6_outputs(242) <= layer5_outputs(4322);
    layer6_outputs(243) <= not(layer5_outputs(3530)) or (layer5_outputs(249));
    layer6_outputs(244) <= (layer5_outputs(4268)) or (layer5_outputs(3768));
    layer6_outputs(245) <= not((layer5_outputs(3957)) or (layer5_outputs(1087)));
    layer6_outputs(246) <= not((layer5_outputs(3876)) or (layer5_outputs(229)));
    layer6_outputs(247) <= not(layer5_outputs(1390)) or (layer5_outputs(2119));
    layer6_outputs(248) <= (layer5_outputs(1413)) xor (layer5_outputs(2238));
    layer6_outputs(249) <= '0';
    layer6_outputs(250) <= not(layer5_outputs(2781)) or (layer5_outputs(2691));
    layer6_outputs(251) <= (layer5_outputs(3807)) xor (layer5_outputs(1906));
    layer6_outputs(252) <= not(layer5_outputs(1537)) or (layer5_outputs(1362));
    layer6_outputs(253) <= not((layer5_outputs(4321)) or (layer5_outputs(4636)));
    layer6_outputs(254) <= not((layer5_outputs(1495)) xor (layer5_outputs(60)));
    layer6_outputs(255) <= not(layer5_outputs(762)) or (layer5_outputs(382));
    layer6_outputs(256) <= (layer5_outputs(241)) and not (layer5_outputs(3445));
    layer6_outputs(257) <= layer5_outputs(1761);
    layer6_outputs(258) <= not(layer5_outputs(2868)) or (layer5_outputs(1891));
    layer6_outputs(259) <= not(layer5_outputs(3853)) or (layer5_outputs(1063));
    layer6_outputs(260) <= not((layer5_outputs(3054)) or (layer5_outputs(4918)));
    layer6_outputs(261) <= layer5_outputs(3581);
    layer6_outputs(262) <= layer5_outputs(3940);
    layer6_outputs(263) <= not(layer5_outputs(1977));
    layer6_outputs(264) <= layer5_outputs(3822);
    layer6_outputs(265) <= not((layer5_outputs(1648)) or (layer5_outputs(2190)));
    layer6_outputs(266) <= (layer5_outputs(751)) and (layer5_outputs(2565));
    layer6_outputs(267) <= (layer5_outputs(780)) and (layer5_outputs(1988));
    layer6_outputs(268) <= (layer5_outputs(2836)) and not (layer5_outputs(4455));
    layer6_outputs(269) <= layer5_outputs(1719);
    layer6_outputs(270) <= '0';
    layer6_outputs(271) <= (layer5_outputs(4857)) and not (layer5_outputs(790));
    layer6_outputs(272) <= layer5_outputs(299);
    layer6_outputs(273) <= layer5_outputs(2633);
    layer6_outputs(274) <= (layer5_outputs(2811)) and not (layer5_outputs(4639));
    layer6_outputs(275) <= not(layer5_outputs(5119)) or (layer5_outputs(4368));
    layer6_outputs(276) <= not(layer5_outputs(4213)) or (layer5_outputs(3457));
    layer6_outputs(277) <= not((layer5_outputs(3925)) and (layer5_outputs(3062)));
    layer6_outputs(278) <= (layer5_outputs(5097)) and not (layer5_outputs(3576));
    layer6_outputs(279) <= not(layer5_outputs(2367)) or (layer5_outputs(1142));
    layer6_outputs(280) <= layer5_outputs(1735);
    layer6_outputs(281) <= not(layer5_outputs(2655)) or (layer5_outputs(1435));
    layer6_outputs(282) <= layer5_outputs(692);
    layer6_outputs(283) <= (layer5_outputs(3421)) or (layer5_outputs(1447));
    layer6_outputs(284) <= (layer5_outputs(2733)) and (layer5_outputs(3428));
    layer6_outputs(285) <= not(layer5_outputs(3105));
    layer6_outputs(286) <= not(layer5_outputs(1382)) or (layer5_outputs(1696));
    layer6_outputs(287) <= '1';
    layer6_outputs(288) <= not((layer5_outputs(3605)) or (layer5_outputs(4002)));
    layer6_outputs(289) <= (layer5_outputs(2883)) and not (layer5_outputs(2278));
    layer6_outputs(290) <= not(layer5_outputs(540)) or (layer5_outputs(1796));
    layer6_outputs(291) <= layer5_outputs(4124);
    layer6_outputs(292) <= not(layer5_outputs(476));
    layer6_outputs(293) <= (layer5_outputs(3201)) and (layer5_outputs(1590));
    layer6_outputs(294) <= layer5_outputs(5011);
    layer6_outputs(295) <= (layer5_outputs(2067)) xor (layer5_outputs(4862));
    layer6_outputs(296) <= (layer5_outputs(4744)) and not (layer5_outputs(3697));
    layer6_outputs(297) <= layer5_outputs(2644);
    layer6_outputs(298) <= not((layer5_outputs(1859)) xor (layer5_outputs(847)));
    layer6_outputs(299) <= not((layer5_outputs(5067)) or (layer5_outputs(3558)));
    layer6_outputs(300) <= not(layer5_outputs(4232));
    layer6_outputs(301) <= not(layer5_outputs(2699));
    layer6_outputs(302) <= not(layer5_outputs(4705));
    layer6_outputs(303) <= (layer5_outputs(2786)) and not (layer5_outputs(4417));
    layer6_outputs(304) <= not((layer5_outputs(20)) xor (layer5_outputs(3825)));
    layer6_outputs(305) <= layer5_outputs(2046);
    layer6_outputs(306) <= not(layer5_outputs(3711));
    layer6_outputs(307) <= layer5_outputs(2723);
    layer6_outputs(308) <= '1';
    layer6_outputs(309) <= not(layer5_outputs(2460)) or (layer5_outputs(3238));
    layer6_outputs(310) <= not((layer5_outputs(2390)) and (layer5_outputs(309)));
    layer6_outputs(311) <= (layer5_outputs(1052)) or (layer5_outputs(802));
    layer6_outputs(312) <= not(layer5_outputs(1008));
    layer6_outputs(313) <= layer5_outputs(3814);
    layer6_outputs(314) <= layer5_outputs(3218);
    layer6_outputs(315) <= not(layer5_outputs(2790));
    layer6_outputs(316) <= not(layer5_outputs(3136)) or (layer5_outputs(1916));
    layer6_outputs(317) <= not(layer5_outputs(3336));
    layer6_outputs(318) <= not(layer5_outputs(1612));
    layer6_outputs(319) <= not(layer5_outputs(657)) or (layer5_outputs(3289));
    layer6_outputs(320) <= (layer5_outputs(2998)) and (layer5_outputs(3740));
    layer6_outputs(321) <= layer5_outputs(861);
    layer6_outputs(322) <= not(layer5_outputs(4889)) or (layer5_outputs(3945));
    layer6_outputs(323) <= not(layer5_outputs(1946));
    layer6_outputs(324) <= not((layer5_outputs(3140)) and (layer5_outputs(3044)));
    layer6_outputs(325) <= (layer5_outputs(39)) and (layer5_outputs(4186));
    layer6_outputs(326) <= not(layer5_outputs(4707)) or (layer5_outputs(1952));
    layer6_outputs(327) <= layer5_outputs(4236);
    layer6_outputs(328) <= layer5_outputs(146);
    layer6_outputs(329) <= (layer5_outputs(4435)) or (layer5_outputs(2344));
    layer6_outputs(330) <= layer5_outputs(65);
    layer6_outputs(331) <= not(layer5_outputs(3066));
    layer6_outputs(332) <= not(layer5_outputs(226));
    layer6_outputs(333) <= (layer5_outputs(139)) and not (layer5_outputs(1359));
    layer6_outputs(334) <= not(layer5_outputs(4152));
    layer6_outputs(335) <= not((layer5_outputs(74)) xor (layer5_outputs(3614)));
    layer6_outputs(336) <= not(layer5_outputs(1904)) or (layer5_outputs(2505));
    layer6_outputs(337) <= not(layer5_outputs(3038)) or (layer5_outputs(3022));
    layer6_outputs(338) <= not(layer5_outputs(1290));
    layer6_outputs(339) <= not(layer5_outputs(2055)) or (layer5_outputs(1504));
    layer6_outputs(340) <= not(layer5_outputs(235));
    layer6_outputs(341) <= (layer5_outputs(4608)) xor (layer5_outputs(705));
    layer6_outputs(342) <= layer5_outputs(2083);
    layer6_outputs(343) <= layer5_outputs(521);
    layer6_outputs(344) <= not(layer5_outputs(1893));
    layer6_outputs(345) <= layer5_outputs(4462);
    layer6_outputs(346) <= not(layer5_outputs(4230));
    layer6_outputs(347) <= not(layer5_outputs(4954));
    layer6_outputs(348) <= (layer5_outputs(1713)) and not (layer5_outputs(3404));
    layer6_outputs(349) <= not((layer5_outputs(909)) and (layer5_outputs(3956)));
    layer6_outputs(350) <= (layer5_outputs(2221)) and (layer5_outputs(2885));
    layer6_outputs(351) <= not(layer5_outputs(1006));
    layer6_outputs(352) <= not(layer5_outputs(2474));
    layer6_outputs(353) <= layer5_outputs(4027);
    layer6_outputs(354) <= layer5_outputs(4062);
    layer6_outputs(355) <= not(layer5_outputs(2992)) or (layer5_outputs(3256));
    layer6_outputs(356) <= not((layer5_outputs(2355)) or (layer5_outputs(4800)));
    layer6_outputs(357) <= not(layer5_outputs(3303)) or (layer5_outputs(1783));
    layer6_outputs(358) <= not(layer5_outputs(4901));
    layer6_outputs(359) <= '1';
    layer6_outputs(360) <= not((layer5_outputs(4133)) and (layer5_outputs(4428)));
    layer6_outputs(361) <= not(layer5_outputs(2799));
    layer6_outputs(362) <= '0';
    layer6_outputs(363) <= (layer5_outputs(3071)) and not (layer5_outputs(3740));
    layer6_outputs(364) <= (layer5_outputs(4223)) and (layer5_outputs(845));
    layer6_outputs(365) <= not((layer5_outputs(3272)) xor (layer5_outputs(148)));
    layer6_outputs(366) <= not(layer5_outputs(2088));
    layer6_outputs(367) <= layer5_outputs(1824);
    layer6_outputs(368) <= not(layer5_outputs(4643));
    layer6_outputs(369) <= (layer5_outputs(314)) and not (layer5_outputs(2894));
    layer6_outputs(370) <= layer5_outputs(3245);
    layer6_outputs(371) <= not(layer5_outputs(4271));
    layer6_outputs(372) <= layer5_outputs(1217);
    layer6_outputs(373) <= layer5_outputs(4810);
    layer6_outputs(374) <= not(layer5_outputs(1812)) or (layer5_outputs(4312));
    layer6_outputs(375) <= layer5_outputs(4677);
    layer6_outputs(376) <= not((layer5_outputs(2702)) xor (layer5_outputs(571)));
    layer6_outputs(377) <= (layer5_outputs(4624)) and not (layer5_outputs(117));
    layer6_outputs(378) <= layer5_outputs(688);
    layer6_outputs(379) <= not((layer5_outputs(3011)) and (layer5_outputs(408)));
    layer6_outputs(380) <= not((layer5_outputs(4602)) and (layer5_outputs(3734)));
    layer6_outputs(381) <= layer5_outputs(548);
    layer6_outputs(382) <= not(layer5_outputs(4881));
    layer6_outputs(383) <= not(layer5_outputs(3304));
    layer6_outputs(384) <= (layer5_outputs(4751)) and (layer5_outputs(2815));
    layer6_outputs(385) <= not((layer5_outputs(5032)) or (layer5_outputs(2540)));
    layer6_outputs(386) <= (layer5_outputs(2779)) and (layer5_outputs(5069));
    layer6_outputs(387) <= not(layer5_outputs(2608));
    layer6_outputs(388) <= layer5_outputs(3978);
    layer6_outputs(389) <= layer5_outputs(2439);
    layer6_outputs(390) <= not(layer5_outputs(3655));
    layer6_outputs(391) <= not(layer5_outputs(4238));
    layer6_outputs(392) <= layer5_outputs(4018);
    layer6_outputs(393) <= not((layer5_outputs(2574)) or (layer5_outputs(4388)));
    layer6_outputs(394) <= not(layer5_outputs(2403)) or (layer5_outputs(2186));
    layer6_outputs(395) <= not((layer5_outputs(1464)) or (layer5_outputs(3587)));
    layer6_outputs(396) <= not((layer5_outputs(2110)) xor (layer5_outputs(4649)));
    layer6_outputs(397) <= layer5_outputs(606);
    layer6_outputs(398) <= not((layer5_outputs(1430)) xor (layer5_outputs(4939)));
    layer6_outputs(399) <= not(layer5_outputs(2139)) or (layer5_outputs(2210));
    layer6_outputs(400) <= layer5_outputs(1923);
    layer6_outputs(401) <= not((layer5_outputs(4356)) or (layer5_outputs(3193)));
    layer6_outputs(402) <= not(layer5_outputs(2127)) or (layer5_outputs(1594));
    layer6_outputs(403) <= not(layer5_outputs(2106));
    layer6_outputs(404) <= (layer5_outputs(4081)) and (layer5_outputs(32));
    layer6_outputs(405) <= (layer5_outputs(3937)) or (layer5_outputs(2042));
    layer6_outputs(406) <= (layer5_outputs(3167)) and not (layer5_outputs(4841));
    layer6_outputs(407) <= not(layer5_outputs(4354));
    layer6_outputs(408) <= not(layer5_outputs(1397));
    layer6_outputs(409) <= not((layer5_outputs(1497)) or (layer5_outputs(1986)));
    layer6_outputs(410) <= not(layer5_outputs(1779)) or (layer5_outputs(2845));
    layer6_outputs(411) <= not(layer5_outputs(141));
    layer6_outputs(412) <= layer5_outputs(4366);
    layer6_outputs(413) <= '1';
    layer6_outputs(414) <= not(layer5_outputs(3680)) or (layer5_outputs(1971));
    layer6_outputs(415) <= layer5_outputs(308);
    layer6_outputs(416) <= (layer5_outputs(1811)) or (layer5_outputs(2567));
    layer6_outputs(417) <= not(layer5_outputs(2451)) or (layer5_outputs(1628));
    layer6_outputs(418) <= layer5_outputs(3567);
    layer6_outputs(419) <= not(layer5_outputs(2149));
    layer6_outputs(420) <= (layer5_outputs(4812)) and not (layer5_outputs(1913));
    layer6_outputs(421) <= not(layer5_outputs(4813));
    layer6_outputs(422) <= layer5_outputs(2057);
    layer6_outputs(423) <= layer5_outputs(917);
    layer6_outputs(424) <= (layer5_outputs(38)) and not (layer5_outputs(546));
    layer6_outputs(425) <= not(layer5_outputs(4703));
    layer6_outputs(426) <= (layer5_outputs(3093)) and not (layer5_outputs(4963));
    layer6_outputs(427) <= (layer5_outputs(28)) and (layer5_outputs(668));
    layer6_outputs(428) <= not((layer5_outputs(3721)) and (layer5_outputs(4554)));
    layer6_outputs(429) <= not(layer5_outputs(1511));
    layer6_outputs(430) <= not((layer5_outputs(2030)) xor (layer5_outputs(1996)));
    layer6_outputs(431) <= not((layer5_outputs(23)) and (layer5_outputs(2988)));
    layer6_outputs(432) <= not((layer5_outputs(1856)) xor (layer5_outputs(1594)));
    layer6_outputs(433) <= layer5_outputs(4199);
    layer6_outputs(434) <= not(layer5_outputs(1850));
    layer6_outputs(435) <= not(layer5_outputs(1209)) or (layer5_outputs(4803));
    layer6_outputs(436) <= (layer5_outputs(3671)) and (layer5_outputs(319));
    layer6_outputs(437) <= not(layer5_outputs(18));
    layer6_outputs(438) <= layer5_outputs(3407);
    layer6_outputs(439) <= layer5_outputs(94);
    layer6_outputs(440) <= (layer5_outputs(602)) and not (layer5_outputs(61));
    layer6_outputs(441) <= (layer5_outputs(2929)) and not (layer5_outputs(1651));
    layer6_outputs(442) <= not(layer5_outputs(2337)) or (layer5_outputs(4869));
    layer6_outputs(443) <= (layer5_outputs(2855)) and (layer5_outputs(266));
    layer6_outputs(444) <= layer5_outputs(1077);
    layer6_outputs(445) <= not(layer5_outputs(1295)) or (layer5_outputs(3364));
    layer6_outputs(446) <= not(layer5_outputs(4528));
    layer6_outputs(447) <= layer5_outputs(296);
    layer6_outputs(448) <= (layer5_outputs(378)) and (layer5_outputs(4450));
    layer6_outputs(449) <= not(layer5_outputs(384));
    layer6_outputs(450) <= not((layer5_outputs(828)) and (layer5_outputs(3663)));
    layer6_outputs(451) <= not(layer5_outputs(1772));
    layer6_outputs(452) <= not(layer5_outputs(4883));
    layer6_outputs(453) <= not(layer5_outputs(3232)) or (layer5_outputs(514));
    layer6_outputs(454) <= (layer5_outputs(3805)) xor (layer5_outputs(340));
    layer6_outputs(455) <= not(layer5_outputs(1548)) or (layer5_outputs(1089));
    layer6_outputs(456) <= layer5_outputs(1338);
    layer6_outputs(457) <= '0';
    layer6_outputs(458) <= not((layer5_outputs(4888)) and (layer5_outputs(619)));
    layer6_outputs(459) <= layer5_outputs(4165);
    layer6_outputs(460) <= not(layer5_outputs(2398));
    layer6_outputs(461) <= not(layer5_outputs(3216));
    layer6_outputs(462) <= (layer5_outputs(4106)) and not (layer5_outputs(1035));
    layer6_outputs(463) <= not((layer5_outputs(2830)) or (layer5_outputs(2974)));
    layer6_outputs(464) <= not((layer5_outputs(4822)) and (layer5_outputs(55)));
    layer6_outputs(465) <= layer5_outputs(1015);
    layer6_outputs(466) <= not(layer5_outputs(3866));
    layer6_outputs(467) <= (layer5_outputs(4745)) and (layer5_outputs(1069));
    layer6_outputs(468) <= '0';
    layer6_outputs(469) <= not(layer5_outputs(2969));
    layer6_outputs(470) <= layer5_outputs(4914);
    layer6_outputs(471) <= not((layer5_outputs(5075)) and (layer5_outputs(1496)));
    layer6_outputs(472) <= not(layer5_outputs(3235));
    layer6_outputs(473) <= layer5_outputs(3673);
    layer6_outputs(474) <= (layer5_outputs(4257)) or (layer5_outputs(598));
    layer6_outputs(475) <= not(layer5_outputs(1555));
    layer6_outputs(476) <= not(layer5_outputs(2765));
    layer6_outputs(477) <= not(layer5_outputs(3582));
    layer6_outputs(478) <= not((layer5_outputs(2697)) and (layer5_outputs(3990)));
    layer6_outputs(479) <= not(layer5_outputs(1279));
    layer6_outputs(480) <= not((layer5_outputs(2500)) or (layer5_outputs(2570)));
    layer6_outputs(481) <= (layer5_outputs(4038)) xor (layer5_outputs(2662));
    layer6_outputs(482) <= '0';
    layer6_outputs(483) <= (layer5_outputs(2272)) or (layer5_outputs(1088));
    layer6_outputs(484) <= not(layer5_outputs(3317)) or (layer5_outputs(1029));
    layer6_outputs(485) <= '1';
    layer6_outputs(486) <= (layer5_outputs(4469)) and not (layer5_outputs(2493));
    layer6_outputs(487) <= not(layer5_outputs(1387)) or (layer5_outputs(3035));
    layer6_outputs(488) <= (layer5_outputs(5033)) xor (layer5_outputs(1910));
    layer6_outputs(489) <= not(layer5_outputs(2251));
    layer6_outputs(490) <= layer5_outputs(1610);
    layer6_outputs(491) <= not(layer5_outputs(1359));
    layer6_outputs(492) <= not((layer5_outputs(4441)) and (layer5_outputs(1118)));
    layer6_outputs(493) <= not((layer5_outputs(4118)) xor (layer5_outputs(2169)));
    layer6_outputs(494) <= not(layer5_outputs(3770));
    layer6_outputs(495) <= not(layer5_outputs(4637));
    layer6_outputs(496) <= not(layer5_outputs(3715)) or (layer5_outputs(575));
    layer6_outputs(497) <= (layer5_outputs(4946)) and not (layer5_outputs(5057));
    layer6_outputs(498) <= (layer5_outputs(3345)) and not (layer5_outputs(1732));
    layer6_outputs(499) <= not(layer5_outputs(1261));
    layer6_outputs(500) <= layer5_outputs(1776);
    layer6_outputs(501) <= (layer5_outputs(125)) or (layer5_outputs(1190));
    layer6_outputs(502) <= layer5_outputs(3077);
    layer6_outputs(503) <= (layer5_outputs(2276)) and not (layer5_outputs(1968));
    layer6_outputs(504) <= not(layer5_outputs(2620));
    layer6_outputs(505) <= layer5_outputs(3687);
    layer6_outputs(506) <= layer5_outputs(1263);
    layer6_outputs(507) <= (layer5_outputs(4365)) and not (layer5_outputs(1592));
    layer6_outputs(508) <= not(layer5_outputs(1676));
    layer6_outputs(509) <= not((layer5_outputs(1791)) or (layer5_outputs(4567)));
    layer6_outputs(510) <= not(layer5_outputs(799));
    layer6_outputs(511) <= not(layer5_outputs(1502));
    layer6_outputs(512) <= not((layer5_outputs(3113)) xor (layer5_outputs(2986)));
    layer6_outputs(513) <= not(layer5_outputs(3658));
    layer6_outputs(514) <= (layer5_outputs(719)) and not (layer5_outputs(2852));
    layer6_outputs(515) <= layer5_outputs(1272);
    layer6_outputs(516) <= (layer5_outputs(1805)) and not (layer5_outputs(256));
    layer6_outputs(517) <= not(layer5_outputs(1680)) or (layer5_outputs(3147));
    layer6_outputs(518) <= layer5_outputs(3579);
    layer6_outputs(519) <= (layer5_outputs(404)) or (layer5_outputs(4131));
    layer6_outputs(520) <= (layer5_outputs(1685)) or (layer5_outputs(3348));
    layer6_outputs(521) <= not(layer5_outputs(532));
    layer6_outputs(522) <= not(layer5_outputs(4041)) or (layer5_outputs(3941));
    layer6_outputs(523) <= layer5_outputs(3019);
    layer6_outputs(524) <= (layer5_outputs(4761)) and not (layer5_outputs(694));
    layer6_outputs(525) <= not((layer5_outputs(2210)) xor (layer5_outputs(5111)));
    layer6_outputs(526) <= not(layer5_outputs(1215));
    layer6_outputs(527) <= layer5_outputs(3431);
    layer6_outputs(528) <= not(layer5_outputs(3668)) or (layer5_outputs(3033));
    layer6_outputs(529) <= (layer5_outputs(1510)) or (layer5_outputs(3264));
    layer6_outputs(530) <= not(layer5_outputs(1252));
    layer6_outputs(531) <= layer5_outputs(906);
    layer6_outputs(532) <= not(layer5_outputs(3229)) or (layer5_outputs(978));
    layer6_outputs(533) <= not(layer5_outputs(5118));
    layer6_outputs(534) <= not((layer5_outputs(4493)) or (layer5_outputs(2440)));
    layer6_outputs(535) <= not(layer5_outputs(3594)) or (layer5_outputs(3578));
    layer6_outputs(536) <= layer5_outputs(163);
    layer6_outputs(537) <= (layer5_outputs(3300)) xor (layer5_outputs(133));
    layer6_outputs(538) <= layer5_outputs(2458);
    layer6_outputs(539) <= layer5_outputs(580);
    layer6_outputs(540) <= not((layer5_outputs(4760)) and (layer5_outputs(1262)));
    layer6_outputs(541) <= not(layer5_outputs(3493));
    layer6_outputs(542) <= layer5_outputs(2231);
    layer6_outputs(543) <= not((layer5_outputs(4043)) xor (layer5_outputs(4170)));
    layer6_outputs(544) <= not(layer5_outputs(4211));
    layer6_outputs(545) <= not(layer5_outputs(1664));
    layer6_outputs(546) <= '1';
    layer6_outputs(547) <= layer5_outputs(4127);
    layer6_outputs(548) <= (layer5_outputs(1207)) xor (layer5_outputs(3481));
    layer6_outputs(549) <= (layer5_outputs(1945)) and (layer5_outputs(4397));
    layer6_outputs(550) <= not(layer5_outputs(2455)) or (layer5_outputs(161));
    layer6_outputs(551) <= not(layer5_outputs(3927)) or (layer5_outputs(3011));
    layer6_outputs(552) <= layer5_outputs(1998);
    layer6_outputs(553) <= (layer5_outputs(329)) and (layer5_outputs(2625));
    layer6_outputs(554) <= (layer5_outputs(474)) and (layer5_outputs(5081));
    layer6_outputs(555) <= not((layer5_outputs(3533)) or (layer5_outputs(4623)));
    layer6_outputs(556) <= not(layer5_outputs(1701)) or (layer5_outputs(608));
    layer6_outputs(557) <= layer5_outputs(3185);
    layer6_outputs(558) <= not((layer5_outputs(2903)) and (layer5_outputs(5030)));
    layer6_outputs(559) <= not((layer5_outputs(3875)) and (layer5_outputs(4920)));
    layer6_outputs(560) <= (layer5_outputs(703)) and not (layer5_outputs(5110));
    layer6_outputs(561) <= (layer5_outputs(3570)) and (layer5_outputs(2391));
    layer6_outputs(562) <= (layer5_outputs(3172)) and not (layer5_outputs(2738));
    layer6_outputs(563) <= (layer5_outputs(4919)) and not (layer5_outputs(2672));
    layer6_outputs(564) <= '0';
    layer6_outputs(565) <= layer5_outputs(283);
    layer6_outputs(566) <= not((layer5_outputs(4936)) or (layer5_outputs(3558)));
    layer6_outputs(567) <= not(layer5_outputs(1505));
    layer6_outputs(568) <= not(layer5_outputs(943));
    layer6_outputs(569) <= '1';
    layer6_outputs(570) <= not(layer5_outputs(1026));
    layer6_outputs(571) <= not(layer5_outputs(3922));
    layer6_outputs(572) <= not((layer5_outputs(587)) and (layer5_outputs(672)));
    layer6_outputs(573) <= (layer5_outputs(3593)) xor (layer5_outputs(2985));
    layer6_outputs(574) <= layer5_outputs(640);
    layer6_outputs(575) <= layer5_outputs(4946);
    layer6_outputs(576) <= not((layer5_outputs(3344)) or (layer5_outputs(2975)));
    layer6_outputs(577) <= not(layer5_outputs(4206)) or (layer5_outputs(5088));
    layer6_outputs(578) <= not((layer5_outputs(38)) and (layer5_outputs(4638)));
    layer6_outputs(579) <= not((layer5_outputs(134)) or (layer5_outputs(3056)));
    layer6_outputs(580) <= layer5_outputs(5050);
    layer6_outputs(581) <= layer5_outputs(3097);
    layer6_outputs(582) <= not((layer5_outputs(2748)) and (layer5_outputs(3682)));
    layer6_outputs(583) <= layer5_outputs(4863);
    layer6_outputs(584) <= not(layer5_outputs(3762));
    layer6_outputs(585) <= not(layer5_outputs(4803));
    layer6_outputs(586) <= not(layer5_outputs(4873));
    layer6_outputs(587) <= (layer5_outputs(91)) or (layer5_outputs(2270));
    layer6_outputs(588) <= (layer5_outputs(750)) and not (layer5_outputs(1899));
    layer6_outputs(589) <= (layer5_outputs(2573)) and not (layer5_outputs(2841));
    layer6_outputs(590) <= not(layer5_outputs(4749));
    layer6_outputs(591) <= not(layer5_outputs(856));
    layer6_outputs(592) <= layer5_outputs(1429);
    layer6_outputs(593) <= not(layer5_outputs(352));
    layer6_outputs(594) <= layer5_outputs(5099);
    layer6_outputs(595) <= (layer5_outputs(1476)) and not (layer5_outputs(49));
    layer6_outputs(596) <= layer5_outputs(3510);
    layer6_outputs(597) <= not(layer5_outputs(203));
    layer6_outputs(598) <= not(layer5_outputs(3387)) or (layer5_outputs(5036));
    layer6_outputs(599) <= (layer5_outputs(4349)) xor (layer5_outputs(2936));
    layer6_outputs(600) <= not(layer5_outputs(1473));
    layer6_outputs(601) <= layer5_outputs(3141);
    layer6_outputs(602) <= not((layer5_outputs(3638)) xor (layer5_outputs(262)));
    layer6_outputs(603) <= not((layer5_outputs(2100)) and (layer5_outputs(1168)));
    layer6_outputs(604) <= layer5_outputs(5046);
    layer6_outputs(605) <= not(layer5_outputs(3821)) or (layer5_outputs(5039));
    layer6_outputs(606) <= (layer5_outputs(969)) or (layer5_outputs(3065));
    layer6_outputs(607) <= not((layer5_outputs(1764)) or (layer5_outputs(698)));
    layer6_outputs(608) <= not(layer5_outputs(3982));
    layer6_outputs(609) <= not(layer5_outputs(717)) or (layer5_outputs(2441));
    layer6_outputs(610) <= layer5_outputs(789);
    layer6_outputs(611) <= not(layer5_outputs(3507));
    layer6_outputs(612) <= not(layer5_outputs(478)) or (layer5_outputs(2105));
    layer6_outputs(613) <= not(layer5_outputs(490)) or (layer5_outputs(990));
    layer6_outputs(614) <= '1';
    layer6_outputs(615) <= not((layer5_outputs(805)) xor (layer5_outputs(3847)));
    layer6_outputs(616) <= (layer5_outputs(946)) and not (layer5_outputs(2307));
    layer6_outputs(617) <= not(layer5_outputs(939));
    layer6_outputs(618) <= not(layer5_outputs(2571));
    layer6_outputs(619) <= layer5_outputs(1378);
    layer6_outputs(620) <= not(layer5_outputs(3646));
    layer6_outputs(621) <= not((layer5_outputs(4157)) xor (layer5_outputs(2478)));
    layer6_outputs(622) <= not((layer5_outputs(1008)) and (layer5_outputs(3757)));
    layer6_outputs(623) <= not(layer5_outputs(3942)) or (layer5_outputs(237));
    layer6_outputs(624) <= layer5_outputs(3170);
    layer6_outputs(625) <= not(layer5_outputs(3966));
    layer6_outputs(626) <= not(layer5_outputs(4680));
    layer6_outputs(627) <= layer5_outputs(1506);
    layer6_outputs(628) <= not((layer5_outputs(1357)) or (layer5_outputs(3722)));
    layer6_outputs(629) <= not((layer5_outputs(3164)) and (layer5_outputs(3852)));
    layer6_outputs(630) <= (layer5_outputs(1421)) and (layer5_outputs(4194));
    layer6_outputs(631) <= (layer5_outputs(542)) and not (layer5_outputs(774));
    layer6_outputs(632) <= (layer5_outputs(4300)) and not (layer5_outputs(4725));
    layer6_outputs(633) <= layer5_outputs(512);
    layer6_outputs(634) <= (layer5_outputs(1599)) and (layer5_outputs(401));
    layer6_outputs(635) <= not(layer5_outputs(525)) or (layer5_outputs(2997));
    layer6_outputs(636) <= not(layer5_outputs(2480));
    layer6_outputs(637) <= (layer5_outputs(4275)) xor (layer5_outputs(349));
    layer6_outputs(638) <= not((layer5_outputs(99)) xor (layer5_outputs(4551)));
    layer6_outputs(639) <= (layer5_outputs(4463)) and (layer5_outputs(4538));
    layer6_outputs(640) <= (layer5_outputs(1129)) and not (layer5_outputs(2736));
    layer6_outputs(641) <= layer5_outputs(3148);
    layer6_outputs(642) <= not((layer5_outputs(1974)) xor (layer5_outputs(1163)));
    layer6_outputs(643) <= (layer5_outputs(973)) and (layer5_outputs(3439));
    layer6_outputs(644) <= layer5_outputs(678);
    layer6_outputs(645) <= layer5_outputs(2101);
    layer6_outputs(646) <= (layer5_outputs(2203)) xor (layer5_outputs(5078));
    layer6_outputs(647) <= (layer5_outputs(1017)) and (layer5_outputs(3038));
    layer6_outputs(648) <= not(layer5_outputs(3822));
    layer6_outputs(649) <= (layer5_outputs(4648)) xor (layer5_outputs(1542));
    layer6_outputs(650) <= not(layer5_outputs(4489));
    layer6_outputs(651) <= not(layer5_outputs(2338));
    layer6_outputs(652) <= layer5_outputs(1556);
    layer6_outputs(653) <= layer5_outputs(4534);
    layer6_outputs(654) <= not(layer5_outputs(955)) or (layer5_outputs(1841));
    layer6_outputs(655) <= (layer5_outputs(432)) and not (layer5_outputs(1095));
    layer6_outputs(656) <= not(layer5_outputs(3521));
    layer6_outputs(657) <= layer5_outputs(3957);
    layer6_outputs(658) <= not(layer5_outputs(4553));
    layer6_outputs(659) <= not(layer5_outputs(4423));
    layer6_outputs(660) <= not((layer5_outputs(2459)) xor (layer5_outputs(4078)));
    layer6_outputs(661) <= '0';
    layer6_outputs(662) <= not(layer5_outputs(4977));
    layer6_outputs(663) <= not(layer5_outputs(2241)) or (layer5_outputs(3052));
    layer6_outputs(664) <= '0';
    layer6_outputs(665) <= not(layer5_outputs(2008));
    layer6_outputs(666) <= (layer5_outputs(1070)) and not (layer5_outputs(2331));
    layer6_outputs(667) <= '0';
    layer6_outputs(668) <= layer5_outputs(2122);
    layer6_outputs(669) <= layer5_outputs(439);
    layer6_outputs(670) <= not((layer5_outputs(4037)) and (layer5_outputs(2166)));
    layer6_outputs(671) <= not(layer5_outputs(405));
    layer6_outputs(672) <= not((layer5_outputs(3436)) or (layer5_outputs(816)));
    layer6_outputs(673) <= (layer5_outputs(1790)) or (layer5_outputs(4750));
    layer6_outputs(674) <= not(layer5_outputs(4536));
    layer6_outputs(675) <= not((layer5_outputs(1994)) and (layer5_outputs(3125)));
    layer6_outputs(676) <= (layer5_outputs(976)) and not (layer5_outputs(4192));
    layer6_outputs(677) <= not(layer5_outputs(4190));
    layer6_outputs(678) <= not((layer5_outputs(2429)) xor (layer5_outputs(360)));
    layer6_outputs(679) <= not((layer5_outputs(981)) or (layer5_outputs(2987)));
    layer6_outputs(680) <= not(layer5_outputs(3002));
    layer6_outputs(681) <= not(layer5_outputs(4721)) or (layer5_outputs(2910));
    layer6_outputs(682) <= not(layer5_outputs(3205));
    layer6_outputs(683) <= not((layer5_outputs(1141)) or (layer5_outputs(215)));
    layer6_outputs(684) <= '0';
    layer6_outputs(685) <= (layer5_outputs(3306)) and not (layer5_outputs(1844));
    layer6_outputs(686) <= layer5_outputs(4974);
    layer6_outputs(687) <= layer5_outputs(33);
    layer6_outputs(688) <= '0';
    layer6_outputs(689) <= (layer5_outputs(3870)) xor (layer5_outputs(1192));
    layer6_outputs(690) <= not((layer5_outputs(3704)) or (layer5_outputs(2952)));
    layer6_outputs(691) <= not(layer5_outputs(1127)) or (layer5_outputs(3334));
    layer6_outputs(692) <= (layer5_outputs(4028)) and not (layer5_outputs(3110));
    layer6_outputs(693) <= '1';
    layer6_outputs(694) <= not(layer5_outputs(2642)) or (layer5_outputs(1244));
    layer6_outputs(695) <= (layer5_outputs(3509)) and not (layer5_outputs(2890));
    layer6_outputs(696) <= not(layer5_outputs(4790)) or (layer5_outputs(2456));
    layer6_outputs(697) <= (layer5_outputs(1589)) and not (layer5_outputs(2025));
    layer6_outputs(698) <= (layer5_outputs(2236)) and not (layer5_outputs(1672));
    layer6_outputs(699) <= not(layer5_outputs(471));
    layer6_outputs(700) <= (layer5_outputs(492)) and not (layer5_outputs(4723));
    layer6_outputs(701) <= (layer5_outputs(3728)) and (layer5_outputs(3815));
    layer6_outputs(702) <= not(layer5_outputs(1513));
    layer6_outputs(703) <= not((layer5_outputs(2199)) and (layer5_outputs(4570)));
    layer6_outputs(704) <= layer5_outputs(3283);
    layer6_outputs(705) <= layer5_outputs(4757);
    layer6_outputs(706) <= layer5_outputs(1292);
    layer6_outputs(707) <= not(layer5_outputs(1800)) or (layer5_outputs(5100));
    layer6_outputs(708) <= layer5_outputs(1837);
    layer6_outputs(709) <= '0';
    layer6_outputs(710) <= not(layer5_outputs(613)) or (layer5_outputs(1843));
    layer6_outputs(711) <= layer5_outputs(1596);
    layer6_outputs(712) <= layer5_outputs(3216);
    layer6_outputs(713) <= layer5_outputs(1538);
    layer6_outputs(714) <= not(layer5_outputs(1057));
    layer6_outputs(715) <= not(layer5_outputs(3279));
    layer6_outputs(716) <= (layer5_outputs(345)) and (layer5_outputs(2674));
    layer6_outputs(717) <= layer5_outputs(1616);
    layer6_outputs(718) <= '1';
    layer6_outputs(719) <= not((layer5_outputs(1977)) xor (layer5_outputs(255)));
    layer6_outputs(720) <= '1';
    layer6_outputs(721) <= (layer5_outputs(3264)) xor (layer5_outputs(2378));
    layer6_outputs(722) <= not(layer5_outputs(4690));
    layer6_outputs(723) <= not((layer5_outputs(3281)) xor (layer5_outputs(393)));
    layer6_outputs(724) <= not(layer5_outputs(1950));
    layer6_outputs(725) <= (layer5_outputs(2457)) xor (layer5_outputs(2538));
    layer6_outputs(726) <= not((layer5_outputs(2685)) or (layer5_outputs(927)));
    layer6_outputs(727) <= layer5_outputs(4838);
    layer6_outputs(728) <= layer5_outputs(2528);
    layer6_outputs(729) <= not((layer5_outputs(2080)) and (layer5_outputs(2233)));
    layer6_outputs(730) <= not((layer5_outputs(48)) and (layer5_outputs(4988)));
    layer6_outputs(731) <= not((layer5_outputs(4105)) or (layer5_outputs(3607)));
    layer6_outputs(732) <= not(layer5_outputs(761)) or (layer5_outputs(756));
    layer6_outputs(733) <= (layer5_outputs(1488)) xor (layer5_outputs(1313));
    layer6_outputs(734) <= layer5_outputs(3684);
    layer6_outputs(735) <= layer5_outputs(3381);
    layer6_outputs(736) <= not(layer5_outputs(579));
    layer6_outputs(737) <= not(layer5_outputs(2492));
    layer6_outputs(738) <= not(layer5_outputs(3423));
    layer6_outputs(739) <= (layer5_outputs(4971)) and not (layer5_outputs(104));
    layer6_outputs(740) <= not((layer5_outputs(3464)) or (layer5_outputs(685)));
    layer6_outputs(741) <= layer5_outputs(4477);
    layer6_outputs(742) <= not(layer5_outputs(1770));
    layer6_outputs(743) <= (layer5_outputs(3053)) and not (layer5_outputs(5));
    layer6_outputs(744) <= not(layer5_outputs(917));
    layer6_outputs(745) <= (layer5_outputs(875)) and not (layer5_outputs(4023));
    layer6_outputs(746) <= not((layer5_outputs(3270)) xor (layer5_outputs(68)));
    layer6_outputs(747) <= layer5_outputs(285);
    layer6_outputs(748) <= not((layer5_outputs(1653)) or (layer5_outputs(1411)));
    layer6_outputs(749) <= layer5_outputs(944);
    layer6_outputs(750) <= not((layer5_outputs(965)) and (layer5_outputs(3522)));
    layer6_outputs(751) <= (layer5_outputs(3989)) and (layer5_outputs(1581));
    layer6_outputs(752) <= layer5_outputs(1405);
    layer6_outputs(753) <= not(layer5_outputs(4341));
    layer6_outputs(754) <= not(layer5_outputs(626));
    layer6_outputs(755) <= (layer5_outputs(3053)) xor (layer5_outputs(1302));
    layer6_outputs(756) <= layer5_outputs(2918);
    layer6_outputs(757) <= not((layer5_outputs(801)) and (layer5_outputs(2688)));
    layer6_outputs(758) <= not((layer5_outputs(1407)) or (layer5_outputs(35)));
    layer6_outputs(759) <= '1';
    layer6_outputs(760) <= (layer5_outputs(2872)) and not (layer5_outputs(2862));
    layer6_outputs(761) <= not((layer5_outputs(4948)) and (layer5_outputs(4179)));
    layer6_outputs(762) <= not(layer5_outputs(2145)) or (layer5_outputs(2263));
    layer6_outputs(763) <= not(layer5_outputs(1116));
    layer6_outputs(764) <= layer5_outputs(1580);
    layer6_outputs(765) <= layer5_outputs(1901);
    layer6_outputs(766) <= not(layer5_outputs(5045));
    layer6_outputs(767) <= not(layer5_outputs(185)) or (layer5_outputs(2453));
    layer6_outputs(768) <= not(layer5_outputs(2775));
    layer6_outputs(769) <= not(layer5_outputs(4062));
    layer6_outputs(770) <= not(layer5_outputs(4740)) or (layer5_outputs(910));
    layer6_outputs(771) <= layer5_outputs(1308);
    layer6_outputs(772) <= not(layer5_outputs(3023)) or (layer5_outputs(5042));
    layer6_outputs(773) <= not(layer5_outputs(4237)) or (layer5_outputs(196));
    layer6_outputs(774) <= not((layer5_outputs(2420)) and (layer5_outputs(2336)));
    layer6_outputs(775) <= layer5_outputs(3020);
    layer6_outputs(776) <= (layer5_outputs(4522)) and not (layer5_outputs(1320));
    layer6_outputs(777) <= layer5_outputs(2488);
    layer6_outputs(778) <= (layer5_outputs(3766)) and not (layer5_outputs(3933));
    layer6_outputs(779) <= not((layer5_outputs(2259)) or (layer5_outputs(740)));
    layer6_outputs(780) <= not(layer5_outputs(4333)) or (layer5_outputs(4234));
    layer6_outputs(781) <= (layer5_outputs(3012)) and not (layer5_outputs(988));
    layer6_outputs(782) <= layer5_outputs(377);
    layer6_outputs(783) <= layer5_outputs(2997);
    layer6_outputs(784) <= not(layer5_outputs(1049));
    layer6_outputs(785) <= not(layer5_outputs(4128)) or (layer5_outputs(3622));
    layer6_outputs(786) <= '1';
    layer6_outputs(787) <= layer5_outputs(1784);
    layer6_outputs(788) <= layer5_outputs(1178);
    layer6_outputs(789) <= (layer5_outputs(1939)) and not (layer5_outputs(1232));
    layer6_outputs(790) <= (layer5_outputs(3742)) or (layer5_outputs(3833));
    layer6_outputs(791) <= not(layer5_outputs(733));
    layer6_outputs(792) <= (layer5_outputs(4932)) and (layer5_outputs(3087));
    layer6_outputs(793) <= not(layer5_outputs(3662)) or (layer5_outputs(4467));
    layer6_outputs(794) <= layer5_outputs(1519);
    layer6_outputs(795) <= (layer5_outputs(4812)) and not (layer5_outputs(4359));
    layer6_outputs(796) <= not(layer5_outputs(3102)) or (layer5_outputs(1338));
    layer6_outputs(797) <= (layer5_outputs(2366)) and (layer5_outputs(629));
    layer6_outputs(798) <= not(layer5_outputs(3130));
    layer6_outputs(799) <= (layer5_outputs(1473)) or (layer5_outputs(2293));
    layer6_outputs(800) <= (layer5_outputs(2014)) and not (layer5_outputs(2125));
    layer6_outputs(801) <= (layer5_outputs(2982)) and (layer5_outputs(2642));
    layer6_outputs(802) <= layer5_outputs(3788);
    layer6_outputs(803) <= (layer5_outputs(1672)) and not (layer5_outputs(3947));
    layer6_outputs(804) <= not(layer5_outputs(2973));
    layer6_outputs(805) <= (layer5_outputs(3565)) or (layer5_outputs(1018));
    layer6_outputs(806) <= (layer5_outputs(96)) or (layer5_outputs(3574));
    layer6_outputs(807) <= not((layer5_outputs(2764)) or (layer5_outputs(3460)));
    layer6_outputs(808) <= layer5_outputs(4563);
    layer6_outputs(809) <= not(layer5_outputs(3907));
    layer6_outputs(810) <= not(layer5_outputs(2904));
    layer6_outputs(811) <= (layer5_outputs(3307)) xor (layer5_outputs(3545));
    layer6_outputs(812) <= (layer5_outputs(1693)) xor (layer5_outputs(2308));
    layer6_outputs(813) <= not(layer5_outputs(2125));
    layer6_outputs(814) <= layer5_outputs(1602);
    layer6_outputs(815) <= not(layer5_outputs(246));
    layer6_outputs(816) <= layer5_outputs(4214);
    layer6_outputs(817) <= layer5_outputs(1850);
    layer6_outputs(818) <= not(layer5_outputs(2767)) or (layer5_outputs(4498));
    layer6_outputs(819) <= not(layer5_outputs(3478)) or (layer5_outputs(4517));
    layer6_outputs(820) <= not(layer5_outputs(4475));
    layer6_outputs(821) <= not((layer5_outputs(1394)) or (layer5_outputs(4013)));
    layer6_outputs(822) <= (layer5_outputs(5019)) or (layer5_outputs(517));
    layer6_outputs(823) <= layer5_outputs(3342);
    layer6_outputs(824) <= not(layer5_outputs(1971)) or (layer5_outputs(812));
    layer6_outputs(825) <= (layer5_outputs(3677)) and not (layer5_outputs(2867));
    layer6_outputs(826) <= not(layer5_outputs(1912)) or (layer5_outputs(2564));
    layer6_outputs(827) <= not(layer5_outputs(3969));
    layer6_outputs(828) <= not(layer5_outputs(817));
    layer6_outputs(829) <= layer5_outputs(4422);
    layer6_outputs(830) <= not(layer5_outputs(3935));
    layer6_outputs(831) <= not(layer5_outputs(536)) or (layer5_outputs(3318));
    layer6_outputs(832) <= layer5_outputs(1784);
    layer6_outputs(833) <= not(layer5_outputs(2803)) or (layer5_outputs(4431));
    layer6_outputs(834) <= '1';
    layer6_outputs(835) <= layer5_outputs(4371);
    layer6_outputs(836) <= (layer5_outputs(4872)) and not (layer5_outputs(1064));
    layer6_outputs(837) <= (layer5_outputs(3424)) or (layer5_outputs(2683));
    layer6_outputs(838) <= (layer5_outputs(2772)) and not (layer5_outputs(3652));
    layer6_outputs(839) <= not(layer5_outputs(1535));
    layer6_outputs(840) <= not(layer5_outputs(3895));
    layer6_outputs(841) <= '0';
    layer6_outputs(842) <= not(layer5_outputs(752)) or (layer5_outputs(5101));
    layer6_outputs(843) <= (layer5_outputs(263)) and (layer5_outputs(844));
    layer6_outputs(844) <= not((layer5_outputs(2474)) and (layer5_outputs(3763)));
    layer6_outputs(845) <= '0';
    layer6_outputs(846) <= layer5_outputs(4509);
    layer6_outputs(847) <= not((layer5_outputs(395)) xor (layer5_outputs(3411)));
    layer6_outputs(848) <= '0';
    layer6_outputs(849) <= (layer5_outputs(111)) xor (layer5_outputs(49));
    layer6_outputs(850) <= not(layer5_outputs(1105));
    layer6_outputs(851) <= (layer5_outputs(5113)) and not (layer5_outputs(3843));
    layer6_outputs(852) <= layer5_outputs(1373);
    layer6_outputs(853) <= not(layer5_outputs(237));
    layer6_outputs(854) <= layer5_outputs(3946);
    layer6_outputs(855) <= not(layer5_outputs(3811));
    layer6_outputs(856) <= (layer5_outputs(788)) and not (layer5_outputs(5114));
    layer6_outputs(857) <= (layer5_outputs(454)) xor (layer5_outputs(1076));
    layer6_outputs(858) <= (layer5_outputs(4225)) and not (layer5_outputs(1586));
    layer6_outputs(859) <= not((layer5_outputs(2187)) and (layer5_outputs(4022)));
    layer6_outputs(860) <= not(layer5_outputs(4797));
    layer6_outputs(861) <= not((layer5_outputs(881)) or (layer5_outputs(3538)));
    layer6_outputs(862) <= not((layer5_outputs(1761)) or (layer5_outputs(4067)));
    layer6_outputs(863) <= '0';
    layer6_outputs(864) <= not(layer5_outputs(3839)) or (layer5_outputs(621));
    layer6_outputs(865) <= not((layer5_outputs(699)) or (layer5_outputs(833)));
    layer6_outputs(866) <= not(layer5_outputs(4313));
    layer6_outputs(867) <= (layer5_outputs(960)) and not (layer5_outputs(214));
    layer6_outputs(868) <= (layer5_outputs(716)) and not (layer5_outputs(442));
    layer6_outputs(869) <= (layer5_outputs(1833)) or (layer5_outputs(3681));
    layer6_outputs(870) <= not(layer5_outputs(459)) or (layer5_outputs(977));
    layer6_outputs(871) <= not((layer5_outputs(4823)) xor (layer5_outputs(3483)));
    layer6_outputs(872) <= (layer5_outputs(4956)) and (layer5_outputs(4217));
    layer6_outputs(873) <= not(layer5_outputs(3915));
    layer6_outputs(874) <= not((layer5_outputs(607)) xor (layer5_outputs(2247)));
    layer6_outputs(875) <= not(layer5_outputs(1204));
    layer6_outputs(876) <= not((layer5_outputs(2546)) or (layer5_outputs(2781)));
    layer6_outputs(877) <= not(layer5_outputs(3237)) or (layer5_outputs(1218));
    layer6_outputs(878) <= not((layer5_outputs(481)) xor (layer5_outputs(2681)));
    layer6_outputs(879) <= layer5_outputs(1601);
    layer6_outputs(880) <= '1';
    layer6_outputs(881) <= not(layer5_outputs(4492));
    layer6_outputs(882) <= '0';
    layer6_outputs(883) <= not(layer5_outputs(1393));
    layer6_outputs(884) <= not(layer5_outputs(5010));
    layer6_outputs(885) <= not(layer5_outputs(696));
    layer6_outputs(886) <= not(layer5_outputs(3885));
    layer6_outputs(887) <= not(layer5_outputs(1043));
    layer6_outputs(888) <= layer5_outputs(4069);
    layer6_outputs(889) <= not(layer5_outputs(3849));
    layer6_outputs(890) <= not((layer5_outputs(413)) and (layer5_outputs(1938)));
    layer6_outputs(891) <= not(layer5_outputs(1362));
    layer6_outputs(892) <= not(layer5_outputs(2570));
    layer6_outputs(893) <= not((layer5_outputs(4003)) or (layer5_outputs(2064)));
    layer6_outputs(894) <= (layer5_outputs(2120)) and not (layer5_outputs(1149));
    layer6_outputs(895) <= (layer5_outputs(2837)) and not (layer5_outputs(1266));
    layer6_outputs(896) <= (layer5_outputs(4905)) and not (layer5_outputs(2666));
    layer6_outputs(897) <= layer5_outputs(3003);
    layer6_outputs(898) <= layer5_outputs(1314);
    layer6_outputs(899) <= layer5_outputs(181);
    layer6_outputs(900) <= not(layer5_outputs(4787));
    layer6_outputs(901) <= layer5_outputs(4422);
    layer6_outputs(902) <= not(layer5_outputs(2545)) or (layer5_outputs(2422));
    layer6_outputs(903) <= layer5_outputs(2364);
    layer6_outputs(904) <= layer5_outputs(351);
    layer6_outputs(905) <= layer5_outputs(1472);
    layer6_outputs(906) <= not(layer5_outputs(3359));
    layer6_outputs(907) <= not((layer5_outputs(89)) and (layer5_outputs(2655)));
    layer6_outputs(908) <= layer5_outputs(4944);
    layer6_outputs(909) <= (layer5_outputs(3721)) and (layer5_outputs(2140));
    layer6_outputs(910) <= (layer5_outputs(3503)) or (layer5_outputs(57));
    layer6_outputs(911) <= not(layer5_outputs(825));
    layer6_outputs(912) <= not(layer5_outputs(1541)) or (layer5_outputs(757));
    layer6_outputs(913) <= not((layer5_outputs(2457)) and (layer5_outputs(1969)));
    layer6_outputs(914) <= not(layer5_outputs(2080));
    layer6_outputs(915) <= not(layer5_outputs(3798));
    layer6_outputs(916) <= layer5_outputs(2552);
    layer6_outputs(917) <= not(layer5_outputs(4917));
    layer6_outputs(918) <= not(layer5_outputs(1213)) or (layer5_outputs(3059));
    layer6_outputs(919) <= not((layer5_outputs(4448)) or (layer5_outputs(3950)));
    layer6_outputs(920) <= layer5_outputs(4465);
    layer6_outputs(921) <= layer5_outputs(3710);
    layer6_outputs(922) <= not(layer5_outputs(2164));
    layer6_outputs(923) <= not(layer5_outputs(4169));
    layer6_outputs(924) <= (layer5_outputs(1527)) and (layer5_outputs(2917));
    layer6_outputs(925) <= (layer5_outputs(97)) and not (layer5_outputs(712));
    layer6_outputs(926) <= not((layer5_outputs(1431)) xor (layer5_outputs(2676)));
    layer6_outputs(927) <= not((layer5_outputs(219)) and (layer5_outputs(1592)));
    layer6_outputs(928) <= not(layer5_outputs(2807));
    layer6_outputs(929) <= layer5_outputs(595);
    layer6_outputs(930) <= not(layer5_outputs(4632));
    layer6_outputs(931) <= layer5_outputs(1187);
    layer6_outputs(932) <= layer5_outputs(986);
    layer6_outputs(933) <= not(layer5_outputs(1745));
    layer6_outputs(934) <= layer5_outputs(3033);
    layer6_outputs(935) <= (layer5_outputs(2820)) and (layer5_outputs(2978));
    layer6_outputs(936) <= not((layer5_outputs(637)) xor (layer5_outputs(2562)));
    layer6_outputs(937) <= not(layer5_outputs(403)) or (layer5_outputs(2175));
    layer6_outputs(938) <= layer5_outputs(2492);
    layer6_outputs(939) <= layer5_outputs(1920);
    layer6_outputs(940) <= not((layer5_outputs(2666)) xor (layer5_outputs(2291)));
    layer6_outputs(941) <= layer5_outputs(2327);
    layer6_outputs(942) <= not(layer5_outputs(967));
    layer6_outputs(943) <= '0';
    layer6_outputs(944) <= not(layer5_outputs(1604));
    layer6_outputs(945) <= (layer5_outputs(4461)) or (layer5_outputs(3471));
    layer6_outputs(946) <= layer5_outputs(4296);
    layer6_outputs(947) <= layer5_outputs(2914);
    layer6_outputs(948) <= layer5_outputs(3954);
    layer6_outputs(949) <= layer5_outputs(3620);
    layer6_outputs(950) <= not((layer5_outputs(4053)) or (layer5_outputs(3745)));
    layer6_outputs(951) <= not(layer5_outputs(1243));
    layer6_outputs(952) <= layer5_outputs(4288);
    layer6_outputs(953) <= layer5_outputs(3000);
    layer6_outputs(954) <= layer5_outputs(4023);
    layer6_outputs(955) <= (layer5_outputs(3746)) and not (layer5_outputs(2242));
    layer6_outputs(956) <= (layer5_outputs(3601)) xor (layer5_outputs(102));
    layer6_outputs(957) <= not((layer5_outputs(2675)) and (layer5_outputs(4966)));
    layer6_outputs(958) <= not(layer5_outputs(1275));
    layer6_outputs(959) <= not(layer5_outputs(2726));
    layer6_outputs(960) <= layer5_outputs(2273);
    layer6_outputs(961) <= not(layer5_outputs(2764));
    layer6_outputs(962) <= layer5_outputs(4648);
    layer6_outputs(963) <= not(layer5_outputs(4406)) or (layer5_outputs(2155));
    layer6_outputs(964) <= not((layer5_outputs(3530)) and (layer5_outputs(3506)));
    layer6_outputs(965) <= not((layer5_outputs(535)) xor (layer5_outputs(2540)));
    layer6_outputs(966) <= (layer5_outputs(2968)) and not (layer5_outputs(3526));
    layer6_outputs(967) <= layer5_outputs(1426);
    layer6_outputs(968) <= (layer5_outputs(4439)) and not (layer5_outputs(1700));
    layer6_outputs(969) <= layer5_outputs(3434);
    layer6_outputs(970) <= (layer5_outputs(3073)) and not (layer5_outputs(826));
    layer6_outputs(971) <= layer5_outputs(2280);
    layer6_outputs(972) <= layer5_outputs(1516);
    layer6_outputs(973) <= not((layer5_outputs(3015)) and (layer5_outputs(4625)));
    layer6_outputs(974) <= layer5_outputs(627);
    layer6_outputs(975) <= (layer5_outputs(3687)) and not (layer5_outputs(2264));
    layer6_outputs(976) <= not(layer5_outputs(4529)) or (layer5_outputs(4731));
    layer6_outputs(977) <= (layer5_outputs(3255)) and not (layer5_outputs(2432));
    layer6_outputs(978) <= (layer5_outputs(266)) and not (layer5_outputs(3735));
    layer6_outputs(979) <= not((layer5_outputs(748)) xor (layer5_outputs(289)));
    layer6_outputs(980) <= (layer5_outputs(4018)) and (layer5_outputs(3596));
    layer6_outputs(981) <= not(layer5_outputs(3905));
    layer6_outputs(982) <= not(layer5_outputs(896));
    layer6_outputs(983) <= '1';
    layer6_outputs(984) <= layer5_outputs(458);
    layer6_outputs(985) <= (layer5_outputs(323)) and (layer5_outputs(3648));
    layer6_outputs(986) <= '0';
    layer6_outputs(987) <= layer5_outputs(311);
    layer6_outputs(988) <= layer5_outputs(892);
    layer6_outputs(989) <= not((layer5_outputs(4277)) and (layer5_outputs(1186)));
    layer6_outputs(990) <= not(layer5_outputs(460));
    layer6_outputs(991) <= (layer5_outputs(3106)) and not (layer5_outputs(4087));
    layer6_outputs(992) <= (layer5_outputs(1394)) and not (layer5_outputs(1094));
    layer6_outputs(993) <= (layer5_outputs(2053)) and not (layer5_outputs(3617));
    layer6_outputs(994) <= not(layer5_outputs(4092));
    layer6_outputs(995) <= not(layer5_outputs(3939));
    layer6_outputs(996) <= not((layer5_outputs(365)) and (layer5_outputs(2259)));
    layer6_outputs(997) <= (layer5_outputs(3587)) and (layer5_outputs(794));
    layer6_outputs(998) <= not(layer5_outputs(838));
    layer6_outputs(999) <= layer5_outputs(1432);
    layer6_outputs(1000) <= (layer5_outputs(1567)) and not (layer5_outputs(1220));
    layer6_outputs(1001) <= not((layer5_outputs(5054)) or (layer5_outputs(3402)));
    layer6_outputs(1002) <= not(layer5_outputs(4759));
    layer6_outputs(1003) <= '1';
    layer6_outputs(1004) <= not(layer5_outputs(1637));
    layer6_outputs(1005) <= (layer5_outputs(3876)) and (layer5_outputs(2903));
    layer6_outputs(1006) <= layer5_outputs(4934);
    layer6_outputs(1007) <= not((layer5_outputs(3669)) or (layer5_outputs(4586)));
    layer6_outputs(1008) <= not(layer5_outputs(317));
    layer6_outputs(1009) <= '1';
    layer6_outputs(1010) <= not(layer5_outputs(3010)) or (layer5_outputs(2090));
    layer6_outputs(1011) <= not(layer5_outputs(4767));
    layer6_outputs(1012) <= (layer5_outputs(4545)) and (layer5_outputs(2725));
    layer6_outputs(1013) <= layer5_outputs(324);
    layer6_outputs(1014) <= not(layer5_outputs(4856));
    layer6_outputs(1015) <= not(layer5_outputs(2107));
    layer6_outputs(1016) <= not(layer5_outputs(2156)) or (layer5_outputs(4628));
    layer6_outputs(1017) <= not(layer5_outputs(707));
    layer6_outputs(1018) <= layer5_outputs(1517);
    layer6_outputs(1019) <= not((layer5_outputs(572)) or (layer5_outputs(4511)));
    layer6_outputs(1020) <= (layer5_outputs(2383)) and not (layer5_outputs(207));
    layer6_outputs(1021) <= layer5_outputs(4777);
    layer6_outputs(1022) <= layer5_outputs(1961);
    layer6_outputs(1023) <= '1';
    layer6_outputs(1024) <= (layer5_outputs(477)) and not (layer5_outputs(4242));
    layer6_outputs(1025) <= not((layer5_outputs(1325)) and (layer5_outputs(4606)));
    layer6_outputs(1026) <= not((layer5_outputs(2674)) xor (layer5_outputs(272)));
    layer6_outputs(1027) <= not(layer5_outputs(3209));
    layer6_outputs(1028) <= not((layer5_outputs(4259)) or (layer5_outputs(1436)));
    layer6_outputs(1029) <= layer5_outputs(2595);
    layer6_outputs(1030) <= not((layer5_outputs(4944)) xor (layer5_outputs(2660)));
    layer6_outputs(1031) <= not(layer5_outputs(3333)) or (layer5_outputs(1079));
    layer6_outputs(1032) <= not(layer5_outputs(1127));
    layer6_outputs(1033) <= not(layer5_outputs(594));
    layer6_outputs(1034) <= (layer5_outputs(1844)) or (layer5_outputs(3856));
    layer6_outputs(1035) <= (layer5_outputs(745)) and not (layer5_outputs(568));
    layer6_outputs(1036) <= not(layer5_outputs(303));
    layer6_outputs(1037) <= not(layer5_outputs(1194)) or (layer5_outputs(1704));
    layer6_outputs(1038) <= not(layer5_outputs(2850)) or (layer5_outputs(2689));
    layer6_outputs(1039) <= (layer5_outputs(4323)) xor (layer5_outputs(1796));
    layer6_outputs(1040) <= layer5_outputs(3499);
    layer6_outputs(1041) <= layer5_outputs(4144);
    layer6_outputs(1042) <= (layer5_outputs(4901)) xor (layer5_outputs(1883));
    layer6_outputs(1043) <= (layer5_outputs(2483)) and not (layer5_outputs(4851));
    layer6_outputs(1044) <= (layer5_outputs(2220)) or (layer5_outputs(2984));
    layer6_outputs(1045) <= not(layer5_outputs(230));
    layer6_outputs(1046) <= (layer5_outputs(2179)) xor (layer5_outputs(4835));
    layer6_outputs(1047) <= layer5_outputs(2096);
    layer6_outputs(1048) <= not(layer5_outputs(4925));
    layer6_outputs(1049) <= not(layer5_outputs(3026));
    layer6_outputs(1050) <= not(layer5_outputs(4870)) or (layer5_outputs(4999));
    layer6_outputs(1051) <= not(layer5_outputs(2200)) or (layer5_outputs(2031));
    layer6_outputs(1052) <= layer5_outputs(3823);
    layer6_outputs(1053) <= layer5_outputs(630);
    layer6_outputs(1054) <= not((layer5_outputs(3090)) or (layer5_outputs(1685)));
    layer6_outputs(1055) <= layer5_outputs(1235);
    layer6_outputs(1056) <= not(layer5_outputs(687));
    layer6_outputs(1057) <= (layer5_outputs(4947)) and not (layer5_outputs(1925));
    layer6_outputs(1058) <= layer5_outputs(491);
    layer6_outputs(1059) <= layer5_outputs(4229);
    layer6_outputs(1060) <= not(layer5_outputs(4305));
    layer6_outputs(1061) <= not(layer5_outputs(1995)) or (layer5_outputs(1446));
    layer6_outputs(1062) <= layer5_outputs(2229);
    layer6_outputs(1063) <= layer5_outputs(4907);
    layer6_outputs(1064) <= not(layer5_outputs(2246)) or (layer5_outputs(3068));
    layer6_outputs(1065) <= layer5_outputs(3438);
    layer6_outputs(1066) <= '0';
    layer6_outputs(1067) <= not((layer5_outputs(606)) or (layer5_outputs(1228)));
    layer6_outputs(1068) <= not((layer5_outputs(4238)) or (layer5_outputs(1294)));
    layer6_outputs(1069) <= not(layer5_outputs(3252));
    layer6_outputs(1070) <= not((layer5_outputs(721)) and (layer5_outputs(1084)));
    layer6_outputs(1071) <= (layer5_outputs(3090)) and not (layer5_outputs(1257));
    layer6_outputs(1072) <= (layer5_outputs(3579)) and not (layer5_outputs(2791));
    layer6_outputs(1073) <= not(layer5_outputs(1310)) or (layer5_outputs(1775));
    layer6_outputs(1074) <= not(layer5_outputs(1016));
    layer6_outputs(1075) <= not((layer5_outputs(1018)) xor (layer5_outputs(3410)));
    layer6_outputs(1076) <= not(layer5_outputs(638));
    layer6_outputs(1077) <= layer5_outputs(2301);
    layer6_outputs(1078) <= not((layer5_outputs(2191)) or (layer5_outputs(2819)));
    layer6_outputs(1079) <= not((layer5_outputs(3767)) or (layer5_outputs(4774)));
    layer6_outputs(1080) <= '0';
    layer6_outputs(1081) <= not((layer5_outputs(2377)) and (layer5_outputs(2852)));
    layer6_outputs(1082) <= not(layer5_outputs(2202)) or (layer5_outputs(1829));
    layer6_outputs(1083) <= not(layer5_outputs(1126)) or (layer5_outputs(2432));
    layer6_outputs(1084) <= not(layer5_outputs(1185)) or (layer5_outputs(3718));
    layer6_outputs(1085) <= not((layer5_outputs(1131)) xor (layer5_outputs(4135)));
    layer6_outputs(1086) <= layer5_outputs(3117);
    layer6_outputs(1087) <= (layer5_outputs(3701)) or (layer5_outputs(1249));
    layer6_outputs(1088) <= not(layer5_outputs(1637));
    layer6_outputs(1089) <= not(layer5_outputs(3641));
    layer6_outputs(1090) <= (layer5_outputs(1489)) and not (layer5_outputs(3305));
    layer6_outputs(1091) <= not((layer5_outputs(422)) xor (layer5_outputs(3909)));
    layer6_outputs(1092) <= (layer5_outputs(3370)) and not (layer5_outputs(3577));
    layer6_outputs(1093) <= not(layer5_outputs(990));
    layer6_outputs(1094) <= not(layer5_outputs(499));
    layer6_outputs(1095) <= not(layer5_outputs(1918));
    layer6_outputs(1096) <= layer5_outputs(185);
    layer6_outputs(1097) <= not((layer5_outputs(1897)) xor (layer5_outputs(481)));
    layer6_outputs(1098) <= layer5_outputs(2810);
    layer6_outputs(1099) <= not((layer5_outputs(3269)) or (layer5_outputs(1752)));
    layer6_outputs(1100) <= not(layer5_outputs(900));
    layer6_outputs(1101) <= (layer5_outputs(4175)) and (layer5_outputs(3918));
    layer6_outputs(1102) <= not(layer5_outputs(1834));
    layer6_outputs(1103) <= (layer5_outputs(1575)) and (layer5_outputs(1530));
    layer6_outputs(1104) <= not(layer5_outputs(1512)) or (layer5_outputs(834));
    layer6_outputs(1105) <= (layer5_outputs(2929)) or (layer5_outputs(1013));
    layer6_outputs(1106) <= not(layer5_outputs(381));
    layer6_outputs(1107) <= not((layer5_outputs(4614)) xor (layer5_outputs(2938)));
    layer6_outputs(1108) <= (layer5_outputs(4427)) or (layer5_outputs(3286));
    layer6_outputs(1109) <= layer5_outputs(1416);
    layer6_outputs(1110) <= layer5_outputs(1881);
    layer6_outputs(1111) <= not(layer5_outputs(63));
    layer6_outputs(1112) <= not(layer5_outputs(4002));
    layer6_outputs(1113) <= not(layer5_outputs(4095));
    layer6_outputs(1114) <= not(layer5_outputs(375));
    layer6_outputs(1115) <= not((layer5_outputs(398)) xor (layer5_outputs(2275)));
    layer6_outputs(1116) <= (layer5_outputs(1042)) xor (layer5_outputs(2261));
    layer6_outputs(1117) <= not(layer5_outputs(15));
    layer6_outputs(1118) <= not(layer5_outputs(3470));
    layer6_outputs(1119) <= not(layer5_outputs(3401)) or (layer5_outputs(2963));
    layer6_outputs(1120) <= layer5_outputs(2127);
    layer6_outputs(1121) <= not(layer5_outputs(2593));
    layer6_outputs(1122) <= (layer5_outputs(2695)) or (layer5_outputs(4214));
    layer6_outputs(1123) <= not(layer5_outputs(4994));
    layer6_outputs(1124) <= (layer5_outputs(457)) and not (layer5_outputs(4902));
    layer6_outputs(1125) <= (layer5_outputs(1970)) and not (layer5_outputs(3710));
    layer6_outputs(1126) <= not(layer5_outputs(3383));
    layer6_outputs(1127) <= not(layer5_outputs(706));
    layer6_outputs(1128) <= not((layer5_outputs(2707)) xor (layer5_outputs(2861)));
    layer6_outputs(1129) <= layer5_outputs(1709);
    layer6_outputs(1130) <= not(layer5_outputs(3029)) or (layer5_outputs(4141));
    layer6_outputs(1131) <= (layer5_outputs(3623)) and (layer5_outputs(2534));
    layer6_outputs(1132) <= not(layer5_outputs(4143));
    layer6_outputs(1133) <= layer5_outputs(4635);
    layer6_outputs(1134) <= layer5_outputs(4379);
    layer6_outputs(1135) <= layer5_outputs(1749);
    layer6_outputs(1136) <= (layer5_outputs(2211)) and (layer5_outputs(4933));
    layer6_outputs(1137) <= layer5_outputs(2314);
    layer6_outputs(1138) <= not(layer5_outputs(3180)) or (layer5_outputs(3829));
    layer6_outputs(1139) <= not((layer5_outputs(224)) or (layer5_outputs(2297)));
    layer6_outputs(1140) <= (layer5_outputs(4516)) xor (layer5_outputs(4806));
    layer6_outputs(1141) <= not(layer5_outputs(1773)) or (layer5_outputs(5026));
    layer6_outputs(1142) <= layer5_outputs(3462);
    layer6_outputs(1143) <= not(layer5_outputs(353));
    layer6_outputs(1144) <= not(layer5_outputs(1981));
    layer6_outputs(1145) <= (layer5_outputs(5061)) and not (layer5_outputs(4938));
    layer6_outputs(1146) <= (layer5_outputs(1198)) and (layer5_outputs(1643));
    layer6_outputs(1147) <= not(layer5_outputs(4715));
    layer6_outputs(1148) <= layer5_outputs(4481);
    layer6_outputs(1149) <= layer5_outputs(2564);
    layer6_outputs(1150) <= (layer5_outputs(1276)) and not (layer5_outputs(4816));
    layer6_outputs(1151) <= (layer5_outputs(2322)) and (layer5_outputs(1049));
    layer6_outputs(1152) <= not(layer5_outputs(1732));
    layer6_outputs(1153) <= not((layer5_outputs(1867)) or (layer5_outputs(2136)));
    layer6_outputs(1154) <= (layer5_outputs(644)) and not (layer5_outputs(2288));
    layer6_outputs(1155) <= layer5_outputs(1913);
    layer6_outputs(1156) <= layer5_outputs(4622);
    layer6_outputs(1157) <= not(layer5_outputs(1060)) or (layer5_outputs(3310));
    layer6_outputs(1158) <= not((layer5_outputs(4051)) xor (layer5_outputs(3355)));
    layer6_outputs(1159) <= not((layer5_outputs(2040)) and (layer5_outputs(5015)));
    layer6_outputs(1160) <= layer5_outputs(3496);
    layer6_outputs(1161) <= not((layer5_outputs(1997)) xor (layer5_outputs(3094)));
    layer6_outputs(1162) <= not(layer5_outputs(4386));
    layer6_outputs(1163) <= (layer5_outputs(840)) and not (layer5_outputs(1418));
    layer6_outputs(1164) <= not(layer5_outputs(995));
    layer6_outputs(1165) <= (layer5_outputs(1159)) xor (layer5_outputs(2072));
    layer6_outputs(1166) <= not(layer5_outputs(1713));
    layer6_outputs(1167) <= not(layer5_outputs(1327)) or (layer5_outputs(1434));
    layer6_outputs(1168) <= layer5_outputs(2169);
    layer6_outputs(1169) <= layer5_outputs(4910);
    layer6_outputs(1170) <= not(layer5_outputs(2319));
    layer6_outputs(1171) <= not((layer5_outputs(2561)) xor (layer5_outputs(1573)));
    layer6_outputs(1172) <= not(layer5_outputs(4380));
    layer6_outputs(1173) <= layer5_outputs(1397);
    layer6_outputs(1174) <= not(layer5_outputs(804)) or (layer5_outputs(2587));
    layer6_outputs(1175) <= (layer5_outputs(773)) and not (layer5_outputs(464));
    layer6_outputs(1176) <= not(layer5_outputs(4630));
    layer6_outputs(1177) <= (layer5_outputs(2109)) and not (layer5_outputs(4242));
    layer6_outputs(1178) <= not((layer5_outputs(4566)) or (layer5_outputs(3318)));
    layer6_outputs(1179) <= '1';
    layer6_outputs(1180) <= not((layer5_outputs(5050)) xor (layer5_outputs(4161)));
    layer6_outputs(1181) <= layer5_outputs(170);
    layer6_outputs(1182) <= not((layer5_outputs(1125)) xor (layer5_outputs(4908)));
    layer6_outputs(1183) <= layer5_outputs(4755);
    layer6_outputs(1184) <= layer5_outputs(3108);
    layer6_outputs(1185) <= layer5_outputs(2399);
    layer6_outputs(1186) <= not(layer5_outputs(2640));
    layer6_outputs(1187) <= not(layer5_outputs(1330));
    layer6_outputs(1188) <= '0';
    layer6_outputs(1189) <= (layer5_outputs(1019)) or (layer5_outputs(4045));
    layer6_outputs(1190) <= layer5_outputs(1955);
    layer6_outputs(1191) <= layer5_outputs(4416);
    layer6_outputs(1192) <= (layer5_outputs(569)) or (layer5_outputs(3064));
    layer6_outputs(1193) <= not(layer5_outputs(1795));
    layer6_outputs(1194) <= not((layer5_outputs(2957)) or (layer5_outputs(3160)));
    layer6_outputs(1195) <= layer5_outputs(3615);
    layer6_outputs(1196) <= not(layer5_outputs(4215));
    layer6_outputs(1197) <= (layer5_outputs(341)) or (layer5_outputs(3712));
    layer6_outputs(1198) <= layer5_outputs(3350);
    layer6_outputs(1199) <= (layer5_outputs(1401)) xor (layer5_outputs(2194));
    layer6_outputs(1200) <= not(layer5_outputs(2947)) or (layer5_outputs(3442));
    layer6_outputs(1201) <= layer5_outputs(1837);
    layer6_outputs(1202) <= '1';
    layer6_outputs(1203) <= not(layer5_outputs(848));
    layer6_outputs(1204) <= (layer5_outputs(3618)) or (layer5_outputs(4552));
    layer6_outputs(1205) <= layer5_outputs(4914);
    layer6_outputs(1206) <= not((layer5_outputs(4300)) or (layer5_outputs(4835)));
    layer6_outputs(1207) <= layer5_outputs(1870);
    layer6_outputs(1208) <= not(layer5_outputs(86));
    layer6_outputs(1209) <= (layer5_outputs(4635)) or (layer5_outputs(3378));
    layer6_outputs(1210) <= not((layer5_outputs(263)) and (layer5_outputs(2061)));
    layer6_outputs(1211) <= (layer5_outputs(3863)) and (layer5_outputs(953));
    layer6_outputs(1212) <= not((layer5_outputs(2199)) xor (layer5_outputs(177)));
    layer6_outputs(1213) <= not(layer5_outputs(466)) or (layer5_outputs(646));
    layer6_outputs(1214) <= not((layer5_outputs(457)) xor (layer5_outputs(4470)));
    layer6_outputs(1215) <= not((layer5_outputs(4539)) and (layer5_outputs(3970)));
    layer6_outputs(1216) <= not(layer5_outputs(3231));
    layer6_outputs(1217) <= layer5_outputs(2236);
    layer6_outputs(1218) <= '1';
    layer6_outputs(1219) <= (layer5_outputs(2499)) and (layer5_outputs(3225));
    layer6_outputs(1220) <= not((layer5_outputs(1060)) xor (layer5_outputs(2531)));
    layer6_outputs(1221) <= (layer5_outputs(3821)) and not (layer5_outputs(1418));
    layer6_outputs(1222) <= layer5_outputs(2386);
    layer6_outputs(1223) <= (layer5_outputs(2291)) and not (layer5_outputs(4112));
    layer6_outputs(1224) <= not(layer5_outputs(2112));
    layer6_outputs(1225) <= not(layer5_outputs(105));
    layer6_outputs(1226) <= not(layer5_outputs(3121));
    layer6_outputs(1227) <= not(layer5_outputs(1626));
    layer6_outputs(1228) <= '0';
    layer6_outputs(1229) <= not(layer5_outputs(5065));
    layer6_outputs(1230) <= not((layer5_outputs(1907)) or (layer5_outputs(59)));
    layer6_outputs(1231) <= (layer5_outputs(2174)) and (layer5_outputs(4160));
    layer6_outputs(1232) <= not((layer5_outputs(4834)) or (layer5_outputs(3190)));
    layer6_outputs(1233) <= (layer5_outputs(3028)) xor (layer5_outputs(2785));
    layer6_outputs(1234) <= layer5_outputs(810);
    layer6_outputs(1235) <= layer5_outputs(2664);
    layer6_outputs(1236) <= not((layer5_outputs(2216)) or (layer5_outputs(2362)));
    layer6_outputs(1237) <= (layer5_outputs(3203)) and (layer5_outputs(1245));
    layer6_outputs(1238) <= not((layer5_outputs(3994)) and (layer5_outputs(3396)));
    layer6_outputs(1239) <= not(layer5_outputs(71));
    layer6_outputs(1240) <= not((layer5_outputs(1889)) xor (layer5_outputs(4105)));
    layer6_outputs(1241) <= not((layer5_outputs(4861)) or (layer5_outputs(413)));
    layer6_outputs(1242) <= not((layer5_outputs(2510)) or (layer5_outputs(1380)));
    layer6_outputs(1243) <= not(layer5_outputs(1780));
    layer6_outputs(1244) <= not(layer5_outputs(3065));
    layer6_outputs(1245) <= layer5_outputs(1431);
    layer6_outputs(1246) <= not(layer5_outputs(3828)) or (layer5_outputs(1256));
    layer6_outputs(1247) <= layer5_outputs(2225);
    layer6_outputs(1248) <= not(layer5_outputs(1902));
    layer6_outputs(1249) <= not(layer5_outputs(2876)) or (layer5_outputs(799));
    layer6_outputs(1250) <= layer5_outputs(576);
    layer6_outputs(1251) <= (layer5_outputs(1017)) and not (layer5_outputs(4843));
    layer6_outputs(1252) <= (layer5_outputs(4163)) xor (layer5_outputs(2863));
    layer6_outputs(1253) <= '1';
    layer6_outputs(1254) <= (layer5_outputs(92)) and not (layer5_outputs(790));
    layer6_outputs(1255) <= (layer5_outputs(659)) and not (layer5_outputs(1239));
    layer6_outputs(1256) <= not((layer5_outputs(2133)) or (layer5_outputs(2942)));
    layer6_outputs(1257) <= (layer5_outputs(2329)) and (layer5_outputs(747));
    layer6_outputs(1258) <= (layer5_outputs(4548)) and not (layer5_outputs(1410));
    layer6_outputs(1259) <= layer5_outputs(1117);
    layer6_outputs(1260) <= layer5_outputs(2159);
    layer6_outputs(1261) <= not((layer5_outputs(2383)) and (layer5_outputs(4839)));
    layer6_outputs(1262) <= layer5_outputs(1754);
    layer6_outputs(1263) <= (layer5_outputs(1337)) or (layer5_outputs(4906));
    layer6_outputs(1264) <= not((layer5_outputs(2390)) or (layer5_outputs(4329)));
    layer6_outputs(1265) <= (layer5_outputs(71)) and not (layer5_outputs(2115));
    layer6_outputs(1266) <= not(layer5_outputs(2182)) or (layer5_outputs(815));
    layer6_outputs(1267) <= layer5_outputs(2884);
    layer6_outputs(1268) <= layer5_outputs(124);
    layer6_outputs(1269) <= not(layer5_outputs(2700)) or (layer5_outputs(3366));
    layer6_outputs(1270) <= layer5_outputs(3678);
    layer6_outputs(1271) <= not(layer5_outputs(3132)) or (layer5_outputs(3748));
    layer6_outputs(1272) <= (layer5_outputs(278)) and not (layer5_outputs(136));
    layer6_outputs(1273) <= (layer5_outputs(1505)) and not (layer5_outputs(3628));
    layer6_outputs(1274) <= not(layer5_outputs(1486));
    layer6_outputs(1275) <= layer5_outputs(2073);
    layer6_outputs(1276) <= not((layer5_outputs(1480)) or (layer5_outputs(4319)));
    layer6_outputs(1277) <= (layer5_outputs(3081)) or (layer5_outputs(1041));
    layer6_outputs(1278) <= not(layer5_outputs(3897)) or (layer5_outputs(4524));
    layer6_outputs(1279) <= '0';
    layer6_outputs(1280) <= (layer5_outputs(4583)) or (layer5_outputs(3990));
    layer6_outputs(1281) <= (layer5_outputs(5046)) and not (layer5_outputs(1867));
    layer6_outputs(1282) <= (layer5_outputs(718)) and (layer5_outputs(746));
    layer6_outputs(1283) <= not((layer5_outputs(764)) or (layer5_outputs(4353)));
    layer6_outputs(1284) <= not(layer5_outputs(3133)) or (layer5_outputs(4874));
    layer6_outputs(1285) <= (layer5_outputs(2812)) and not (layer5_outputs(4900));
    layer6_outputs(1286) <= (layer5_outputs(4651)) and not (layer5_outputs(374));
    layer6_outputs(1287) <= layer5_outputs(76);
    layer6_outputs(1288) <= not(layer5_outputs(1482));
    layer6_outputs(1289) <= layer5_outputs(3647);
    layer6_outputs(1290) <= layer5_outputs(2996);
    layer6_outputs(1291) <= not(layer5_outputs(783)) or (layer5_outputs(1006));
    layer6_outputs(1292) <= (layer5_outputs(1892)) or (layer5_outputs(2913));
    layer6_outputs(1293) <= (layer5_outputs(3344)) and (layer5_outputs(982));
    layer6_outputs(1294) <= not(layer5_outputs(2277)) or (layer5_outputs(2937));
    layer6_outputs(1295) <= layer5_outputs(818);
    layer6_outputs(1296) <= not((layer5_outputs(4799)) and (layer5_outputs(560)));
    layer6_outputs(1297) <= layer5_outputs(2468);
    layer6_outputs(1298) <= layer5_outputs(3487);
    layer6_outputs(1299) <= (layer5_outputs(2349)) and not (layer5_outputs(1512));
    layer6_outputs(1300) <= not(layer5_outputs(3024)) or (layer5_outputs(3798));
    layer6_outputs(1301) <= not(layer5_outputs(259));
    layer6_outputs(1302) <= layer5_outputs(4288);
    layer6_outputs(1303) <= (layer5_outputs(3478)) and not (layer5_outputs(1146));
    layer6_outputs(1304) <= not(layer5_outputs(4655));
    layer6_outputs(1305) <= layer5_outputs(3359);
    layer6_outputs(1306) <= (layer5_outputs(4876)) and not (layer5_outputs(3838));
    layer6_outputs(1307) <= not(layer5_outputs(4284)) or (layer5_outputs(2417));
    layer6_outputs(1308) <= (layer5_outputs(3055)) and not (layer5_outputs(429));
    layer6_outputs(1309) <= not(layer5_outputs(4085));
    layer6_outputs(1310) <= (layer5_outputs(3176)) or (layer5_outputs(3871));
    layer6_outputs(1311) <= not((layer5_outputs(3724)) or (layer5_outputs(1759)));
    layer6_outputs(1312) <= not(layer5_outputs(2792));
    layer6_outputs(1313) <= layer5_outputs(3405);
    layer6_outputs(1314) <= (layer5_outputs(987)) or (layer5_outputs(212));
    layer6_outputs(1315) <= not(layer5_outputs(2325));
    layer6_outputs(1316) <= (layer5_outputs(1327)) and not (layer5_outputs(603));
    layer6_outputs(1317) <= not((layer5_outputs(3432)) xor (layer5_outputs(3286)));
    layer6_outputs(1318) <= layer5_outputs(3414);
    layer6_outputs(1319) <= not(layer5_outputs(2991)) or (layer5_outputs(1967));
    layer6_outputs(1320) <= not(layer5_outputs(3946)) or (layer5_outputs(2267));
    layer6_outputs(1321) <= layer5_outputs(744);
    layer6_outputs(1322) <= not((layer5_outputs(4446)) xor (layer5_outputs(3455)));
    layer6_outputs(1323) <= layer5_outputs(3722);
    layer6_outputs(1324) <= (layer5_outputs(4898)) and (layer5_outputs(1767));
    layer6_outputs(1325) <= not((layer5_outputs(1056)) or (layer5_outputs(1513)));
    layer6_outputs(1326) <= not((layer5_outputs(3779)) and (layer5_outputs(2419)));
    layer6_outputs(1327) <= layer5_outputs(2710);
    layer6_outputs(1328) <= (layer5_outputs(346)) and not (layer5_outputs(2464));
    layer6_outputs(1329) <= (layer5_outputs(2099)) and not (layer5_outputs(2609));
    layer6_outputs(1330) <= not((layer5_outputs(2269)) and (layer5_outputs(1861)));
    layer6_outputs(1331) <= layer5_outputs(522);
    layer6_outputs(1332) <= '0';
    layer6_outputs(1333) <= not((layer5_outputs(4961)) or (layer5_outputs(819)));
    layer6_outputs(1334) <= not(layer5_outputs(942));
    layer6_outputs(1335) <= not(layer5_outputs(1482));
    layer6_outputs(1336) <= (layer5_outputs(4012)) and not (layer5_outputs(1617));
    layer6_outputs(1337) <= layer5_outputs(1334);
    layer6_outputs(1338) <= '1';
    layer6_outputs(1339) <= not(layer5_outputs(4399));
    layer6_outputs(1340) <= not((layer5_outputs(2400)) or (layer5_outputs(1679)));
    layer6_outputs(1341) <= not(layer5_outputs(3496)) or (layer5_outputs(3855));
    layer6_outputs(1342) <= (layer5_outputs(2543)) xor (layer5_outputs(711));
    layer6_outputs(1343) <= (layer5_outputs(4255)) and not (layer5_outputs(3695));
    layer6_outputs(1344) <= '1';
    layer6_outputs(1345) <= layer5_outputs(4808);
    layer6_outputs(1346) <= not(layer5_outputs(5018));
    layer6_outputs(1347) <= not(layer5_outputs(882));
    layer6_outputs(1348) <= not(layer5_outputs(1610));
    layer6_outputs(1349) <= not((layer5_outputs(4008)) and (layer5_outputs(2989)));
    layer6_outputs(1350) <= not(layer5_outputs(1756));
    layer6_outputs(1351) <= (layer5_outputs(3511)) or (layer5_outputs(880));
    layer6_outputs(1352) <= not(layer5_outputs(739));
    layer6_outputs(1353) <= (layer5_outputs(2758)) or (layer5_outputs(732));
    layer6_outputs(1354) <= (layer5_outputs(2359)) xor (layer5_outputs(3518));
    layer6_outputs(1355) <= not((layer5_outputs(3008)) or (layer5_outputs(4660)));
    layer6_outputs(1356) <= not(layer5_outputs(3240));
    layer6_outputs(1357) <= '1';
    layer6_outputs(1358) <= (layer5_outputs(4189)) and not (layer5_outputs(728));
    layer6_outputs(1359) <= (layer5_outputs(2663)) or (layer5_outputs(144));
    layer6_outputs(1360) <= (layer5_outputs(1616)) xor (layer5_outputs(3508));
    layer6_outputs(1361) <= not((layer5_outputs(3491)) xor (layer5_outputs(3356)));
    layer6_outputs(1362) <= not(layer5_outputs(625)) or (layer5_outputs(1585));
    layer6_outputs(1363) <= not(layer5_outputs(4764));
    layer6_outputs(1364) <= not(layer5_outputs(1652));
    layer6_outputs(1365) <= (layer5_outputs(1682)) and not (layer5_outputs(1528));
    layer6_outputs(1366) <= not(layer5_outputs(3425));
    layer6_outputs(1367) <= not(layer5_outputs(3182));
    layer6_outputs(1368) <= '0';
    layer6_outputs(1369) <= layer5_outputs(360);
    layer6_outputs(1370) <= '1';
    layer6_outputs(1371) <= not((layer5_outputs(704)) xor (layer5_outputs(11)));
    layer6_outputs(1372) <= layer5_outputs(3921);
    layer6_outputs(1373) <= not((layer5_outputs(485)) and (layer5_outputs(3555)));
    layer6_outputs(1374) <= '0';
    layer6_outputs(1375) <= layer5_outputs(550);
    layer6_outputs(1376) <= not(layer5_outputs(2912)) or (layer5_outputs(4828));
    layer6_outputs(1377) <= not(layer5_outputs(4006));
    layer6_outputs(1378) <= not(layer5_outputs(1839));
    layer6_outputs(1379) <= not((layer5_outputs(601)) and (layer5_outputs(4048)));
    layer6_outputs(1380) <= layer5_outputs(2189);
    layer6_outputs(1381) <= (layer5_outputs(557)) or (layer5_outputs(4027));
    layer6_outputs(1382) <= not(layer5_outputs(2741)) or (layer5_outputs(970));
    layer6_outputs(1383) <= layer5_outputs(2091);
    layer6_outputs(1384) <= layer5_outputs(4937);
    layer6_outputs(1385) <= layer5_outputs(3447);
    layer6_outputs(1386) <= not(layer5_outputs(4464));
    layer6_outputs(1387) <= not(layer5_outputs(2641));
    layer6_outputs(1388) <= layer5_outputs(3048);
    layer6_outputs(1389) <= not((layer5_outputs(4709)) or (layer5_outputs(4678)));
    layer6_outputs(1390) <= layer5_outputs(1544);
    layer6_outputs(1391) <= not((layer5_outputs(3308)) or (layer5_outputs(1356)));
    layer6_outputs(1392) <= not((layer5_outputs(3918)) and (layer5_outputs(3802)));
    layer6_outputs(1393) <= not((layer5_outputs(1003)) or (layer5_outputs(1125)));
    layer6_outputs(1394) <= layer5_outputs(1841);
    layer6_outputs(1395) <= layer5_outputs(2634);
    layer6_outputs(1396) <= not((layer5_outputs(2050)) or (layer5_outputs(553)));
    layer6_outputs(1397) <= layer5_outputs(1328);
    layer6_outputs(1398) <= (layer5_outputs(3340)) and (layer5_outputs(2235));
    layer6_outputs(1399) <= not(layer5_outputs(2275));
    layer6_outputs(1400) <= layer5_outputs(539);
    layer6_outputs(1401) <= not(layer5_outputs(4621));
    layer6_outputs(1402) <= layer5_outputs(401);
    layer6_outputs(1403) <= not(layer5_outputs(4140)) or (layer5_outputs(2747));
    layer6_outputs(1404) <= not(layer5_outputs(2320));
    layer6_outputs(1405) <= '1';
    layer6_outputs(1406) <= not(layer5_outputs(178)) or (layer5_outputs(4252));
    layer6_outputs(1407) <= layer5_outputs(3869);
    layer6_outputs(1408) <= (layer5_outputs(5104)) and not (layer5_outputs(1774));
    layer6_outputs(1409) <= '0';
    layer6_outputs(1410) <= (layer5_outputs(3066)) and not (layer5_outputs(4310));
    layer6_outputs(1411) <= layer5_outputs(1678);
    layer6_outputs(1412) <= not((layer5_outputs(852)) xor (layer5_outputs(3634)));
    layer6_outputs(1413) <= layer5_outputs(2557);
    layer6_outputs(1414) <= not((layer5_outputs(2831)) and (layer5_outputs(1476)));
    layer6_outputs(1415) <= not(layer5_outputs(4033)) or (layer5_outputs(5093));
    layer6_outputs(1416) <= (layer5_outputs(1260)) xor (layer5_outputs(4226));
    layer6_outputs(1417) <= not((layer5_outputs(4468)) and (layer5_outputs(3632)));
    layer6_outputs(1418) <= layer5_outputs(131);
    layer6_outputs(1419) <= '0';
    layer6_outputs(1420) <= not(layer5_outputs(3262));
    layer6_outputs(1421) <= layer5_outputs(740);
    layer6_outputs(1422) <= not(layer5_outputs(1527));
    layer6_outputs(1423) <= not(layer5_outputs(1895)) or (layer5_outputs(136));
    layer6_outputs(1424) <= layer5_outputs(158);
    layer6_outputs(1425) <= not(layer5_outputs(230));
    layer6_outputs(1426) <= not(layer5_outputs(2990));
    layer6_outputs(1427) <= not(layer5_outputs(1924));
    layer6_outputs(1428) <= not((layer5_outputs(4686)) or (layer5_outputs(4637)));
    layer6_outputs(1429) <= not((layer5_outputs(4128)) xor (layer5_outputs(4070)));
    layer6_outputs(1430) <= not(layer5_outputs(4615));
    layer6_outputs(1431) <= (layer5_outputs(4298)) or (layer5_outputs(3716));
    layer6_outputs(1432) <= not(layer5_outputs(793));
    layer6_outputs(1433) <= (layer5_outputs(3010)) or (layer5_outputs(575));
    layer6_outputs(1434) <= layer5_outputs(4466);
    layer6_outputs(1435) <= not(layer5_outputs(4102)) or (layer5_outputs(2274));
    layer6_outputs(1436) <= (layer5_outputs(126)) and (layer5_outputs(2298));
    layer6_outputs(1437) <= layer5_outputs(2485);
    layer6_outputs(1438) <= not(layer5_outputs(4749));
    layer6_outputs(1439) <= (layer5_outputs(1973)) and not (layer5_outputs(2261));
    layer6_outputs(1440) <= '0';
    layer6_outputs(1441) <= not(layer5_outputs(4838));
    layer6_outputs(1442) <= not((layer5_outputs(2284)) or (layer5_outputs(2467)));
    layer6_outputs(1443) <= layer5_outputs(3087);
    layer6_outputs(1444) <= not((layer5_outputs(4065)) and (layer5_outputs(2240)));
    layer6_outputs(1445) <= layer5_outputs(1605);
    layer6_outputs(1446) <= layer5_outputs(1263);
    layer6_outputs(1447) <= not(layer5_outputs(3915)) or (layer5_outputs(685));
    layer6_outputs(1448) <= not(layer5_outputs(2915));
    layer6_outputs(1449) <= not(layer5_outputs(5090)) or (layer5_outputs(544));
    layer6_outputs(1450) <= (layer5_outputs(2801)) and not (layer5_outputs(36));
    layer6_outputs(1451) <= (layer5_outputs(574)) xor (layer5_outputs(3171));
    layer6_outputs(1452) <= not((layer5_outputs(4728)) and (layer5_outputs(3733)));
    layer6_outputs(1453) <= '1';
    layer6_outputs(1454) <= (layer5_outputs(1163)) and not (layer5_outputs(4129));
    layer6_outputs(1455) <= not(layer5_outputs(2007));
    layer6_outputs(1456) <= not(layer5_outputs(2871));
    layer6_outputs(1457) <= (layer5_outputs(1923)) and not (layer5_outputs(1389));
    layer6_outputs(1458) <= '1';
    layer6_outputs(1459) <= not(layer5_outputs(3565));
    layer6_outputs(1460) <= (layer5_outputs(3254)) and not (layer5_outputs(2983));
    layer6_outputs(1461) <= (layer5_outputs(4184)) or (layer5_outputs(4568));
    layer6_outputs(1462) <= (layer5_outputs(4383)) xor (layer5_outputs(2047));
    layer6_outputs(1463) <= layer5_outputs(3233);
    layer6_outputs(1464) <= not(layer5_outputs(4141));
    layer6_outputs(1465) <= layer5_outputs(2372);
    layer6_outputs(1466) <= not(layer5_outputs(3705));
    layer6_outputs(1467) <= (layer5_outputs(1949)) or (layer5_outputs(4735));
    layer6_outputs(1468) <= layer5_outputs(1352);
    layer6_outputs(1469) <= not((layer5_outputs(4840)) xor (layer5_outputs(4187)));
    layer6_outputs(1470) <= not(layer5_outputs(920));
    layer6_outputs(1471) <= layer5_outputs(467);
    layer6_outputs(1472) <= layer5_outputs(2032);
    layer6_outputs(1473) <= not((layer5_outputs(2173)) and (layer5_outputs(1694)));
    layer6_outputs(1474) <= (layer5_outputs(4512)) and not (layer5_outputs(1540));
    layer6_outputs(1475) <= (layer5_outputs(4162)) and not (layer5_outputs(4916));
    layer6_outputs(1476) <= (layer5_outputs(3316)) and not (layer5_outputs(2813));
    layer6_outputs(1477) <= (layer5_outputs(1216)) and not (layer5_outputs(5063));
    layer6_outputs(1478) <= (layer5_outputs(5007)) xor (layer5_outputs(1037));
    layer6_outputs(1479) <= '0';
    layer6_outputs(1480) <= not(layer5_outputs(2541)) or (layer5_outputs(731));
    layer6_outputs(1481) <= not(layer5_outputs(4408));
    layer6_outputs(1482) <= (layer5_outputs(429)) and not (layer5_outputs(180));
    layer6_outputs(1483) <= not(layer5_outputs(2243)) or (layer5_outputs(3320));
    layer6_outputs(1484) <= layer5_outputs(2691);
    layer6_outputs(1485) <= layer5_outputs(3499);
    layer6_outputs(1486) <= not((layer5_outputs(2634)) and (layer5_outputs(1061)));
    layer6_outputs(1487) <= not(layer5_outputs(4802)) or (layer5_outputs(934));
    layer6_outputs(1488) <= not(layer5_outputs(2758));
    layer6_outputs(1489) <= not(layer5_outputs(3398));
    layer6_outputs(1490) <= not(layer5_outputs(2009));
    layer6_outputs(1491) <= '1';
    layer6_outputs(1492) <= not(layer5_outputs(564));
    layer6_outputs(1493) <= not((layer5_outputs(453)) or (layer5_outputs(3258)));
    layer6_outputs(1494) <= (layer5_outputs(1947)) and not (layer5_outputs(3269));
    layer6_outputs(1495) <= not(layer5_outputs(729));
    layer6_outputs(1496) <= '0';
    layer6_outputs(1497) <= not((layer5_outputs(3872)) xor (layer5_outputs(2328)));
    layer6_outputs(1498) <= (layer5_outputs(3176)) or (layer5_outputs(4883));
    layer6_outputs(1499) <= not(layer5_outputs(870)) or (layer5_outputs(1858));
    layer6_outputs(1500) <= not(layer5_outputs(1832)) or (layer5_outputs(3652));
    layer6_outputs(1501) <= (layer5_outputs(249)) xor (layer5_outputs(3074));
    layer6_outputs(1502) <= '0';
    layer6_outputs(1503) <= layer5_outputs(157);
    layer6_outputs(1504) <= '1';
    layer6_outputs(1505) <= not(layer5_outputs(3026));
    layer6_outputs(1506) <= (layer5_outputs(2866)) and (layer5_outputs(4447));
    layer6_outputs(1507) <= not(layer5_outputs(815));
    layer6_outputs(1508) <= not(layer5_outputs(964));
    layer6_outputs(1509) <= not(layer5_outputs(271));
    layer6_outputs(1510) <= not(layer5_outputs(109));
    layer6_outputs(1511) <= not(layer5_outputs(4430));
    layer6_outputs(1512) <= not(layer5_outputs(1978)) or (layer5_outputs(330));
    layer6_outputs(1513) <= not((layer5_outputs(4864)) and (layer5_outputs(4219)));
    layer6_outputs(1514) <= not(layer5_outputs(3027));
    layer6_outputs(1515) <= (layer5_outputs(482)) and not (layer5_outputs(758));
    layer6_outputs(1516) <= not(layer5_outputs(4837));
    layer6_outputs(1517) <= layer5_outputs(3391);
    layer6_outputs(1518) <= not(layer5_outputs(1714)) or (layer5_outputs(1499));
    layer6_outputs(1519) <= (layer5_outputs(3606)) and (layer5_outputs(3455));
    layer6_outputs(1520) <= (layer5_outputs(4540)) and (layer5_outputs(3813));
    layer6_outputs(1521) <= not(layer5_outputs(4716)) or (layer5_outputs(423));
    layer6_outputs(1522) <= (layer5_outputs(2838)) and (layer5_outputs(2484));
    layer6_outputs(1523) <= not(layer5_outputs(3229));
    layer6_outputs(1524) <= layer5_outputs(16);
    layer6_outputs(1525) <= (layer5_outputs(2778)) xor (layer5_outputs(1231));
    layer6_outputs(1526) <= '0';
    layer6_outputs(1527) <= '1';
    layer6_outputs(1528) <= layer5_outputs(3292);
    layer6_outputs(1529) <= not(layer5_outputs(4770)) or (layer5_outputs(4584));
    layer6_outputs(1530) <= not(layer5_outputs(502));
    layer6_outputs(1531) <= layer5_outputs(4286);
    layer6_outputs(1532) <= layer5_outputs(4143);
    layer6_outputs(1533) <= layer5_outputs(3524);
    layer6_outputs(1534) <= (layer5_outputs(4871)) xor (layer5_outputs(3728));
    layer6_outputs(1535) <= not(layer5_outputs(2761));
    layer6_outputs(1536) <= (layer5_outputs(5058)) and not (layer5_outputs(4547));
    layer6_outputs(1537) <= layer5_outputs(1248);
    layer6_outputs(1538) <= layer5_outputs(842);
    layer6_outputs(1539) <= not(layer5_outputs(498)) or (layer5_outputs(601));
    layer6_outputs(1540) <= (layer5_outputs(242)) xor (layer5_outputs(3906));
    layer6_outputs(1541) <= not(layer5_outputs(2029)) or (layer5_outputs(3115));
    layer6_outputs(1542) <= not(layer5_outputs(3964));
    layer6_outputs(1543) <= (layer5_outputs(679)) or (layer5_outputs(3940));
    layer6_outputs(1544) <= not((layer5_outputs(2102)) or (layer5_outputs(3987)));
    layer6_outputs(1545) <= (layer5_outputs(3930)) and (layer5_outputs(922));
    layer6_outputs(1546) <= not(layer5_outputs(3474)) or (layer5_outputs(3058));
    layer6_outputs(1547) <= (layer5_outputs(4764)) and (layer5_outputs(1655));
    layer6_outputs(1548) <= not((layer5_outputs(670)) or (layer5_outputs(1676)));
    layer6_outputs(1549) <= (layer5_outputs(2833)) and not (layer5_outputs(2887));
    layer6_outputs(1550) <= layer5_outputs(2286);
    layer6_outputs(1551) <= not(layer5_outputs(3354));
    layer6_outputs(1552) <= layer5_outputs(346);
    layer6_outputs(1553) <= not((layer5_outputs(1533)) and (layer5_outputs(674)));
    layer6_outputs(1554) <= (layer5_outputs(1350)) and (layer5_outputs(3983));
    layer6_outputs(1555) <= layer5_outputs(171);
    layer6_outputs(1556) <= layer5_outputs(3867);
    layer6_outputs(1557) <= not(layer5_outputs(2743));
    layer6_outputs(1558) <= (layer5_outputs(2930)) xor (layer5_outputs(3604));
    layer6_outputs(1559) <= layer5_outputs(2780);
    layer6_outputs(1560) <= not((layer5_outputs(5052)) or (layer5_outputs(663)));
    layer6_outputs(1561) <= layer5_outputs(2500);
    layer6_outputs(1562) <= not(layer5_outputs(1398)) or (layer5_outputs(5085));
    layer6_outputs(1563) <= '1';
    layer6_outputs(1564) <= '0';
    layer6_outputs(1565) <= not(layer5_outputs(2640));
    layer6_outputs(1566) <= layer5_outputs(167);
    layer6_outputs(1567) <= not(layer5_outputs(1048));
    layer6_outputs(1568) <= not((layer5_outputs(943)) or (layer5_outputs(3329)));
    layer6_outputs(1569) <= (layer5_outputs(1509)) and not (layer5_outputs(104));
    layer6_outputs(1570) <= (layer5_outputs(2196)) xor (layer5_outputs(4436));
    layer6_outputs(1571) <= (layer5_outputs(2416)) or (layer5_outputs(568));
    layer6_outputs(1572) <= '0';
    layer6_outputs(1573) <= not((layer5_outputs(2507)) xor (layer5_outputs(3132)));
    layer6_outputs(1574) <= (layer5_outputs(2021)) and (layer5_outputs(3243));
    layer6_outputs(1575) <= (layer5_outputs(1868)) or (layer5_outputs(2027));
    layer6_outputs(1576) <= not(layer5_outputs(2849)) or (layer5_outputs(2178));
    layer6_outputs(1577) <= layer5_outputs(2393);
    layer6_outputs(1578) <= layer5_outputs(4989);
    layer6_outputs(1579) <= '1';
    layer6_outputs(1580) <= not(layer5_outputs(784));
    layer6_outputs(1581) <= not((layer5_outputs(1233)) and (layer5_outputs(813)));
    layer6_outputs(1582) <= (layer5_outputs(1349)) or (layer5_outputs(3894));
    layer6_outputs(1583) <= layer5_outputs(190);
    layer6_outputs(1584) <= (layer5_outputs(3764)) or (layer5_outputs(2697));
    layer6_outputs(1585) <= layer5_outputs(4881);
    layer6_outputs(1586) <= not(layer5_outputs(259));
    layer6_outputs(1587) <= not((layer5_outputs(5062)) and (layer5_outputs(3997)));
    layer6_outputs(1588) <= not((layer5_outputs(4107)) or (layer5_outputs(4483)));
    layer6_outputs(1589) <= not(layer5_outputs(1115)) or (layer5_outputs(3705));
    layer6_outputs(1590) <= (layer5_outputs(1445)) and not (layer5_outputs(618));
    layer6_outputs(1591) <= '1';
    layer6_outputs(1592) <= not(layer5_outputs(2602)) or (layer5_outputs(4010));
    layer6_outputs(1593) <= not((layer5_outputs(3713)) xor (layer5_outputs(3907)));
    layer6_outputs(1594) <= not(layer5_outputs(2584)) or (layer5_outputs(4597));
    layer6_outputs(1595) <= (layer5_outputs(632)) and (layer5_outputs(534));
    layer6_outputs(1596) <= layer5_outputs(4199);
    layer6_outputs(1597) <= not(layer5_outputs(983));
    layer6_outputs(1598) <= not(layer5_outputs(3873)) or (layer5_outputs(2828));
    layer6_outputs(1599) <= not((layer5_outputs(1364)) and (layer5_outputs(3787)));
    layer6_outputs(1600) <= not(layer5_outputs(3717)) or (layer5_outputs(2397));
    layer6_outputs(1601) <= (layer5_outputs(715)) and not (layer5_outputs(755));
    layer6_outputs(1602) <= not((layer5_outputs(4188)) and (layer5_outputs(4885)));
    layer6_outputs(1603) <= '1';
    layer6_outputs(1604) <= (layer5_outputs(558)) or (layer5_outputs(4780));
    layer6_outputs(1605) <= (layer5_outputs(2411)) and (layer5_outputs(2153));
    layer6_outputs(1606) <= not(layer5_outputs(4201));
    layer6_outputs(1607) <= layer5_outputs(2146);
    layer6_outputs(1608) <= layer5_outputs(4418);
    layer6_outputs(1609) <= (layer5_outputs(2978)) and (layer5_outputs(2104));
    layer6_outputs(1610) <= not((layer5_outputs(77)) or (layer5_outputs(1295)));
    layer6_outputs(1611) <= not(layer5_outputs(4761)) or (layer5_outputs(675));
    layer6_outputs(1612) <= not(layer5_outputs(1134));
    layer6_outputs(1613) <= (layer5_outputs(5040)) and (layer5_outputs(106));
    layer6_outputs(1614) <= (layer5_outputs(1354)) and (layer5_outputs(1806));
    layer6_outputs(1615) <= (layer5_outputs(1956)) and not (layer5_outputs(885));
    layer6_outputs(1616) <= (layer5_outputs(262)) and (layer5_outputs(3843));
    layer6_outputs(1617) <= (layer5_outputs(3339)) or (layer5_outputs(4641));
    layer6_outputs(1618) <= not(layer5_outputs(4445));
    layer6_outputs(1619) <= not(layer5_outputs(487));
    layer6_outputs(1620) <= not(layer5_outputs(4805));
    layer6_outputs(1621) <= layer5_outputs(1291);
    layer6_outputs(1622) <= layer5_outputs(506);
    layer6_outputs(1623) <= (layer5_outputs(3647)) and (layer5_outputs(1153));
    layer6_outputs(1624) <= not(layer5_outputs(1782));
    layer6_outputs(1625) <= (layer5_outputs(796)) and (layer5_outputs(1823));
    layer6_outputs(1626) <= layer5_outputs(677);
    layer6_outputs(1627) <= '1';
    layer6_outputs(1628) <= (layer5_outputs(3188)) and (layer5_outputs(459));
    layer6_outputs(1629) <= (layer5_outputs(694)) and not (layer5_outputs(4548));
    layer6_outputs(1630) <= not(layer5_outputs(661));
    layer6_outputs(1631) <= (layer5_outputs(3775)) and (layer5_outputs(4520));
    layer6_outputs(1632) <= '1';
    layer6_outputs(1633) <= layer5_outputs(1699);
    layer6_outputs(1634) <= not((layer5_outputs(1299)) or (layer5_outputs(3049)));
    layer6_outputs(1635) <= not(layer5_outputs(4795)) or (layer5_outputs(4384));
    layer6_outputs(1636) <= (layer5_outputs(300)) or (layer5_outputs(1028));
    layer6_outputs(1637) <= (layer5_outputs(860)) and not (layer5_outputs(231));
    layer6_outputs(1638) <= not((layer5_outputs(2134)) or (layer5_outputs(359)));
    layer6_outputs(1639) <= not(layer5_outputs(4506));
    layer6_outputs(1640) <= (layer5_outputs(3645)) and (layer5_outputs(4389));
    layer6_outputs(1641) <= not((layer5_outputs(5067)) or (layer5_outputs(4202)));
    layer6_outputs(1642) <= layer5_outputs(128);
    layer6_outputs(1643) <= (layer5_outputs(1255)) and not (layer5_outputs(4706));
    layer6_outputs(1644) <= (layer5_outputs(114)) xor (layer5_outputs(3894));
    layer6_outputs(1645) <= '0';
    layer6_outputs(1646) <= not(layer5_outputs(3914));
    layer6_outputs(1647) <= layer5_outputs(4048);
    layer6_outputs(1648) <= not((layer5_outputs(1497)) xor (layer5_outputs(2401)));
    layer6_outputs(1649) <= layer5_outputs(2647);
    layer6_outputs(1650) <= not(layer5_outputs(2519)) or (layer5_outputs(3683));
    layer6_outputs(1651) <= (layer5_outputs(2371)) or (layer5_outputs(2805));
    layer6_outputs(1652) <= not((layer5_outputs(5004)) and (layer5_outputs(591)));
    layer6_outputs(1653) <= (layer5_outputs(596)) xor (layer5_outputs(4354));
    layer6_outputs(1654) <= (layer5_outputs(336)) and not (layer5_outputs(2581));
    layer6_outputs(1655) <= '1';
    layer6_outputs(1656) <= layer5_outputs(1589);
    layer6_outputs(1657) <= '0';
    layer6_outputs(1658) <= layer5_outputs(159);
    layer6_outputs(1659) <= (layer5_outputs(3559)) and (layer5_outputs(3585));
    layer6_outputs(1660) <= not(layer5_outputs(3244));
    layer6_outputs(1661) <= not(layer5_outputs(2515)) or (layer5_outputs(3836));
    layer6_outputs(1662) <= not(layer5_outputs(4858));
    layer6_outputs(1663) <= not(layer5_outputs(3428)) or (layer5_outputs(4082));
    layer6_outputs(1664) <= not(layer5_outputs(3402)) or (layer5_outputs(3832));
    layer6_outputs(1665) <= layer5_outputs(573);
    layer6_outputs(1666) <= (layer5_outputs(4245)) xor (layer5_outputs(886));
    layer6_outputs(1667) <= not(layer5_outputs(1836));
    layer6_outputs(1668) <= layer5_outputs(1918);
    layer6_outputs(1669) <= not((layer5_outputs(1051)) or (layer5_outputs(6)));
    layer6_outputs(1670) <= layer5_outputs(3893);
    layer6_outputs(1671) <= '1';
    layer6_outputs(1672) <= (layer5_outputs(623)) and not (layer5_outputs(959));
    layer6_outputs(1673) <= not(layer5_outputs(1002));
    layer6_outputs(1674) <= not(layer5_outputs(1936)) or (layer5_outputs(3519));
    layer6_outputs(1675) <= layer5_outputs(1888);
    layer6_outputs(1676) <= (layer5_outputs(1936)) and not (layer5_outputs(212));
    layer6_outputs(1677) <= not(layer5_outputs(5118));
    layer6_outputs(1678) <= not(layer5_outputs(2928)) or (layer5_outputs(4387));
    layer6_outputs(1679) <= not(layer5_outputs(4490));
    layer6_outputs(1680) <= (layer5_outputs(441)) and not (layer5_outputs(1151));
    layer6_outputs(1681) <= layer5_outputs(5004);
    layer6_outputs(1682) <= layer5_outputs(4618);
    layer6_outputs(1683) <= not((layer5_outputs(4891)) and (layer5_outputs(2231)));
    layer6_outputs(1684) <= layer5_outputs(4393);
    layer6_outputs(1685) <= not(layer5_outputs(3965)) or (layer5_outputs(407));
    layer6_outputs(1686) <= not(layer5_outputs(2406)) or (layer5_outputs(2937));
    layer6_outputs(1687) <= '0';
    layer6_outputs(1688) <= not((layer5_outputs(2774)) and (layer5_outputs(906)));
    layer6_outputs(1689) <= '1';
    layer6_outputs(1690) <= not((layer5_outputs(2223)) xor (layer5_outputs(1624)));
    layer6_outputs(1691) <= not(layer5_outputs(2710));
    layer6_outputs(1692) <= not((layer5_outputs(2476)) or (layer5_outputs(3682)));
    layer6_outputs(1693) <= not(layer5_outputs(4406));
    layer6_outputs(1694) <= not(layer5_outputs(4622)) or (layer5_outputs(1628));
    layer6_outputs(1695) <= not(layer5_outputs(3145));
    layer6_outputs(1696) <= layer5_outputs(1443);
    layer6_outputs(1697) <= layer5_outputs(4929);
    layer6_outputs(1698) <= not((layer5_outputs(993)) and (layer5_outputs(2430)));
    layer6_outputs(1699) <= layer5_outputs(3208);
    layer6_outputs(1700) <= layer5_outputs(2212);
    layer6_outputs(1701) <= not((layer5_outputs(2103)) and (layer5_outputs(1966)));
    layer6_outputs(1702) <= not(layer5_outputs(617));
    layer6_outputs(1703) <= layer5_outputs(3848);
    layer6_outputs(1704) <= not((layer5_outputs(933)) xor (layer5_outputs(3138)));
    layer6_outputs(1705) <= layer5_outputs(5102);
    layer6_outputs(1706) <= (layer5_outputs(4613)) and not (layer5_outputs(25));
    layer6_outputs(1707) <= not(layer5_outputs(1040)) or (layer5_outputs(851));
    layer6_outputs(1708) <= not(layer5_outputs(3104));
    layer6_outputs(1709) <= '1';
    layer6_outputs(1710) <= not(layer5_outputs(754));
    layer6_outputs(1711) <= (layer5_outputs(4234)) xor (layer5_outputs(4734));
    layer6_outputs(1712) <= not(layer5_outputs(5100));
    layer6_outputs(1713) <= not(layer5_outputs(3854)) or (layer5_outputs(4487));
    layer6_outputs(1714) <= layer5_outputs(3845);
    layer6_outputs(1715) <= not(layer5_outputs(2248)) or (layer5_outputs(2469));
    layer6_outputs(1716) <= not(layer5_outputs(3352));
    layer6_outputs(1717) <= layer5_outputs(4216);
    layer6_outputs(1718) <= not((layer5_outputs(4125)) xor (layer5_outputs(5076)));
    layer6_outputs(1719) <= not((layer5_outputs(483)) and (layer5_outputs(4610)));
    layer6_outputs(1720) <= '0';
    layer6_outputs(1721) <= layer5_outputs(464);
    layer6_outputs(1722) <= not((layer5_outputs(337)) and (layer5_outputs(2181)));
    layer6_outputs(1723) <= '0';
    layer6_outputs(1724) <= (layer5_outputs(3844)) or (layer5_outputs(1755));
    layer6_outputs(1725) <= '0';
    layer6_outputs(1726) <= not(layer5_outputs(2537));
    layer6_outputs(1727) <= not(layer5_outputs(4321));
    layer6_outputs(1728) <= layer5_outputs(4854);
    layer6_outputs(1729) <= not(layer5_outputs(2458)) or (layer5_outputs(2676));
    layer6_outputs(1730) <= layer5_outputs(628);
    layer6_outputs(1731) <= not(layer5_outputs(4145)) or (layer5_outputs(736));
    layer6_outputs(1732) <= '0';
    layer6_outputs(1733) <= layer5_outputs(4690);
    layer6_outputs(1734) <= not(layer5_outputs(939));
    layer6_outputs(1735) <= not(layer5_outputs(4916));
    layer6_outputs(1736) <= (layer5_outputs(2696)) and not (layer5_outputs(2471));
    layer6_outputs(1737) <= layer5_outputs(233);
    layer6_outputs(1738) <= not((layer5_outputs(4584)) or (layer5_outputs(1110)));
    layer6_outputs(1739) <= layer5_outputs(1937);
    layer6_outputs(1740) <= not(layer5_outputs(3898)) or (layer5_outputs(2267));
    layer6_outputs(1741) <= layer5_outputs(1560);
    layer6_outputs(1742) <= not(layer5_outputs(839));
    layer6_outputs(1743) <= not((layer5_outputs(4670)) or (layer5_outputs(4533)));
    layer6_outputs(1744) <= not((layer5_outputs(2266)) xor (layer5_outputs(1534)));
    layer6_outputs(1745) <= not(layer5_outputs(1668)) or (layer5_outputs(1197));
    layer6_outputs(1746) <= (layer5_outputs(2966)) or (layer5_outputs(4410));
    layer6_outputs(1747) <= not(layer5_outputs(4632));
    layer6_outputs(1748) <= not((layer5_outputs(3922)) and (layer5_outputs(2152)));
    layer6_outputs(1749) <= layer5_outputs(1419);
    layer6_outputs(1750) <= not((layer5_outputs(2358)) or (layer5_outputs(2299)));
    layer6_outputs(1751) <= layer5_outputs(260);
    layer6_outputs(1752) <= layer5_outputs(963);
    layer6_outputs(1753) <= not((layer5_outputs(2053)) xor (layer5_outputs(4746)));
    layer6_outputs(1754) <= layer5_outputs(2103);
    layer6_outputs(1755) <= '0';
    layer6_outputs(1756) <= not(layer5_outputs(4638));
    layer6_outputs(1757) <= not(layer5_outputs(198));
    layer6_outputs(1758) <= not((layer5_outputs(3099)) or (layer5_outputs(46)));
    layer6_outputs(1759) <= not(layer5_outputs(2743));
    layer6_outputs(1760) <= not(layer5_outputs(4697));
    layer6_outputs(1761) <= layer5_outputs(2672);
    layer6_outputs(1762) <= (layer5_outputs(3441)) and (layer5_outputs(614));
    layer6_outputs(1763) <= (layer5_outputs(2946)) and not (layer5_outputs(2242));
    layer6_outputs(1764) <= '1';
    layer6_outputs(1765) <= not(layer5_outputs(2496)) or (layer5_outputs(4555));
    layer6_outputs(1766) <= layer5_outputs(3467);
    layer6_outputs(1767) <= not(layer5_outputs(1414));
    layer6_outputs(1768) <= not(layer5_outputs(3509));
    layer6_outputs(1769) <= not(layer5_outputs(4602)) or (layer5_outputs(517));
    layer6_outputs(1770) <= not(layer5_outputs(655));
    layer6_outputs(1771) <= not((layer5_outputs(149)) or (layer5_outputs(3465)));
    layer6_outputs(1772) <= (layer5_outputs(1859)) or (layer5_outputs(810));
    layer6_outputs(1773) <= layer5_outputs(183);
    layer6_outputs(1774) <= not((layer5_outputs(817)) and (layer5_outputs(1370)));
    layer6_outputs(1775) <= not(layer5_outputs(3054));
    layer6_outputs(1776) <= not(layer5_outputs(765));
    layer6_outputs(1777) <= (layer5_outputs(4705)) and (layer5_outputs(2227));
    layer6_outputs(1778) <= layer5_outputs(4178);
    layer6_outputs(1779) <= layer5_outputs(548);
    layer6_outputs(1780) <= not(layer5_outputs(1443));
    layer6_outputs(1781) <= (layer5_outputs(986)) or (layer5_outputs(2341));
    layer6_outputs(1782) <= not(layer5_outputs(4921));
    layer6_outputs(1783) <= '1';
    layer6_outputs(1784) <= layer5_outputs(3047);
    layer6_outputs(1785) <= not((layer5_outputs(4750)) or (layer5_outputs(2297)));
    layer6_outputs(1786) <= not(layer5_outputs(1766)) or (layer5_outputs(2579));
    layer6_outputs(1787) <= layer5_outputs(4396);
    layer6_outputs(1788) <= not(layer5_outputs(2780)) or (layer5_outputs(4626));
    layer6_outputs(1789) <= not(layer5_outputs(3492));
    layer6_outputs(1790) <= layer5_outputs(2592);
    layer6_outputs(1791) <= layer5_outputs(3725);
    layer6_outputs(1792) <= layer5_outputs(1025);
    layer6_outputs(1793) <= layer5_outputs(4395);
    layer6_outputs(1794) <= (layer5_outputs(738)) and not (layer5_outputs(928));
    layer6_outputs(1795) <= '0';
    layer6_outputs(1796) <= not(layer5_outputs(2052));
    layer6_outputs(1797) <= not(layer5_outputs(1423));
    layer6_outputs(1798) <= not(layer5_outputs(1650));
    layer6_outputs(1799) <= (layer5_outputs(2558)) and not (layer5_outputs(1333));
    layer6_outputs(1800) <= not(layer5_outputs(101));
    layer6_outputs(1801) <= not((layer5_outputs(3137)) or (layer5_outputs(0)));
    layer6_outputs(1802) <= '0';
    layer6_outputs(1803) <= not(layer5_outputs(1727));
    layer6_outputs(1804) <= (layer5_outputs(2054)) and not (layer5_outputs(2766));
    layer6_outputs(1805) <= not((layer5_outputs(2901)) and (layer5_outputs(3594)));
    layer6_outputs(1806) <= (layer5_outputs(4645)) xor (layer5_outputs(578));
    layer6_outputs(1807) <= not(layer5_outputs(2557));
    layer6_outputs(1808) <= layer5_outputs(1190);
    layer6_outputs(1809) <= layer5_outputs(3774);
    layer6_outputs(1810) <= not(layer5_outputs(4500));
    layer6_outputs(1811) <= (layer5_outputs(1185)) and not (layer5_outputs(2201));
    layer6_outputs(1812) <= not(layer5_outputs(4281));
    layer6_outputs(1813) <= not((layer5_outputs(2484)) xor (layer5_outputs(2099)));
    layer6_outputs(1814) <= (layer5_outputs(432)) or (layer5_outputs(3880));
    layer6_outputs(1815) <= '0';
    layer6_outputs(1816) <= not((layer5_outputs(915)) and (layer5_outputs(1595)));
    layer6_outputs(1817) <= '1';
    layer6_outputs(1818) <= (layer5_outputs(3146)) or (layer5_outputs(4077));
    layer6_outputs(1819) <= layer5_outputs(2768);
    layer6_outputs(1820) <= not(layer5_outputs(4438)) or (layer5_outputs(4719));
    layer6_outputs(1821) <= layer5_outputs(131);
    layer6_outputs(1822) <= not(layer5_outputs(4246));
    layer6_outputs(1823) <= layer5_outputs(733);
    layer6_outputs(1824) <= layer5_outputs(2949);
    layer6_outputs(1825) <= not((layer5_outputs(4666)) and (layer5_outputs(908)));
    layer6_outputs(1826) <= layer5_outputs(1754);
    layer6_outputs(1827) <= '0';
    layer6_outputs(1828) <= layer5_outputs(3950);
    layer6_outputs(1829) <= (layer5_outputs(2891)) and (layer5_outputs(2750));
    layer6_outputs(1830) <= '1';
    layer6_outputs(1831) <= not((layer5_outputs(4194)) or (layer5_outputs(2641)));
    layer6_outputs(1832) <= (layer5_outputs(3995)) xor (layer5_outputs(2032));
    layer6_outputs(1833) <= not(layer5_outputs(293));
    layer6_outputs(1834) <= layer5_outputs(1521);
    layer6_outputs(1835) <= not(layer5_outputs(4064)) or (layer5_outputs(584));
    layer6_outputs(1836) <= layer5_outputs(757);
    layer6_outputs(1837) <= not((layer5_outputs(1640)) or (layer5_outputs(142)));
    layer6_outputs(1838) <= not(layer5_outputs(837));
    layer6_outputs(1839) <= (layer5_outputs(90)) and not (layer5_outputs(5029));
    layer6_outputs(1840) <= layer5_outputs(3806);
    layer6_outputs(1841) <= '0';
    layer6_outputs(1842) <= layer5_outputs(3928);
    layer6_outputs(1843) <= not(layer5_outputs(376));
    layer6_outputs(1844) <= layer5_outputs(1335);
    layer6_outputs(1845) <= not(layer5_outputs(2351));
    layer6_outputs(1846) <= layer5_outputs(5048);
    layer6_outputs(1847) <= '1';
    layer6_outputs(1848) <= not((layer5_outputs(1461)) or (layer5_outputs(4038)));
    layer6_outputs(1849) <= not(layer5_outputs(3323));
    layer6_outputs(1850) <= not((layer5_outputs(2405)) or (layer5_outputs(3384)));
    layer6_outputs(1851) <= not(layer5_outputs(4167));
    layer6_outputs(1852) <= not(layer5_outputs(1449)) or (layer5_outputs(516));
    layer6_outputs(1853) <= layer5_outputs(2963);
    layer6_outputs(1854) <= (layer5_outputs(323)) and not (layer5_outputs(1104));
    layer6_outputs(1855) <= layer5_outputs(3667);
    layer6_outputs(1856) <= not(layer5_outputs(2847));
    layer6_outputs(1857) <= not(layer5_outputs(1673));
    layer6_outputs(1858) <= (layer5_outputs(380)) xor (layer5_outputs(1597));
    layer6_outputs(1859) <= (layer5_outputs(3126)) xor (layer5_outputs(526));
    layer6_outputs(1860) <= (layer5_outputs(2144)) and not (layer5_outputs(362));
    layer6_outputs(1861) <= (layer5_outputs(2305)) and (layer5_outputs(4000));
    layer6_outputs(1862) <= layer5_outputs(3497);
    layer6_outputs(1863) <= not(layer5_outputs(1231));
    layer6_outputs(1864) <= (layer5_outputs(2276)) and (layer5_outputs(2208));
    layer6_outputs(1865) <= not((layer5_outputs(2713)) and (layer5_outputs(5031)));
    layer6_outputs(1866) <= '0';
    layer6_outputs(1867) <= (layer5_outputs(1422)) and (layer5_outputs(531));
    layer6_outputs(1868) <= not(layer5_outputs(4719));
    layer6_outputs(1869) <= (layer5_outputs(615)) xor (layer5_outputs(173));
    layer6_outputs(1870) <= layer5_outputs(57);
    layer6_outputs(1871) <= (layer5_outputs(2331)) and not (layer5_outputs(3556));
    layer6_outputs(1872) <= '0';
    layer6_outputs(1873) <= layer5_outputs(4100);
    layer6_outputs(1874) <= not((layer5_outputs(5098)) and (layer5_outputs(3769)));
    layer6_outputs(1875) <= not(layer5_outputs(2296));
    layer6_outputs(1876) <= layer5_outputs(4552);
    layer6_outputs(1877) <= (layer5_outputs(113)) and (layer5_outputs(4898));
    layer6_outputs(1878) <= layer5_outputs(2490);
    layer6_outputs(1879) <= not(layer5_outputs(1666));
    layer6_outputs(1880) <= not(layer5_outputs(4326));
    layer6_outputs(1881) <= layer5_outputs(3846);
    layer6_outputs(1882) <= not(layer5_outputs(1503));
    layer6_outputs(1883) <= not(layer5_outputs(64));
    layer6_outputs(1884) <= not(layer5_outputs(2197));
    layer6_outputs(1885) <= not(layer5_outputs(2213));
    layer6_outputs(1886) <= not((layer5_outputs(2728)) and (layer5_outputs(777)));
    layer6_outputs(1887) <= (layer5_outputs(3901)) and not (layer5_outputs(437));
    layer6_outputs(1888) <= '1';
    layer6_outputs(1889) <= (layer5_outputs(4829)) and (layer5_outputs(347));
    layer6_outputs(1890) <= not((layer5_outputs(4241)) and (layer5_outputs(3322)));
    layer6_outputs(1891) <= (layer5_outputs(4904)) and not (layer5_outputs(3249));
    layer6_outputs(1892) <= layer5_outputs(2592);
    layer6_outputs(1893) <= not(layer5_outputs(3985));
    layer6_outputs(1894) <= not((layer5_outputs(4399)) xor (layer5_outputs(4789)));
    layer6_outputs(1895) <= not(layer5_outputs(5003));
    layer6_outputs(1896) <= not((layer5_outputs(4960)) xor (layer5_outputs(3514)));
    layer6_outputs(1897) <= layer5_outputs(3453);
    layer6_outputs(1898) <= layer5_outputs(515);
    layer6_outputs(1899) <= (layer5_outputs(5022)) xor (layer5_outputs(2723));
    layer6_outputs(1900) <= layer5_outputs(4392);
    layer6_outputs(1901) <= not(layer5_outputs(1080)) or (layer5_outputs(4867));
    layer6_outputs(1902) <= (layer5_outputs(232)) or (layer5_outputs(2544));
    layer6_outputs(1903) <= layer5_outputs(2363);
    layer6_outputs(1904) <= not((layer5_outputs(5021)) xor (layer5_outputs(1145)));
    layer6_outputs(1905) <= (layer5_outputs(1019)) and not (layer5_outputs(3042));
    layer6_outputs(1906) <= layer5_outputs(907);
    layer6_outputs(1907) <= not((layer5_outputs(2410)) or (layer5_outputs(919)));
    layer6_outputs(1908) <= not(layer5_outputs(3300));
    layer6_outputs(1909) <= not((layer5_outputs(56)) or (layer5_outputs(4052)));
    layer6_outputs(1910) <= (layer5_outputs(738)) and (layer5_outputs(2265));
    layer6_outputs(1911) <= not(layer5_outputs(2177)) or (layer5_outputs(4736));
    layer6_outputs(1912) <= (layer5_outputs(4007)) xor (layer5_outputs(178));
    layer6_outputs(1913) <= not((layer5_outputs(4136)) xor (layer5_outputs(3350)));
    layer6_outputs(1914) <= not((layer5_outputs(4316)) or (layer5_outputs(2817)));
    layer6_outputs(1915) <= layer5_outputs(2606);
    layer6_outputs(1916) <= (layer5_outputs(964)) and (layer5_outputs(3103));
    layer6_outputs(1917) <= not((layer5_outputs(287)) xor (layer5_outputs(3017)));
    layer6_outputs(1918) <= layer5_outputs(968);
    layer6_outputs(1919) <= layer5_outputs(2737);
    layer6_outputs(1920) <= layer5_outputs(876);
    layer6_outputs(1921) <= not((layer5_outputs(651)) or (layer5_outputs(3593)));
    layer6_outputs(1922) <= layer5_outputs(4267);
    layer6_outputs(1923) <= not(layer5_outputs(2932)) or (layer5_outputs(2178));
    layer6_outputs(1924) <= not((layer5_outputs(766)) or (layer5_outputs(3348)));
    layer6_outputs(1925) <= not(layer5_outputs(2019)) or (layer5_outputs(1046));
    layer6_outputs(1926) <= not(layer5_outputs(651));
    layer6_outputs(1927) <= layer5_outputs(1395);
    layer6_outputs(1928) <= not(layer5_outputs(4556));
    layer6_outputs(1929) <= layer5_outputs(963);
    layer6_outputs(1930) <= '0';
    layer6_outputs(1931) <= not((layer5_outputs(313)) or (layer5_outputs(3298)));
    layer6_outputs(1932) <= (layer5_outputs(3276)) xor (layer5_outputs(3431));
    layer6_outputs(1933) <= layer5_outputs(4976);
    layer6_outputs(1934) <= not(layer5_outputs(1893)) or (layer5_outputs(4403));
    layer6_outputs(1935) <= (layer5_outputs(1905)) xor (layer5_outputs(4817));
    layer6_outputs(1936) <= not(layer5_outputs(68));
    layer6_outputs(1937) <= not(layer5_outputs(4860));
    layer6_outputs(1938) <= not(layer5_outputs(1798));
    layer6_outputs(1939) <= layer5_outputs(4167);
    layer6_outputs(1940) <= not(layer5_outputs(4724));
    layer6_outputs(1941) <= not(layer5_outputs(4293));
    layer6_outputs(1942) <= not(layer5_outputs(1345));
    layer6_outputs(1943) <= layer5_outputs(2192);
    layer6_outputs(1944) <= not((layer5_outputs(770)) and (layer5_outputs(1440)));
    layer6_outputs(1945) <= not(layer5_outputs(1233)) or (layer5_outputs(3780));
    layer6_outputs(1946) <= not((layer5_outputs(2294)) or (layer5_outputs(2536)));
    layer6_outputs(1947) <= not((layer5_outputs(1825)) or (layer5_outputs(179)));
    layer6_outputs(1948) <= not(layer5_outputs(3098));
    layer6_outputs(1949) <= layer5_outputs(2775);
    layer6_outputs(1950) <= not((layer5_outputs(529)) xor (layer5_outputs(356)));
    layer6_outputs(1951) <= (layer5_outputs(199)) xor (layer5_outputs(674));
    layer6_outputs(1952) <= (layer5_outputs(3727)) and (layer5_outputs(411));
    layer6_outputs(1953) <= layer5_outputs(3706);
    layer6_outputs(1954) <= not((layer5_outputs(2010)) and (layer5_outputs(5059)));
    layer6_outputs(1955) <= not((layer5_outputs(4657)) and (layer5_outputs(2808)));
    layer6_outputs(1956) <= not((layer5_outputs(2157)) or (layer5_outputs(1985)));
    layer6_outputs(1957) <= (layer5_outputs(470)) or (layer5_outputs(1899));
    layer6_outputs(1958) <= (layer5_outputs(4691)) and (layer5_outputs(1311));
    layer6_outputs(1959) <= (layer5_outputs(4930)) xor (layer5_outputs(5068));
    layer6_outputs(1960) <= not((layer5_outputs(3173)) or (layer5_outputs(147)));
    layer6_outputs(1961) <= not(layer5_outputs(400));
    layer6_outputs(1962) <= '0';
    layer6_outputs(1963) <= not(layer5_outputs(2046));
    layer6_outputs(1964) <= layer5_outputs(3343);
    layer6_outputs(1965) <= not(layer5_outputs(416));
    layer6_outputs(1966) <= (layer5_outputs(4453)) and not (layer5_outputs(2846));
    layer6_outputs(1967) <= (layer5_outputs(462)) and not (layer5_outputs(378));
    layer6_outputs(1968) <= (layer5_outputs(2239)) or (layer5_outputs(240));
    layer6_outputs(1969) <= not(layer5_outputs(971));
    layer6_outputs(1970) <= layer5_outputs(3627);
    layer6_outputs(1971) <= not(layer5_outputs(4001));
    layer6_outputs(1972) <= (layer5_outputs(4375)) and not (layer5_outputs(3675));
    layer6_outputs(1973) <= not(layer5_outputs(1428));
    layer6_outputs(1974) <= not((layer5_outputs(3158)) xor (layer5_outputs(524)));
    layer6_outputs(1975) <= not((layer5_outputs(2819)) or (layer5_outputs(624)));
    layer6_outputs(1976) <= not(layer5_outputs(3395));
    layer6_outputs(1977) <= not(layer5_outputs(4222));
    layer6_outputs(1978) <= not(layer5_outputs(2027));
    layer6_outputs(1979) <= not((layer5_outputs(2941)) or (layer5_outputs(3743)));
    layer6_outputs(1980) <= not(layer5_outputs(93));
    layer6_outputs(1981) <= not(layer5_outputs(2453));
    layer6_outputs(1982) <= (layer5_outputs(4668)) and (layer5_outputs(2370));
    layer6_outputs(1983) <= not(layer5_outputs(194));
    layer6_outputs(1984) <= layer5_outputs(4057);
    layer6_outputs(1985) <= not(layer5_outputs(4833)) or (layer5_outputs(2341));
    layer6_outputs(1986) <= not(layer5_outputs(3916));
    layer6_outputs(1987) <= (layer5_outputs(2924)) or (layer5_outputs(1126));
    layer6_outputs(1988) <= not(layer5_outputs(3237));
    layer6_outputs(1989) <= not((layer5_outputs(772)) xor (layer5_outputs(350)));
    layer6_outputs(1990) <= '1';
    layer6_outputs(1991) <= (layer5_outputs(3174)) and (layer5_outputs(4330));
    layer6_outputs(1992) <= (layer5_outputs(1073)) and not (layer5_outputs(5001));
    layer6_outputs(1993) <= not(layer5_outputs(216));
    layer6_outputs(1994) <= (layer5_outputs(1425)) and not (layer5_outputs(2180));
    layer6_outputs(1995) <= '0';
    layer6_outputs(1996) <= (layer5_outputs(1157)) and (layer5_outputs(615));
    layer6_outputs(1997) <= '0';
    layer6_outputs(1998) <= '1';
    layer6_outputs(1999) <= not(layer5_outputs(2586)) or (layer5_outputs(4363));
    layer6_outputs(2000) <= not(layer5_outputs(1062));
    layer6_outputs(2001) <= not(layer5_outputs(3765)) or (layer5_outputs(2433));
    layer6_outputs(2002) <= not((layer5_outputs(3660)) or (layer5_outputs(4518)));
    layer6_outputs(2003) <= (layer5_outputs(367)) or (layer5_outputs(1043));
    layer6_outputs(2004) <= (layer5_outputs(2948)) and not (layer5_outputs(3502));
    layer6_outputs(2005) <= (layer5_outputs(3651)) and not (layer5_outputs(2452));
    layer6_outputs(2006) <= layer5_outputs(1808);
    layer6_outputs(2007) <= layer5_outputs(1124);
    layer6_outputs(2008) <= not((layer5_outputs(4104)) xor (layer5_outputs(3975)));
    layer6_outputs(2009) <= (layer5_outputs(1519)) and not (layer5_outputs(2654));
    layer6_outputs(2010) <= (layer5_outputs(2381)) and not (layer5_outputs(886));
    layer6_outputs(2011) <= (layer5_outputs(710)) or (layer5_outputs(931));
    layer6_outputs(2012) <= not((layer5_outputs(631)) xor (layer5_outputs(1882)));
    layer6_outputs(2013) <= not(layer5_outputs(1031));
    layer6_outputs(2014) <= not(layer5_outputs(1054));
    layer6_outputs(2015) <= not(layer5_outputs(1437)) or (layer5_outputs(3691));
    layer6_outputs(2016) <= layer5_outputs(3127);
    layer6_outputs(2017) <= not(layer5_outputs(2303)) or (layer5_outputs(977));
    layer6_outputs(2018) <= (layer5_outputs(4004)) and not (layer5_outputs(4549));
    layer6_outputs(2019) <= (layer5_outputs(291)) and not (layer5_outputs(2408));
    layer6_outputs(2020) <= layer5_outputs(4770);
    layer6_outputs(2021) <= not(layer5_outputs(2200)) or (layer5_outputs(3288));
    layer6_outputs(2022) <= (layer5_outputs(4614)) and not (layer5_outputs(4384));
    layer6_outputs(2023) <= (layer5_outputs(2062)) or (layer5_outputs(1874));
    layer6_outputs(2024) <= not(layer5_outputs(586));
    layer6_outputs(2025) <= not(layer5_outputs(7));
    layer6_outputs(2026) <= not(layer5_outputs(883)) or (layer5_outputs(903));
    layer6_outputs(2027) <= not(layer5_outputs(5092)) or (layer5_outputs(2281));
    layer6_outputs(2028) <= (layer5_outputs(2769)) and (layer5_outputs(4684));
    layer6_outputs(2029) <= (layer5_outputs(5018)) and not (layer5_outputs(1792));
    layer6_outputs(2030) <= layer5_outputs(2473);
    layer6_outputs(2031) <= layer5_outputs(1389);
    layer6_outputs(2032) <= not((layer5_outputs(227)) and (layer5_outputs(594)));
    layer6_outputs(2033) <= (layer5_outputs(3520)) and not (layer5_outputs(2176));
    layer6_outputs(2034) <= layer5_outputs(1156);
    layer6_outputs(2035) <= not((layer5_outputs(670)) xor (layer5_outputs(1283)));
    layer6_outputs(2036) <= '0';
    layer6_outputs(2037) <= (layer5_outputs(2092)) and not (layer5_outputs(1618));
    layer6_outputs(2038) <= layer5_outputs(5112);
    layer6_outputs(2039) <= (layer5_outputs(4029)) and (layer5_outputs(4539));
    layer6_outputs(2040) <= not(layer5_outputs(3256)) or (layer5_outputs(1269));
    layer6_outputs(2041) <= not(layer5_outputs(325)) or (layer5_outputs(53));
    layer6_outputs(2042) <= layer5_outputs(3500);
    layer6_outputs(2043) <= layer5_outputs(308);
    layer6_outputs(2044) <= layer5_outputs(103);
    layer6_outputs(2045) <= layer5_outputs(1499);
    layer6_outputs(2046) <= '0';
    layer6_outputs(2047) <= layer5_outputs(2539);
    layer6_outputs(2048) <= not(layer5_outputs(1440));
    layer6_outputs(2049) <= (layer5_outputs(1393)) and not (layer5_outputs(3421));
    layer6_outputs(2050) <= layer5_outputs(5105);
    layer6_outputs(2051) <= not(layer5_outputs(1407));
    layer6_outputs(2052) <= not(layer5_outputs(4959)) or (layer5_outputs(4180));
    layer6_outputs(2053) <= not(layer5_outputs(1635)) or (layer5_outputs(1916));
    layer6_outputs(2054) <= not((layer5_outputs(835)) xor (layer5_outputs(897)));
    layer6_outputs(2055) <= not(layer5_outputs(3999));
    layer6_outputs(2056) <= not((layer5_outputs(72)) or (layer5_outputs(66)));
    layer6_outputs(2057) <= not(layer5_outputs(2313));
    layer6_outputs(2058) <= not(layer5_outputs(1557));
    layer6_outputs(2059) <= not((layer5_outputs(2324)) xor (layer5_outputs(4558)));
    layer6_outputs(2060) <= not(layer5_outputs(5022));
    layer6_outputs(2061) <= '0';
    layer6_outputs(2062) <= (layer5_outputs(1108)) xor (layer5_outputs(2150));
    layer6_outputs(2063) <= not(layer5_outputs(928));
    layer6_outputs(2064) <= '1';
    layer6_outputs(2065) <= (layer5_outputs(2462)) xor (layer5_outputs(1717));
    layer6_outputs(2066) <= (layer5_outputs(2832)) xor (layer5_outputs(3312));
    layer6_outputs(2067) <= layer5_outputs(4709);
    layer6_outputs(2068) <= not(layer5_outputs(541)) or (layer5_outputs(4932));
    layer6_outputs(2069) <= (layer5_outputs(3809)) and not (layer5_outputs(2350));
    layer6_outputs(2070) <= layer5_outputs(562);
    layer6_outputs(2071) <= (layer5_outputs(1142)) xor (layer5_outputs(1229));
    layer6_outputs(2072) <= layer5_outputs(1865);
    layer6_outputs(2073) <= layer5_outputs(1835);
    layer6_outputs(2074) <= not(layer5_outputs(3474));
    layer6_outputs(2075) <= not((layer5_outputs(1558)) xor (layer5_outputs(3360)));
    layer6_outputs(2076) <= (layer5_outputs(1031)) and not (layer5_outputs(1379));
    layer6_outputs(2077) <= layer5_outputs(4988);
    layer6_outputs(2078) <= not(layer5_outputs(1999));
    layer6_outputs(2079) <= not(layer5_outputs(1187)) or (layer5_outputs(1583));
    layer6_outputs(2080) <= layer5_outputs(213);
    layer6_outputs(2081) <= not(layer5_outputs(117));
    layer6_outputs(2082) <= layer5_outputs(1009);
    layer6_outputs(2083) <= not((layer5_outputs(2719)) and (layer5_outputs(3330)));
    layer6_outputs(2084) <= (layer5_outputs(4224)) and not (layer5_outputs(3134));
    layer6_outputs(2085) <= not((layer5_outputs(2782)) xor (layer5_outputs(4444)));
    layer6_outputs(2086) <= not(layer5_outputs(5024)) or (layer5_outputs(3826));
    layer6_outputs(2087) <= (layer5_outputs(4671)) and not (layer5_outputs(4036));
    layer6_outputs(2088) <= layer5_outputs(2815);
    layer6_outputs(2089) <= not(layer5_outputs(991));
    layer6_outputs(2090) <= not((layer5_outputs(2896)) or (layer5_outputs(3280)));
    layer6_outputs(2091) <= (layer5_outputs(1100)) and (layer5_outputs(3954));
    layer6_outputs(2092) <= not((layer5_outputs(3896)) xor (layer5_outputs(354)));
    layer6_outputs(2093) <= not((layer5_outputs(3588)) and (layer5_outputs(2637)));
    layer6_outputs(2094) <= (layer5_outputs(1349)) and (layer5_outputs(2969));
    layer6_outputs(2095) <= not((layer5_outputs(4794)) xor (layer5_outputs(3481)));
    layer6_outputs(2096) <= not(layer5_outputs(4689)) or (layer5_outputs(1702));
    layer6_outputs(2097) <= not((layer5_outputs(1102)) or (layer5_outputs(4492)));
    layer6_outputs(2098) <= layer5_outputs(2415);
    layer6_outputs(2099) <= layer5_outputs(1036);
    layer6_outputs(2100) <= (layer5_outputs(3267)) and not (layer5_outputs(3498));
    layer6_outputs(2101) <= (layer5_outputs(5029)) and not (layer5_outputs(633));
    layer6_outputs(2102) <= not((layer5_outputs(3846)) or (layer5_outputs(800)));
    layer6_outputs(2103) <= layer5_outputs(4217);
    layer6_outputs(2104) <= (layer5_outputs(4494)) and (layer5_outputs(5106));
    layer6_outputs(2105) <= not(layer5_outputs(396)) or (layer5_outputs(1326));
    layer6_outputs(2106) <= not(layer5_outputs(3482));
    layer6_outputs(2107) <= not(layer5_outputs(3621));
    layer6_outputs(2108) <= layer5_outputs(17);
    layer6_outputs(2109) <= (layer5_outputs(1058)) and not (layer5_outputs(1165));
    layer6_outputs(2110) <= layer5_outputs(4670);
    layer6_outputs(2111) <= layer5_outputs(3953);
    layer6_outputs(2112) <= layer5_outputs(4348);
    layer6_outputs(2113) <= (layer5_outputs(465)) or (layer5_outputs(2033));
    layer6_outputs(2114) <= not((layer5_outputs(5040)) and (layer5_outputs(1863)));
    layer6_outputs(2115) <= (layer5_outputs(3771)) and (layer5_outputs(2566));
    layer6_outputs(2116) <= layer5_outputs(1423);
    layer6_outputs(2117) <= not((layer5_outputs(4679)) and (layer5_outputs(4419)));
    layer6_outputs(2118) <= not(layer5_outputs(4779)) or (layer5_outputs(3905));
    layer6_outputs(2119) <= not((layer5_outputs(3446)) xor (layer5_outputs(4599)));
    layer6_outputs(2120) <= not(layer5_outputs(4673));
    layer6_outputs(2121) <= layer5_outputs(4267);
    layer6_outputs(2122) <= not(layer5_outputs(192));
    layer6_outputs(2123) <= not(layer5_outputs(994));
    layer6_outputs(2124) <= layer5_outputs(2724);
    layer6_outputs(2125) <= not(layer5_outputs(3473)) or (layer5_outputs(2223));
    layer6_outputs(2126) <= '0';
    layer6_outputs(2127) <= not((layer5_outputs(3817)) and (layer5_outputs(4876)));
    layer6_outputs(2128) <= not(layer5_outputs(1412));
    layer6_outputs(2129) <= layer5_outputs(902);
    layer6_outputs(2130) <= not(layer5_outputs(5051));
    layer6_outputs(2131) <= not(layer5_outputs(2579));
    layer6_outputs(2132) <= (layer5_outputs(3838)) and (layer5_outputs(4599));
    layer6_outputs(2133) <= not(layer5_outputs(1678));
    layer6_outputs(2134) <= '1';
    layer6_outputs(2135) <= not(layer5_outputs(4276));
    layer6_outputs(2136) <= (layer5_outputs(2720)) or (layer5_outputs(1520));
    layer6_outputs(2137) <= '0';
    layer6_outputs(2138) <= layer5_outputs(2167);
    layer6_outputs(2139) <= not((layer5_outputs(4212)) and (layer5_outputs(4250)));
    layer6_outputs(2140) <= layer5_outputs(106);
    layer6_outputs(2141) <= '0';
    layer6_outputs(2142) <= not((layer5_outputs(495)) xor (layer5_outputs(4987)));
    layer6_outputs(2143) <= layer5_outputs(4339);
    layer6_outputs(2144) <= not((layer5_outputs(1175)) xor (layer5_outputs(417)));
    layer6_outputs(2145) <= (layer5_outputs(3714)) or (layer5_outputs(4478));
    layer6_outputs(2146) <= '1';
    layer6_outputs(2147) <= '1';
    layer6_outputs(2148) <= (layer5_outputs(579)) and not (layer5_outputs(4867));
    layer6_outputs(2149) <= not((layer5_outputs(3270)) xor (layer5_outputs(2421)));
    layer6_outputs(2150) <= not(layer5_outputs(1120)) or (layer5_outputs(2683));
    layer6_outputs(2151) <= layer5_outputs(2576);
    layer6_outputs(2152) <= layer5_outputs(3527);
    layer6_outputs(2153) <= not(layer5_outputs(2255));
    layer6_outputs(2154) <= not(layer5_outputs(427)) or (layer5_outputs(1942));
    layer6_outputs(2155) <= not(layer5_outputs(1725)) or (layer5_outputs(3072));
    layer6_outputs(2156) <= not((layer5_outputs(2698)) xor (layer5_outputs(4633)));
    layer6_outputs(2157) <= not((layer5_outputs(118)) and (layer5_outputs(2771)));
    layer6_outputs(2158) <= not(layer5_outputs(3436)) or (layer5_outputs(4609));
    layer6_outputs(2159) <= not((layer5_outputs(3482)) and (layer5_outputs(4050)));
    layer6_outputs(2160) <= not(layer5_outputs(1949));
    layer6_outputs(2161) <= not((layer5_outputs(2366)) or (layer5_outputs(165)));
    layer6_outputs(2162) <= layer5_outputs(3732);
    layer6_outputs(2163) <= (layer5_outputs(3001)) xor (layer5_outputs(450));
    layer6_outputs(2164) <= not((layer5_outputs(3707)) xor (layer5_outputs(1491)));
    layer6_outputs(2165) <= not(layer5_outputs(2907)) or (layer5_outputs(3450));
    layer6_outputs(2166) <= not(layer5_outputs(4222));
    layer6_outputs(2167) <= layer5_outputs(2482);
    layer6_outputs(2168) <= (layer5_outputs(364)) and (layer5_outputs(2115));
    layer6_outputs(2169) <= not((layer5_outputs(2763)) or (layer5_outputs(22)));
    layer6_outputs(2170) <= layer5_outputs(4859);
    layer6_outputs(2171) <= (layer5_outputs(2300)) and not (layer5_outputs(3020));
    layer6_outputs(2172) <= not(layer5_outputs(4650));
    layer6_outputs(2173) <= not(layer5_outputs(113));
    layer6_outputs(2174) <= (layer5_outputs(484)) and not (layer5_outputs(3477));
    layer6_outputs(2175) <= not(layer5_outputs(4742));
    layer6_outputs(2176) <= not(layer5_outputs(1807));
    layer6_outputs(2177) <= layer5_outputs(3248);
    layer6_outputs(2178) <= not(layer5_outputs(357));
    layer6_outputs(2179) <= not((layer5_outputs(4053)) and (layer5_outputs(2408)));
    layer6_outputs(2180) <= '1';
    layer6_outputs(2181) <= not(layer5_outputs(53));
    layer6_outputs(2182) <= not(layer5_outputs(1096));
    layer6_outputs(2183) <= '1';
    layer6_outputs(2184) <= '1';
    layer6_outputs(2185) <= not(layer5_outputs(1285));
    layer6_outputs(2186) <= not(layer5_outputs(4957));
    layer6_outputs(2187) <= not((layer5_outputs(1344)) and (layer5_outputs(2305)));
    layer6_outputs(2188) <= (layer5_outputs(4762)) xor (layer5_outputs(4767));
    layer6_outputs(2189) <= (layer5_outputs(969)) and not (layer5_outputs(434));
    layer6_outputs(2190) <= '1';
    layer6_outputs(2191) <= not(layer5_outputs(4056));
    layer6_outputs(2192) <= (layer5_outputs(15)) and not (layer5_outputs(1705));
    layer6_outputs(2193) <= layer5_outputs(4680);
    layer6_outputs(2194) <= not(layer5_outputs(208)) or (layer5_outputs(2621));
    layer6_outputs(2195) <= not(layer5_outputs(5095)) or (layer5_outputs(1137));
    layer6_outputs(2196) <= '1';
    layer6_outputs(2197) <= not(layer5_outputs(2721));
    layer6_outputs(2198) <= not(layer5_outputs(3842));
    layer6_outputs(2199) <= not((layer5_outputs(2315)) xor (layer5_outputs(2475)));
    layer6_outputs(2200) <= layer5_outputs(2481);
    layer6_outputs(2201) <= (layer5_outputs(1543)) and not (layer5_outputs(4760));
    layer6_outputs(2202) <= '1';
    layer6_outputs(2203) <= layer5_outputs(2521);
    layer6_outputs(2204) <= not(layer5_outputs(3253));
    layer6_outputs(2205) <= (layer5_outputs(3287)) or (layer5_outputs(2033));
    layer6_outputs(2206) <= layer5_outputs(468);
    layer6_outputs(2207) <= layer5_outputs(1695);
    layer6_outputs(2208) <= (layer5_outputs(267)) and not (layer5_outputs(36));
    layer6_outputs(2209) <= (layer5_outputs(3186)) and not (layer5_outputs(3943));
    layer6_outputs(2210) <= not(layer5_outputs(1355));
    layer6_outputs(2211) <= (layer5_outputs(2412)) or (layer5_outputs(728));
    layer6_outputs(2212) <= not((layer5_outputs(1011)) xor (layer5_outputs(188)));
    layer6_outputs(2213) <= layer5_outputs(2285);
    layer6_outputs(2214) <= (layer5_outputs(2429)) and (layer5_outputs(2848));
    layer6_outputs(2215) <= not(layer5_outputs(551));
    layer6_outputs(2216) <= layer5_outputs(2709);
    layer6_outputs(2217) <= (layer5_outputs(2720)) and not (layer5_outputs(737));
    layer6_outputs(2218) <= (layer5_outputs(3466)) xor (layer5_outputs(2610));
    layer6_outputs(2219) <= not(layer5_outputs(3519)) or (layer5_outputs(3424));
    layer6_outputs(2220) <= not(layer5_outputs(3952)) or (layer5_outputs(1530));
    layer6_outputs(2221) <= (layer5_outputs(4796)) and not (layer5_outputs(3630));
    layer6_outputs(2222) <= (layer5_outputs(1944)) xor (layer5_outputs(2881));
    layer6_outputs(2223) <= layer5_outputs(2532);
    layer6_outputs(2224) <= not(layer5_outputs(476)) or (layer5_outputs(2824));
    layer6_outputs(2225) <= not(layer5_outputs(1170));
    layer6_outputs(2226) <= layer5_outputs(353);
    layer6_outputs(2227) <= not(layer5_outputs(4337));
    layer6_outputs(2228) <= not((layer5_outputs(322)) or (layer5_outputs(4831)));
    layer6_outputs(2229) <= '1';
    layer6_outputs(2230) <= not(layer5_outputs(4672));
    layer6_outputs(2231) <= layer5_outputs(2014);
    layer6_outputs(2232) <= not((layer5_outputs(287)) and (layer5_outputs(3061)));
    layer6_outputs(2233) <= not(layer5_outputs(3440));
    layer6_outputs(2234) <= (layer5_outputs(2755)) and (layer5_outputs(4676));
    layer6_outputs(2235) <= layer5_outputs(184);
    layer6_outputs(2236) <= (layer5_outputs(2095)) xor (layer5_outputs(4656));
    layer6_outputs(2237) <= not((layer5_outputs(2578)) and (layer5_outputs(3021)));
    layer6_outputs(2238) <= not((layer5_outputs(4652)) or (layer5_outputs(951)));
    layer6_outputs(2239) <= layer5_outputs(1717);
    layer6_outputs(2240) <= layer5_outputs(3635);
    layer6_outputs(2241) <= (layer5_outputs(2789)) or (layer5_outputs(4146));
    layer6_outputs(2242) <= (layer5_outputs(3037)) or (layer5_outputs(748));
    layer6_outputs(2243) <= not((layer5_outputs(5008)) or (layer5_outputs(556)));
    layer6_outputs(2244) <= layer5_outputs(277);
    layer6_outputs(2245) <= layer5_outputs(181);
    layer6_outputs(2246) <= not(layer5_outputs(5071)) or (layer5_outputs(3541));
    layer6_outputs(2247) <= (layer5_outputs(3704)) or (layer5_outputs(945));
    layer6_outputs(2248) <= not(layer5_outputs(4221)) or (layer5_outputs(1757));
    layer6_outputs(2249) <= layer5_outputs(4530);
    layer6_outputs(2250) <= '0';
    layer6_outputs(2251) <= layer5_outputs(2329);
    layer6_outputs(2252) <= not(layer5_outputs(4487));
    layer6_outputs(2253) <= not(layer5_outputs(72)) or (layer5_outputs(1344));
    layer6_outputs(2254) <= not(layer5_outputs(275));
    layer6_outputs(2255) <= (layer5_outputs(1406)) xor (layer5_outputs(3855));
    layer6_outputs(2256) <= (layer5_outputs(4470)) and not (layer5_outputs(980));
    layer6_outputs(2257) <= not(layer5_outputs(4139)) or (layer5_outputs(1131));
    layer6_outputs(2258) <= (layer5_outputs(3765)) and not (layer5_outputs(2525));
    layer6_outputs(2259) <= layer5_outputs(3650);
    layer6_outputs(2260) <= not(layer5_outputs(1319));
    layer6_outputs(2261) <= not(layer5_outputs(558));
    layer6_outputs(2262) <= (layer5_outputs(2847)) or (layer5_outputs(952));
    layer6_outputs(2263) <= (layer5_outputs(4504)) and not (layer5_outputs(295));
    layer6_outputs(2264) <= not(layer5_outputs(3403)) or (layer5_outputs(4579));
    layer6_outputs(2265) <= not(layer5_outputs(4449)) or (layer5_outputs(4493));
    layer6_outputs(2266) <= not(layer5_outputs(4605));
    layer6_outputs(2267) <= not(layer5_outputs(1630));
    layer6_outputs(2268) <= not(layer5_outputs(4553));
    layer6_outputs(2269) <= layer5_outputs(3937);
    layer6_outputs(2270) <= (layer5_outputs(151)) xor (layer5_outputs(4941));
    layer6_outputs(2271) <= not(layer5_outputs(2890));
    layer6_outputs(2272) <= not(layer5_outputs(2667));
    layer6_outputs(2273) <= not((layer5_outputs(3283)) and (layer5_outputs(3552)));
    layer6_outputs(2274) <= not((layer5_outputs(4784)) xor (layer5_outputs(32)));
    layer6_outputs(2275) <= not(layer5_outputs(2614));
    layer6_outputs(2276) <= (layer5_outputs(1790)) xor (layer5_outputs(3601));
    layer6_outputs(2277) <= layer5_outputs(4526);
    layer6_outputs(2278) <= '1';
    layer6_outputs(2279) <= (layer5_outputs(1238)) and (layer5_outputs(4717));
    layer6_outputs(2280) <= not(layer5_outputs(1315));
    layer6_outputs(2281) <= (layer5_outputs(4138)) and (layer5_outputs(2699));
    layer6_outputs(2282) <= (layer5_outputs(3781)) and (layer5_outputs(4893));
    layer6_outputs(2283) <= not((layer5_outputs(3335)) or (layer5_outputs(2445)));
    layer6_outputs(2284) <= not(layer5_outputs(318));
    layer6_outputs(2285) <= layer5_outputs(1745);
    layer6_outputs(2286) <= not(layer5_outputs(2648)) or (layer5_outputs(2071));
    layer6_outputs(2287) <= (layer5_outputs(1682)) and not (layer5_outputs(4798));
    layer6_outputs(2288) <= (layer5_outputs(4805)) and not (layer5_outputs(126));
    layer6_outputs(2289) <= not(layer5_outputs(1922));
    layer6_outputs(2290) <= (layer5_outputs(3996)) and (layer5_outputs(3615));
    layer6_outputs(2291) <= (layer5_outputs(3571)) and (layer5_outputs(2035));
    layer6_outputs(2292) <= layer5_outputs(3653);
    layer6_outputs(2293) <= not(layer5_outputs(3847));
    layer6_outputs(2294) <= not((layer5_outputs(1980)) xor (layer5_outputs(2660)));
    layer6_outputs(2295) <= not((layer5_outputs(162)) and (layer5_outputs(4390)));
    layer6_outputs(2296) <= not(layer5_outputs(3086));
    layer6_outputs(2297) <= (layer5_outputs(1862)) and not (layer5_outputs(1385));
    layer6_outputs(2298) <= (layer5_outputs(2706)) and not (layer5_outputs(4530));
    layer6_outputs(2299) <= (layer5_outputs(1067)) and (layer5_outputs(1422));
    layer6_outputs(2300) <= not(layer5_outputs(2669));
    layer6_outputs(2301) <= not((layer5_outputs(2729)) and (layer5_outputs(4137)));
    layer6_outputs(2302) <= not(layer5_outputs(254));
    layer6_outputs(2303) <= not(layer5_outputs(1737));
    layer6_outputs(2304) <= layer5_outputs(1332);
    layer6_outputs(2305) <= not(layer5_outputs(1312)) or (layer5_outputs(3115));
    layer6_outputs(2306) <= not((layer5_outputs(2222)) or (layer5_outputs(5039)));
    layer6_outputs(2307) <= layer5_outputs(5042);
    layer6_outputs(2308) <= layer5_outputs(2440);
    layer6_outputs(2309) <= layer5_outputs(4196);
    layer6_outputs(2310) <= layer5_outputs(2250);
    layer6_outputs(2311) <= not(layer5_outputs(1207)) or (layer5_outputs(1724));
    layer6_outputs(2312) <= (layer5_outputs(3744)) xor (layer5_outputs(3397));
    layer6_outputs(2313) <= layer5_outputs(4371);
    layer6_outputs(2314) <= (layer5_outputs(3714)) or (layer5_outputs(325));
    layer6_outputs(2315) <= (layer5_outputs(1541)) xor (layer5_outputs(3858));
    layer6_outputs(2316) <= not(layer5_outputs(3214)) or (layer5_outputs(2157));
    layer6_outputs(2317) <= (layer5_outputs(2786)) and not (layer5_outputs(1528));
    layer6_outputs(2318) <= not(layer5_outputs(1483));
    layer6_outputs(2319) <= not(layer5_outputs(3562));
    layer6_outputs(2320) <= layer5_outputs(2703);
    layer6_outputs(2321) <= layer5_outputs(683);
    layer6_outputs(2322) <= (layer5_outputs(4845)) and not (layer5_outputs(2026));
    layer6_outputs(2323) <= not(layer5_outputs(2438));
    layer6_outputs(2324) <= '0';
    layer6_outputs(2325) <= not(layer5_outputs(4344)) or (layer5_outputs(3168));
    layer6_outputs(2326) <= (layer5_outputs(2603)) and not (layer5_outputs(1108));
    layer6_outputs(2327) <= not(layer5_outputs(426));
    layer6_outputs(2328) <= layer5_outputs(3835);
    layer6_outputs(2329) <= '0';
    layer6_outputs(2330) <= not((layer5_outputs(1860)) xor (layer5_outputs(2803)));
    layer6_outputs(2331) <= '0';
    layer6_outputs(2332) <= layer5_outputs(188);
    layer6_outputs(2333) <= not((layer5_outputs(3919)) or (layer5_outputs(4022)));
    layer6_outputs(2334) <= (layer5_outputs(3181)) and not (layer5_outputs(19));
    layer6_outputs(2335) <= (layer5_outputs(3469)) and not (layer5_outputs(4086));
    layer6_outputs(2336) <= layer5_outputs(4885);
    layer6_outputs(2337) <= (layer5_outputs(2020)) and not (layer5_outputs(4269));
    layer6_outputs(2338) <= not(layer5_outputs(555));
    layer6_outputs(2339) <= layer5_outputs(4078);
    layer6_outputs(2340) <= layer5_outputs(2684);
    layer6_outputs(2341) <= not(layer5_outputs(2765));
    layer6_outputs(2342) <= (layer5_outputs(1046)) and not (layer5_outputs(331));
    layer6_outputs(2343) <= layer5_outputs(1619);
    layer6_outputs(2344) <= layer5_outputs(676);
    layer6_outputs(2345) <= (layer5_outputs(65)) and not (layer5_outputs(3616));
    layer6_outputs(2346) <= (layer5_outputs(251)) and not (layer5_outputs(865));
    layer6_outputs(2347) <= not(layer5_outputs(4469));
    layer6_outputs(2348) <= not(layer5_outputs(2135)) or (layer5_outputs(3494));
    layer6_outputs(2349) <= (layer5_outputs(357)) or (layer5_outputs(4839));
    layer6_outputs(2350) <= (layer5_outputs(2330)) or (layer5_outputs(310));
    layer6_outputs(2351) <= (layer5_outputs(108)) or (layer5_outputs(1200));
    layer6_outputs(2352) <= not(layer5_outputs(4557));
    layer6_outputs(2353) <= (layer5_outputs(4363)) and not (layer5_outputs(5056));
    layer6_outputs(2354) <= layer5_outputs(3358);
    layer6_outputs(2355) <= (layer5_outputs(198)) or (layer5_outputs(1367));
    layer6_outputs(2356) <= layer5_outputs(1293);
    layer6_outputs(2357) <= not(layer5_outputs(4634)) or (layer5_outputs(3837));
    layer6_outputs(2358) <= (layer5_outputs(968)) and not (layer5_outputs(1377));
    layer6_outputs(2359) <= (layer5_outputs(2893)) and (layer5_outputs(3050));
    layer6_outputs(2360) <= not(layer5_outputs(2612)) or (layer5_outputs(2527));
    layer6_outputs(2361) <= '0';
    layer6_outputs(2362) <= not((layer5_outputs(107)) xor (layer5_outputs(82)));
    layer6_outputs(2363) <= not(layer5_outputs(1055));
    layer6_outputs(2364) <= not((layer5_outputs(3723)) xor (layer5_outputs(3332)));
    layer6_outputs(2365) <= not(layer5_outputs(3445));
    layer6_outputs(2366) <= not(layer5_outputs(909)) or (layer5_outputs(273));
    layer6_outputs(2367) <= '1';
    layer6_outputs(2368) <= not((layer5_outputs(3221)) and (layer5_outputs(4254)));
    layer6_outputs(2369) <= not(layer5_outputs(1946));
    layer6_outputs(2370) <= (layer5_outputs(4796)) and not (layer5_outputs(693));
    layer6_outputs(2371) <= layer5_outputs(1480);
    layer6_outputs(2372) <= (layer5_outputs(2142)) and not (layer5_outputs(2587));
    layer6_outputs(2373) <= not(layer5_outputs(1921)) or (layer5_outputs(3195));
    layer6_outputs(2374) <= (layer5_outputs(4401)) and not (layer5_outputs(4032));
    layer6_outputs(2375) <= (layer5_outputs(1884)) and not (layer5_outputs(4644));
    layer6_outputs(2376) <= not((layer5_outputs(643)) xor (layer5_outputs(2628)));
    layer6_outputs(2377) <= '0';
    layer6_outputs(2378) <= layer5_outputs(1557);
    layer6_outputs(2379) <= layer5_outputs(2434);
    layer6_outputs(2380) <= not((layer5_outputs(282)) and (layer5_outputs(218)));
    layer6_outputs(2381) <= not(layer5_outputs(879)) or (layer5_outputs(1350));
    layer6_outputs(2382) <= '0';
    layer6_outputs(2383) <= layer5_outputs(3228);
    layer6_outputs(2384) <= layer5_outputs(4456);
    layer6_outputs(2385) <= not(layer5_outputs(3703));
    layer6_outputs(2386) <= not(layer5_outputs(3899));
    layer6_outputs(2387) <= not(layer5_outputs(3206)) or (layer5_outputs(921));
    layer6_outputs(2388) <= layer5_outputs(859);
    layer6_outputs(2389) <= not(layer5_outputs(2009)) or (layer5_outputs(4576));
    layer6_outputs(2390) <= '1';
    layer6_outputs(2391) <= (layer5_outputs(5077)) and not (layer5_outputs(3434));
    layer6_outputs(2392) <= '0';
    layer6_outputs(2393) <= (layer5_outputs(4984)) or (layer5_outputs(4564));
    layer6_outputs(2394) <= not(layer5_outputs(4675));
    layer6_outputs(2395) <= not(layer5_outputs(1011));
    layer6_outputs(2396) <= (layer5_outputs(498)) and not (layer5_outputs(2548));
    layer6_outputs(2397) <= layer5_outputs(2224);
    layer6_outputs(2398) <= not(layer5_outputs(4075)) or (layer5_outputs(3896));
    layer6_outputs(2399) <= not(layer5_outputs(3415));
    layer6_outputs(2400) <= not(layer5_outputs(4123));
    layer6_outputs(2401) <= layer5_outputs(4331);
    layer6_outputs(2402) <= not(layer5_outputs(4735));
    layer6_outputs(2403) <= layer5_outputs(3875);
    layer6_outputs(2404) <= layer5_outputs(3036);
    layer6_outputs(2405) <= not(layer5_outputs(1470)) or (layer5_outputs(2362));
    layer6_outputs(2406) <= (layer5_outputs(3793)) or (layer5_outputs(2712));
    layer6_outputs(2407) <= not(layer5_outputs(1558));
    layer6_outputs(2408) <= not(layer5_outputs(2930));
    layer6_outputs(2409) <= not(layer5_outputs(3583));
    layer6_outputs(2410) <= (layer5_outputs(4925)) and (layer5_outputs(3183));
    layer6_outputs(2411) <= (layer5_outputs(3031)) and (layer5_outputs(853));
    layer6_outputs(2412) <= not(layer5_outputs(4434)) or (layer5_outputs(2512));
    layer6_outputs(2413) <= (layer5_outputs(4092)) and not (layer5_outputs(1273));
    layer6_outputs(2414) <= (layer5_outputs(4414)) and (layer5_outputs(2763));
    layer6_outputs(2415) <= (layer5_outputs(1860)) xor (layer5_outputs(1351));
    layer6_outputs(2416) <= not((layer5_outputs(1021)) and (layer5_outputs(2415)));
    layer6_outputs(2417) <= layer5_outputs(406);
    layer6_outputs(2418) <= not(layer5_outputs(386)) or (layer5_outputs(3708));
    layer6_outputs(2419) <= (layer5_outputs(2042)) xor (layer5_outputs(3515));
    layer6_outputs(2420) <= not(layer5_outputs(5093)) or (layer5_outputs(4249));
    layer6_outputs(2421) <= not(layer5_outputs(4820)) or (layer5_outputs(1718));
    layer6_outputs(2422) <= not((layer5_outputs(406)) or (layer5_outputs(2493)));
    layer6_outputs(2423) <= not((layer5_outputs(4915)) and (layer5_outputs(4997)));
    layer6_outputs(2424) <= (layer5_outputs(2608)) xor (layer5_outputs(2023));
    layer6_outputs(2425) <= not((layer5_outputs(973)) and (layer5_outputs(3480)));
    layer6_outputs(2426) <= not((layer5_outputs(2913)) and (layer5_outputs(272)));
    layer6_outputs(2427) <= not(layer5_outputs(996));
    layer6_outputs(2428) <= not(layer5_outputs(2972)) or (layer5_outputs(2566));
    layer6_outputs(2429) <= '0';
    layer6_outputs(2430) <= (layer5_outputs(1251)) xor (layer5_outputs(1942));
    layer6_outputs(2431) <= (layer5_outputs(3057)) or (layer5_outputs(4797));
    layer6_outputs(2432) <= not(layer5_outputs(1956));
    layer6_outputs(2433) <= not((layer5_outputs(3149)) and (layer5_outputs(653)));
    layer6_outputs(2434) <= (layer5_outputs(4100)) or (layer5_outputs(3599));
    layer6_outputs(2435) <= not((layer5_outputs(1471)) or (layer5_outputs(1078)));
    layer6_outputs(2436) <= not((layer5_outputs(4029)) and (layer5_outputs(3751)));
    layer6_outputs(2437) <= not((layer5_outputs(3183)) xor (layer5_outputs(543)));
    layer6_outputs(2438) <= layer5_outputs(2143);
    layer6_outputs(2439) <= not(layer5_outputs(4891));
    layer6_outputs(2440) <= not((layer5_outputs(2185)) and (layer5_outputs(3533)));
    layer6_outputs(2441) <= not(layer5_outputs(861));
    layer6_outputs(2442) <= layer5_outputs(3039);
    layer6_outputs(2443) <= layer5_outputs(297);
    layer6_outputs(2444) <= not(layer5_outputs(3916));
    layer6_outputs(2445) <= layer5_outputs(1316);
    layer6_outputs(2446) <= layer5_outputs(5053);
    layer6_outputs(2447) <= not((layer5_outputs(2117)) xor (layer5_outputs(3389)));
    layer6_outputs(2448) <= (layer5_outputs(3454)) and (layer5_outputs(510));
    layer6_outputs(2449) <= (layer5_outputs(1424)) and (layer5_outputs(172));
    layer6_outputs(2450) <= not(layer5_outputs(1218));
    layer6_outputs(2451) <= '1';
    layer6_outputs(2452) <= (layer5_outputs(4111)) xor (layer5_outputs(701));
    layer6_outputs(2453) <= (layer5_outputs(4869)) or (layer5_outputs(3136));
    layer6_outputs(2454) <= not(layer5_outputs(1728)) or (layer5_outputs(4778));
    layer6_outputs(2455) <= layer5_outputs(1524);
    layer6_outputs(2456) <= (layer5_outputs(411)) xor (layer5_outputs(3177));
    layer6_outputs(2457) <= not((layer5_outputs(1490)) or (layer5_outputs(1345)));
    layer6_outputs(2458) <= not(layer5_outputs(1198));
    layer6_outputs(2459) <= not(layer5_outputs(4081));
    layer6_outputs(2460) <= not(layer5_outputs(2012));
    layer6_outputs(2461) <= not(layer5_outputs(3532)) or (layer5_outputs(1038));
    layer6_outputs(2462) <= not(layer5_outputs(105));
    layer6_outputs(2463) <= not(layer5_outputs(4051));
    layer6_outputs(2464) <= layer5_outputs(3945);
    layer6_outputs(2465) <= layer5_outputs(4457);
    layer6_outputs(2466) <= (layer5_outputs(4036)) and not (layer5_outputs(4134));
    layer6_outputs(2467) <= not(layer5_outputs(2902));
    layer6_outputs(2468) <= layer5_outputs(667);
    layer6_outputs(2469) <= layer5_outputs(4067);
    layer6_outputs(2470) <= (layer5_outputs(2821)) and not (layer5_outputs(4099));
    layer6_outputs(2471) <= '1';
    layer6_outputs(2472) <= layer5_outputs(612);
    layer6_outputs(2473) <= (layer5_outputs(2326)) and not (layer5_outputs(1247));
    layer6_outputs(2474) <= not(layer5_outputs(891)) or (layer5_outputs(2563));
    layer6_outputs(2475) <= (layer5_outputs(1048)) and not (layer5_outputs(2495));
    layer6_outputs(2476) <= (layer5_outputs(4071)) and (layer5_outputs(4785));
    layer6_outputs(2477) <= (layer5_outputs(4197)) and (layer5_outputs(286));
    layer6_outputs(2478) <= '1';
    layer6_outputs(2479) <= (layer5_outputs(1022)) and not (layer5_outputs(267));
    layer6_outputs(2480) <= not(layer5_outputs(4744));
    layer6_outputs(2481) <= not(layer5_outputs(2951));
    layer6_outputs(2482) <= not((layer5_outputs(3327)) or (layer5_outputs(1920)));
    layer6_outputs(2483) <= not(layer5_outputs(3027)) or (layer5_outputs(3052));
    layer6_outputs(2484) <= not((layer5_outputs(3091)) xor (layer5_outputs(1012)));
    layer6_outputs(2485) <= '1';
    layer6_outputs(2486) <= not(layer5_outputs(2105)) or (layer5_outputs(942));
    layer6_outputs(2487) <= (layer5_outputs(4887)) and (layer5_outputs(3298));
    layer6_outputs(2488) <= (layer5_outputs(1098)) or (layer5_outputs(835));
    layer6_outputs(2489) <= not(layer5_outputs(115)) or (layer5_outputs(1804));
    layer6_outputs(2490) <= layer5_outputs(732);
    layer6_outputs(2491) <= layer5_outputs(337);
    layer6_outputs(2492) <= not(layer5_outputs(3145)) or (layer5_outputs(1993));
    layer6_outputs(2493) <= not(layer5_outputs(3390));
    layer6_outputs(2494) <= not(layer5_outputs(955));
    layer6_outputs(2495) <= layer5_outputs(3723);
    layer6_outputs(2496) <= (layer5_outputs(3790)) and (layer5_outputs(4130));
    layer6_outputs(2497) <= (layer5_outputs(2848)) or (layer5_outputs(538));
    layer6_outputs(2498) <= not(layer5_outputs(3830));
    layer6_outputs(2499) <= layer5_outputs(975);
    layer6_outputs(2500) <= '1';
    layer6_outputs(2501) <= not(layer5_outputs(2698)) or (layer5_outputs(1003));
    layer6_outputs(2502) <= layer5_outputs(473);
    layer6_outputs(2503) <= not(layer5_outputs(3869));
    layer6_outputs(2504) <= not(layer5_outputs(4516));
    layer6_outputs(2505) <= not(layer5_outputs(4987)) or (layer5_outputs(1688));
    layer6_outputs(2506) <= not(layer5_outputs(1336));
    layer6_outputs(2507) <= (layer5_outputs(2694)) or (layer5_outputs(1089));
    layer6_outputs(2508) <= (layer5_outputs(2502)) xor (layer5_outputs(820));
    layer6_outputs(2509) <= not(layer5_outputs(3450));
    layer6_outputs(2510) <= not(layer5_outputs(3088));
    layer6_outputs(2511) <= layer5_outputs(595);
    layer6_outputs(2512) <= layer5_outputs(638);
    layer6_outputs(2513) <= layer5_outputs(246);
    layer6_outputs(2514) <= (layer5_outputs(3778)) xor (layer5_outputs(4232));
    layer6_outputs(2515) <= layer5_outputs(3962);
    layer6_outputs(2516) <= not(layer5_outputs(4031));
    layer6_outputs(2517) <= layer5_outputs(946);
    layer6_outputs(2518) <= (layer5_outputs(1881)) and not (layer5_outputs(2795));
    layer6_outputs(2519) <= (layer5_outputs(4310)) and not (layer5_outputs(3627));
    layer6_outputs(2520) <= '0';
    layer6_outputs(2521) <= (layer5_outputs(13)) and not (layer5_outputs(5013));
    layer6_outputs(2522) <= (layer5_outputs(3811)) and not (layer5_outputs(3495));
    layer6_outputs(2523) <= layer5_outputs(29);
    layer6_outputs(2524) <= not(layer5_outputs(3013)) or (layer5_outputs(3077));
    layer6_outputs(2525) <= (layer5_outputs(4864)) xor (layer5_outputs(1830));
    layer6_outputs(2526) <= layer5_outputs(611);
    layer6_outputs(2527) <= layer5_outputs(3139);
    layer6_outputs(2528) <= (layer5_outputs(1206)) xor (layer5_outputs(2443));
    layer6_outputs(2529) <= '1';
    layer6_outputs(2530) <= layer5_outputs(475);
    layer6_outputs(2531) <= (layer5_outputs(1531)) and not (layer5_outputs(1133));
    layer6_outputs(2532) <= not((layer5_outputs(4164)) or (layer5_outputs(1193)));
    layer6_outputs(2533) <= layer5_outputs(3550);
    layer6_outputs(2534) <= not((layer5_outputs(2272)) or (layer5_outputs(2431)));
    layer6_outputs(2535) <= not((layer5_outputs(2664)) and (layer5_outputs(2312)));
    layer6_outputs(2536) <= not(layer5_outputs(874));
    layer6_outputs(2537) <= not((layer5_outputs(4977)) xor (layer5_outputs(4451)));
    layer6_outputs(2538) <= not(layer5_outputs(803));
    layer6_outputs(2539) <= (layer5_outputs(1027)) and not (layer5_outputs(2814));
    layer6_outputs(2540) <= not((layer5_outputs(3741)) or (layer5_outputs(4802)));
    layer6_outputs(2541) <= not(layer5_outputs(4997));
    layer6_outputs(2542) <= (layer5_outputs(1283)) or (layer5_outputs(2111));
    layer6_outputs(2543) <= (layer5_outputs(1584)) and (layer5_outputs(112));
    layer6_outputs(2544) <= layer5_outputs(1113);
    layer6_outputs(2545) <= not(layer5_outputs(3963));
    layer6_outputs(2546) <= '0';
    layer6_outputs(2547) <= not(layer5_outputs(3141));
    layer6_outputs(2548) <= '1';
    layer6_outputs(2549) <= not((layer5_outputs(4915)) and (layer5_outputs(2506)));
    layer6_outputs(2550) <= (layer5_outputs(531)) xor (layer5_outputs(5023));
    layer6_outputs(2551) <= not(layer5_outputs(1)) or (layer5_outputs(5003));
    layer6_outputs(2552) <= '1';
    layer6_outputs(2553) <= layer5_outputs(316);
    layer6_outputs(2554) <= (layer5_outputs(940)) and not (layer5_outputs(2509));
    layer6_outputs(2555) <= (layer5_outputs(3472)) and not (layer5_outputs(4971));
    layer6_outputs(2556) <= not(layer5_outputs(5038)) or (layer5_outputs(2377));
    layer6_outputs(2557) <= not((layer5_outputs(2631)) or (layer5_outputs(3190)));
    layer6_outputs(2558) <= not(layer5_outputs(3349));
    layer6_outputs(2559) <= not(layer5_outputs(1686)) or (layer5_outputs(4879));
    layer6_outputs(2560) <= not(layer5_outputs(79));
    layer6_outputs(2561) <= not((layer5_outputs(3271)) or (layer5_outputs(2026)));
    layer6_outputs(2562) <= (layer5_outputs(2093)) and not (layer5_outputs(2695));
    layer6_outputs(2563) <= not(layer5_outputs(2054)) or (layer5_outputs(544));
    layer6_outputs(2564) <= layer5_outputs(967);
    layer6_outputs(2565) <= not(layer5_outputs(3964));
    layer6_outputs(2566) <= not((layer5_outputs(2871)) xor (layer5_outputs(4973)));
    layer6_outputs(2567) <= (layer5_outputs(1148)) and (layer5_outputs(1926));
    layer6_outputs(2568) <= layer5_outputs(2785);
    layer6_outputs(2569) <= not(layer5_outputs(2846)) or (layer5_outputs(5113));
    layer6_outputs(2570) <= not((layer5_outputs(974)) and (layer5_outputs(1534)));
    layer6_outputs(2571) <= '0';
    layer6_outputs(2572) <= (layer5_outputs(5009)) and not (layer5_outputs(4456));
    layer6_outputs(2573) <= '0';
    layer6_outputs(2574) <= (layer5_outputs(4940)) and not (layer5_outputs(2589));
    layer6_outputs(2575) <= layer5_outputs(2056);
    layer6_outputs(2576) <= not(layer5_outputs(3444));
    layer6_outputs(2577) <= not(layer5_outputs(4882)) or (layer5_outputs(4856));
    layer6_outputs(2578) <= layer5_outputs(2933);
    layer6_outputs(2579) <= (layer5_outputs(3313)) and not (layer5_outputs(4647));
    layer6_outputs(2580) <= layer5_outputs(4858);
    layer6_outputs(2581) <= layer5_outputs(4005);
    layer6_outputs(2582) <= not(layer5_outputs(2204));
    layer6_outputs(2583) <= layer5_outputs(3865);
    layer6_outputs(2584) <= layer5_outputs(4950);
    layer6_outputs(2585) <= not((layer5_outputs(4985)) and (layer5_outputs(1324)));
    layer6_outputs(2586) <= not(layer5_outputs(1258));
    layer6_outputs(2587) <= not(layer5_outputs(2086));
    layer6_outputs(2588) <= layer5_outputs(4254);
    layer6_outputs(2589) <= not(layer5_outputs(5087)) or (layer5_outputs(3153));
    layer6_outputs(2590) <= (layer5_outputs(4000)) and not (layer5_outputs(2376));
    layer6_outputs(2591) <= not(layer5_outputs(4968));
    layer6_outputs(2592) <= not(layer5_outputs(783));
    layer6_outputs(2593) <= not((layer5_outputs(4372)) or (layer5_outputs(3022)));
    layer6_outputs(2594) <= not(layer5_outputs(3791));
    layer6_outputs(2595) <= not(layer5_outputs(207));
    layer6_outputs(2596) <= '1';
    layer6_outputs(2597) <= layer5_outputs(2616);
    layer6_outputs(2598) <= not(layer5_outputs(3037));
    layer6_outputs(2599) <= (layer5_outputs(3570)) or (layer5_outputs(891));
    layer6_outputs(2600) <= (layer5_outputs(4527)) and not (layer5_outputs(1064));
    layer6_outputs(2601) <= layer5_outputs(1093);
    layer6_outputs(2602) <= '1';
    layer6_outputs(2603) <= layer5_outputs(3803);
    layer6_outputs(2604) <= layer5_outputs(561);
    layer6_outputs(2605) <= not((layer5_outputs(133)) or (layer5_outputs(1742)));
    layer6_outputs(2606) <= layer5_outputs(4010);
    layer6_outputs(2607) <= not(layer5_outputs(2355));
    layer6_outputs(2608) <= not(layer5_outputs(244));
    layer6_outputs(2609) <= (layer5_outputs(4416)) and not (layer5_outputs(3859));
    layer6_outputs(2610) <= layer5_outputs(4913);
    layer6_outputs(2611) <= not(layer5_outputs(2859));
    layer6_outputs(2612) <= layer5_outputs(1598);
    layer6_outputs(2613) <= (layer5_outputs(2993)) and not (layer5_outputs(2744));
    layer6_outputs(2614) <= not(layer5_outputs(3531));
    layer6_outputs(2615) <= layer5_outputs(5059);
    layer6_outputs(2616) <= not((layer5_outputs(3082)) or (layer5_outputs(4147)));
    layer6_outputs(2617) <= not(layer5_outputs(1601)) or (layer5_outputs(4810));
    layer6_outputs(2618) <= (layer5_outputs(3075)) xor (layer5_outputs(1081));
    layer6_outputs(2619) <= not(layer5_outputs(3842)) or (layer5_outputs(956));
    layer6_outputs(2620) <= not(layer5_outputs(4983));
    layer6_outputs(2621) <= layer5_outputs(2112);
    layer6_outputs(2622) <= layer5_outputs(2129);
    layer6_outputs(2623) <= layer5_outputs(4030);
    layer6_outputs(2624) <= not((layer5_outputs(1241)) xor (layer5_outputs(854)));
    layer6_outputs(2625) <= layer5_outputs(3817);
    layer6_outputs(2626) <= (layer5_outputs(856)) and not (layer5_outputs(4765));
    layer6_outputs(2627) <= layer5_outputs(160);
    layer6_outputs(2628) <= (layer5_outputs(4589)) and not (layer5_outputs(2613));
    layer6_outputs(2629) <= not((layer5_outputs(1930)) or (layer5_outputs(2714)));
    layer6_outputs(2630) <= (layer5_outputs(742)) and (layer5_outputs(1114));
    layer6_outputs(2631) <= (layer5_outputs(3738)) or (layer5_outputs(1284));
    layer6_outputs(2632) <= not(layer5_outputs(4397)) or (layer5_outputs(3642));
    layer6_outputs(2633) <= not((layer5_outputs(5049)) and (layer5_outputs(1606)));
    layer6_outputs(2634) <= '0';
    layer6_outputs(2635) <= not(layer5_outputs(427)) or (layer5_outputs(2426));
    layer6_outputs(2636) <= '0';
    layer6_outputs(2637) <= '0';
    layer6_outputs(2638) <= not((layer5_outputs(2870)) xor (layer5_outputs(3486)));
    layer6_outputs(2639) <= layer5_outputs(778);
    layer6_outputs(2640) <= (layer5_outputs(1982)) and (layer5_outputs(2679));
    layer6_outputs(2641) <= not(layer5_outputs(30)) or (layer5_outputs(2737));
    layer6_outputs(2642) <= not(layer5_outputs(1326));
    layer6_outputs(2643) <= layer5_outputs(4168);
    layer6_outputs(2644) <= (layer5_outputs(3330)) or (layer5_outputs(4306));
    layer6_outputs(2645) <= '0';
    layer6_outputs(2646) <= layer5_outputs(3632);
    layer6_outputs(2647) <= (layer5_outputs(3619)) and not (layer5_outputs(2853));
    layer6_outputs(2648) <= '1';
    layer6_outputs(2649) <= not(layer5_outputs(2878));
    layer6_outputs(2650) <= not(layer5_outputs(4226)) or (layer5_outputs(2576));
    layer6_outputs(2651) <= (layer5_outputs(824)) or (layer5_outputs(1805));
    layer6_outputs(2652) <= layer5_outputs(2472);
    layer6_outputs(2653) <= layer5_outputs(3755);
    layer6_outputs(2654) <= (layer5_outputs(371)) and not (layer5_outputs(2000));
    layer6_outputs(2655) <= not(layer5_outputs(3575)) or (layer5_outputs(14));
    layer6_outputs(2656) <= layer5_outputs(2472);
    layer6_outputs(2657) <= not((layer5_outputs(775)) and (layer5_outputs(2425)));
    layer6_outputs(2658) <= not((layer5_outputs(5026)) xor (layer5_outputs(3697)));
    layer6_outputs(2659) <= not(layer5_outputs(21)) or (layer5_outputs(1980));
    layer6_outputs(2660) <= not(layer5_outputs(681));
    layer6_outputs(2661) <= '1';
    layer6_outputs(2662) <= (layer5_outputs(5035)) and (layer5_outputs(2379));
    layer6_outputs(2663) <= not((layer5_outputs(1687)) xor (layer5_outputs(3377)));
    layer6_outputs(2664) <= (layer5_outputs(132)) xor (layer5_outputs(1776));
    layer6_outputs(2665) <= not(layer5_outputs(3189));
    layer6_outputs(2666) <= not(layer5_outputs(83)) or (layer5_outputs(4003));
    layer6_outputs(2667) <= (layer5_outputs(4474)) and (layer5_outputs(1447));
    layer6_outputs(2668) <= not(layer5_outputs(2281));
    layer6_outputs(2669) <= (layer5_outputs(2237)) and not (layer5_outputs(604));
    layer6_outputs(2670) <= layer5_outputs(3441);
    layer6_outputs(2671) <= layer5_outputs(4499);
    layer6_outputs(2672) <= (layer5_outputs(2193)) and (layer5_outputs(794));
    layer6_outputs(2673) <= not((layer5_outputs(1309)) or (layer5_outputs(2854)));
    layer6_outputs(2674) <= layer5_outputs(1741);
    layer6_outputs(2675) <= not(layer5_outputs(4287));
    layer6_outputs(2676) <= (layer5_outputs(1030)) and not (layer5_outputs(1852));
    layer6_outputs(2677) <= (layer5_outputs(2420)) and not (layer5_outputs(5008));
    layer6_outputs(2678) <= not((layer5_outputs(2416)) and (layer5_outputs(3274)));
    layer6_outputs(2679) <= (layer5_outputs(2679)) xor (layer5_outputs(4380));
    layer6_outputs(2680) <= layer5_outputs(2538);
    layer6_outputs(2681) <= not((layer5_outputs(374)) and (layer5_outputs(2633)));
    layer6_outputs(2682) <= not(layer5_outputs(1935));
    layer6_outputs(2683) <= layer5_outputs(532);
    layer6_outputs(2684) <= (layer5_outputs(709)) and not (layer5_outputs(622));
    layer6_outputs(2685) <= not(layer5_outputs(4325));
    layer6_outputs(2686) <= not(layer5_outputs(5041));
    layer6_outputs(2687) <= (layer5_outputs(1002)) and not (layer5_outputs(921));
    layer6_outputs(2688) <= (layer5_outputs(4777)) and not (layer5_outputs(2604));
    layer6_outputs(2689) <= (layer5_outputs(4071)) and not (layer5_outputs(749));
    layer6_outputs(2690) <= not((layer5_outputs(1976)) or (layer5_outputs(3864)));
    layer6_outputs(2691) <= '0';
    layer6_outputs(2692) <= (layer5_outputs(4667)) and not (layer5_outputs(722));
    layer6_outputs(2693) <= layer5_outputs(1908);
    layer6_outputs(2694) <= not(layer5_outputs(1261));
    layer6_outputs(2695) <= layer5_outputs(2463);
    layer6_outputs(2696) <= (layer5_outputs(4658)) and not (layer5_outputs(1600));
    layer6_outputs(2697) <= layer5_outputs(2247);
    layer6_outputs(2698) <= not(layer5_outputs(4240));
    layer6_outputs(2699) <= not(layer5_outputs(4986));
    layer6_outputs(2700) <= (layer5_outputs(5091)) and (layer5_outputs(547));
    layer6_outputs(2701) <= '0';
    layer6_outputs(2702) <= (layer5_outputs(4734)) and not (layer5_outputs(35));
    layer6_outputs(2703) <= (layer5_outputs(3159)) xor (layer5_outputs(2617));
    layer6_outputs(2704) <= not(layer5_outputs(1096));
    layer6_outputs(2705) <= not((layer5_outputs(2794)) xor (layer5_outputs(3693)));
    layer6_outputs(2706) <= (layer5_outputs(4511)) and not (layer5_outputs(2490));
    layer6_outputs(2707) <= not((layer5_outputs(3214)) and (layer5_outputs(2687)));
    layer6_outputs(2708) <= (layer5_outputs(1525)) xor (layer5_outputs(897));
    layer6_outputs(2709) <= not(layer5_outputs(4103)) or (layer5_outputs(1155));
    layer6_outputs(2710) <= not(layer5_outputs(2085));
    layer6_outputs(2711) <= (layer5_outputs(2163)) and not (layer5_outputs(142));
    layer6_outputs(2712) <= layer5_outputs(2049);
    layer6_outputs(2713) <= layer5_outputs(3196);
    layer6_outputs(2714) <= not(layer5_outputs(1508));
    layer6_outputs(2715) <= not(layer5_outputs(1372));
    layer6_outputs(2716) <= '1';
    layer6_outputs(2717) <= (layer5_outputs(2865)) and (layer5_outputs(1878));
    layer6_outputs(2718) <= not(layer5_outputs(2584));
    layer6_outputs(2719) <= not(layer5_outputs(1736));
    layer6_outputs(2720) <= not((layer5_outputs(335)) or (layer5_outputs(2427)));
    layer6_outputs(2721) <= not((layer5_outputs(1622)) and (layer5_outputs(1250)));
    layer6_outputs(2722) <= (layer5_outputs(4804)) xor (layer5_outputs(2834));
    layer6_outputs(2723) <= not((layer5_outputs(424)) or (layer5_outputs(2773)));
    layer6_outputs(2724) <= not(layer5_outputs(2005)) or (layer5_outputs(3763));
    layer6_outputs(2725) <= layer5_outputs(3729);
    layer6_outputs(2726) <= not(layer5_outputs(840)) or (layer5_outputs(4951));
    layer6_outputs(2727) <= not((layer5_outputs(1056)) and (layer5_outputs(3226)));
    layer6_outputs(2728) <= '0';
    layer6_outputs(2729) <= not(layer5_outputs(1174));
    layer6_outputs(2730) <= layer5_outputs(760);
    layer6_outputs(2731) <= not(layer5_outputs(4593));
    layer6_outputs(2732) <= not(layer5_outputs(4341)) or (layer5_outputs(381));
    layer6_outputs(2733) <= not(layer5_outputs(28));
    layer6_outputs(2734) <= not(layer5_outputs(2328)) or (layer5_outputs(1972));
    layer6_outputs(2735) <= not(layer5_outputs(4396));
    layer6_outputs(2736) <= (layer5_outputs(3760)) or (layer5_outputs(731));
    layer6_outputs(2737) <= (layer5_outputs(4428)) and not (layer5_outputs(3881));
    layer6_outputs(2738) <= layer5_outputs(2771);
    layer6_outputs(2739) <= not((layer5_outputs(625)) or (layer5_outputs(1130)));
    layer6_outputs(2740) <= not(layer5_outputs(734));
    layer6_outputs(2741) <= (layer5_outputs(4611)) and (layer5_outputs(1765));
    layer6_outputs(2742) <= (layer5_outputs(4114)) xor (layer5_outputs(2515));
    layer6_outputs(2743) <= (layer5_outputs(3354)) or (layer5_outputs(1385));
    layer6_outputs(2744) <= not(layer5_outputs(4824));
    layer6_outputs(2745) <= not(layer5_outputs(3142));
    layer6_outputs(2746) <= not((layer5_outputs(4846)) xor (layer5_outputs(3239)));
    layer6_outputs(2747) <= layer5_outputs(3758);
    layer6_outputs(2748) <= (layer5_outputs(4662)) and not (layer5_outputs(398));
    layer6_outputs(2749) <= not((layer5_outputs(1542)) or (layer5_outputs(4788)));
    layer6_outputs(2750) <= not(layer5_outputs(4361));
    layer6_outputs(2751) <= (layer5_outputs(4476)) and (layer5_outputs(646));
    layer6_outputs(2752) <= '1';
    layer6_outputs(2753) <= not(layer5_outputs(3621));
    layer6_outputs(2754) <= not(layer5_outputs(1444)) or (layer5_outputs(868));
    layer6_outputs(2755) <= (layer5_outputs(1572)) and not (layer5_outputs(3351));
    layer6_outputs(2756) <= (layer5_outputs(418)) and not (layer5_outputs(3685));
    layer6_outputs(2757) <= layer5_outputs(339);
    layer6_outputs(2758) <= not(layer5_outputs(4659));
    layer6_outputs(2759) <= (layer5_outputs(735)) and (layer5_outputs(1538));
    layer6_outputs(2760) <= not((layer5_outputs(741)) or (layer5_outputs(3118)));
    layer6_outputs(2761) <= not(layer5_outputs(929));
    layer6_outputs(2762) <= layer5_outputs(3986);
    layer6_outputs(2763) <= not(layer5_outputs(3043)) or (layer5_outputs(1485));
    layer6_outputs(2764) <= (layer5_outputs(1817)) and not (layer5_outputs(2895));
    layer6_outputs(2765) <= (layer5_outputs(1715)) and not (layer5_outputs(5047));
    layer6_outputs(2766) <= (layer5_outputs(1723)) xor (layer5_outputs(340));
    layer6_outputs(2767) <= not(layer5_outputs(4096)) or (layer5_outputs(84));
    layer6_outputs(2768) <= not((layer5_outputs(4769)) and (layer5_outputs(189)));
    layer6_outputs(2769) <= (layer5_outputs(5089)) or (layer5_outputs(191));
    layer6_outputs(2770) <= layer5_outputs(1914);
    layer6_outputs(2771) <= not(layer5_outputs(4574));
    layer6_outputs(2772) <= not(layer5_outputs(4054));
    layer6_outputs(2773) <= layer5_outputs(3063);
    layer6_outputs(2774) <= not((layer5_outputs(4309)) or (layer5_outputs(684)));
    layer6_outputs(2775) <= not(layer5_outputs(1307));
    layer6_outputs(2776) <= not((layer5_outputs(2752)) and (layer5_outputs(309)));
    layer6_outputs(2777) <= not(layer5_outputs(4449));
    layer6_outputs(2778) <= not((layer5_outputs(2762)) or (layer5_outputs(1143)));
    layer6_outputs(2779) <= not(layer5_outputs(194));
    layer6_outputs(2780) <= not(layer5_outputs(1175)) or (layer5_outputs(4753));
    layer6_outputs(2781) <= not(layer5_outputs(3375));
    layer6_outputs(2782) <= not((layer5_outputs(3322)) and (layer5_outputs(2154)));
    layer6_outputs(2783) <= layer5_outputs(539);
    layer6_outputs(2784) <= (layer5_outputs(1282)) and not (layer5_outputs(2682));
    layer6_outputs(2785) <= not(layer5_outputs(3326));
    layer6_outputs(2786) <= not(layer5_outputs(1944));
    layer6_outputs(2787) <= (layer5_outputs(3143)) and not (layer5_outputs(394));
    layer6_outputs(2788) <= not(layer5_outputs(2479)) or (layer5_outputs(2685));
    layer6_outputs(2789) <= not(layer5_outputs(3576)) or (layer5_outputs(2656));
    layer6_outputs(2790) <= layer5_outputs(3804);
    layer6_outputs(2791) <= not(layer5_outputs(1461));
    layer6_outputs(2792) <= not(layer5_outputs(2189));
    layer6_outputs(2793) <= not((layer5_outputs(3198)) or (layer5_outputs(2165)));
    layer6_outputs(2794) <= (layer5_outputs(3744)) or (layer5_outputs(4419));
    layer6_outputs(2795) <= (layer5_outputs(4766)) or (layer5_outputs(4825));
    layer6_outputs(2796) <= not((layer5_outputs(2353)) and (layer5_outputs(4317)));
    layer6_outputs(2797) <= not(layer5_outputs(4096)) or (layer5_outputs(155));
    layer6_outputs(2798) <= (layer5_outputs(1262)) and not (layer5_outputs(2138));
    layer6_outputs(2799) <= (layer5_outputs(3663)) and (layer5_outputs(2018));
    layer6_outputs(2800) <= layer5_outputs(2449);
    layer6_outputs(2801) <= not((layer5_outputs(2348)) or (layer5_outputs(5096)));
    layer6_outputs(2802) <= not(layer5_outputs(2198));
    layer6_outputs(2803) <= layer5_outputs(1236);
    layer6_outputs(2804) <= not(layer5_outputs(4720));
    layer6_outputs(2805) <= not((layer5_outputs(4671)) xor (layer5_outputs(3395)));
    layer6_outputs(2806) <= not(layer5_outputs(3988)) or (layer5_outputs(4558));
    layer6_outputs(2807) <= layer5_outputs(707);
    layer6_outputs(2808) <= layer5_outputs(2206);
    layer6_outputs(2809) <= (layer5_outputs(463)) xor (layer5_outputs(2772));
    layer6_outputs(2810) <= (layer5_outputs(4535)) and not (layer5_outputs(1925));
    layer6_outputs(2811) <= not(layer5_outputs(1498));
    layer6_outputs(2812) <= layer5_outputs(1159);
    layer6_outputs(2813) <= not((layer5_outputs(3934)) or (layer5_outputs(1188)));
    layer6_outputs(2814) <= (layer5_outputs(2447)) or (layer5_outputs(1919));
    layer6_outputs(2815) <= layer5_outputs(849);
    layer6_outputs(2816) <= (layer5_outputs(4879)) and not (layer5_outputs(3329));
    layer6_outputs(2817) <= not(layer5_outputs(811));
    layer6_outputs(2818) <= not(layer5_outputs(1855));
    layer6_outputs(2819) <= (layer5_outputs(3820)) xor (layer5_outputs(5047));
    layer6_outputs(2820) <= not(layer5_outputs(4415));
    layer6_outputs(2821) <= (layer5_outputs(4927)) and (layer5_outputs(4277));
    layer6_outputs(2822) <= not((layer5_outputs(4581)) and (layer5_outputs(395)));
    layer6_outputs(2823) <= not(layer5_outputs(2501)) or (layer5_outputs(3716));
    layer6_outputs(2824) <= not(layer5_outputs(1205));
    layer6_outputs(2825) <= not(layer5_outputs(4462)) or (layer5_outputs(2072));
    layer6_outputs(2826) <= layer5_outputs(182);
    layer6_outputs(2827) <= (layer5_outputs(307)) or (layer5_outputs(2821));
    layer6_outputs(2828) <= not((layer5_outputs(8)) and (layer5_outputs(1492)));
    layer6_outputs(2829) <= layer5_outputs(1691);
    layer6_outputs(2830) <= (layer5_outputs(270)) and not (layer5_outputs(4775));
    layer6_outputs(2831) <= not((layer5_outputs(1901)) and (layer5_outputs(3968)));
    layer6_outputs(2832) <= not((layer5_outputs(934)) or (layer5_outputs(1189)));
    layer6_outputs(2833) <= not((layer5_outputs(4774)) and (layer5_outputs(1342)));
    layer6_outputs(2834) <= not(layer5_outputs(753));
    layer6_outputs(2835) <= not(layer5_outputs(2693)) or (layer5_outputs(435));
    layer6_outputs(2836) <= not(layer5_outputs(1090));
    layer6_outputs(2837) <= not((layer5_outputs(1222)) xor (layer5_outputs(1718)));
    layer6_outputs(2838) <= not((layer5_outputs(2114)) or (layer5_outputs(1399)));
    layer6_outputs(2839) <= not(layer5_outputs(2258));
    layer6_outputs(2840) <= not(layer5_outputs(4595)) or (layer5_outputs(51));
    layer6_outputs(2841) <= '0';
    layer6_outputs(2842) <= (layer5_outputs(3226)) and not (layer5_outputs(3003));
    layer6_outputs(2843) <= (layer5_outputs(4563)) and (layer5_outputs(460));
    layer6_outputs(2844) <= not(layer5_outputs(2706));
    layer6_outputs(2845) <= not(layer5_outputs(4308));
    layer6_outputs(2846) <= (layer5_outputs(884)) or (layer5_outputs(4230));
    layer6_outputs(2847) <= layer5_outputs(1485);
    layer6_outputs(2848) <= layer5_outputs(1166);
    layer6_outputs(2849) <= not((layer5_outputs(864)) xor (layer5_outputs(1865)));
    layer6_outputs(2850) <= (layer5_outputs(3335)) and not (layer5_outputs(509));
    layer6_outputs(2851) <= not(layer5_outputs(4964)) or (layer5_outputs(2361));
    layer6_outputs(2852) <= not(layer5_outputs(4074));
    layer6_outputs(2853) <= (layer5_outputs(3575)) and not (layer5_outputs(3169));
    layer6_outputs(2854) <= '1';
    layer6_outputs(2855) <= layer5_outputs(3726);
    layer6_outputs(2856) <= layer5_outputs(2108);
    layer6_outputs(2857) <= not(layer5_outputs(4534));
    layer6_outputs(2858) <= not(layer5_outputs(1645));
    layer6_outputs(2859) <= layer5_outputs(1346);
    layer6_outputs(2860) <= layer5_outputs(4345);
    layer6_outputs(2861) <= (layer5_outputs(4852)) and (layer5_outputs(826));
    layer6_outputs(2862) <= (layer5_outputs(2036)) or (layer5_outputs(1962));
    layer6_outputs(2863) <= layer5_outputs(5052);
    layer6_outputs(2864) <= (layer5_outputs(3791)) and (layer5_outputs(2626));
    layer6_outputs(2865) <= not(layer5_outputs(697)) or (layer5_outputs(2993));
    layer6_outputs(2866) <= layer5_outputs(1549);
    layer6_outputs(2867) <= not(layer5_outputs(501)) or (layer5_outputs(4890));
    layer6_outputs(2868) <= layer5_outputs(4340);
    layer6_outputs(2869) <= (layer5_outputs(1181)) and not (layer5_outputs(1647));
    layer6_outputs(2870) <= not((layer5_outputs(590)) and (layer5_outputs(2487)));
    layer6_outputs(2871) <= not(layer5_outputs(1794)) or (layer5_outputs(4021));
    layer6_outputs(2872) <= (layer5_outputs(2311)) or (layer5_outputs(745));
    layer6_outputs(2873) <= (layer5_outputs(525)) and not (layer5_outputs(268));
    layer6_outputs(2874) <= not(layer5_outputs(4282));
    layer6_outputs(2875) <= layer5_outputs(3973);
    layer6_outputs(2876) <= (layer5_outputs(1932)) or (layer5_outputs(2740));
    layer6_outputs(2877) <= not(layer5_outputs(4714));
    layer6_outputs(2878) <= not(layer5_outputs(4562));
    layer6_outputs(2879) <= not(layer5_outputs(434));
    layer6_outputs(2880) <= layer5_outputs(753);
    layer6_outputs(2881) <= not(layer5_outputs(4429)) or (layer5_outputs(4261));
    layer6_outputs(2882) <= (layer5_outputs(3926)) and not (layer5_outputs(1720));
    layer6_outputs(2883) <= not(layer5_outputs(3384));
    layer6_outputs(2884) <= layer5_outputs(1857);
    layer6_outputs(2885) <= '0';
    layer6_outputs(2886) <= not(layer5_outputs(3948));
    layer6_outputs(2887) <= (layer5_outputs(2043)) and not (layer5_outputs(3101));
    layer6_outputs(2888) <= layer5_outputs(1059);
    layer6_outputs(2889) <= layer5_outputs(4335);
    layer6_outputs(2890) <= '1';
    layer6_outputs(2891) <= layer5_outputs(3100);
    layer6_outputs(2892) <= not((layer5_outputs(4712)) and (layer5_outputs(4902)));
    layer6_outputs(2893) <= layer5_outputs(541);
    layer6_outputs(2894) <= (layer5_outputs(1034)) and not (layer5_outputs(686));
    layer6_outputs(2895) <= not(layer5_outputs(970)) or (layer5_outputs(4225));
    layer6_outputs(2896) <= (layer5_outputs(3780)) xor (layer5_outputs(1504));
    layer6_outputs(2897) <= layer5_outputs(4624);
    layer6_outputs(2898) <= layer5_outputs(3356);
    layer6_outputs(2899) <= not(layer5_outputs(4082)) or (layer5_outputs(2615));
    layer6_outputs(2900) <= layer5_outputs(1674);
    layer6_outputs(2901) <= (layer5_outputs(4708)) and not (layer5_outputs(366));
    layer6_outputs(2902) <= not(layer5_outputs(4210));
    layer6_outputs(2903) <= (layer5_outputs(895)) and not (layer5_outputs(1769));
    layer6_outputs(2904) <= not(layer5_outputs(1895));
    layer6_outputs(2905) <= (layer5_outputs(328)) or (layer5_outputs(2318));
    layer6_outputs(2906) <= (layer5_outputs(952)) xor (layer5_outputs(4577));
    layer6_outputs(2907) <= not(layer5_outputs(1729));
    layer6_outputs(2908) <= not((layer5_outputs(926)) or (layer5_outputs(3399)));
    layer6_outputs(2909) <= layer5_outputs(2840);
    layer6_outputs(2910) <= (layer5_outputs(3898)) and not (layer5_outputs(648));
    layer6_outputs(2911) <= not(layer5_outputs(4224));
    layer6_outputs(2912) <= layer5_outputs(3153);
    layer6_outputs(2913) <= layer5_outputs(3416);
    layer6_outputs(2914) <= (layer5_outputs(4035)) and not (layer5_outputs(3948));
    layer6_outputs(2915) <= (layer5_outputs(2287)) or (layer5_outputs(2694));
    layer6_outputs(2916) <= (layer5_outputs(1669)) xor (layer5_outputs(274));
    layer6_outputs(2917) <= layer5_outputs(2314);
    layer6_outputs(2918) <= '0';
    layer6_outputs(2919) <= (layer5_outputs(3311)) or (layer5_outputs(3926));
    layer6_outputs(2920) <= layer5_outputs(2647);
    layer6_outputs(2921) <= not(layer5_outputs(4337)) or (layer5_outputs(3960));
    layer6_outputs(2922) <= not(layer5_outputs(4781)) or (layer5_outputs(2353));
    layer6_outputs(2923) <= not(layer5_outputs(4498));
    layer6_outputs(2924) <= not((layer5_outputs(2678)) and (layer5_outputs(709)));
    layer6_outputs(2925) <= not(layer5_outputs(5055));
    layer6_outputs(2926) <= not(layer5_outputs(3912));
    layer6_outputs(2927) <= layer5_outputs(832);
    layer6_outputs(2928) <= not(layer5_outputs(439));
    layer6_outputs(2929) <= layer5_outputs(3369);
    layer6_outputs(2930) <= (layer5_outputs(2107)) and (layer5_outputs(3924));
    layer6_outputs(2931) <= '0';
    layer6_outputs(2932) <= (layer5_outputs(4351)) and not (layer5_outputs(3584));
    layer6_outputs(2933) <= '1';
    layer6_outputs(2934) <= not(layer5_outputs(4504));
    layer6_outputs(2935) <= not(layer5_outputs(5056)) or (layer5_outputs(4355));
    layer6_outputs(2936) <= layer5_outputs(352);
    layer6_outputs(2937) <= not(layer5_outputs(239)) or (layer5_outputs(549));
    layer6_outputs(2938) <= not(layer5_outputs(2491));
    layer6_outputs(2939) <= (layer5_outputs(2160)) or (layer5_outputs(397));
    layer6_outputs(2940) <= (layer5_outputs(3440)) and not (layer5_outputs(664));
    layer6_outputs(2941) <= layer5_outputs(444);
    layer6_outputs(2942) <= layer5_outputs(2074);
    layer6_outputs(2943) <= '1';
    layer6_outputs(2944) <= not((layer5_outputs(3778)) or (layer5_outputs(3088)));
    layer6_outputs(2945) <= layer5_outputs(1254);
    layer6_outputs(2946) <= layer5_outputs(4488);
    layer6_outputs(2947) <= not(layer5_outputs(3622)) or (layer5_outputs(3536));
    layer6_outputs(2948) <= layer5_outputs(260);
    layer6_outputs(2949) <= not(layer5_outputs(2347));
    layer6_outputs(2950) <= not((layer5_outputs(4978)) and (layer5_outputs(4801)));
    layer6_outputs(2951) <= not(layer5_outputs(1630));
    layer6_outputs(2952) <= not((layer5_outputs(2987)) and (layer5_outputs(3005)));
    layer6_outputs(2953) <= '1';
    layer6_outputs(2954) <= not((layer5_outputs(4884)) or (layer5_outputs(3372)));
    layer6_outputs(2955) <= (layer5_outputs(2845)) and not (layer5_outputs(81));
    layer6_outputs(2956) <= not(layer5_outputs(1880));
    layer6_outputs(2957) <= not(layer5_outputs(1514));
    layer6_outputs(2958) <= not(layer5_outputs(4755));
    layer6_outputs(2959) <= not(layer5_outputs(1659)) or (layer5_outputs(656));
    layer6_outputs(2960) <= (layer5_outputs(614)) and not (layer5_outputs(4699));
    layer6_outputs(2961) <= not(layer5_outputs(4490));
    layer6_outputs(2962) <= not(layer5_outputs(2048));
    layer6_outputs(2963) <= layer5_outputs(2582);
    layer6_outputs(2964) <= (layer5_outputs(3549)) or (layer5_outputs(1933));
    layer6_outputs(2965) <= not(layer5_outputs(3975));
    layer6_outputs(2966) <= '0';
    layer6_outputs(2967) <= not(layer5_outputs(4496)) or (layer5_outputs(1689));
    layer6_outputs(2968) <= (layer5_outputs(1401)) xor (layer5_outputs(3771));
    layer6_outputs(2969) <= (layer5_outputs(2797)) or (layer5_outputs(93));
    layer6_outputs(2970) <= layer5_outputs(3472);
    layer6_outputs(2971) <= (layer5_outputs(4087)) and (layer5_outputs(3548));
    layer6_outputs(2972) <= '0';
    layer6_outputs(2973) <= layer5_outputs(354);
    layer6_outputs(2974) <= not(layer5_outputs(4370));
    layer6_outputs(2975) <= not((layer5_outputs(1357)) xor (layer5_outputs(1803)));
    layer6_outputs(2976) <= (layer5_outputs(1571)) or (layer5_outputs(2711));
    layer6_outputs(2977) <= not(layer5_outputs(1753)) or (layer5_outputs(2794));
    layer6_outputs(2978) <= (layer5_outputs(4843)) and not (layer5_outputs(3743));
    layer6_outputs(2979) <= (layer5_outputs(1103)) and (layer5_outputs(4158));
    layer6_outputs(2980) <= (layer5_outputs(4169)) or (layer5_outputs(4276));
    layer6_outputs(2981) <= layer5_outputs(2131);
    layer6_outputs(2982) <= not(layer5_outputs(5086));
    layer6_outputs(2983) <= (layer5_outputs(3733)) and not (layer5_outputs(19));
    layer6_outputs(2984) <= not(layer5_outputs(4642)) or (layer5_outputs(1703));
    layer6_outputs(2985) <= (layer5_outputs(4969)) and not (layer5_outputs(720));
    layer6_outputs(2986) <= (layer5_outputs(1234)) and (layer5_outputs(1744));
    layer6_outputs(2987) <= not(layer5_outputs(1989));
    layer6_outputs(2988) <= not(layer5_outputs(1192));
    layer6_outputs(2989) <= not(layer5_outputs(3850));
    layer6_outputs(2990) <= not(layer5_outputs(3257)) or (layer5_outputs(4631));
    layer6_outputs(2991) <= not(layer5_outputs(52));
    layer6_outputs(2992) <= layer5_outputs(3970);
    layer6_outputs(2993) <= not(layer5_outputs(4623));
    layer6_outputs(2994) <= (layer5_outputs(2717)) and (layer5_outputs(3790));
    layer6_outputs(2995) <= (layer5_outputs(768)) and not (layer5_outputs(4068));
    layer6_outputs(2996) <= not(layer5_outputs(3608));
    layer6_outputs(2997) <= layer5_outputs(1983);
    layer6_outputs(2998) <= not(layer5_outputs(4135));
    layer6_outputs(2999) <= not(layer5_outputs(4888));
    layer6_outputs(3000) <= (layer5_outputs(334)) and not (layer5_outputs(5072));
    layer6_outputs(3001) <= (layer5_outputs(658)) or (layer5_outputs(480));
    layer6_outputs(3002) <= (layer5_outputs(2212)) and (layer5_outputs(3325));
    layer6_outputs(3003) <= layer5_outputs(455);
    layer6_outputs(3004) <= (layer5_outputs(431)) and not (layer5_outputs(0));
    layer6_outputs(3005) <= not(layer5_outputs(59)) or (layer5_outputs(4362));
    layer6_outputs(3006) <= (layer5_outputs(1738)) and not (layer5_outputs(2700));
    layer6_outputs(3007) <= not((layer5_outputs(1156)) xor (layer5_outputs(2008)));
    layer6_outputs(3008) <= (layer5_outputs(1370)) xor (layer5_outputs(4091));
    layer6_outputs(3009) <= not((layer5_outputs(3273)) or (layer5_outputs(2073)));
    layer6_outputs(3010) <= layer5_outputs(2282);
    layer6_outputs(3011) <= not(layer5_outputs(210)) or (layer5_outputs(2232));
    layer6_outputs(3012) <= not(layer5_outputs(3947));
    layer6_outputs(3013) <= (layer5_outputs(4564)) and (layer5_outputs(2529));
    layer6_outputs(3014) <= (layer5_outputs(3084)) and not (layer5_outputs(4124));
    layer6_outputs(3015) <= (layer5_outputs(4816)) or (layer5_outputs(944));
    layer6_outputs(3016) <= not(layer5_outputs(358));
    layer6_outputs(3017) <= (layer5_outputs(4459)) and (layer5_outputs(2658));
    layer6_outputs(3018) <= not((layer5_outputs(4239)) xor (layer5_outputs(492)));
    layer6_outputs(3019) <= not(layer5_outputs(2335));
    layer6_outputs(3020) <= (layer5_outputs(5044)) and not (layer5_outputs(4996));
    layer6_outputs(3021) <= not(layer5_outputs(2248));
    layer6_outputs(3022) <= not(layer5_outputs(3737));
    layer6_outputs(3023) <= not((layer5_outputs(2921)) and (layer5_outputs(4400)));
    layer6_outputs(3024) <= (layer5_outputs(2590)) and not (layer5_outputs(4791));
    layer6_outputs(3025) <= layer5_outputs(1777);
    layer6_outputs(3026) <= not(layer5_outputs(1208));
    layer6_outputs(3027) <= not((layer5_outputs(55)) or (layer5_outputs(2884)));
    layer6_outputs(3028) <= not((layer5_outputs(2777)) and (layer5_outputs(116)));
    layer6_outputs(3029) <= (layer5_outputs(3586)) xor (layer5_outputs(2944));
    layer6_outputs(3030) <= layer5_outputs(73);
    layer6_outputs(3031) <= not(layer5_outputs(1044));
    layer6_outputs(3032) <= (layer5_outputs(923)) and (layer5_outputs(4391));
    layer6_outputs(3033) <= not(layer5_outputs(4452));
    layer6_outputs(3034) <= '0';
    layer6_outputs(3035) <= layer5_outputs(893);
    layer6_outputs(3036) <= layer5_outputs(4800);
    layer6_outputs(3037) <= (layer5_outputs(200)) and not (layer5_outputs(3161));
    layer6_outputs(3038) <= not((layer5_outputs(3222)) xor (layer5_outputs(3195)));
    layer6_outputs(3039) <= layer5_outputs(3614);
    layer6_outputs(3040) <= not(layer5_outputs(1237)) or (layer5_outputs(368));
    layer6_outputs(3041) <= (layer5_outputs(417)) or (layer5_outputs(482));
    layer6_outputs(3042) <= layer5_outputs(4153);
    layer6_outputs(3043) <= not((layer5_outputs(130)) or (layer5_outputs(513)));
    layer6_outputs(3044) <= not(layer5_outputs(4191));
    layer6_outputs(3045) <= not(layer5_outputs(393));
    layer6_outputs(3046) <= not((layer5_outputs(2211)) and (layer5_outputs(2371)));
    layer6_outputs(3047) <= not(layer5_outputs(312)) or (layer5_outputs(1093));
    layer6_outputs(3048) <= not(layer5_outputs(1335));
    layer6_outputs(3049) <= not(layer5_outputs(542));
    layer6_outputs(3050) <= (layer5_outputs(3808)) and not (layer5_outputs(236));
    layer6_outputs(3051) <= (layer5_outputs(2548)) or (layer5_outputs(858));
    layer6_outputs(3052) <= (layer5_outputs(2460)) and not (layer5_outputs(4861));
    layer6_outputs(3053) <= not(layer5_outputs(1990));
    layer6_outputs(3054) <= (layer5_outputs(1128)) and (layer5_outputs(1866));
    layer6_outputs(3055) <= not(layer5_outputs(3520));
    layer6_outputs(3056) <= layer5_outputs(1613);
    layer6_outputs(3057) <= layer5_outputs(2000);
    layer6_outputs(3058) <= layer5_outputs(3048);
    layer6_outputs(3059) <= not((layer5_outputs(1472)) or (layer5_outputs(1300)));
    layer6_outputs(3060) <= layer5_outputs(630);
    layer6_outputs(3061) <= (layer5_outputs(2060)) and (layer5_outputs(4453));
    layer6_outputs(3062) <= '1';
    layer6_outputs(3063) <= layer5_outputs(3640);
    layer6_outputs(3064) <= '0';
    layer6_outputs(3065) <= layer5_outputs(552);
    layer6_outputs(3066) <= layer5_outputs(3659);
    layer6_outputs(3067) <= (layer5_outputs(2863)) and (layer5_outputs(3676));
    layer6_outputs(3068) <= not(layer5_outputs(1170)) or (layer5_outputs(4728));
    layer6_outputs(3069) <= not(layer5_outputs(4285)) or (layer5_outputs(4763));
    layer6_outputs(3070) <= layer5_outputs(1442);
    layer6_outputs(3071) <= (layer5_outputs(1996)) and (layer5_outputs(5082));
    layer6_outputs(3072) <= '0';
    layer6_outputs(3073) <= not(layer5_outputs(2860));
    layer6_outputs(3074) <= layer5_outputs(1903);
    layer6_outputs(3075) <= (layer5_outputs(2909)) and not (layer5_outputs(1675));
    layer6_outputs(3076) <= layer5_outputs(144);
    layer6_outputs(3077) <= not(layer5_outputs(4743)) or (layer5_outputs(1911));
    layer6_outputs(3078) <= not(layer5_outputs(1384)) or (layer5_outputs(4619));
    layer6_outputs(3079) <= not((layer5_outputs(5016)) and (layer5_outputs(4086)));
    layer6_outputs(3080) <= layer5_outputs(2238);
    layer6_outputs(3081) <= not(layer5_outputs(3369));
    layer6_outputs(3082) <= not((layer5_outputs(2185)) or (layer5_outputs(3072)));
    layer6_outputs(3083) <= layer5_outputs(2221);
    layer6_outputs(3084) <= (layer5_outputs(2552)) and not (layer5_outputs(4605));
    layer6_outputs(3085) <= not((layer5_outputs(2950)) or (layer5_outputs(4591)));
    layer6_outputs(3086) <= not(layer5_outputs(4153));
    layer6_outputs(3087) <= not((layer5_outputs(47)) or (layer5_outputs(3958)));
    layer6_outputs(3088) <= not(layer5_outputs(4617));
    layer6_outputs(3089) <= layer5_outputs(52);
    layer6_outputs(3090) <= not(layer5_outputs(2085));
    layer6_outputs(3091) <= not((layer5_outputs(572)) xor (layer5_outputs(4676)));
    layer6_outputs(3092) <= layer5_outputs(2630);
    layer6_outputs(3093) <= (layer5_outputs(3636)) and not (layer5_outputs(563));
    layer6_outputs(3094) <= not(layer5_outputs(493));
    layer6_outputs(3095) <= not(layer5_outputs(4413)) or (layer5_outputs(1880));
    layer6_outputs(3096) <= not((layer5_outputs(1748)) and (layer5_outputs(4114)));
    layer6_outputs(3097) <= not((layer5_outputs(2439)) and (layer5_outputs(430)));
    layer6_outputs(3098) <= (layer5_outputs(1876)) and not (layer5_outputs(2704));
    layer6_outputs(3099) <= layer5_outputs(1605);
    layer6_outputs(3100) <= (layer5_outputs(3538)) xor (layer5_outputs(850));
    layer6_outputs(3101) <= (layer5_outputs(3965)) and not (layer5_outputs(2062));
    layer6_outputs(3102) <= not((layer5_outputs(4557)) xor (layer5_outputs(1675)));
    layer6_outputs(3103) <= (layer5_outputs(98)) and not (layer5_outputs(2365));
    layer6_outputs(3104) <= not(layer5_outputs(2280));
    layer6_outputs(3105) <= (layer5_outputs(2533)) xor (layer5_outputs(751));
    layer6_outputs(3106) <= not(layer5_outputs(3291));
    layer6_outputs(3107) <= layer5_outputs(4270);
    layer6_outputs(3108) <= (layer5_outputs(4999)) and not (layer5_outputs(1477));
    layer6_outputs(3109) <= not(layer5_outputs(1448)) or (layer5_outputs(2028));
    layer6_outputs(3110) <= not(layer5_outputs(1803)) or (layer5_outputs(980));
    layer6_outputs(3111) <= (layer5_outputs(2832)) or (layer5_outputs(217));
    layer6_outputs(3112) <= not(layer5_outputs(2118)) or (layer5_outputs(4441));
    layer6_outputs(3113) <= '0';
    layer6_outputs(3114) <= not(layer5_outputs(3260)) or (layer5_outputs(767));
    layer6_outputs(3115) <= not(layer5_outputs(3258)) or (layer5_outputs(1777));
    layer6_outputs(3116) <= (layer5_outputs(271)) and not (layer5_outputs(2316));
    layer6_outputs(3117) <= not((layer5_outputs(3391)) and (layer5_outputs(1436)));
    layer6_outputs(3118) <= layer5_outputs(2394);
    layer6_outputs(3119) <= (layer5_outputs(1124)) xor (layer5_outputs(1376));
    layer6_outputs(3120) <= '1';
    layer6_outputs(3121) <= not(layer5_outputs(1408));
    layer6_outputs(3122) <= not(layer5_outputs(4461)) or (layer5_outputs(3636));
    layer6_outputs(3123) <= not((layer5_outputs(3920)) and (layer5_outputs(3569)));
    layer6_outputs(3124) <= layer5_outputs(2396);
    layer6_outputs(3125) <= (layer5_outputs(4097)) and not (layer5_outputs(743));
    layer6_outputs(3126) <= layer5_outputs(868);
    layer6_outputs(3127) <= not(layer5_outputs(3952));
    layer6_outputs(3128) <= (layer5_outputs(2981)) and (layer5_outputs(4014));
    layer6_outputs(3129) <= not((layer5_outputs(3644)) xor (layer5_outputs(4350)));
    layer6_outputs(3130) <= not(layer5_outputs(382));
    layer6_outputs(3131) <= not(layer5_outputs(3980));
    layer6_outputs(3132) <= layer5_outputs(1194);
    layer6_outputs(3133) <= not(layer5_outputs(1801));
    layer6_outputs(3134) <= not(layer5_outputs(4357)) or (layer5_outputs(1038));
    layer6_outputs(3135) <= not(layer5_outputs(3789));
    layer6_outputs(3136) <= (layer5_outputs(1712)) and not (layer5_outputs(2392));
    layer6_outputs(3137) <= not(layer5_outputs(45));
    layer6_outputs(3138) <= not(layer5_outputs(4465)) or (layer5_outputs(2234));
    layer6_outputs(3139) <= layer5_outputs(4781);
    layer6_outputs(3140) <= not(layer5_outputs(4875));
    layer6_outputs(3141) <= layer5_outputs(4575);
    layer6_outputs(3142) <= not(layer5_outputs(3812));
    layer6_outputs(3143) <= not(layer5_outputs(3611));
    layer6_outputs(3144) <= layer5_outputs(4421);
    layer6_outputs(3145) <= not(layer5_outputs(823));
    layer6_outputs(3146) <= '1';
    layer6_outputs(3147) <= not((layer5_outputs(2724)) and (layer5_outputs(286)));
    layer6_outputs(3148) <= layer5_outputs(3900);
    layer6_outputs(3149) <= not((layer5_outputs(4505)) and (layer5_outputs(3040)));
    layer6_outputs(3150) <= not(layer5_outputs(2286)) or (layer5_outputs(1353));
    layer6_outputs(3151) <= (layer5_outputs(356)) xor (layer5_outputs(755));
    layer6_outputs(3152) <= not((layer5_outputs(1353)) xor (layer5_outputs(2981)));
    layer6_outputs(3153) <= (layer5_outputs(2226)) xor (layer5_outputs(4601));
    layer6_outputs(3154) <= not((layer5_outputs(348)) or (layer5_outputs(4184)));
    layer6_outputs(3155) <= (layer5_outputs(3541)) and not (layer5_outputs(754));
    layer6_outputs(3156) <= not(layer5_outputs(3566));
    layer6_outputs(3157) <= not((layer5_outputs(4506)) or (layer5_outputs(1974)));
    layer6_outputs(3158) <= (layer5_outputs(70)) and not (layer5_outputs(3152));
    layer6_outputs(3159) <= not(layer5_outputs(3487)) or (layer5_outputs(2220));
    layer6_outputs(3160) <= not((layer5_outputs(2842)) xor (layer5_outputs(4732)));
    layer6_outputs(3161) <= (layer5_outputs(169)) or (layer5_outputs(2998));
    layer6_outputs(3162) <= layer5_outputs(3980);
    layer6_outputs(3163) <= layer5_outputs(3678);
    layer6_outputs(3164) <= not((layer5_outputs(163)) or (layer5_outputs(3460)));
    layer6_outputs(3165) <= (layer5_outputs(4689)) or (layer5_outputs(948));
    layer6_outputs(3166) <= '1';
    layer6_outputs(3167) <= '1';
    layer6_outputs(3168) <= (layer5_outputs(1580)) or (layer5_outputs(4342));
    layer6_outputs(3169) <= not(layer5_outputs(4596));
    layer6_outputs(3170) <= layer5_outputs(3315);
    layer6_outputs(3171) <= not((layer5_outputs(2337)) xor (layer5_outputs(2994)));
    layer6_outputs(3172) <= layer5_outputs(4544);
    layer6_outputs(3173) <= (layer5_outputs(366)) and not (layer5_outputs(3543));
    layer6_outputs(3174) <= layer5_outputs(2293);
    layer6_outputs(3175) <= (layer5_outputs(1367)) xor (layer5_outputs(4981));
    layer6_outputs(3176) <= not(layer5_outputs(54));
    layer6_outputs(3177) <= not(layer5_outputs(2715)) or (layer5_outputs(2436));
    layer6_outputs(3178) <= not((layer5_outputs(2182)) and (layer5_outputs(1840)));
    layer6_outputs(3179) <= not(layer5_outputs(1789));
    layer6_outputs(3180) <= layer5_outputs(3938);
    layer6_outputs(3181) <= not((layer5_outputs(2709)) or (layer5_outputs(1184)));
    layer6_outputs(3182) <= not((layer5_outputs(3833)) or (layer5_outputs(1246)));
    layer6_outputs(3183) <= not((layer5_outputs(2990)) and (layer5_outputs(4951)));
    layer6_outputs(3184) <= not(layer5_outputs(3051));
    layer6_outputs(3185) <= not(layer5_outputs(2675)) or (layer5_outputs(1532));
    layer6_outputs(3186) <= layer5_outputs(2363);
    layer6_outputs(3187) <= (layer5_outputs(4588)) and not (layer5_outputs(1617));
    layer6_outputs(3188) <= not((layer5_outputs(2701)) or (layer5_outputs(3995)));
    layer6_outputs(3189) <= not(layer5_outputs(4438));
    layer6_outputs(3190) <= '0';
    layer6_outputs(3191) <= not((layer5_outputs(4451)) or (layer5_outputs(1940)));
    layer6_outputs(3192) <= layer5_outputs(4312);
    layer6_outputs(3193) <= not((layer5_outputs(3776)) or (layer5_outputs(4996)));
    layer6_outputs(3194) <= not(layer5_outputs(2456));
    layer6_outputs(3195) <= (layer5_outputs(3362)) and not (layer5_outputs(1196));
    layer6_outputs(3196) <= (layer5_outputs(3605)) and (layer5_outputs(545));
    layer6_outputs(3197) <= layer5_outputs(1183);
    layer6_outputs(3198) <= not(layer5_outputs(661)) or (layer5_outputs(279));
    layer6_outputs(3199) <= not(layer5_outputs(2407));
    layer6_outputs(3200) <= (layer5_outputs(1331)) or (layer5_outputs(3036));
    layer6_outputs(3201) <= not(layer5_outputs(1520)) or (layer5_outputs(4652));
    layer6_outputs(3202) <= layer5_outputs(3111);
    layer6_outputs(3203) <= layer5_outputs(3489);
    layer6_outputs(3204) <= (layer5_outputs(3083)) and not (layer5_outputs(4514));
    layer6_outputs(3205) <= not((layer5_outputs(3371)) and (layer5_outputs(4847)));
    layer6_outputs(3206) <= not((layer5_outputs(4346)) xor (layer5_outputs(3154)));
    layer6_outputs(3207) <= (layer5_outputs(2886)) xor (layer5_outputs(203));
    layer6_outputs(3208) <= layer5_outputs(4837);
    layer6_outputs(3209) <= not(layer5_outputs(5007));
    layer6_outputs(3210) <= not((layer5_outputs(3210)) or (layer5_outputs(1264)));
    layer6_outputs(3211) <= not(layer5_outputs(538)) or (layer5_outputs(4895));
    layer6_outputs(3212) <= not((layer5_outputs(3355)) xor (layer5_outputs(3631)));
    layer6_outputs(3213) <= not((layer5_outputs(1495)) and (layer5_outputs(2715)));
    layer6_outputs(3214) <= '1';
    layer6_outputs(3215) <= layer5_outputs(1119);
    layer6_outputs(3216) <= layer5_outputs(4284);
    layer6_outputs(3217) <= '0';
    layer6_outputs(3218) <= not(layer5_outputs(3667));
    layer6_outputs(3219) <= layer5_outputs(2857);
    layer6_outputs(3220) <= not(layer5_outputs(2601));
    layer6_outputs(3221) <= (layer5_outputs(160)) and (layer5_outputs(1566));
    layer6_outputs(3222) <= not(layer5_outputs(3707)) or (layer5_outputs(2079));
    layer6_outputs(3223) <= not(layer5_outputs(3613)) or (layer5_outputs(4756));
    layer6_outputs(3224) <= not((layer5_outputs(62)) or (layer5_outputs(3432)));
    layer6_outputs(3225) <= layer5_outputs(4617);
    layer6_outputs(3226) <= not(layer5_outputs(1027));
    layer6_outputs(3227) <= not(layer5_outputs(2346));
    layer6_outputs(3228) <= not(layer5_outputs(3829)) or (layer5_outputs(3666));
    layer6_outputs(3229) <= not((layer5_outputs(3851)) and (layer5_outputs(1424)));
    layer6_outputs(3230) <= not(layer5_outputs(2354)) or (layer5_outputs(3479));
    layer6_outputs(3231) <= not((layer5_outputs(2900)) xor (layer5_outputs(2555)));
    layer6_outputs(3232) <= (layer5_outputs(2652)) and not (layer5_outputs(666));
    layer6_outputs(3233) <= (layer5_outputs(4974)) or (layer5_outputs(989));
    layer6_outputs(3234) <= '0';
    layer6_outputs(3235) <= (layer5_outputs(3553)) xor (layer5_outputs(3992));
    layer6_outputs(3236) <= layer5_outputs(1467);
    layer6_outputs(3237) <= (layer5_outputs(296)) and not (layer5_outputs(1669));
    layer6_outputs(3238) <= not(layer5_outputs(1398)) or (layer5_outputs(409));
    layer6_outputs(3239) <= '1';
    layer6_outputs(3240) <= '1';
    layer6_outputs(3241) <= not(layer5_outputs(3903));
    layer6_outputs(3242) <= (layer5_outputs(2361)) and (layer5_outputs(1109));
    layer6_outputs(3243) <= (layer5_outputs(2986)) or (layer5_outputs(3886));
    layer6_outputs(3244) <= not(layer5_outputs(2205)) or (layer5_outputs(1164));
    layer6_outputs(3245) <= not(layer5_outputs(3073)) or (layer5_outputs(4476));
    layer6_outputs(3246) <= not((layer5_outputs(1223)) or (layer5_outputs(930)));
    layer6_outputs(3247) <= layer5_outputs(4664);
    layer6_outputs(3248) <= (layer5_outputs(2814)) or (layer5_outputs(164));
    layer6_outputs(3249) <= (layer5_outputs(3864)) or (layer5_outputs(2389));
    layer6_outputs(3250) <= layer5_outputs(1169);
    layer6_outputs(3251) <= (layer5_outputs(4307)) and (layer5_outputs(4804));
    layer6_outputs(3252) <= not(layer5_outputs(445));
    layer6_outputs(3253) <= not(layer5_outputs(2041)) or (layer5_outputs(1374));
    layer6_outputs(3254) <= not(layer5_outputs(809)) or (layer5_outputs(958));
    layer6_outputs(3255) <= (layer5_outputs(4969)) and not (layer5_outputs(3696));
    layer6_outputs(3256) <= (layer5_outputs(565)) or (layer5_outputs(3761));
    layer6_outputs(3257) <= not(layer5_outputs(663)) or (layer5_outputs(1704));
    layer6_outputs(3258) <= not(layer5_outputs(2735)) or (layer5_outputs(1769));
    layer6_outputs(3259) <= not(layer5_outputs(404));
    layer6_outputs(3260) <= not(layer5_outputs(4318));
    layer6_outputs(3261) <= layer5_outputs(4737);
    layer6_outputs(3262) <= not(layer5_outputs(3302));
    layer6_outputs(3263) <= (layer5_outputs(3623)) and not (layer5_outputs(2443));
    layer6_outputs(3264) <= not((layer5_outputs(851)) or (layer5_outputs(888)));
    layer6_outputs(3265) <= layer5_outputs(3598);
    layer6_outputs(3266) <= not((layer5_outputs(3160)) xor (layer5_outputs(1607)));
    layer6_outputs(3267) <= (layer5_outputs(4423)) or (layer5_outputs(201));
    layer6_outputs(3268) <= not(layer5_outputs(807));
    layer6_outputs(3269) <= '1';
    layer6_outputs(3270) <= not(layer5_outputs(3736));
    layer6_outputs(3271) <= not((layer5_outputs(578)) or (layer5_outputs(1161)));
    layer6_outputs(3272) <= (layer5_outputs(2727)) and not (layer5_outputs(4088));
    layer6_outputs(3273) <= (layer5_outputs(2746)) and not (layer5_outputs(1613));
    layer6_outputs(3274) <= not(layer5_outputs(4298));
    layer6_outputs(3275) <= layer5_outputs(4306);
    layer6_outputs(3276) <= not(layer5_outputs(1161));
    layer6_outputs(3277) <= (layer5_outputs(3972)) or (layer5_outputs(559));
    layer6_outputs(3278) <= layer5_outputs(3014);
    layer6_outputs(3279) <= (layer5_outputs(2224)) and (layer5_outputs(2233));
    layer6_outputs(3280) <= (layer5_outputs(1123)) and not (layer5_outputs(2751));
    layer6_outputs(3281) <= not(layer5_outputs(304));
    layer6_outputs(3282) <= (layer5_outputs(2844)) and (layer5_outputs(3987));
    layer6_outputs(3283) <= layer5_outputs(2089);
    layer6_outputs(3284) <= layer5_outputs(1660);
    layer6_outputs(3285) <= not(layer5_outputs(1437));
    layer6_outputs(3286) <= not(layer5_outputs(175)) or (layer5_outputs(4328));
    layer6_outputs(3287) <= not(layer5_outputs(5109));
    layer6_outputs(3288) <= layer5_outputs(132);
    layer6_outputs(3289) <= layer5_outputs(4477);
    layer6_outputs(3290) <= layer5_outputs(1402);
    layer6_outputs(3291) <= (layer5_outputs(869)) or (layer5_outputs(3));
    layer6_outputs(3292) <= not((layer5_outputs(499)) or (layer5_outputs(1639)));
    layer6_outputs(3293) <= not(layer5_outputs(3211));
    layer6_outputs(3294) <= '0';
    layer6_outputs(3295) <= '0';
    layer6_outputs(3296) <= (layer5_outputs(4519)) and not (layer5_outputs(5077));
    layer6_outputs(3297) <= not(layer5_outputs(2350)) or (layer5_outputs(3670));
    layer6_outputs(3298) <= layer5_outputs(3457);
    layer6_outputs(3299) <= (layer5_outputs(1827)) and not (layer5_outputs(4480));
    layer6_outputs(3300) <= layer5_outputs(3076);
    layer6_outputs(3301) <= '0';
    layer6_outputs(3302) <= not(layer5_outputs(1877));
    layer6_outputs(3303) <= (layer5_outputs(189)) xor (layer5_outputs(1270));
    layer6_outputs(3304) <= (layer5_outputs(3338)) and not (layer5_outputs(3572));
    layer6_outputs(3305) <= (layer5_outputs(966)) and (layer5_outputs(3677));
    layer6_outputs(3306) <= not(layer5_outputs(1271));
    layer6_outputs(3307) <= not((layer5_outputs(324)) or (layer5_outputs(1730)));
    layer6_outputs(3308) <= layer5_outputs(470);
    layer6_outputs(3309) <= (layer5_outputs(3336)) or (layer5_outputs(536));
    layer6_outputs(3310) <= not(layer5_outputs(4576)) or (layer5_outputs(4765));
    layer6_outputs(3311) <= '1';
    layer6_outputs(3312) <= '0';
    layer6_outputs(3313) <= (layer5_outputs(4235)) and not (layer5_outputs(1748));
    layer6_outputs(3314) <= not(layer5_outputs(3931));
    layer6_outputs(3315) <= '0';
    layer6_outputs(3316) <= '1';
    layer6_outputs(3317) <= not(layer5_outputs(3079)) or (layer5_outputs(5034));
    layer6_outputs(3318) <= not(layer5_outputs(4653)) or (layer5_outputs(947));
    layer6_outputs(3319) <= (layer5_outputs(2726)) and not (layer5_outputs(1188));
    layer6_outputs(3320) <= (layer5_outputs(1084)) xor (layer5_outputs(474));
    layer6_outputs(3321) <= not((layer5_outputs(1819)) and (layer5_outputs(2568)));
    layer6_outputs(3322) <= not(layer5_outputs(887)) or (layer5_outputs(3603));
    layer6_outputs(3323) <= not(layer5_outputs(4243));
    layer6_outputs(3324) <= not((layer5_outputs(521)) and (layer5_outputs(3206)));
    layer6_outputs(3325) <= layer5_outputs(4253);
    layer6_outputs(3326) <= layer5_outputs(3518);
    layer6_outputs(3327) <= not(layer5_outputs(583));
    layer6_outputs(3328) <= not(layer5_outputs(1303));
    layer6_outputs(3329) <= not((layer5_outputs(1400)) xor (layer5_outputs(4931)));
    layer6_outputs(3330) <= layer5_outputs(3261);
    layer6_outputs(3331) <= not(layer5_outputs(3735));
    layer6_outputs(3332) <= (layer5_outputs(4863)) xor (layer5_outputs(1820));
    layer6_outputs(3333) <= layer5_outputs(3807);
    layer6_outputs(3334) <= not(layer5_outputs(3689));
    layer6_outputs(3335) <= (layer5_outputs(148)) and not (layer5_outputs(966));
    layer6_outputs(3336) <= not(layer5_outputs(415));
    layer6_outputs(3337) <= not(layer5_outputs(2546)) or (layer5_outputs(1846));
    layer6_outputs(3338) <= not(layer5_outputs(69));
    layer6_outputs(3339) <= '0';
    layer6_outputs(3340) <= (layer5_outputs(2284)) or (layer5_outputs(2308));
    layer6_outputs(3341) <= not(layer5_outputs(2788)) or (layer5_outputs(3196));
    layer6_outputs(3342) <= layer5_outputs(3092);
    layer6_outputs(3343) <= (layer5_outputs(4531)) and not (layer5_outputs(3019));
    layer6_outputs(3344) <= not(layer5_outputs(2719)) or (layer5_outputs(3967));
    layer6_outputs(3345) <= layer5_outputs(4650);
    layer6_outputs(3346) <= layer5_outputs(4345);
    layer6_outputs(3347) <= (layer5_outputs(3788)) and not (layer5_outputs(3418));
    layer6_outputs(3348) <= not(layer5_outputs(2991)) or (layer5_outputs(2749));
    layer6_outputs(3349) <= (layer5_outputs(1523)) xor (layer5_outputs(2652));
    layer6_outputs(3350) <= layer5_outputs(3297);
    layer6_outputs(3351) <= (layer5_outputs(1969)) xor (layer5_outputs(1309));
    layer6_outputs(3352) <= (layer5_outputs(3074)) and (layer5_outputs(4076));
    layer6_outputs(3353) <= not((layer5_outputs(2394)) xor (layer5_outputs(3944)));
    layer6_outputs(3354) <= not(layer5_outputs(885));
    layer6_outputs(3355) <= not(layer5_outputs(1128)) or (layer5_outputs(1014));
    layer6_outputs(3356) <= (layer5_outputs(756)) xor (layer5_outputs(4831));
    layer6_outputs(3357) <= not((layer5_outputs(4740)) and (layer5_outputs(1382)));
    layer6_outputs(3358) <= (layer5_outputs(91)) and (layer5_outputs(4994));
    layer6_outputs(3359) <= (layer5_outputs(2800)) or (layer5_outputs(4933));
    layer6_outputs(3360) <= not(layer5_outputs(2506));
    layer6_outputs(3361) <= not(layer5_outputs(2665));
    layer6_outputs(3362) <= not((layer5_outputs(4201)) or (layer5_outputs(4725)));
    layer6_outputs(3363) <= not(layer5_outputs(2101));
    layer6_outputs(3364) <= layer5_outputs(4892);
    layer6_outputs(3365) <= '0';
    layer6_outputs(3366) <= not((layer5_outputs(1173)) or (layer5_outputs(4698)));
    layer6_outputs(3367) <= not(layer5_outputs(3841)) or (layer5_outputs(2773));
    layer6_outputs(3368) <= (layer5_outputs(3515)) or (layer5_outputs(2104));
    layer6_outputs(3369) <= layer5_outputs(2648);
    layer6_outputs(3370) <= not((layer5_outputs(4089)) xor (layer5_outputs(4945)));
    layer6_outputs(3371) <= (layer5_outputs(4653)) or (layer5_outputs(2834));
    layer6_outputs(3372) <= not(layer5_outputs(4685)) or (layer5_outputs(1954));
    layer6_outputs(3373) <= (layer5_outputs(3172)) xor (layer5_outputs(4730));
    layer6_outputs(3374) <= not(layer5_outputs(4188));
    layer6_outputs(3375) <= '1';
    layer6_outputs(3376) <= not(layer5_outputs(3938)) or (layer5_outputs(3961));
    layer6_outputs(3377) <= layer5_outputs(373);
    layer6_outputs(3378) <= layer5_outputs(3251);
    layer6_outputs(3379) <= not((layer5_outputs(214)) xor (layer5_outputs(959)));
    layer6_outputs(3380) <= not(layer5_outputs(1342));
    layer6_outputs(3381) <= not((layer5_outputs(2572)) or (layer5_outputs(4515)));
    layer6_outputs(3382) <= (layer5_outputs(598)) xor (layer5_outputs(2774));
    layer6_outputs(3383) <= not(layer5_outputs(1025)) or (layer5_outputs(276));
    layer6_outputs(3384) <= layer5_outputs(2885);
    layer6_outputs(3385) <= not(layer5_outputs(2910)) or (layer5_outputs(691));
    layer6_outputs(3386) <= not(layer5_outputs(4426));
    layer6_outputs(3387) <= not(layer5_outputs(438)) or (layer5_outputs(2306));
    layer6_outputs(3388) <= (layer5_outputs(4880)) xor (layer5_outputs(786));
    layer6_outputs(3389) <= (layer5_outputs(208)) and (layer5_outputs(1176));
    layer6_outputs(3390) <= layer5_outputs(787);
    layer6_outputs(3391) <= not(layer5_outputs(1104));
    layer6_outputs(3392) <= not(layer5_outputs(4542));
    layer6_outputs(3393) <= '0';
    layer6_outputs(3394) <= not(layer5_outputs(1414));
    layer6_outputs(3395) <= (layer5_outputs(2137)) and not (layer5_outputs(1065));
    layer6_outputs(3396) <= not((layer5_outputs(4058)) and (layer5_outputs(3797)));
    layer6_outputs(3397) <= '0';
    layer6_outputs(3398) <= (layer5_outputs(4258)) and not (layer5_outputs(1199));
    layer6_outputs(3399) <= (layer5_outputs(1744)) and not (layer5_outputs(2889));
    layer6_outputs(3400) <= (layer5_outputs(5115)) and (layer5_outputs(2454));
    layer6_outputs(3401) <= not((layer5_outputs(902)) and (layer5_outputs(3057)));
    layer6_outputs(3402) <= not((layer5_outputs(4149)) or (layer5_outputs(2522)));
    layer6_outputs(3403) <= not((layer5_outputs(923)) and (layer5_outputs(83)));
    layer6_outputs(3404) <= layer5_outputs(3988);
    layer6_outputs(3405) <= layer5_outputs(5078);
    layer6_outputs(3406) <= (layer5_outputs(2347)) and not (layer5_outputs(2692));
    layer6_outputs(3407) <= not(layer5_outputs(2982));
    layer6_outputs(3408) <= layer5_outputs(1289);
    layer6_outputs(3409) <= not(layer5_outputs(1444));
    layer6_outputs(3410) <= layer5_outputs(4610);
    layer6_outputs(3411) <= layer5_outputs(2906);
    layer6_outputs(3412) <= layer5_outputs(3184);
    layer6_outputs(3413) <= not((layer5_outputs(4289)) or (layer5_outputs(3703)));
    layer6_outputs(3414) <= layer5_outputs(1062);
    layer6_outputs(3415) <= not(layer5_outputs(1466)) or (layer5_outputs(2002));
    layer6_outputs(3416) <= layer5_outputs(4155);
    layer6_outputs(3417) <= not(layer5_outputs(1800));
    layer6_outputs(3418) <= not(layer5_outputs(843)) or (layer5_outputs(1259));
    layer6_outputs(3419) <= layer5_outputs(3977);
    layer6_outputs(3420) <= not(layer5_outputs(1892));
    layer6_outputs(3421) <= not(layer5_outputs(1552));
    layer6_outputs(3422) <= '0';
    layer6_outputs(3423) <= (layer5_outputs(3337)) and not (layer5_outputs(1734));
    layer6_outputs(3424) <= layer5_outputs(863);
    layer6_outputs(3425) <= (layer5_outputs(2256)) or (layer5_outputs(4121));
    layer6_outputs(3426) <= not(layer5_outputs(261));
    layer6_outputs(3427) <= layer5_outputs(1215);
    layer6_outputs(3428) <= (layer5_outputs(138)) and not (layer5_outputs(1532));
    layer6_outputs(3429) <= (layer5_outputs(3777)) and not (layer5_outputs(455));
    layer6_outputs(3430) <= (layer5_outputs(4619)) and (layer5_outputs(235));
    layer6_outputs(3431) <= (layer5_outputs(2332)) and not (layer5_outputs(569));
    layer6_outputs(3432) <= (layer5_outputs(107)) and (layer5_outputs(1328));
    layer6_outputs(3433) <= (layer5_outputs(4691)) and not (layer5_outputs(1280));
    layer6_outputs(3434) <= not(layer5_outputs(3931)) or (layer5_outputs(2097));
    layer6_outputs(3435) <= layer5_outputs(1429);
    layer6_outputs(3436) <= not(layer5_outputs(4679));
    layer6_outputs(3437) <= not((layer5_outputs(899)) and (layer5_outputs(823)));
    layer6_outputs(3438) <= not(layer5_outputs(2489)) or (layer5_outputs(2759));
    layer6_outputs(3439) <= layer5_outputs(3690);
    layer6_outputs(3440) <= layer5_outputs(3100);
    layer6_outputs(3441) <= layer5_outputs(451);
    layer6_outputs(3442) <= layer5_outputs(2184);
    layer6_outputs(3443) <= layer5_outputs(4501);
    layer6_outputs(3444) <= '1';
    layer6_outputs(3445) <= (layer5_outputs(1646)) or (layer5_outputs(847));
    layer6_outputs(3446) <= (layer5_outputs(2452)) or (layer5_outputs(3372));
    layer6_outputs(3447) <= layer5_outputs(448);
    layer6_outputs(3448) <= layer5_outputs(1433);
    layer6_outputs(3449) <= not(layer5_outputs(869));
    layer6_outputs(3450) <= layer5_outputs(2759);
    layer6_outputs(3451) <= layer5_outputs(2635);
    layer6_outputs(3452) <= layer5_outputs(936);
    layer6_outputs(3453) <= not(layer5_outputs(580)) or (layer5_outputs(2605));
    layer6_outputs(3454) <= not(layer5_outputs(4193));
    layer6_outputs(3455) <= not((layer5_outputs(80)) xor (layer5_outputs(2999)));
    layer6_outputs(3456) <= layer5_outputs(1415);
    layer6_outputs(3457) <= (layer5_outputs(3971)) xor (layer5_outputs(2972));
    layer6_outputs(3458) <= (layer5_outputs(2162)) xor (layer5_outputs(1333));
    layer6_outputs(3459) <= not(layer5_outputs(587)) or (layer5_outputs(553));
    layer6_outputs(3460) <= not((layer5_outputs(4559)) or (layer5_outputs(1462)));
    layer6_outputs(3461) <= (layer5_outputs(2045)) and not (layer5_outputs(2707));
    layer6_outputs(3462) <= not(layer5_outputs(4228));
    layer6_outputs(3463) <= not((layer5_outputs(3532)) or (layer5_outputs(2077)));
    layer6_outputs(3464) <= (layer5_outputs(2653)) xor (layer5_outputs(4521));
    layer6_outputs(3465) <= not(layer5_outputs(1547));
    layer6_outputs(3466) <= layer5_outputs(4006);
    layer6_outputs(3467) <= (layer5_outputs(1898)) and (layer5_outputs(4611));
    layer6_outputs(3468) <= not(layer5_outputs(2559));
    layer6_outputs(3469) <= not((layer5_outputs(4686)) or (layer5_outputs(2962)));
    layer6_outputs(3470) <= (layer5_outputs(703)) and (layer5_outputs(2556));
    layer6_outputs(3471) <= not(layer5_outputs(2271));
    layer6_outputs(3472) <= layer5_outputs(500);
    layer6_outputs(3473) <= (layer5_outputs(585)) xor (layer5_outputs(1292));
    layer6_outputs(3474) <= (layer5_outputs(4491)) and not (layer5_outputs(2933));
    layer6_outputs(3475) <= not((layer5_outputs(2477)) xor (layer5_outputs(792)));
    layer6_outputs(3476) <= not(layer5_outputs(1176));
    layer6_outputs(3477) <= not(layer5_outputs(3488)) or (layer5_outputs(4950));
    layer6_outputs(3478) <= not(layer5_outputs(1851));
    layer6_outputs(3479) <= not((layer5_outputs(3241)) and (layer5_outputs(1180)));
    layer6_outputs(3480) <= not(layer5_outputs(2424)) or (layer5_outputs(2316));
    layer6_outputs(3481) <= layer5_outputs(315);
    layer6_outputs(3482) <= not(layer5_outputs(4166)) or (layer5_outputs(1930));
    layer6_outputs(3483) <= not((layer5_outputs(1078)) or (layer5_outputs(2523)));
    layer6_outputs(3484) <= '0';
    layer6_outputs(3485) <= (layer5_outputs(421)) xor (layer5_outputs(4274));
    layer6_outputs(3486) <= layer5_outputs(2547);
    layer6_outputs(3487) <= layer5_outputs(3392);
    layer6_outputs(3488) <= '1';
    layer6_outputs(3489) <= layer5_outputs(4561);
    layer6_outputs(3490) <= layer5_outputs(3974);
    layer6_outputs(3491) <= '1';
    layer6_outputs(3492) <= (layer5_outputs(2604)) xor (layer5_outputs(4641));
    layer6_outputs(3493) <= not(layer5_outputs(4155)) or (layer5_outputs(1733));
    layer6_outputs(3494) <= layer5_outputs(4597);
    layer6_outputs(3495) <= (layer5_outputs(3971)) or (layer5_outputs(3546));
    layer6_outputs(3496) <= (layer5_outputs(3637)) and not (layer5_outputs(423));
    layer6_outputs(3497) <= layer5_outputs(2227);
    layer6_outputs(3498) <= not(layer5_outputs(3998)) or (layer5_outputs(1792));
    layer6_outputs(3499) <= not((layer5_outputs(1466)) and (layer5_outputs(3539)));
    layer6_outputs(3500) <= (layer5_outputs(4364)) or (layer5_outputs(1396));
    layer6_outputs(3501) <= not((layer5_outputs(2673)) and (layer5_outputs(2898)));
    layer6_outputs(3502) <= not(layer5_outputs(5069));
    layer6_outputs(3503) <= (layer5_outputs(2567)) or (layer5_outputs(839));
    layer6_outputs(3504) <= not((layer5_outputs(1223)) or (layer5_outputs(505)));
    layer6_outputs(3505) <= not(layer5_outputs(1852)) or (layer5_outputs(1417));
    layer6_outputs(3506) <= layer5_outputs(426);
    layer6_outputs(3507) <= (layer5_outputs(786)) and (layer5_outputs(2388));
    layer6_outputs(3508) <= not(layer5_outputs(97));
    layer6_outputs(3509) <= not(layer5_outputs(2037)) or (layer5_outputs(1224));
    layer6_outputs(3510) <= (layer5_outputs(197)) and not (layer5_outputs(253));
    layer6_outputs(3511) <= not(layer5_outputs(3257));
    layer6_outputs(3512) <= not(layer5_outputs(778));
    layer6_outputs(3513) <= layer5_outputs(5027);
    layer6_outputs(3514) <= (layer5_outputs(1817)) and (layer5_outputs(4256));
    layer6_outputs(3515) <= not(layer5_outputs(3911));
    layer6_outputs(3516) <= '0';
    layer6_outputs(3517) <= (layer5_outputs(4980)) and not (layer5_outputs(2744));
    layer6_outputs(3518) <= not(layer5_outputs(205));
    layer6_outputs(3519) <= not(layer5_outputs(3772));
    layer6_outputs(3520) <= not(layer5_outputs(899)) or (layer5_outputs(4324));
    layer6_outputs(3521) <= (layer5_outputs(23)) and not (layer5_outputs(1772));
    layer6_outputs(3522) <= not(layer5_outputs(138));
    layer6_outputs(3523) <= (layer5_outputs(4340)) or (layer5_outputs(854));
    layer6_outputs(3524) <= not(layer5_outputs(5107));
    layer6_outputs(3525) <= not(layer5_outputs(2555)) or (layer5_outputs(1979));
    layer6_outputs(3526) <= (layer5_outputs(2559)) and not (layer5_outputs(10));
    layer6_outputs(3527) <= (layer5_outputs(4049)) and not (layer5_outputs(1600));
    layer6_outputs(3528) <= not(layer5_outputs(4512));
    layer6_outputs(3529) <= not((layer5_outputs(3170)) or (layer5_outputs(4400)));
    layer6_outputs(3530) <= not(layer5_outputs(2953));
    layer6_outputs(3531) <= not(layer5_outputs(992));
    layer6_outputs(3532) <= not(layer5_outputs(1099));
    layer6_outputs(3533) <= not(layer5_outputs(4682));
    layer6_outputs(3534) <= not(layer5_outputs(3007));
    layer6_outputs(3535) <= not(layer5_outputs(285));
    layer6_outputs(3536) <= layer5_outputs(2005);
    layer6_outputs(3537) <= not(layer5_outputs(1493));
    layer6_outputs(3538) <= not(layer5_outputs(843));
    layer6_outputs(3539) <= not(layer5_outputs(5111)) or (layer5_outputs(678));
    layer6_outputs(3540) <= not((layer5_outputs(4055)) and (layer5_outputs(2590)));
    layer6_outputs(3541) <= not((layer5_outputs(4958)) and (layer5_outputs(947)));
    layer6_outputs(3542) <= '0';
    layer6_outputs(3543) <= not(layer5_outputs(2208));
    layer6_outputs(3544) <= not(layer5_outputs(4266));
    layer6_outputs(3545) <= layer5_outputs(74);
    layer6_outputs(3546) <= layer5_outputs(3430);
    layer6_outputs(3547) <= not(layer5_outputs(3367));
    layer6_outputs(3548) <= not(layer5_outputs(958));
    layer6_outputs(3549) <= not(layer5_outputs(2618));
    layer6_outputs(3550) <= (layer5_outputs(736)) or (layer5_outputs(456));
    layer6_outputs(3551) <= (layer5_outputs(894)) and not (layer5_outputs(2121));
    layer6_outputs(3552) <= layer5_outputs(2019);
    layer6_outputs(3553) <= not(layer5_outputs(4159));
    layer6_outputs(3554) <= not(layer5_outputs(300)) or (layer5_outputs(729));
    layer6_outputs(3555) <= not(layer5_outputs(3712)) or (layer5_outputs(4832));
    layer6_outputs(3556) <= not(layer5_outputs(2964));
    layer6_outputs(3557) <= not(layer5_outputs(1068));
    layer6_outputs(3558) <= '1';
    layer6_outputs(3559) <= layer5_outputs(4041);
    layer6_outputs(3560) <= not(layer5_outputs(2262)) or (layer5_outputs(593));
    layer6_outputs(3561) <= (layer5_outputs(1462)) and not (layer5_outputs(4639));
    layer6_outputs(3562) <= (layer5_outputs(1508)) and not (layer5_outputs(1662));
    layer6_outputs(3563) <= (layer5_outputs(2491)) or (layer5_outputs(4771));
    layer6_outputs(3564) <= not(layer5_outputs(4221));
    layer6_outputs(3565) <= not(layer5_outputs(1656)) or (layer5_outputs(137));
    layer6_outputs(3566) <= (layer5_outputs(4865)) and not (layer5_outputs(1202));
    layer6_outputs(3567) <= layer5_outputs(4116);
    layer6_outputs(3568) <= not(layer5_outputs(2971)) or (layer5_outputs(3890));
    layer6_outputs(3569) <= not(layer5_outputs(2162));
    layer6_outputs(3570) <= (layer5_outputs(4017)) xor (layer5_outputs(590));
    layer6_outputs(3571) <= layer5_outputs(2345);
    layer6_outputs(3572) <= layer5_outputs(1993);
    layer6_outputs(3573) <= not((layer5_outputs(490)) or (layer5_outputs(4007)));
    layer6_outputs(3574) <= layer5_outputs(582);
    layer6_outputs(3575) <= (layer5_outputs(2007)) xor (layer5_outputs(974));
    layer6_outputs(3576) <= not((layer5_outputs(2071)) or (layer5_outputs(3412)));
    layer6_outputs(3577) <= not(layer5_outputs(4020));
    layer6_outputs(3578) <= layer5_outputs(3346);
    layer6_outputs(3579) <= (layer5_outputs(1828)) and not (layer5_outputs(1183));
    layer6_outputs(3580) <= not((layer5_outputs(637)) or (layer5_outputs(604)));
    layer6_outputs(3581) <= (layer5_outputs(2581)) or (layer5_outputs(243));
    layer6_outputs(3582) <= not(layer5_outputs(3104)) or (layer5_outputs(1839));
    layer6_outputs(3583) <= not((layer5_outputs(180)) or (layer5_outputs(4019)));
    layer6_outputs(3584) <= not(layer5_outputs(2627));
    layer6_outputs(3585) <= layer5_outputs(1515);
    layer6_outputs(3586) <= not(layer5_outputs(2058)) or (layer5_outputs(4791));
    layer6_outputs(3587) <= not(layer5_outputs(1413)) or (layer5_outputs(3973));
    layer6_outputs(3588) <= '0';
    layer6_outputs(3589) <= (layer5_outputs(2849)) and not (layer5_outputs(4142));
    layer6_outputs(3590) <= '0';
    layer6_outputs(3591) <= '0';
    layer6_outputs(3592) <= not(layer5_outputs(4606)) or (layer5_outputs(3212));
    layer6_outputs(3593) <= not((layer5_outputs(5103)) and (layer5_outputs(1760)));
    layer6_outputs(3594) <= (layer5_outputs(3325)) and (layer5_outputs(2880));
    layer6_outputs(3595) <= (layer5_outputs(2955)) or (layer5_outputs(3857));
    layer6_outputs(3596) <= layer5_outputs(298);
    layer6_outputs(3597) <= (layer5_outputs(4173)) and not (layer5_outputs(3089));
    layer6_outputs(3598) <= (layer5_outputs(2911)) and not (layer5_outputs(2728));
    layer6_outputs(3599) <= (layer5_outputs(2330)) and not (layer5_outputs(2040));
    layer6_outputs(3600) <= (layer5_outputs(3230)) and not (layer5_outputs(4229));
    layer6_outputs(3601) <= not((layer5_outputs(2829)) or (layer5_outputs(1133)));
    layer6_outputs(3602) <= not(layer5_outputs(2379)) or (layer5_outputs(1000));
    layer6_outputs(3603) <= not(layer5_outputs(1114));
    layer6_outputs(3604) <= (layer5_outputs(1051)) and not (layer5_outputs(1879));
    layer6_outputs(3605) <= not(layer5_outputs(3858));
    layer6_outputs(3606) <= (layer5_outputs(3749)) and not (layer5_outputs(4532));
    layer6_outputs(3607) <= not((layer5_outputs(4550)) and (layer5_outputs(4773)));
    layer6_outputs(3608) <= not(layer5_outputs(2649)) or (layer5_outputs(1004));
    layer6_outputs(3609) <= not(layer5_outputs(2696));
    layer6_outputs(3610) <= not(layer5_outputs(3178)) or (layer5_outputs(4377));
    layer6_outputs(3611) <= not(layer5_outputs(3420)) or (layer5_outputs(1253));
    layer6_outputs(3612) <= not(layer5_outputs(3853)) or (layer5_outputs(2856));
    layer6_outputs(3613) <= layer5_outputs(452);
    layer6_outputs(3614) <= (layer5_outputs(282)) and not (layer5_outputs(4666));
    layer6_outputs(3615) <= layer5_outputs(3223);
    layer6_outputs(3616) <= (layer5_outputs(2816)) and not (layer5_outputs(920));
    layer6_outputs(3617) <= '0';
    layer6_outputs(3618) <= (layer5_outputs(1318)) and not (layer5_outputs(4008));
    layer6_outputs(3619) <= not(layer5_outputs(3985));
    layer6_outputs(3620) <= not(layer5_outputs(3873));
    layer6_outputs(3621) <= (layer5_outputs(3809)) and (layer5_outputs(1347));
    layer6_outputs(3622) <= (layer5_outputs(4291)) xor (layer5_outputs(3386));
    layer6_outputs(3623) <= '1';
    layer6_outputs(3624) <= layer5_outputs(3130);
    layer6_outputs(3625) <= not(layer5_outputs(4440));
    layer6_outputs(3626) <= not(layer5_outputs(4906));
    layer6_outputs(3627) <= layer5_outputs(621);
    layer6_outputs(3628) <= layer5_outputs(1667);
    layer6_outputs(3629) <= (layer5_outputs(258)) xor (layer5_outputs(1210));
    layer6_outputs(3630) <= layer5_outputs(2992);
    layer6_outputs(3631) <= layer5_outputs(1872);
    layer6_outputs(3632) <= not(layer5_outputs(3783));
    layer6_outputs(3633) <= (layer5_outputs(1943)) or (layer5_outputs(2503));
    layer6_outputs(3634) <= (layer5_outputs(4893)) and not (layer5_outputs(3793));
    layer6_outputs(3635) <= not(layer5_outputs(1169)) or (layer5_outputs(4730));
    layer6_outputs(3636) <= (layer5_outputs(3544)) and not (layer5_outputs(2022));
    layer6_outputs(3637) <= layer5_outputs(1869);
    layer6_outputs(3638) <= layer5_outputs(3400);
    layer6_outputs(3639) <= layer5_outputs(4015);
    layer6_outputs(3640) <= layer5_outputs(3816);
    layer6_outputs(3641) <= layer5_outputs(5009);
    layer6_outputs(3642) <= not(layer5_outputs(3451));
    layer6_outputs(3643) <= not(layer5_outputs(1620)) or (layer5_outputs(2732));
    layer6_outputs(3644) <= (layer5_outputs(4163)) and (layer5_outputs(1885));
    layer6_outputs(3645) <= layer5_outputs(1291);
    layer6_outputs(3646) <= layer5_outputs(3749);
    layer6_outputs(3647) <= '0';
    layer6_outputs(3648) <= not(layer5_outputs(81)) or (layer5_outputs(2134));
    layer6_outputs(3649) <= layer5_outputs(827);
    layer6_outputs(3650) <= (layer5_outputs(254)) and not (layer5_outputs(1102));
    layer6_outputs(3651) <= (layer5_outputs(1515)) and not (layer5_outputs(3059));
    layer6_outputs(3652) <= not(layer5_outputs(4)) or (layer5_outputs(4244));
    layer6_outputs(3653) <= (layer5_outputs(2140)) xor (layer5_outputs(552));
    layer6_outputs(3654) <= not((layer5_outputs(739)) xor (layer5_outputs(3017)));
    layer6_outputs(3655) <= not(layer5_outputs(2004)) or (layer5_outputs(3649));
    layer6_outputs(3656) <= layer5_outputs(2075);
    layer6_outputs(3657) <= layer5_outputs(4785);
    layer6_outputs(3658) <= layer5_outputs(4070);
    layer6_outputs(3659) <= not(layer5_outputs(1268));
    layer6_outputs(3660) <= not((layer5_outputs(4415)) xor (layer5_outputs(95)));
    layer6_outputs(3661) <= not((layer5_outputs(3341)) or (layer5_outputs(984)));
    layer6_outputs(3662) <= not(layer5_outputs(1028)) or (layer5_outputs(305));
    layer6_outputs(3663) <= (layer5_outputs(4182)) and not (layer5_outputs(1341));
    layer6_outputs(3664) <= (layer5_outputs(1502)) and (layer5_outputs(1455));
    layer6_outputs(3665) <= not((layer5_outputs(771)) or (layer5_outputs(2503)));
    layer6_outputs(3666) <= not(layer5_outputs(878));
    layer6_outputs(3667) <= not((layer5_outputs(4215)) xor (layer5_outputs(1391)));
    layer6_outputs(3668) <= layer5_outputs(1885);
    layer6_outputs(3669) <= not(layer5_outputs(4868)) or (layer5_outputs(779));
    layer6_outputs(3670) <= not(layer5_outputs(1992));
    layer6_outputs(3671) <= not(layer5_outputs(2246));
    layer6_outputs(3672) <= not((layer5_outputs(3645)) and (layer5_outputs(1988)));
    layer6_outputs(3673) <= layer5_outputs(3407);
    layer6_outputs(3674) <= (layer5_outputs(3831)) and not (layer5_outputs(1134));
    layer6_outputs(3675) <= not(layer5_outputs(3517)) or (layer5_outputs(3932));
    layer6_outputs(3676) <= not(layer5_outputs(2681));
    layer6_outputs(3677) <= not(layer5_outputs(2522));
    layer6_outputs(3678) <= not(layer5_outputs(4320));
    layer6_outputs(3679) <= not(layer5_outputs(950));
    layer6_outputs(3680) <= (layer5_outputs(4953)) and (layer5_outputs(547));
    layer6_outputs(3681) <= (layer5_outputs(3529)) and (layer5_outputs(2025));
    layer6_outputs(3682) <= layer5_outputs(2143);
    layer6_outputs(3683) <= (layer5_outputs(2323)) xor (layer5_outputs(642));
    layer6_outputs(3684) <= not(layer5_outputs(2172));
    layer6_outputs(3685) <= (layer5_outputs(4818)) or (layer5_outputs(2769));
    layer6_outputs(3686) <= (layer5_outputs(2995)) or (layer5_outputs(2010));
    layer6_outputs(3687) <= not(layer5_outputs(2906));
    layer6_outputs(3688) <= not(layer5_outputs(2818)) or (layer5_outputs(3613));
    layer6_outputs(3689) <= (layer5_outputs(4590)) and (layer5_outputs(2961));
    layer6_outputs(3690) <= not(layer5_outputs(3223)) or (layer5_outputs(1549));
    layer6_outputs(3691) <= (layer5_outputs(3969)) xor (layer5_outputs(4034));
    layer6_outputs(3692) <= layer5_outputs(822);
    layer6_outputs(3693) <= layer5_outputs(3804);
    layer6_outputs(3694) <= layer5_outputs(4889);
    layer6_outputs(3695) <= not((layer5_outputs(1864)) and (layer5_outputs(2296)));
    layer6_outputs(3696) <= '0';
    layer6_outputs(3697) <= (layer5_outputs(845)) and (layer5_outputs(1459));
    layer6_outputs(3698) <= not(layer5_outputs(1266));
    layer6_outputs(3699) <= not(layer5_outputs(3737));
    layer6_outputs(3700) <= layer5_outputs(2526);
    layer6_outputs(3701) <= not((layer5_outputs(380)) xor (layer5_outputs(24)));
    layer6_outputs(3702) <= '0';
    layer6_outputs(3703) <= (layer5_outputs(2057)) and not (layer5_outputs(3471));
    layer6_outputs(3704) <= layer5_outputs(1455);
    layer6_outputs(3705) <= not(layer5_outputs(2225));
    layer6_outputs(3706) <= not(layer5_outputs(1827));
    layer6_outputs(3707) <= (layer5_outputs(3254)) and (layer5_outputs(290));
    layer6_outputs(3708) <= '0';
    layer6_outputs(3709) <= not(layer5_outputs(3368)) or (layer5_outputs(3299));
    layer6_outputs(3710) <= (layer5_outputs(1642)) and (layer5_outputs(2093));
    layer6_outputs(3711) <= not(layer5_outputs(1576));
    layer6_outputs(3712) <= layer5_outputs(2144);
    layer6_outputs(3713) <= (layer5_outputs(5065)) or (layer5_outputs(1245));
    layer6_outputs(3714) <= (layer5_outputs(846)) and (layer5_outputs(3220));
    layer6_outputs(3715) <= not(layer5_outputs(3305));
    layer6_outputs(3716) <= not(layer5_outputs(1360));
    layer6_outputs(3717) <= not(layer5_outputs(925));
    layer6_outputs(3718) <= (layer5_outputs(4303)) and not (layer5_outputs(1007));
    layer6_outputs(3719) <= (layer5_outputs(4039)) xor (layer5_outputs(1259));
    layer6_outputs(3720) <= (layer5_outputs(1929)) and not (layer5_outputs(1689));
    layer6_outputs(3721) <= not(layer5_outputs(2807));
    layer6_outputs(3722) <= layer5_outputs(4523);
    layer6_outputs(3723) <= not((layer5_outputs(1213)) xor (layer5_outputs(3302)));
    layer6_outputs(3724) <= not(layer5_outputs(2462));
    layer6_outputs(3725) <= '0';
    layer6_outputs(3726) <= '0';
    layer6_outputs(3727) <= layer5_outputs(3840);
    layer6_outputs(3728) <= (layer5_outputs(4369)) and not (layer5_outputs(5070));
    layer6_outputs(3729) <= '1';
    layer6_outputs(3730) <= not((layer5_outputs(867)) or (layer5_outputs(215)));
    layer6_outputs(3731) <= not(layer5_outputs(4640));
    layer6_outputs(3732) <= '1';
    layer6_outputs(3733) <= not(layer5_outputs(924));
    layer6_outputs(3734) <= (layer5_outputs(4714)) and not (layer5_outputs(3531));
    layer6_outputs(3735) <= (layer5_outputs(781)) and (layer5_outputs(328));
    layer6_outputs(3736) <= (layer5_outputs(2265)) or (layer5_outputs(3361));
    layer6_outputs(3737) <= (layer5_outputs(3341)) and not (layer5_outputs(2270));
    layer6_outputs(3738) <= (layer5_outputs(197)) and (layer5_outputs(1768));
    layer6_outputs(3739) <= (layer5_outputs(1976)) xor (layer5_outputs(4886));
    layer6_outputs(3740) <= not(layer5_outputs(2091));
    layer6_outputs(3741) <= not(layer5_outputs(4112));
    layer6_outputs(3742) <= not((layer5_outputs(3504)) or (layer5_outputs(4960)));
    layer6_outputs(3743) <= layer5_outputs(4573);
    layer6_outputs(3744) <= not(layer5_outputs(3292));
    layer6_outputs(3745) <= not(layer5_outputs(4794)) or (layer5_outputs(1463));
    layer6_outputs(3746) <= (layer5_outputs(5013)) xor (layer5_outputs(193));
    layer6_outputs(3747) <= not(layer5_outputs(1409));
    layer6_outputs(3748) <= not((layer5_outputs(3480)) and (layer5_outputs(1781)));
    layer6_outputs(3749) <= (layer5_outputs(4283)) xor (layer5_outputs(3865));
    layer6_outputs(3750) <= not(layer5_outputs(1306)) or (layer5_outputs(4347));
    layer6_outputs(3751) <= not(layer5_outputs(2438));
    layer6_outputs(3752) <= not((layer5_outputs(634)) xor (layer5_outputs(2602)));
    layer6_outputs(3753) <= not(layer5_outputs(570));
    layer6_outputs(3754) <= not((layer5_outputs(4547)) or (layer5_outputs(4328)));
    layer6_outputs(3755) <= not(layer5_outputs(1055));
    layer6_outputs(3756) <= not(layer5_outputs(1193));
    layer6_outputs(3757) <= not((layer5_outputs(4776)) or (layer5_outputs(217)));
    layer6_outputs(3758) <= (layer5_outputs(2136)) and (layer5_outputs(4694));
    layer6_outputs(3759) <= (layer5_outputs(146)) and (layer5_outputs(2349));
    layer6_outputs(3760) <= (layer5_outputs(1855)) xor (layer5_outputs(3133));
    layer6_outputs(3761) <= not(layer5_outputs(3549));
    layer6_outputs(3762) <= not((layer5_outputs(4464)) or (layer5_outputs(4640)));
    layer6_outputs(3763) <= not((layer5_outputs(560)) and (layer5_outputs(2921)));
    layer6_outputs(3764) <= layer5_outputs(3510);
    layer6_outputs(3765) <= layer5_outputs(4983);
    layer6_outputs(3766) <= not(layer5_outputs(3156));
    layer6_outputs(3767) <= (layer5_outputs(3688)) and not (layer5_outputs(2801));
    layer6_outputs(3768) <= not((layer5_outputs(3698)) or (layer5_outputs(2919)));
    layer6_outputs(3769) <= not(layer5_outputs(4855));
    layer6_outputs(3770) <= not(layer5_outputs(3700));
    layer6_outputs(3771) <= (layer5_outputs(662)) and (layer5_outputs(3949));
    layer6_outputs(3772) <= not(layer5_outputs(1509));
    layer6_outputs(3773) <= not(layer5_outputs(3008)) or (layer5_outputs(402));
    layer6_outputs(3774) <= layer5_outputs(2155);
    layer6_outputs(3775) <= not(layer5_outputs(327));
    layer6_outputs(3776) <= not(layer5_outputs(3314));
    layer6_outputs(3777) <= layer5_outputs(2520);
    layer6_outputs(3778) <= (layer5_outputs(2124)) and (layer5_outputs(487));
    layer6_outputs(3779) <= (layer5_outputs(2677)) or (layer5_outputs(3617));
    layer6_outputs(3780) <= '0';
    layer6_outputs(3781) <= not(layer5_outputs(1274));
    layer6_outputs(3782) <= (layer5_outputs(824)) or (layer5_outputs(2285));
    layer6_outputs(3783) <= not((layer5_outputs(2739)) xor (layer5_outputs(603)));
    layer6_outputs(3784) <= not(layer5_outputs(1166));
    layer6_outputs(3785) <= (layer5_outputs(1369)) and (layer5_outputs(1778));
    layer6_outputs(3786) <= (layer5_outputs(2731)) xor (layer5_outputs(1314));
    layer6_outputs(3787) <= (layer5_outputs(1130)) and not (layer5_outputs(1366));
    layer6_outputs(3788) <= (layer5_outputs(3023)) and (layer5_outputs(2623));
    layer6_outputs(3789) <= not((layer5_outputs(1688)) xor (layer5_outputs(1870)));
    layer6_outputs(3790) <= not(layer5_outputs(3024));
    layer6_outputs(3791) <= (layer5_outputs(3081)) and not (layer5_outputs(1240));
    layer6_outputs(3792) <= layer5_outputs(4665);
    layer6_outputs(3793) <= (layer5_outputs(3803)) and not (layer5_outputs(42));
    layer6_outputs(3794) <= not(layer5_outputs(4937));
    layer6_outputs(3795) <= not(layer5_outputs(714)) or (layer5_outputs(4404));
    layer6_outputs(3796) <= not(layer5_outputs(2258)) or (layer5_outputs(416));
    layer6_outputs(3797) <= (layer5_outputs(2809)) and not (layer5_outputs(1158));
    layer6_outputs(3798) <= not(layer5_outputs(3374));
    layer6_outputs(3799) <= not(layer5_outputs(2061));
    layer6_outputs(3800) <= (layer5_outputs(3373)) or (layer5_outputs(5057));
    layer6_outputs(3801) <= layer5_outputs(341);
    layer6_outputs(3802) <= not(layer5_outputs(1965)) or (layer5_outputs(1334));
    layer6_outputs(3803) <= not((layer5_outputs(5106)) and (layer5_outputs(4180)));
    layer6_outputs(3804) <= layer5_outputs(2041);
    layer6_outputs(3805) <= not((layer5_outputs(4061)) xor (layer5_outputs(4643)));
    layer6_outputs(3806) <= layer5_outputs(3637);
    layer6_outputs(3807) <= (layer5_outputs(3700)) or (layer5_outputs(1749));
    layer6_outputs(3808) <= not(layer5_outputs(4412));
    layer6_outputs(3809) <= not(layer5_outputs(1531));
    layer6_outputs(3810) <= layer5_outputs(2262);
    layer6_outputs(3811) <= not(layer5_outputs(1390)) or (layer5_outputs(3650));
    layer6_outputs(3812) <= not(layer5_outputs(129)) or (layer5_outputs(3255));
    layer6_outputs(3813) <= layer5_outputs(4696);
    layer6_outputs(3814) <= not(layer5_outputs(4920));
    layer6_outputs(3815) <= not(layer5_outputs(4627));
    layer6_outputs(3816) <= not((layer5_outputs(3819)) or (layer5_outputs(4251)));
    layer6_outputs(3817) <= not(layer5_outputs(1957)) or (layer5_outputs(2721));
    layer6_outputs(3818) <= not(layer5_outputs(1591)) or (layer5_outputs(747));
    layer6_outputs(3819) <= (layer5_outputs(4982)) and (layer5_outputs(4305));
    layer6_outputs(3820) <= layer5_outputs(3469);
    layer6_outputs(3821) <= not(layer5_outputs(769));
    layer6_outputs(3822) <= '1';
    layer6_outputs(3823) <= layer5_outputs(4058);
    layer6_outputs(3824) <= not((layer5_outputs(4116)) or (layer5_outputs(1410)));
    layer6_outputs(3825) <= not((layer5_outputs(2436)) or (layer5_outputs(3782)));
    layer6_outputs(3826) <= not((layer5_outputs(4219)) or (layer5_outputs(2370)));
    layer6_outputs(3827) <= not(layer5_outputs(2762));
    layer6_outputs(3828) <= (layer5_outputs(4830)) and not (layer5_outputs(1372));
    layer6_outputs(3829) <= (layer5_outputs(4094)) and not (layer5_outputs(2554));
    layer6_outputs(3830) <= not((layer5_outputs(1609)) or (layer5_outputs(1667)));
    layer6_outputs(3831) <= not((layer5_outputs(581)) and (layer5_outputs(503)));
    layer6_outputs(3832) <= not(layer5_outputs(3806)) or (layer5_outputs(1848));
    layer6_outputs(3833) <= layer5_outputs(3485);
    layer6_outputs(3834) <= not(layer5_outputs(82));
    layer6_outputs(3835) <= layer5_outputs(1400);
    layer6_outputs(3836) <= layer5_outputs(4702);
    layer6_outputs(3837) <= not(layer5_outputs(3030));
    layer6_outputs(3838) <= (layer5_outputs(2750)) xor (layer5_outputs(436));
    layer6_outputs(3839) <= not(layer5_outputs(24));
    layer6_outputs(3840) <= '0';
    layer6_outputs(3841) <= (layer5_outputs(1189)) and (layer5_outputs(1559));
    layer6_outputs(3842) <= not(layer5_outputs(204));
    layer6_outputs(3843) <= (layer5_outputs(3265)) and not (layer5_outputs(2070));
    layer6_outputs(3844) <= (layer5_outputs(1415)) xor (layer5_outputs(3498));
    layer6_outputs(3845) <= not(layer5_outputs(44)) or (layer5_outputs(2158));
    layer6_outputs(3846) <= (layer5_outputs(5112)) and not (layer5_outputs(1574));
    layer6_outputs(3847) <= not((layer5_outputs(4722)) or (layer5_outputs(1432)));
    layer6_outputs(3848) <= (layer5_outputs(1321)) and not (layer5_outputs(4104));
    layer6_outputs(3849) <= not(layer5_outputs(2368));
    layer6_outputs(3850) <= (layer5_outputs(4717)) and (layer5_outputs(2106));
    layer6_outputs(3851) <= layer5_outputs(1806);
    layer6_outputs(3852) <= not((layer5_outputs(3917)) and (layer5_outputs(1374)));
    layer6_outputs(3853) <= not((layer5_outputs(3155)) xor (layer5_outputs(305)));
    layer6_outputs(3854) <= not((layer5_outputs(3194)) and (layer5_outputs(2858)));
    layer6_outputs(3855) <= not((layer5_outputs(4304)) and (layer5_outputs(1698)));
    layer6_outputs(3856) <= layer5_outputs(4873);
    layer6_outputs(3857) <= '0';
    layer6_outputs(3858) <= not((layer5_outputs(686)) xor (layer5_outputs(3263)));
    layer6_outputs(3859) <= (layer5_outputs(2909)) and not (layer5_outputs(1989));
    layer6_outputs(3860) <= not((layer5_outputs(2572)) xor (layer5_outputs(1700)));
    layer6_outputs(3861) <= layer5_outputs(4264);
    layer6_outputs(3862) <= (layer5_outputs(727)) or (layer5_outputs(1228));
    layer6_outputs(3863) <= layer5_outputs(4463);
    layer6_outputs(3864) <= not(layer5_outputs(1756)) or (layer5_outputs(937));
    layer6_outputs(3865) <= not(layer5_outputs(4402));
    layer6_outputs(3866) <= layer5_outputs(2444);
    layer6_outputs(3867) <= not(layer5_outputs(2283));
    layer6_outputs(3868) <= (layer5_outputs(4266)) and not (layer5_outputs(1090));
    layer6_outputs(3869) <= '0';
    layer6_outputs(3870) <= (layer5_outputs(5058)) and not (layer5_outputs(5074));
    layer6_outputs(3871) <= not(layer5_outputs(2434)) or (layer5_outputs(3899));
    layer6_outputs(3872) <= layer5_outputs(4699);
    layer6_outputs(3873) <= (layer5_outputs(2324)) and not (layer5_outputs(4327));
    layer6_outputs(3874) <= not((layer5_outputs(4126)) and (layer5_outputs(2979)));
    layer6_outputs(3875) <= not((layer5_outputs(2395)) xor (layer5_outputs(2011)));
    layer6_outputs(3876) <= not(layer5_outputs(1994)) or (layer5_outputs(2273));
    layer6_outputs(3877) <= (layer5_outputs(4301)) xor (layer5_outputs(529));
    layer6_outputs(3878) <= layer5_outputs(750);
    layer6_outputs(3879) <= layer5_outputs(4555);
    layer6_outputs(3880) <= (layer5_outputs(1654)) and (layer5_outputs(1569));
    layer6_outputs(3881) <= not(layer5_outputs(2682)) or (layer5_outputs(3935));
    layer6_outputs(3882) <= not(layer5_outputs(2454)) or (layer5_outputs(1325));
    layer6_outputs(3883) <= (layer5_outputs(281)) and (layer5_outputs(4842));
    layer6_outputs(3884) <= '1';
    layer6_outputs(3885) <= layer5_outputs(2818);
    layer6_outputs(3886) <= (layer5_outputs(508)) and not (layer5_outputs(4871));
    layer6_outputs(3887) <= layer5_outputs(4032);
    layer6_outputs(3888) <= not(layer5_outputs(4959));
    layer6_outputs(3889) <= (layer5_outputs(2702)) or (layer5_outputs(385));
    layer6_outputs(3890) <= (layer5_outputs(978)) xor (layer5_outputs(3365));
    layer6_outputs(3891) <= (layer5_outputs(2730)) and (layer5_outputs(319));
    layer6_outputs(3892) <= not((layer5_outputs(1220)) or (layer5_outputs(4585)));
    layer6_outputs(3893) <= layer5_outputs(806);
    layer6_outputs(3894) <= not(layer5_outputs(4874));
    layer6_outputs(3895) <= (layer5_outputs(2497)) xor (layer5_outputs(3225));
    layer6_outputs(3896) <= not((layer5_outputs(472)) xor (layer5_outputs(4573)));
    layer6_outputs(3897) <= layer5_outputs(4046);
    layer6_outputs(3898) <= (layer5_outputs(3639)) or (layer5_outputs(3296));
    layer6_outputs(3899) <= (layer5_outputs(2920)) and (layer5_outputs(591));
    layer6_outputs(3900) <= (layer5_outputs(3927)) xor (layer5_outputs(3238));
    layer6_outputs(3901) <= not(layer5_outputs(3562));
    layer6_outputs(3902) <= not(layer5_outputs(3776));
    layer6_outputs(3903) <= layer5_outputs(4083);
    layer6_outputs(3904) <= not(layer5_outputs(4954)) or (layer5_outputs(4571));
    layer6_outputs(3905) <= not((layer5_outputs(1970)) xor (layer5_outputs(56)));
    layer6_outputs(3906) <= not(layer5_outputs(289));
    layer6_outputs(3907) <= not(layer5_outputs(1206));
    layer6_outputs(3908) <= not((layer5_outputs(4326)) xor (layer5_outputs(3769)));
    layer6_outputs(3909) <= '1';
    layer6_outputs(3910) <= not(layer5_outputs(4183));
    layer6_outputs(3911) <= not((layer5_outputs(853)) or (layer5_outputs(1545)));
    layer6_outputs(3912) <= not((layer5_outputs(4929)) or (layer5_outputs(983)));
    layer6_outputs(3913) <= (layer5_outputs(1659)) or (layer5_outputs(3409));
    layer6_outputs(3914) <= not(layer5_outputs(710)) or (layer5_outputs(3295));
    layer6_outputs(3915) <= not(layer5_outputs(1868)) or (layer5_outputs(4695));
    layer6_outputs(3916) <= (layer5_outputs(2428)) and not (layer5_outputs(2449));
    layer6_outputs(3917) <= not(layer5_outputs(4156)) or (layer5_outputs(2190));
    layer6_outputs(3918) <= layer5_outputs(2141);
    layer6_outputs(3919) <= (layer5_outputs(776)) and not (layer5_outputs(2643));
    layer6_outputs(3920) <= not(layer5_outputs(3490));
    layer6_outputs(3921) <= (layer5_outputs(2941)) and not (layer5_outputs(227));
    layer6_outputs(3922) <= not(layer5_outputs(4425));
    layer6_outputs(3923) <= not(layer5_outputs(2283));
    layer6_outputs(3924) <= not(layer5_outputs(1638));
    layer6_outputs(3925) <= not(layer5_outputs(895)) or (layer5_outputs(3923));
    layer6_outputs(3926) <= (layer5_outputs(1230)) and (layer5_outputs(3006));
    layer6_outputs(3927) <= layer5_outputs(1118);
    layer6_outputs(3928) <= layer5_outputs(2442);
    layer6_outputs(3929) <= not(layer5_outputs(2507)) or (layer5_outputs(2321));
    layer6_outputs(3930) <= not(layer5_outputs(3785));
    layer6_outputs(3931) <= (layer5_outputs(2455)) xor (layer5_outputs(1905));
    layer6_outputs(3932) <= (layer5_outputs(4117)) or (layer5_outputs(617));
    layer6_outputs(3933) <= not(layer5_outputs(2417));
    layer6_outputs(3934) <= not(layer5_outputs(483));
    layer6_outputs(3935) <= layer5_outputs(1536);
    layer6_outputs(3936) <= layer5_outputs(3423);
    layer6_outputs(3937) <= not((layer5_outputs(2413)) or (layer5_outputs(186)));
    layer6_outputs(3938) <= layer5_outputs(2017);
    layer6_outputs(3939) <= not(layer5_outputs(3618)) or (layer5_outputs(2397));
    layer6_outputs(3940) <= not(layer5_outputs(4877));
    layer6_outputs(3941) <= (layer5_outputs(4241)) xor (layer5_outputs(2629));
    layer6_outputs(3942) <= not(layer5_outputs(2553)) or (layer5_outputs(4279));
    layer6_outputs(3943) <= layer5_outputs(1481);
    layer6_outputs(3944) <= not(layer5_outputs(4683)) or (layer5_outputs(4211));
    layer6_outputs(3945) <= (layer5_outputs(1888)) and not (layer5_outputs(2444));
    layer6_outputs(3946) <= '1';
    layer6_outputs(3947) <= not(layer5_outputs(4826));
    layer6_outputs(3948) <= not(layer5_outputs(4065));
    layer6_outputs(3949) <= not((layer5_outputs(2508)) or (layer5_outputs(2520)));
    layer6_outputs(3950) <= layer5_outputs(3756);
    layer6_outputs(3951) <= layer5_outputs(1200);
    layer6_outputs(3952) <= (layer5_outputs(3902)) xor (layer5_outputs(8));
    layer6_outputs(3953) <= (layer5_outputs(3598)) and (layer5_outputs(3409));
    layer6_outputs(3954) <= not(layer5_outputs(4325)) or (layer5_outputs(1001));
    layer6_outputs(3955) <= (layer5_outputs(2745)) xor (layer5_outputs(3583));
    layer6_outputs(3956) <= layer5_outputs(3299);
    layer6_outputs(3957) <= layer5_outputs(608);
    layer6_outputs(3958) <= (layer5_outputs(4054)) or (layer5_outputs(3848));
    layer6_outputs(3959) <= not(layer5_outputs(3638));
    layer6_outputs(3960) <= (layer5_outputs(3930)) and (layer5_outputs(4024));
    layer6_outputs(3961) <= not((layer5_outputs(850)) and (layer5_outputs(1375)));
    layer6_outputs(3962) <= (layer5_outputs(295)) and (layer5_outputs(3561));
    layer6_outputs(3963) <= not(layer5_outputs(173)) or (layer5_outputs(3679));
    layer6_outputs(3964) <= not((layer5_outputs(4815)) or (layer5_outputs(4661)));
    layer6_outputs(3965) <= not(layer5_outputs(931)) or (layer5_outputs(4212));
    layer6_outputs(3966) <= not(layer5_outputs(468)) or (layer5_outputs(359));
    layer6_outputs(3967) <= not(layer5_outputs(3360));
    layer6_outputs(3968) <= (layer5_outputs(231)) and not (layer5_outputs(567));
    layer6_outputs(3969) <= not((layer5_outputs(3517)) or (layer5_outputs(4975)));
    layer6_outputs(3970) <= layer5_outputs(219);
    layer6_outputs(3971) <= not((layer5_outputs(5084)) and (layer5_outputs(3837)));
    layer6_outputs(3972) <= not(layer5_outputs(3502));
    layer6_outputs(3973) <= layer5_outputs(3025);
    layer6_outputs(3974) <= not((layer5_outputs(42)) xor (layer5_outputs(1063)));
    layer6_outputs(3975) <= layer5_outputs(2386);
    layer6_outputs(3976) <= layer5_outputs(2545);
    layer6_outputs(3977) <= '1';
    layer6_outputs(3978) <= not((layer5_outputs(4982)) xor (layer5_outputs(4747)));
    layer6_outputs(3979) <= (layer5_outputs(1024)) and not (layer5_outputs(4261));
    layer6_outputs(3980) <= (layer5_outputs(3408)) xor (layer5_outputs(924));
    layer6_outputs(3981) <= not(layer5_outputs(2643));
    layer6_outputs(3982) <= (layer5_outputs(831)) and (layer5_outputs(5048));
    layer6_outputs(3983) <= layer5_outputs(2289);
    layer6_outputs(3984) <= not((layer5_outputs(1710)) xor (layer5_outputs(206)));
    layer6_outputs(3985) <= (layer5_outputs(702)) or (layer5_outputs(2081));
    layer6_outputs(3986) <= layer5_outputs(896);
    layer6_outputs(3987) <= not(layer5_outputs(4113));
    layer6_outputs(3988) <= not(layer5_outputs(1105));
    layer6_outputs(3989) <= layer5_outputs(911);
    layer6_outputs(3990) <= not((layer5_outputs(3191)) or (layer5_outputs(3381)));
    layer6_outputs(3991) <= not(layer5_outputs(1998));
    layer6_outputs(3992) <= '1';
    layer6_outputs(3993) <= (layer5_outputs(92)) and not (layer5_outputs(176));
    layer6_outputs(3994) <= '0';
    layer6_outputs(3995) <= not(layer5_outputs(1274)) or (layer5_outputs(1317));
    layer6_outputs(3996) <= not(layer5_outputs(4537));
    layer6_outputs(3997) <= (layer5_outputs(3119)) and not (layer5_outputs(1091));
    layer6_outputs(3998) <= '1';
    layer6_outputs(3999) <= (layer5_outputs(9)) xor (layer5_outputs(3267));
    layer6_outputs(4000) <= not((layer5_outputs(3250)) and (layer5_outputs(2195)));
    layer6_outputs(4001) <= (layer5_outputs(4675)) xor (layer5_outputs(4825));
    layer6_outputs(4002) <= (layer5_outputs(721)) and not (layer5_outputs(2536));
    layer6_outputs(4003) <= layer5_outputs(2166);
    layer6_outputs(4004) <= '1';
    layer6_outputs(4005) <= (layer5_outputs(1179)) and (layer5_outputs(4314));
    layer6_outputs(4006) <= layer5_outputs(1665);
    layer6_outputs(4007) <= not((layer5_outputs(849)) and (layer5_outputs(4766)));
    layer6_outputs(4008) <= not(layer5_outputs(1714));
    layer6_outputs(4009) <= not((layer5_outputs(2278)) xor (layer5_outputs(2289)));
    layer6_outputs(4010) <= (layer5_outputs(4703)) xor (layer5_outputs(4110));
    layer6_outputs(4011) <= (layer5_outputs(3014)) and not (layer5_outputs(4569));
    layer6_outputs(4012) <= layer5_outputs(5019);
    layer6_outputs(4013) <= not((layer5_outputs(3199)) xor (layer5_outputs(3175)));
    layer6_outputs(4014) <= '1';
    layer6_outputs(4015) <= not(layer5_outputs(535));
    layer6_outputs(4016) <= not(layer5_outputs(2748)) or (layer5_outputs(122));
    layer6_outputs(4017) <= layer5_outputs(1961);
    layer6_outputs(4018) <= not(layer5_outputs(1082));
    layer6_outputs(4019) <= layer5_outputs(4255);
    layer6_outputs(4020) <= layer5_outputs(4729);
    layer6_outputs(4021) <= layer5_outputs(3910);
    layer6_outputs(4022) <= (layer5_outputs(3665)) and not (layer5_outputs(3446));
    layer6_outputs(4023) <= layer5_outputs(3511);
    layer6_outputs(4024) <= not(layer5_outputs(880));
    layer6_outputs(4025) <= layer5_outputs(4043);
    layer6_outputs(4026) <= '1';
    layer6_outputs(4027) <= not((layer5_outputs(1910)) and (layer5_outputs(4773)));
    layer6_outputs(4028) <= '0';
    layer6_outputs(4029) <= not(layer5_outputs(1300));
    layer6_outputs(4030) <= (layer5_outputs(2867)) and not (layer5_outputs(2498));
    layer6_outputs(4031) <= layer5_outputs(1560);
    layer6_outputs(4032) <= (layer5_outputs(3872)) and not (layer5_outputs(292));
    layer6_outputs(4033) <= not((layer5_outputs(1739)) xor (layer5_outputs(4033)));
    layer6_outputs(4034) <= not(layer5_outputs(3039));
    layer6_outputs(4035) <= not(layer5_outputs(5116));
    layer6_outputs(4036) <= (layer5_outputs(2796)) and not (layer5_outputs(3157));
    layer6_outputs(4037) <= not((layer5_outputs(2523)) and (layer5_outputs(4646)));
    layer6_outputs(4038) <= (layer5_outputs(3135)) or (layer5_outputs(742));
    layer6_outputs(4039) <= layer5_outputs(3045);
    layer6_outputs(4040) <= not(layer5_outputs(2974)) or (layer5_outputs(3109));
    layer6_outputs(4041) <= (layer5_outputs(4271)) and not (layer5_outputs(4541));
    layer6_outputs(4042) <= (layer5_outputs(5012)) and (layer5_outputs(288));
    layer6_outputs(4043) <= not(layer5_outputs(362));
    layer6_outputs(4044) <= not((layer5_outputs(1501)) xor (layer5_outputs(157)));
    layer6_outputs(4045) <= (layer5_outputs(4853)) and not (layer5_outputs(4409));
    layer6_outputs(4046) <= (layer5_outputs(795)) and not (layer5_outputs(479));
    layer6_outputs(4047) <= not(layer5_outputs(4636));
    layer6_outputs(4048) <= layer5_outputs(583);
    layer6_outputs(4049) <= layer5_outputs(936);
    layer6_outputs(4050) <= (layer5_outputs(1963)) or (layer5_outputs(3669));
    layer6_outputs(4051) <= layer5_outputs(2219);
    layer6_outputs(4052) <= not(layer5_outputs(3784)) or (layer5_outputs(3453));
    layer6_outputs(4053) <= (layer5_outputs(3411)) or (layer5_outputs(5027));
    layer6_outputs(4054) <= not(layer5_outputs(4779));
    layer6_outputs(4055) <= not(layer5_outputs(1908)) or (layer5_outputs(1692));
    layer6_outputs(4056) <= not(layer5_outputs(1579)) or (layer5_outputs(4248));
    layer6_outputs(4057) <= (layer5_outputs(3719)) and not (layer5_outputs(2752));
    layer6_outputs(4058) <= not(layer5_outputs(1109));
    layer6_outputs(4059) <= layer5_outputs(1097);
    layer6_outputs(4060) <= not(layer5_outputs(523));
    layer6_outputs(4061) <= not(layer5_outputs(4185));
    layer6_outputs(4062) <= layer5_outputs(2184);
    layer6_outputs(4063) <= (layer5_outputs(3750)) and (layer5_outputs(877));
    layer6_outputs(4064) <= not(layer5_outputs(4009));
    layer6_outputs(4065) <= layer5_outputs(2686);
    layer6_outputs(4066) <= not((layer5_outputs(3976)) xor (layer5_outputs(4459)));
    layer6_outputs(4067) <= layer5_outputs(4592);
    layer6_outputs(4068) <= (layer5_outputs(3542)) or (layer5_outputs(2840));
    layer6_outputs(4069) <= (layer5_outputs(4688)) and (layer5_outputs(2094));
    layer6_outputs(4070) <= layer5_outputs(1567);
    layer6_outputs(4071) <= not(layer5_outputs(1770)) or (layer5_outputs(2896));
    layer6_outputs(4072) <= not(layer5_outputs(789));
    layer6_outputs(4073) <= not(layer5_outputs(4647)) or (layer5_outputs(2447));
    layer6_outputs(4074) <= not(layer5_outputs(2217)) or (layer5_outputs(4949));
    layer6_outputs(4075) <= not(layer5_outputs(1101));
    layer6_outputs(4076) <= (layer5_outputs(4278)) and (layer5_outputs(3845));
    layer6_outputs(4077) <= not(layer5_outputs(4272));
    layer6_outputs(4078) <= not(layer5_outputs(4084));
    layer6_outputs(4079) <= (layer5_outputs(797)) and not (layer5_outputs(2888));
    layer6_outputs(4080) <= layer5_outputs(2835);
    layer6_outputs(4081) <= not((layer5_outputs(1705)) and (layer5_outputs(2250)));
    layer6_outputs(4082) <= layer5_outputs(1201);
    layer6_outputs(4083) <= not((layer5_outputs(702)) and (layer5_outputs(2015)));
    layer6_outputs(4084) <= (layer5_outputs(4181)) and not (layer5_outputs(3069));
    layer6_outputs(4085) <= (layer5_outputs(2435)) and not (layer5_outputs(4536));
    layer6_outputs(4086) <= layer5_outputs(1439);
    layer6_outputs(4087) <= not(layer5_outputs(3342)) or (layer5_outputs(4407));
    layer6_outputs(4088) <= not((layer5_outputs(410)) xor (layer5_outputs(2335)));
    layer6_outputs(4089) <= layer5_outputs(3444);
    layer6_outputs(4090) <= (layer5_outputs(1286)) or (layer5_outputs(119));
    layer6_outputs(4091) <= not(layer5_outputs(3456)) or (layer5_outputs(4297));
    layer6_outputs(4092) <= layer5_outputs(2999);
    layer6_outputs(4093) <= (layer5_outputs(2560)) and not (layer5_outputs(4786));
    layer6_outputs(4094) <= (layer5_outputs(2732)) or (layer5_outputs(4975));
    layer6_outputs(4095) <= layer5_outputs(997);
    layer6_outputs(4096) <= not(layer5_outputs(1588)) or (layer5_outputs(4949));
    layer6_outputs(4097) <= not(layer5_outputs(1510));
    layer6_outputs(4098) <= not(layer5_outputs(2838));
    layer6_outputs(4099) <= (layer5_outputs(3290)) xor (layer5_outputs(1402));
    layer6_outputs(4100) <= layer5_outputs(3149);
    layer6_outputs(4101) <= layer5_outputs(1647);
    layer6_outputs(4102) <= layer5_outputs(1638);
    layer6_outputs(4103) <= (layer5_outputs(241)) and not (layer5_outputs(3689));
    layer6_outputs(4104) <= not(layer5_outputs(3888)) or (layer5_outputs(2960));
    layer6_outputs(4105) <= not((layer5_outputs(3923)) and (layer5_outputs(3217)));
    layer6_outputs(4106) <= layer5_outputs(1680);
    layer6_outputs(4107) <= '0';
    layer6_outputs(4108) <= layer5_outputs(1854);
    layer6_outputs(4109) <= not(layer5_outputs(3849));
    layer6_outputs(4110) <= layer5_outputs(5020);
    layer6_outputs(4111) <= (layer5_outputs(1478)) and not (layer5_outputs(3246));
    layer6_outputs(4112) <= not(layer5_outputs(4503)) or (layer5_outputs(4545));
    layer6_outputs(4113) <= not(layer5_outputs(1831)) or (layer5_outputs(1746));
    layer6_outputs(4114) <= not(layer5_outputs(1614));
    layer6_outputs(4115) <= '1';
    layer6_outputs(4116) <= (layer5_outputs(229)) or (layer5_outputs(4698));
    layer6_outputs(4117) <= (layer5_outputs(3070)) and not (layer5_outputs(1959));
    layer6_outputs(4118) <= not(layer5_outputs(4776));
    layer6_outputs(4119) <= not(layer5_outputs(1926)) or (layer5_outputs(31));
    layer6_outputs(4120) <= not(layer5_outputs(4684));
    layer6_outputs(4121) <= not(layer5_outputs(2241)) or (layer5_outputs(3426));
    layer6_outputs(4122) <= layer5_outputs(264);
    layer6_outputs(4123) <= not(layer5_outputs(792));
    layer6_outputs(4124) <= layer5_outputs(2657);
    layer6_outputs(4125) <= (layer5_outputs(2518)) or (layer5_outputs(507));
    layer6_outputs(4126) <= not(layer5_outputs(78)) or (layer5_outputs(110));
    layer6_outputs(4127) <= layer5_outputs(3197);
    layer6_outputs(4128) <= (layer5_outputs(2183)) and not (layer5_outputs(4037));
    layer6_outputs(4129) <= layer5_outputs(3211);
    layer6_outputs(4130) <= layer5_outputs(1562);
    layer6_outputs(4131) <= (layer5_outputs(689)) and (layer5_outputs(1072));
    layer6_outputs(4132) <= layer5_outputs(994);
    layer6_outputs(4133) <= not(layer5_outputs(2187));
    layer6_outputs(4134) <= layer5_outputs(3089);
    layer6_outputs(4135) <= (layer5_outputs(3278)) and not (layer5_outputs(3171));
    layer6_outputs(4136) <= layer5_outputs(2782);
    layer6_outputs(4137) <= layer5_outputs(4815);
    layer6_outputs(4138) <= layer5_outputs(3835);
    layer6_outputs(4139) <= not(layer5_outputs(1917));
    layer6_outputs(4140) <= layer5_outputs(3815);
    layer6_outputs(4141) <= not((layer5_outputs(2516)) and (layer5_outputs(612)));
    layer6_outputs(4142) <= not(layer5_outputs(4700));
    layer6_outputs(4143) <= not(layer5_outputs(4737));
    layer6_outputs(4144) <= (layer5_outputs(1305)) xor (layer5_outputs(1693));
    layer6_outputs(4145) <= layer5_outputs(3840);
    layer6_outputs(4146) <= '0';
    layer6_outputs(4147) <= not(layer5_outputs(4798));
    layer6_outputs(4148) <= not(layer5_outputs(2749)) or (layer5_outputs(2495));
    layer6_outputs(4149) <= (layer5_outputs(671)) and not (layer5_outputs(3380));
    layer6_outputs(4150) <= layer5_outputs(4278);
    layer6_outputs(4151) <= not(layer5_outputs(1830));
    layer6_outputs(4152) <= (layer5_outputs(150)) or (layer5_outputs(2589));
    layer6_outputs(4153) <= not(layer5_outputs(4436)) or (layer5_outputs(4600));
    layer6_outputs(4154) <= not(layer5_outputs(238));
    layer6_outputs(4155) <= not((layer5_outputs(559)) or (layer5_outputs(1249)));
    layer6_outputs(4156) <= (layer5_outputs(1294)) and not (layer5_outputs(1241));
    layer6_outputs(4157) <= (layer5_outputs(1596)) and not (layer5_outputs(4272));
    layer6_outputs(4158) <= (layer5_outputs(2087)) and (layer5_outputs(1351));
    layer6_outputs(4159) <= not(layer5_outputs(5051));
    layer6_outputs(4160) <= not((layer5_outputs(1147)) xor (layer5_outputs(1115)));
    layer6_outputs(4161) <= not((layer5_outputs(4848)) and (layer5_outputs(2534)));
    layer6_outputs(4162) <= not((layer5_outputs(4918)) xor (layer5_outputs(2435)));
    layer6_outputs(4163) <= (layer5_outputs(191)) xor (layer5_outputs(3173));
    layer6_outputs(4164) <= not(layer5_outputs(989)) or (layer5_outputs(3696));
    layer6_outputs(4165) <= layer5_outputs(3961);
    layer6_outputs(4166) <= '0';
    layer6_outputs(4167) <= layer5_outputs(4426);
    layer6_outputs(4168) <= not((layer5_outputs(1561)) xor (layer5_outputs(1331)));
    layer6_outputs(4169) <= layer5_outputs(4757);
    layer6_outputs(4170) <= not((layer5_outputs(3337)) and (layer5_outputs(720)));
    layer6_outputs(4171) <= '1';
    layer6_outputs(4172) <= not((layer5_outputs(3800)) and (layer5_outputs(3067)));
    layer6_outputs(4173) <= not(layer5_outputs(1563));
    layer6_outputs(4174) <= (layer5_outputs(2638)) or (layer5_outputs(4290));
    layer6_outputs(4175) <= layer5_outputs(2915);
    layer6_outputs(4176) <= (layer5_outputs(1536)) and (layer5_outputs(4460));
    layer6_outputs(4177) <= layer5_outputs(1122);
    layer6_outputs(4178) <= not((layer5_outputs(3850)) or (layer5_outputs(1856)));
    layer6_outputs(4179) <= (layer5_outputs(4374)) and (layer5_outputs(1015));
    layer6_outputs(4180) <= '1';
    layer6_outputs(4181) <= not(layer5_outputs(422));
    layer6_outputs(4182) <= layer5_outputs(4466);
    layer6_outputs(4183) <= (layer5_outputs(2860)) and (layer5_outputs(1750));
    layer6_outputs(4184) <= (layer5_outputs(4118)) xor (layer5_outputs(1731));
    layer6_outputs(4185) <= (layer5_outputs(2365)) xor (layer5_outputs(2413));
    layer6_outputs(4186) <= layer5_outputs(5070);
    layer6_outputs(4187) <= not(layer5_outputs(3626)) or (layer5_outputs(2479));
    layer6_outputs(4188) <= not(layer5_outputs(4357)) or (layer5_outputs(458));
    layer6_outputs(4189) <= not(layer5_outputs(3009));
    layer6_outputs(4190) <= layer5_outputs(3760);
    layer6_outputs(4191) <= layer5_outputs(960);
    layer6_outputs(4192) <= (layer5_outputs(597)) and not (layer5_outputs(2960));
    layer6_outputs(4193) <= layer5_outputs(1281);
    layer6_outputs(4194) <= not(layer5_outputs(4535)) or (layer5_outputs(1636));
    layer6_outputs(4195) <= layer5_outputs(1369);
    layer6_outputs(4196) <= (layer5_outputs(1598)) and (layer5_outputs(3694));
    layer6_outputs(4197) <= layer5_outputs(1371);
    layer6_outputs(4198) <= (layer5_outputs(837)) and (layer5_outputs(2597));
    layer6_outputs(4199) <= not((layer5_outputs(363)) or (layer5_outputs(4122)));
    layer6_outputs(4200) <= layer5_outputs(2468);
    layer6_outputs(4201) <= (layer5_outputs(444)) or (layer5_outputs(3399));
    layer6_outputs(4202) <= layer5_outputs(4073);
    layer6_outputs(4203) <= layer5_outputs(4809);
    layer6_outputs(4204) <= not((layer5_outputs(1219)) or (layer5_outputs(4280)));
    layer6_outputs(4205) <= layer5_outputs(3527);
    layer6_outputs(4206) <= layer5_outputs(3554);
    layer6_outputs(4207) <= layer5_outputs(2388);
    layer6_outputs(4208) <= not(layer5_outputs(2861));
    layer6_outputs(4209) <= layer5_outputs(677);
    layer6_outputs(4210) <= (layer5_outputs(3367)) and not (layer5_outputs(1284));
    layer6_outputs(4211) <= '0';
    layer6_outputs(4212) <= not(layer5_outputs(2542));
    layer6_outputs(4213) <= (layer5_outputs(3745)) or (layer5_outputs(3163));
    layer6_outputs(4214) <= not(layer5_outputs(3430));
    layer6_outputs(4215) <= not(layer5_outputs(4517));
    layer6_outputs(4216) <= not(layer5_outputs(3690)) or (layer5_outputs(2793));
    layer6_outputs(4217) <= not((layer5_outputs(631)) xor (layer5_outputs(3708)));
    layer6_outputs(4218) <= not((layer5_outputs(1982)) or (layer5_outputs(2798)));
    layer6_outputs(4219) <= not(layer5_outputs(1545));
    layer6_outputs(4220) <= not((layer5_outputs(1738)) or (layer5_outputs(1222)));
    layer6_outputs(4221) <= not(layer5_outputs(1984));
    layer6_outputs(4222) <= not((layer5_outputs(813)) and (layer5_outputs(2146)));
    layer6_outputs(4223) <= '1';
    layer6_outputs(4224) <= (layer5_outputs(2063)) and not (layer5_outputs(1029));
    layer6_outputs(4225) <= not((layer5_outputs(6)) and (layer5_outputs(3882)));
    layer6_outputs(4226) <= '1';
    layer6_outputs(4227) <= '1';
    layer6_outputs(4228) <= (layer5_outputs(1690)) and not (layer5_outputs(478));
    layer6_outputs(4229) <= not((layer5_outputs(2690)) and (layer5_outputs(3361)));
    layer6_outputs(4230) <= not((layer5_outputs(1319)) or (layer5_outputs(4589)));
    layer6_outputs(4231) <= '0';
    layer6_outputs(4232) <= (layer5_outputs(3293)) xor (layer5_outputs(2580));
    layer6_outputs(4233) <= not(layer5_outputs(4311));
    layer6_outputs(4234) <= not(layer5_outputs(2167));
    layer6_outputs(4235) <= not(layer5_outputs(1040));
    layer6_outputs(4236) <= layer5_outputs(1458);
    layer6_outputs(4237) <= not(layer5_outputs(3580));
    layer6_outputs(4238) <= layer5_outputs(2651);
    layer6_outputs(4239) <= layer5_outputs(33);
    layer6_outputs(4240) <= not((layer5_outputs(2016)) xor (layer5_outputs(4028)));
    layer6_outputs(4241) <= not(layer5_outputs(4875)) or (layer5_outputs(4454));
    layer6_outputs(4242) <= not((layer5_outputs(4200)) xor (layer5_outputs(2203)));
    layer6_outputs(4243) <= layer5_outputs(1603);
    layer6_outputs(4244) <= (layer5_outputs(2970)) or (layer5_outputs(4607));
    layer6_outputs(4245) <= not(layer5_outputs(1807));
    layer6_outputs(4246) <= (layer5_outputs(313)) and not (layer5_outputs(1711));
    layer6_outputs(4247) <= not(layer5_outputs(957));
    layer6_outputs(4248) <= layer5_outputs(79);
    layer6_outputs(4249) <= '0';
    layer6_outputs(4250) <= layer5_outputs(609);
    layer6_outputs(4251) <= (layer5_outputs(4497)) and not (layer5_outputs(448));
    layer6_outputs(4252) <= not(layer5_outputs(1763));
    layer6_outputs(4253) <= not(layer5_outputs(2851));
    layer6_outputs(4254) <= (layer5_outputs(2925)) and not (layer5_outputs(2650));
    layer6_outputs(4255) <= not(layer5_outputs(653));
    layer6_outputs(4256) <= not(layer5_outputs(956));
    layer6_outputs(4257) <= '0';
    layer6_outputs(4258) <= (layer5_outputs(3320)) and not (layer5_outputs(29));
    layer6_outputs(4259) <= '0';
    layer6_outputs(4260) <= not(layer5_outputs(3827)) or (layer5_outputs(766));
    layer6_outputs(4261) <= not((layer5_outputs(1361)) xor (layer5_outputs(283)));
    layer6_outputs(4262) <= '0';
    layer6_outputs(4263) <= layer5_outputs(1269);
    layer6_outputs(4264) <= not(layer5_outputs(3007));
    layer6_outputs(4265) <= not(layer5_outputs(953)) or (layer5_outputs(2839));
    layer6_outputs(4266) <= layer5_outputs(5030);
    layer6_outputs(4267) <= layer5_outputs(2254);
    layer6_outputs(4268) <= layer5_outputs(2605);
    layer6_outputs(4269) <= not((layer5_outputs(2797)) and (layer5_outputs(3561)));
    layer6_outputs(4270) <= not(layer5_outputs(4283));
    layer6_outputs(4271) <= not((layer5_outputs(496)) or (layer5_outputs(3128)));
    layer6_outputs(4272) <= not((layer5_outputs(2754)) and (layer5_outputs(690)));
    layer6_outputs(4273) <= not((layer5_outputs(2381)) xor (layer5_outputs(4063)));
    layer6_outputs(4274) <= not((layer5_outputs(4970)) or (layer5_outputs(1147)));
    layer6_outputs(4275) <= layer5_outputs(4912);
    layer6_outputs(4276) <= layer5_outputs(2881);
    layer6_outputs(4277) <= not((layer5_outputs(2544)) xor (layer5_outputs(2958)));
    layer6_outputs(4278) <= (layer5_outputs(1953)) or (layer5_outputs(4877));
    layer6_outputs(4279) <= layer5_outputs(4672);
    layer6_outputs(4280) <= not(layer5_outputs(4631));
    layer6_outputs(4281) <= not((layer5_outputs(4533)) or (layer5_outputs(1643)));
    layer6_outputs(4282) <= layer5_outputs(4220);
    layer6_outputs(4283) <= not(layer5_outputs(1554)) or (layer5_outputs(3165));
    layer6_outputs(4284) <= not(layer5_outputs(1387)) or (layer5_outputs(2527));
    layer6_outputs(4285) <= not((layer5_outputs(4289)) or (layer5_outputs(2620)));
    layer6_outputs(4286) <= not(layer5_outputs(659)) or (layer5_outputs(3654));
    layer6_outputs(4287) <= (layer5_outputs(4674)) xor (layer5_outputs(715));
    layer6_outputs(4288) <= not(layer5_outputs(3507));
    layer6_outputs(4289) <= '0';
    layer6_outputs(4290) <= layer5_outputs(4962);
    layer6_outputs(4291) <= not(layer5_outputs(2044)) or (layer5_outputs(584));
    layer6_outputs(4292) <= (layer5_outputs(3236)) and (layer5_outputs(2927));
    layer6_outputs(4293) <= (layer5_outputs(1595)) and (layer5_outputs(4237));
    layer6_outputs(4294) <= not(layer5_outputs(4655)) or (layer5_outputs(504));
    layer6_outputs(4295) <= not(layer5_outputs(5107));
    layer6_outputs(4296) <= layer5_outputs(4430);
    layer6_outputs(4297) <= not(layer5_outputs(2111));
    layer6_outputs(4298) <= '0';
    layer6_outputs(4299) <= (layer5_outputs(2851)) and (layer5_outputs(2421));
    layer6_outputs(4300) <= (layer5_outputs(447)) xor (layer5_outputs(1632));
    layer6_outputs(4301) <= (layer5_outputs(495)) and (layer5_outputs(744));
    layer6_outputs(4302) <= (layer5_outputs(4775)) and not (layer5_outputs(62));
    layer6_outputs(4303) <= not(layer5_outputs(152)) or (layer5_outputs(3904));
    layer6_outputs(4304) <= layer5_outputs(4976);
    layer6_outputs(4305) <= (layer5_outputs(1725)) and not (layer5_outputs(4207));
    layer6_outputs(4306) <= layer5_outputs(3799);
    layer6_outputs(4307) <= not(layer5_outputs(3326));
    layer6_outputs(4308) <= (layer5_outputs(2051)) and not (layer5_outputs(1132));
    layer6_outputs(4309) <= not(layer5_outputs(3786)) or (layer5_outputs(998));
    layer6_outputs(4310) <= not(layer5_outputs(1896)) or (layer5_outputs(2943));
    layer6_outputs(4311) <= layer5_outputs(3042);
    layer6_outputs(4312) <= '0';
    layer6_outputs(4313) <= not((layer5_outputs(635)) or (layer5_outputs(2356)));
    layer6_outputs(4314) <= not(layer5_outputs(2588));
    layer6_outputs(4315) <= (layer5_outputs(2657)) or (layer5_outputs(4269));
    layer6_outputs(4316) <= layer5_outputs(2205);
    layer6_outputs(4317) <= not((layer5_outputs(4601)) or (layer5_outputs(3581)));
    layer6_outputs(4318) <= not((layer5_outputs(3686)) xor (layer5_outputs(588)));
    layer6_outputs(4319) <= layer5_outputs(1454);
    layer6_outputs(4320) <= layer5_outputs(2670);
    layer6_outputs(4321) <= not(layer5_outputs(3729));
    layer6_outputs(4322) <= layer5_outputs(2646);
    layer6_outputs(4323) <= not(layer5_outputs(109)) or (layer5_outputs(3484));
    layer6_outputs(4324) <= (layer5_outputs(3758)) and not (layer5_outputs(515));
    layer6_outputs(4325) <= layer5_outputs(3098);
    layer6_outputs(4326) <= not(layer5_outputs(265)) or (layer5_outputs(150));
    layer6_outputs(4327) <= '1';
    layer6_outputs(4328) <= layer5_outputs(4440);
    layer6_outputs(4329) <= layer5_outputs(3390);
    layer6_outputs(4330) <= layer5_outputs(2302);
    layer6_outputs(4331) <= not((layer5_outputs(797)) xor (layer5_outputs(3580)));
    layer6_outputs(4332) <= (layer5_outputs(4662)) or (layer5_outputs(3470));
    layer6_outputs(4333) <= not((layer5_outputs(2181)) xor (layer5_outputs(3228)));
    layer6_outputs(4334) <= not(layer5_outputs(4722));
    layer6_outputs(4335) <= (layer5_outputs(1361)) or (layer5_outputs(2869));
    layer6_outputs(4336) <= layer5_outputs(3862);
    layer6_outputs(4337) <= '1';
    layer6_outputs(4338) <= not(layer5_outputs(3131)) or (layer5_outputs(893));
    layer6_outputs(4339) <= not(layer5_outputs(4523)) or (layer5_outputs(2405));
    layer6_outputs(4340) <= (layer5_outputs(2373)) and (layer5_outputs(1352));
    layer6_outputs(4341) <= not((layer5_outputs(2)) or (layer5_outputs(2875)));
    layer6_outputs(4342) <= not(layer5_outputs(2823)) or (layer5_outputs(3321));
    layer6_outputs(4343) <= '1';
    layer6_outputs(4344) <= layer5_outputs(4998);
    layer6_outputs(4345) <= not(layer5_outputs(4707));
    layer6_outputs(4346) <= layer5_outputs(2955);
    layer6_outputs(4347) <= layer5_outputs(2686);
    layer6_outputs(4348) <= layer5_outputs(402);
    layer6_outputs(4349) <= (layer5_outputs(4115)) or (layer5_outputs(830));
    layer6_outputs(4350) <= layer5_outputs(4425);
    layer6_outputs(4351) <= layer5_outputs(4265);
    layer6_outputs(4352) <= (layer5_outputs(3080)) or (layer5_outputs(4210));
    layer6_outputs(4353) <= (layer5_outputs(2636)) and not (layer5_outputs(4045));
    layer6_outputs(4354) <= not(layer5_outputs(3294));
    layer6_outputs(4355) <= not(layer5_outputs(2742));
    layer6_outputs(4356) <= layer5_outputs(1033);
    layer6_outputs(4357) <= not(layer5_outputs(1719));
    layer6_outputs(4358) <= '1';
    layer6_outputs(4359) <= (layer5_outputs(1392)) or (layer5_outputs(1564));
    layer6_outputs(4360) <= not(layer5_outputs(101));
    layer6_outputs(4361) <= layer5_outputs(4434);
    layer6_outputs(4362) <= not(layer5_outputs(3955));
    layer6_outputs(4363) <= layer5_outputs(4339);
    layer6_outputs(4364) <= not((layer5_outputs(1611)) or (layer5_outputs(3908)));
    layer6_outputs(4365) <= not(layer5_outputs(2188)) or (layer5_outputs(2795));
    layer6_outputs(4366) <= not((layer5_outputs(327)) xor (layer5_outputs(3227)));
    layer6_outputs(4367) <= (layer5_outputs(4262)) or (layer5_outputs(4710));
    layer6_outputs(4368) <= (layer5_outputs(1780)) and (layer5_outputs(1987));
    layer6_outputs(4369) <= not(layer5_outputs(2244)) or (layer5_outputs(3174));
    layer6_outputs(4370) <= not(layer5_outputs(2074));
    layer6_outputs(4371) <= '0';
    layer6_outputs(4372) <= not((layer5_outputs(303)) xor (layer5_outputs(2302)));
    layer6_outputs(4373) <= not(layer5_outputs(1785));
    layer6_outputs(4374) <= not(layer5_outputs(2825));
    layer6_outputs(4375) <= '0';
    layer6_outputs(4376) <= layer5_outputs(12);
    layer6_outputs(4377) <= not(layer5_outputs(3505));
    layer6_outputs(4378) <= '0';
    layer6_outputs(4379) <= not(layer5_outputs(3673));
    layer6_outputs(4380) <= layer5_outputs(2418);
    layer6_outputs(4381) <= layer5_outputs(3085);
    layer6_outputs(4382) <= not(layer5_outputs(2001)) or (layer5_outputs(3500));
    layer6_outputs(4383) <= '1';
    layer6_outputs(4384) <= not(layer5_outputs(2268)) or (layer5_outputs(2753));
    layer6_outputs(4385) <= not(layer5_outputs(4718));
    layer6_outputs(4386) <= layer5_outputs(1277);
    layer6_outputs(4387) <= (layer5_outputs(2228)) and (layer5_outputs(2804));
    layer6_outputs(4388) <= layer5_outputs(1122);
    layer6_outputs(4389) <= not((layer5_outputs(46)) or (layer5_outputs(2245)));
    layer6_outputs(4390) <= (layer5_outputs(1795)) or (layer5_outputs(2841));
    layer6_outputs(4391) <= layer5_outputs(2601);
    layer6_outputs(4392) <= (layer5_outputs(3387)) and not (layer5_outputs(4073));
    layer6_outputs(4393) <= layer5_outputs(3107);
    layer6_outputs(4394) <= layer5_outputs(2624);
    layer6_outputs(4395) <= layer5_outputs(4849);
    layer6_outputs(4396) <= not(layer5_outputs(4688));
    layer6_outputs(4397) <= not(layer5_outputs(3382));
    layer6_outputs(4398) <= layer5_outputs(643);
    layer6_outputs(4399) <= not(layer5_outputs(1363)) or (layer5_outputs(3512));
    layer6_outputs(4400) <= '0';
    layer6_outputs(4401) <= '1';
    layer6_outputs(4402) <= not(layer5_outputs(524));
    layer6_outputs(4403) <= not(layer5_outputs(3285)) or (layer5_outputs(1758));
    layer6_outputs(4404) <= not((layer5_outputs(4173)) xor (layer5_outputs(1456)));
    layer6_outputs(4405) <= (layer5_outputs(3419)) and (layer5_outputs(2967));
    layer6_outputs(4406) <= layer5_outputs(1494);
    layer6_outputs(4407) <= layer5_outputs(2940);
    layer6_outputs(4408) <= not((layer5_outputs(2983)) or (layer5_outputs(3550)));
    layer6_outputs(4409) <= (layer5_outputs(4228)) and not (layer5_outputs(2175));
    layer6_outputs(4410) <= (layer5_outputs(2427)) xor (layer5_outputs(3194));
    layer6_outputs(4411) <= not(layer5_outputs(1375));
    layer6_outputs(4412) <= layer5_outputs(3543);
    layer6_outputs(4413) <= layer5_outputs(3539);
    layer6_outputs(4414) <= (layer5_outputs(3220)) and not (layer5_outputs(1191));
    layer6_outputs(4415) <= not(layer5_outputs(493));
    layer6_outputs(4416) <= layer5_outputs(1201);
    layer6_outputs(4417) <= (layer5_outputs(3106)) xor (layer5_outputs(613));
    layer6_outputs(4418) <= (layer5_outputs(3168)) xor (layer5_outputs(4503));
    layer6_outputs(4419) <= (layer5_outputs(1135)) or (layer5_outputs(3476));
    layer6_outputs(4420) <= (layer5_outputs(3977)) and not (layer5_outputs(5035));
    layer6_outputs(4421) <= (layer5_outputs(4372)) xor (layer5_outputs(396));
    layer6_outputs(4422) <= (layer5_outputs(668)) and not (layer5_outputs(2949));
    layer6_outputs(4423) <= (layer5_outputs(3874)) and not (layer5_outputs(3943));
    layer6_outputs(4424) <= not((layer5_outputs(5073)) and (layer5_outputs(2260)));
    layer6_outputs(4425) <= layer5_outputs(2150);
    layer6_outputs(4426) <= (layer5_outputs(879)) and (layer5_outputs(4192));
    layer6_outputs(4427) <= '0';
    layer6_outputs(4428) <= (layer5_outputs(2235)) and not (layer5_outputs(2031));
    layer6_outputs(4429) <= layer5_outputs(3271);
    layer6_outputs(4430) <= '1';
    layer6_outputs(4431) <= layer5_outputs(3067);
    layer6_outputs(4432) <= not((layer5_outputs(1928)) xor (layer5_outputs(2003)));
    layer6_outputs(4433) <= (layer5_outputs(4739)) and not (layer5_outputs(2478));
    layer6_outputs(4434) <= (layer5_outputs(2798)) and not (layer5_outputs(918));
    layer6_outputs(4435) <= layer5_outputs(602);
    layer6_outputs(4436) <= (layer5_outputs(2573)) and (layer5_outputs(3404));
    layer6_outputs(4437) <= not(layer5_outputs(4485));
    layer6_outputs(4438) <= (layer5_outputs(3516)) and not (layer5_outputs(564));
    layer6_outputs(4439) <= not(layer5_outputs(1381)) or (layer5_outputs(1886));
    layer6_outputs(4440) <= '0';
    layer6_outputs(4441) <= layer5_outputs(1267);
    layer6_outputs(4442) <= layer5_outputs(466);
    layer6_outputs(4443) <= (layer5_outputs(2292)) or (layer5_outputs(2654));
    layer6_outputs(4444) <= not(layer5_outputs(708));
    layer6_outputs(4445) <= layer5_outputs(767);
    layer6_outputs(4446) <= not(layer5_outputs(2348));
    layer6_outputs(4447) <= (layer5_outputs(1260)) and (layer5_outputs(752));
    layer6_outputs(4448) <= not((layer5_outputs(3334)) or (layer5_outputs(1632)));
    layer6_outputs(4449) <= not(layer5_outputs(4485));
    layer6_outputs(4450) <= not((layer5_outputs(4824)) or (layer5_outputs(4382)));
    layer6_outputs(4451) <= not(layer5_outputs(2923));
    layer6_outputs(4452) <= not(layer5_outputs(4402));
    layer6_outputs(4453) <= (layer5_outputs(3268)) and (layer5_outputs(759));
    layer6_outputs(4454) <= not(layer5_outputs(4733));
    layer6_outputs(4455) <= (layer5_outputs(408)) and not (layer5_outputs(4458));
    layer6_outputs(4456) <= (layer5_outputs(4387)) and (layer5_outputs(2122));
    layer6_outputs(4457) <= layer5_outputs(3555);
    layer6_outputs(4458) <= not(layer5_outputs(1771));
    layer6_outputs(4459) <= (layer5_outputs(343)) and not (layer5_outputs(3936));
    layer6_outputs(4460) <= not(layer5_outputs(1526)) or (layer5_outputs(1890));
    layer6_outputs(4461) <= not(layer5_outputs(4924)) or (layer5_outputs(809));
    layer6_outputs(4462) <= (layer5_outputs(2168)) and (layer5_outputs(5006));
    layer6_outputs(4463) <= not(layer5_outputs(3786));
    layer6_outputs(4464) <= (layer5_outputs(2704)) and not (layer5_outputs(4984));
    layer6_outputs(4465) <= layer5_outputs(1793);
    layer6_outputs(4466) <= layer5_outputs(4486);
    layer6_outputs(4467) <= (layer5_outputs(2535)) and not (layer5_outputs(3766));
    layer6_outputs(4468) <= (layer5_outputs(4373)) or (layer5_outputs(120));
    layer6_outputs(4469) <= (layer5_outputs(791)) and not (layer5_outputs(3597));
    layer6_outputs(4470) <= not(layer5_outputs(2760));
    layer6_outputs(4471) <= not(layer5_outputs(4701));
    layer6_outputs(4472) <= (layer5_outputs(2757)) xor (layer5_outputs(675));
    layer6_outputs(4473) <= (layer5_outputs(3165)) xor (layer5_outputs(1225));
    layer6_outputs(4474) <= not((layer5_outputs(4912)) or (layer5_outputs(4549)));
    layer6_outputs(4475) <= not(layer5_outputs(3783));
    layer6_outputs(4476) <= layer5_outputs(4287);
    layer6_outputs(4477) <= not((layer5_outputs(3582)) xor (layer5_outputs(2799)));
    layer6_outputs(4478) <= not(layer5_outputs(2206));
    layer6_outputs(4479) <= layer5_outputs(4150);
    layer6_outputs(4480) <= (layer5_outputs(3123)) xor (layer5_outputs(3417));
    layer6_outputs(4481) <= layer5_outputs(1599);
    layer6_outputs(4482) <= (layer5_outputs(51)) and (layer5_outputs(1690));
    layer6_outputs(4483) <= not(layer5_outputs(2423));
    layer6_outputs(4484) <= not(layer5_outputs(3827));
    layer6_outputs(4485) <= not(layer5_outputs(2433));
    layer6_outputs(4486) <= not(layer5_outputs(808)) or (layer5_outputs(1896));
    layer6_outputs(4487) <= (layer5_outputs(894)) and (layer5_outputs(2600));
    layer6_outputs(4488) <= layer5_outputs(2309);
    layer6_outputs(4489) <= not(layer5_outputs(4694));
    layer6_outputs(4490) <= (layer5_outputs(3878)) and (layer5_outputs(302));
    layer6_outputs(4491) <= not(layer5_outputs(639));
    layer6_outputs(4492) <= (layer5_outputs(3770)) and not (layer5_outputs(447));
    layer6_outputs(4493) <= not(layer5_outputs(4151));
    layer6_outputs(4494) <= (layer5_outputs(1815)) xor (layer5_outputs(862));
    layer6_outputs(4495) <= (layer5_outputs(1656)) xor (layer5_outputs(2126));
    layer6_outputs(4496) <= (layer5_outputs(611)) and (layer5_outputs(1958));
    layer6_outputs(4497) <= layer5_outputs(877);
    layer6_outputs(4498) <= layer5_outputs(2159);
    layer6_outputs(4499) <= (layer5_outputs(2402)) and not (layer5_outputs(2209));
    layer6_outputs(4500) <= '0';
    layer6_outputs(4501) <= layer5_outputs(4119);
    layer6_outputs(4502) <= layer5_outputs(4125);
    layer6_outputs(4503) <= layer5_outputs(9);
    layer6_outputs(4504) <= not(layer5_outputs(1391));
    layer6_outputs(4505) <= layer5_outputs(1157);
    layer6_outputs(4506) <= (layer5_outputs(846)) and not (layer5_outputs(1377));
    layer6_outputs(4507) <= '1';
    layer6_outputs(4508) <= layer5_outputs(1952);
    layer6_outputs(4509) <= layer5_outputs(4753);
    layer6_outputs(4510) <= (layer5_outputs(4374)) or (layer5_outputs(3559));
    layer6_outputs(4511) <= (layer5_outputs(2354)) and (layer5_outputs(4144));
    layer6_outputs(4512) <= (layer5_outputs(2756)) and not (layer5_outputs(2158));
    layer6_outputs(4513) <= '1';
    layer6_outputs(4514) <= not(layer5_outputs(3045)) or (layer5_outputs(1927));
    layer6_outputs(4515) <= '0';
    layer6_outputs(4516) <= layer5_outputs(4615);
    layer6_outputs(4517) <= layer5_outputs(4585);
    layer6_outputs(4518) <= (layer5_outputs(660)) or (layer5_outputs(1951));
    layer6_outputs(4519) <= (layer5_outputs(2426)) xor (layer5_outputs(566));
    layer6_outputs(4520) <= layer5_outputs(2693);
    layer6_outputs(4521) <= layer5_outputs(159);
    layer6_outputs(4522) <= layer5_outputs(4336);
    layer6_outputs(4523) <= (layer5_outputs(2859)) and (layer5_outputs(3932));
    layer6_outputs(4524) <= (layer5_outputs(1636)) or (layer5_outputs(4317));
    layer6_outputs(4525) <= (layer5_outputs(1180)) and (layer5_outputs(4294));
    layer6_outputs(4526) <= not((layer5_outputs(700)) and (layer5_outputs(2029)));
    layer6_outputs(4527) <= (layer5_outputs(4738)) or (layer5_outputs(3169));
    layer6_outputs(4528) <= not(layer5_outputs(2934));
    layer6_outputs(4529) <= (layer5_outputs(4634)) and not (layer5_outputs(1950));
    layer6_outputs(4530) <= layer5_outputs(326);
    layer6_outputs(4531) <= not(layer5_outputs(3966));
    layer6_outputs(4532) <= layer5_outputs(2360);
    layer6_outputs(4533) <= layer5_outputs(1347);
    layer6_outputs(4534) <= not(layer5_outputs(75));
    layer6_outputs(4535) <= layer5_outputs(4844);
    layer6_outputs(4536) <= not(layer5_outputs(4353));
    layer6_outputs(4537) <= not(layer5_outputs(2113)) or (layer5_outputs(2598));
    layer6_outputs(4538) <= not(layer5_outputs(1702));
    layer6_outputs(4539) <= layer5_outputs(1503);
    layer6_outputs(4540) <= '1';
    layer6_outputs(4541) <= (layer5_outputs(2922)) or (layer5_outputs(3281));
    layer6_outputs(4542) <= not(layer5_outputs(4245)) or (layer5_outputs(315));
    layer6_outputs(4543) <= (layer5_outputs(4896)) or (layer5_outputs(1758));
    layer6_outputs(4544) <= (layer5_outputs(326)) and not (layer5_outputs(63));
    layer6_outputs(4545) <= (layer5_outputs(4508)) and (layer5_outputs(3416));
    layer6_outputs(4546) <= not((layer5_outputs(1191)) xor (layer5_outputs(5011)));
    layer6_outputs(4547) <= not(layer5_outputs(1818));
    layer6_outputs(4548) <= layer5_outputs(3005);
    layer6_outputs(4549) <= (layer5_outputs(2392)) or (layer5_outputs(1087));
    layer6_outputs(4550) <= (layer5_outputs(4227)) and not (layer5_outputs(2646));
    layer6_outputs(4551) <= not(layer5_outputs(871));
    layer6_outputs(4552) <= not(layer5_outputs(1229));
    layer6_outputs(4553) <= (layer5_outputs(4132)) or (layer5_outputs(3091));
    layer6_outputs(4554) <= layer5_outputs(4290);
    layer6_outputs(4555) <= not(layer5_outputs(2742));
    layer6_outputs(4556) <= '0';
    layer6_outputs(4557) <= '0';
    layer6_outputs(4558) <= layer5_outputs(4186);
    layer6_outputs(4559) <= (layer5_outputs(502)) or (layer5_outputs(4157));
    layer6_outputs(4560) <= not(layer5_outputs(463));
    layer6_outputs(4561) <= (layer5_outputs(1958)) xor (layer5_outputs(1902));
    layer6_outputs(4562) <= not(layer5_outputs(1082)) or (layer5_outputs(3592));
    layer6_outputs(4563) <= layer5_outputs(1739);
    layer6_outputs(4564) <= layer5_outputs(802);
    layer6_outputs(4565) <= layer5_outputs(278);
    layer6_outputs(4566) <= (layer5_outputs(2116)) and not (layer5_outputs(2722));
    layer6_outputs(4567) <= not(layer5_outputs(667));
    layer6_outputs(4568) <= layer5_outputs(1523);
    layer6_outputs(4569) <= (layer5_outputs(2942)) and not (layer5_outputs(1494));
    layer6_outputs(4570) <= not(layer5_outputs(3557)) or (layer5_outputs(1703));
    layer6_outputs(4571) <= not((layer5_outputs(3086)) and (layer5_outputs(245)));
    layer6_outputs(4572) <= layer5_outputs(4811);
    layer6_outputs(4573) <= (layer5_outputs(2892)) and (layer5_outputs(211));
    layer6_outputs(4574) <= not(layer5_outputs(1957));
    layer6_outputs(4575) <= not(layer5_outputs(3034));
    layer6_outputs(4576) <= layer5_outputs(3787);
    layer6_outputs(4577) <= not(layer5_outputs(3437)) or (layer5_outputs(933));
    layer6_outputs(4578) <= (layer5_outputs(2279)) and not (layer5_outputs(75));
    layer6_outputs(4579) <= not((layer5_outputs(5072)) or (layer5_outputs(3301)));
    layer6_outputs(4580) <= not(layer5_outputs(4348));
    layer6_outputs(4581) <= layer5_outputs(2254);
    layer6_outputs(4582) <= not(layer5_outputs(281)) or (layer5_outputs(4578));
    layer6_outputs(4583) <= (layer5_outputs(1388)) xor (layer5_outputs(1651));
    layer6_outputs(4584) <= not((layer5_outputs(2508)) xor (layer5_outputs(2135)));
    layer6_outputs(4585) <= not(layer5_outputs(1023));
    layer6_outputs(4586) <= not(layer5_outputs(865));
    layer6_outputs(4587) <= not(layer5_outputs(1697));
    layer6_outputs(4588) <= layer5_outputs(243);
    layer6_outputs(4589) <= not(layer5_outputs(4649));
    layer6_outputs(4590) <= layer5_outputs(820);
    layer6_outputs(4591) <= layer5_outputs(4099);
    layer6_outputs(4592) <= (layer5_outputs(4274)) or (layer5_outputs(2307));
    layer6_outputs(4593) <= not(layer5_outputs(2855)) or (layer5_outputs(3188));
    layer6_outputs(4594) <= not(layer5_outputs(410));
    layer6_outputs(4595) <= (layer5_outputs(4110)) and (layer5_outputs(1760));
    layer6_outputs(4596) <= not(layer5_outputs(4821));
    layer6_outputs(4597) <= not(layer5_outputs(152)) or (layer5_outputs(4149));
    layer6_outputs(4598) <= not(layer5_outputs(3123));
    layer6_outputs(4599) <= not(layer5_outputs(3688)) or (layer5_outputs(2627));
    layer6_outputs(4600) <= not(layer5_outputs(2012)) or (layer5_outputs(1384));
    layer6_outputs(4601) <= not(layer5_outputs(293)) or (layer5_outputs(4343));
    layer6_outputs(4602) <= layer5_outputs(3732);
    layer6_outputs(4603) <= not(layer5_outputs(640));
    layer6_outputs(4604) <= not(layer5_outputs(4754)) or (layer5_outputs(3917));
    layer6_outputs(4605) <= (layer5_outputs(3591)) or (layer5_outputs(3978));
    layer6_outputs(4606) <= (layer5_outputs(743)) and not (layer5_outputs(3552));
    layer6_outputs(4607) <= not(layer5_outputs(1092)) or (layer5_outputs(1937));
    layer6_outputs(4608) <= '1';
    layer6_outputs(4609) <= not((layer5_outputs(1564)) or (layer5_outputs(2894)));
    layer6_outputs(4610) <= not(layer5_outputs(311));
    layer6_outputs(4611) <= not(layer5_outputs(3810));
    layer6_outputs(4612) <= (layer5_outputs(716)) and not (layer5_outputs(2839));
    layer6_outputs(4613) <= layer5_outputs(69);
    layer6_outputs(4614) <= (layer5_outputs(592)) and not (layer5_outputs(1894));
    layer6_outputs(4615) <= not(layer5_outputs(2996));
    layer6_outputs(4616) <= not(layer5_outputs(318));
    layer6_outputs(4617) <= layer5_outputs(5068);
    layer6_outputs(4618) <= not(layer5_outputs(3215)) or (layer5_outputs(2600));
    layer6_outputs(4619) <= (layer5_outputs(4695)) and (layer5_outputs(1934));
    layer6_outputs(4620) <= not((layer5_outputs(3046)) and (layer5_outputs(545)));
    layer6_outputs(4621) <= not((layer5_outputs(1909)) and (layer5_outputs(3060)));
    layer6_outputs(4622) <= (layer5_outputs(4862)) and (layer5_outputs(4809));
    layer6_outputs(4623) <= (layer5_outputs(1339)) xor (layer5_outputs(3979));
    layer6_outputs(4624) <= not((layer5_outputs(3839)) or (layer5_outputs(647)));
    layer6_outputs(4625) <= not((layer5_outputs(2255)) or (layer5_outputs(4344)));
    layer6_outputs(4626) <= not(layer5_outputs(89));
    layer6_outputs(4627) <= (layer5_outputs(3789)) and not (layer5_outputs(3656));
    layer6_outputs(4628) <= layer5_outputs(2684);
    layer6_outputs(4629) <= layer5_outputs(3959);
    layer6_outputs(4630) <= not(layer5_outputs(310));
    layer6_outputs(4631) <= not(layer5_outputs(3963));
    layer6_outputs(4632) <= not(layer5_outputs(1196)) or (layer5_outputs(1587));
    layer6_outputs(4633) <= not(layer5_outputs(4111)) or (layer5_outputs(3466));
    layer6_outputs(4634) <= layer5_outputs(2035);
    layer6_outputs(4635) <= not(layer5_outputs(1644));
    layer6_outputs(4636) <= not(layer5_outputs(2118));
    layer6_outputs(4637) <= layer5_outputs(3959);
    layer6_outputs(4638) <= not((layer5_outputs(972)) and (layer5_outputs(4332)));
    layer6_outputs(4639) <= layer5_outputs(4247);
    layer6_outputs(4640) <= '0';
    layer6_outputs(4641) <= not(layer5_outputs(2087)) or (layer5_outputs(3813));
    layer6_outputs(4642) <= (layer5_outputs(2116)) or (layer5_outputs(3097));
    layer6_outputs(4643) <= (layer5_outputs(5021)) and (layer5_outputs(3119));
    layer6_outputs(4644) <= layer5_outputs(4181);
    layer6_outputs(4645) <= '0';
    layer6_outputs(4646) <= not(layer5_outputs(3831)) or (layer5_outputs(3208));
    layer6_outputs(4647) <= not((layer5_outputs(5066)) or (layer5_outputs(2530)));
    layer6_outputs(4648) <= (layer5_outputs(3290)) and not (layer5_outputs(3834));
    layer6_outputs(4649) <= not((layer5_outputs(50)) or (layer5_outputs(1789)));
    layer6_outputs(4650) <= not((layer5_outputs(4500)) or (layer5_outputs(4713)));
    layer6_outputs(4651) <= not((layer5_outputs(4030)) xor (layer5_outputs(2179)));
    layer6_outputs(4652) <= layer5_outputs(2380);
    layer6_outputs(4653) <= layer5_outputs(162);
    layer6_outputs(4654) <= not(layer5_outputs(1879));
    layer6_outputs(4655) <= not(layer5_outputs(174));
    layer6_outputs(4656) <= (layer5_outputs(652)) and not (layer5_outputs(3857));
    layer6_outputs(4657) <= layer5_outputs(1438);
    layer6_outputs(4658) <= not(layer5_outputs(4908));
    layer6_outputs(4659) <= not(layer5_outputs(4302));
    layer6_outputs(4660) <= not(layer5_outputs(5089));
    layer6_outputs(4661) <= not(layer5_outputs(127));
    layer6_outputs(4662) <= (layer5_outputs(1782)) and not (layer5_outputs(4338));
    layer6_outputs(4663) <= not(layer5_outputs(2483)) or (layer5_outputs(3150));
    layer6_outputs(4664) <= not((layer5_outputs(3628)) xor (layer5_outputs(489)));
    layer6_outputs(4665) <= layer5_outputs(3577);
    layer6_outputs(4666) <= not(layer5_outputs(2117)) or (layer5_outputs(1318));
    layer6_outputs(4667) <= not((layer5_outputs(2437)) or (layer5_outputs(1488)));
    layer6_outputs(4668) <= not(layer5_outputs(3681)) or (layer5_outputs(1210));
    layer6_outputs(4669) <= (layer5_outputs(4529)) and (layer5_outputs(16));
    layer6_outputs(4670) <= not((layer5_outputs(1238)) or (layer5_outputs(414)));
    layer6_outputs(4671) <= not(layer5_outputs(4495)) or (layer5_outputs(11));
    layer6_outputs(4672) <= not(layer5_outputs(2783));
    layer6_outputs(4673) <= (layer5_outputs(1767)) and not (layer5_outputs(2746));
    layer6_outputs(4674) <= (layer5_outputs(1681)) xor (layer5_outputs(27));
    layer6_outputs(4675) <= (layer5_outputs(609)) and (layer5_outputs(1582));
    layer6_outputs(4676) <= (layer5_outputs(1323)) and (layer5_outputs(1386));
    layer6_outputs(4677) <= not((layer5_outputs(3114)) and (layer5_outputs(1119)));
    layer6_outputs(4678) <= layer5_outputs(1650);
    layer6_outputs(4679) <= not((layer5_outputs(3792)) or (layer5_outputs(2295)));
    layer6_outputs(4680) <= not(layer5_outputs(3451));
    layer6_outputs(4681) <= layer5_outputs(1154);
    layer6_outputs(4682) <= (layer5_outputs(2477)) or (layer5_outputs(704));
    layer6_outputs(4683) <= (layer5_outputs(1529)) xor (layer5_outputs(5034));
    layer6_outputs(4684) <= not(layer5_outputs(1293));
    layer6_outputs(4685) <= not(layer5_outputs(3676));
    layer6_outputs(4686) <= (layer5_outputs(124)) and (layer5_outputs(2128));
    layer6_outputs(4687) <= (layer5_outputs(1634)) and (layer5_outputs(1237));
    layer6_outputs(4688) <= layer5_outputs(1563);
    layer6_outputs(4689) <= not(layer5_outputs(4926));
    layer6_outputs(4690) <= layer5_outputs(2789);
    layer6_outputs(4691) <= layer5_outputs(13);
    layer6_outputs(4692) <= (layer5_outputs(399)) and not (layer5_outputs(4658));
    layer6_outputs(4693) <= '1';
    layer6_outputs(4694) <= not((layer5_outputs(4068)) or (layer5_outputs(618)));
    layer6_outputs(4695) <= not((layer5_outputs(4247)) and (layer5_outputs(2488)));
    layer6_outputs(4696) <= '0';
    layer6_outputs(4697) <= not((layer5_outputs(2513)) or (layer5_outputs(3717)));
    layer6_outputs(4698) <= (layer5_outputs(3213)) and not (layer5_outputs(2975));
    layer6_outputs(4699) <= (layer5_outputs(4618)) and (layer5_outputs(225));
    layer6_outputs(4700) <= (layer5_outputs(1066)) and (layer5_outputs(4204));
    layer6_outputs(4701) <= not((layer5_outputs(2406)) or (layer5_outputs(456)));
    layer6_outputs(4702) <= (layer5_outputs(2708)) and not (layer5_outputs(5080));
    layer6_outputs(4703) <= not((layer5_outputs(1358)) or (layer5_outputs(1818)));
    layer6_outputs(4704) <= not((layer5_outputs(489)) or (layer5_outputs(2875)));
    layer6_outputs(4705) <= (layer5_outputs(153)) and not (layer5_outputs(250));
    layer6_outputs(4706) <= not((layer5_outputs(2108)) xor (layer5_outputs(2791)));
    layer6_outputs(4707) <= layer5_outputs(730);
    layer6_outputs(4708) <= layer5_outputs(3660);
    layer6_outputs(4709) <= (layer5_outputs(1779)) and not (layer5_outputs(403));
    layer6_outputs(4710) <= (layer5_outputs(3437)) xor (layer5_outputs(3720));
    layer6_outputs(4711) <= '0';
    layer6_outputs(4712) <= not((layer5_outputs(1072)) and (layer5_outputs(3902)));
    layer6_outputs(4713) <= layer5_outputs(3516);
    layer6_outputs(4714) <= layer5_outputs(1710);
    layer6_outputs(4715) <= layer5_outputs(4378);
    layer6_outputs(4716) <= not((layer5_outputs(3398)) xor (layer5_outputs(2058)));
    layer6_outputs(4717) <= layer5_outputs(2916);
    layer6_outputs(4718) <= (layer5_outputs(1845)) and not (layer5_outputs(2787));
    layer6_outputs(4719) <= not(layer5_outputs(1552));
    layer6_outputs(4720) <= (layer5_outputs(220)) and not (layer5_outputs(1615));
    layer6_outputs(4721) <= layer5_outputs(2899);
    layer6_outputs(4722) <= (layer5_outputs(1661)) and (layer5_outputs(5014));
    layer6_outputs(4723) <= (layer5_outputs(2599)) xor (layer5_outputs(2897));
    layer6_outputs(4724) <= not(layer5_outputs(312));
    layer6_outputs(4725) <= (layer5_outputs(4913)) and not (layer5_outputs(1236));
    layer6_outputs(4726) <= not(layer5_outputs(818));
    layer6_outputs(4727) <= not(layer5_outputs(2094));
    layer6_outputs(4728) <= not((layer5_outputs(4365)) xor (layer5_outputs(2613)));
    layer6_outputs(4729) <= not((layer5_outputs(2256)) and (layer5_outputs(3345)));
    layer6_outputs(4730) <= not((layer5_outputs(2333)) and (layer5_outputs(2944)));
    layer6_outputs(4731) <= not(layer5_outputs(4335));
    layer6_outputs(4732) <= layer5_outputs(4738);
    layer6_outputs(4733) <= layer5_outputs(2214);
    layer6_outputs(4734) <= '1';
    layer6_outputs(4735) <= not(layer5_outputs(4079));
    layer6_outputs(4736) <= not(layer5_outputs(3161)) or (layer5_outputs(1547));
    layer6_outputs(4737) <= '1';
    layer6_outputs(4738) <= not(layer5_outputs(2943)) or (layer5_outputs(2532));
    layer6_outputs(4739) <= not(layer5_outputs(831)) or (layer5_outputs(1975));
    layer6_outputs(4740) <= not((layer5_outputs(649)) and (layer5_outputs(975)));
    layer6_outputs(4741) <= not(layer5_outputs(347)) or (layer5_outputs(1783));
    layer6_outputs(4742) <= (layer5_outputs(4571)) and not (layer5_outputs(4582));
    layer6_outputs(4743) <= not(layer5_outputs(4388)) or (layer5_outputs(4));
    layer6_outputs(4744) <= not(layer5_outputs(4303));
    layer6_outputs(4745) <= not(layer5_outputs(4080)) or (layer5_outputs(1024));
    layer6_outputs(4746) <= '0';
    layer6_outputs(4747) <= (layer5_outputs(3009)) or (layer5_outputs(3477));
    layer6_outputs(4748) <= '0';
    layer6_outputs(4749) <= not(layer5_outputs(3157));
    layer6_outputs(4750) <= not((layer5_outputs(102)) or (layer5_outputs(3856)));
    layer6_outputs(4751) <= not(layer5_outputs(1203));
    layer6_outputs(4752) <= not(layer5_outputs(3998));
    layer6_outputs(4753) <= not((layer5_outputs(488)) and (layer5_outputs(3609)));
    layer6_outputs(4754) <= (layer5_outputs(4748)) xor (layer5_outputs(4401));
    layer6_outputs(4755) <= not(layer5_outputs(1280));
    layer6_outputs(4756) <= (layer5_outputs(949)) and (layer5_outputs(5038));
    layer6_outputs(4757) <= not(layer5_outputs(30));
    layer6_outputs(4758) <= '0';
    layer6_outputs(4759) <= layer5_outputs(526);
    layer6_outputs(4760) <= (layer5_outputs(1240)) and (layer5_outputs(1216));
    layer6_outputs(4761) <= (layer5_outputs(4367)) or (layer5_outputs(2596));
    layer6_outputs(4762) <= not((layer5_outputs(2170)) and (layer5_outputs(2505)));
    layer6_outputs(4763) <= (layer5_outputs(1388)) or (layer5_outputs(4088));
    layer6_outputs(4764) <= not(layer5_outputs(425));
    layer6_outputs(4765) <= not((layer5_outputs(2437)) xor (layer5_outputs(2514)));
    layer6_outputs(4766) <= layer5_outputs(3275);
    layer6_outputs(4767) <= not(layer5_outputs(164));
    layer6_outputs(4768) <= '0';
    layer6_outputs(4769) <= not((layer5_outputs(4712)) and (layer5_outputs(1853)));
    layer6_outputs(4770) <= not(layer5_outputs(1550));
    layer6_outputs(4771) <= layer5_outputs(1304);
    layer6_outputs(4772) <= not((layer5_outputs(3706)) xor (layer5_outputs(3151)));
    layer6_outputs(4773) <= not(layer5_outputs(4919));
    layer6_outputs(4774) <= not(layer5_outputs(1548)) or (layer5_outputs(938));
    layer6_outputs(4775) <= (layer5_outputs(2292)) and not (layer5_outputs(2712));
    layer6_outputs(4776) <= (layer5_outputs(3425)) and not (layer5_outputs(644));
    layer6_outputs(4777) <= (layer5_outputs(1968)) or (layer5_outputs(4973));
    layer6_outputs(4778) <= (layer5_outputs(889)) or (layer5_outputs(4515));
    layer6_outputs(4779) <= (layer5_outputs(2524)) and not (layer5_outputs(3554));
    layer6_outputs(4780) <= not(layer5_outputs(3825));
    layer6_outputs(4781) <= not((layer5_outputs(624)) xor (layer5_outputs(3525)));
    layer6_outputs(4782) <= not(layer5_outputs(4052));
    layer6_outputs(4783) <= not((layer5_outputs(3389)) and (layer5_outputs(3748)));
    layer6_outputs(4784) <= not(layer5_outputs(4243));
    layer6_outputs(4785) <= layer5_outputs(4019);
    layer6_outputs(4786) <= (layer5_outputs(734)) xor (layer5_outputs(4398));
    layer6_outputs(4787) <= not(layer5_outputs(3563));
    layer6_outputs(4788) <= not(layer5_outputs(2312));
    layer6_outputs(4789) <= not((layer5_outputs(3222)) or (layer5_outputs(4375)));
    layer6_outputs(4790) <= '1';
    layer6_outputs(4791) <= '1';
    layer6_outputs(4792) <= layer5_outputs(2731);
    layer6_outputs(4793) <= not(layer5_outputs(3376));
    layer6_outputs(4794) <= layer5_outputs(277);
    layer6_outputs(4795) <= not(layer5_outputs(1648)) or (layer5_outputs(4479));
    layer6_outputs(4796) <= layer5_outputs(1069);
    layer6_outputs(4797) <= not((layer5_outputs(915)) and (layer5_outputs(2473)));
    layer6_outputs(4798) <= not((layer5_outputs(205)) and (layer5_outputs(626)));
    layer6_outputs(4799) <= not(layer5_outputs(1173));
    layer6_outputs(4800) <= not(layer5_outputs(571));
    layer6_outputs(4801) <= layer5_outputs(3883);
    layer6_outputs(4802) <= layer5_outputs(4543);
    layer6_outputs(4803) <= layer5_outputs(2945);
    layer6_outputs(4804) <= not(layer5_outputs(233));
    layer6_outputs(4805) <= '1';
    layer6_outputs(4806) <= layer5_outputs(4189);
    layer6_outputs(4807) <= not((layer5_outputs(3371)) xor (layer5_outputs(1625)));
    layer6_outputs(4808) <= not((layer5_outputs(4227)) or (layer5_outputs(4370)));
    layer6_outputs(4809) <= not((layer5_outputs(2382)) or (layer5_outputs(3167)));
    layer6_outputs(4810) <= (layer5_outputs(486)) and not (layer5_outputs(4550));
    layer6_outputs(4811) <= not(layer5_outputs(1788));
    layer6_outputs(4812) <= not((layer5_outputs(2310)) or (layer5_outputs(1047)));
    layer6_outputs(4813) <= (layer5_outputs(379)) xor (layer5_outputs(166));
    layer6_outputs(4814) <= not(layer5_outputs(195)) or (layer5_outputs(2580));
    layer6_outputs(4815) <= not((layer5_outputs(1585)) xor (layer5_outputs(3648)));
    layer6_outputs(4816) <= not(layer5_outputs(1248));
    layer6_outputs(4817) <= not((layer5_outputs(2480)) or (layer5_outputs(3504)));
    layer6_outputs(4818) <= layer5_outputs(5098);
    layer6_outputs(4819) <= layer5_outputs(3468);
    layer6_outputs(4820) <= layer5_outputs(344);
    layer6_outputs(4821) <= not((layer5_outputs(2149)) xor (layer5_outputs(4939)));
    layer6_outputs(4822) <= not(layer5_outputs(3162));
    layer6_outputs(4823) <= (layer5_outputs(1863)) and not (layer5_outputs(976));
    layer6_outputs(4824) <= not((layer5_outputs(4468)) and (layer5_outputs(345)));
    layer6_outputs(4825) <= not((layer5_outputs(1317)) xor (layer5_outputs(3150)));
    layer6_outputs(4826) <= (layer5_outputs(3362)) and not (layer5_outputs(1786));
    layer6_outputs(4827) <= layer5_outputs(1743);
    layer6_outputs(4828) <= (layer5_outputs(5075)) xor (layer5_outputs(1095));
    layer6_outputs(4829) <= not((layer5_outputs(156)) and (layer5_outputs(2364)));
    layer6_outputs(4830) <= not(layer5_outputs(4832));
    layer6_outputs(4831) <= not((layer5_outputs(914)) xor (layer5_outputs(4726)));
    layer6_outputs(4832) <= not((layer5_outputs(5083)) and (layer5_outputs(37)));
    layer6_outputs(4833) <= not(layer5_outputs(1474));
    layer6_outputs(4834) <= layer5_outputs(4185);
    layer6_outputs(4835) <= not(layer5_outputs(4841));
    layer6_outputs(4836) <= not(layer5_outputs(2954)) or (layer5_outputs(3120));
    layer6_outputs(4837) <= (layer5_outputs(3492)) or (layer5_outputs(314));
    layer6_outputs(4838) <= layer5_outputs(1);
    layer6_outputs(4839) <= not(layer5_outputs(3293)) or (layer5_outputs(3107));
    layer6_outputs(4840) <= (layer5_outputs(565)) and (layer5_outputs(4386));
    layer6_outputs(4841) <= layer5_outputs(2897);
    layer6_outputs(4842) <= not(layer5_outputs(723));
    layer6_outputs(4843) <= layer5_outputs(2024);
    layer6_outputs(4844) <= not(layer5_outputs(3994));
    layer6_outputs(4845) <= layer5_outputs(2448);
    layer6_outputs(4846) <= (layer5_outputs(2404)) or (layer5_outputs(4472));
    layer6_outputs(4847) <= not((layer5_outputs(3217)) xor (layer5_outputs(3529)));
    layer6_outputs(4848) <= not(layer5_outputs(3526)) or (layer5_outputs(1022));
    layer6_outputs(4849) <= layer5_outputs(3321);
    layer6_outputs(4850) <= (layer5_outputs(4510)) xor (layer5_outputs(2023));
    layer6_outputs(4851) <= (layer5_outputs(3385)) and not (layer5_outputs(332));
    layer6_outputs(4852) <= layer5_outputs(2518);
    layer6_outputs(4853) <= not(layer5_outputs(418));
    layer6_outputs(4854) <= not(layer5_outputs(4452)) or (layer5_outputs(665));
    layer6_outputs(4855) <= not((layer5_outputs(3282)) or (layer5_outputs(1684)));
    layer6_outputs(4856) <= not((layer5_outputs(4842)) and (layer5_outputs(4031)));
    layer6_outputs(4857) <= not((layer5_outputs(3925)) or (layer5_outputs(4751)));
    layer6_outputs(4858) <= (layer5_outputs(4782)) or (layer5_outputs(1787));
    layer6_outputs(4859) <= layer5_outputs(2269);
    layer6_outputs(4860) <= not(layer5_outputs(1116));
    layer6_outputs(4861) <= layer5_outputs(4060);
    layer6_outputs(4862) <= not((layer5_outputs(588)) xor (layer5_outputs(2783)));
    layer6_outputs(4863) <= not(layer5_outputs(2900));
    layer6_outputs(4864) <= (layer5_outputs(4544)) xor (layer5_outputs(2217));
    layer6_outputs(4865) <= (layer5_outputs(514)) or (layer5_outputs(634));
    layer6_outputs(4866) <= layer5_outputs(848);
    layer6_outputs(4867) <= not((layer5_outputs(1518)) xor (layer5_outputs(18)));
    layer6_outputs(4868) <= (layer5_outputs(25)) xor (layer5_outputs(3691));
    layer6_outputs(4869) <= layer5_outputs(650);
    layer6_outputs(4870) <= not((layer5_outputs(2645)) xor (layer5_outputs(5063)));
    layer6_outputs(4871) <= (layer5_outputs(1574)) and not (layer5_outputs(903));
    layer6_outputs(4872) <= layer5_outputs(4315);
    layer6_outputs(4873) <= (layer5_outputs(294)) xor (layer5_outputs(2400));
    layer6_outputs(4874) <= (layer5_outputs(4294)) xor (layer5_outputs(3643));
    layer6_outputs(4875) <= layer5_outputs(2373);
    layer6_outputs(4876) <= layer5_outputs(3754);
    layer6_outputs(4877) <= not(layer5_outputs(2793));
    layer6_outputs(4878) <= not(layer5_outputs(3929)) or (layer5_outputs(4501));
    layer6_outputs(4879) <= (layer5_outputs(2714)) and (layer5_outputs(116));
    layer6_outputs(4880) <= (layer5_outputs(1654)) and not (layer5_outputs(3046));
    layer6_outputs(4881) <= not(layer5_outputs(636)) or (layer5_outputs(1570));
    layer6_outputs(4882) <= '1';
    layer6_outputs(4883) <= not(layer5_outputs(4138));
    layer6_outputs(4884) <= not(layer5_outputs(2827)) or (layer5_outputs(3413));
    layer6_outputs(4885) <= (layer5_outputs(388)) and (layer5_outputs(3184));
    layer6_outputs(4886) <= (layer5_outputs(4324)) xor (layer5_outputs(4567));
    layer6_outputs(4887) <= not(layer5_outputs(428)) or (layer5_outputs(1578));
    layer6_outputs(4888) <= (layer5_outputs(898)) and not (layer5_outputs(4146));
    layer6_outputs(4889) <= (layer5_outputs(486)) and (layer5_outputs(3207));
    layer6_outputs(4890) <= (layer5_outputs(1816)) xor (layer5_outputs(764));
    layer6_outputs(4891) <= layer5_outputs(1983);
    layer6_outputs(4892) <= '1';
    layer6_outputs(4893) <= (layer5_outputs(4385)) and not (layer5_outputs(3734));
    layer6_outputs(4894) <= layer5_outputs(4942);
    layer6_outputs(4895) <= layer5_outputs(2588);
    layer6_outputs(4896) <= not((layer5_outputs(2152)) or (layer5_outputs(1962)));
    layer6_outputs(4897) <= not(layer5_outputs(2968));
    layer6_outputs(4898) <= not(layer5_outputs(165));
    layer6_outputs(4899) <= (layer5_outputs(4299)) xor (layer5_outputs(3711));
    layer6_outputs(4900) <= not(layer5_outputs(4236));
    layer6_outputs(4901) <= layer5_outputs(1518);
    layer6_outputs(4902) <= layer5_outputs(253);
    layer6_outputs(4903) <= layer5_outputs(833);
    layer6_outputs(4904) <= not(layer5_outputs(2151)) or (layer5_outputs(3560));
    layer6_outputs(4905) <= not(layer5_outputs(2985));
    layer6_outputs(4906) <= layer5_outputs(4411);
    layer6_outputs(4907) <= not(layer5_outputs(2808)) or (layer5_outputs(4855));
    layer6_outputs(4908) <= (layer5_outputs(7)) and not (layer5_outputs(1540));
    layer6_outputs(4909) <= not(layer5_outputs(2372));
    layer6_outputs(4910) <= layer5_outputs(1559);
    layer6_outputs(4911) <= (layer5_outputs(2905)) and (layer5_outputs(1083));
    layer6_outputs(4912) <= layer5_outputs(3556);
    layer6_outputs(4913) <= layer5_outputs(3834);
    layer6_outputs(4914) <= (layer5_outputs(657)) and (layer5_outputs(620));
    layer6_outputs(4915) <= (layer5_outputs(3308)) or (layer5_outputs(4772));
    layer6_outputs(4916) <= layer5_outputs(2649);
    layer6_outputs(4917) <= not((layer5_outputs(2877)) and (layer5_outputs(4301)));
    layer6_outputs(4918) <= '0';
    layer6_outputs(4919) <= not((layer5_outputs(228)) and (layer5_outputs(712)));
    layer6_outputs(4920) <= (layer5_outputs(370)) and not (layer5_outputs(1460));
    layer6_outputs(4921) <= not(layer5_outputs(3968));
    layer6_outputs(4922) <= not(layer5_outputs(2916)) or (layer5_outputs(3661));
    layer6_outputs(4923) <= (layer5_outputs(1677)) and not (layer5_outputs(1799));
    layer6_outputs(4924) <= not((layer5_outputs(645)) and (layer5_outputs(890)));
    layer6_outputs(4925) <= layer5_outputs(4499);
    layer6_outputs(4926) <= not(layer5_outputs(4183));
    layer6_outputs(4927) <= not(layer5_outputs(1857)) or (layer5_outputs(1297));
    layer6_outputs(4928) <= '1';
    layer6_outputs(4929) <= layer5_outputs(2953);
    layer6_outputs(4930) <= not(layer5_outputs(1964)) or (layer5_outputs(4854));
    layer6_outputs(4931) <= not(layer5_outputs(330));
    layer6_outputs(4932) <= not(layer5_outputs(4834));
    layer6_outputs(4933) <= not(layer5_outputs(1221));
    layer6_outputs(4934) <= layer5_outputs(2198);
    layer6_outputs(4935) <= not(layer5_outputs(3109));
    layer6_outputs(4936) <= (layer5_outputs(177)) or (layer5_outputs(3147));
    layer6_outputs(4937) <= layer5_outputs(4315);
    layer6_outputs(4938) <= not(layer5_outputs(3540));
    layer6_outputs(4939) <= (layer5_outputs(1734)) xor (layer5_outputs(1307));
    layer6_outputs(4940) <= '0';
    layer6_outputs(4941) <= not((layer5_outputs(1587)) or (layer5_outputs(174)));
    layer6_outputs(4942) <= layer5_outputs(3227);
    layer6_outputs(4943) <= not((layer5_outputs(2711)) or (layer5_outputs(3284)));
    layer6_outputs(4944) <= not(layer5_outputs(3429)) or (layer5_outputs(3859));
    layer6_outputs(4945) <= (layer5_outputs(1762)) and not (layer5_outputs(3756));
    layer6_outputs(4946) <= not((layer5_outputs(368)) and (layer5_outputs(1641)));
    layer6_outputs(4947) <= (layer5_outputs(1235)) and (layer5_outputs(3262));
    layer6_outputs(4948) <= (layer5_outputs(3435)) or (layer5_outputs(4410));
    layer6_outputs(4949) <= not(layer5_outputs(4260));
    layer6_outputs(4950) <= (layer5_outputs(2877)) and not (layer5_outputs(449));
    layer6_outputs(4951) <= not((layer5_outputs(4162)) and (layer5_outputs(4291)));
    layer6_outputs(4952) <= layer5_outputs(1211);
    layer6_outputs(4953) <= layer5_outputs(3692);
    layer6_outputs(4954) <= layer5_outputs(248);
    layer6_outputs(4955) <= (layer5_outputs(2082)) or (layer5_outputs(1922));
    layer6_outputs(4956) <= not(layer5_outputs(780)) or (layer5_outputs(1723));
    layer6_outputs(4957) <= (layer5_outputs(40)) or (layer5_outputs(4903));
    layer6_outputs(4958) <= layer5_outputs(2300);
    layer6_outputs(4959) <= (layer5_outputs(962)) and not (layer5_outputs(4367));
    layer6_outputs(4960) <= layer5_outputs(1861);
    layer6_outputs(4961) <= (layer5_outputs(3491)) and not (layer5_outputs(1727));
    layer6_outputs(4962) <= (layer5_outputs(3175)) and not (layer5_outputs(4171));
    layer6_outputs(4963) <= not(layer5_outputs(3154));
    layer6_outputs(4964) <= (layer5_outputs(4565)) and not (layer5_outputs(1451));
    layer6_outputs(4965) <= not((layer5_outputs(2804)) and (layer5_outputs(2656)));
    layer6_outputs(4966) <= (layer5_outputs(1683)) and not (layer5_outputs(4295));
    layer6_outputs(4967) <= not(layer5_outputs(1132));
    layer6_outputs(4968) <= layer5_outputs(47);
    layer6_outputs(4969) <= layer5_outputs(1211);
    layer6_outputs(4970) <= not((layer5_outputs(2218)) xor (layer5_outputs(4319)));
    layer6_outputs(4971) <= not(layer5_outputs(1329));
    layer6_outputs(4972) <= not((layer5_outputs(1073)) or (layer5_outputs(2659)));
    layer6_outputs(4973) <= '1';
    layer6_outputs(4974) <= (layer5_outputs(4518)) xor (layer5_outputs(2549));
    layer6_outputs(4975) <= '1';
    layer6_outputs(4976) <= not(layer5_outputs(4187)) or (layer5_outputs(5037));
    layer6_outputs(4977) <= not((layer5_outputs(683)) xor (layer5_outputs(3832)));
    layer6_outputs(4978) <= not(layer5_outputs(496));
    layer6_outputs(4979) <= layer5_outputs(4446);
    layer6_outputs(4980) <= (layer5_outputs(3495)) and (layer5_outputs(4799));
    layer6_outputs(4981) <= layer5_outputs(2450);
    layer6_outputs(4982) <= (layer5_outputs(2922)) and not (layer5_outputs(3794));
    layer6_outputs(4983) <= not(layer5_outputs(1151)) or (layer5_outputs(4502));
    layer6_outputs(4984) <= not((layer5_outputs(412)) and (layer5_outputs(2214)));
    layer6_outputs(4985) <= not((layer5_outputs(4681)) and (layer5_outputs(4176)));
    layer6_outputs(4986) <= (layer5_outputs(1117)) and (layer5_outputs(4177));
    layer6_outputs(4987) <= (layer5_outputs(3694)) xor (layer5_outputs(1111));
    layer6_outputs(4988) <= (layer5_outputs(3782)) and not (layer5_outputs(4592));
    layer6_outputs(4989) <= not(layer5_outputs(4016));
    layer6_outputs(4990) <= layer5_outputs(4819);
    layer6_outputs(4991) <= '0';
    layer6_outputs(4992) <= not(layer5_outputs(98)) or (layer5_outputs(1511));
    layer6_outputs(4993) <= (layer5_outputs(4673)) and not (layer5_outputs(120));
    layer6_outputs(4994) <= (layer5_outputs(656)) and not (layer5_outputs(2828));
    layer6_outputs(4995) <= layer5_outputs(5061);
    layer6_outputs(4996) <= layer5_outputs(3540);
    layer6_outputs(4997) <= layer5_outputs(1120);
    layer6_outputs(4998) <= (layer5_outputs(3339)) and not (layer5_outputs(1065));
    layer6_outputs(4999) <= not(layer5_outputs(1364));
    layer6_outputs(5000) <= layer5_outputs(3025);
    layer6_outputs(5001) <= not(layer5_outputs(777)) or (layer5_outputs(3836));
    layer6_outputs(5002) <= (layer5_outputs(763)) and (layer5_outputs(788));
    layer6_outputs(5003) <= '1';
    layer6_outputs(5004) <= (layer5_outputs(2612)) or (layer5_outputs(2039));
    layer6_outputs(5005) <= not(layer5_outputs(859));
    layer6_outputs(5006) <= layer5_outputs(3868);
    layer6_outputs(5007) <= layer5_outputs(4021);
    layer6_outputs(5008) <= layer5_outputs(905);
    layer6_outputs(5009) <= not((layer5_outputs(1947)) or (layer5_outputs(2147)));
    layer6_outputs(5010) <= not(layer5_outputs(1835));
    layer6_outputs(5011) <= (layer5_outputs(4233)) and (layer5_outputs(1490));
    layer6_outputs(5012) <= (layer5_outputs(497)) and not (layer5_outputs(1849));
    layer6_outputs(5013) <= not(layer5_outputs(3612)) or (layer5_outputs(2806));
    layer6_outputs(5014) <= (layer5_outputs(4376)) and not (layer5_outputs(2204));
    layer6_outputs(5015) <= not(layer5_outputs(365)) or (layer5_outputs(2251));
    layer6_outputs(5016) <= not(layer5_outputs(3266));
    layer6_outputs(5017) <= (layer5_outputs(1113)) or (layer5_outputs(2401));
    layer6_outputs(5018) <= not(layer5_outputs(187)) or (layer5_outputs(3567));
    layer6_outputs(5019) <= layer5_outputs(4878);
    layer6_outputs(5020) <= not((layer5_outputs(3187)) xor (layer5_outputs(1619)));
    layer6_outputs(5021) <= not(layer5_outputs(2)) or (layer5_outputs(1026));
    layer6_outputs(5022) <= not(layer5_outputs(1081));
    layer6_outputs(5023) <= not(layer5_outputs(4060)) or (layer5_outputs(2191));
    layer6_outputs(5024) <= (layer5_outputs(3536)) or (layer5_outputs(573));
    layer6_outputs(5025) <= layer5_outputs(4113);
    layer6_outputs(5026) <= not(layer5_outputs(4034));
    layer6_outputs(5027) <= not((layer5_outputs(4409)) or (layer5_outputs(3096)));
    layer6_outputs(5028) <= not(layer5_outputs(1340));
    layer6_outputs(5029) <= (layer5_outputs(1677)) or (layer5_outputs(2562));
    layer6_outputs(5030) <= layer5_outputs(3874);
    layer6_outputs(5031) <= (layer5_outputs(1227)) or (layer5_outputs(4172));
    layer6_outputs(5032) <= (layer5_outputs(4793)) or (layer5_outputs(218));
    layer6_outputs(5033) <= layer5_outputs(3242);
    layer6_outputs(5034) <= (layer5_outputs(1831)) and (layer5_outputs(4204));
    layer6_outputs(5035) <= (layer5_outputs(4257)) and not (layer5_outputs(4264));
    layer6_outputs(5036) <= not(layer5_outputs(4663));
    layer6_outputs(5037) <= not(layer5_outputs(2018));
    layer6_outputs(5038) <= (layer5_outputs(2378)) and (layer5_outputs(549));
    layer6_outputs(5039) <= layer5_outputs(627);
    layer6_outputs(5040) <= not((layer5_outputs(4928)) or (layer5_outputs(4829)));
    layer6_outputs(5041) <= '0';
    layer6_outputs(5042) <= not((layer5_outputs(2065)) and (layer5_outputs(2504)));
    layer6_outputs(5043) <= (layer5_outputs(2168)) xor (layer5_outputs(3201));
    layer6_outputs(5044) <= layer5_outputs(2409);
    layer6_outputs(5045) <= (layer5_outputs(1506)) xor (layer5_outputs(2820));
    layer6_outputs(5046) <= (layer5_outputs(1474)) or (layer5_outputs(4013));
    layer6_outputs(5047) <= (layer5_outputs(3866)) and not (layer5_outputs(155));
    layer6_outputs(5048) <= not(layer5_outputs(3275)) or (layer5_outputs(3117));
    layer6_outputs(5049) <= not(layer5_outputs(1454)) or (layer5_outputs(2931));
    layer6_outputs(5050) <= not((layer5_outputs(3709)) xor (layer5_outputs(4850)));
    layer6_outputs(5051) <= not(layer5_outputs(961));
    layer6_outputs(5052) <= not((layer5_outputs(67)) xor (layer5_outputs(39)));
    layer6_outputs(5053) <= layer5_outputs(2489);
    layer6_outputs(5054) <= (layer5_outputs(1086)) and (layer5_outputs(2260));
    layer6_outputs(5055) <= not(layer5_outputs(4293));
    layer6_outputs(5056) <= (layer5_outputs(2745)) and not (layer5_outputs(2777));
    layer6_outputs(5057) <= layer5_outputs(998);
    layer6_outputs(5058) <= layer5_outputs(758);
    layer6_outputs(5059) <= (layer5_outputs(2129)) and (layer5_outputs(3657));
    layer6_outputs(5060) <= not(layer5_outputs(2825));
    layer6_outputs(5061) <= not(layer5_outputs(3204)) or (layer5_outputs(3801));
    layer6_outputs(5062) <= layer5_outputs(3852);
    layer6_outputs(5063) <= (layer5_outputs(4677)) xor (layer5_outputs(1094));
    layer6_outputs(5064) <= not(layer5_outputs(3991)) or (layer5_outputs(2530));
    layer6_outputs(5065) <= (layer5_outputs(586)) and (layer5_outputs(2977));
    layer6_outputs(5066) <= not(layer5_outputs(1139));
    layer6_outputs(5067) <= not(layer5_outputs(2100));
    layer6_outputs(5068) <= not(layer5_outputs(355));
    layer6_outputs(5069) <= (layer5_outputs(5109)) or (layer5_outputs(3944));
    layer6_outputs(5070) <= (layer5_outputs(1866)) and not (layer5_outputs(4467));
    layer6_outputs(5071) <= not((layer5_outputs(3448)) or (layer5_outputs(234)));
    layer6_outputs(5072) <= '0';
    layer6_outputs(5073) <= (layer5_outputs(2063)) and not (layer5_outputs(5017));
    layer6_outputs(5074) <= layer5_outputs(4156);
    layer6_outputs(5075) <= not((layer5_outputs(4992)) or (layer5_outputs(4741)));
    layer6_outputs(5076) <= not((layer5_outputs(454)) or (layer5_outputs(2635)));
    layer6_outputs(5077) <= '0';
    layer6_outputs(5078) <= '0';
    layer6_outputs(5079) <= layer5_outputs(722);
    layer6_outputs(5080) <= layer5_outputs(737);
    layer6_outputs(5081) <= (layer5_outputs(4454)) xor (layer5_outputs(3612));
    layer6_outputs(5082) <= (layer5_outputs(4756)) or (layer5_outputs(1172));
    layer6_outputs(5083) <= layer5_outputs(5043);
    layer6_outputs(5084) <= not((layer5_outputs(4721)) or (layer5_outputs(1453)));
    layer6_outputs(5085) <= layer5_outputs(1984);
    layer6_outputs(5086) <= not(layer5_outputs(430));
    layer6_outputs(5087) <= (layer5_outputs(1652)) and not (layer5_outputs(1138));
    layer6_outputs(5088) <= not(layer5_outputs(3602));
    layer6_outputs(5089) <= (layer5_outputs(1243)) and not (layer5_outputs(2624));
    layer6_outputs(5090) <= not(layer5_outputs(1464));
    layer6_outputs(5091) <= not(layer5_outputs(2215)) or (layer5_outputs(1301));
    layer6_outputs(5092) <= not(layer5_outputs(2833)) or (layer5_outputs(911));
    layer6_outputs(5093) <= not(layer5_outputs(1471));
    layer6_outputs(5094) <= (layer5_outputs(4200)) and not (layer5_outputs(4793));
    layer6_outputs(5095) <= layer5_outputs(4379);
    layer6_outputs(5096) <= not((layer5_outputs(1246)) or (layer5_outputs(3626)));
    layer6_outputs(5097) <= (layer5_outputs(1253)) xor (layer5_outputs(2360));
    layer6_outputs(5098) <= not(layer5_outputs(2810));
    layer6_outputs(5099) <= not(layer5_outputs(2487));
    layer6_outputs(5100) <= not(layer5_outputs(5028));
    layer6_outputs(5101) <= (layer5_outputs(1907)) and not (layer5_outputs(926));
    layer6_outputs(5102) <= not(layer5_outputs(3279));
    layer6_outputs(5103) <= not(layer5_outputs(1933));
    layer6_outputs(5104) <= not((layer5_outputs(4857)) and (layer5_outputs(882)));
    layer6_outputs(5105) <= not(layer5_outputs(257)) or (layer5_outputs(405));
    layer6_outputs(5106) <= not(layer5_outputs(1935));
    layer6_outputs(5107) <= (layer5_outputs(3983)) and not (layer5_outputs(1995));
    layer6_outputs(5108) <= layer5_outputs(2614);
    layer6_outputs(5109) <= not(layer5_outputs(2718)) or (layer5_outputs(4664));
    layer6_outputs(5110) <= not(layer5_outputs(320));
    layer6_outputs(5111) <= not(layer5_outputs(3242));
    layer6_outputs(5112) <= not(layer5_outputs(2202));
    layer6_outputs(5113) <= layer5_outputs(2028);
    layer6_outputs(5114) <= not(layer5_outputs(4450));
    layer6_outputs(5115) <= (layer5_outputs(3030)) and not (layer5_outputs(5085));
    layer6_outputs(5116) <= not((layer5_outputs(179)) or (layer5_outputs(5043)));
    layer6_outputs(5117) <= not(layer5_outputs(442)) or (layer5_outputs(1614));
    layer6_outputs(5118) <= (layer5_outputs(3095)) or (layer5_outputs(1575));
    layer6_outputs(5119) <= layer5_outputs(4887);
    layer7_outputs(0) <= not(layer6_outputs(391));
    layer7_outputs(1) <= not((layer6_outputs(4139)) xor (layer6_outputs(2622)));
    layer7_outputs(2) <= (layer6_outputs(1740)) xor (layer6_outputs(1085));
    layer7_outputs(3) <= layer6_outputs(2574);
    layer7_outputs(4) <= (layer6_outputs(3657)) xor (layer6_outputs(2348));
    layer7_outputs(5) <= layer6_outputs(3410);
    layer7_outputs(6) <= (layer6_outputs(4894)) xor (layer6_outputs(2367));
    layer7_outputs(7) <= (layer6_outputs(4966)) and (layer6_outputs(3647));
    layer7_outputs(8) <= layer6_outputs(1854);
    layer7_outputs(9) <= layer6_outputs(1719);
    layer7_outputs(10) <= (layer6_outputs(725)) xor (layer6_outputs(4398));
    layer7_outputs(11) <= not(layer6_outputs(295));
    layer7_outputs(12) <= not(layer6_outputs(2754));
    layer7_outputs(13) <= layer6_outputs(3104);
    layer7_outputs(14) <= '1';
    layer7_outputs(15) <= layer6_outputs(5);
    layer7_outputs(16) <= not(layer6_outputs(1519));
    layer7_outputs(17) <= not(layer6_outputs(2892));
    layer7_outputs(18) <= not(layer6_outputs(920));
    layer7_outputs(19) <= not(layer6_outputs(4628)) or (layer6_outputs(2536));
    layer7_outputs(20) <= not(layer6_outputs(4697)) or (layer6_outputs(2062));
    layer7_outputs(21) <= not(layer6_outputs(1433));
    layer7_outputs(22) <= (layer6_outputs(1674)) and not (layer6_outputs(3562));
    layer7_outputs(23) <= not(layer6_outputs(2012));
    layer7_outputs(24) <= not(layer6_outputs(1002)) or (layer6_outputs(2031));
    layer7_outputs(25) <= not(layer6_outputs(2326)) or (layer6_outputs(4783));
    layer7_outputs(26) <= '1';
    layer7_outputs(27) <= not((layer6_outputs(3384)) xor (layer6_outputs(4874)));
    layer7_outputs(28) <= (layer6_outputs(3379)) and not (layer6_outputs(491));
    layer7_outputs(29) <= not(layer6_outputs(4372));
    layer7_outputs(30) <= (layer6_outputs(455)) and not (layer6_outputs(969));
    layer7_outputs(31) <= (layer6_outputs(2995)) and not (layer6_outputs(2406));
    layer7_outputs(32) <= not(layer6_outputs(349));
    layer7_outputs(33) <= not(layer6_outputs(3103));
    layer7_outputs(34) <= not((layer6_outputs(4918)) and (layer6_outputs(1855)));
    layer7_outputs(35) <= not(layer6_outputs(4650));
    layer7_outputs(36) <= not(layer6_outputs(373));
    layer7_outputs(37) <= not(layer6_outputs(4535));
    layer7_outputs(38) <= layer6_outputs(1137);
    layer7_outputs(39) <= not(layer6_outputs(1517));
    layer7_outputs(40) <= not(layer6_outputs(4132));
    layer7_outputs(41) <= (layer6_outputs(4559)) or (layer6_outputs(519));
    layer7_outputs(42) <= not(layer6_outputs(5014));
    layer7_outputs(43) <= not(layer6_outputs(3864));
    layer7_outputs(44) <= (layer6_outputs(251)) xor (layer6_outputs(3168));
    layer7_outputs(45) <= not((layer6_outputs(4789)) and (layer6_outputs(4910)));
    layer7_outputs(46) <= not((layer6_outputs(2640)) and (layer6_outputs(784)));
    layer7_outputs(47) <= layer6_outputs(2214);
    layer7_outputs(48) <= layer6_outputs(2097);
    layer7_outputs(49) <= not(layer6_outputs(3457));
    layer7_outputs(50) <= layer6_outputs(4931);
    layer7_outputs(51) <= not(layer6_outputs(2919));
    layer7_outputs(52) <= not(layer6_outputs(2278));
    layer7_outputs(53) <= not((layer6_outputs(1512)) or (layer6_outputs(799)));
    layer7_outputs(54) <= not((layer6_outputs(1869)) and (layer6_outputs(3337)));
    layer7_outputs(55) <= (layer6_outputs(308)) or (layer6_outputs(903));
    layer7_outputs(56) <= (layer6_outputs(4834)) and not (layer6_outputs(2511));
    layer7_outputs(57) <= not(layer6_outputs(3567));
    layer7_outputs(58) <= not(layer6_outputs(4900));
    layer7_outputs(59) <= not((layer6_outputs(3184)) or (layer6_outputs(3358)));
    layer7_outputs(60) <= not((layer6_outputs(4491)) or (layer6_outputs(1884)));
    layer7_outputs(61) <= (layer6_outputs(3739)) xor (layer6_outputs(1660));
    layer7_outputs(62) <= layer6_outputs(2926);
    layer7_outputs(63) <= not((layer6_outputs(1248)) xor (layer6_outputs(2698)));
    layer7_outputs(64) <= not(layer6_outputs(1825));
    layer7_outputs(65) <= layer6_outputs(898);
    layer7_outputs(66) <= layer6_outputs(2731);
    layer7_outputs(67) <= not(layer6_outputs(2126)) or (layer6_outputs(3496));
    layer7_outputs(68) <= not(layer6_outputs(3893)) or (layer6_outputs(1621));
    layer7_outputs(69) <= not((layer6_outputs(1604)) or (layer6_outputs(2232)));
    layer7_outputs(70) <= (layer6_outputs(2949)) xor (layer6_outputs(1826));
    layer7_outputs(71) <= (layer6_outputs(4253)) or (layer6_outputs(3855));
    layer7_outputs(72) <= layer6_outputs(4887);
    layer7_outputs(73) <= not(layer6_outputs(1223)) or (layer6_outputs(5059));
    layer7_outputs(74) <= (layer6_outputs(710)) xor (layer6_outputs(1254));
    layer7_outputs(75) <= not((layer6_outputs(401)) and (layer6_outputs(1702)));
    layer7_outputs(76) <= not(layer6_outputs(4838)) or (layer6_outputs(3495));
    layer7_outputs(77) <= not((layer6_outputs(1141)) or (layer6_outputs(1071)));
    layer7_outputs(78) <= not(layer6_outputs(5085));
    layer7_outputs(79) <= not(layer6_outputs(4039));
    layer7_outputs(80) <= not(layer6_outputs(4835)) or (layer6_outputs(1968));
    layer7_outputs(81) <= not(layer6_outputs(3510));
    layer7_outputs(82) <= not(layer6_outputs(1970));
    layer7_outputs(83) <= not(layer6_outputs(350));
    layer7_outputs(84) <= layer6_outputs(3011);
    layer7_outputs(85) <= not(layer6_outputs(1160));
    layer7_outputs(86) <= layer6_outputs(2656);
    layer7_outputs(87) <= not(layer6_outputs(1731));
    layer7_outputs(88) <= not((layer6_outputs(3995)) xor (layer6_outputs(4219)));
    layer7_outputs(89) <= not((layer6_outputs(171)) xor (layer6_outputs(1622)));
    layer7_outputs(90) <= layer6_outputs(625);
    layer7_outputs(91) <= not(layer6_outputs(1194));
    layer7_outputs(92) <= not(layer6_outputs(4807));
    layer7_outputs(93) <= (layer6_outputs(1065)) xor (layer6_outputs(1757));
    layer7_outputs(94) <= layer6_outputs(1714);
    layer7_outputs(95) <= '1';
    layer7_outputs(96) <= not((layer6_outputs(4864)) and (layer6_outputs(358)));
    layer7_outputs(97) <= not(layer6_outputs(3403));
    layer7_outputs(98) <= not(layer6_outputs(3151)) or (layer6_outputs(1898));
    layer7_outputs(99) <= layer6_outputs(2788);
    layer7_outputs(100) <= (layer6_outputs(2387)) and not (layer6_outputs(887));
    layer7_outputs(101) <= layer6_outputs(80);
    layer7_outputs(102) <= not(layer6_outputs(5080));
    layer7_outputs(103) <= not(layer6_outputs(196));
    layer7_outputs(104) <= not(layer6_outputs(4357));
    layer7_outputs(105) <= not(layer6_outputs(2732));
    layer7_outputs(106) <= not(layer6_outputs(3896));
    layer7_outputs(107) <= not(layer6_outputs(3129)) or (layer6_outputs(2200));
    layer7_outputs(108) <= (layer6_outputs(2766)) and not (layer6_outputs(2604));
    layer7_outputs(109) <= not((layer6_outputs(1889)) and (layer6_outputs(4744)));
    layer7_outputs(110) <= not((layer6_outputs(286)) and (layer6_outputs(173)));
    layer7_outputs(111) <= not(layer6_outputs(4933)) or (layer6_outputs(4714));
    layer7_outputs(112) <= layer6_outputs(2404);
    layer7_outputs(113) <= not((layer6_outputs(3463)) xor (layer6_outputs(970)));
    layer7_outputs(114) <= not((layer6_outputs(3985)) or (layer6_outputs(1317)));
    layer7_outputs(115) <= not(layer6_outputs(1920)) or (layer6_outputs(937));
    layer7_outputs(116) <= not((layer6_outputs(154)) and (layer6_outputs(905)));
    layer7_outputs(117) <= layer6_outputs(2339);
    layer7_outputs(118) <= (layer6_outputs(4524)) and not (layer6_outputs(1909));
    layer7_outputs(119) <= not(layer6_outputs(2948));
    layer7_outputs(120) <= not(layer6_outputs(2683));
    layer7_outputs(121) <= not(layer6_outputs(4124));
    layer7_outputs(122) <= not(layer6_outputs(986));
    layer7_outputs(123) <= (layer6_outputs(2720)) and not (layer6_outputs(4043));
    layer7_outputs(124) <= not(layer6_outputs(2136)) or (layer6_outputs(4801));
    layer7_outputs(125) <= (layer6_outputs(2021)) and not (layer6_outputs(357));
    layer7_outputs(126) <= (layer6_outputs(2466)) xor (layer6_outputs(2644));
    layer7_outputs(127) <= (layer6_outputs(4583)) and (layer6_outputs(757));
    layer7_outputs(128) <= not((layer6_outputs(1723)) and (layer6_outputs(2858)));
    layer7_outputs(129) <= layer6_outputs(2505);
    layer7_outputs(130) <= (layer6_outputs(2449)) and (layer6_outputs(968));
    layer7_outputs(131) <= layer6_outputs(5002);
    layer7_outputs(132) <= not((layer6_outputs(3761)) and (layer6_outputs(2258)));
    layer7_outputs(133) <= not(layer6_outputs(1715));
    layer7_outputs(134) <= (layer6_outputs(2517)) or (layer6_outputs(4791));
    layer7_outputs(135) <= not(layer6_outputs(2438));
    layer7_outputs(136) <= (layer6_outputs(4998)) and (layer6_outputs(2415));
    layer7_outputs(137) <= layer6_outputs(1932);
    layer7_outputs(138) <= (layer6_outputs(5066)) or (layer6_outputs(1489));
    layer7_outputs(139) <= not((layer6_outputs(3669)) xor (layer6_outputs(4305)));
    layer7_outputs(140) <= not(layer6_outputs(5086));
    layer7_outputs(141) <= (layer6_outputs(2674)) or (layer6_outputs(3467));
    layer7_outputs(142) <= not(layer6_outputs(2080));
    layer7_outputs(143) <= not((layer6_outputs(2992)) xor (layer6_outputs(2218)));
    layer7_outputs(144) <= (layer6_outputs(235)) or (layer6_outputs(2883));
    layer7_outputs(145) <= '0';
    layer7_outputs(146) <= layer6_outputs(3442);
    layer7_outputs(147) <= (layer6_outputs(1670)) and (layer6_outputs(4589));
    layer7_outputs(148) <= (layer6_outputs(3327)) xor (layer6_outputs(4087));
    layer7_outputs(149) <= '1';
    layer7_outputs(150) <= not(layer6_outputs(2129));
    layer7_outputs(151) <= not((layer6_outputs(3504)) xor (layer6_outputs(2777)));
    layer7_outputs(152) <= not((layer6_outputs(680)) xor (layer6_outputs(4861)));
    layer7_outputs(153) <= '0';
    layer7_outputs(154) <= layer6_outputs(3430);
    layer7_outputs(155) <= not(layer6_outputs(2576));
    layer7_outputs(156) <= not(layer6_outputs(1456));
    layer7_outputs(157) <= not(layer6_outputs(4921));
    layer7_outputs(158) <= not((layer6_outputs(4070)) xor (layer6_outputs(4198)));
    layer7_outputs(159) <= not(layer6_outputs(3143));
    layer7_outputs(160) <= (layer6_outputs(4747)) xor (layer6_outputs(2900));
    layer7_outputs(161) <= not(layer6_outputs(4757));
    layer7_outputs(162) <= (layer6_outputs(5045)) or (layer6_outputs(1947));
    layer7_outputs(163) <= not((layer6_outputs(158)) or (layer6_outputs(167)));
    layer7_outputs(164) <= not((layer6_outputs(3349)) and (layer6_outputs(1192)));
    layer7_outputs(165) <= layer6_outputs(2441);
    layer7_outputs(166) <= not(layer6_outputs(5118));
    layer7_outputs(167) <= not(layer6_outputs(3294)) or (layer6_outputs(3177));
    layer7_outputs(168) <= not(layer6_outputs(358));
    layer7_outputs(169) <= not(layer6_outputs(3423));
    layer7_outputs(170) <= not(layer6_outputs(956));
    layer7_outputs(171) <= layer6_outputs(4877);
    layer7_outputs(172) <= not((layer6_outputs(2248)) xor (layer6_outputs(2220)));
    layer7_outputs(173) <= layer6_outputs(3068);
    layer7_outputs(174) <= not((layer6_outputs(4640)) or (layer6_outputs(4551)));
    layer7_outputs(175) <= layer6_outputs(3743);
    layer7_outputs(176) <= not(layer6_outputs(2500));
    layer7_outputs(177) <= not(layer6_outputs(3280));
    layer7_outputs(178) <= (layer6_outputs(647)) and not (layer6_outputs(3239));
    layer7_outputs(179) <= not(layer6_outputs(899));
    layer7_outputs(180) <= not(layer6_outputs(4565)) or (layer6_outputs(776));
    layer7_outputs(181) <= layer6_outputs(596);
    layer7_outputs(182) <= (layer6_outputs(516)) and not (layer6_outputs(793));
    layer7_outputs(183) <= not(layer6_outputs(4039));
    layer7_outputs(184) <= not((layer6_outputs(3427)) xor (layer6_outputs(3849)));
    layer7_outputs(185) <= (layer6_outputs(604)) xor (layer6_outputs(4825));
    layer7_outputs(186) <= not(layer6_outputs(2438)) or (layer6_outputs(4467));
    layer7_outputs(187) <= layer6_outputs(3749);
    layer7_outputs(188) <= not(layer6_outputs(3266)) or (layer6_outputs(1808));
    layer7_outputs(189) <= not(layer6_outputs(922));
    layer7_outputs(190) <= (layer6_outputs(1793)) and (layer6_outputs(2394));
    layer7_outputs(191) <= (layer6_outputs(2872)) and not (layer6_outputs(175));
    layer7_outputs(192) <= not((layer6_outputs(4560)) xor (layer6_outputs(3339)));
    layer7_outputs(193) <= not((layer6_outputs(268)) xor (layer6_outputs(176)));
    layer7_outputs(194) <= not(layer6_outputs(3131));
    layer7_outputs(195) <= layer6_outputs(569);
    layer7_outputs(196) <= not(layer6_outputs(4796));
    layer7_outputs(197) <= layer6_outputs(998);
    layer7_outputs(198) <= (layer6_outputs(3149)) xor (layer6_outputs(2323));
    layer7_outputs(199) <= not(layer6_outputs(4224)) or (layer6_outputs(670));
    layer7_outputs(200) <= not(layer6_outputs(239));
    layer7_outputs(201) <= not(layer6_outputs(3180)) or (layer6_outputs(125));
    layer7_outputs(202) <= not((layer6_outputs(3942)) and (layer6_outputs(4809)));
    layer7_outputs(203) <= (layer6_outputs(230)) or (layer6_outputs(4430));
    layer7_outputs(204) <= not((layer6_outputs(1709)) xor (layer6_outputs(1318)));
    layer7_outputs(205) <= (layer6_outputs(4590)) xor (layer6_outputs(992));
    layer7_outputs(206) <= layer6_outputs(2297);
    layer7_outputs(207) <= (layer6_outputs(3930)) and (layer6_outputs(2235));
    layer7_outputs(208) <= layer6_outputs(1113);
    layer7_outputs(209) <= (layer6_outputs(548)) and not (layer6_outputs(106));
    layer7_outputs(210) <= layer6_outputs(3946);
    layer7_outputs(211) <= not(layer6_outputs(3134)) or (layer6_outputs(1499));
    layer7_outputs(212) <= layer6_outputs(3233);
    layer7_outputs(213) <= not((layer6_outputs(4991)) xor (layer6_outputs(2024)));
    layer7_outputs(214) <= (layer6_outputs(4640)) or (layer6_outputs(3130));
    layer7_outputs(215) <= layer6_outputs(2358);
    layer7_outputs(216) <= not(layer6_outputs(1499));
    layer7_outputs(217) <= layer6_outputs(1236);
    layer7_outputs(218) <= not(layer6_outputs(1068));
    layer7_outputs(219) <= layer6_outputs(3450);
    layer7_outputs(220) <= layer6_outputs(1837);
    layer7_outputs(221) <= not(layer6_outputs(1714));
    layer7_outputs(222) <= not(layer6_outputs(3699));
    layer7_outputs(223) <= (layer6_outputs(1812)) and not (layer6_outputs(330));
    layer7_outputs(224) <= (layer6_outputs(4486)) or (layer6_outputs(2351));
    layer7_outputs(225) <= not((layer6_outputs(2902)) or (layer6_outputs(2334)));
    layer7_outputs(226) <= not(layer6_outputs(3965)) or (layer6_outputs(52));
    layer7_outputs(227) <= not(layer6_outputs(8));
    layer7_outputs(228) <= layer6_outputs(4372);
    layer7_outputs(229) <= layer6_outputs(4793);
    layer7_outputs(230) <= (layer6_outputs(1110)) xor (layer6_outputs(1215));
    layer7_outputs(231) <= not(layer6_outputs(4801));
    layer7_outputs(232) <= layer6_outputs(3548);
    layer7_outputs(233) <= (layer6_outputs(3177)) and (layer6_outputs(339));
    layer7_outputs(234) <= not(layer6_outputs(3069));
    layer7_outputs(235) <= not(layer6_outputs(17)) or (layer6_outputs(816));
    layer7_outputs(236) <= (layer6_outputs(3820)) and not (layer6_outputs(3894));
    layer7_outputs(237) <= not(layer6_outputs(4683));
    layer7_outputs(238) <= layer6_outputs(1613);
    layer7_outputs(239) <= not((layer6_outputs(2363)) xor (layer6_outputs(1303)));
    layer7_outputs(240) <= not(layer6_outputs(4374));
    layer7_outputs(241) <= not(layer6_outputs(2650)) or (layer6_outputs(4994));
    layer7_outputs(242) <= (layer6_outputs(533)) and not (layer6_outputs(2950));
    layer7_outputs(243) <= not((layer6_outputs(3157)) and (layer6_outputs(4111)));
    layer7_outputs(244) <= (layer6_outputs(4533)) and not (layer6_outputs(4642));
    layer7_outputs(245) <= not(layer6_outputs(1061));
    layer7_outputs(246) <= not(layer6_outputs(3997)) or (layer6_outputs(1944));
    layer7_outputs(247) <= (layer6_outputs(4679)) and not (layer6_outputs(2269));
    layer7_outputs(248) <= layer6_outputs(919);
    layer7_outputs(249) <= layer6_outputs(218);
    layer7_outputs(250) <= (layer6_outputs(4363)) and (layer6_outputs(1674));
    layer7_outputs(251) <= not(layer6_outputs(3191));
    layer7_outputs(252) <= not(layer6_outputs(3770));
    layer7_outputs(253) <= not(layer6_outputs(1953)) or (layer6_outputs(47));
    layer7_outputs(254) <= (layer6_outputs(1871)) and not (layer6_outputs(4994));
    layer7_outputs(255) <= layer6_outputs(969);
    layer7_outputs(256) <= (layer6_outputs(3101)) and not (layer6_outputs(3026));
    layer7_outputs(257) <= (layer6_outputs(2546)) and (layer6_outputs(3953));
    layer7_outputs(258) <= not(layer6_outputs(4586));
    layer7_outputs(259) <= layer6_outputs(615);
    layer7_outputs(260) <= layer6_outputs(68);
    layer7_outputs(261) <= layer6_outputs(3470);
    layer7_outputs(262) <= not((layer6_outputs(2109)) xor (layer6_outputs(4966)));
    layer7_outputs(263) <= (layer6_outputs(5029)) xor (layer6_outputs(473));
    layer7_outputs(264) <= not(layer6_outputs(3607));
    layer7_outputs(265) <= (layer6_outputs(3231)) xor (layer6_outputs(3042));
    layer7_outputs(266) <= layer6_outputs(4338);
    layer7_outputs(267) <= layer6_outputs(832);
    layer7_outputs(268) <= (layer6_outputs(3695)) and not (layer6_outputs(4490));
    layer7_outputs(269) <= layer6_outputs(4180);
    layer7_outputs(270) <= not(layer6_outputs(2364)) or (layer6_outputs(566));
    layer7_outputs(271) <= layer6_outputs(4641);
    layer7_outputs(272) <= layer6_outputs(2796);
    layer7_outputs(273) <= not(layer6_outputs(1012));
    layer7_outputs(274) <= layer6_outputs(726);
    layer7_outputs(275) <= not(layer6_outputs(18));
    layer7_outputs(276) <= layer6_outputs(1510);
    layer7_outputs(277) <= not(layer6_outputs(4074));
    layer7_outputs(278) <= layer6_outputs(1476);
    layer7_outputs(279) <= layer6_outputs(2393);
    layer7_outputs(280) <= (layer6_outputs(2817)) and not (layer6_outputs(319));
    layer7_outputs(281) <= not(layer6_outputs(4810));
    layer7_outputs(282) <= layer6_outputs(4053);
    layer7_outputs(283) <= not(layer6_outputs(2017));
    layer7_outputs(284) <= layer6_outputs(2315);
    layer7_outputs(285) <= not((layer6_outputs(3194)) or (layer6_outputs(3633)));
    layer7_outputs(286) <= not((layer6_outputs(3663)) and (layer6_outputs(2957)));
    layer7_outputs(287) <= not(layer6_outputs(4462));
    layer7_outputs(288) <= layer6_outputs(4870);
    layer7_outputs(289) <= (layer6_outputs(729)) and not (layer6_outputs(3719));
    layer7_outputs(290) <= layer6_outputs(733);
    layer7_outputs(291) <= not((layer6_outputs(2572)) and (layer6_outputs(253)));
    layer7_outputs(292) <= not(layer6_outputs(5019));
    layer7_outputs(293) <= layer6_outputs(1380);
    layer7_outputs(294) <= layer6_outputs(1707);
    layer7_outputs(295) <= (layer6_outputs(4511)) and (layer6_outputs(3492));
    layer7_outputs(296) <= (layer6_outputs(2756)) xor (layer6_outputs(1672));
    layer7_outputs(297) <= (layer6_outputs(3139)) and (layer6_outputs(3752));
    layer7_outputs(298) <= layer6_outputs(3061);
    layer7_outputs(299) <= not(layer6_outputs(1694));
    layer7_outputs(300) <= not((layer6_outputs(1161)) and (layer6_outputs(1868)));
    layer7_outputs(301) <= not(layer6_outputs(2755));
    layer7_outputs(302) <= not(layer6_outputs(3102));
    layer7_outputs(303) <= not(layer6_outputs(4905));
    layer7_outputs(304) <= '0';
    layer7_outputs(305) <= not((layer6_outputs(1940)) and (layer6_outputs(1228)));
    layer7_outputs(306) <= layer6_outputs(301);
    layer7_outputs(307) <= not((layer6_outputs(2714)) xor (layer6_outputs(1060)));
    layer7_outputs(308) <= not(layer6_outputs(4010));
    layer7_outputs(309) <= layer6_outputs(1922);
    layer7_outputs(310) <= (layer6_outputs(1974)) and not (layer6_outputs(3070));
    layer7_outputs(311) <= (layer6_outputs(2772)) or (layer6_outputs(3203));
    layer7_outputs(312) <= (layer6_outputs(4891)) xor (layer6_outputs(4219));
    layer7_outputs(313) <= (layer6_outputs(2171)) xor (layer6_outputs(2766));
    layer7_outputs(314) <= not((layer6_outputs(3190)) xor (layer6_outputs(3332)));
    layer7_outputs(315) <= not((layer6_outputs(4227)) or (layer6_outputs(1776)));
    layer7_outputs(316) <= (layer6_outputs(2321)) and (layer6_outputs(1881));
    layer7_outputs(317) <= (layer6_outputs(3988)) and (layer6_outputs(4896));
    layer7_outputs(318) <= (layer6_outputs(1036)) xor (layer6_outputs(2087));
    layer7_outputs(319) <= not(layer6_outputs(1149));
    layer7_outputs(320) <= layer6_outputs(4228);
    layer7_outputs(321) <= layer6_outputs(4146);
    layer7_outputs(322) <= (layer6_outputs(4357)) xor (layer6_outputs(3412));
    layer7_outputs(323) <= not((layer6_outputs(1880)) and (layer6_outputs(2582)));
    layer7_outputs(324) <= not(layer6_outputs(409));
    layer7_outputs(325) <= layer6_outputs(4474);
    layer7_outputs(326) <= layer6_outputs(4777);
    layer7_outputs(327) <= layer6_outputs(465);
    layer7_outputs(328) <= not(layer6_outputs(689)) or (layer6_outputs(3010));
    layer7_outputs(329) <= not(layer6_outputs(1608));
    layer7_outputs(330) <= not(layer6_outputs(4803));
    layer7_outputs(331) <= layer6_outputs(1177);
    layer7_outputs(332) <= (layer6_outputs(2224)) and not (layer6_outputs(531));
    layer7_outputs(333) <= (layer6_outputs(3079)) xor (layer6_outputs(3364));
    layer7_outputs(334) <= not(layer6_outputs(2414));
    layer7_outputs(335) <= not((layer6_outputs(1144)) or (layer6_outputs(2689)));
    layer7_outputs(336) <= layer6_outputs(1707);
    layer7_outputs(337) <= (layer6_outputs(1386)) or (layer6_outputs(425));
    layer7_outputs(338) <= layer6_outputs(3485);
    layer7_outputs(339) <= not(layer6_outputs(260));
    layer7_outputs(340) <= layer6_outputs(582);
    layer7_outputs(341) <= (layer6_outputs(4763)) xor (layer6_outputs(4382));
    layer7_outputs(342) <= not(layer6_outputs(3108));
    layer7_outputs(343) <= not((layer6_outputs(4404)) or (layer6_outputs(4352)));
    layer7_outputs(344) <= not(layer6_outputs(2646));
    layer7_outputs(345) <= not((layer6_outputs(1184)) xor (layer6_outputs(4742)));
    layer7_outputs(346) <= (layer6_outputs(2811)) or (layer6_outputs(1878));
    layer7_outputs(347) <= layer6_outputs(3097);
    layer7_outputs(348) <= (layer6_outputs(3954)) xor (layer6_outputs(2508));
    layer7_outputs(349) <= (layer6_outputs(2340)) and not (layer6_outputs(3360));
    layer7_outputs(350) <= layer6_outputs(1216);
    layer7_outputs(351) <= layer6_outputs(4538);
    layer7_outputs(352) <= not((layer6_outputs(1083)) xor (layer6_outputs(3489)));
    layer7_outputs(353) <= (layer6_outputs(4755)) and not (layer6_outputs(2125));
    layer7_outputs(354) <= not(layer6_outputs(3888));
    layer7_outputs(355) <= not(layer6_outputs(4758));
    layer7_outputs(356) <= (layer6_outputs(4743)) xor (layer6_outputs(1187));
    layer7_outputs(357) <= layer6_outputs(3248);
    layer7_outputs(358) <= not(layer6_outputs(375));
    layer7_outputs(359) <= layer6_outputs(2584);
    layer7_outputs(360) <= (layer6_outputs(2993)) and (layer6_outputs(2440));
    layer7_outputs(361) <= not((layer6_outputs(1500)) xor (layer6_outputs(2934)));
    layer7_outputs(362) <= not(layer6_outputs(1792)) or (layer6_outputs(2948));
    layer7_outputs(363) <= (layer6_outputs(2150)) and not (layer6_outputs(1251));
    layer7_outputs(364) <= not(layer6_outputs(3660)) or (layer6_outputs(3199));
    layer7_outputs(365) <= not(layer6_outputs(4996));
    layer7_outputs(366) <= layer6_outputs(474);
    layer7_outputs(367) <= (layer6_outputs(1964)) xor (layer6_outputs(648));
    layer7_outputs(368) <= not(layer6_outputs(287));
    layer7_outputs(369) <= not(layer6_outputs(1120));
    layer7_outputs(370) <= (layer6_outputs(2649)) and (layer6_outputs(5009));
    layer7_outputs(371) <= not(layer6_outputs(220)) or (layer6_outputs(4121));
    layer7_outputs(372) <= (layer6_outputs(1116)) xor (layer6_outputs(3333));
    layer7_outputs(373) <= layer6_outputs(3361);
    layer7_outputs(374) <= (layer6_outputs(3449)) and not (layer6_outputs(1593));
    layer7_outputs(375) <= not((layer6_outputs(3510)) or (layer6_outputs(2161)));
    layer7_outputs(376) <= not((layer6_outputs(1261)) and (layer6_outputs(2699)));
    layer7_outputs(377) <= (layer6_outputs(4059)) and not (layer6_outputs(3908));
    layer7_outputs(378) <= not(layer6_outputs(2511));
    layer7_outputs(379) <= not((layer6_outputs(1302)) or (layer6_outputs(3132)));
    layer7_outputs(380) <= layer6_outputs(3207);
    layer7_outputs(381) <= (layer6_outputs(832)) and (layer6_outputs(3302));
    layer7_outputs(382) <= (layer6_outputs(2852)) and not (layer6_outputs(1799));
    layer7_outputs(383) <= (layer6_outputs(3355)) or (layer6_outputs(2935));
    layer7_outputs(384) <= not((layer6_outputs(4395)) or (layer6_outputs(3350)));
    layer7_outputs(385) <= not(layer6_outputs(1617));
    layer7_outputs(386) <= not(layer6_outputs(4581));
    layer7_outputs(387) <= (layer6_outputs(3445)) xor (layer6_outputs(376));
    layer7_outputs(388) <= not((layer6_outputs(4911)) xor (layer6_outputs(138)));
    layer7_outputs(389) <= layer6_outputs(1150);
    layer7_outputs(390) <= not(layer6_outputs(3082)) or (layer6_outputs(2460));
    layer7_outputs(391) <= not((layer6_outputs(3814)) or (layer6_outputs(2232)));
    layer7_outputs(392) <= layer6_outputs(1153);
    layer7_outputs(393) <= not(layer6_outputs(3997)) or (layer6_outputs(1779));
    layer7_outputs(394) <= (layer6_outputs(2301)) and not (layer6_outputs(3751));
    layer7_outputs(395) <= (layer6_outputs(2168)) and (layer6_outputs(2801));
    layer7_outputs(396) <= (layer6_outputs(4413)) and not (layer6_outputs(3906));
    layer7_outputs(397) <= (layer6_outputs(4193)) and (layer6_outputs(997));
    layer7_outputs(398) <= not(layer6_outputs(4959));
    layer7_outputs(399) <= layer6_outputs(411);
    layer7_outputs(400) <= not((layer6_outputs(4755)) or (layer6_outputs(3552)));
    layer7_outputs(401) <= layer6_outputs(3357);
    layer7_outputs(402) <= '1';
    layer7_outputs(403) <= not((layer6_outputs(489)) xor (layer6_outputs(4170)));
    layer7_outputs(404) <= layer6_outputs(4095);
    layer7_outputs(405) <= layer6_outputs(2663);
    layer7_outputs(406) <= not(layer6_outputs(3677));
    layer7_outputs(407) <= not((layer6_outputs(1393)) and (layer6_outputs(240)));
    layer7_outputs(408) <= not((layer6_outputs(1075)) xor (layer6_outputs(1900)));
    layer7_outputs(409) <= not((layer6_outputs(393)) or (layer6_outputs(1711)));
    layer7_outputs(410) <= not(layer6_outputs(2479));
    layer7_outputs(411) <= not((layer6_outputs(2685)) or (layer6_outputs(3288)));
    layer7_outputs(412) <= '0';
    layer7_outputs(413) <= layer6_outputs(3348);
    layer7_outputs(414) <= not(layer6_outputs(5078)) or (layer6_outputs(2409));
    layer7_outputs(415) <= layer6_outputs(1163);
    layer7_outputs(416) <= (layer6_outputs(1618)) and (layer6_outputs(375));
    layer7_outputs(417) <= (layer6_outputs(1804)) and not (layer6_outputs(951));
    layer7_outputs(418) <= layer6_outputs(1985);
    layer7_outputs(419) <= not((layer6_outputs(1190)) xor (layer6_outputs(337)));
    layer7_outputs(420) <= '0';
    layer7_outputs(421) <= (layer6_outputs(3311)) and not (layer6_outputs(5001));
    layer7_outputs(422) <= layer6_outputs(2159);
    layer7_outputs(423) <= (layer6_outputs(5023)) xor (layer6_outputs(4256));
    layer7_outputs(424) <= not((layer6_outputs(1298)) and (layer6_outputs(1882)));
    layer7_outputs(425) <= layer6_outputs(2487);
    layer7_outputs(426) <= (layer6_outputs(1389)) and (layer6_outputs(400));
    layer7_outputs(427) <= layer6_outputs(4207);
    layer7_outputs(428) <= (layer6_outputs(4281)) and (layer6_outputs(283));
    layer7_outputs(429) <= not(layer6_outputs(4588));
    layer7_outputs(430) <= not((layer6_outputs(3282)) or (layer6_outputs(4131)));
    layer7_outputs(431) <= not((layer6_outputs(3958)) or (layer6_outputs(404)));
    layer7_outputs(432) <= (layer6_outputs(4566)) xor (layer6_outputs(2252));
    layer7_outputs(433) <= not(layer6_outputs(3809));
    layer7_outputs(434) <= (layer6_outputs(1366)) xor (layer6_outputs(4172));
    layer7_outputs(435) <= not(layer6_outputs(2591));
    layer7_outputs(436) <= (layer6_outputs(1708)) xor (layer6_outputs(1930));
    layer7_outputs(437) <= layer6_outputs(560);
    layer7_outputs(438) <= not(layer6_outputs(2579)) or (layer6_outputs(867));
    layer7_outputs(439) <= layer6_outputs(3668);
    layer7_outputs(440) <= (layer6_outputs(160)) or (layer6_outputs(1372));
    layer7_outputs(441) <= not((layer6_outputs(4642)) and (layer6_outputs(978)));
    layer7_outputs(442) <= layer6_outputs(2132);
    layer7_outputs(443) <= layer6_outputs(2493);
    layer7_outputs(444) <= layer6_outputs(1802);
    layer7_outputs(445) <= not((layer6_outputs(363)) xor (layer6_outputs(3641)));
    layer7_outputs(446) <= not(layer6_outputs(3461));
    layer7_outputs(447) <= layer6_outputs(644);
    layer7_outputs(448) <= (layer6_outputs(2971)) xor (layer6_outputs(2498));
    layer7_outputs(449) <= not(layer6_outputs(4260));
    layer7_outputs(450) <= not(layer6_outputs(5089));
    layer7_outputs(451) <= not(layer6_outputs(4391));
    layer7_outputs(452) <= not((layer6_outputs(2382)) and (layer6_outputs(3920)));
    layer7_outputs(453) <= layer6_outputs(2032);
    layer7_outputs(454) <= not((layer6_outputs(1568)) or (layer6_outputs(4289)));
    layer7_outputs(455) <= not(layer6_outputs(2719)) or (layer6_outputs(1867));
    layer7_outputs(456) <= not(layer6_outputs(3468));
    layer7_outputs(457) <= not((layer6_outputs(877)) or (layer6_outputs(2827)));
    layer7_outputs(458) <= layer6_outputs(3854);
    layer7_outputs(459) <= not((layer6_outputs(958)) xor (layer6_outputs(4380)));
    layer7_outputs(460) <= not((layer6_outputs(1343)) or (layer6_outputs(787)));
    layer7_outputs(461) <= layer6_outputs(413);
    layer7_outputs(462) <= (layer6_outputs(3887)) xor (layer6_outputs(5021));
    layer7_outputs(463) <= layer6_outputs(2225);
    layer7_outputs(464) <= not(layer6_outputs(1849));
    layer7_outputs(465) <= layer6_outputs(1861);
    layer7_outputs(466) <= (layer6_outputs(274)) and not (layer6_outputs(2586));
    layer7_outputs(467) <= '1';
    layer7_outputs(468) <= not((layer6_outputs(4630)) and (layer6_outputs(2496)));
    layer7_outputs(469) <= layer6_outputs(256);
    layer7_outputs(470) <= layer6_outputs(4061);
    layer7_outputs(471) <= layer6_outputs(4882);
    layer7_outputs(472) <= not(layer6_outputs(2031));
    layer7_outputs(473) <= layer6_outputs(3099);
    layer7_outputs(474) <= (layer6_outputs(4190)) and not (layer6_outputs(3909));
    layer7_outputs(475) <= not(layer6_outputs(1739));
    layer7_outputs(476) <= not((layer6_outputs(1315)) xor (layer6_outputs(700)));
    layer7_outputs(477) <= layer6_outputs(2918);
    layer7_outputs(478) <= layer6_outputs(2806);
    layer7_outputs(479) <= not(layer6_outputs(4275)) or (layer6_outputs(4120));
    layer7_outputs(480) <= '1';
    layer7_outputs(481) <= (layer6_outputs(1430)) and (layer6_outputs(262));
    layer7_outputs(482) <= not(layer6_outputs(3756)) or (layer6_outputs(2009));
    layer7_outputs(483) <= (layer6_outputs(1173)) xor (layer6_outputs(1521));
    layer7_outputs(484) <= not(layer6_outputs(5034));
    layer7_outputs(485) <= layer6_outputs(1260);
    layer7_outputs(486) <= not((layer6_outputs(994)) xor (layer6_outputs(1522)));
    layer7_outputs(487) <= not(layer6_outputs(3536));
    layer7_outputs(488) <= layer6_outputs(2335);
    layer7_outputs(489) <= not(layer6_outputs(3323));
    layer7_outputs(490) <= not(layer6_outputs(5090));
    layer7_outputs(491) <= not(layer6_outputs(2367));
    layer7_outputs(492) <= (layer6_outputs(12)) xor (layer6_outputs(4473));
    layer7_outputs(493) <= not((layer6_outputs(3380)) and (layer6_outputs(3981)));
    layer7_outputs(494) <= not(layer6_outputs(2557));
    layer7_outputs(495) <= not((layer6_outputs(2532)) and (layer6_outputs(3593)));
    layer7_outputs(496) <= not(layer6_outputs(1809));
    layer7_outputs(497) <= not((layer6_outputs(3089)) xor (layer6_outputs(765)));
    layer7_outputs(498) <= (layer6_outputs(3905)) xor (layer6_outputs(1340));
    layer7_outputs(499) <= layer6_outputs(1480);
    layer7_outputs(500) <= not((layer6_outputs(3302)) and (layer6_outputs(3194)));
    layer7_outputs(501) <= layer6_outputs(4437);
    layer7_outputs(502) <= not(layer6_outputs(639)) or (layer6_outputs(2568));
    layer7_outputs(503) <= layer6_outputs(3515);
    layer7_outputs(504) <= layer6_outputs(3263);
    layer7_outputs(505) <= layer6_outputs(55);
    layer7_outputs(506) <= layer6_outputs(20);
    layer7_outputs(507) <= (layer6_outputs(4526)) and not (layer6_outputs(380));
    layer7_outputs(508) <= '0';
    layer7_outputs(509) <= not(layer6_outputs(1811));
    layer7_outputs(510) <= layer6_outputs(1819);
    layer7_outputs(511) <= not(layer6_outputs(3624)) or (layer6_outputs(2664));
    layer7_outputs(512) <= not(layer6_outputs(91));
    layer7_outputs(513) <= not((layer6_outputs(3781)) and (layer6_outputs(344)));
    layer7_outputs(514) <= not((layer6_outputs(2811)) or (layer6_outputs(5106)));
    layer7_outputs(515) <= not(layer6_outputs(4650));
    layer7_outputs(516) <= not((layer6_outputs(2814)) and (layer6_outputs(3902)));
    layer7_outputs(517) <= not(layer6_outputs(2914)) or (layer6_outputs(3441));
    layer7_outputs(518) <= (layer6_outputs(4047)) and not (layer6_outputs(3724));
    layer7_outputs(519) <= layer6_outputs(719);
    layer7_outputs(520) <= not(layer6_outputs(3571));
    layer7_outputs(521) <= (layer6_outputs(3899)) or (layer6_outputs(4044));
    layer7_outputs(522) <= layer6_outputs(4724);
    layer7_outputs(523) <= not(layer6_outputs(2191)) or (layer6_outputs(2553));
    layer7_outputs(524) <= not(layer6_outputs(207));
    layer7_outputs(525) <= layer6_outputs(3542);
    layer7_outputs(526) <= not(layer6_outputs(3124));
    layer7_outputs(527) <= not((layer6_outputs(4903)) or (layer6_outputs(3819)));
    layer7_outputs(528) <= not(layer6_outputs(2615));
    layer7_outputs(529) <= not((layer6_outputs(3737)) xor (layer6_outputs(3111)));
    layer7_outputs(530) <= layer6_outputs(4387);
    layer7_outputs(531) <= not(layer6_outputs(2931)) or (layer6_outputs(2423));
    layer7_outputs(532) <= not(layer6_outputs(3407));
    layer7_outputs(533) <= not((layer6_outputs(862)) or (layer6_outputs(3586)));
    layer7_outputs(534) <= not((layer6_outputs(690)) and (layer6_outputs(407)));
    layer7_outputs(535) <= not((layer6_outputs(3693)) xor (layer6_outputs(807)));
    layer7_outputs(536) <= (layer6_outputs(1586)) and (layer6_outputs(568));
    layer7_outputs(537) <= '1';
    layer7_outputs(538) <= not(layer6_outputs(3686)) or (layer6_outputs(3802));
    layer7_outputs(539) <= layer6_outputs(3728);
    layer7_outputs(540) <= (layer6_outputs(4001)) xor (layer6_outputs(3025));
    layer7_outputs(541) <= not((layer6_outputs(5041)) xor (layer6_outputs(11)));
    layer7_outputs(542) <= layer6_outputs(211);
    layer7_outputs(543) <= not(layer6_outputs(1827)) or (layer6_outputs(1354));
    layer7_outputs(544) <= not((layer6_outputs(1635)) or (layer6_outputs(364)));
    layer7_outputs(545) <= not(layer6_outputs(2444));
    layer7_outputs(546) <= (layer6_outputs(1851)) and not (layer6_outputs(293));
    layer7_outputs(547) <= layer6_outputs(3155);
    layer7_outputs(548) <= layer6_outputs(3549);
    layer7_outputs(549) <= not(layer6_outputs(3664));
    layer7_outputs(550) <= not(layer6_outputs(1034));
    layer7_outputs(551) <= not(layer6_outputs(1210));
    layer7_outputs(552) <= not(layer6_outputs(3889));
    layer7_outputs(553) <= not((layer6_outputs(3814)) and (layer6_outputs(2857)));
    layer7_outputs(554) <= not(layer6_outputs(5017));
    layer7_outputs(555) <= '0';
    layer7_outputs(556) <= layer6_outputs(3818);
    layer7_outputs(557) <= not((layer6_outputs(2227)) or (layer6_outputs(775)));
    layer7_outputs(558) <= not((layer6_outputs(822)) or (layer6_outputs(3648)));
    layer7_outputs(559) <= not((layer6_outputs(3503)) and (layer6_outputs(3625)));
    layer7_outputs(560) <= (layer6_outputs(3675)) and not (layer6_outputs(1569));
    layer7_outputs(561) <= (layer6_outputs(4847)) or (layer6_outputs(141));
    layer7_outputs(562) <= not((layer6_outputs(3026)) and (layer6_outputs(901)));
    layer7_outputs(563) <= layer6_outputs(570);
    layer7_outputs(564) <= not((layer6_outputs(497)) and (layer6_outputs(72)));
    layer7_outputs(565) <= not(layer6_outputs(3867));
    layer7_outputs(566) <= not((layer6_outputs(1453)) and (layer6_outputs(1991)));
    layer7_outputs(567) <= not((layer6_outputs(3159)) or (layer6_outputs(3534)));
    layer7_outputs(568) <= (layer6_outputs(265)) xor (layer6_outputs(2817));
    layer7_outputs(569) <= not((layer6_outputs(666)) or (layer6_outputs(4245)));
    layer7_outputs(570) <= layer6_outputs(1194);
    layer7_outputs(571) <= not((layer6_outputs(944)) or (layer6_outputs(2690)));
    layer7_outputs(572) <= not(layer6_outputs(2411));
    layer7_outputs(573) <= '1';
    layer7_outputs(574) <= (layer6_outputs(3068)) xor (layer6_outputs(888));
    layer7_outputs(575) <= '0';
    layer7_outputs(576) <= not(layer6_outputs(3127)) or (layer6_outputs(2309));
    layer7_outputs(577) <= not(layer6_outputs(2069)) or (layer6_outputs(3442));
    layer7_outputs(578) <= not((layer6_outputs(3197)) or (layer6_outputs(2147)));
    layer7_outputs(579) <= (layer6_outputs(4538)) and not (layer6_outputs(4445));
    layer7_outputs(580) <= (layer6_outputs(2547)) and (layer6_outputs(1703));
    layer7_outputs(581) <= '0';
    layer7_outputs(582) <= (layer6_outputs(2357)) or (layer6_outputs(3574));
    layer7_outputs(583) <= layer6_outputs(1103);
    layer7_outputs(584) <= not((layer6_outputs(3396)) or (layer6_outputs(1244)));
    layer7_outputs(585) <= not(layer6_outputs(2436));
    layer7_outputs(586) <= (layer6_outputs(2911)) xor (layer6_outputs(316));
    layer7_outputs(587) <= not(layer6_outputs(3035));
    layer7_outputs(588) <= layer6_outputs(1127);
    layer7_outputs(589) <= not((layer6_outputs(3680)) or (layer6_outputs(4071)));
    layer7_outputs(590) <= '0';
    layer7_outputs(591) <= not(layer6_outputs(4548));
    layer7_outputs(592) <= layer6_outputs(4127);
    layer7_outputs(593) <= '1';
    layer7_outputs(594) <= not((layer6_outputs(3295)) or (layer6_outputs(54)));
    layer7_outputs(595) <= not(layer6_outputs(4517)) or (layer6_outputs(1450));
    layer7_outputs(596) <= not(layer6_outputs(3156));
    layer7_outputs(597) <= not(layer6_outputs(3765));
    layer7_outputs(598) <= not((layer6_outputs(65)) and (layer6_outputs(1905)));
    layer7_outputs(599) <= '0';
    layer7_outputs(600) <= layer6_outputs(4448);
    layer7_outputs(601) <= layer6_outputs(1190);
    layer7_outputs(602) <= not(layer6_outputs(2738));
    layer7_outputs(603) <= not(layer6_outputs(5016));
    layer7_outputs(604) <= layer6_outputs(2273);
    layer7_outputs(605) <= '1';
    layer7_outputs(606) <= (layer6_outputs(2008)) xor (layer6_outputs(576));
    layer7_outputs(607) <= not(layer6_outputs(361));
    layer7_outputs(608) <= (layer6_outputs(1242)) and not (layer6_outputs(4731));
    layer7_outputs(609) <= (layer6_outputs(78)) xor (layer6_outputs(2063));
    layer7_outputs(610) <= layer6_outputs(1453);
    layer7_outputs(611) <= not((layer6_outputs(2774)) xor (layer6_outputs(3990)));
    layer7_outputs(612) <= not(layer6_outputs(2934));
    layer7_outputs(613) <= '0';
    layer7_outputs(614) <= layer6_outputs(131);
    layer7_outputs(615) <= (layer6_outputs(335)) and not (layer6_outputs(4672));
    layer7_outputs(616) <= (layer6_outputs(3148)) xor (layer6_outputs(582));
    layer7_outputs(617) <= not(layer6_outputs(4927));
    layer7_outputs(618) <= (layer6_outputs(3488)) or (layer6_outputs(973));
    layer7_outputs(619) <= not((layer6_outputs(2685)) and (layer6_outputs(2710)));
    layer7_outputs(620) <= (layer6_outputs(199)) and (layer6_outputs(4780));
    layer7_outputs(621) <= (layer6_outputs(4199)) xor (layer6_outputs(1768));
    layer7_outputs(622) <= not((layer6_outputs(3040)) and (layer6_outputs(2130)));
    layer7_outputs(623) <= not(layer6_outputs(3824));
    layer7_outputs(624) <= (layer6_outputs(3872)) and not (layer6_outputs(433));
    layer7_outputs(625) <= (layer6_outputs(4838)) or (layer6_outputs(4158));
    layer7_outputs(626) <= (layer6_outputs(377)) and not (layer6_outputs(2567));
    layer7_outputs(627) <= (layer6_outputs(4754)) or (layer6_outputs(2613));
    layer7_outputs(628) <= not(layer6_outputs(2156)) or (layer6_outputs(112));
    layer7_outputs(629) <= not(layer6_outputs(3341)) or (layer6_outputs(701));
    layer7_outputs(630) <= not(layer6_outputs(4184));
    layer7_outputs(631) <= not(layer6_outputs(410));
    layer7_outputs(632) <= not((layer6_outputs(1789)) and (layer6_outputs(3380)));
    layer7_outputs(633) <= not(layer6_outputs(1636));
    layer7_outputs(634) <= not(layer6_outputs(2542));
    layer7_outputs(635) <= not((layer6_outputs(2137)) xor (layer6_outputs(838)));
    layer7_outputs(636) <= layer6_outputs(2105);
    layer7_outputs(637) <= (layer6_outputs(394)) or (layer6_outputs(216));
    layer7_outputs(638) <= layer6_outputs(4306);
    layer7_outputs(639) <= '0';
    layer7_outputs(640) <= not((layer6_outputs(4976)) xor (layer6_outputs(607)));
    layer7_outputs(641) <= layer6_outputs(2980);
    layer7_outputs(642) <= layer6_outputs(229);
    layer7_outputs(643) <= '1';
    layer7_outputs(644) <= (layer6_outputs(3639)) and not (layer6_outputs(2108));
    layer7_outputs(645) <= not(layer6_outputs(2239));
    layer7_outputs(646) <= not(layer6_outputs(4662));
    layer7_outputs(647) <= not(layer6_outputs(3810));
    layer7_outputs(648) <= not(layer6_outputs(1727));
    layer7_outputs(649) <= not((layer6_outputs(4291)) xor (layer6_outputs(3581)));
    layer7_outputs(650) <= layer6_outputs(2513);
    layer7_outputs(651) <= not(layer6_outputs(1355)) or (layer6_outputs(1312));
    layer7_outputs(652) <= (layer6_outputs(3605)) and not (layer6_outputs(99));
    layer7_outputs(653) <= not(layer6_outputs(3931));
    layer7_outputs(654) <= layer6_outputs(1981);
    layer7_outputs(655) <= not(layer6_outputs(3820)) or (layer6_outputs(4235));
    layer7_outputs(656) <= layer6_outputs(4919);
    layer7_outputs(657) <= not(layer6_outputs(4530));
    layer7_outputs(658) <= not(layer6_outputs(4703));
    layer7_outputs(659) <= (layer6_outputs(2843)) and not (layer6_outputs(3091));
    layer7_outputs(660) <= not((layer6_outputs(4231)) or (layer6_outputs(1412)));
    layer7_outputs(661) <= layer6_outputs(4578);
    layer7_outputs(662) <= (layer6_outputs(3888)) xor (layer6_outputs(635));
    layer7_outputs(663) <= '1';
    layer7_outputs(664) <= not(layer6_outputs(3285)) or (layer6_outputs(4797));
    layer7_outputs(665) <= not(layer6_outputs(2102));
    layer7_outputs(666) <= layer6_outputs(704);
    layer7_outputs(667) <= not(layer6_outputs(2999)) or (layer6_outputs(4788));
    layer7_outputs(668) <= (layer6_outputs(2742)) or (layer6_outputs(654));
    layer7_outputs(669) <= not(layer6_outputs(4059)) or (layer6_outputs(1145));
    layer7_outputs(670) <= not(layer6_outputs(3630));
    layer7_outputs(671) <= not(layer6_outputs(1925));
    layer7_outputs(672) <= not(layer6_outputs(4092));
    layer7_outputs(673) <= not(layer6_outputs(976)) or (layer6_outputs(312));
    layer7_outputs(674) <= (layer6_outputs(3590)) and not (layer6_outputs(2905));
    layer7_outputs(675) <= not(layer6_outputs(898));
    layer7_outputs(676) <= not(layer6_outputs(4457)) or (layer6_outputs(2220));
    layer7_outputs(677) <= not(layer6_outputs(379)) or (layer6_outputs(3382));
    layer7_outputs(678) <= '0';
    layer7_outputs(679) <= not((layer6_outputs(2929)) and (layer6_outputs(17)));
    layer7_outputs(680) <= layer6_outputs(4261);
    layer7_outputs(681) <= not(layer6_outputs(1364)) or (layer6_outputs(3317));
    layer7_outputs(682) <= (layer6_outputs(3581)) xor (layer6_outputs(3640));
    layer7_outputs(683) <= not((layer6_outputs(4104)) xor (layer6_outputs(398)));
    layer7_outputs(684) <= (layer6_outputs(4491)) and not (layer6_outputs(3572));
    layer7_outputs(685) <= layer6_outputs(332);
    layer7_outputs(686) <= not((layer6_outputs(4441)) xor (layer6_outputs(2494)));
    layer7_outputs(687) <= not(layer6_outputs(2408));
    layer7_outputs(688) <= (layer6_outputs(3107)) and (layer6_outputs(2874));
    layer7_outputs(689) <= not(layer6_outputs(5000));
    layer7_outputs(690) <= not(layer6_outputs(791));
    layer7_outputs(691) <= layer6_outputs(5056);
    layer7_outputs(692) <= layer6_outputs(2570);
    layer7_outputs(693) <= not((layer6_outputs(196)) xor (layer6_outputs(1454)));
    layer7_outputs(694) <= not(layer6_outputs(3938));
    layer7_outputs(695) <= layer6_outputs(4309);
    layer7_outputs(696) <= layer6_outputs(4343);
    layer7_outputs(697) <= (layer6_outputs(286)) xor (layer6_outputs(2234));
    layer7_outputs(698) <= (layer6_outputs(4443)) or (layer6_outputs(1041));
    layer7_outputs(699) <= layer6_outputs(2437);
    layer7_outputs(700) <= not(layer6_outputs(2355));
    layer7_outputs(701) <= not(layer6_outputs(501)) or (layer6_outputs(5071));
    layer7_outputs(702) <= not(layer6_outputs(3075));
    layer7_outputs(703) <= not(layer6_outputs(739)) or (layer6_outputs(3416));
    layer7_outputs(704) <= not(layer6_outputs(2717));
    layer7_outputs(705) <= not(layer6_outputs(3119));
    layer7_outputs(706) <= layer6_outputs(3956);
    layer7_outputs(707) <= layer6_outputs(2800);
    layer7_outputs(708) <= not((layer6_outputs(2806)) xor (layer6_outputs(1828)));
    layer7_outputs(709) <= not(layer6_outputs(4687));
    layer7_outputs(710) <= not(layer6_outputs(3408)) or (layer6_outputs(1370));
    layer7_outputs(711) <= not((layer6_outputs(2167)) and (layer6_outputs(537)));
    layer7_outputs(712) <= '1';
    layer7_outputs(713) <= not((layer6_outputs(2910)) xor (layer6_outputs(3259)));
    layer7_outputs(714) <= layer6_outputs(2818);
    layer7_outputs(715) <= (layer6_outputs(3001)) xor (layer6_outputs(933));
    layer7_outputs(716) <= (layer6_outputs(1956)) and not (layer6_outputs(1833));
    layer7_outputs(717) <= not(layer6_outputs(3077));
    layer7_outputs(718) <= layer6_outputs(4661);
    layer7_outputs(719) <= not(layer6_outputs(2006));
    layer7_outputs(720) <= not((layer6_outputs(4989)) xor (layer6_outputs(1845)));
    layer7_outputs(721) <= not((layer6_outputs(2238)) xor (layer6_outputs(2162)));
    layer7_outputs(722) <= layer6_outputs(1958);
    layer7_outputs(723) <= not((layer6_outputs(1748)) and (layer6_outputs(498)));
    layer7_outputs(724) <= (layer6_outputs(3729)) or (layer6_outputs(4026));
    layer7_outputs(725) <= not(layer6_outputs(4571));
    layer7_outputs(726) <= not((layer6_outputs(3409)) xor (layer6_outputs(1488)));
    layer7_outputs(727) <= not(layer6_outputs(584));
    layer7_outputs(728) <= not((layer6_outputs(2779)) or (layer6_outputs(2221)));
    layer7_outputs(729) <= not((layer6_outputs(1663)) xor (layer6_outputs(557)));
    layer7_outputs(730) <= not(layer6_outputs(1665));
    layer7_outputs(731) <= layer6_outputs(4910);
    layer7_outputs(732) <= (layer6_outputs(3334)) or (layer6_outputs(64));
    layer7_outputs(733) <= not(layer6_outputs(2886));
    layer7_outputs(734) <= (layer6_outputs(1544)) and not (layer6_outputs(124));
    layer7_outputs(735) <= layer6_outputs(1786);
    layer7_outputs(736) <= not((layer6_outputs(2513)) and (layer6_outputs(4911)));
    layer7_outputs(737) <= layer6_outputs(1454);
    layer7_outputs(738) <= not((layer6_outputs(2509)) and (layer6_outputs(1810)));
    layer7_outputs(739) <= layer6_outputs(4840);
    layer7_outputs(740) <= not(layer6_outputs(4049));
    layer7_outputs(741) <= not(layer6_outputs(2450));
    layer7_outputs(742) <= (layer6_outputs(1152)) xor (layer6_outputs(4980));
    layer7_outputs(743) <= (layer6_outputs(707)) and not (layer6_outputs(1829));
    layer7_outputs(744) <= not(layer6_outputs(427));
    layer7_outputs(745) <= not(layer6_outputs(4884));
    layer7_outputs(746) <= layer6_outputs(2651);
    layer7_outputs(747) <= (layer6_outputs(1913)) and (layer6_outputs(2531));
    layer7_outputs(748) <= layer6_outputs(2631);
    layer7_outputs(749) <= (layer6_outputs(3720)) and not (layer6_outputs(2732));
    layer7_outputs(750) <= (layer6_outputs(4422)) and (layer6_outputs(2267));
    layer7_outputs(751) <= not(layer6_outputs(822));
    layer7_outputs(752) <= '1';
    layer7_outputs(753) <= (layer6_outputs(3081)) and (layer6_outputs(980));
    layer7_outputs(754) <= (layer6_outputs(1612)) and not (layer6_outputs(4601));
    layer7_outputs(755) <= not(layer6_outputs(738));
    layer7_outputs(756) <= not((layer6_outputs(532)) xor (layer6_outputs(5046)));
    layer7_outputs(757) <= layer6_outputs(4759);
    layer7_outputs(758) <= (layer6_outputs(386)) xor (layer6_outputs(3557));
    layer7_outputs(759) <= not(layer6_outputs(1863));
    layer7_outputs(760) <= (layer6_outputs(1340)) xor (layer6_outputs(1755));
    layer7_outputs(761) <= (layer6_outputs(4028)) and (layer6_outputs(4707));
    layer7_outputs(762) <= (layer6_outputs(3115)) or (layer6_outputs(2870));
    layer7_outputs(763) <= not(layer6_outputs(1708));
    layer7_outputs(764) <= not(layer6_outputs(3867));
    layer7_outputs(765) <= layer6_outputs(3138);
    layer7_outputs(766) <= not(layer6_outputs(2946));
    layer7_outputs(767) <= (layer6_outputs(714)) or (layer6_outputs(4852));
    layer7_outputs(768) <= not(layer6_outputs(2020)) or (layer6_outputs(368));
    layer7_outputs(769) <= not(layer6_outputs(4280));
    layer7_outputs(770) <= not((layer6_outputs(2465)) xor (layer6_outputs(4677)));
    layer7_outputs(771) <= not(layer6_outputs(4297)) or (layer6_outputs(2361));
    layer7_outputs(772) <= (layer6_outputs(2522)) xor (layer6_outputs(2005));
    layer7_outputs(773) <= not(layer6_outputs(2995)) or (layer6_outputs(1425));
    layer7_outputs(774) <= layer6_outputs(5103);
    layer7_outputs(775) <= (layer6_outputs(3074)) and not (layer6_outputs(1976));
    layer7_outputs(776) <= (layer6_outputs(3614)) or (layer6_outputs(1691));
    layer7_outputs(777) <= (layer6_outputs(4210)) and not (layer6_outputs(316));
    layer7_outputs(778) <= layer6_outputs(552);
    layer7_outputs(779) <= layer6_outputs(4846);
    layer7_outputs(780) <= (layer6_outputs(4056)) and (layer6_outputs(1800));
    layer7_outputs(781) <= not((layer6_outputs(3014)) xor (layer6_outputs(3654)));
    layer7_outputs(782) <= layer6_outputs(679);
    layer7_outputs(783) <= (layer6_outputs(861)) and not (layer6_outputs(1115));
    layer7_outputs(784) <= layer6_outputs(868);
    layer7_outputs(785) <= not(layer6_outputs(1429));
    layer7_outputs(786) <= (layer6_outputs(276)) and (layer6_outputs(2670));
    layer7_outputs(787) <= layer6_outputs(4103);
    layer7_outputs(788) <= not(layer6_outputs(3883));
    layer7_outputs(789) <= (layer6_outputs(1018)) and (layer6_outputs(2135));
    layer7_outputs(790) <= (layer6_outputs(1845)) xor (layer6_outputs(4937));
    layer7_outputs(791) <= not(layer6_outputs(2849));
    layer7_outputs(792) <= not((layer6_outputs(22)) and (layer6_outputs(2628)));
    layer7_outputs(793) <= (layer6_outputs(4898)) or (layer6_outputs(3116));
    layer7_outputs(794) <= '0';
    layer7_outputs(795) <= not(layer6_outputs(5031));
    layer7_outputs(796) <= layer6_outputs(3680);
    layer7_outputs(797) <= layer6_outputs(264);
    layer7_outputs(798) <= (layer6_outputs(3631)) and not (layer6_outputs(226));
    layer7_outputs(799) <= layer6_outputs(2196);
    layer7_outputs(800) <= layer6_outputs(4021);
    layer7_outputs(801) <= not(layer6_outputs(4433));
    layer7_outputs(802) <= not(layer6_outputs(2956));
    layer7_outputs(803) <= not((layer6_outputs(5068)) and (layer6_outputs(4867)));
    layer7_outputs(804) <= (layer6_outputs(1515)) xor (layer6_outputs(1324));
    layer7_outputs(805) <= layer6_outputs(318);
    layer7_outputs(806) <= layer6_outputs(4706);
    layer7_outputs(807) <= not(layer6_outputs(5034)) or (layer6_outputs(1852));
    layer7_outputs(808) <= not(layer6_outputs(4657));
    layer7_outputs(809) <= layer6_outputs(1816);
    layer7_outputs(810) <= layer6_outputs(2521);
    layer7_outputs(811) <= layer6_outputs(558);
    layer7_outputs(812) <= layer6_outputs(388);
    layer7_outputs(813) <= not(layer6_outputs(1501));
    layer7_outputs(814) <= (layer6_outputs(77)) and not (layer6_outputs(5031));
    layer7_outputs(815) <= (layer6_outputs(1822)) and (layer6_outputs(4864));
    layer7_outputs(816) <= not(layer6_outputs(720)) or (layer6_outputs(3319));
    layer7_outputs(817) <= (layer6_outputs(4758)) and (layer6_outputs(448));
    layer7_outputs(818) <= not(layer6_outputs(979));
    layer7_outputs(819) <= not(layer6_outputs(4554));
    layer7_outputs(820) <= not(layer6_outputs(5065)) or (layer6_outputs(1349));
    layer7_outputs(821) <= layer6_outputs(4779);
    layer7_outputs(822) <= (layer6_outputs(1935)) xor (layer6_outputs(4871));
    layer7_outputs(823) <= layer6_outputs(3305);
    layer7_outputs(824) <= layer6_outputs(4280);
    layer7_outputs(825) <= layer6_outputs(1823);
    layer7_outputs(826) <= not(layer6_outputs(1754)) or (layer6_outputs(3591));
    layer7_outputs(827) <= (layer6_outputs(4423)) and not (layer6_outputs(4351));
    layer7_outputs(828) <= layer6_outputs(1150);
    layer7_outputs(829) <= not(layer6_outputs(2853));
    layer7_outputs(830) <= not(layer6_outputs(2906));
    layer7_outputs(831) <= (layer6_outputs(3659)) xor (layer6_outputs(4355));
    layer7_outputs(832) <= layer6_outputs(3938);
    layer7_outputs(833) <= not(layer6_outputs(3039));
    layer7_outputs(834) <= not(layer6_outputs(381));
    layer7_outputs(835) <= not(layer6_outputs(3230));
    layer7_outputs(836) <= not(layer6_outputs(2065));
    layer7_outputs(837) <= layer6_outputs(4610);
    layer7_outputs(838) <= layer6_outputs(2422);
    layer7_outputs(839) <= layer6_outputs(732);
    layer7_outputs(840) <= not((layer6_outputs(1235)) or (layer6_outputs(4523)));
    layer7_outputs(841) <= (layer6_outputs(1994)) and (layer6_outputs(3052));
    layer7_outputs(842) <= not((layer6_outputs(2868)) xor (layer6_outputs(1051)));
    layer7_outputs(843) <= layer6_outputs(36);
    layer7_outputs(844) <= not(layer6_outputs(5007));
    layer7_outputs(845) <= not(layer6_outputs(4090)) or (layer6_outputs(917));
    layer7_outputs(846) <= (layer6_outputs(150)) xor (layer6_outputs(3934));
    layer7_outputs(847) <= (layer6_outputs(205)) or (layer6_outputs(108));
    layer7_outputs(848) <= not((layer6_outputs(2081)) and (layer6_outputs(86)));
    layer7_outputs(849) <= not(layer6_outputs(3162));
    layer7_outputs(850) <= layer6_outputs(3453);
    layer7_outputs(851) <= not(layer6_outputs(4588));
    layer7_outputs(852) <= not(layer6_outputs(3506));
    layer7_outputs(853) <= not((layer6_outputs(3195)) and (layer6_outputs(4163)));
    layer7_outputs(854) <= (layer6_outputs(4893)) xor (layer6_outputs(660));
    layer7_outputs(855) <= '1';
    layer7_outputs(856) <= not(layer6_outputs(4812));
    layer7_outputs(857) <= (layer6_outputs(2904)) and not (layer6_outputs(4414));
    layer7_outputs(858) <= (layer6_outputs(235)) and not (layer6_outputs(3611));
    layer7_outputs(859) <= layer6_outputs(2182);
    layer7_outputs(860) <= not(layer6_outputs(4444));
    layer7_outputs(861) <= not(layer6_outputs(2502));
    layer7_outputs(862) <= layer6_outputs(1738);
    layer7_outputs(863) <= not(layer6_outputs(3700));
    layer7_outputs(864) <= not(layer6_outputs(989));
    layer7_outputs(865) <= layer6_outputs(3410);
    layer7_outputs(866) <= not(layer6_outputs(3648)) or (layer6_outputs(3247));
    layer7_outputs(867) <= (layer6_outputs(3065)) and (layer6_outputs(2058));
    layer7_outputs(868) <= not(layer6_outputs(2400));
    layer7_outputs(869) <= not((layer6_outputs(1581)) xor (layer6_outputs(1161)));
    layer7_outputs(870) <= not(layer6_outputs(2029)) or (layer6_outputs(3683));
    layer7_outputs(871) <= not(layer6_outputs(405));
    layer7_outputs(872) <= (layer6_outputs(5083)) or (layer6_outputs(4804));
    layer7_outputs(873) <= layer6_outputs(3040);
    layer7_outputs(874) <= layer6_outputs(2174);
    layer7_outputs(875) <= not(layer6_outputs(3969));
    layer7_outputs(876) <= (layer6_outputs(1541)) xor (layer6_outputs(5101));
    layer7_outputs(877) <= not((layer6_outputs(4058)) or (layer6_outputs(3220)));
    layer7_outputs(878) <= not((layer6_outputs(4771)) and (layer6_outputs(3856)));
    layer7_outputs(879) <= '1';
    layer7_outputs(880) <= not(layer6_outputs(2135));
    layer7_outputs(881) <= (layer6_outputs(3433)) and not (layer6_outputs(1304));
    layer7_outputs(882) <= not(layer6_outputs(645));
    layer7_outputs(883) <= layer6_outputs(112);
    layer7_outputs(884) <= not(layer6_outputs(2293)) or (layer6_outputs(4922));
    layer7_outputs(885) <= not(layer6_outputs(2675));
    layer7_outputs(886) <= not(layer6_outputs(3861)) or (layer6_outputs(629));
    layer7_outputs(887) <= layer6_outputs(92);
    layer7_outputs(888) <= layer6_outputs(1583);
    layer7_outputs(889) <= (layer6_outputs(2690)) and not (layer6_outputs(2684));
    layer7_outputs(890) <= not((layer6_outputs(3599)) and (layer6_outputs(74)));
    layer7_outputs(891) <= not(layer6_outputs(599));
    layer7_outputs(892) <= not((layer6_outputs(4320)) and (layer6_outputs(4012)));
    layer7_outputs(893) <= not(layer6_outputs(1945));
    layer7_outputs(894) <= not((layer6_outputs(331)) and (layer6_outputs(3589)));
    layer7_outputs(895) <= (layer6_outputs(4497)) and not (layer6_outputs(2818));
    layer7_outputs(896) <= layer6_outputs(794);
    layer7_outputs(897) <= layer6_outputs(4125);
    layer7_outputs(898) <= layer6_outputs(745);
    layer7_outputs(899) <= layer6_outputs(5054);
    layer7_outputs(900) <= not(layer6_outputs(490));
    layer7_outputs(901) <= layer6_outputs(2530);
    layer7_outputs(902) <= (layer6_outputs(5024)) xor (layer6_outputs(2543));
    layer7_outputs(903) <= layer6_outputs(3518);
    layer7_outputs(904) <= not((layer6_outputs(1273)) or (layer6_outputs(4096)));
    layer7_outputs(905) <= (layer6_outputs(2998)) and not (layer6_outputs(2593));
    layer7_outputs(906) <= not(layer6_outputs(3967));
    layer7_outputs(907) <= layer6_outputs(4646);
    layer7_outputs(908) <= not(layer6_outputs(622)) or (layer6_outputs(823));
    layer7_outputs(909) <= layer6_outputs(56);
    layer7_outputs(910) <= layer6_outputs(1649);
    layer7_outputs(911) <= (layer6_outputs(2624)) xor (layer6_outputs(535));
    layer7_outputs(912) <= not((layer6_outputs(4832)) and (layer6_outputs(2853)));
    layer7_outputs(913) <= not(layer6_outputs(272));
    layer7_outputs(914) <= not(layer6_outputs(2454));
    layer7_outputs(915) <= layer6_outputs(3792);
    layer7_outputs(916) <= layer6_outputs(1685);
    layer7_outputs(917) <= not((layer6_outputs(971)) xor (layer6_outputs(3835)));
    layer7_outputs(918) <= layer6_outputs(3512);
    layer7_outputs(919) <= layer6_outputs(2682);
    layer7_outputs(920) <= layer6_outputs(2540);
    layer7_outputs(921) <= (layer6_outputs(4617)) or (layer6_outputs(1342));
    layer7_outputs(922) <= layer6_outputs(1544);
    layer7_outputs(923) <= not(layer6_outputs(1775));
    layer7_outputs(924) <= not((layer6_outputs(1963)) xor (layer6_outputs(2175)));
    layer7_outputs(925) <= not(layer6_outputs(980)) or (layer6_outputs(1139));
    layer7_outputs(926) <= layer6_outputs(770);
    layer7_outputs(927) <= not(layer6_outputs(1388));
    layer7_outputs(928) <= layer6_outputs(1229);
    layer7_outputs(929) <= '0';
    layer7_outputs(930) <= layer6_outputs(986);
    layer7_outputs(931) <= (layer6_outputs(2294)) xor (layer6_outputs(3920));
    layer7_outputs(932) <= (layer6_outputs(4977)) xor (layer6_outputs(4533));
    layer7_outputs(933) <= not(layer6_outputs(2702));
    layer7_outputs(934) <= not((layer6_outputs(4855)) or (layer6_outputs(3433)));
    layer7_outputs(935) <= (layer6_outputs(4112)) and not (layer6_outputs(2372));
    layer7_outputs(936) <= not((layer6_outputs(3146)) or (layer6_outputs(244)));
    layer7_outputs(937) <= layer6_outputs(1431);
    layer7_outputs(938) <= layer6_outputs(3668);
    layer7_outputs(939) <= not((layer6_outputs(3376)) or (layer6_outputs(4094)));
    layer7_outputs(940) <= layer6_outputs(5051);
    layer7_outputs(941) <= (layer6_outputs(3053)) and not (layer6_outputs(4658));
    layer7_outputs(942) <= layer6_outputs(4904);
    layer7_outputs(943) <= (layer6_outputs(586)) and not (layer6_outputs(4973));
    layer7_outputs(944) <= layer6_outputs(1385);
    layer7_outputs(945) <= layer6_outputs(3865);
    layer7_outputs(946) <= layer6_outputs(1557);
    layer7_outputs(947) <= not((layer6_outputs(2761)) or (layer6_outputs(854)));
    layer7_outputs(948) <= not(layer6_outputs(2546));
    layer7_outputs(949) <= '1';
    layer7_outputs(950) <= layer6_outputs(829);
    layer7_outputs(951) <= not(layer6_outputs(2383));
    layer7_outputs(952) <= not(layer6_outputs(3513));
    layer7_outputs(953) <= '1';
    layer7_outputs(954) <= layer6_outputs(1332);
    layer7_outputs(955) <= (layer6_outputs(1297)) xor (layer6_outputs(2411));
    layer7_outputs(956) <= not(layer6_outputs(4323));
    layer7_outputs(957) <= not((layer6_outputs(3606)) or (layer6_outputs(2421)));
    layer7_outputs(958) <= (layer6_outputs(1754)) xor (layer6_outputs(3533));
    layer7_outputs(959) <= not((layer6_outputs(1457)) xor (layer6_outputs(548)));
    layer7_outputs(960) <= '1';
    layer7_outputs(961) <= (layer6_outputs(4277)) xor (layer6_outputs(3966));
    layer7_outputs(962) <= (layer6_outputs(3017)) and not (layer6_outputs(2959));
    layer7_outputs(963) <= not((layer6_outputs(618)) xor (layer6_outputs(3565)));
    layer7_outputs(964) <= layer6_outputs(711);
    layer7_outputs(965) <= not(layer6_outputs(2432));
    layer7_outputs(966) <= layer6_outputs(4529);
    layer7_outputs(967) <= not((layer6_outputs(402)) or (layer6_outputs(259)));
    layer7_outputs(968) <= not(layer6_outputs(4498));
    layer7_outputs(969) <= not(layer6_outputs(677));
    layer7_outputs(970) <= not(layer6_outputs(3830)) or (layer6_outputs(3905));
    layer7_outputs(971) <= not(layer6_outputs(3983)) or (layer6_outputs(2181));
    layer7_outputs(972) <= not(layer6_outputs(1352));
    layer7_outputs(973) <= (layer6_outputs(4550)) and not (layer6_outputs(827));
    layer7_outputs(974) <= layer6_outputs(4256);
    layer7_outputs(975) <= (layer6_outputs(3946)) and not (layer6_outputs(1022));
    layer7_outputs(976) <= layer6_outputs(502);
    layer7_outputs(977) <= not(layer6_outputs(4478));
    layer7_outputs(978) <= not(layer6_outputs(2237)) or (layer6_outputs(2194));
    layer7_outputs(979) <= (layer6_outputs(343)) and not (layer6_outputs(1657));
    layer7_outputs(980) <= not(layer6_outputs(1639)) or (layer6_outputs(166));
    layer7_outputs(981) <= '1';
    layer7_outputs(982) <= (layer6_outputs(3382)) and (layer6_outputs(1564));
    layer7_outputs(983) <= (layer6_outputs(2599)) and not (layer6_outputs(2542));
    layer7_outputs(984) <= not(layer6_outputs(4420));
    layer7_outputs(985) <= not((layer6_outputs(3661)) and (layer6_outputs(4449)));
    layer7_outputs(986) <= '1';
    layer7_outputs(987) <= not(layer6_outputs(4904));
    layer7_outputs(988) <= (layer6_outputs(458)) and not (layer6_outputs(4286));
    layer7_outputs(989) <= (layer6_outputs(1479)) and not (layer6_outputs(2285));
    layer7_outputs(990) <= not(layer6_outputs(4958)) or (layer6_outputs(311));
    layer7_outputs(991) <= (layer6_outputs(268)) or (layer6_outputs(4221));
    layer7_outputs(992) <= not(layer6_outputs(1416));
    layer7_outputs(993) <= not(layer6_outputs(4086));
    layer7_outputs(994) <= layer6_outputs(2664);
    layer7_outputs(995) <= not(layer6_outputs(3799));
    layer7_outputs(996) <= '1';
    layer7_outputs(997) <= not(layer6_outputs(3881));
    layer7_outputs(998) <= layer6_outputs(3564);
    layer7_outputs(999) <= not(layer6_outputs(580));
    layer7_outputs(1000) <= '0';
    layer7_outputs(1001) <= (layer6_outputs(539)) xor (layer6_outputs(1282));
    layer7_outputs(1002) <= not(layer6_outputs(1398));
    layer7_outputs(1003) <= not((layer6_outputs(23)) and (layer6_outputs(1656)));
    layer7_outputs(1004) <= layer6_outputs(3800);
    layer7_outputs(1005) <= layer6_outputs(3198);
    layer7_outputs(1006) <= (layer6_outputs(5040)) and not (layer6_outputs(2987));
    layer7_outputs(1007) <= layer6_outputs(835);
    layer7_outputs(1008) <= not(layer6_outputs(1513));
    layer7_outputs(1009) <= (layer6_outputs(107)) xor (layer6_outputs(4213));
    layer7_outputs(1010) <= layer6_outputs(1954);
    layer7_outputs(1011) <= (layer6_outputs(797)) and not (layer6_outputs(165));
    layer7_outputs(1012) <= layer6_outputs(1222);
    layer7_outputs(1013) <= (layer6_outputs(665)) xor (layer6_outputs(4913));
    layer7_outputs(1014) <= not(layer6_outputs(3827));
    layer7_outputs(1015) <= not(layer6_outputs(5013));
    layer7_outputs(1016) <= not((layer6_outputs(4856)) xor (layer6_outputs(544)));
    layer7_outputs(1017) <= not(layer6_outputs(556));
    layer7_outputs(1018) <= not(layer6_outputs(2371)) or (layer6_outputs(2658));
    layer7_outputs(1019) <= not((layer6_outputs(1341)) xor (layer6_outputs(1158)));
    layer7_outputs(1020) <= not((layer6_outputs(21)) or (layer6_outputs(3125)));
    layer7_outputs(1021) <= layer6_outputs(3351);
    layer7_outputs(1022) <= not(layer6_outputs(984));
    layer7_outputs(1023) <= not((layer6_outputs(1467)) xor (layer6_outputs(2933)));
    layer7_outputs(1024) <= not((layer6_outputs(3552)) or (layer6_outputs(3780)));
    layer7_outputs(1025) <= '0';
    layer7_outputs(1026) <= layer6_outputs(4404);
    layer7_outputs(1027) <= not(layer6_outputs(751));
    layer7_outputs(1028) <= (layer6_outputs(2354)) xor (layer6_outputs(3722));
    layer7_outputs(1029) <= (layer6_outputs(3705)) and (layer6_outputs(389));
    layer7_outputs(1030) <= layer6_outputs(1609);
    layer7_outputs(1031) <= (layer6_outputs(3388)) and not (layer6_outputs(5070));
    layer7_outputs(1032) <= layer6_outputs(3855);
    layer7_outputs(1033) <= not(layer6_outputs(1076)) or (layer6_outputs(508));
    layer7_outputs(1034) <= not((layer6_outputs(4246)) xor (layer6_outputs(3756)));
    layer7_outputs(1035) <= layer6_outputs(490);
    layer7_outputs(1036) <= layer6_outputs(4003);
    layer7_outputs(1037) <= (layer6_outputs(128)) and not (layer6_outputs(4188));
    layer7_outputs(1038) <= (layer6_outputs(47)) and not (layer6_outputs(3009));
    layer7_outputs(1039) <= layer6_outputs(1856);
    layer7_outputs(1040) <= not(layer6_outputs(2639));
    layer7_outputs(1041) <= layer6_outputs(1299);
    layer7_outputs(1042) <= not((layer6_outputs(616)) and (layer6_outputs(1945)));
    layer7_outputs(1043) <= not((layer6_outputs(3553)) xor (layer6_outputs(2415)));
    layer7_outputs(1044) <= layer6_outputs(686);
    layer7_outputs(1045) <= not(layer6_outputs(4781));
    layer7_outputs(1046) <= not((layer6_outputs(440)) or (layer6_outputs(3507)));
    layer7_outputs(1047) <= (layer6_outputs(2397)) and not (layer6_outputs(4136));
    layer7_outputs(1048) <= layer6_outputs(3858);
    layer7_outputs(1049) <= not((layer6_outputs(1612)) and (layer6_outputs(3805)));
    layer7_outputs(1050) <= not(layer6_outputs(4596));
    layer7_outputs(1051) <= not(layer6_outputs(1117));
    layer7_outputs(1052) <= not((layer6_outputs(1838)) and (layer6_outputs(298)));
    layer7_outputs(1053) <= not(layer6_outputs(4343));
    layer7_outputs(1054) <= not(layer6_outputs(1234));
    layer7_outputs(1055) <= not(layer6_outputs(4072));
    layer7_outputs(1056) <= not(layer6_outputs(4248));
    layer7_outputs(1057) <= (layer6_outputs(361)) and not (layer6_outputs(2393));
    layer7_outputs(1058) <= not(layer6_outputs(1009));
    layer7_outputs(1059) <= not((layer6_outputs(2742)) and (layer6_outputs(2881)));
    layer7_outputs(1060) <= (layer6_outputs(2462)) xor (layer6_outputs(1563));
    layer7_outputs(1061) <= layer6_outputs(4695);
    layer7_outputs(1062) <= not(layer6_outputs(1952)) or (layer6_outputs(2946));
    layer7_outputs(1063) <= not((layer6_outputs(252)) or (layer6_outputs(4995)));
    layer7_outputs(1064) <= (layer6_outputs(4704)) and (layer6_outputs(2792));
    layer7_outputs(1065) <= not(layer6_outputs(1778)) or (layer6_outputs(520));
    layer7_outputs(1066) <= not(layer6_outputs(2222));
    layer7_outputs(1067) <= not((layer6_outputs(4839)) and (layer6_outputs(1749)));
    layer7_outputs(1068) <= not(layer6_outputs(3143));
    layer7_outputs(1069) <= layer6_outputs(1276);
    layer7_outputs(1070) <= not(layer6_outputs(3388));
    layer7_outputs(1071) <= not(layer6_outputs(3056));
    layer7_outputs(1072) <= (layer6_outputs(1695)) and not (layer6_outputs(4680));
    layer7_outputs(1073) <= (layer6_outputs(3413)) or (layer6_outputs(2575));
    layer7_outputs(1074) <= not(layer6_outputs(4592));
    layer7_outputs(1075) <= not((layer6_outputs(5012)) xor (layer6_outputs(694)));
    layer7_outputs(1076) <= layer6_outputs(4169);
    layer7_outputs(1077) <= layer6_outputs(1933);
    layer7_outputs(1078) <= not((layer6_outputs(1725)) xor (layer6_outputs(3110)));
    layer7_outputs(1079) <= layer6_outputs(1687);
    layer7_outputs(1080) <= not(layer6_outputs(1244));
    layer7_outputs(1081) <= (layer6_outputs(4440)) xor (layer6_outputs(439));
    layer7_outputs(1082) <= layer6_outputs(1200);
    layer7_outputs(1083) <= (layer6_outputs(3071)) and not (layer6_outputs(4805));
    layer7_outputs(1084) <= not(layer6_outputs(1124));
    layer7_outputs(1085) <= (layer6_outputs(1237)) xor (layer6_outputs(266));
    layer7_outputs(1086) <= (layer6_outputs(479)) and (layer6_outputs(2085));
    layer7_outputs(1087) <= not(layer6_outputs(2802));
    layer7_outputs(1088) <= layer6_outputs(5104);
    layer7_outputs(1089) <= layer6_outputs(1673);
    layer7_outputs(1090) <= (layer6_outputs(4307)) or (layer6_outputs(981));
    layer7_outputs(1091) <= layer6_outputs(1185);
    layer7_outputs(1092) <= (layer6_outputs(3318)) and not (layer6_outputs(2365));
    layer7_outputs(1093) <= not(layer6_outputs(4262));
    layer7_outputs(1094) <= not((layer6_outputs(4743)) xor (layer6_outputs(4271)));
    layer7_outputs(1095) <= not(layer6_outputs(1682));
    layer7_outputs(1096) <= not(layer6_outputs(3760));
    layer7_outputs(1097) <= not((layer6_outputs(982)) xor (layer6_outputs(4573)));
    layer7_outputs(1098) <= (layer6_outputs(1739)) and (layer6_outputs(3563));
    layer7_outputs(1099) <= not(layer6_outputs(4784));
    layer7_outputs(1100) <= layer6_outputs(3558);
    layer7_outputs(1101) <= (layer6_outputs(3257)) xor (layer6_outputs(2653));
    layer7_outputs(1102) <= layer6_outputs(4543);
    layer7_outputs(1103) <= layer6_outputs(3414);
    layer7_outputs(1104) <= not(layer6_outputs(4102));
    layer7_outputs(1105) <= not(layer6_outputs(1042));
    layer7_outputs(1106) <= layer6_outputs(5099);
    layer7_outputs(1107) <= not(layer6_outputs(3478));
    layer7_outputs(1108) <= '0';
    layer7_outputs(1109) <= (layer6_outputs(4305)) and not (layer6_outputs(2402));
    layer7_outputs(1110) <= (layer6_outputs(2880)) or (layer6_outputs(4647));
    layer7_outputs(1111) <= not(layer6_outputs(2473));
    layer7_outputs(1112) <= not((layer6_outputs(156)) or (layer6_outputs(718)));
    layer7_outputs(1113) <= not((layer6_outputs(3146)) xor (layer6_outputs(4282)));
    layer7_outputs(1114) <= not(layer6_outputs(2265));
    layer7_outputs(1115) <= layer6_outputs(4329);
    layer7_outputs(1116) <= not(layer6_outputs(4413)) or (layer6_outputs(2787));
    layer7_outputs(1117) <= (layer6_outputs(2643)) xor (layer6_outputs(951));
    layer7_outputs(1118) <= (layer6_outputs(3527)) and (layer6_outputs(4859));
    layer7_outputs(1119) <= layer6_outputs(1096);
    layer7_outputs(1120) <= not(layer6_outputs(3345)) or (layer6_outputs(1492));
    layer7_outputs(1121) <= (layer6_outputs(4379)) xor (layer6_outputs(3790));
    layer7_outputs(1122) <= layer6_outputs(4335);
    layer7_outputs(1123) <= layer6_outputs(704);
    layer7_outputs(1124) <= not(layer6_outputs(4016));
    layer7_outputs(1125) <= not((layer6_outputs(4298)) and (layer6_outputs(3656)));
    layer7_outputs(1126) <= (layer6_outputs(62)) xor (layer6_outputs(3435));
    layer7_outputs(1127) <= not(layer6_outputs(3497));
    layer7_outputs(1128) <= layer6_outputs(3210);
    layer7_outputs(1129) <= not(layer6_outputs(2802));
    layer7_outputs(1130) <= not(layer6_outputs(49));
    layer7_outputs(1131) <= not((layer6_outputs(3765)) xor (layer6_outputs(4383)));
    layer7_outputs(1132) <= not((layer6_outputs(499)) and (layer6_outputs(1006)));
    layer7_outputs(1133) <= not((layer6_outputs(3246)) xor (layer6_outputs(4198)));
    layer7_outputs(1134) <= layer6_outputs(3579);
    layer7_outputs(1135) <= not(layer6_outputs(2661));
    layer7_outputs(1136) <= not(layer6_outputs(101)) or (layer6_outputs(2647));
    layer7_outputs(1137) <= not((layer6_outputs(2889)) xor (layer6_outputs(100)));
    layer7_outputs(1138) <= not((layer6_outputs(2121)) and (layer6_outputs(4293)));
    layer7_outputs(1139) <= '1';
    layer7_outputs(1140) <= not(layer6_outputs(3758)) or (layer6_outputs(4342));
    layer7_outputs(1141) <= not(layer6_outputs(775));
    layer7_outputs(1142) <= (layer6_outputs(2613)) and not (layer6_outputs(2302));
    layer7_outputs(1143) <= (layer6_outputs(4726)) xor (layer6_outputs(3592));
    layer7_outputs(1144) <= not(layer6_outputs(935));
    layer7_outputs(1145) <= (layer6_outputs(4177)) and not (layer6_outputs(2207));
    layer7_outputs(1146) <= not((layer6_outputs(3730)) xor (layer6_outputs(2834)));
    layer7_outputs(1147) <= not(layer6_outputs(2365));
    layer7_outputs(1148) <= layer6_outputs(2335);
    layer7_outputs(1149) <= (layer6_outputs(4339)) xor (layer6_outputs(1712));
    layer7_outputs(1150) <= (layer6_outputs(1062)) and not (layer6_outputs(2428));
    layer7_outputs(1151) <= (layer6_outputs(1475)) xor (layer6_outputs(226));
    layer7_outputs(1152) <= (layer6_outputs(350)) xor (layer6_outputs(111));
    layer7_outputs(1153) <= layer6_outputs(1074);
    layer7_outputs(1154) <= not((layer6_outputs(3019)) and (layer6_outputs(2865)));
    layer7_outputs(1155) <= (layer6_outputs(1196)) xor (layer6_outputs(1133));
    layer7_outputs(1156) <= not(layer6_outputs(640));
    layer7_outputs(1157) <= not(layer6_outputs(2896));
    layer7_outputs(1158) <= not((layer6_outputs(1716)) xor (layer6_outputs(1941)));
    layer7_outputs(1159) <= not(layer6_outputs(3173));
    layer7_outputs(1160) <= layer6_outputs(2254);
    layer7_outputs(1161) <= (layer6_outputs(2381)) and not (layer6_outputs(2745));
    layer7_outputs(1162) <= not(layer6_outputs(4852));
    layer7_outputs(1163) <= not(layer6_outputs(2245));
    layer7_outputs(1164) <= not(layer6_outputs(927));
    layer7_outputs(1165) <= layer6_outputs(1358);
    layer7_outputs(1166) <= not(layer6_outputs(2627));
    layer7_outputs(1167) <= not((layer6_outputs(4164)) xor (layer6_outputs(4418)));
    layer7_outputs(1168) <= (layer6_outputs(3051)) and not (layer6_outputs(4932));
    layer7_outputs(1169) <= not((layer6_outputs(2048)) or (layer6_outputs(2478)));
    layer7_outputs(1170) <= (layer6_outputs(4217)) or (layer6_outputs(4239));
    layer7_outputs(1171) <= not(layer6_outputs(3597)) or (layer6_outputs(4187));
    layer7_outputs(1172) <= not(layer6_outputs(1596));
    layer7_outputs(1173) <= not((layer6_outputs(3426)) xor (layer6_outputs(1663)));
    layer7_outputs(1174) <= not(layer6_outputs(824));
    layer7_outputs(1175) <= (layer6_outputs(2936)) and (layer6_outputs(202));
    layer7_outputs(1176) <= not(layer6_outputs(532));
    layer7_outputs(1177) <= layer6_outputs(4385);
    layer7_outputs(1178) <= (layer6_outputs(3305)) xor (layer6_outputs(2265));
    layer7_outputs(1179) <= not((layer6_outputs(482)) or (layer6_outputs(2724)));
    layer7_outputs(1180) <= not(layer6_outputs(5017));
    layer7_outputs(1181) <= layer6_outputs(305);
    layer7_outputs(1182) <= not((layer6_outputs(3462)) or (layer6_outputs(2317)));
    layer7_outputs(1183) <= layer6_outputs(2519);
    layer7_outputs(1184) <= layer6_outputs(3753);
    layer7_outputs(1185) <= not(layer6_outputs(4263)) or (layer6_outputs(4638));
    layer7_outputs(1186) <= (layer6_outputs(2877)) and (layer6_outputs(1199));
    layer7_outputs(1187) <= '0';
    layer7_outputs(1188) <= not(layer6_outputs(2619));
    layer7_outputs(1189) <= not((layer6_outputs(4564)) xor (layer6_outputs(2654)));
    layer7_outputs(1190) <= (layer6_outputs(688)) xor (layer6_outputs(3222));
    layer7_outputs(1191) <= '0';
    layer7_outputs(1192) <= not(layer6_outputs(1706));
    layer7_outputs(1193) <= not(layer6_outputs(89));
    layer7_outputs(1194) <= (layer6_outputs(1760)) and not (layer6_outputs(3231));
    layer7_outputs(1195) <= layer6_outputs(1790);
    layer7_outputs(1196) <= not((layer6_outputs(676)) and (layer6_outputs(142)));
    layer7_outputs(1197) <= (layer6_outputs(2782)) and not (layer6_outputs(4948));
    layer7_outputs(1198) <= not(layer6_outputs(2632));
    layer7_outputs(1199) <= not((layer6_outputs(3689)) and (layer6_outputs(4118)));
    layer7_outputs(1200) <= not((layer6_outputs(3448)) xor (layer6_outputs(2927)));
    layer7_outputs(1201) <= layer6_outputs(4214);
    layer7_outputs(1202) <= not(layer6_outputs(1524)) or (layer6_outputs(1367));
    layer7_outputs(1203) <= (layer6_outputs(1995)) and (layer6_outputs(3179));
    layer7_outputs(1204) <= not(layer6_outputs(691));
    layer7_outputs(1205) <= not(layer6_outputs(3386));
    layer7_outputs(1206) <= not(layer6_outputs(4585));
    layer7_outputs(1207) <= (layer6_outputs(1452)) and (layer6_outputs(3460));
    layer7_outputs(1208) <= layer6_outputs(651);
    layer7_outputs(1209) <= not(layer6_outputs(2333));
    layer7_outputs(1210) <= '0';
    layer7_outputs(1211) <= not(layer6_outputs(4654));
    layer7_outputs(1212) <= layer6_outputs(3803);
    layer7_outputs(1213) <= layer6_outputs(1636);
    layer7_outputs(1214) <= not(layer6_outputs(1287)) or (layer6_outputs(224));
    layer7_outputs(1215) <= (layer6_outputs(993)) xor (layer6_outputs(2099));
    layer7_outputs(1216) <= not(layer6_outputs(2212));
    layer7_outputs(1217) <= not(layer6_outputs(4594));
    layer7_outputs(1218) <= not(layer6_outputs(1105));
    layer7_outputs(1219) <= layer6_outputs(1892);
    layer7_outputs(1220) <= not(layer6_outputs(2300));
    layer7_outputs(1221) <= layer6_outputs(3105);
    layer7_outputs(1222) <= (layer6_outputs(3094)) and not (layer6_outputs(2663));
    layer7_outputs(1223) <= layer6_outputs(2926);
    layer7_outputs(1224) <= not((layer6_outputs(3921)) and (layer6_outputs(2662)));
    layer7_outputs(1225) <= not(layer6_outputs(3564));
    layer7_outputs(1226) <= not(layer6_outputs(2552)) or (layer6_outputs(3687));
    layer7_outputs(1227) <= not(layer6_outputs(2441)) or (layer6_outputs(1170));
    layer7_outputs(1228) <= not((layer6_outputs(3123)) or (layer6_outputs(959)));
    layer7_outputs(1229) <= not(layer6_outputs(4337));
    layer7_outputs(1230) <= not(layer6_outputs(1575));
    layer7_outputs(1231) <= layer6_outputs(4608);
    layer7_outputs(1232) <= not((layer6_outputs(5014)) or (layer6_outputs(1735)));
    layer7_outputs(1233) <= layer6_outputs(389);
    layer7_outputs(1234) <= layer6_outputs(1053);
    layer7_outputs(1235) <= not(layer6_outputs(2032));
    layer7_outputs(1236) <= not(layer6_outputs(3113)) or (layer6_outputs(3983));
    layer7_outputs(1237) <= (layer6_outputs(3878)) xor (layer6_outputs(4165));
    layer7_outputs(1238) <= not(layer6_outputs(2172)) or (layer6_outputs(4235));
    layer7_outputs(1239) <= not((layer6_outputs(1927)) and (layer6_outputs(3812)));
    layer7_outputs(1240) <= not((layer6_outputs(2678)) or (layer6_outputs(73)));
    layer7_outputs(1241) <= (layer6_outputs(313)) xor (layer6_outputs(1280));
    layer7_outputs(1242) <= not(layer6_outputs(1619));
    layer7_outputs(1243) <= layer6_outputs(4117);
    layer7_outputs(1244) <= not(layer6_outputs(4502));
    layer7_outputs(1245) <= layer6_outputs(506);
    layer7_outputs(1246) <= not(layer6_outputs(550));
    layer7_outputs(1247) <= layer6_outputs(3226);
    layer7_outputs(1248) <= (layer6_outputs(3757)) and not (layer6_outputs(4631));
    layer7_outputs(1249) <= not(layer6_outputs(1623)) or (layer6_outputs(1892));
    layer7_outputs(1250) <= not(layer6_outputs(1310));
    layer7_outputs(1251) <= layer6_outputs(1793);
    layer7_outputs(1252) <= layer6_outputs(763);
    layer7_outputs(1253) <= layer6_outputs(1230);
    layer7_outputs(1254) <= not(layer6_outputs(4285));
    layer7_outputs(1255) <= (layer6_outputs(5055)) and not (layer6_outputs(90));
    layer7_outputs(1256) <= not(layer6_outputs(2462));
    layer7_outputs(1257) <= not((layer6_outputs(2815)) or (layer6_outputs(3438)));
    layer7_outputs(1258) <= not(layer6_outputs(302));
    layer7_outputs(1259) <= (layer6_outputs(1846)) and not (layer6_outputs(4395));
    layer7_outputs(1260) <= not(layer6_outputs(1916)) or (layer6_outputs(2828));
    layer7_outputs(1261) <= (layer6_outputs(3327)) xor (layer6_outputs(4070));
    layer7_outputs(1262) <= (layer6_outputs(4587)) and not (layer6_outputs(1116));
    layer7_outputs(1263) <= '1';
    layer7_outputs(1264) <= not(layer6_outputs(1982));
    layer7_outputs(1265) <= layer6_outputs(57);
    layer7_outputs(1266) <= not(layer6_outputs(4780)) or (layer6_outputs(2829));
    layer7_outputs(1267) <= (layer6_outputs(2727)) or (layer6_outputs(4854));
    layer7_outputs(1268) <= not(layer6_outputs(1046));
    layer7_outputs(1269) <= not(layer6_outputs(2651));
    layer7_outputs(1270) <= not(layer6_outputs(3744));
    layer7_outputs(1271) <= (layer6_outputs(4023)) and not (layer6_outputs(2565));
    layer7_outputs(1272) <= (layer6_outputs(2939)) and (layer6_outputs(4173));
    layer7_outputs(1273) <= (layer6_outputs(355)) and not (layer6_outputs(4099));
    layer7_outputs(1274) <= not(layer6_outputs(941));
    layer7_outputs(1275) <= not((layer6_outputs(1117)) xor (layer6_outputs(4426)));
    layer7_outputs(1276) <= layer6_outputs(4097);
    layer7_outputs(1277) <= layer6_outputs(4939);
    layer7_outputs(1278) <= not((layer6_outputs(4682)) or (layer6_outputs(359)));
    layer7_outputs(1279) <= not((layer6_outputs(5039)) xor (layer6_outputs(1253)));
    layer7_outputs(1280) <= not((layer6_outputs(4781)) xor (layer6_outputs(2375)));
    layer7_outputs(1281) <= not((layer6_outputs(5002)) xor (layer6_outputs(2164)));
    layer7_outputs(1282) <= layer6_outputs(2290);
    layer7_outputs(1283) <= not(layer6_outputs(4077)) or (layer6_outputs(1465));
    layer7_outputs(1284) <= not((layer6_outputs(4216)) xor (layer6_outputs(4274)));
    layer7_outputs(1285) <= layer6_outputs(1597);
    layer7_outputs(1286) <= (layer6_outputs(2719)) xor (layer6_outputs(2014));
    layer7_outputs(1287) <= not(layer6_outputs(3228));
    layer7_outputs(1288) <= (layer6_outputs(1691)) and (layer6_outputs(2977));
    layer7_outputs(1289) <= not((layer6_outputs(1891)) xor (layer6_outputs(848)));
    layer7_outputs(1290) <= not(layer6_outputs(1483)) or (layer6_outputs(1376));
    layer7_outputs(1291) <= (layer6_outputs(1747)) and not (layer6_outputs(4914));
    layer7_outputs(1292) <= (layer6_outputs(4034)) and (layer6_outputs(2765));
    layer7_outputs(1293) <= not(layer6_outputs(4983));
    layer7_outputs(1294) <= (layer6_outputs(352)) or (layer6_outputs(5062));
    layer7_outputs(1295) <= not(layer6_outputs(1871)) or (layer6_outputs(2386));
    layer7_outputs(1296) <= not((layer6_outputs(1366)) and (layer6_outputs(3739)));
    layer7_outputs(1297) <= layer6_outputs(3732);
    layer7_outputs(1298) <= not(layer6_outputs(953)) or (layer6_outputs(4892));
    layer7_outputs(1299) <= layer6_outputs(1445);
    layer7_outputs(1300) <= not(layer6_outputs(2094));
    layer7_outputs(1301) <= not(layer6_outputs(3651));
    layer7_outputs(1302) <= not(layer6_outputs(2404));
    layer7_outputs(1303) <= '0';
    layer7_outputs(1304) <= layer6_outputs(1323);
    layer7_outputs(1305) <= layer6_outputs(4768);
    layer7_outputs(1306) <= not((layer6_outputs(785)) xor (layer6_outputs(1097)));
    layer7_outputs(1307) <= layer6_outputs(4303);
    layer7_outputs(1308) <= layer6_outputs(2936);
    layer7_outputs(1309) <= not((layer6_outputs(261)) or (layer6_outputs(2520)));
    layer7_outputs(1310) <= layer6_outputs(4975);
    layer7_outputs(1311) <= layer6_outputs(120);
    layer7_outputs(1312) <= (layer6_outputs(1850)) xor (layer6_outputs(4232));
    layer7_outputs(1313) <= not(layer6_outputs(1740));
    layer7_outputs(1314) <= (layer6_outputs(1073)) and (layer6_outputs(3097));
    layer7_outputs(1315) <= (layer6_outputs(2190)) and not (layer6_outputs(3345));
    layer7_outputs(1316) <= not(layer6_outputs(4202)) or (layer6_outputs(513));
    layer7_outputs(1317) <= (layer6_outputs(1584)) and not (layer6_outputs(432));
    layer7_outputs(1318) <= layer6_outputs(3161);
    layer7_outputs(1319) <= not(layer6_outputs(2389));
    layer7_outputs(1320) <= not(layer6_outputs(1180)) or (layer6_outputs(512));
    layer7_outputs(1321) <= not((layer6_outputs(1130)) xor (layer6_outputs(2384)));
    layer7_outputs(1322) <= (layer6_outputs(4159)) or (layer6_outputs(5095));
    layer7_outputs(1323) <= not((layer6_outputs(3523)) xor (layer6_outputs(1411)));
    layer7_outputs(1324) <= not((layer6_outputs(3972)) xor (layer6_outputs(7)));
    layer7_outputs(1325) <= (layer6_outputs(1182)) xor (layer6_outputs(595));
    layer7_outputs(1326) <= not(layer6_outputs(1962)) or (layer6_outputs(728));
    layer7_outputs(1327) <= layer6_outputs(3640);
    layer7_outputs(1328) <= not(layer6_outputs(422));
    layer7_outputs(1329) <= not(layer6_outputs(2835));
    layer7_outputs(1330) <= not(layer6_outputs(1550));
    layer7_outputs(1331) <= '1';
    layer7_outputs(1332) <= not(layer6_outputs(3731));
    layer7_outputs(1333) <= not(layer6_outputs(55));
    layer7_outputs(1334) <= not((layer6_outputs(4309)) xor (layer6_outputs(2303)));
    layer7_outputs(1335) <= (layer6_outputs(4606)) or (layer6_outputs(1983));
    layer7_outputs(1336) <= not((layer6_outputs(903)) and (layer6_outputs(2638)));
    layer7_outputs(1337) <= (layer6_outputs(2831)) and not (layer6_outputs(3268));
    layer7_outputs(1338) <= (layer6_outputs(668)) xor (layer6_outputs(4138));
    layer7_outputs(1339) <= not(layer6_outputs(3863)) or (layer6_outputs(2747));
    layer7_outputs(1340) <= layer6_outputs(3858);
    layer7_outputs(1341) <= not(layer6_outputs(1318));
    layer7_outputs(1342) <= not(layer6_outputs(360));
    layer7_outputs(1343) <= layer6_outputs(4999);
    layer7_outputs(1344) <= not(layer6_outputs(760));
    layer7_outputs(1345) <= not(layer6_outputs(1162)) or (layer6_outputs(679));
    layer7_outputs(1346) <= layer6_outputs(4548);
    layer7_outputs(1347) <= (layer6_outputs(201)) and not (layer6_outputs(2753));
    layer7_outputs(1348) <= (layer6_outputs(2158)) xor (layer6_outputs(3647));
    layer7_outputs(1349) <= layer6_outputs(3267);
    layer7_outputs(1350) <= not(layer6_outputs(3560)) or (layer6_outputs(2708));
    layer7_outputs(1351) <= (layer6_outputs(4664)) and not (layer6_outputs(2055));
    layer7_outputs(1352) <= layer6_outputs(2874);
    layer7_outputs(1353) <= (layer6_outputs(2764)) or (layer6_outputs(2298));
    layer7_outputs(1354) <= not((layer6_outputs(281)) xor (layer6_outputs(4982)));
    layer7_outputs(1355) <= (layer6_outputs(3270)) and not (layer6_outputs(808));
    layer7_outputs(1356) <= not(layer6_outputs(3006));
    layer7_outputs(1357) <= not(layer6_outputs(193));
    layer7_outputs(1358) <= not((layer6_outputs(1980)) and (layer6_outputs(172)));
    layer7_outputs(1359) <= not(layer6_outputs(2768)) or (layer6_outputs(4723));
    layer7_outputs(1360) <= (layer6_outputs(3474)) and not (layer6_outputs(846));
    layer7_outputs(1361) <= not(layer6_outputs(1873));
    layer7_outputs(1362) <= (layer6_outputs(3841)) and not (layer6_outputs(1279));
    layer7_outputs(1363) <= layer6_outputs(1170);
    layer7_outputs(1364) <= not(layer6_outputs(636));
    layer7_outputs(1365) <= layer6_outputs(374);
    layer7_outputs(1366) <= not(layer6_outputs(5095));
    layer7_outputs(1367) <= layer6_outputs(4661);
    layer7_outputs(1368) <= not(layer6_outputs(1422)) or (layer6_outputs(351));
    layer7_outputs(1369) <= not(layer6_outputs(1999)) or (layer6_outputs(2385));
    layer7_outputs(1370) <= (layer6_outputs(2750)) xor (layer6_outputs(3723));
    layer7_outputs(1371) <= not((layer6_outputs(3563)) xor (layer6_outputs(1166)));
    layer7_outputs(1372) <= not((layer6_outputs(4140)) xor (layer6_outputs(992)));
    layer7_outputs(1373) <= layer6_outputs(755);
    layer7_outputs(1374) <= (layer6_outputs(4993)) and not (layer6_outputs(2825));
    layer7_outputs(1375) <= '0';
    layer7_outputs(1376) <= layer6_outputs(3063);
    layer7_outputs(1377) <= not((layer6_outputs(4624)) and (layer6_outputs(1647)));
    layer7_outputs(1378) <= not(layer6_outputs(3879));
    layer7_outputs(1379) <= not(layer6_outputs(4688));
    layer7_outputs(1380) <= not((layer6_outputs(476)) xor (layer6_outputs(5032)));
    layer7_outputs(1381) <= not(layer6_outputs(3944)) or (layer6_outputs(1256));
    layer7_outputs(1382) <= (layer6_outputs(2291)) xor (layer6_outputs(1817));
    layer7_outputs(1383) <= not(layer6_outputs(2794));
    layer7_outputs(1384) <= not(layer6_outputs(1680));
    layer7_outputs(1385) <= not(layer6_outputs(245));
    layer7_outputs(1386) <= layer6_outputs(1041);
    layer7_outputs(1387) <= not(layer6_outputs(2018)) or (layer6_outputs(632));
    layer7_outputs(1388) <= not((layer6_outputs(4259)) xor (layer6_outputs(3303)));
    layer7_outputs(1389) <= layer6_outputs(1005);
    layer7_outputs(1390) <= not(layer6_outputs(3233)) or (layer6_outputs(1965));
    layer7_outputs(1391) <= not(layer6_outputs(520));
    layer7_outputs(1392) <= not(layer6_outputs(4586));
    layer7_outputs(1393) <= not(layer6_outputs(4152)) or (layer6_outputs(3400));
    layer7_outputs(1394) <= not((layer6_outputs(3646)) or (layer6_outputs(1059)));
    layer7_outputs(1395) <= not(layer6_outputs(518));
    layer7_outputs(1396) <= layer6_outputs(82);
    layer7_outputs(1397) <= not((layer6_outputs(1445)) xor (layer6_outputs(2075)));
    layer7_outputs(1398) <= not(layer6_outputs(4672));
    layer7_outputs(1399) <= layer6_outputs(183);
    layer7_outputs(1400) <= not(layer6_outputs(3104));
    layer7_outputs(1401) <= not((layer6_outputs(1876)) xor (layer6_outputs(2577)));
    layer7_outputs(1402) <= not(layer6_outputs(90));
    layer7_outputs(1403) <= layer6_outputs(1494);
    layer7_outputs(1404) <= not(layer6_outputs(2673)) or (layer6_outputs(3576));
    layer7_outputs(1405) <= layer6_outputs(2749);
    layer7_outputs(1406) <= not((layer6_outputs(2470)) xor (layer6_outputs(1093)));
    layer7_outputs(1407) <= not(layer6_outputs(655));
    layer7_outputs(1408) <= (layer6_outputs(4123)) and not (layer6_outputs(2470));
    layer7_outputs(1409) <= not(layer6_outputs(1229));
    layer7_outputs(1410) <= not(layer6_outputs(3073)) or (layer6_outputs(338));
    layer7_outputs(1411) <= not((layer6_outputs(325)) xor (layer6_outputs(2165)));
    layer7_outputs(1412) <= not(layer6_outputs(4735));
    layer7_outputs(1413) <= not(layer6_outputs(4954)) or (layer6_outputs(4355));
    layer7_outputs(1414) <= not(layer6_outputs(3060));
    layer7_outputs(1415) <= (layer6_outputs(3439)) xor (layer6_outputs(663));
    layer7_outputs(1416) <= (layer6_outputs(779)) and not (layer6_outputs(780));
    layer7_outputs(1417) <= not((layer6_outputs(4920)) xor (layer6_outputs(1328)));
    layer7_outputs(1418) <= not((layer6_outputs(536)) xor (layer6_outputs(5027)));
    layer7_outputs(1419) <= not(layer6_outputs(433));
    layer7_outputs(1420) <= layer6_outputs(2131);
    layer7_outputs(1421) <= layer6_outputs(180);
    layer7_outputs(1422) <= not((layer6_outputs(1148)) xor (layer6_outputs(2420)));
    layer7_outputs(1423) <= not((layer6_outputs(2898)) xor (layer6_outputs(1084)));
    layer7_outputs(1424) <= layer6_outputs(1638);
    layer7_outputs(1425) <= not(layer6_outputs(1911)) or (layer6_outputs(3709));
    layer7_outputs(1426) <= (layer6_outputs(143)) xor (layer6_outputs(269));
    layer7_outputs(1427) <= not(layer6_outputs(1551));
    layer7_outputs(1428) <= not(layer6_outputs(3294));
    layer7_outputs(1429) <= (layer6_outputs(1066)) xor (layer6_outputs(1559));
    layer7_outputs(1430) <= layer6_outputs(1114);
    layer7_outputs(1431) <= (layer6_outputs(3733)) and not (layer6_outputs(2056));
    layer7_outputs(1432) <= (layer6_outputs(2614)) and (layer6_outputs(3422));
    layer7_outputs(1433) <= not(layer6_outputs(4015)) or (layer6_outputs(1800));
    layer7_outputs(1434) <= (layer6_outputs(1104)) and not (layer6_outputs(909));
    layer7_outputs(1435) <= layer6_outputs(1519);
    layer7_outputs(1436) <= layer6_outputs(4142);
    layer7_outputs(1437) <= not(layer6_outputs(2155));
    layer7_outputs(1438) <= layer6_outputs(935);
    layer7_outputs(1439) <= not(layer6_outputs(4860));
    layer7_outputs(1440) <= not((layer6_outputs(2073)) xor (layer6_outputs(3373)));
    layer7_outputs(1441) <= not((layer6_outputs(3836)) and (layer6_outputs(3235)));
    layer7_outputs(1442) <= not((layer6_outputs(1741)) xor (layer6_outputs(1176)));
    layer7_outputs(1443) <= layer6_outputs(897);
    layer7_outputs(1444) <= (layer6_outputs(649)) and not (layer6_outputs(1616));
    layer7_outputs(1445) <= (layer6_outputs(1833)) xor (layer6_outputs(706));
    layer7_outputs(1446) <= not(layer6_outputs(408));
    layer7_outputs(1447) <= layer6_outputs(3853);
    layer7_outputs(1448) <= not(layer6_outputs(4612));
    layer7_outputs(1449) <= not((layer6_outputs(372)) xor (layer6_outputs(3268)));
    layer7_outputs(1450) <= (layer6_outputs(239)) and (layer6_outputs(3641));
    layer7_outputs(1451) <= layer6_outputs(3363);
    layer7_outputs(1452) <= not(layer6_outputs(5049));
    layer7_outputs(1453) <= not(layer6_outputs(725));
    layer7_outputs(1454) <= layer6_outputs(2783);
    layer7_outputs(1455) <= layer6_outputs(202);
    layer7_outputs(1456) <= not(layer6_outputs(950)) or (layer6_outputs(2459));
    layer7_outputs(1457) <= not(layer6_outputs(4222));
    layer7_outputs(1458) <= not(layer6_outputs(45)) or (layer6_outputs(1980));
    layer7_outputs(1459) <= (layer6_outputs(1615)) or (layer6_outputs(1460));
    layer7_outputs(1460) <= (layer6_outputs(1645)) and not (layer6_outputs(4191));
    layer7_outputs(1461) <= (layer6_outputs(1341)) and not (layer6_outputs(4200));
    layer7_outputs(1462) <= (layer6_outputs(3129)) xor (layer6_outputs(3760));
    layer7_outputs(1463) <= layer6_outputs(2870);
    layer7_outputs(1464) <= not((layer6_outputs(1143)) and (layer6_outputs(1197)));
    layer7_outputs(1465) <= layer6_outputs(431);
    layer7_outputs(1466) <= not(layer6_outputs(3720)) or (layer6_outputs(2771));
    layer7_outputs(1467) <= not(layer6_outputs(4827));
    layer7_outputs(1468) <= not(layer6_outputs(1642));
    layer7_outputs(1469) <= not((layer6_outputs(2352)) xor (layer6_outputs(4034)));
    layer7_outputs(1470) <= not(layer6_outputs(5111));
    layer7_outputs(1471) <= not(layer6_outputs(3482));
    layer7_outputs(1472) <= (layer6_outputs(2553)) or (layer6_outputs(784));
    layer7_outputs(1473) <= not((layer6_outputs(639)) xor (layer6_outputs(1641)));
    layer7_outputs(1474) <= not((layer6_outputs(1501)) or (layer6_outputs(754)));
    layer7_outputs(1475) <= '1';
    layer7_outputs(1476) <= (layer6_outputs(4313)) and not (layer6_outputs(2739));
    layer7_outputs(1477) <= '1';
    layer7_outputs(1478) <= not(layer6_outputs(3060));
    layer7_outputs(1479) <= (layer6_outputs(3636)) and not (layer6_outputs(2154));
    layer7_outputs(1480) <= layer6_outputs(1471);
    layer7_outputs(1481) <= (layer6_outputs(2370)) and not (layer6_outputs(2959));
    layer7_outputs(1482) <= not((layer6_outputs(4373)) or (layer6_outputs(262)));
    layer7_outputs(1483) <= (layer6_outputs(4626)) and not (layer6_outputs(2408));
    layer7_outputs(1484) <= not(layer6_outputs(4908));
    layer7_outputs(1485) <= not((layer6_outputs(2823)) or (layer6_outputs(3754)));
    layer7_outputs(1486) <= not(layer6_outputs(3975));
    layer7_outputs(1487) <= not((layer6_outputs(254)) or (layer6_outputs(4480)));
    layer7_outputs(1488) <= not((layer6_outputs(1191)) or (layer6_outputs(4819)));
    layer7_outputs(1489) <= not(layer6_outputs(3443));
    layer7_outputs(1490) <= (layer6_outputs(2810)) xor (layer6_outputs(5047));
    layer7_outputs(1491) <= not(layer6_outputs(368));
    layer7_outputs(1492) <= not((layer6_outputs(4407)) or (layer6_outputs(895)));
    layer7_outputs(1493) <= not((layer6_outputs(3991)) and (layer6_outputs(1214)));
    layer7_outputs(1494) <= (layer6_outputs(554)) and (layer6_outputs(4949));
    layer7_outputs(1495) <= (layer6_outputs(4080)) xor (layer6_outputs(1996));
    layer7_outputs(1496) <= not(layer6_outputs(4637));
    layer7_outputs(1497) <= not(layer6_outputs(3028)) or (layer6_outputs(3871));
    layer7_outputs(1498) <= (layer6_outputs(4497)) xor (layer6_outputs(4501));
    layer7_outputs(1499) <= not(layer6_outputs(3036));
    layer7_outputs(1500) <= not(layer6_outputs(4652));
    layer7_outputs(1501) <= (layer6_outputs(3747)) and not (layer6_outputs(2602));
    layer7_outputs(1502) <= (layer6_outputs(1761)) xor (layer6_outputs(1326));
    layer7_outputs(1503) <= not((layer6_outputs(3975)) and (layer6_outputs(3671)));
    layer7_outputs(1504) <= not(layer6_outputs(4173));
    layer7_outputs(1505) <= (layer6_outputs(3608)) or (layer6_outputs(3005));
    layer7_outputs(1506) <= not(layer6_outputs(1296));
    layer7_outputs(1507) <= not(layer6_outputs(699));
    layer7_outputs(1508) <= layer6_outputs(719);
    layer7_outputs(1509) <= (layer6_outputs(4725)) or (layer6_outputs(478));
    layer7_outputs(1510) <= not(layer6_outputs(374));
    layer7_outputs(1511) <= not(layer6_outputs(2608));
    layer7_outputs(1512) <= layer6_outputs(1875);
    layer7_outputs(1513) <= not(layer6_outputs(1509));
    layer7_outputs(1514) <= not(layer6_outputs(1578));
    layer7_outputs(1515) <= layer6_outputs(3044);
    layer7_outputs(1516) <= layer6_outputs(3391);
    layer7_outputs(1517) <= (layer6_outputs(1409)) and (layer6_outputs(1138));
    layer7_outputs(1518) <= layer6_outputs(2504);
    layer7_outputs(1519) <= layer6_outputs(1486);
    layer7_outputs(1520) <= (layer6_outputs(2667)) and not (layer6_outputs(4569));
    layer7_outputs(1521) <= not(layer6_outputs(4114)) or (layer6_outputs(3140));
    layer7_outputs(1522) <= not(layer6_outputs(1325));
    layer7_outputs(1523) <= '1';
    layer7_outputs(1524) <= '1';
    layer7_outputs(1525) <= (layer6_outputs(1587)) or (layer6_outputs(1321));
    layer7_outputs(1526) <= layer6_outputs(3397);
    layer7_outputs(1527) <= not((layer6_outputs(4623)) xor (layer6_outputs(4394)));
    layer7_outputs(1528) <= layer6_outputs(4698);
    layer7_outputs(1529) <= layer6_outputs(354);
    layer7_outputs(1530) <= (layer6_outputs(1345)) and not (layer6_outputs(2529));
    layer7_outputs(1531) <= (layer6_outputs(678)) or (layer6_outputs(943));
    layer7_outputs(1532) <= not(layer6_outputs(3407)) or (layer6_outputs(3076));
    layer7_outputs(1533) <= not(layer6_outputs(1259));
    layer7_outputs(1534) <= not((layer6_outputs(1885)) and (layer6_outputs(195)));
    layer7_outputs(1535) <= layer6_outputs(3016);
    layer7_outputs(1536) <= layer6_outputs(1648);
    layer7_outputs(1537) <= layer6_outputs(3457);
    layer7_outputs(1538) <= (layer6_outputs(4054)) or (layer6_outputs(4532));
    layer7_outputs(1539) <= not(layer6_outputs(5051));
    layer7_outputs(1540) <= (layer6_outputs(1890)) and not (layer6_outputs(3539));
    layer7_outputs(1541) <= not(layer6_outputs(2117));
    layer7_outputs(1542) <= not((layer6_outputs(4440)) xor (layer6_outputs(4237)));
    layer7_outputs(1543) <= layer6_outputs(14);
    layer7_outputs(1544) <= not(layer6_outputs(447));
    layer7_outputs(1545) <= '0';
    layer7_outputs(1546) <= layer6_outputs(2125);
    layer7_outputs(1547) <= not(layer6_outputs(2096));
    layer7_outputs(1548) <= not((layer6_outputs(3100)) and (layer6_outputs(3704)));
    layer7_outputs(1549) <= layer6_outputs(4477);
    layer7_outputs(1550) <= layer6_outputs(2605);
    layer7_outputs(1551) <= not(layer6_outputs(5026));
    layer7_outputs(1552) <= not(layer6_outputs(2120));
    layer7_outputs(1553) <= not(layer6_outputs(4708));
    layer7_outputs(1554) <= not(layer6_outputs(4474)) or (layer6_outputs(2890));
    layer7_outputs(1555) <= (layer6_outputs(2175)) and not (layer6_outputs(1095));
    layer7_outputs(1556) <= layer6_outputs(4818);
    layer7_outputs(1557) <= (layer6_outputs(3286)) or (layer6_outputs(3371));
    layer7_outputs(1558) <= (layer6_outputs(745)) and not (layer6_outputs(169));
    layer7_outputs(1559) <= not((layer6_outputs(4076)) or (layer6_outputs(830)));
    layer7_outputs(1560) <= layer6_outputs(2279);
    layer7_outputs(1561) <= (layer6_outputs(736)) xor (layer6_outputs(4861));
    layer7_outputs(1562) <= not((layer6_outputs(4716)) xor (layer6_outputs(2273)));
    layer7_outputs(1563) <= not(layer6_outputs(873));
    layer7_outputs(1564) <= not(layer6_outputs(3710)) or (layer6_outputs(3316));
    layer7_outputs(1565) <= layer6_outputs(3512);
    layer7_outputs(1566) <= not(layer6_outputs(4990));
    layer7_outputs(1567) <= not((layer6_outputs(1493)) and (layer6_outputs(1494)));
    layer7_outputs(1568) <= not(layer6_outputs(1486));
    layer7_outputs(1569) <= not(layer6_outputs(2620));
    layer7_outputs(1570) <= not((layer6_outputs(637)) or (layer6_outputs(2550)));
    layer7_outputs(1571) <= layer6_outputs(326);
    layer7_outputs(1572) <= layer6_outputs(1115);
    layer7_outputs(1573) <= (layer6_outputs(1847)) and not (layer6_outputs(981));
    layer7_outputs(1574) <= layer6_outputs(2517);
    layer7_outputs(1575) <= not(layer6_outputs(3547)) or (layer6_outputs(238));
    layer7_outputs(1576) <= layer6_outputs(3998);
    layer7_outputs(1577) <= not((layer6_outputs(52)) or (layer6_outputs(712)));
    layer7_outputs(1578) <= layer6_outputs(237);
    layer7_outputs(1579) <= not(layer6_outputs(2062));
    layer7_outputs(1580) <= (layer6_outputs(515)) xor (layer6_outputs(3786));
    layer7_outputs(1581) <= not(layer6_outputs(1586));
    layer7_outputs(1582) <= not(layer6_outputs(3714));
    layer7_outputs(1583) <= layer6_outputs(4688);
    layer7_outputs(1584) <= not(layer6_outputs(2130)) or (layer6_outputs(163));
    layer7_outputs(1585) <= layer6_outputs(915);
    layer7_outputs(1586) <= (layer6_outputs(2098)) xor (layer6_outputs(4855));
    layer7_outputs(1587) <= not((layer6_outputs(1307)) or (layer6_outputs(2846)));
    layer7_outputs(1588) <= '0';
    layer7_outputs(1589) <= layer6_outputs(195);
    layer7_outputs(1590) <= layer6_outputs(3350);
    layer7_outputs(1591) <= (layer6_outputs(4554)) and not (layer6_outputs(1175));
    layer7_outputs(1592) <= not((layer6_outputs(3917)) and (layer6_outputs(946)));
    layer7_outputs(1593) <= layer6_outputs(2864);
    layer7_outputs(1594) <= (layer6_outputs(1664)) xor (layer6_outputs(1507));
    layer7_outputs(1595) <= not(layer6_outputs(1236));
    layer7_outputs(1596) <= not(layer6_outputs(2297));
    layer7_outputs(1597) <= layer6_outputs(2905);
    layer7_outputs(1598) <= layer6_outputs(2384);
    layer7_outputs(1599) <= layer6_outputs(1118);
    layer7_outputs(1600) <= not(layer6_outputs(3736));
    layer7_outputs(1601) <= layer6_outputs(2353);
    layer7_outputs(1602) <= not(layer6_outputs(4182));
    layer7_outputs(1603) <= not((layer6_outputs(1734)) and (layer6_outputs(2988)));
    layer7_outputs(1604) <= not((layer6_outputs(2287)) xor (layer6_outputs(4624)));
    layer7_outputs(1605) <= '1';
    layer7_outputs(1606) <= not(layer6_outputs(1438));
    layer7_outputs(1607) <= (layer6_outputs(246)) and (layer6_outputs(2122));
    layer7_outputs(1608) <= not(layer6_outputs(2675));
    layer7_outputs(1609) <= (layer6_outputs(1135)) xor (layer6_outputs(2398));
    layer7_outputs(1610) <= layer6_outputs(140);
    layer7_outputs(1611) <= not(layer6_outputs(2033)) or (layer6_outputs(2590));
    layer7_outputs(1612) <= not(layer6_outputs(4097));
    layer7_outputs(1613) <= (layer6_outputs(2424)) or (layer6_outputs(3328));
    layer7_outputs(1614) <= layer6_outputs(3112);
    layer7_outputs(1615) <= not(layer6_outputs(779)) or (layer6_outputs(2850));
    layer7_outputs(1616) <= not(layer6_outputs(4570));
    layer7_outputs(1617) <= (layer6_outputs(3554)) and not (layer6_outputs(3613));
    layer7_outputs(1618) <= (layer6_outputs(587)) or (layer6_outputs(4941));
    layer7_outputs(1619) <= not((layer6_outputs(4225)) xor (layer6_outputs(4316)));
    layer7_outputs(1620) <= not((layer6_outputs(3493)) xor (layer6_outputs(3224)));
    layer7_outputs(1621) <= (layer6_outputs(1561)) and not (layer6_outputs(4531));
    layer7_outputs(1622) <= layer6_outputs(2570);
    layer7_outputs(1623) <= (layer6_outputs(3306)) xor (layer6_outputs(794));
    layer7_outputs(1624) <= layer6_outputs(1019);
    layer7_outputs(1625) <= not(layer6_outputs(3234));
    layer7_outputs(1626) <= layer6_outputs(3801);
    layer7_outputs(1627) <= layer6_outputs(2270);
    layer7_outputs(1628) <= (layer6_outputs(3790)) and not (layer6_outputs(1457));
    layer7_outputs(1629) <= not(layer6_outputs(1379)) or (layer6_outputs(297));
    layer7_outputs(1630) <= (layer6_outputs(3885)) or (layer6_outputs(3538));
    layer7_outputs(1631) <= not(layer6_outputs(5117)) or (layer6_outputs(444));
    layer7_outputs(1632) <= not((layer6_outputs(3251)) xor (layer6_outputs(781)));
    layer7_outputs(1633) <= not(layer6_outputs(2713));
    layer7_outputs(1634) <= not(layer6_outputs(634));
    layer7_outputs(1635) <= not((layer6_outputs(4040)) xor (layer6_outputs(656)));
    layer7_outputs(1636) <= layer6_outputs(2538);
    layer7_outputs(1637) <= (layer6_outputs(2591)) and not (layer6_outputs(3204));
    layer7_outputs(1638) <= layer6_outputs(1465);
    layer7_outputs(1639) <= not(layer6_outputs(4659));
    layer7_outputs(1640) <= not(layer6_outputs(2087));
    layer7_outputs(1641) <= not(layer6_outputs(518));
    layer7_outputs(1642) <= layer6_outputs(3282);
    layer7_outputs(1643) <= layer6_outputs(2437);
    layer7_outputs(1644) <= not(layer6_outputs(3936));
    layer7_outputs(1645) <= layer6_outputs(3035);
    layer7_outputs(1646) <= layer6_outputs(4347);
    layer7_outputs(1647) <= not((layer6_outputs(4738)) or (layer6_outputs(426)));
    layer7_outputs(1648) <= layer6_outputs(2938);
    layer7_outputs(1649) <= layer6_outputs(1647);
    layer7_outputs(1650) <= layer6_outputs(1738);
    layer7_outputs(1651) <= not((layer6_outputs(1331)) xor (layer6_outputs(4180)));
    layer7_outputs(1652) <= layer6_outputs(2358);
    layer7_outputs(1653) <= not(layer6_outputs(2350));
    layer7_outputs(1654) <= not(layer6_outputs(3843)) or (layer6_outputs(4294));
    layer7_outputs(1655) <= not(layer6_outputs(583));
    layer7_outputs(1656) <= not(layer6_outputs(4591));
    layer7_outputs(1657) <= layer6_outputs(70);
    layer7_outputs(1658) <= layer6_outputs(482);
    layer7_outputs(1659) <= layer6_outputs(4792);
    layer7_outputs(1660) <= not((layer6_outputs(4348)) xor (layer6_outputs(113)));
    layer7_outputs(1661) <= not(layer6_outputs(4542));
    layer7_outputs(1662) <= not(layer6_outputs(3041));
    layer7_outputs(1663) <= not(layer6_outputs(2255));
    layer7_outputs(1664) <= layer6_outputs(4411);
    layer7_outputs(1665) <= (layer6_outputs(416)) or (layer6_outputs(2236));
    layer7_outputs(1666) <= layer6_outputs(4792);
    layer7_outputs(1667) <= not(layer6_outputs(858));
    layer7_outputs(1668) <= not(layer6_outputs(4350));
    layer7_outputs(1669) <= (layer6_outputs(1052)) and not (layer6_outputs(412));
    layer7_outputs(1670) <= not((layer6_outputs(3080)) xor (layer6_outputs(4449)));
    layer7_outputs(1671) <= (layer6_outputs(4340)) and not (layer6_outputs(1462));
    layer7_outputs(1672) <= layer6_outputs(780);
    layer7_outputs(1673) <= not((layer6_outputs(2231)) xor (layer6_outputs(876)));
    layer7_outputs(1674) <= not((layer6_outputs(1038)) or (layer6_outputs(572)));
    layer7_outputs(1675) <= layer6_outputs(3505);
    layer7_outputs(1676) <= layer6_outputs(965);
    layer7_outputs(1677) <= layer6_outputs(3452);
    layer7_outputs(1678) <= not(layer6_outputs(864));
    layer7_outputs(1679) <= layer6_outputs(2463);
    layer7_outputs(1680) <= not((layer6_outputs(3468)) and (layer6_outputs(3621)));
    layer7_outputs(1681) <= (layer6_outputs(2046)) xor (layer6_outputs(1266));
    layer7_outputs(1682) <= not((layer6_outputs(3534)) xor (layer6_outputs(3586)));
    layer7_outputs(1683) <= not((layer6_outputs(2219)) or (layer6_outputs(1761)));
    layer7_outputs(1684) <= (layer6_outputs(2909)) and not (layer6_outputs(2842));
    layer7_outputs(1685) <= not((layer6_outputs(5035)) or (layer6_outputs(3827)));
    layer7_outputs(1686) <= not(layer6_outputs(421));
    layer7_outputs(1687) <= (layer6_outputs(4323)) and not (layer6_outputs(3238));
    layer7_outputs(1688) <= not(layer6_outputs(578));
    layer7_outputs(1689) <= not(layer6_outputs(1221)) or (layer6_outputs(4737));
    layer7_outputs(1690) <= not((layer6_outputs(4094)) xor (layer6_outputs(1252)));
    layer7_outputs(1691) <= not(layer6_outputs(4784));
    layer7_outputs(1692) <= not(layer6_outputs(2223));
    layer7_outputs(1693) <= not(layer6_outputs(4454));
    layer7_outputs(1694) <= not(layer6_outputs(3549)) or (layer6_outputs(4806));
    layer7_outputs(1695) <= (layer6_outputs(2933)) xor (layer6_outputs(1966));
    layer7_outputs(1696) <= '1';
    layer7_outputs(1697) <= (layer6_outputs(1536)) and not (layer6_outputs(2563));
    layer7_outputs(1698) <= (layer6_outputs(5042)) xor (layer6_outputs(657));
    layer7_outputs(1699) <= (layer6_outputs(1896)) and not (layer6_outputs(3901));
    layer7_outputs(1700) <= layer6_outputs(193);
    layer7_outputs(1701) <= not(layer6_outputs(2468));
    layer7_outputs(1702) <= not(layer6_outputs(3385));
    layer7_outputs(1703) <= not(layer6_outputs(378));
    layer7_outputs(1704) <= layer6_outputs(137);
    layer7_outputs(1705) <= (layer6_outputs(524)) and not (layer6_outputs(4884));
    layer7_outputs(1706) <= layer6_outputs(3596);
    layer7_outputs(1707) <= not(layer6_outputs(397));
    layer7_outputs(1708) <= layer6_outputs(4888);
    layer7_outputs(1709) <= layer6_outputs(929);
    layer7_outputs(1710) <= (layer6_outputs(2259)) and (layer6_outputs(2468));
    layer7_outputs(1711) <= (layer6_outputs(1931)) and not (layer6_outputs(1264));
    layer7_outputs(1712) <= layer6_outputs(644);
    layer7_outputs(1713) <= layer6_outputs(2881);
    layer7_outputs(1714) <= (layer6_outputs(114)) xor (layer6_outputs(4019));
    layer7_outputs(1715) <= not((layer6_outputs(4868)) xor (layer6_outputs(1357)));
    layer7_outputs(1716) <= not(layer6_outputs(3074));
    layer7_outputs(1717) <= (layer6_outputs(3812)) and not (layer6_outputs(1472));
    layer7_outputs(1718) <= (layer6_outputs(1189)) and not (layer6_outputs(4425));
    layer7_outputs(1719) <= layer6_outputs(2076);
    layer7_outputs(1720) <= layer6_outputs(1401);
    layer7_outputs(1721) <= not(layer6_outputs(603)) or (layer6_outputs(2642));
    layer7_outputs(1722) <= (layer6_outputs(41)) and not (layer6_outputs(2427));
    layer7_outputs(1723) <= layer6_outputs(189);
    layer7_outputs(1724) <= (layer6_outputs(4431)) and not (layer6_outputs(3336));
    layer7_outputs(1725) <= (layer6_outputs(1773)) or (layer6_outputs(3121));
    layer7_outputs(1726) <= (layer6_outputs(5004)) xor (layer6_outputs(1520));
    layer7_outputs(1727) <= not((layer6_outputs(4786)) xor (layer6_outputs(1285)));
    layer7_outputs(1728) <= not(layer6_outputs(4594));
    layer7_outputs(1729) <= layer6_outputs(4177);
    layer7_outputs(1730) <= layer6_outputs(1956);
    layer7_outputs(1731) <= layer6_outputs(1668);
    layer7_outputs(1732) <= not(layer6_outputs(2558)) or (layer6_outputs(4429));
    layer7_outputs(1733) <= layer6_outputs(1122);
    layer7_outputs(1734) <= layer6_outputs(764);
    layer7_outputs(1735) <= layer6_outputs(1876);
    layer7_outputs(1736) <= not((layer6_outputs(4856)) and (layer6_outputs(2403)));
    layer7_outputs(1737) <= not(layer6_outputs(716)) or (layer6_outputs(1109));
    layer7_outputs(1738) <= layer6_outputs(4584);
    layer7_outputs(1739) <= (layer6_outputs(2876)) or (layer6_outputs(868));
    layer7_outputs(1740) <= not(layer6_outputs(2611));
    layer7_outputs(1741) <= not((layer6_outputs(4333)) xor (layer6_outputs(1550)));
    layer7_outputs(1742) <= (layer6_outputs(3467)) xor (layer6_outputs(4964));
    layer7_outputs(1743) <= (layer6_outputs(293)) and not (layer6_outputs(2427));
    layer7_outputs(1744) <= not(layer6_outputs(4787));
    layer7_outputs(1745) <= layer6_outputs(4330);
    layer7_outputs(1746) <= (layer6_outputs(2447)) and not (layer6_outputs(785));
    layer7_outputs(1747) <= layer6_outputs(4893);
    layer7_outputs(1748) <= not(layer6_outputs(2704));
    layer7_outputs(1749) <= not(layer6_outputs(3066));
    layer7_outputs(1750) <= not(layer6_outputs(1039)) or (layer6_outputs(559));
    layer7_outputs(1751) <= (layer6_outputs(3484)) and not (layer6_outputs(1893));
    layer7_outputs(1752) <= (layer6_outputs(4271)) and not (layer6_outputs(798));
    layer7_outputs(1753) <= (layer6_outputs(3387)) xor (layer6_outputs(89));
    layer7_outputs(1754) <= (layer6_outputs(646)) or (layer6_outputs(4351));
    layer7_outputs(1755) <= not(layer6_outputs(2616));
    layer7_outputs(1756) <= not(layer6_outputs(4844));
    layer7_outputs(1757) <= not(layer6_outputs(1167));
    layer7_outputs(1758) <= (layer6_outputs(2955)) xor (layer6_outputs(4731));
    layer7_outputs(1759) <= layer6_outputs(4503);
    layer7_outputs(1760) <= (layer6_outputs(575)) and (layer6_outputs(3923));
    layer7_outputs(1761) <= not(layer6_outputs(3435));
    layer7_outputs(1762) <= layer6_outputs(3055);
    layer7_outputs(1763) <= not((layer6_outputs(2126)) xor (layer6_outputs(881)));
    layer7_outputs(1764) <= not((layer6_outputs(3638)) or (layer6_outputs(1013)));
    layer7_outputs(1765) <= not(layer6_outputs(2306));
    layer7_outputs(1766) <= not(layer6_outputs(2674));
    layer7_outputs(1767) <= (layer6_outputs(3825)) and (layer6_outputs(4988));
    layer7_outputs(1768) <= not(layer6_outputs(2649)) or (layer6_outputs(4740));
    layer7_outputs(1769) <= (layer6_outputs(480)) and not (layer6_outputs(1591));
    layer7_outputs(1770) <= not(layer6_outputs(4114));
    layer7_outputs(1771) <= (layer6_outputs(2966)) and (layer6_outputs(277));
    layer7_outputs(1772) <= not(layer6_outputs(1741));
    layer7_outputs(1773) <= (layer6_outputs(735)) and (layer6_outputs(1864));
    layer7_outputs(1774) <= not(layer6_outputs(683));
    layer7_outputs(1775) <= layer6_outputs(1905);
    layer7_outputs(1776) <= not((layer6_outputs(1862)) and (layer6_outputs(4420)));
    layer7_outputs(1777) <= layer6_outputs(2026);
    layer7_outputs(1778) <= (layer6_outputs(2081)) xor (layer6_outputs(434));
    layer7_outputs(1779) <= not(layer6_outputs(948));
    layer7_outputs(1780) <= layer6_outputs(802);
    layer7_outputs(1781) <= layer6_outputs(4341);
    layer7_outputs(1782) <= (layer6_outputs(1419)) and not (layer6_outputs(3702));
    layer7_outputs(1783) <= not((layer6_outputs(4819)) xor (layer6_outputs(2724)));
    layer7_outputs(1784) <= '1';
    layer7_outputs(1785) <= not((layer6_outputs(4771)) or (layer6_outputs(2019)));
    layer7_outputs(1786) <= layer6_outputs(4846);
    layer7_outputs(1787) <= not((layer6_outputs(3773)) xor (layer6_outputs(4762)));
    layer7_outputs(1788) <= layer6_outputs(2323);
    layer7_outputs(1789) <= layer6_outputs(3580);
    layer7_outputs(1790) <= not(layer6_outputs(2207));
    layer7_outputs(1791) <= '1';
    layer7_outputs(1792) <= not((layer6_outputs(2773)) and (layer6_outputs(3445)));
    layer7_outputs(1793) <= not(layer6_outputs(4332));
    layer7_outputs(1794) <= layer6_outputs(3738);
    layer7_outputs(1795) <= layer6_outputs(4248);
    layer7_outputs(1796) <= not(layer6_outputs(724));
    layer7_outputs(1797) <= not(layer6_outputs(3278)) or (layer6_outputs(1869));
    layer7_outputs(1798) <= not(layer6_outputs(3049));
    layer7_outputs(1799) <= not(layer6_outputs(762));
    layer7_outputs(1800) <= layer6_outputs(1045);
    layer7_outputs(1801) <= (layer6_outputs(3834)) and not (layer6_outputs(3254));
    layer7_outputs(1802) <= not((layer6_outputs(2572)) xor (layer6_outputs(4631)));
    layer7_outputs(1803) <= (layer6_outputs(2745)) xor (layer6_outputs(1098));
    layer7_outputs(1804) <= not(layer6_outputs(4349));
    layer7_outputs(1805) <= not((layer6_outputs(1028)) or (layer6_outputs(2243)));
    layer7_outputs(1806) <= not((layer6_outputs(4121)) and (layer6_outputs(4084)));
    layer7_outputs(1807) <= not(layer6_outputs(1848));
    layer7_outputs(1808) <= (layer6_outputs(4344)) and not (layer6_outputs(4072));
    layer7_outputs(1809) <= not(layer6_outputs(767));
    layer7_outputs(1810) <= not(layer6_outputs(2866));
    layer7_outputs(1811) <= (layer6_outputs(881)) and (layer6_outputs(4565));
    layer7_outputs(1812) <= not(layer6_outputs(4292));
    layer7_outputs(1813) <= (layer6_outputs(2376)) and not (layer6_outputs(1021));
    layer7_outputs(1814) <= (layer6_outputs(3688)) xor (layer6_outputs(1526));
    layer7_outputs(1815) <= not((layer6_outputs(4800)) or (layer6_outputs(348)));
    layer7_outputs(1816) <= (layer6_outputs(3371)) xor (layer6_outputs(2399));
    layer7_outputs(1817) <= '0';
    layer7_outputs(1818) <= not(layer6_outputs(1978));
    layer7_outputs(1819) <= (layer6_outputs(1321)) xor (layer6_outputs(833));
    layer7_outputs(1820) <= layer6_outputs(505);
    layer7_outputs(1821) <= (layer6_outputs(3859)) and (layer6_outputs(4318));
    layer7_outputs(1822) <= layer6_outputs(2680);
    layer7_outputs(1823) <= layer6_outputs(5099);
    layer7_outputs(1824) <= (layer6_outputs(1637)) or (layer6_outputs(440));
    layer7_outputs(1825) <= not(layer6_outputs(504)) or (layer6_outputs(1312));
    layer7_outputs(1826) <= (layer6_outputs(1657)) and not (layer6_outputs(3022));
    layer7_outputs(1827) <= not(layer6_outputs(930));
    layer7_outputs(1828) <= (layer6_outputs(1306)) and not (layer6_outputs(2706));
    layer7_outputs(1829) <= layer6_outputs(672);
    layer7_outputs(1830) <= layer6_outputs(4967);
    layer7_outputs(1831) <= layer6_outputs(3664);
    layer7_outputs(1832) <= layer6_outputs(936);
    layer7_outputs(1833) <= not((layer6_outputs(2631)) xor (layer6_outputs(3259)));
    layer7_outputs(1834) <= layer6_outputs(2887);
    layer7_outputs(1835) <= not((layer6_outputs(4272)) and (layer6_outputs(4794)));
    layer7_outputs(1836) <= not((layer6_outputs(3583)) or (layer6_outputs(1705)));
    layer7_outputs(1837) <= (layer6_outputs(4896)) and (layer6_outputs(3491));
    layer7_outputs(1838) <= layer6_outputs(959);
    layer7_outputs(1839) <= layer6_outputs(1735);
    layer7_outputs(1840) <= not(layer6_outputs(2458));
    layer7_outputs(1841) <= not((layer6_outputs(4251)) and (layer6_outputs(4306)));
    layer7_outputs(1842) <= not(layer6_outputs(1420));
    layer7_outputs(1843) <= not(layer6_outputs(908));
    layer7_outputs(1844) <= (layer6_outputs(1361)) and not (layer6_outputs(4844));
    layer7_outputs(1845) <= (layer6_outputs(4376)) or (layer6_outputs(2551));
    layer7_outputs(1846) <= not(layer6_outputs(4660));
    layer7_outputs(1847) <= not(layer6_outputs(4008));
    layer7_outputs(1848) <= not((layer6_outputs(117)) or (layer6_outputs(619)));
    layer7_outputs(1849) <= layer6_outputs(4278);
    layer7_outputs(1850) <= layer6_outputs(3071);
    layer7_outputs(1851) <= not((layer6_outputs(1831)) xor (layer6_outputs(540)));
    layer7_outputs(1852) <= not((layer6_outputs(1548)) xor (layer6_outputs(1698)));
    layer7_outputs(1853) <= not(layer6_outputs(2573));
    layer7_outputs(1854) <= not(layer6_outputs(4873));
    layer7_outputs(1855) <= not(layer6_outputs(793));
    layer7_outputs(1856) <= (layer6_outputs(5080)) and not (layer6_outputs(4233));
    layer7_outputs(1857) <= layer6_outputs(1025);
    layer7_outputs(1858) <= not(layer6_outputs(1958));
    layer7_outputs(1859) <= not((layer6_outputs(1363)) xor (layer6_outputs(3277)));
    layer7_outputs(1860) <= not(layer6_outputs(469));
    layer7_outputs(1861) <= (layer6_outputs(3602)) xor (layer6_outputs(4104));
    layer7_outputs(1862) <= not(layer6_outputs(4137));
    layer7_outputs(1863) <= layer6_outputs(3261);
    layer7_outputs(1864) <= layer6_outputs(74);
    layer7_outputs(1865) <= not((layer6_outputs(3352)) xor (layer6_outputs(4812)));
    layer7_outputs(1866) <= not(layer6_outputs(4301)) or (layer6_outputs(1294));
    layer7_outputs(1867) <= layer6_outputs(475);
    layer7_outputs(1868) <= layer6_outputs(4254);
    layer7_outputs(1869) <= layer6_outputs(75);
    layer7_outputs(1870) <= layer6_outputs(1401);
    layer7_outputs(1871) <= (layer6_outputs(4150)) or (layer6_outputs(4416));
    layer7_outputs(1872) <= not(layer6_outputs(3004));
    layer7_outputs(1873) <= not(layer6_outputs(50));
    layer7_outputs(1874) <= not((layer6_outputs(58)) xor (layer6_outputs(1089)));
    layer7_outputs(1875) <= (layer6_outputs(413)) xor (layer6_outputs(2140));
    layer7_outputs(1876) <= not((layer6_outputs(5083)) xor (layer6_outputs(3924)));
    layer7_outputs(1877) <= layer6_outputs(3252);
    layer7_outputs(1878) <= not(layer6_outputs(4638));
    layer7_outputs(1879) <= not((layer6_outputs(32)) or (layer6_outputs(3755)));
    layer7_outputs(1880) <= not(layer6_outputs(3774)) or (layer6_outputs(2671));
    layer7_outputs(1881) <= (layer6_outputs(2050)) or (layer6_outputs(4621));
    layer7_outputs(1882) <= layer6_outputs(3452);
    layer7_outputs(1883) <= not((layer6_outputs(1595)) and (layer6_outputs(831)));
    layer7_outputs(1884) <= layer6_outputs(3347);
    layer7_outputs(1885) <= (layer6_outputs(3455)) and not (layer6_outputs(3733));
    layer7_outputs(1886) <= (layer6_outputs(3168)) and not (layer6_outputs(854));
    layer7_outputs(1887) <= (layer6_outputs(2856)) and (layer6_outputs(4361));
    layer7_outputs(1888) <= (layer6_outputs(2693)) xor (layer6_outputs(2313));
    layer7_outputs(1889) <= not(layer6_outputs(3771));
    layer7_outputs(1890) <= not(layer6_outputs(4938));
    layer7_outputs(1891) <= not(layer6_outputs(326));
    layer7_outputs(1892) <= (layer6_outputs(4406)) and not (layer6_outputs(3837));
    layer7_outputs(1893) <= (layer6_outputs(4261)) and not (layer6_outputs(4499));
    layer7_outputs(1894) <= layer6_outputs(4288);
    layer7_outputs(1895) <= layer6_outputs(948);
    layer7_outputs(1896) <= not(layer6_outputs(209));
    layer7_outputs(1897) <= layer6_outputs(4850);
    layer7_outputs(1898) <= layer6_outputs(3865);
    layer7_outputs(1899) <= not((layer6_outputs(3383)) xor (layer6_outputs(2872)));
    layer7_outputs(1900) <= layer6_outputs(35);
    layer7_outputs(1901) <= (layer6_outputs(3484)) and not (layer6_outputs(2498));
    layer7_outputs(1902) <= not((layer6_outputs(1931)) and (layer6_outputs(54)));
    layer7_outputs(1903) <= layer6_outputs(4257);
    layer7_outputs(1904) <= not((layer6_outputs(4857)) xor (layer6_outputs(800)));
    layer7_outputs(1905) <= layer6_outputs(3346);
    layer7_outputs(1906) <= layer6_outputs(4729);
    layer7_outputs(1907) <= not((layer6_outputs(1814)) and (layer6_outputs(3241)));
    layer7_outputs(1908) <= layer6_outputs(4891);
    layer7_outputs(1909) <= '0';
    layer7_outputs(1910) <= not(layer6_outputs(347));
    layer7_outputs(1911) <= layer6_outputs(883);
    layer7_outputs(1912) <= layer6_outputs(1216);
    layer7_outputs(1913) <= not((layer6_outputs(1582)) or (layer6_outputs(783)));
    layer7_outputs(1914) <= layer6_outputs(4709);
    layer7_outputs(1915) <= (layer6_outputs(2901)) xor (layer6_outputs(3535));
    layer7_outputs(1916) <= not(layer6_outputs(477));
    layer7_outputs(1917) <= layer6_outputs(1530);
    layer7_outputs(1918) <= (layer6_outputs(416)) xor (layer6_outputs(3600));
    layer7_outputs(1919) <= layer6_outputs(463);
    layer7_outputs(1920) <= not((layer6_outputs(2556)) and (layer6_outputs(2119)));
    layer7_outputs(1921) <= (layer6_outputs(4327)) and not (layer6_outputs(597));
    layer7_outputs(1922) <= layer6_outputs(2483);
    layer7_outputs(1923) <= (layer6_outputs(2329)) and not (layer6_outputs(194));
    layer7_outputs(1924) <= layer6_outputs(1570);
    layer7_outputs(1925) <= (layer6_outputs(4482)) and not (layer6_outputs(5091));
    layer7_outputs(1926) <= layer6_outputs(2057);
    layer7_outputs(1927) <= (layer6_outputs(343)) and (layer6_outputs(4940));
    layer7_outputs(1928) <= not((layer6_outputs(2138)) xor (layer6_outputs(1781)));
    layer7_outputs(1929) <= (layer6_outputs(3421)) and not (layer6_outputs(2078));
    layer7_outputs(1930) <= not((layer6_outputs(1609)) xor (layer6_outputs(4546)));
    layer7_outputs(1931) <= not((layer6_outputs(2229)) xor (layer6_outputs(5096)));
    layer7_outputs(1932) <= (layer6_outputs(396)) xor (layer6_outputs(206));
    layer7_outputs(1933) <= (layer6_outputs(594)) and (layer6_outputs(1753));
    layer7_outputs(1934) <= (layer6_outputs(3059)) and not (layer6_outputs(3486));
    layer7_outputs(1935) <= not(layer6_outputs(4675));
    layer7_outputs(1936) <= (layer6_outputs(1018)) and (layer6_outputs(336));
    layer7_outputs(1937) <= (layer6_outputs(4203)) xor (layer6_outputs(1061));
    layer7_outputs(1938) <= layer6_outputs(2328);
    layer7_outputs(1939) <= not((layer6_outputs(1512)) xor (layer6_outputs(4745)));
    layer7_outputs(1940) <= layer6_outputs(3449);
    layer7_outputs(1941) <= not(layer6_outputs(2453));
    layer7_outputs(1942) <= (layer6_outputs(4346)) and not (layer6_outputs(4179));
    layer7_outputs(1943) <= not((layer6_outputs(1460)) and (layer6_outputs(1203)));
    layer7_outputs(1944) <= not((layer6_outputs(2994)) xor (layer6_outputs(2765)));
    layer7_outputs(1945) <= not(layer6_outputs(660)) or (layer6_outputs(2607));
    layer7_outputs(1946) <= (layer6_outputs(998)) or (layer6_outputs(4250));
    layer7_outputs(1947) <= not((layer6_outputs(2223)) and (layer6_outputs(4206)));
    layer7_outputs(1948) <= not(layer6_outputs(1780)) or (layer6_outputs(3315));
    layer7_outputs(1949) <= not(layer6_outputs(1278));
    layer7_outputs(1950) <= not((layer6_outputs(2574)) xor (layer6_outputs(2286)));
    layer7_outputs(1951) <= not((layer6_outputs(653)) or (layer6_outputs(3030)));
    layer7_outputs(1952) <= layer6_outputs(4426);
    layer7_outputs(1953) <= not((layer6_outputs(3471)) or (layer6_outputs(4037)));
    layer7_outputs(1954) <= not(layer6_outputs(1794));
    layer7_outputs(1955) <= not(layer6_outputs(4985));
    layer7_outputs(1956) <= not(layer6_outputs(5048));
    layer7_outputs(1957) <= not(layer6_outputs(1745));
    layer7_outputs(1958) <= (layer6_outputs(3064)) and (layer6_outputs(2283));
    layer7_outputs(1959) <= not(layer6_outputs(1232));
    layer7_outputs(1960) <= (layer6_outputs(812)) and not (layer6_outputs(1553));
    layer7_outputs(1961) <= (layer6_outputs(1180)) and (layer6_outputs(3529));
    layer7_outputs(1962) <= not(layer6_outputs(3155));
    layer7_outputs(1963) <= not(layer6_outputs(3226));
    layer7_outputs(1964) <= '0';
    layer7_outputs(1965) <= not(layer6_outputs(3540));
    layer7_outputs(1966) <= layer6_outputs(1387);
    layer7_outputs(1967) <= layer6_outputs(976);
    layer7_outputs(1968) <= (layer6_outputs(4345)) and not (layer6_outputs(2395));
    layer7_outputs(1969) <= (layer6_outputs(4669)) xor (layer6_outputs(197));
    layer7_outputs(1970) <= not(layer6_outputs(4067));
    layer7_outputs(1971) <= layer6_outputs(398);
    layer7_outputs(1972) <= not((layer6_outputs(2277)) xor (layer6_outputs(4456)));
    layer7_outputs(1973) <= layer6_outputs(2312);
    layer7_outputs(1974) <= not(layer6_outputs(3574));
    layer7_outputs(1975) <= not(layer6_outputs(2527));
    layer7_outputs(1976) <= not(layer6_outputs(3662));
    layer7_outputs(1977) <= (layer6_outputs(2605)) and (layer6_outputs(3206));
    layer7_outputs(1978) <= not(layer6_outputs(1777)) or (layer6_outputs(1934));
    layer7_outputs(1979) <= not(layer6_outputs(3999)) or (layer6_outputs(1574));
    layer7_outputs(1980) <= layer6_outputs(2345);
    layer7_outputs(1981) <= not((layer6_outputs(2028)) and (layer6_outputs(632)));
    layer7_outputs(1982) <= (layer6_outputs(4834)) and not (layer6_outputs(183));
    layer7_outputs(1983) <= not(layer6_outputs(5110));
    layer7_outputs(1984) <= not(layer6_outputs(2105));
    layer7_outputs(1985) <= not((layer6_outputs(2002)) xor (layer6_outputs(4969)));
    layer7_outputs(1986) <= not(layer6_outputs(1525));
    layer7_outputs(1987) <= not(layer6_outputs(2616));
    layer7_outputs(1988) <= not(layer6_outputs(3283));
    layer7_outputs(1989) <= layer6_outputs(4618);
    layer7_outputs(1990) <= not((layer6_outputs(4361)) and (layer6_outputs(1815)));
    layer7_outputs(1991) <= (layer6_outputs(3928)) xor (layer6_outputs(1734));
    layer7_outputs(1992) <= not(layer6_outputs(1866));
    layer7_outputs(1993) <= (layer6_outputs(4407)) xor (layer6_outputs(4611));
    layer7_outputs(1994) <= not(layer6_outputs(1782));
    layer7_outputs(1995) <= layer6_outputs(1885);
    layer7_outputs(1996) <= not(layer6_outputs(894)) or (layer6_outputs(4738));
    layer7_outputs(1997) <= layer6_outputs(4270);
    layer7_outputs(1998) <= not((layer6_outputs(4552)) or (layer6_outputs(1331)));
    layer7_outputs(1999) <= layer6_outputs(1387);
    layer7_outputs(2000) <= layer6_outputs(4877);
    layer7_outputs(2001) <= not((layer6_outputs(4616)) and (layer6_outputs(1360)));
    layer7_outputs(2002) <= not(layer6_outputs(4901));
    layer7_outputs(2003) <= (layer6_outputs(3655)) or (layer6_outputs(1008));
    layer7_outputs(2004) <= not(layer6_outputs(961));
    layer7_outputs(2005) <= not(layer6_outputs(4310));
    layer7_outputs(2006) <= (layer6_outputs(2701)) and not (layer6_outputs(4869));
    layer7_outputs(2007) <= '1';
    layer7_outputs(2008) <= (layer6_outputs(2063)) and not (layer6_outputs(4968));
    layer7_outputs(2009) <= not((layer6_outputs(1081)) xor (layer6_outputs(4615)));
    layer7_outputs(2010) <= (layer6_outputs(2079)) and not (layer6_outputs(1715));
    layer7_outputs(2011) <= (layer6_outputs(1006)) and not (layer6_outputs(1100));
    layer7_outputs(2012) <= layer6_outputs(4670);
    layer7_outputs(2013) <= layer6_outputs(3254);
    layer7_outputs(2014) <= not(layer6_outputs(674));
    layer7_outputs(2015) <= not((layer6_outputs(3084)) xor (layer6_outputs(528)));
    layer7_outputs(2016) <= not((layer6_outputs(3832)) or (layer6_outputs(3314)));
    layer7_outputs(2017) <= not((layer6_outputs(2969)) or (layer6_outputs(1765)));
    layer7_outputs(2018) <= not(layer6_outputs(4156));
    layer7_outputs(2019) <= not(layer6_outputs(2145)) or (layer6_outputs(1305));
    layer7_outputs(2020) <= not(layer6_outputs(1629));
    layer7_outputs(2021) <= (layer6_outputs(1526)) xor (layer6_outputs(4244));
    layer7_outputs(2022) <= not((layer6_outputs(4556)) xor (layer6_outputs(2633)));
    layer7_outputs(2023) <= not(layer6_outputs(4251));
    layer7_outputs(2024) <= (layer6_outputs(3314)) xor (layer6_outputs(2960));
    layer7_outputs(2025) <= (layer6_outputs(2471)) xor (layer6_outputs(2382));
    layer7_outputs(2026) <= (layer6_outputs(4878)) and (layer6_outputs(3956));
    layer7_outputs(2027) <= layer6_outputs(4811);
    layer7_outputs(2028) <= not(layer6_outputs(3770));
    layer7_outputs(2029) <= not(layer6_outputs(1782));
    layer7_outputs(2030) <= layer6_outputs(1347);
    layer7_outputs(2031) <= layer6_outputs(4338);
    layer7_outputs(2032) <= not((layer6_outputs(3612)) xor (layer6_outputs(3937)));
    layer7_outputs(2033) <= not(layer6_outputs(2104)) or (layer6_outputs(3841));
    layer7_outputs(2034) <= layer6_outputs(3390);
    layer7_outputs(2035) <= (layer6_outputs(4970)) xor (layer6_outputs(2156));
    layer7_outputs(2036) <= not((layer6_outputs(3597)) and (layer6_outputs(1436)));
    layer7_outputs(2037) <= not(layer6_outputs(4944));
    layer7_outputs(2038) <= (layer6_outputs(4125)) xor (layer6_outputs(4448));
    layer7_outputs(2039) <= not((layer6_outputs(4902)) and (layer6_outputs(3191)));
    layer7_outputs(2040) <= not(layer6_outputs(2216));
    layer7_outputs(2041) <= not(layer6_outputs(1415));
    layer7_outputs(2042) <= not((layer6_outputs(4568)) xor (layer6_outputs(4024)));
    layer7_outputs(2043) <= layer6_outputs(4979);
    layer7_outputs(2044) <= (layer6_outputs(952)) or (layer6_outputs(1631));
    layer7_outputs(2045) <= not((layer6_outputs(5073)) xor (layer6_outputs(2276)));
    layer7_outputs(2046) <= (layer6_outputs(271)) and not (layer6_outputs(4937));
    layer7_outputs(2047) <= not((layer6_outputs(3909)) and (layer6_outputs(2301)));
    layer7_outputs(2048) <= not(layer6_outputs(2407)) or (layer6_outputs(2305));
    layer7_outputs(2049) <= (layer6_outputs(3594)) or (layer6_outputs(4957));
    layer7_outputs(2050) <= layer6_outputs(1652);
    layer7_outputs(2051) <= not(layer6_outputs(3192)) or (layer6_outputs(5036));
    layer7_outputs(2052) <= (layer6_outputs(772)) xor (layer6_outputs(414));
    layer7_outputs(2053) <= (layer6_outputs(1730)) and not (layer6_outputs(4445));
    layer7_outputs(2054) <= not(layer6_outputs(506));
    layer7_outputs(2055) <= not(layer6_outputs(1705));
    layer7_outputs(2056) <= not(layer6_outputs(4495));
    layer7_outputs(2057) <= not(layer6_outputs(3437));
    layer7_outputs(2058) <= not(layer6_outputs(1713)) or (layer6_outputs(2));
    layer7_outputs(2059) <= not((layer6_outputs(2592)) xor (layer6_outputs(3661)));
    layer7_outputs(2060) <= (layer6_outputs(5015)) xor (layer6_outputs(2337));
    layer7_outputs(2061) <= (layer6_outputs(1994)) xor (layer6_outputs(4105));
    layer7_outputs(2062) <= not((layer6_outputs(157)) or (layer6_outputs(687)));
    layer7_outputs(2063) <= not(layer6_outputs(2830)) or (layer6_outputs(801));
    layer7_outputs(2064) <= layer6_outputs(1594);
    layer7_outputs(2065) <= '0';
    layer7_outputs(2066) <= layer6_outputs(4443);
    layer7_outputs(2067) <= not(layer6_outputs(4321));
    layer7_outputs(2068) <= not(layer6_outputs(12));
    layer7_outputs(2069) <= layer6_outputs(1665);
    layer7_outputs(2070) <= layer6_outputs(4205);
    layer7_outputs(2071) <= not(layer6_outputs(2603));
    layer7_outputs(2072) <= not(layer6_outputs(177)) or (layer6_outputs(715));
    layer7_outputs(2073) <= not((layer6_outputs(983)) xor (layer6_outputs(1057)));
    layer7_outputs(2074) <= layer6_outputs(2526);
    layer7_outputs(2075) <= layer6_outputs(3399);
    layer7_outputs(2076) <= layer6_outputs(1878);
    layer7_outputs(2077) <= layer6_outputs(4200);
    layer7_outputs(2078) <= not(layer6_outputs(1047));
    layer7_outputs(2079) <= (layer6_outputs(1919)) or (layer6_outputs(1064));
    layer7_outputs(2080) <= not(layer6_outputs(721)) or (layer6_outputs(2170));
    layer7_outputs(2081) <= (layer6_outputs(3728)) xor (layer6_outputs(2813));
    layer7_outputs(2082) <= layer6_outputs(3917);
    layer7_outputs(2083) <= '1';
    layer7_outputs(2084) <= not(layer6_outputs(921));
    layer7_outputs(2085) <= layer6_outputs(256);
    layer7_outputs(2086) <= not((layer6_outputs(313)) xor (layer6_outputs(2704)));
    layer7_outputs(2087) <= (layer6_outputs(4463)) and not (layer6_outputs(2177));
    layer7_outputs(2088) <= not(layer6_outputs(2467));
    layer7_outputs(2089) <= (layer6_outputs(2558)) xor (layer6_outputs(4284));
    layer7_outputs(2090) <= layer6_outputs(3797);
    layer7_outputs(2091) <= not(layer6_outputs(1992));
    layer7_outputs(2092) <= not((layer6_outputs(4400)) and (layer6_outputs(1910)));
    layer7_outputs(2093) <= not(layer6_outputs(1258));
    layer7_outputs(2094) <= layer6_outputs(3349);
    layer7_outputs(2095) <= (layer6_outputs(2466)) xor (layer6_outputs(759));
    layer7_outputs(2096) <= layer6_outputs(1045);
    layer7_outputs(2097) <= (layer6_outputs(2501)) and not (layer6_outputs(467));
    layer7_outputs(2098) <= not((layer6_outputs(3792)) xor (layer6_outputs(3874)));
    layer7_outputs(2099) <= (layer6_outputs(2089)) xor (layer6_outputs(2266));
    layer7_outputs(2100) <= not(layer6_outputs(4505));
    layer7_outputs(2101) <= layer6_outputs(568);
    layer7_outputs(2102) <= not(layer6_outputs(1484));
    layer7_outputs(2103) <= not((layer6_outputs(889)) xor (layer6_outputs(4853)));
    layer7_outputs(2104) <= (layer6_outputs(1590)) xor (layer6_outputs(3963));
    layer7_outputs(2105) <= (layer6_outputs(2269)) xor (layer6_outputs(4830));
    layer7_outputs(2106) <= not(layer6_outputs(1167));
    layer7_outputs(2107) <= (layer6_outputs(3393)) and not (layer6_outputs(1627));
    layer7_outputs(2108) <= (layer6_outputs(4328)) xor (layer6_outputs(3939));
    layer7_outputs(2109) <= not(layer6_outputs(149));
    layer7_outputs(2110) <= not(layer6_outputs(828));
    layer7_outputs(2111) <= (layer6_outputs(435)) or (layer6_outputs(1689));
    layer7_outputs(2112) <= not((layer6_outputs(4836)) or (layer6_outputs(1427)));
    layer7_outputs(2113) <= (layer6_outputs(462)) and not (layer6_outputs(3055));
    layer7_outputs(2114) <= not((layer6_outputs(3643)) xor (layer6_outputs(1652)));
    layer7_outputs(2115) <= (layer6_outputs(602)) and (layer6_outputs(1744));
    layer7_outputs(2116) <= layer6_outputs(1681);
    layer7_outputs(2117) <= not(layer6_outputs(4862)) or (layer6_outputs(1732));
    layer7_outputs(2118) <= layer6_outputs(1810);
    layer7_outputs(2119) <= (layer6_outputs(1024)) and not (layer6_outputs(2302));
    layer7_outputs(2120) <= '0';
    layer7_outputs(2121) <= (layer6_outputs(3133)) and not (layer6_outputs(2293));
    layer7_outputs(2122) <= not((layer6_outputs(1923)) xor (layer6_outputs(3528)));
    layer7_outputs(2123) <= layer6_outputs(2923);
    layer7_outputs(2124) <= layer6_outputs(3752);
    layer7_outputs(2125) <= not(layer6_outputs(2194));
    layer7_outputs(2126) <= layer6_outputs(3573);
    layer7_outputs(2127) <= not(layer6_outputs(1339));
    layer7_outputs(2128) <= layer6_outputs(3577);
    layer7_outputs(2129) <= layer6_outputs(3412);
    layer7_outputs(2130) <= not((layer6_outputs(415)) and (layer6_outputs(2635)));
    layer7_outputs(2131) <= layer6_outputs(938);
    layer7_outputs(2132) <= layer6_outputs(4202);
    layer7_outputs(2133) <= not((layer6_outputs(2536)) xor (layer6_outputs(4883)));
    layer7_outputs(2134) <= not(layer6_outputs(3506));
    layer7_outputs(2135) <= not(layer6_outputs(41));
    layer7_outputs(2136) <= not(layer6_outputs(588)) or (layer6_outputs(844));
    layer7_outputs(2137) <= not((layer6_outputs(3462)) and (layer6_outputs(790)));
    layer7_outputs(2138) <= not(layer6_outputs(2961));
    layer7_outputs(2139) <= not((layer6_outputs(3705)) and (layer6_outputs(186)));
    layer7_outputs(2140) <= '0';
    layer7_outputs(2141) <= (layer6_outputs(3624)) or (layer6_outputs(1330));
    layer7_outputs(2142) <= (layer6_outputs(2543)) and not (layer6_outputs(109));
    layer7_outputs(2143) <= (layer6_outputs(5067)) and (layer6_outputs(72));
    layer7_outputs(2144) <= not((layer6_outputs(580)) and (layer6_outputs(4155)));
    layer7_outputs(2145) <= layer6_outputs(529);
    layer7_outputs(2146) <= (layer6_outputs(3324)) and not (layer6_outputs(335));
    layer7_outputs(2147) <= not(layer6_outputs(2256)) or (layer6_outputs(3083));
    layer7_outputs(2148) <= layer6_outputs(289);
    layer7_outputs(2149) <= layer6_outputs(3360);
    layer7_outputs(2150) <= not(layer6_outputs(429));
    layer7_outputs(2151) <= layer6_outputs(1939);
    layer7_outputs(2152) <= not(layer6_outputs(2343));
    layer7_outputs(2153) <= not((layer6_outputs(3532)) xor (layer6_outputs(3853)));
    layer7_outputs(2154) <= (layer6_outputs(2244)) xor (layer6_outputs(2569));
    layer7_outputs(2155) <= not(layer6_outputs(438));
    layer7_outputs(2156) <= not(layer6_outputs(1164));
    layer7_outputs(2157) <= layer6_outputs(1339);
    layer7_outputs(2158) <= not(layer6_outputs(4131));
    layer7_outputs(2159) <= not(layer6_outputs(1441)) or (layer6_outputs(2525));
    layer7_outputs(2160) <= (layer6_outputs(4873)) xor (layer6_outputs(2110));
    layer7_outputs(2161) <= (layer6_outputs(4795)) and (layer6_outputs(312));
    layer7_outputs(2162) <= not(layer6_outputs(2070));
    layer7_outputs(2163) <= layer6_outputs(1911);
    layer7_outputs(2164) <= layer6_outputs(1644);
    layer7_outputs(2165) <= '0';
    layer7_outputs(2166) <= (layer6_outputs(1605)) and not (layer6_outputs(3300));
    layer7_outputs(2167) <= not(layer6_outputs(1111));
    layer7_outputs(2168) <= (layer6_outputs(819)) xor (layer6_outputs(2184));
    layer7_outputs(2169) <= (layer6_outputs(2741)) and (layer6_outputs(4720));
    layer7_outputs(2170) <= not(layer6_outputs(1490));
    layer7_outputs(2171) <= layer6_outputs(1728);
    layer7_outputs(2172) <= (layer6_outputs(4238)) xor (layer6_outputs(2235));
    layer7_outputs(2173) <= not(layer6_outputs(3630));
    layer7_outputs(2174) <= not(layer6_outputs(2378));
    layer7_outputs(2175) <= (layer6_outputs(2938)) xor (layer6_outputs(1959));
    layer7_outputs(2176) <= layer6_outputs(3824);
    layer7_outputs(2177) <= layer6_outputs(1458);
    layer7_outputs(2178) <= not(layer6_outputs(1753)) or (layer6_outputs(497));
    layer7_outputs(2179) <= layer6_outputs(2545);
    layer7_outputs(2180) <= not(layer6_outputs(2514));
    layer7_outputs(2181) <= not(layer6_outputs(2890)) or (layer6_outputs(1004));
    layer7_outputs(2182) <= not(layer6_outputs(2413));
    layer7_outputs(2183) <= layer6_outputs(3584);
    layer7_outputs(2184) <= not((layer6_outputs(597)) xor (layer6_outputs(76)));
    layer7_outputs(2185) <= layer6_outputs(4143);
    layer7_outputs(2186) <= not(layer6_outputs(1030));
    layer7_outputs(2187) <= (layer6_outputs(2590)) and not (layer6_outputs(4178));
    layer7_outputs(2188) <= layer6_outputs(3981);
    layer7_outputs(2189) <= layer6_outputs(3392);
    layer7_outputs(2190) <= (layer6_outputs(759)) or (layer6_outputs(1037));
    layer7_outputs(2191) <= not((layer6_outputs(2396)) and (layer6_outputs(1743)));
    layer7_outputs(2192) <= (layer6_outputs(1224)) and not (layer6_outputs(4176));
    layer7_outputs(2193) <= (layer6_outputs(577)) or (layer6_outputs(2705));
    layer7_outputs(2194) <= layer6_outputs(1432);
    layer7_outputs(2195) <= (layer6_outputs(1013)) and not (layer6_outputs(666));
    layer7_outputs(2196) <= (layer6_outputs(2092)) and not (layer6_outputs(4865));
    layer7_outputs(2197) <= (layer6_outputs(1770)) and not (layer6_outputs(3280));
    layer7_outputs(2198) <= not(layer6_outputs(2209));
    layer7_outputs(2199) <= not(layer6_outputs(4626));
    layer7_outputs(2200) <= not(layer6_outputs(3478));
    layer7_outputs(2201) <= '0';
    layer7_outputs(2202) <= (layer6_outputs(4583)) and not (layer6_outputs(1857));
    layer7_outputs(2203) <= layer6_outputs(4240);
    layer7_outputs(2204) <= (layer6_outputs(3344)) and not (layer6_outputs(2308));
    layer7_outputs(2205) <= not((layer6_outputs(2141)) xor (layer6_outputs(470)));
    layer7_outputs(2206) <= not((layer6_outputs(3777)) xor (layer6_outputs(2356)));
    layer7_outputs(2207) <= not((layer6_outputs(4567)) and (layer6_outputs(1709)));
    layer7_outputs(2208) <= layer6_outputs(987);
    layer7_outputs(2209) <= not(layer6_outputs(3490));
    layer7_outputs(2210) <= layer6_outputs(266);
    layer7_outputs(2211) <= not(layer6_outputs(3170));
    layer7_outputs(2212) <= not((layer6_outputs(3913)) xor (layer6_outputs(152)));
    layer7_outputs(2213) <= not(layer6_outputs(4393));
    layer7_outputs(2214) <= not(layer6_outputs(3053));
    layer7_outputs(2215) <= layer6_outputs(3033);
    layer7_outputs(2216) <= layer6_outputs(1466);
    layer7_outputs(2217) <= not(layer6_outputs(1669)) or (layer6_outputs(423));
    layer7_outputs(2218) <= not(layer6_outputs(3613));
    layer7_outputs(2219) <= not(layer6_outputs(292));
    layer7_outputs(2220) <= not(layer6_outputs(4536));
    layer7_outputs(2221) <= layer6_outputs(1122);
    layer7_outputs(2222) <= (layer6_outputs(3551)) and not (layer6_outputs(4507));
    layer7_outputs(2223) <= not((layer6_outputs(4625)) or (layer6_outputs(2869)));
    layer7_outputs(2224) <= not(layer6_outputs(2264)) or (layer6_outputs(4022));
    layer7_outputs(2225) <= not(layer6_outputs(4839));
    layer7_outputs(2226) <= (layer6_outputs(3994)) xor (layer6_outputs(730));
    layer7_outputs(2227) <= not((layer6_outputs(1398)) or (layer6_outputs(4489)));
    layer7_outputs(2228) <= not((layer6_outputs(2176)) or (layer6_outputs(11)));
    layer7_outputs(2229) <= not(layer6_outputs(3114)) or (layer6_outputs(3594));
    layer7_outputs(2230) <= layer6_outputs(399);
    layer7_outputs(2231) <= not(layer6_outputs(847));
    layer7_outputs(2232) <= layer6_outputs(3834);
    layer7_outputs(2233) <= not(layer6_outputs(3522));
    layer7_outputs(2234) <= (layer6_outputs(3016)) and not (layer6_outputs(650));
    layer7_outputs(2235) <= (layer6_outputs(4986)) and (layer6_outputs(2693));
    layer7_outputs(2236) <= not(layer6_outputs(2478));
    layer7_outputs(2237) <= not(layer6_outputs(1300));
    layer7_outputs(2238) <= layer6_outputs(3420);
    layer7_outputs(2239) <= not(layer6_outputs(1522));
    layer7_outputs(2240) <= layer6_outputs(4678);
    layer7_outputs(2241) <= layer6_outputs(3929);
    layer7_outputs(2242) <= not((layer6_outputs(1443)) or (layer6_outputs(1241)));
    layer7_outputs(2243) <= not(layer6_outputs(1497));
    layer7_outputs(2244) <= (layer6_outputs(858)) or (layer6_outputs(453));
    layer7_outputs(2245) <= '0';
    layer7_outputs(2246) <= '0';
    layer7_outputs(2247) <= (layer6_outputs(906)) xor (layer6_outputs(960));
    layer7_outputs(2248) <= '0';
    layer7_outputs(2249) <= not(layer6_outputs(3267));
    layer7_outputs(2250) <= layer6_outputs(1860);
    layer7_outputs(2251) <= not(layer6_outputs(4212)) or (layer6_outputs(3787));
    layer7_outputs(2252) <= layer6_outputs(2143);
    layer7_outputs(2253) <= not(layer6_outputs(993));
    layer7_outputs(2254) <= (layer6_outputs(817)) and (layer6_outputs(3675));
    layer7_outputs(2255) <= layer6_outputs(1965);
    layer7_outputs(2256) <= not(layer6_outputs(788));
    layer7_outputs(2257) <= not(layer6_outputs(3838));
    layer7_outputs(2258) <= layer6_outputs(1696);
    layer7_outputs(2259) <= not(layer6_outputs(5100)) or (layer6_outputs(1027));
    layer7_outputs(2260) <= (layer6_outputs(430)) or (layer6_outputs(4501));
    layer7_outputs(2261) <= not((layer6_outputs(1769)) xor (layer6_outputs(4496)));
    layer7_outputs(2262) <= not(layer6_outputs(218));
    layer7_outputs(2263) <= (layer6_outputs(1976)) or (layer6_outputs(3152));
    layer7_outputs(2264) <= not(layer6_outputs(4073));
    layer7_outputs(2265) <= '1';
    layer7_outputs(2266) <= (layer6_outputs(4769)) and (layer6_outputs(2211));
    layer7_outputs(2267) <= (layer6_outputs(3202)) and not (layer6_outputs(2878));
    layer7_outputs(2268) <= layer6_outputs(2945);
    layer7_outputs(2269) <= (layer6_outputs(2311)) or (layer6_outputs(1054));
    layer7_outputs(2270) <= layer6_outputs(234);
    layer7_outputs(2271) <= (layer6_outputs(4067)) xor (layer6_outputs(1873));
    layer7_outputs(2272) <= not(layer6_outputs(2492));
    layer7_outputs(2273) <= layer6_outputs(882);
    layer7_outputs(2274) <= (layer6_outputs(37)) and not (layer6_outputs(204));
    layer7_outputs(2275) <= not(layer6_outputs(1595));
    layer7_outputs(2276) <= (layer6_outputs(2425)) xor (layer6_outputs(3918));
    layer7_outputs(2277) <= not(layer6_outputs(4580));
    layer7_outputs(2278) <= layer6_outputs(4914);
    layer7_outputs(2279) <= not(layer6_outputs(4160));
    layer7_outputs(2280) <= (layer6_outputs(61)) and not (layer6_outputs(4694));
    layer7_outputs(2281) <= not(layer6_outputs(4116));
    layer7_outputs(2282) <= layer6_outputs(4603);
    layer7_outputs(2283) <= layer6_outputs(3850);
    layer7_outputs(2284) <= layer6_outputs(1724);
    layer7_outputs(2285) <= layer6_outputs(110);
    layer7_outputs(2286) <= '1';
    layer7_outputs(2287) <= (layer6_outputs(4602)) or (layer6_outputs(1073));
    layer7_outputs(2288) <= (layer6_outputs(2798)) xor (layer6_outputs(1314));
    layer7_outputs(2289) <= layer6_outputs(988);
    layer7_outputs(2290) <= layer6_outputs(219);
    layer7_outputs(2291) <= not(layer6_outputs(5020));
    layer7_outputs(2292) <= not((layer6_outputs(3206)) and (layer6_outputs(1035)));
    layer7_outputs(2293) <= (layer6_outputs(2004)) xor (layer6_outputs(3123));
    layer7_outputs(2294) <= not(layer6_outputs(314));
    layer7_outputs(2295) <= layer6_outputs(4451);
    layer7_outputs(2296) <= not(layer6_outputs(1542)) or (layer6_outputs(4162));
    layer7_outputs(2297) <= layer6_outputs(2424);
    layer7_outputs(2298) <= (layer6_outputs(534)) and (layer6_outputs(2611));
    layer7_outputs(2299) <= not(layer6_outputs(4353));
    layer7_outputs(2300) <= '1';
    layer7_outputs(2301) <= not(layer6_outputs(2917));
    layer7_outputs(2302) <= (layer6_outputs(1532)) xor (layer6_outputs(164));
    layer7_outputs(2303) <= layer6_outputs(662);
    layer7_outputs(2304) <= (layer6_outputs(1034)) or (layer6_outputs(1382));
    layer7_outputs(2305) <= layer6_outputs(3128);
    layer7_outputs(2306) <= (layer6_outputs(2912)) xor (layer6_outputs(1205));
    layer7_outputs(2307) <= not(layer6_outputs(1113));
    layer7_outputs(2308) <= not(layer6_outputs(4830)) or (layer6_outputs(2177));
    layer7_outputs(2309) <= not((layer6_outputs(1451)) or (layer6_outputs(1774)));
    layer7_outputs(2310) <= not(layer6_outputs(803));
    layer7_outputs(2311) <= not((layer6_outputs(1213)) or (layer6_outputs(1762)));
    layer7_outputs(2312) <= not(layer6_outputs(777));
    layer7_outputs(2313) <= not((layer6_outputs(1461)) xor (layer6_outputs(721)));
    layer7_outputs(2314) <= not(layer6_outputs(3639)) or (layer6_outputs(1619));
    layer7_outputs(2315) <= (layer6_outputs(3171)) and not (layer6_outputs(1593));
    layer7_outputs(2316) <= not((layer6_outputs(2965)) or (layer6_outputs(4971)));
    layer7_outputs(2317) <= layer6_outputs(3565);
    layer7_outputs(2318) <= not((layer6_outputs(2812)) or (layer6_outputs(2131)));
    layer7_outputs(2319) <= not(layer6_outputs(2071));
    layer7_outputs(2320) <= layer6_outputs(4152);
    layer7_outputs(2321) <= not(layer6_outputs(1988));
    layer7_outputs(2322) <= (layer6_outputs(1664)) xor (layer6_outputs(4050));
    layer7_outputs(2323) <= '0';
    layer7_outputs(2324) <= not(layer6_outputs(2615));
    layer7_outputs(2325) <= not((layer6_outputs(2838)) xor (layer6_outputs(3973)));
    layer7_outputs(2326) <= not(layer6_outputs(2578)) or (layer6_outputs(4558));
    layer7_outputs(2327) <= not((layer6_outputs(1610)) or (layer6_outputs(4093)));
    layer7_outputs(2328) <= layer6_outputs(1409);
    layer7_outputs(2329) <= layer6_outputs(563);
    layer7_outputs(2330) <= not(layer6_outputs(902));
    layer7_outputs(2331) <= layer6_outputs(1157);
    layer7_outputs(2332) <= layer6_outputs(2821);
    layer7_outputs(2333) <= not(layer6_outputs(1760));
    layer7_outputs(2334) <= layer6_outputs(3008);
    layer7_outputs(2335) <= (layer6_outputs(1999)) and (layer6_outputs(1806));
    layer7_outputs(2336) <= not(layer6_outputs(144));
    layer7_outputs(2337) <= (layer6_outputs(3354)) or (layer6_outputs(3498));
    layer7_outputs(2338) <= not(layer6_outputs(3178));
    layer7_outputs(2339) <= not(layer6_outputs(492));
    layer7_outputs(2340) <= not(layer6_outputs(2744));
    layer7_outputs(2341) <= (layer6_outputs(481)) xor (layer6_outputs(4168));
    layer7_outputs(2342) <= not(layer6_outputs(4391));
    layer7_outputs(2343) <= not(layer6_outputs(2612));
    layer7_outputs(2344) <= not(layer6_outputs(2475)) or (layer6_outputs(2465));
    layer7_outputs(2345) <= (layer6_outputs(4041)) and not (layer6_outputs(3645));
    layer7_outputs(2346) <= not((layer6_outputs(5075)) xor (layer6_outputs(4933)));
    layer7_outputs(2347) <= not(layer6_outputs(5114));
    layer7_outputs(2348) <= not((layer6_outputs(1396)) xor (layer6_outputs(4858)));
    layer7_outputs(2349) <= not(layer6_outputs(1362)) or (layer6_outputs(1692));
    layer7_outputs(2350) <= not((layer6_outputs(3575)) and (layer6_outputs(5086)));
    layer7_outputs(2351) <= '1';
    layer7_outputs(2352) <= layer6_outputs(4415);
    layer7_outputs(2353) <= layer6_outputs(291);
    layer7_outputs(2354) <= (layer6_outputs(3338)) xor (layer6_outputs(1393));
    layer7_outputs(2355) <= not(layer6_outputs(1083));
    layer7_outputs(2356) <= not(layer6_outputs(3187)) or (layer6_outputs(1015));
    layer7_outputs(2357) <= layer6_outputs(2827);
    layer7_outputs(2358) <= not((layer6_outputs(3128)) xor (layer6_outputs(25)));
    layer7_outputs(2359) <= not(layer6_outputs(1291)) or (layer6_outputs(1545));
    layer7_outputs(2360) <= layer6_outputs(565);
    layer7_outputs(2361) <= (layer6_outputs(1325)) and not (layer6_outputs(2930));
    layer7_outputs(2362) <= (layer6_outputs(2831)) and not (layer6_outputs(4364));
    layer7_outputs(2363) <= layer6_outputs(1458);
    layer7_outputs(2364) <= not(layer6_outputs(3208));
    layer7_outputs(2365) <= layer6_outputs(1702);
    layer7_outputs(2366) <= not(layer6_outputs(2771));
    layer7_outputs(2367) <= not(layer6_outputs(2960)) or (layer6_outputs(1646));
    layer7_outputs(2368) <= (layer6_outputs(5010)) and not (layer6_outputs(3992));
    layer7_outputs(2369) <= layer6_outputs(2862);
    layer7_outputs(2370) <= not(layer6_outputs(1881)) or (layer6_outputs(731));
    layer7_outputs(2371) <= (layer6_outputs(4750)) and not (layer6_outputs(3851));
    layer7_outputs(2372) <= '0';
    layer7_outputs(2373) <= layer6_outputs(4129);
    layer7_outputs(2374) <= (layer6_outputs(3329)) xor (layer6_outputs(2102));
    layer7_outputs(2375) <= (layer6_outputs(230)) or (layer6_outputs(4287));
    layer7_outputs(2376) <= (layer6_outputs(3543)) or (layer6_outputs(4629));
    layer7_outputs(2377) <= layer6_outputs(3249);
    layer7_outputs(2378) <= (layer6_outputs(162)) and (layer6_outputs(385));
    layer7_outputs(2379) <= layer6_outputs(1623);
    layer7_outputs(2380) <= '0';
    layer7_outputs(2381) <= not(layer6_outputs(388));
    layer7_outputs(2382) <= layer6_outputs(1768);
    layer7_outputs(2383) <= layer6_outputs(2714);
    layer7_outputs(2384) <= (layer6_outputs(2412)) or (layer6_outputs(337));
    layer7_outputs(2385) <= not(layer6_outputs(643)) or (layer6_outputs(3595));
    layer7_outputs(2386) <= layer6_outputs(213);
    layer7_outputs(2387) <= not(layer6_outputs(2132));
    layer7_outputs(2388) <= layer6_outputs(1349);
    layer7_outputs(2389) <= layer6_outputs(3336);
    layer7_outputs(2390) <= not(layer6_outputs(579)) or (layer6_outputs(608));
    layer7_outputs(2391) <= layer6_outputs(3908);
    layer7_outputs(2392) <= layer6_outputs(712);
    layer7_outputs(2393) <= (layer6_outputs(3027)) or (layer6_outputs(4451));
    layer7_outputs(2394) <= (layer6_outputs(592)) and not (layer6_outputs(2287));
    layer7_outputs(2395) <= (layer6_outputs(1916)) and not (layer6_outputs(4265));
    layer7_outputs(2396) <= '0';
    layer7_outputs(2397) <= not(layer6_outputs(2668));
    layer7_outputs(2398) <= not((layer6_outputs(1723)) xor (layer6_outputs(2715)));
    layer7_outputs(2399) <= not(layer6_outputs(4925));
    layer7_outputs(2400) <= layer6_outputs(1670);
    layer7_outputs(2401) <= (layer6_outputs(723)) and (layer6_outputs(2009));
    layer7_outputs(2402) <= not((layer6_outputs(4653)) xor (layer6_outputs(4468)));
    layer7_outputs(2403) <= (layer6_outputs(754)) and not (layer6_outputs(3309));
    layer7_outputs(2404) <= not((layer6_outputs(1611)) or (layer6_outputs(1182)));
    layer7_outputs(2405) <= not(layer6_outputs(2702)) or (layer6_outputs(4081));
    layer7_outputs(2406) <= not((layer6_outputs(4469)) and (layer6_outputs(247)));
    layer7_outputs(2407) <= not(layer6_outputs(814));
    layer7_outputs(2408) <= layer6_outputs(2555);
    layer7_outputs(2409) <= not(layer6_outputs(3902));
    layer7_outputs(2410) <= not((layer6_outputs(4055)) xor (layer6_outputs(4646)));
    layer7_outputs(2411) <= (layer6_outputs(4334)) and not (layer6_outputs(3465));
    layer7_outputs(2412) <= not(layer6_outputs(3042));
    layer7_outputs(2413) <= layer6_outputs(2606);
    layer7_outputs(2414) <= not(layer6_outputs(1972)) or (layer6_outputs(1620));
    layer7_outputs(2415) <= (layer6_outputs(3501)) and (layer6_outputs(188));
    layer7_outputs(2416) <= not((layer6_outputs(3885)) xor (layer6_outputs(713)));
    layer7_outputs(2417) <= (layer6_outputs(4842)) xor (layer6_outputs(795));
    layer7_outputs(2418) <= not(layer6_outputs(4159));
    layer7_outputs(2419) <= (layer6_outputs(2694)) and not (layer6_outputs(2339));
    layer7_outputs(2420) <= layer6_outputs(3901);
    layer7_outputs(2421) <= (layer6_outputs(1430)) xor (layer6_outputs(2118));
    layer7_outputs(2422) <= not(layer6_outputs(2708));
    layer7_outputs(2423) <= (layer6_outputs(3217)) and (layer6_outputs(2417));
    layer7_outputs(2424) <= '1';
    layer7_outputs(2425) <= (layer6_outputs(4709)) and (layer6_outputs(3381));
    layer7_outputs(2426) <= layer6_outputs(2989);
    layer7_outputs(2427) <= not(layer6_outputs(2976));
    layer7_outputs(2428) <= not(layer6_outputs(2088));
    layer7_outputs(2429) <= not(layer6_outputs(558));
    layer7_outputs(2430) <= not(layer6_outputs(2119));
    layer7_outputs(2431) <= layer6_outputs(139);
    layer7_outputs(2432) <= not(layer6_outputs(2842));
    layer7_outputs(2433) <= not((layer6_outputs(1957)) xor (layer6_outputs(3001)));
    layer7_outputs(2434) <= not(layer6_outputs(2630));
    layer7_outputs(2435) <= (layer6_outputs(2648)) and (layer6_outputs(3000));
    layer7_outputs(2436) <= layer6_outputs(3892);
    layer7_outputs(2437) <= not(layer6_outputs(3548));
    layer7_outputs(2438) <= not(layer6_outputs(1666));
    layer7_outputs(2439) <= (layer6_outputs(1343)) or (layer6_outputs(3978));
    layer7_outputs(2440) <= not((layer6_outputs(494)) xor (layer6_outputs(2477)));
    layer7_outputs(2441) <= not(layer6_outputs(2800));
    layer7_outputs(2442) <= '0';
    layer7_outputs(2443) <= not((layer6_outputs(1239)) or (layer6_outputs(4657)));
    layer7_outputs(2444) <= layer6_outputs(3384);
    layer7_outputs(2445) <= not((layer6_outputs(964)) xor (layer6_outputs(4736)));
    layer7_outputs(2446) <= '0';
    layer7_outputs(2447) <= not(layer6_outputs(4562));
    layer7_outputs(2448) <= not(layer6_outputs(2991));
    layer7_outputs(2449) <= not((layer6_outputs(234)) xor (layer6_outputs(2485)));
    layer7_outputs(2450) <= (layer6_outputs(1485)) and not (layer6_outputs(3829));
    layer7_outputs(2451) <= (layer6_outputs(2295)) and not (layer6_outputs(4960));
    layer7_outputs(2452) <= layer6_outputs(4314);
    layer7_outputs(2453) <= not(layer6_outputs(1406));
    layer7_outputs(2454) <= (layer6_outputs(1973)) and not (layer6_outputs(290));
    layer7_outputs(2455) <= not(layer6_outputs(3229)) or (layer6_outputs(4441));
    layer7_outputs(2456) <= layer6_outputs(5105);
    layer7_outputs(2457) <= not(layer6_outputs(5003));
    layer7_outputs(2458) <= layer6_outputs(2836);
    layer7_outputs(2459) <= (layer6_outputs(3090)) or (layer6_outputs(348));
    layer7_outputs(2460) <= not(layer6_outputs(3919));
    layer7_outputs(2461) <= layer6_outputs(1992);
    layer7_outputs(2462) <= (layer6_outputs(98)) xor (layer6_outputs(5117));
    layer7_outputs(2463) <= (layer6_outputs(5119)) xor (layer6_outputs(2425));
    layer7_outputs(2464) <= not(layer6_outputs(702));
    layer7_outputs(2465) <= not(layer6_outputs(1334)) or (layer6_outputs(1791));
    layer7_outputs(2466) <= not(layer6_outputs(626));
    layer7_outputs(2467) <= not(layer6_outputs(1492));
    layer7_outputs(2468) <= not(layer6_outputs(2036));
    layer7_outputs(2469) <= '1';
    layer7_outputs(2470) <= not(layer6_outputs(479)) or (layer6_outputs(2068));
    layer7_outputs(2471) <= (layer6_outputs(4054)) or (layer6_outputs(3275));
    layer7_outputs(2472) <= (layer6_outputs(1287)) xor (layer6_outputs(2210));
    layer7_outputs(2473) <= not((layer6_outputs(2860)) and (layer6_outputs(4824)));
    layer7_outputs(2474) <= (layer6_outputs(1464)) and not (layer6_outputs(1692));
    layer7_outputs(2475) <= not(layer6_outputs(3211));
    layer7_outputs(2476) <= not((layer6_outputs(3340)) or (layer6_outputs(5049)));
    layer7_outputs(2477) <= not(layer6_outputs(3069));
    layer7_outputs(2478) <= not(layer6_outputs(829)) or (layer6_outputs(2016));
    layer7_outputs(2479) <= (layer6_outputs(1363)) and not (layer6_outputs(5100));
    layer7_outputs(2480) <= (layer6_outputs(2275)) and not (layer6_outputs(1095));
    layer7_outputs(2481) <= not((layer6_outputs(861)) xor (layer6_outputs(1304)));
    layer7_outputs(2482) <= '1';
    layer7_outputs(2483) <= not(layer6_outputs(4078));
    layer7_outputs(2484) <= not(layer6_outputs(2877)) or (layer6_outputs(2097));
    layer7_outputs(2485) <= '0';
    layer7_outputs(2486) <= not((layer6_outputs(178)) or (layer6_outputs(2352)));
    layer7_outputs(2487) <= not(layer6_outputs(1088));
    layer7_outputs(2488) <= (layer6_outputs(3891)) and not (layer6_outputs(4119));
    layer7_outputs(2489) <= (layer6_outputs(2864)) or (layer6_outputs(1729));
    layer7_outputs(2490) <= (layer6_outputs(800)) and not (layer6_outputs(4972));
    layer7_outputs(2491) <= not(layer6_outputs(4711)) or (layer6_outputs(2460));
    layer7_outputs(2492) <= not((layer6_outputs(1063)) and (layer6_outputs(1153)));
    layer7_outputs(2493) <= (layer6_outputs(4794)) and not (layer6_outputs(5101));
    layer7_outputs(2494) <= not((layer6_outputs(1154)) xor (layer6_outputs(4350)));
    layer7_outputs(2495) <= layer6_outputs(1087);
    layer7_outputs(2496) <= (layer6_outputs(3735)) and (layer6_outputs(4332));
    layer7_outputs(2497) <= '1';
    layer7_outputs(2498) <= not((layer6_outputs(1094)) xor (layer6_outputs(191)));
    layer7_outputs(2499) <= '0';
    layer7_outputs(2500) <= layer6_outputs(1922);
    layer7_outputs(2501) <= layer6_outputs(1954);
    layer7_outputs(2502) <= (layer6_outputs(2262)) and not (layer6_outputs(655));
    layer7_outputs(2503) <= not(layer6_outputs(4130)) or (layer6_outputs(3704));
    layer7_outputs(2504) <= (layer6_outputs(2825)) or (layer6_outputs(2476));
    layer7_outputs(2505) <= not(layer6_outputs(663)) or (layer6_outputs(4662));
    layer7_outputs(2506) <= layer6_outputs(272);
    layer7_outputs(2507) <= not(layer6_outputs(4929));
    layer7_outputs(2508) <= layer6_outputs(2665);
    layer7_outputs(2509) <= layer6_outputs(2208);
    layer7_outputs(2510) <= not(layer6_outputs(3974));
    layer7_outputs(2511) <= not(layer6_outputs(1531));
    layer7_outputs(2512) <= not(layer6_outputs(3768));
    layer7_outputs(2513) <= layer6_outputs(2248);
    layer7_outputs(2514) <= layer6_outputs(135);
    layer7_outputs(2515) <= (layer6_outputs(559)) or (layer6_outputs(2795));
    layer7_outputs(2516) <= not(layer6_outputs(3559));
    layer7_outputs(2517) <= layer6_outputs(555);
    layer7_outputs(2518) <= not((layer6_outputs(1824)) xor (layer6_outputs(1633)));
    layer7_outputs(2519) <= layer6_outputs(504);
    layer7_outputs(2520) <= (layer6_outputs(2431)) and (layer6_outputs(3823));
    layer7_outputs(2521) <= not((layer6_outputs(2787)) xor (layer6_outputs(66)));
    layer7_outputs(2522) <= layer6_outputs(3606);
    layer7_outputs(2523) <= not(layer6_outputs(1668));
    layer7_outputs(2524) <= not(layer6_outputs(3454));
    layer7_outputs(2525) <= not(layer6_outputs(184)) or (layer6_outputs(3106));
    layer7_outputs(2526) <= layer6_outputs(962);
    layer7_outputs(2527) <= (layer6_outputs(4614)) or (layer6_outputs(4105));
    layer7_outputs(2528) <= (layer6_outputs(2037)) and not (layer6_outputs(3041));
    layer7_outputs(2529) <= not(layer6_outputs(3049)) or (layer6_outputs(1196));
    layer7_outputs(2530) <= layer6_outputs(4505);
    layer7_outputs(2531) <= layer6_outputs(3145);
    layer7_outputs(2532) <= not(layer6_outputs(1630));
    layer7_outputs(2533) <= layer6_outputs(5108);
    layer7_outputs(2534) <= not((layer6_outputs(4536)) and (layer6_outputs(1592)));
    layer7_outputs(2535) <= not((layer6_outputs(2015)) xor (layer6_outputs(273)));
    layer7_outputs(2536) <= (layer6_outputs(2984)) xor (layer6_outputs(1373));
    layer7_outputs(2537) <= not(layer6_outputs(369));
    layer7_outputs(2538) <= layer6_outputs(3256);
    layer7_outputs(2539) <= (layer6_outputs(4516)) xor (layer6_outputs(4143));
    layer7_outputs(2540) <= layer6_outputs(2573);
    layer7_outputs(2541) <= not(layer6_outputs(3237));
    layer7_outputs(2542) <= '1';
    layer7_outputs(2543) <= (layer6_outputs(4732)) and not (layer6_outputs(2071));
    layer7_outputs(2544) <= not((layer6_outputs(1425)) and (layer6_outputs(4328)));
    layer7_outputs(2545) <= not((layer6_outputs(3772)) xor (layer6_outputs(4245)));
    layer7_outputs(2546) <= layer6_outputs(2019);
    layer7_outputs(2547) <= not(layer6_outputs(924)) or (layer6_outputs(5064));
    layer7_outputs(2548) <= not(layer6_outputs(173));
    layer7_outputs(2549) <= layer6_outputs(3751);
    layer7_outputs(2550) <= (layer6_outputs(1385)) or (layer6_outputs(2401));
    layer7_outputs(2551) <= layer6_outputs(686);
    layer7_outputs(2552) <= (layer6_outputs(3)) and not (layer6_outputs(345));
    layer7_outputs(2553) <= layer6_outputs(3417);
    layer7_outputs(2554) <= (layer6_outputs(1099)) and not (layer6_outputs(1558));
    layer7_outputs(2555) <= not((layer6_outputs(122)) xor (layer6_outputs(3010)));
    layer7_outputs(2556) <= layer6_outputs(3524);
    layer7_outputs(2557) <= not((layer6_outputs(2908)) xor (layer6_outputs(4987)));
    layer7_outputs(2558) <= not(layer6_outputs(69));
    layer7_outputs(2559) <= (layer6_outputs(2134)) xor (layer6_outputs(2495));
    layer7_outputs(2560) <= layer6_outputs(4084);
    layer7_outputs(2561) <= not(layer6_outputs(2701)) or (layer6_outputs(2545));
    layer7_outputs(2562) <= (layer6_outputs(1967)) and not (layer6_outputs(1985));
    layer7_outputs(2563) <= (layer6_outputs(1961)) or (layer6_outputs(1853));
    layer7_outputs(2564) <= (layer6_outputs(151)) xor (layer6_outputs(2845));
    layer7_outputs(2565) <= layer6_outputs(3188);
    layer7_outputs(2566) <= layer6_outputs(1797);
    layer7_outputs(2567) <= (layer6_outputs(1081)) or (layer6_outputs(3089));
    layer7_outputs(2568) <= not(layer6_outputs(1757));
    layer7_outputs(2569) <= not(layer6_outputs(356)) or (layer6_outputs(5097));
    layer7_outputs(2570) <= (layer6_outputs(1979)) xor (layer6_outputs(4135));
    layer7_outputs(2571) <= (layer6_outputs(4019)) xor (layer6_outputs(4439));
    layer7_outputs(2572) <= '1';
    layer7_outputs(2573) <= layer6_outputs(1314);
    layer7_outputs(2574) <= not(layer6_outputs(3394));
    layer7_outputs(2575) <= not(layer6_outputs(624));
    layer7_outputs(2576) <= layer6_outputs(892);
    layer7_outputs(2577) <= layer6_outputs(3446);
    layer7_outputs(2578) <= layer6_outputs(2185);
    layer7_outputs(2579) <= layer6_outputs(1877);
    layer7_outputs(2580) <= layer6_outputs(1964);
    layer7_outputs(2581) <= not(layer6_outputs(4678));
    layer7_outputs(2582) <= layer6_outputs(4012);
    layer7_outputs(2583) <= layer6_outputs(488);
    layer7_outputs(2584) <= layer6_outputs(2523);
    layer7_outputs(2585) <= not((layer6_outputs(4163)) or (layer6_outputs(299)));
    layer7_outputs(2586) <= layer6_outputs(4164);
    layer7_outputs(2587) <= (layer6_outputs(1879)) xor (layer6_outputs(3110));
    layer7_outputs(2588) <= not(layer6_outputs(787));
    layer7_outputs(2589) <= not((layer6_outputs(4031)) and (layer6_outputs(2485)));
    layer7_outputs(2590) <= layer6_outputs(1718);
    layer7_outputs(2591) <= not(layer6_outputs(4897));
    layer7_outputs(2592) <= not(layer6_outputs(276));
    layer7_outputs(2593) <= (layer6_outputs(884)) xor (layer6_outputs(1906));
    layer7_outputs(2594) <= not((layer6_outputs(3229)) and (layer6_outputs(4778)));
    layer7_outputs(2595) <= not(layer6_outputs(3461));
    layer7_outputs(2596) <= (layer6_outputs(4831)) and not (layer6_outputs(1921));
    layer7_outputs(2597) <= layer6_outputs(3942);
    layer7_outputs(2598) <= layer6_outputs(3605);
    layer7_outputs(2599) <= (layer6_outputs(3925)) and not (layer6_outputs(2920));
    layer7_outputs(2600) <= not(layer6_outputs(3403));
    layer7_outputs(2601) <= layer6_outputs(4512);
    layer7_outputs(2602) <= layer6_outputs(4513);
    layer7_outputs(2603) <= not((layer6_outputs(492)) xor (layer6_outputs(1369)));
    layer7_outputs(2604) <= not(layer6_outputs(3793));
    layer7_outputs(2605) <= layer6_outputs(45);
    layer7_outputs(2606) <= not(layer6_outputs(4167));
    layer7_outputs(2607) <= '0';
    layer7_outputs(2608) <= not((layer6_outputs(511)) and (layer6_outputs(1797)));
    layer7_outputs(2609) <= layer6_outputs(3425);
    layer7_outputs(2610) <= not(layer6_outputs(3178));
    layer7_outputs(2611) <= not(layer6_outputs(4514));
    layer7_outputs(2612) <= not(layer6_outputs(1308)) or (layer6_outputs(2213));
    layer7_outputs(2613) <= (layer6_outputs(2537)) and (layer6_outputs(192));
    layer7_outputs(2614) <= '1';
    layer7_outputs(2615) <= (layer6_outputs(4401)) or (layer6_outputs(2154));
    layer7_outputs(2616) <= layer6_outputs(4265);
    layer7_outputs(2617) <= layer6_outputs(273);
    layer7_outputs(2618) <= not(layer6_outputs(491));
    layer7_outputs(2619) <= layer6_outputs(554);
    layer7_outputs(2620) <= layer6_outputs(3644);
    layer7_outputs(2621) <= layer6_outputs(4837);
    layer7_outputs(2622) <= (layer6_outputs(1283)) and not (layer6_outputs(620));
    layer7_outputs(2623) <= not((layer6_outputs(3021)) xor (layer6_outputs(138)));
    layer7_outputs(2624) <= (layer6_outputs(2075)) xor (layer6_outputs(1837));
    layer7_outputs(2625) <= (layer6_outputs(3105)) and (layer6_outputs(1188));
    layer7_outputs(2626) <= not(layer6_outputs(3660)) or (layer6_outputs(4101));
    layer7_outputs(2627) <= layer6_outputs(641);
    layer7_outputs(2628) <= (layer6_outputs(4821)) or (layer6_outputs(904));
    layer7_outputs(2629) <= not((layer6_outputs(4542)) xor (layer6_outputs(3193)));
    layer7_outputs(2630) <= not(layer6_outputs(2906));
    layer7_outputs(2631) <= not(layer6_outputs(4316));
    layer7_outputs(2632) <= (layer6_outputs(92)) and not (layer6_outputs(2055));
    layer7_outputs(2633) <= not(layer6_outputs(2839));
    layer7_outputs(2634) <= (layer6_outputs(4161)) and not (layer6_outputs(1615));
    layer7_outputs(2635) <= not((layer6_outputs(4345)) and (layer6_outputs(503)));
    layer7_outputs(2636) <= layer6_outputs(2697);
    layer7_outputs(2637) <= not(layer6_outputs(4275));
    layer7_outputs(2638) <= not(layer6_outputs(189));
    layer7_outputs(2639) <= (layer6_outputs(249)) and not (layer6_outputs(2776));
    layer7_outputs(2640) <= not((layer6_outputs(2656)) xor (layer6_outputs(1428)));
    layer7_outputs(2641) <= (layer6_outputs(601)) or (layer6_outputs(4885));
    layer7_outputs(2642) <= layer6_outputs(522);
    layer7_outputs(2643) <= layer6_outputs(4916);
    layer7_outputs(2644) <= not(layer6_outputs(4664));
    layer7_outputs(2645) <= (layer6_outputs(2257)) xor (layer6_outputs(3871));
    layer7_outputs(2646) <= layer6_outputs(4541);
    layer7_outputs(2647) <= layer6_outputs(4726);
    layer7_outputs(2648) <= not(layer6_outputs(4006));
    layer7_outputs(2649) <= not(layer6_outputs(685));
    layer7_outputs(2650) <= layer6_outputs(2174);
    layer7_outputs(2651) <= not(layer6_outputs(3821));
    layer7_outputs(2652) <= not(layer6_outputs(3292));
    layer7_outputs(2653) <= not(layer6_outputs(1751));
    layer7_outputs(2654) <= not(layer6_outputs(4435));
    layer7_outputs(2655) <= layer6_outputs(4615);
    layer7_outputs(2656) <= not(layer6_outputs(1696));
    layer7_outputs(2657) <= not((layer6_outputs(975)) and (layer6_outputs(259)));
    layer7_outputs(2658) <= not((layer6_outputs(2989)) xor (layer6_outputs(3243)));
    layer7_outputs(2659) <= not(layer6_outputs(586)) or (layer6_outputs(4154));
    layer7_outputs(2660) <= not(layer6_outputs(2514));
    layer7_outputs(2661) <= (layer6_outputs(669)) and not (layer6_outputs(4436));
    layer7_outputs(2662) <= (layer6_outputs(665)) and not (layer6_outputs(4778));
    layer7_outputs(2663) <= layer6_outputs(139);
    layer7_outputs(2664) <= not((layer6_outputs(1903)) and (layer6_outputs(2003)));
    layer7_outputs(2665) <= not(layer6_outputs(200));
    layer7_outputs(2666) <= not((layer6_outputs(3829)) or (layer6_outputs(3746)));
    layer7_outputs(2667) <= (layer6_outputs(4620)) and (layer6_outputs(210));
    layer7_outputs(2668) <= not((layer6_outputs(5063)) xor (layer6_outputs(429)));
    layer7_outputs(2669) <= (layer6_outputs(2038)) and not (layer6_outputs(2012));
    layer7_outputs(2670) <= not(layer6_outputs(4017));
    layer7_outputs(2671) <= '0';
    layer7_outputs(2672) <= (layer6_outputs(3982)) or (layer6_outputs(1977));
    layer7_outputs(2673) <= not(layer6_outputs(796));
    layer7_outputs(2674) <= (layer6_outputs(3803)) or (layer6_outputs(2322));
    layer7_outputs(2675) <= not((layer6_outputs(4018)) or (layer6_outputs(3489)));
    layer7_outputs(2676) <= (layer6_outputs(876)) and not (layer6_outputs(1688));
    layer7_outputs(2677) <= not((layer6_outputs(3934)) and (layer6_outputs(4924)));
    layer7_outputs(2678) <= not(layer6_outputs(2785));
    layer7_outputs(2679) <= layer6_outputs(2961);
    layer7_outputs(2680) <= not((layer6_outputs(2053)) or (layer6_outputs(801)));
    layer7_outputs(2681) <= (layer6_outputs(1172)) and not (layer6_outputs(4165));
    layer7_outputs(2682) <= (layer6_outputs(213)) and (layer6_outputs(1105));
    layer7_outputs(2683) <= layer6_outputs(1400);
    layer7_outputs(2684) <= not(layer6_outputs(3859));
    layer7_outputs(2685) <= not(layer6_outputs(1245)) or (layer6_outputs(3391));
    layer7_outputs(2686) <= layer6_outputs(3524);
    layer7_outputs(2687) <= not(layer6_outputs(3497));
    layer7_outputs(2688) <= not(layer6_outputs(3172));
    layer7_outputs(2689) <= not(layer6_outputs(3272));
    layer7_outputs(2690) <= layer6_outputs(3278);
    layer7_outputs(2691) <= layer6_outputs(417);
    layer7_outputs(2692) <= not(layer6_outputs(1718));
    layer7_outputs(2693) <= not(layer6_outputs(3615)) or (layer6_outputs(4000));
    layer7_outputs(2694) <= not(layer6_outputs(4197)) or (layer6_outputs(3307));
    layer7_outputs(2695) <= not(layer6_outputs(4302)) or (layer6_outputs(3772));
    layer7_outputs(2696) <= not((layer6_outputs(4531)) xor (layer6_outputs(3474)));
    layer7_outputs(2697) <= not(layer6_outputs(3511)) or (layer6_outputs(4368));
    layer7_outputs(2698) <= not(layer6_outputs(4471));
    layer7_outputs(2699) <= not(layer6_outputs(872));
    layer7_outputs(2700) <= layer6_outputs(2507);
    layer7_outputs(2701) <= layer6_outputs(2703);
    layer7_outputs(2702) <= not(layer6_outputs(4346));
    layer7_outputs(2703) <= not(layer6_outputs(855));
    layer7_outputs(2704) <= not(layer6_outputs(1189));
    layer7_outputs(2705) <= not(layer6_outputs(4078));
    layer7_outputs(2706) <= not((layer6_outputs(2557)) xor (layer6_outputs(4056)));
    layer7_outputs(2707) <= (layer6_outputs(3019)) and (layer6_outputs(2539));
    layer7_outputs(2708) <= layer6_outputs(4060);
    layer7_outputs(2709) <= (layer6_outputs(2794)) and not (layer6_outputs(93));
    layer7_outputs(2710) <= not(layer6_outputs(3092));
    layer7_outputs(2711) <= (layer6_outputs(3626)) or (layer6_outputs(4732));
    layer7_outputs(2712) <= not(layer6_outputs(1516));
    layer7_outputs(2713) <= '1';
    layer7_outputs(2714) <= not(layer6_outputs(1375)) or (layer6_outputs(2064));
    layer7_outputs(2715) <= not((layer6_outputs(2185)) xor (layer6_outputs(96)));
    layer7_outputs(2716) <= not(layer6_outputs(1455));
    layer7_outputs(2717) <= not((layer6_outputs(1646)) xor (layer6_outputs(5114)));
    layer7_outputs(2718) <= layer6_outputs(4848);
    layer7_outputs(2719) <= not(layer6_outputs(4183)) or (layer6_outputs(1967));
    layer7_outputs(2720) <= not(layer6_outputs(2360));
    layer7_outputs(2721) <= (layer6_outputs(2299)) and not (layer6_outputs(174));
    layer7_outputs(2722) <= (layer6_outputs(2847)) and not (layer6_outputs(2778));
    layer7_outputs(2723) <= layer6_outputs(3321);
    layer7_outputs(2724) <= layer6_outputs(4197);
    layer7_outputs(2725) <= (layer6_outputs(351)) xor (layer6_outputs(3783));
    layer7_outputs(2726) <= not(layer6_outputs(364));
    layer7_outputs(2727) <= (layer6_outputs(3689)) xor (layer6_outputs(2879));
    layer7_outputs(2728) <= not(layer6_outputs(3721)) or (layer6_outputs(188));
    layer7_outputs(2729) <= not(layer6_outputs(1573));
    layer7_outputs(2730) <= (layer6_outputs(2221)) xor (layer6_outputs(3342));
    layer7_outputs(2731) <= layer6_outputs(2982);
    layer7_outputs(2732) <= layer6_outputs(592);
    layer7_outputs(2733) <= (layer6_outputs(294)) and not (layer6_outputs(4480));
    layer7_outputs(2734) <= '0';
    layer7_outputs(2735) <= not(layer6_outputs(3570));
    layer7_outputs(2736) <= not(layer6_outputs(88));
    layer7_outputs(2737) <= (layer6_outputs(1756)) and not (layer6_outputs(2793));
    layer7_outputs(2738) <= not(layer6_outputs(1262));
    layer7_outputs(2739) <= layer6_outputs(4671);
    layer7_outputs(2740) <= not(layer6_outputs(938));
    layer7_outputs(2741) <= layer6_outputs(3703);
    layer7_outputs(2742) <= not((layer6_outputs(3184)) xor (layer6_outputs(3766)));
    layer7_outputs(2743) <= (layer6_outputs(1203)) or (layer6_outputs(1887));
    layer7_outputs(2744) <= not(layer6_outputs(2962));
    layer7_outputs(2745) <= layer6_outputs(3043);
    layer7_outputs(2746) <= not(layer6_outputs(2001)) or (layer6_outputs(1156));
    layer7_outputs(2747) <= not((layer6_outputs(369)) xor (layer6_outputs(4793)));
    layer7_outputs(2748) <= (layer6_outputs(287)) and not (layer6_outputs(229));
    layer7_outputs(2749) <= (layer6_outputs(4106)) and not (layer6_outputs(1981));
    layer7_outputs(2750) <= layer6_outputs(859);
    layer7_outputs(2751) <= (layer6_outputs(2116)) xor (layer6_outputs(4107));
    layer7_outputs(2752) <= not(layer6_outputs(2058));
    layer7_outputs(2753) <= not((layer6_outputs(3005)) xor (layer6_outputs(3475)));
    layer7_outputs(2754) <= layer6_outputs(3691);
    layer7_outputs(2755) <= not(layer6_outputs(4196));
    layer7_outputs(2756) <= (layer6_outputs(3471)) xor (layer6_outputs(42));
    layer7_outputs(2757) <= (layer6_outputs(1023)) xor (layer6_outputs(630));
    layer7_outputs(2758) <= not((layer6_outputs(4317)) or (layer6_outputs(2741)));
    layer7_outputs(2759) <= not(layer6_outputs(1143));
    layer7_outputs(2760) <= layer6_outputs(1146);
    layer7_outputs(2761) <= not((layer6_outputs(4728)) and (layer6_outputs(4375)));
    layer7_outputs(2762) <= not(layer6_outputs(3261));
    layer7_outputs(2763) <= (layer6_outputs(4603)) and not (layer6_outputs(300));
    layer7_outputs(2764) <= not((layer6_outputs(1128)) xor (layer6_outputs(561)));
    layer7_outputs(2765) <= not((layer6_outputs(3711)) or (layer6_outputs(2263)));
    layer7_outputs(2766) <= not(layer6_outputs(3745));
    layer7_outputs(2767) <= '1';
    layer7_outputs(2768) <= (layer6_outputs(3284)) or (layer6_outputs(3979));
    layer7_outputs(2769) <= not(layer6_outputs(5112));
    layer7_outputs(2770) <= not(layer6_outputs(4992)) or (layer6_outputs(810));
    layer7_outputs(2771) <= layer6_outputs(1684);
    layer7_outputs(2772) <= not((layer6_outputs(3696)) xor (layer6_outputs(1635)));
    layer7_outputs(2773) <= layer6_outputs(3095);
    layer7_outputs(2774) <= not(layer6_outputs(3013));
    layer7_outputs(2775) <= not(layer6_outputs(23)) or (layer6_outputs(2016));
    layer7_outputs(2776) <= not((layer6_outputs(2133)) and (layer6_outputs(5077)));
    layer7_outputs(2777) <= not(layer6_outputs(1077)) or (layer6_outputs(2965));
    layer7_outputs(2778) <= not((layer6_outputs(673)) or (layer6_outputs(1862)));
    layer7_outputs(2779) <= not(layer6_outputs(3844));
    layer7_outputs(2780) <= layer6_outputs(4216);
    layer7_outputs(2781) <= layer6_outputs(1726);
    layer7_outputs(2782) <= (layer6_outputs(2240)) or (layer6_outputs(4719));
    layer7_outputs(2783) <= not((layer6_outputs(1917)) or (layer6_outputs(1003)));
    layer7_outputs(2784) <= not(layer6_outputs(1330));
    layer7_outputs(2785) <= not((layer6_outputs(241)) xor (layer6_outputs(4053)));
    layer7_outputs(2786) <= '1';
    layer7_outputs(2787) <= not(layer6_outputs(3903));
    layer7_outputs(2788) <= layer6_outputs(5085);
    layer7_outputs(2789) <= (layer6_outputs(885)) or (layer6_outputs(3118));
    layer7_outputs(2790) <= not(layer6_outputs(3794));
    layer7_outputs(2791) <= layer6_outputs(1347);
    layer7_outputs(2792) <= (layer6_outputs(1960)) xor (layer6_outputs(437));
    layer7_outputs(2793) <= not(layer6_outputs(2895)) or (layer6_outputs(4201));
    layer7_outputs(2794) <= not((layer6_outputs(4567)) and (layer6_outputs(1186)));
    layer7_outputs(2795) <= layer6_outputs(891);
    layer7_outputs(2796) <= layer6_outputs(3464);
    layer7_outputs(2797) <= not((layer6_outputs(3916)) or (layer6_outputs(2442)));
    layer7_outputs(2798) <= layer6_outputs(2791);
    layer7_outputs(2799) <= (layer6_outputs(1400)) and not (layer6_outputs(3078));
    layer7_outputs(2800) <= not(layer6_outputs(2111));
    layer7_outputs(2801) <= not(layer6_outputs(437));
    layer7_outputs(2802) <= not((layer6_outputs(43)) xor (layer6_outputs(206)));
    layer7_outputs(2803) <= (layer6_outputs(2452)) and (layer6_outputs(3167));
    layer7_outputs(2804) <= not(layer6_outputs(4028));
    layer7_outputs(2805) <= (layer6_outputs(3004)) and not (layer6_outputs(2450));
    layer7_outputs(2806) <= not(layer6_outputs(2779));
    layer7_outputs(2807) <= not(layer6_outputs(3414));
    layer7_outputs(2808) <= not(layer6_outputs(4412));
    layer7_outputs(2809) <= layer6_outputs(2457);
    layer7_outputs(2810) <= (layer6_outputs(3299)) xor (layer6_outputs(2073));
    layer7_outputs(2811) <= not(layer6_outputs(2458));
    layer7_outputs(2812) <= layer6_outputs(2990);
    layer7_outputs(2813) <= not((layer6_outputs(4096)) and (layer6_outputs(4995)));
    layer7_outputs(2814) <= (layer6_outputs(3359)) xor (layer6_outputs(1015));
    layer7_outputs(2815) <= not(layer6_outputs(278)) or (layer6_outputs(978));
    layer7_outputs(2816) <= (layer6_outputs(2321)) and (layer6_outputs(3771));
    layer7_outputs(2817) <= layer6_outputs(1353);
    layer7_outputs(2818) <= not(layer6_outputs(464));
    layer7_outputs(2819) <= layer6_outputs(2621);
    layer7_outputs(2820) <= layer6_outputs(1839);
    layer7_outputs(2821) <= not(layer6_outputs(1537));
    layer7_outputs(2822) <= not(layer6_outputs(3577));
    layer7_outputs(2823) <= (layer6_outputs(2436)) and not (layer6_outputs(1614));
    layer7_outputs(2824) <= not(layer6_outputs(3684)) or (layer6_outputs(2966));
    layer7_outputs(2825) <= not(layer6_outputs(5109));
    layer7_outputs(2826) <= layer6_outputs(2809);
    layer7_outputs(2827) <= layer6_outputs(1414);
    layer7_outputs(2828) <= not(layer6_outputs(403));
    layer7_outputs(2829) <= not(layer6_outputs(4549));
    layer7_outputs(2830) <= not((layer6_outputs(346)) and (layer6_outputs(623)));
    layer7_outputs(2831) <= not((layer6_outputs(5042)) and (layer6_outputs(2713)));
    layer7_outputs(2832) <= layer6_outputs(2276);
    layer7_outputs(2833) <= layer6_outputs(1438);
    layer7_outputs(2834) <= not(layer6_outputs(4629)) or (layer6_outputs(2925));
    layer7_outputs(2835) <= (layer6_outputs(333)) and (layer6_outputs(3793));
    layer7_outputs(2836) <= not((layer6_outputs(2722)) xor (layer6_outputs(2841)));
    layer7_outputs(2837) <= not(layer6_outputs(4192));
    layer7_outputs(2838) <= (layer6_outputs(2045)) or (layer6_outputs(3205));
    layer7_outputs(2839) <= not(layer6_outputs(908)) or (layer6_outputs(3154));
    layer7_outputs(2840) <= (layer6_outputs(3618)) and not (layer6_outputs(1926));
    layer7_outputs(2841) <= layer6_outputs(2950);
    layer7_outputs(2842) <= not(layer6_outputs(1528));
    layer7_outputs(2843) <= (layer6_outputs(889)) and not (layer6_outputs(25));
    layer7_outputs(2844) <= layer6_outputs(902);
    layer7_outputs(2845) <= layer6_outputs(1843);
    layer7_outputs(2846) <= not(layer6_outputs(1527));
    layer7_outputs(2847) <= not(layer6_outputs(1163));
    layer7_outputs(2848) <= layer6_outputs(1067);
    layer7_outputs(2849) <= layer6_outputs(3438);
    layer7_outputs(2850) <= (layer6_outputs(1971)) xor (layer6_outputs(419));
    layer7_outputs(2851) <= not(layer6_outputs(3131));
    layer7_outputs(2852) <= not(layer6_outputs(283)) or (layer6_outputs(3390));
    layer7_outputs(2853) <= layer6_outputs(1155);
    layer7_outputs(2854) <= layer6_outputs(4630);
    layer7_outputs(2855) <= not(layer6_outputs(4962)) or (layer6_outputs(2349));
    layer7_outputs(2856) <= layer6_outputs(2319);
    layer7_outputs(2857) <= not(layer6_outputs(1016));
    layer7_outputs(2858) <= not(layer6_outputs(4915));
    layer7_outputs(2859) <= not((layer6_outputs(3828)) or (layer6_outputs(2949)));
    layer7_outputs(2860) <= not(layer6_outputs(1548));
    layer7_outputs(2861) <= '1';
    layer7_outputs(2862) <= not((layer6_outputs(3701)) and (layer6_outputs(1106)));
    layer7_outputs(2863) <= not(layer6_outputs(1751));
    layer7_outputs(2864) <= layer6_outputs(2261);
    layer7_outputs(2865) <= layer6_outputs(4126);
    layer7_outputs(2866) <= (layer6_outputs(722)) and not (layer6_outputs(3022));
    layer7_outputs(2867) <= not(layer6_outputs(146));
    layer7_outputs(2868) <= layer6_outputs(1598);
    layer7_outputs(2869) <= (layer6_outputs(1192)) and (layer6_outputs(1178));
    layer7_outputs(2870) <= not(layer6_outputs(4031)) or (layer6_outputs(1802));
    layer7_outputs(2871) <= not(layer6_outputs(599));
    layer7_outputs(2872) <= not((layer6_outputs(1603)) and (layer6_outputs(1224)));
    layer7_outputs(2873) <= (layer6_outputs(243)) and not (layer6_outputs(1639));
    layer7_outputs(2874) <= not((layer6_outputs(2440)) and (layer6_outputs(1510)));
    layer7_outputs(2875) <= not(layer6_outputs(1405)) or (layer6_outputs(2875));
    layer7_outputs(2876) <= '1';
    layer7_outputs(2877) <= (layer6_outputs(4946)) or (layer6_outputs(1957));
    layer7_outputs(2878) <= layer6_outputs(1334);
    layer7_outputs(2879) <= (layer6_outputs(2198)) or (layer6_outputs(4288));
    layer7_outputs(2880) <= (layer6_outputs(700)) and not (layer6_outputs(4783));
    layer7_outputs(2881) <= not((layer6_outputs(2897)) and (layer6_outputs(2022)));
    layer7_outputs(2882) <= (layer6_outputs(1032)) and (layer6_outputs(4849));
    layer7_outputs(2883) <= not(layer6_outputs(4885));
    layer7_outputs(2884) <= not(layer6_outputs(2491)) or (layer6_outputs(1285));
    layer7_outputs(2885) <= not(layer6_outputs(3912));
    layer7_outputs(2886) <= (layer6_outputs(4869)) or (layer6_outputs(1487));
    layer7_outputs(2887) <= (layer6_outputs(4331)) and not (layer6_outputs(1489));
    layer7_outputs(2888) <= not((layer6_outputs(3788)) xor (layer6_outputs(2801)));
    layer7_outputs(2889) <= layer6_outputs(3958);
    layer7_outputs(2890) <= not(layer6_outputs(3530));
    layer7_outputs(2891) <= (layer6_outputs(1697)) xor (layer6_outputs(2585));
    layer7_outputs(2892) <= layer6_outputs(2803);
    layer7_outputs(2893) <= layer6_outputs(3568);
    layer7_outputs(2894) <= not(layer6_outputs(1126));
    layer7_outputs(2895) <= not(layer6_outputs(2326)) or (layer6_outputs(3072));
    layer7_outputs(2896) <= layer6_outputs(1033);
    layer7_outputs(2897) <= (layer6_outputs(1686)) and (layer6_outputs(2324));
    layer7_outputs(2898) <= not(layer6_outputs(2074));
    layer7_outputs(2899) <= (layer6_outputs(1109)) and (layer6_outputs(1402));
    layer7_outputs(2900) <= not(layer6_outputs(170));
    layer7_outputs(2901) <= (layer6_outputs(104)) and not (layer6_outputs(1579));
    layer7_outputs(2902) <= (layer6_outputs(1515)) and not (layer6_outputs(1928));
    layer7_outputs(2903) <= not(layer6_outputs(1053));
    layer7_outputs(2904) <= layer6_outputs(966);
    layer7_outputs(2905) <= not(layer6_outputs(3693)) or (layer6_outputs(1995));
    layer7_outputs(2906) <= not(layer6_outputs(3133));
    layer7_outputs(2907) <= not(layer6_outputs(1035));
    layer7_outputs(2908) <= not((layer6_outputs(2192)) xor (layer6_outputs(2469)));
    layer7_outputs(2909) <= layer6_outputs(4989);
    layer7_outputs(2910) <= not(layer6_outputs(4667));
    layer7_outputs(2911) <= layer6_outputs(4463);
    layer7_outputs(2912) <= not(layer6_outputs(1062));
    layer7_outputs(2913) <= not((layer6_outputs(1730)) and (layer6_outputs(4488)));
    layer7_outputs(2914) <= not(layer6_outputs(4502));
    layer7_outputs(2915) <= (layer6_outputs(2066)) or (layer6_outputs(4648));
    layer7_outputs(2916) <= not(layer6_outputs(2007));
    layer7_outputs(2917) <= not(layer6_outputs(1474));
    layer7_outputs(2918) <= not((layer6_outputs(4703)) and (layer6_outputs(4033)));
    layer7_outputs(2919) <= (layer6_outputs(261)) and not (layer6_outputs(3032));
    layer7_outputs(2920) <= layer6_outputs(2962);
    layer7_outputs(2921) <= not((layer6_outputs(4061)) or (layer6_outputs(2134)));
    layer7_outputs(2922) <= (layer6_outputs(2092)) and (layer6_outputs(493));
    layer7_outputs(2923) <= not(layer6_outputs(1301));
    layer7_outputs(2924) <= not(layer6_outputs(681));
    layer7_outputs(2925) <= layer6_outputs(2764);
    layer7_outputs(2926) <= (layer6_outputs(2757)) xor (layer6_outputs(4663));
    layer7_outputs(2927) <= not(layer6_outputs(3950)) or (layer6_outputs(3629));
    layer7_outputs(2928) <= not((layer6_outputs(4392)) xor (layer6_outputs(2348)));
    layer7_outputs(2929) <= layer6_outputs(4464);
    layer7_outputs(2930) <= not(layer6_outputs(4336));
    layer7_outputs(2931) <= layer6_outputs(341);
    layer7_outputs(2932) <= not((layer6_outputs(1474)) and (layer6_outputs(2157)));
    layer7_outputs(2933) <= (layer6_outputs(3964)) and not (layer6_outputs(3227));
    layer7_outputs(2934) <= not((layer6_outputs(2751)) or (layer6_outputs(153)));
    layer7_outputs(2935) <= layer6_outputs(3409);
    layer7_outputs(2936) <= not(layer6_outputs(2082));
    layer7_outputs(2937) <= layer6_outputs(807);
    layer7_outputs(2938) <= layer6_outputs(2814);
    layer7_outputs(2939) <= (layer6_outputs(366)) xor (layer6_outputs(897));
    layer7_outputs(2940) <= not(layer6_outputs(5081));
    layer7_outputs(2941) <= not(layer6_outputs(3813));
    layer7_outputs(2942) <= not((layer6_outputs(462)) or (layer6_outputs(1490)));
    layer7_outputs(2943) <= not(layer6_outputs(2072));
    layer7_outputs(2944) <= not(layer6_outputs(877)) or (layer6_outputs(2803));
    layer7_outputs(2945) <= not(layer6_outputs(2388));
    layer7_outputs(2946) <= not((layer6_outputs(1132)) or (layer6_outputs(29)));
    layer7_outputs(2947) <= not(layer6_outputs(621));
    layer7_outputs(2948) <= (layer6_outputs(4221)) and (layer6_outputs(631));
    layer7_outputs(2949) <= not((layer6_outputs(2298)) or (layer6_outputs(4386)));
    layer7_outputs(2950) <= not((layer6_outputs(3719)) xor (layer6_outputs(4702)));
    layer7_outputs(2951) <= (layer6_outputs(478)) xor (layer6_outputs(2280));
    layer7_outputs(2952) <= layer6_outputs(4390);
    layer7_outputs(2953) <= layer6_outputs(2049);
    layer7_outputs(2954) <= layer6_outputs(3039);
    layer7_outputs(2955) <= layer6_outputs(1096);
    layer7_outputs(2956) <= layer6_outputs(3245);
    layer7_outputs(2957) <= not((layer6_outputs(584)) xor (layer6_outputs(1699)));
    layer7_outputs(2958) <= not(layer6_outputs(4211));
    layer7_outputs(2959) <= (layer6_outputs(4302)) xor (layer6_outputs(366));
    layer7_outputs(2960) <= not((layer6_outputs(3244)) and (layer6_outputs(3672)));
    layer7_outputs(2961) <= layer6_outputs(2264);
    layer7_outputs(2962) <= not((layer6_outputs(4492)) xor (layer6_outputs(2224)));
    layer7_outputs(2963) <= not((layer6_outputs(1783)) or (layer6_outputs(1172)));
    layer7_outputs(2964) <= not((layer6_outputs(2014)) or (layer6_outputs(2626)));
    layer7_outputs(2965) <= (layer6_outputs(3098)) and not (layer6_outputs(2490));
    layer7_outputs(2966) <= layer6_outputs(2083);
    layer7_outputs(2967) <= not(layer6_outputs(2403));
    layer7_outputs(2968) <= not(layer6_outputs(3729));
    layer7_outputs(2969) <= not((layer6_outputs(3667)) xor (layer6_outputs(3287)));
    layer7_outputs(2970) <= not(layer6_outputs(2776));
    layer7_outputs(2971) <= not(layer6_outputs(1567)) or (layer6_outputs(4729));
    layer7_outputs(2972) <= (layer6_outputs(4514)) and (layer6_outputs(643));
    layer7_outputs(2973) <= (layer6_outputs(114)) xor (layer6_outputs(4287));
    layer7_outputs(2974) <= not(layer6_outputs(3088)) or (layer6_outputs(3866));
    layer7_outputs(2975) <= layer6_outputs(5033);
    layer7_outputs(2976) <= not(layer6_outputs(730)) or (layer6_outputs(2244));
    layer7_outputs(2977) <= not(layer6_outputs(2029)) or (layer6_outputs(2023));
    layer7_outputs(2978) <= (layer6_outputs(1164)) and not (layer6_outputs(990));
    layer7_outputs(2979) <= not(layer6_outputs(2472));
    layer7_outputs(2980) <= not((layer6_outputs(4540)) and (layer6_outputs(1867)));
    layer7_outputs(2981) <= layer6_outputs(1263);
    layer7_outputs(2982) <= not(layer6_outputs(3609));
    layer7_outputs(2983) <= not((layer6_outputs(3370)) xor (layer6_outputs(2751)));
    layer7_outputs(2984) <= (layer6_outputs(1131)) and not (layer6_outputs(653));
    layer7_outputs(2985) <= (layer6_outputs(1805)) xor (layer6_outputs(4438));
    layer7_outputs(2986) <= layer6_outputs(4748);
    layer7_outputs(2987) <= (layer6_outputs(2343)) and not (layer6_outputs(616));
    layer7_outputs(2988) <= not((layer6_outputs(4246)) xor (layer6_outputs(4108)));
    layer7_outputs(2989) <= layer6_outputs(3296);
    layer7_outputs(2990) <= layer6_outputs(619);
    layer7_outputs(2991) <= (layer6_outputs(1686)) and not (layer6_outputs(1974));
    layer7_outputs(2992) <= not((layer6_outputs(153)) xor (layer6_outputs(1880)));
    layer7_outputs(2993) <= layer6_outputs(1252);
    layer7_outputs(2994) <= not(layer6_outputs(836));
    layer7_outputs(2995) <= not(layer6_outputs(1434));
    layer7_outputs(2996) <= (layer6_outputs(208)) xor (layer6_outputs(4912));
    layer7_outputs(2997) <= not(layer6_outputs(3432));
    layer7_outputs(2998) <= (layer6_outputs(169)) or (layer6_outputs(2917));
    layer7_outputs(2999) <= layer6_outputs(591);
    layer7_outputs(3000) <= (layer6_outputs(396)) xor (layer6_outputs(4847));
    layer7_outputs(3001) <= layer6_outputs(3816);
    layer7_outputs(3002) <= not(layer6_outputs(4442));
    layer7_outputs(3003) <= (layer6_outputs(2709)) or (layer6_outputs(4255));
    layer7_outputs(3004) <= not((layer6_outputs(974)) and (layer6_outputs(2618)));
    layer7_outputs(3005) <= (layer6_outputs(1897)) and (layer6_outputs(4472));
    layer7_outputs(3006) <= not((layer6_outputs(3115)) or (layer6_outputs(107)));
    layer7_outputs(3007) <= layer6_outputs(654);
    layer7_outputs(3008) <= layer6_outputs(4593);
    layer7_outputs(3009) <= not(layer6_outputs(2209));
    layer7_outputs(3010) <= layer6_outputs(3011);
    layer7_outputs(3011) <= (layer6_outputs(3949)) xor (layer6_outputs(1655));
    layer7_outputs(3012) <= not((layer6_outputs(3165)) xor (layer6_outputs(2481)));
    layer7_outputs(3013) <= layer6_outputs(4186);
    layer7_outputs(3014) <= (layer6_outputs(1003)) or (layer6_outputs(3214));
    layer7_outputs(3015) <= not(layer6_outputs(4705));
    layer7_outputs(3016) <= not(layer6_outputs(86)) or (layer6_outputs(3588));
    layer7_outputs(3017) <= layer6_outputs(33);
    layer7_outputs(3018) <= not(layer6_outputs(3379));
    layer7_outputs(3019) <= (layer6_outputs(1057)) or (layer6_outputs(2002));
    layer7_outputs(3020) <= not(layer6_outputs(1789)) or (layer6_outputs(2596));
    layer7_outputs(3021) <= (layer6_outputs(4050)) and not (layer6_outputs(4363));
    layer7_outputs(3022) <= not(layer6_outputs(5097)) or (layer6_outputs(2268));
    layer7_outputs(3023) <= not((layer6_outputs(224)) and (layer6_outputs(2617)));
    layer7_outputs(3024) <= layer6_outputs(439);
    layer7_outputs(3025) <= not((layer6_outputs(2682)) or (layer6_outputs(4243)));
    layer7_outputs(3026) <= (layer6_outputs(4974)) and not (layer6_outputs(4128));
    layer7_outputs(3027) <= not((layer6_outputs(4192)) xor (layer6_outputs(2895)));
    layer7_outputs(3028) <= (layer6_outputs(617)) and (layer6_outputs(282));
    layer7_outputs(3029) <= not(layer6_outputs(4790));
    layer7_outputs(3030) <= not(layer6_outputs(3590));
    layer7_outputs(3031) <= not((layer6_outputs(4961)) or (layer6_outputs(2699)));
    layer7_outputs(3032) <= not(layer6_outputs(1786));
    layer7_outputs(3033) <= (layer6_outputs(3180)) or (layer6_outputs(3852));
    layer7_outputs(3034) <= not((layer6_outputs(2165)) or (layer6_outputs(1374)));
    layer7_outputs(3035) <= not(layer6_outputs(2219));
    layer7_outputs(3036) <= layer6_outputs(2025);
    layer7_outputs(3037) <= not(layer6_outputs(4934));
    layer7_outputs(3038) <= (layer6_outputs(3293)) xor (layer6_outputs(3519));
    layer7_outputs(3039) <= (layer6_outputs(2262)) or (layer6_outputs(3656));
    layer7_outputs(3040) <= (layer6_outputs(4652)) or (layer6_outputs(3084));
    layer7_outputs(3041) <= not(layer6_outputs(3573));
    layer7_outputs(3042) <= not(layer6_outputs(1012)) or (layer6_outputs(1541));
    layer7_outputs(3043) <= (layer6_outputs(3768)) and not (layer6_outputs(3228));
    layer7_outputs(3044) <= layer6_outputs(758);
    layer7_outputs(3045) <= not(layer6_outputs(2919));
    layer7_outputs(3046) <= not(layer6_outputs(2166));
    layer7_outputs(3047) <= not((layer6_outputs(4975)) or (layer6_outputs(460)));
    layer7_outputs(3048) <= (layer6_outputs(1925)) and (layer6_outputs(1446));
    layer7_outputs(3049) <= not(layer6_outputs(1470));
    layer7_outputs(3050) <= not(layer6_outputs(133));
    layer7_outputs(3051) <= not(layer6_outputs(2907));
    layer7_outputs(3052) <= not(layer6_outputs(1259));
    layer7_outputs(3053) <= not(layer6_outputs(3127));
    layer7_outputs(3054) <= not((layer6_outputs(531)) xor (layer6_outputs(2240)));
    layer7_outputs(3055) <= (layer6_outputs(3740)) and not (layer6_outputs(727));
    layer7_outputs(3056) <= layer6_outputs(2808);
    layer7_outputs(3057) <= layer6_outputs(3096);
    layer7_outputs(3058) <= not(layer6_outputs(1891));
    layer7_outputs(3059) <= not(layer6_outputs(3363)) or (layer6_outputs(4017));
    layer7_outputs(3060) <= (layer6_outputs(4667)) and (layer6_outputs(786));
    layer7_outputs(3061) <= not(layer6_outputs(1681));
    layer7_outputs(3062) <= not((layer6_outputs(3046)) and (layer6_outputs(2443)));
    layer7_outputs(3063) <= (layer6_outputs(3428)) or (layer6_outputs(2160));
    layer7_outputs(3064) <= not((layer6_outputs(4403)) and (layer6_outputs(1337)));
    layer7_outputs(3065) <= not((layer6_outputs(2258)) and (layer6_outputs(2392)));
    layer7_outputs(3066) <= (layer6_outputs(3831)) and (layer6_outputs(4233));
    layer7_outputs(3067) <= '1';
    layer7_outputs(3068) <= (layer6_outputs(3331)) xor (layer6_outputs(1108));
    layer7_outputs(3069) <= layer6_outputs(4141);
    layer7_outputs(3070) <= layer6_outputs(3583);
    layer7_outputs(3071) <= (layer6_outputs(1104)) and not (layer6_outputs(954));
    layer7_outputs(3072) <= layer6_outputs(1475);
    layer7_outputs(3073) <= not((layer6_outputs(1546)) and (layer6_outputs(278)));
    layer7_outputs(3074) <= not(layer6_outputs(2059));
    layer7_outputs(3075) <= not(layer6_outputs(3061));
    layer7_outputs(3076) <= layer6_outputs(2051);
    layer7_outputs(3077) <= not(layer6_outputs(4713));
    layer7_outputs(3078) <= (layer6_outputs(4095)) or (layer6_outputs(4452));
    layer7_outputs(3079) <= layer6_outputs(1679);
    layer7_outputs(3080) <= (layer6_outputs(3169)) xor (layer6_outputs(3560));
    layer7_outputs(3081) <= (layer6_outputs(4785)) xor (layer6_outputs(2932));
    layer7_outputs(3082) <= (layer6_outputs(4082)) and not (layer6_outputs(3387));
    layer7_outputs(3083) <= (layer6_outputs(4010)) and not (layer6_outputs(3138));
    layer7_outputs(3084) <= (layer6_outputs(674)) and (layer6_outputs(2320));
    layer7_outputs(3085) <= (layer6_outputs(3950)) and (layer6_outputs(3469));
    layer7_outputs(3086) <= not(layer6_outputs(1899));
    layer7_outputs(3087) <= layer6_outputs(2781);
    layer7_outputs(3088) <= layer6_outputs(34);
    layer7_outputs(3089) <= not((layer6_outputs(3343)) or (layer6_outputs(4018)));
    layer7_outputs(3090) <= not((layer6_outputs(3181)) or (layer6_outputs(2824)));
    layer7_outputs(3091) <= not((layer6_outputs(2972)) xor (layer6_outputs(1552)));
    layer7_outputs(3092) <= layer6_outputs(3174);
    layer7_outputs(3093) <= not(layer6_outputs(4209));
    layer7_outputs(3094) <= not(layer6_outputs(2834));
    layer7_outputs(3095) <= not(layer6_outputs(1989));
    layer7_outputs(3096) <= not((layer6_outputs(382)) or (layer6_outputs(2967)));
    layer7_outputs(3097) <= not((layer6_outputs(1043)) and (layer6_outputs(724)));
    layer7_outputs(3098) <= not(layer6_outputs(1381));
    layer7_outputs(3099) <= (layer6_outputs(1026)) or (layer6_outputs(914));
    layer7_outputs(3100) <= not((layer6_outputs(4682)) xor (layer6_outputs(2740)));
    layer7_outputs(3101) <= not(layer6_outputs(4236));
    layer7_outputs(3102) <= not(layer6_outputs(3122)) or (layer6_outputs(1376));
    layer7_outputs(3103) <= layer6_outputs(2153);
    layer7_outputs(3104) <= not((layer6_outputs(3450)) or (layer6_outputs(3023)));
    layer7_outputs(3105) <= '0';
    layer7_outputs(3106) <= not(layer6_outputs(2510));
    layer7_outputs(3107) <= (layer6_outputs(3593)) and not (layer6_outputs(2362));
    layer7_outputs(3108) <= (layer6_outputs(2898)) xor (layer6_outputs(3348));
    layer7_outputs(3109) <= not(layer6_outputs(2530));
    layer7_outputs(3110) <= (layer6_outputs(1293)) or (layer6_outputs(843));
    layer7_outputs(3111) <= not(layer6_outputs(546));
    layer7_outputs(3112) <= (layer6_outputs(3535)) xor (layer6_outputs(1732));
    layer7_outputs(3113) <= (layer6_outputs(2196)) xor (layer6_outputs(1854));
    layer7_outputs(3114) <= not(layer6_outputs(1436)) or (layer6_outputs(417));
    layer7_outputs(3115) <= (layer6_outputs(1320)) or (layer6_outputs(2867));
    layer7_outputs(3116) <= layer6_outputs(1553);
    layer7_outputs(3117) <= (layer6_outputs(4791)) or (layer6_outputs(3500));
    layer7_outputs(3118) <= not(layer6_outputs(1847)) or (layer6_outputs(2686));
    layer7_outputs(3119) <= layer6_outputs(2085);
    layer7_outputs(3120) <= (layer6_outputs(1556)) xor (layer6_outputs(4014));
    layer7_outputs(3121) <= (layer6_outputs(4144)) xor (layer6_outputs(4713));
    layer7_outputs(3122) <= (layer6_outputs(4227)) or (layer6_outputs(2617));
    layer7_outputs(3123) <= layer6_outputs(753);
    layer7_outputs(3124) <= not(layer6_outputs(4576));
    layer7_outputs(3125) <= layer6_outputs(85);
    layer7_outputs(3126) <= layer6_outputs(1559);
    layer7_outputs(3127) <= not(layer6_outputs(4044));
    layer7_outputs(3128) <= layer6_outputs(3522);
    layer7_outputs(3129) <= (layer6_outputs(3503)) xor (layer6_outputs(5005));
    layer7_outputs(3130) <= (layer6_outputs(1574)) or (layer6_outputs(170));
    layer7_outputs(3131) <= not((layer6_outputs(675)) and (layer6_outputs(73)));
    layer7_outputs(3132) <= (layer6_outputs(4974)) and (layer6_outputs(2840));
    layer7_outputs(3133) <= not(layer6_outputs(250));
    layer7_outputs(3134) <= layer6_outputs(1722);
    layer7_outputs(3135) <= not(layer6_outputs(955));
    layer7_outputs(3136) <= not(layer6_outputs(2862));
    layer7_outputs(3137) <= not(layer6_outputs(843));
    layer7_outputs(3138) <= not(layer6_outputs(22)) or (layer6_outputs(3525));
    layer7_outputs(3139) <= layer6_outputs(500);
    layer7_outputs(3140) <= not(layer6_outputs(4759));
    layer7_outputs(3141) <= not(layer6_outputs(3943)) or (layer6_outputs(285));
    layer7_outputs(3142) <= (layer6_outputs(4013)) xor (layer6_outputs(4875));
    layer7_outputs(3143) <= not(layer6_outputs(496));
    layer7_outputs(3144) <= (layer6_outputs(469)) or (layer6_outputs(201));
    layer7_outputs(3145) <= not(layer6_outputs(2859));
    layer7_outputs(3146) <= (layer6_outputs(827)) xor (layer6_outputs(2230));
    layer7_outputs(3147) <= not(layer6_outputs(3258)) or (layer6_outputs(514));
    layer7_outputs(3148) <= not(layer6_outputs(2692));
    layer7_outputs(3149) <= not(layer6_outputs(461));
    layer7_outputs(3150) <= not(layer6_outputs(2723));
    layer7_outputs(3151) <= not(layer6_outputs(2314)) or (layer6_outputs(3562));
    layer7_outputs(3152) <= not(layer6_outputs(3944)) or (layer6_outputs(1677));
    layer7_outputs(3153) <= not((layer6_outputs(573)) or (layer6_outputs(1355)));
    layer7_outputs(3154) <= not(layer6_outputs(1213));
    layer7_outputs(3155) <= layer6_outputs(1106);
    layer7_outputs(3156) <= not((layer6_outputs(3424)) or (layer6_outputs(255)));
    layer7_outputs(3157) <= not(layer6_outputs(3238));
    layer7_outputs(3158) <= (layer6_outputs(750)) and not (layer6_outputs(3507));
    layer7_outputs(3159) <= not(layer6_outputs(2359));
    layer7_outputs(3160) <= not(layer6_outputs(1275));
    layer7_outputs(3161) <= (layer6_outputs(4442)) and not (layer6_outputs(1949));
    layer7_outputs(3162) <= (layer6_outputs(1008)) xor (layer6_outputs(2603));
    layer7_outputs(3163) <= not((layer6_outputs(4189)) and (layer6_outputs(4734)));
    layer7_outputs(3164) <= not(layer6_outputs(483));
    layer7_outputs(3165) <= not(layer6_outputs(1212)) or (layer6_outputs(1212));
    layer7_outputs(3166) <= layer6_outputs(815);
    layer7_outputs(3167) <= (layer6_outputs(5038)) and not (layer6_outputs(4775));
    layer7_outputs(3168) <= not(layer6_outputs(4566));
    layer7_outputs(3169) <= not(layer6_outputs(5113)) or (layer6_outputs(1947));
    layer7_outputs(3170) <= not(layer6_outputs(4274)) or (layer6_outputs(4848));
    layer7_outputs(3171) <= layer6_outputs(696);
    layer7_outputs(3172) <= (layer6_outputs(3696)) and not (layer6_outputs(3924));
    layer7_outputs(3173) <= not(layer6_outputs(4860));
    layer7_outputs(3174) <= not(layer6_outputs(4366)) or (layer6_outputs(1784));
    layer7_outputs(3175) <= not((layer6_outputs(4378)) xor (layer6_outputs(3172)));
    layer7_outputs(3176) <= not(layer6_outputs(4081));
    layer7_outputs(3177) <= not((layer6_outputs(2201)) xor (layer6_outputs(392)));
    layer7_outputs(3178) <= layer6_outputs(2186);
    layer7_outputs(3179) <= not(layer6_outputs(650));
    layer7_outputs(3180) <= not(layer6_outputs(1989)) or (layer6_outputs(1272));
    layer7_outputs(3181) <= not((layer6_outputs(2955)) or (layer6_outputs(2291)));
    layer7_outputs(3182) <= layer6_outputs(4998);
    layer7_outputs(3183) <= (layer6_outputs(753)) or (layer6_outputs(1661));
    layer7_outputs(3184) <= not((layer6_outputs(1449)) or (layer6_outputs(4371)));
    layer7_outputs(3185) <= not(layer6_outputs(929));
    layer7_outputs(3186) <= (layer6_outputs(2442)) xor (layer6_outputs(2188));
    layer7_outputs(3187) <= (layer6_outputs(2018)) and not (layer6_outputs(484));
    layer7_outputs(3188) <= not(layer6_outputs(4952));
    layer7_outputs(3189) <= layer6_outputs(4295);
    layer7_outputs(3190) <= layer6_outputs(2077);
    layer7_outputs(3191) <= (layer6_outputs(4996)) and not (layer6_outputs(10));
    layer7_outputs(3192) <= not(layer6_outputs(4810)) or (layer6_outputs(583));
    layer7_outputs(3193) <= (layer6_outputs(1901)) xor (layer6_outputs(175));
    layer7_outputs(3194) <= layer6_outputs(1897);
    layer7_outputs(3195) <= not(layer6_outputs(1123));
    layer7_outputs(3196) <= not(layer6_outputs(4958));
    layer7_outputs(3197) <= not(layer6_outputs(4495)) or (layer6_outputs(3204));
    layer7_outputs(3198) <= (layer6_outputs(3477)) and not (layer6_outputs(3189));
    layer7_outputs(3199) <= not(layer6_outputs(2238));
    layer7_outputs(3200) <= not(layer6_outputs(4816));
    layer7_outputs(3201) <= layer6_outputs(4811);
    layer7_outputs(3202) <= not(layer6_outputs(4785));
    layer7_outputs(3203) <= not((layer6_outputs(3741)) xor (layer6_outputs(4060)));
    layer7_outputs(3204) <= not((layer6_outputs(4545)) xor (layer6_outputs(2580)));
    layer7_outputs(3205) <= not((layer6_outputs(693)) or (layer6_outputs(3694)));
    layer7_outputs(3206) <= (layer6_outputs(3826)) and not (layer6_outputs(113));
    layer7_outputs(3207) <= (layer6_outputs(2482)) and not (layer6_outputs(4001));
    layer7_outputs(3208) <= not(layer6_outputs(4691));
    layer7_outputs(3209) <= not(layer6_outputs(792));
    layer7_outputs(3210) <= not(layer6_outputs(1138)) or (layer6_outputs(1169));
    layer7_outputs(3211) <= not((layer6_outputs(1650)) and (layer6_outputs(562)));
    layer7_outputs(3212) <= not(layer6_outputs(148));
    layer7_outputs(3213) <= not((layer6_outputs(4042)) and (layer6_outputs(103)));
    layer7_outputs(3214) <= (layer6_outputs(4229)) xor (layer6_outputs(2385));
    layer7_outputs(3215) <= layer6_outputs(3961);
    layer7_outputs(3216) <= not(layer6_outputs(2871));
    layer7_outputs(3217) <= not(layer6_outputs(1835));
    layer7_outputs(3218) <= layer6_outputs(2076);
    layer7_outputs(3219) <= not(layer6_outputs(1562));
    layer7_outputs(3220) <= not(layer6_outputs(1842));
    layer7_outputs(3221) <= layer6_outputs(1719);
    layer7_outputs(3222) <= not((layer6_outputs(4674)) xor (layer6_outputs(1648)));
    layer7_outputs(3223) <= layer6_outputs(1534);
    layer7_outputs(3224) <= layer6_outputs(2884);
    layer7_outputs(3225) <= not(layer6_outputs(3021));
    layer7_outputs(3226) <= layer6_outputs(4360);
    layer7_outputs(3227) <= not((layer6_outputs(2490)) or (layer6_outputs(2435)));
    layer7_outputs(3228) <= (layer6_outputs(3785)) xor (layer6_outputs(102));
    layer7_outputs(3229) <= layer6_outputs(3531);
    layer7_outputs(3230) <= (layer6_outputs(2770)) and not (layer6_outputs(945));
    layer7_outputs(3231) <= not(layer6_outputs(3864));
    layer7_outputs(3232) <= (layer6_outputs(3876)) xor (layer6_outputs(4469));
    layer7_outputs(3233) <= not(layer6_outputs(743));
    layer7_outputs(3234) <= '0';
    layer7_outputs(3235) <= layer6_outputs(4318);
    layer7_outputs(3236) <= (layer6_outputs(4076)) xor (layer6_outputs(2230));
    layer7_outputs(3237) <= layer6_outputs(4775);
    layer7_outputs(3238) <= not((layer6_outputs(4313)) and (layer6_outputs(4696)));
    layer7_outputs(3239) <= layer6_outputs(4721);
    layer7_outputs(3240) <= not((layer6_outputs(2640)) xor (layer6_outputs(267)));
    layer7_outputs(3241) <= not(layer6_outputs(896));
    layer7_outputs(3242) <= not(layer6_outputs(1020));
    layer7_outputs(3243) <= not(layer6_outputs(4705));
    layer7_outputs(3244) <= (layer6_outputs(3017)) and (layer6_outputs(4308));
    layer7_outputs(3245) <= (layer6_outputs(3024)) xor (layer6_outputs(3255));
    layer7_outputs(3246) <= not(layer6_outputs(2621));
    layer7_outputs(3247) <= layer6_outputs(49);
    layer7_outputs(3248) <= not(layer6_outputs(2488));
    layer7_outputs(3249) <= layer6_outputs(3723);
    layer7_outputs(3250) <= (layer6_outputs(2756)) xor (layer6_outputs(1570));
    layer7_outputs(3251) <= not(layer6_outputs(355)) or (layer6_outputs(306));
    layer7_outputs(3252) <= not(layer6_outputs(917));
    layer7_outputs(3253) <= (layer6_outputs(3296)) and (layer6_outputs(4553));
    layer7_outputs(3254) <= not((layer6_outputs(4551)) or (layer6_outputs(809)));
    layer7_outputs(3255) <= layer6_outputs(2821);
    layer7_outputs(3256) <= not((layer6_outputs(2533)) xor (layer6_outputs(4916)));
    layer7_outputs(3257) <= (layer6_outputs(1040)) xor (layer6_outputs(222));
    layer7_outputs(3258) <= layer6_outputs(2474);
    layer7_outputs(3259) <= (layer6_outputs(2217)) and not (layer6_outputs(1771));
    layer7_outputs(3260) <= layer6_outputs(5110);
    layer7_outputs(3261) <= not(layer6_outputs(4353));
    layer7_outputs(3262) <= layer6_outputs(744);
    layer7_outputs(3263) <= (layer6_outputs(2328)) xor (layer6_outputs(932));
    layer7_outputs(3264) <= not((layer6_outputs(4561)) and (layer6_outputs(4897)));
    layer7_outputs(3265) <= (layer6_outputs(4492)) and not (layer6_outputs(4644));
    layer7_outputs(3266) <= not(layer6_outputs(2942));
    layer7_outputs(3267) <= layer6_outputs(432);
    layer7_outputs(3268) <= not(layer6_outputs(2620));
    layer7_outputs(3269) <= (layer6_outputs(4814)) and (layer6_outputs(2654));
    layer7_outputs(3270) <= (layer6_outputs(2484)) and not (layer6_outputs(397));
    layer7_outputs(3271) <= (layer6_outputs(2373)) and not (layer6_outputs(2422));
    layer7_outputs(3272) <= not(layer6_outputs(4418));
    layer7_outputs(3273) <= layer6_outputs(2077);
    layer7_outputs(3274) <= (layer6_outputs(4088)) xor (layer6_outputs(3795));
    layer7_outputs(3275) <= not((layer6_outputs(1531)) or (layer6_outputs(2726)));
    layer7_outputs(3276) <= layer6_outputs(2082);
    layer7_outputs(3277) <= not(layer6_outputs(1987));
    layer7_outputs(3278) <= layer6_outputs(79);
    layer7_outputs(3279) <= not(layer6_outputs(4217));
    layer7_outputs(3280) <= not(layer6_outputs(1118)) or (layer6_outputs(4396));
    layer7_outputs(3281) <= '0';
    layer7_outputs(3282) <= (layer6_outputs(1629)) or (layer6_outputs(300));
    layer7_outputs(3283) <= not(layer6_outputs(1234));
    layer7_outputs(3284) <= not(layer6_outputs(2792)) or (layer6_outputs(2569));
    layer7_outputs(3285) <= not(layer6_outputs(2718)) or (layer6_outputs(240));
    layer7_outputs(3286) <= (layer6_outputs(121)) xor (layer6_outputs(3550));
    layer7_outputs(3287) <= layer6_outputs(1776);
    layer7_outputs(3288) <= not(layer6_outputs(931));
    layer7_outputs(3289) <= layer6_outputs(849);
    layer7_outputs(3290) <= layer6_outputs(2187);
    layer7_outputs(3291) <= (layer6_outputs(3642)) xor (layer6_outputs(68));
    layer7_outputs(3292) <= layer6_outputs(714);
    layer7_outputs(3293) <= not(layer6_outputs(1982)) or (layer6_outputs(4038));
    layer7_outputs(3294) <= layer6_outputs(5010);
    layer7_outputs(3295) <= not(layer6_outputs(3057));
    layer7_outputs(3296) <= not(layer6_outputs(4534)) or (layer6_outputs(4598));
    layer7_outputs(3297) <= not((layer6_outputs(3588)) xor (layer6_outputs(4402)));
    layer7_outputs(3298) <= layer6_outputs(3100);
    layer7_outputs(3299) <= not(layer6_outputs(4604));
    layer7_outputs(3300) <= not(layer6_outputs(3383));
    layer7_outputs(3301) <= not(layer6_outputs(3570)) or (layer6_outputs(4692));
    layer7_outputs(3302) <= (layer6_outputs(872)) or (layer6_outputs(851));
    layer7_outputs(3303) <= layer6_outputs(1390);
    layer7_outputs(3304) <= layer6_outputs(1971);
    layer7_outputs(3305) <= not(layer6_outputs(930));
    layer7_outputs(3306) <= (layer6_outputs(2633)) and not (layer6_outputs(4360));
    layer7_outputs(3307) <= layer6_outputs(2733);
    layer7_outputs(3308) <= not(layer6_outputs(219));
    layer7_outputs(3309) <= not((layer6_outputs(4047)) or (layer6_outputs(428)));
    layer7_outputs(3310) <= layer6_outputs(3376);
    layer7_outputs(3311) <= (layer6_outputs(2652)) xor (layer6_outputs(746));
    layer7_outputs(3312) <= not((layer6_outputs(3286)) xor (layer6_outputs(2678)));
    layer7_outputs(3313) <= not(layer6_outputs(1201));
    layer7_outputs(3314) <= not(layer6_outputs(601)) or (layer6_outputs(4294));
    layer7_outputs(3315) <= not(layer6_outputs(997));
    layer7_outputs(3316) <= not((layer6_outputs(4225)) xor (layer6_outputs(2216)));
    layer7_outputs(3317) <= layer6_outputs(658);
    layer7_outputs(3318) <= not(layer6_outputs(2767));
    layer7_outputs(3319) <= not(layer6_outputs(1710));
    layer7_outputs(3320) <= not(layer6_outputs(5103));
    layer7_outputs(3321) <= layer6_outputs(4210);
    layer7_outputs(3322) <= (layer6_outputs(865)) and not (layer6_outputs(4715));
    layer7_outputs(3323) <= (layer6_outputs(813)) and not (layer6_outputs(1752));
    layer7_outputs(3324) <= not(layer6_outputs(2274)) or (layer6_outputs(4358));
    layer7_outputs(3325) <= (layer6_outputs(2151)) and (layer6_outputs(5011));
    layer7_outputs(3326) <= layer6_outputs(3045);
    layer7_outputs(3327) <= (layer6_outputs(156)) xor (layer6_outputs(134));
    layer7_outputs(3328) <= layer6_outputs(2250);
    layer7_outputs(3329) <= layer6_outputs(2304);
    layer7_outputs(3330) <= not(layer6_outputs(192));
    layer7_outputs(3331) <= layer6_outputs(2975);
    layer7_outputs(3332) <= '1';
    layer7_outputs(3333) <= (layer6_outputs(3614)) xor (layer6_outputs(1585));
    layer7_outputs(3334) <= '0';
    layer7_outputs(3335) <= not((layer6_outputs(95)) xor (layer6_outputs(4037)));
    layer7_outputs(3336) <= not((layer6_outputs(2095)) xor (layer6_outputs(2304)));
    layer7_outputs(3337) <= not(layer6_outputs(3796)) or (layer6_outputs(2944));
    layer7_outputs(3338) <= not(layer6_outputs(1488)) or (layer6_outputs(761));
    layer7_outputs(3339) <= layer6_outputs(1826);
    layer7_outputs(3340) <= layer6_outputs(4925);
    layer7_outputs(3341) <= not((layer6_outputs(4040)) or (layer6_outputs(3617)));
    layer7_outputs(3342) <= not(layer6_outputs(3340));
    layer7_outputs(3343) <= (layer6_outputs(3915)) and not (layer6_outputs(4022));
    layer7_outputs(3344) <= not((layer6_outputs(2316)) xor (layer6_outputs(1422)));
    layer7_outputs(3345) <= layer6_outputs(3967);
    layer7_outputs(3346) <= not(layer6_outputs(2587)) or (layer6_outputs(1435));
    layer7_outputs(3347) <= not(layer6_outputs(2181));
    layer7_outputs(3348) <= not(layer6_outputs(135)) or (layer6_outputs(4113));
    layer7_outputs(3349) <= (layer6_outputs(1599)) or (layer6_outputs(349));
    layer7_outputs(3350) <= not(layer6_outputs(1569)) or (layer6_outputs(2911));
    layer7_outputs(3351) <= (layer6_outputs(2968)) xor (layer6_outputs(251));
    layer7_outputs(3352) <= not(layer6_outputs(3676)) or (layer6_outputs(5053));
    layer7_outputs(3353) <= not((layer6_outputs(3473)) xor (layer6_outputs(4569)));
    layer7_outputs(3354) <= not((layer6_outputs(5009)) xor (layer6_outputs(4267)));
    layer7_outputs(3355) <= not(layer6_outputs(1267));
    layer7_outputs(3356) <= not(layer6_outputs(2034));
    layer7_outputs(3357) <= not(layer6_outputs(2399));
    layer7_outputs(3358) <= layer6_outputs(1516);
    layer7_outputs(3359) <= not((layer6_outputs(618)) xor (layer6_outputs(1071)));
    layer7_outputs(3360) <= layer6_outputs(2528);
    layer7_outputs(3361) <= not((layer6_outputs(3990)) xor (layer6_outputs(4307)));
    layer7_outputs(3362) <= not(layer6_outputs(79)) or (layer6_outputs(4752));
    layer7_outputs(3363) <= layer6_outputs(4283);
    layer7_outputs(3364) <= (layer6_outputs(165)) xor (layer6_outputs(1737));
    layer7_outputs(3365) <= layer6_outputs(1306);
    layer7_outputs(3366) <= not((layer6_outputs(5005)) xor (layer6_outputs(3884)));
    layer7_outputs(3367) <= layer6_outputs(3025);
    layer7_outputs(3368) <= not(layer6_outputs(301));
    layer7_outputs(3369) <= layer6_outputs(3712);
    layer7_outputs(3370) <= layer6_outputs(1834);
    layer7_outputs(3371) <= not((layer6_outputs(1322)) xor (layer6_outputs(38)));
    layer7_outputs(3372) <= '1';
    layer7_outputs(3373) <= (layer6_outputs(3431)) and not (layer6_outputs(198));
    layer7_outputs(3374) <= layer6_outputs(3922);
    layer7_outputs(3375) <= layer6_outputs(3260);
    layer7_outputs(3376) <= not(layer6_outputs(1215));
    layer7_outputs(3377) <= not((layer6_outputs(1431)) xor (layer6_outputs(305)));
    layer7_outputs(3378) <= (layer6_outputs(2243)) and not (layer6_outputs(3568));
    layer7_outputs(3379) <= not((layer6_outputs(1257)) xor (layer6_outputs(2272)));
    layer7_outputs(3380) <= layer6_outputs(16);
    layer7_outputs(3381) <= '0';
    layer7_outputs(3382) <= not((layer6_outputs(570)) and (layer6_outputs(1504)));
    layer7_outputs(3383) <= layer6_outputs(4947);
    layer7_outputs(3384) <= (layer6_outputs(1140)) or (layer6_outputs(4204));
    layer7_outputs(3385) <= not((layer6_outputs(879)) or (layer6_outputs(1256)));
    layer7_outputs(3386) <= layer6_outputs(4069);
    layer7_outputs(3387) <= layer6_outputs(2969);
    layer7_outputs(3388) <= layer6_outputs(3029);
    layer7_outputs(3389) <= not((layer6_outputs(963)) and (layer6_outputs(4032)));
    layer7_outputs(3390) <= not(layer6_outputs(2241));
    layer7_outputs(3391) <= layer6_outputs(1491);
    layer7_outputs(3392) <= not(layer6_outputs(2648));
    layer7_outputs(3393) <= (layer6_outputs(3870)) and (layer6_outputs(4459));
    layer7_outputs(3394) <= not((layer6_outputs(1711)) and (layer6_outputs(3914)));
    layer7_outputs(3395) <= layer6_outputs(4676);
    layer7_outputs(3396) <= layer6_outputs(2217);
    layer7_outputs(3397) <= not((layer6_outputs(67)) xor (layer6_outputs(2562)));
    layer7_outputs(3398) <= not(layer6_outputs(4527));
    layer7_outputs(3399) <= not((layer6_outputs(436)) and (layer6_outputs(2146)));
    layer7_outputs(3400) <= not(layer6_outputs(2920));
    layer7_outputs(3401) <= layer6_outputs(1785);
    layer7_outputs(3402) <= (layer6_outputs(185)) and not (layer6_outputs(659));
    layer7_outputs(3403) <= not(layer6_outputs(3135));
    layer7_outputs(3404) <= not((layer6_outputs(4926)) and (layer6_outputs(3331)));
    layer7_outputs(3405) <= layer6_outputs(1921);
    layer7_outputs(3406) <= not(layer6_outputs(176)) or (layer6_outputs(4145));
    layer7_outputs(3407) <= not(layer6_outputs(51)) or (layer6_outputs(39));
    layer7_outputs(3408) <= not((layer6_outputs(3298)) xor (layer6_outputs(1344)));
    layer7_outputs(3409) <= not((layer6_outputs(1941)) or (layer6_outputs(2008)));
    layer7_outputs(3410) <= (layer6_outputs(3353)) xor (layer6_outputs(1894));
    layer7_outputs(3411) <= not(layer6_outputs(5065));
    layer7_outputs(3412) <= not(layer6_outputs(1479));
    layer7_outputs(3413) <= layer6_outputs(4987);
    layer7_outputs(3414) <= (layer6_outputs(4128)) xor (layer6_outputs(1784));
    layer7_outputs(3415) <= layer6_outputs(748);
    layer7_outputs(3416) <= not((layer6_outputs(2228)) xor (layer6_outputs(4126)));
    layer7_outputs(3417) <= not(layer6_outputs(1411)) or (layer6_outputs(1495));
    layer7_outputs(3418) <= layer6_outputs(30);
    layer7_outputs(3419) <= not(layer6_outputs(2684));
    layer7_outputs(3420) <= (layer6_outputs(1079)) and not (layer6_outputs(3099));
    layer7_outputs(3421) <= not((layer6_outputs(4532)) or (layer6_outputs(967)));
    layer7_outputs(3422) <= (layer6_outputs(2759)) xor (layer6_outputs(460));
    layer7_outputs(3423) <= not((layer6_outputs(4561)) or (layer6_outputs(4045)));
    layer7_outputs(3424) <= layer6_outputs(4088);
    layer7_outputs(3425) <= not((layer6_outputs(2001)) xor (layer6_outputs(1288)));
    layer7_outputs(3426) <= layer6_outputs(2472);
    layer7_outputs(3427) <= not(layer6_outputs(628));
    layer7_outputs(3428) <= (layer6_outputs(5081)) and (layer6_outputs(3627));
    layer7_outputs(3429) <= layer6_outputs(1736);
    layer7_outputs(3430) <= layer6_outputs(3694);
    layer7_outputs(3431) <= (layer6_outputs(5109)) and not (layer6_outputs(906));
    layer7_outputs(3432) <= layer6_outputs(4633);
    layer7_outputs(3433) <= layer6_outputs(180);
    layer7_outputs(3434) <= layer6_outputs(354);
    layer7_outputs(3435) <= not(layer6_outputs(1429));
    layer7_outputs(3436) <= not((layer6_outputs(4715)) xor (layer6_outputs(3289)));
    layer7_outputs(3437) <= not(layer6_outputs(3718)) or (layer6_outputs(3623));
    layer7_outputs(3438) <= not(layer6_outputs(972));
    layer7_outputs(3439) <= not((layer6_outputs(4820)) xor (layer6_outputs(3221)));
    layer7_outputs(3440) <= (layer6_outputs(327)) and not (layer6_outputs(2499));
    layer7_outputs(3441) <= layer6_outputs(1565);
    layer7_outputs(3442) <= layer6_outputs(117);
    layer7_outputs(3443) <= layer6_outputs(378);
    layer7_outputs(3444) <= (layer6_outputs(3692)) and not (layer6_outputs(3514));
    layer7_outputs(3445) <= (layer6_outputs(4876)) and not (layer6_outputs(3587));
    layer7_outputs(3446) <= layer6_outputs(4196);
    layer7_outputs(3447) <= layer6_outputs(811);
    layer7_outputs(3448) <= not(layer6_outputs(1801));
    layer7_outputs(3449) <= not(layer6_outputs(2011));
    layer7_outputs(3450) <= not(layer6_outputs(3945));
    layer7_outputs(3451) <= layer6_outputs(818);
    layer7_outputs(3452) <= layer6_outputs(31);
    layer7_outputs(3453) <= not(layer6_outputs(1315)) or (layer6_outputs(4774));
    layer7_outputs(3454) <= not((layer6_outputs(1162)) xor (layer6_outputs(412)));
    layer7_outputs(3455) <= not(layer6_outputs(1814));
    layer7_outputs(3456) <= not((layer6_outputs(3687)) xor (layer6_outputs(3281)));
    layer7_outputs(3457) <= (layer6_outputs(187)) and (layer6_outputs(1653));
    layer7_outputs(3458) <= not(layer6_outputs(3402)) or (layer6_outputs(414));
    layer7_outputs(3459) <= not(layer6_outputs(3541));
    layer7_outputs(3460) <= not(layer6_outputs(4748));
    layer7_outputs(3461) <= not(layer6_outputs(886));
    layer7_outputs(3462) <= layer6_outputs(1132);
    layer7_outputs(3463) <= layer6_outputs(1262);
    layer7_outputs(3464) <= '1';
    layer7_outputs(3465) <= not(layer6_outputs(3090));
    layer7_outputs(3466) <= layer6_outputs(1219);
    layer7_outputs(3467) <= not((layer6_outputs(3140)) xor (layer6_outputs(3547)));
    layer7_outputs(3468) <= (layer6_outputs(2229)) xor (layer6_outputs(2967));
    layer7_outputs(3469) <= layer6_outputs(1333);
    layer7_outputs(3470) <= not(layer6_outputs(3686));
    layer7_outputs(3471) <= layer6_outputs(4181);
    layer7_outputs(3472) <= not(layer6_outputs(2716)) or (layer6_outputs(1451));
    layer7_outputs(3473) <= not(layer6_outputs(211)) or (layer6_outputs(2197));
    layer7_outputs(3474) <= not(layer6_outputs(2681));
    layer7_outputs(3475) <= layer6_outputs(4359);
    layer7_outputs(3476) <= not((layer6_outputs(2805)) and (layer6_outputs(4997)));
    layer7_outputs(3477) <= not((layer6_outputs(5015)) or (layer6_outputs(2529)));
    layer7_outputs(3478) <= not(layer6_outputs(1110)) or (layer6_outputs(418));
    layer7_outputs(3479) <= not((layer6_outputs(4568)) xor (layer6_outputs(3418)));
    layer7_outputs(3480) <= (layer6_outputs(110)) xor (layer6_outputs(4656));
    layer7_outputs(3481) <= not((layer6_outputs(1010)) xor (layer6_outputs(3043)));
    layer7_outputs(3482) <= (layer6_outputs(1727)) xor (layer6_outputs(4863));
    layer7_outputs(3483) <= (layer6_outputs(2237)) and not (layer6_outputs(4889));
    layer7_outputs(3484) <= (layer6_outputs(1859)) or (layer6_outputs(3553));
    layer7_outputs(3485) <= layer6_outputs(913);
    layer7_outputs(3486) <= (layer6_outputs(2199)) xor (layer6_outputs(3145));
    layer7_outputs(3487) <= not(layer6_outputs(3469)) or (layer6_outputs(542));
    layer7_outputs(3488) <= not(layer6_outputs(1299));
    layer7_outputs(3489) <= not(layer6_outputs(1919));
    layer7_outputs(3490) <= (layer6_outputs(1928)) or (layer6_outputs(3335));
    layer7_outputs(3491) <= (layer6_outputs(1103)) xor (layer6_outputs(3434));
    layer7_outputs(3492) <= not((layer6_outputs(2183)) xor (layer6_outputs(1742)));
    layer7_outputs(3493) <= not(layer6_outputs(3976)) or (layer6_outputs(4670));
    layer7_outputs(3494) <= layer6_outputs(1025);
    layer7_outputs(3495) <= not(layer6_outputs(4263)) or (layer6_outputs(623));
    layer7_outputs(3496) <= not(layer6_outputs(3799));
    layer7_outputs(3497) <= not(layer6_outputs(4965));
    layer7_outputs(3498) <= not(layer6_outputs(1000));
    layer7_outputs(3499) <= (layer6_outputs(2894)) and (layer6_outputs(2629));
    layer7_outputs(3500) <= layer6_outputs(3116);
    layer7_outputs(3501) <= layer6_outputs(3378);
    layer7_outputs(3502) <= not(layer6_outputs(2271)) or (layer6_outputs(141));
    layer7_outputs(3503) <= not(layer6_outputs(3247));
    layer7_outputs(3504) <= not(layer6_outputs(1968));
    layer7_outputs(3505) <= layer6_outputs(3708);
    layer7_outputs(3506) <= not(layer6_outputs(1588)) or (layer6_outputs(1943));
    layer7_outputs(3507) <= not((layer6_outputs(3281)) or (layer6_outputs(3980)));
    layer7_outputs(3508) <= layer6_outputs(2896);
    layer7_outputs(3509) <= not(layer6_outputs(2118)) or (layer6_outputs(1130));
    layer7_outputs(3510) <= not(layer6_outputs(4906));
    layer7_outputs(3511) <= layer6_outputs(2657);
    layer7_outputs(3512) <= not((layer6_outputs(816)) xor (layer6_outputs(1700)));
    layer7_outputs(3513) <= (layer6_outputs(4843)) and not (layer6_outputs(689));
    layer7_outputs(3514) <= (layer6_outputs(2665)) xor (layer6_outputs(4422));
    layer7_outputs(3515) <= not(layer6_outputs(3186));
    layer7_outputs(3516) <= (layer6_outputs(4478)) or (layer6_outputs(3628));
    layer7_outputs(3517) <= layer6_outputs(1721);
    layer7_outputs(3518) <= (layer6_outputs(4948)) and not (layer6_outputs(2104));
    layer7_outputs(3519) <= not((layer6_outputs(640)) and (layer6_outputs(3408)));
    layer7_outputs(3520) <= not((layer6_outputs(837)) xor (layer6_outputs(4007)));
    layer7_outputs(3521) <= not(layer6_outputs(1166));
    layer7_outputs(3522) <= (layer6_outputs(1766)) or (layer6_outputs(4365));
    layer7_outputs(3523) <= (layer6_outputs(907)) and not (layer6_outputs(2050));
    layer7_outputs(3524) <= not(layer6_outputs(3777));
    layer7_outputs(3525) <= (layer6_outputs(3034)) and not (layer6_outputs(1239));
    layer7_outputs(3526) <= not((layer6_outputs(3811)) xor (layer6_outputs(4208)));
    layer7_outputs(3527) <= (layer6_outputs(4117)) and (layer6_outputs(2540));
    layer7_outputs(3528) <= (layer6_outputs(4595)) and (layer6_outputs(425));
    layer7_outputs(3529) <= not(layer6_outputs(605)) or (layer6_outputs(564));
    layer7_outputs(3530) <= not(layer6_outputs(2013));
    layer7_outputs(3531) <= layer6_outputs(3072);
    layer7_outputs(3532) <= not(layer6_outputs(3750));
    layer7_outputs(3533) <= not((layer6_outputs(2676)) and (layer6_outputs(4746)));
    layer7_outputs(3534) <= not(layer6_outputs(1368)) or (layer6_outputs(3375));
    layer7_outputs(3535) <= (layer6_outputs(4452)) xor (layer6_outputs(4304));
    layer7_outputs(3536) <= layer6_outputs(505);
    layer7_outputs(3537) <= layer6_outputs(3796);
    layer7_outputs(3538) <= (layer6_outputs(1608)) xor (layer6_outputs(1904));
    layer7_outputs(3539) <= not((layer6_outputs(773)) and (layer6_outputs(3406)));
    layer7_outputs(3540) <= not(layer6_outputs(581));
    layer7_outputs(3541) <= not((layer6_outputs(3845)) xor (layer6_outputs(937)));
    layer7_outputs(3542) <= not(layer6_outputs(3847));
    layer7_outputs(3543) <= not(layer6_outputs(3397));
    layer7_outputs(3544) <= layer6_outputs(2312);
    layer7_outputs(3545) <= (layer6_outputs(3653)) xor (layer6_outputs(247));
    layer7_outputs(3546) <= layer6_outputs(1448);
    layer7_outputs(3547) <= (layer6_outputs(4508)) and not (layer6_outputs(4544));
    layer7_outputs(3548) <= '0';
    layer7_outputs(3549) <= not((layer6_outputs(5039)) and (layer6_outputs(3276)));
    layer7_outputs(3550) <= (layer6_outputs(1266)) or (layer6_outputs(4086));
    layer7_outputs(3551) <= layer6_outputs(1470);
    layer7_outputs(3552) <= (layer6_outputs(28)) and (layer6_outputs(4681));
    layer7_outputs(3553) <= not(layer6_outputs(2035));
    layer7_outputs(3554) <= (layer6_outputs(977)) and not (layer6_outputs(4115));
    layer7_outputs(3555) <= layer6_outputs(4206);
    layer7_outputs(3556) <= not(layer6_outputs(99));
    layer7_outputs(3557) <= not(layer6_outputs(1912));
    layer7_outputs(3558) <= not(layer6_outputs(3200));
    layer7_outputs(3559) <= layer6_outputs(4905);
    layer7_outputs(3560) <= layer6_outputs(3726);
    layer7_outputs(3561) <= not(layer6_outputs(5008));
    layer7_outputs(3562) <= (layer6_outputs(1934)) and not (layer6_outputs(2353));
    layer7_outputs(3563) <= (layer6_outputs(595)) and not (layer6_outputs(834));
    layer7_outputs(3564) <= not(layer6_outputs(4476));
    layer7_outputs(3565) <= not(layer6_outputs(637));
    layer7_outputs(3566) <= (layer6_outputs(4665)) xor (layer6_outputs(3516));
    layer7_outputs(3567) <= not(layer6_outputs(1986)) or (layer6_outputs(702));
    layer7_outputs(3568) <= '1';
    layer7_outputs(3569) <= not(layer6_outputs(828));
    layer7_outputs(3570) <= layer6_outputs(883);
    layer7_outputs(3571) <= (layer6_outputs(2098)) xor (layer6_outputs(1205));
    layer7_outputs(3572) <= layer6_outputs(2362);
    layer7_outputs(3573) <= not(layer6_outputs(1171));
    layer7_outputs(3574) <= not(layer6_outputs(4635));
    layer7_outputs(3575) <= layer6_outputs(645);
    layer7_outputs(3576) <= not(layer6_outputs(1785));
    layer7_outputs(3577) <= not(layer6_outputs(4808));
    layer7_outputs(3578) <= not(layer6_outputs(1188));
    layer7_outputs(3579) <= (layer6_outputs(3649)) or (layer6_outputs(1690));
    layer7_outputs(3580) <= (layer6_outputs(1713)) xor (layer6_outputs(709));
    layer7_outputs(3581) <= not((layer6_outputs(3620)) xor (layer6_outputs(4854)));
    layer7_outputs(3582) <= not((layer6_outputs(4692)) or (layer6_outputs(2554)));
    layer7_outputs(3583) <= not((layer6_outputs(3795)) xor (layer6_outputs(2725)));
    layer7_outputs(3584) <= layer6_outputs(3356);
    layer7_outputs(3585) <= not(layer6_outputs(1193));
    layer7_outputs(3586) <= (layer6_outputs(132)) and not (layer6_outputs(1937));
    layer7_outputs(3587) <= layer6_outputs(330);
    layer7_outputs(3588) <= layer6_outputs(1277);
    layer7_outputs(3589) <= layer6_outputs(3731);
    layer7_outputs(3590) <= not(layer6_outputs(4409)) or (layer6_outputs(4655));
    layer7_outputs(3591) <= not(layer6_outputs(633)) or (layer6_outputs(2028));
    layer7_outputs(3592) <= (layer6_outputs(3374)) xor (layer6_outputs(3971));
    layer7_outputs(3593) <= not((layer6_outputs(4234)) or (layer6_outputs(534)));
    layer7_outputs(3594) <= not(layer6_outputs(1717));
    layer7_outputs(3595) <= layer6_outputs(3807);
    layer7_outputs(3596) <= not(layer6_outputs(3674));
    layer7_outputs(3597) <= (layer6_outputs(805)) xor (layer6_outputs(5025));
    layer7_outputs(3598) <= layer6_outputs(2544);
    layer7_outputs(3599) <= not((layer6_outputs(1912)) or (layer6_outputs(2860)));
    layer7_outputs(3600) <= (layer6_outputs(2993)) xor (layer6_outputs(121));
    layer7_outputs(3601) <= layer6_outputs(4510);
    layer7_outputs(3602) <= (layer6_outputs(1918)) and not (layer6_outputs(2749));
    layer7_outputs(3603) <= (layer6_outputs(4960)) xor (layer6_outputs(336));
    layer7_outputs(3604) <= layer6_outputs(231);
    layer7_outputs(3605) <= (layer6_outputs(2869)) and not (layer6_outputs(2319));
    layer7_outputs(3606) <= not(layer6_outputs(4611));
    layer7_outputs(3607) <= (layer6_outputs(3353)) xor (layer6_outputs(1221));
    layer7_outputs(3608) <= not((layer6_outputs(1107)) and (layer6_outputs(696)));
    layer7_outputs(3609) <= layer6_outputs(1302);
    layer7_outputs(3610) <= not((layer6_outputs(4886)) xor (layer6_outputs(5018)));
    layer7_outputs(3611) <= not(layer6_outputs(3389));
    layer7_outputs(3612) <= not((layer6_outputs(4458)) or (layer6_outputs(3364)));
    layer7_outputs(3613) <= (layer6_outputs(2350)) or (layer6_outputs(1491));
    layer7_outputs(3614) <= '0';
    layer7_outputs(3615) <= not(layer6_outputs(4429));
    layer7_outputs(3616) <= layer6_outputs(1223);
    layer7_outputs(3617) <= not(layer6_outputs(2065));
    layer7_outputs(3618) <= (layer6_outputs(2163)) and not (layer6_outputs(1626));
    layer7_outputs(3619) <= not(layer6_outputs(395));
    layer7_outputs(3620) <= not((layer6_outputs(968)) xor (layer6_outputs(3659)));
    layer7_outputs(3621) <= layer6_outputs(604);
    layer7_outputs(3622) <= not((layer6_outputs(3740)) or (layer6_outputs(2316)));
    layer7_outputs(3623) <= (layer6_outputs(1509)) and (layer6_outputs(865));
    layer7_outputs(3624) <= (layer6_outputs(4362)) xor (layer6_outputs(4367));
    layer7_outputs(3625) <= not(layer6_outputs(4179));
    layer7_outputs(3626) <= layer6_outputs(3008);
    layer7_outputs(3627) <= layer6_outputs(3356);
    layer7_outputs(3628) <= not(layer6_outputs(1952)) or (layer6_outputs(642));
    layer7_outputs(3629) <= not(layer6_outputs(4215));
    layer7_outputs(3630) <= layer6_outputs(3769);
    layer7_outputs(3631) <= not(layer6_outputs(1311));
    layer7_outputs(3632) <= (layer6_outputs(4677)) and not (layer6_outputs(2011));
    layer7_outputs(3633) <= not(layer6_outputs(1508));
    layer7_outputs(3634) <= not(layer6_outputs(424));
    layer7_outputs(3635) <= layer6_outputs(4693);
    layer7_outputs(3636) <= (layer6_outputs(146)) or (layer6_outputs(3698));
    layer7_outputs(3637) <= layer6_outputs(4525);
    layer7_outputs(3638) <= not(layer6_outputs(1563)) or (layer6_outputs(1378));
    layer7_outputs(3639) <= not(layer6_outputs(4907));
    layer7_outputs(3640) <= not(layer6_outputs(2112));
    layer7_outputs(3641) <= layer6_outputs(4387);
    layer7_outputs(3642) <= layer6_outputs(633);
    layer7_outputs(3643) <= layer6_outputs(2226);
    layer7_outputs(3644) <= '0';
    layer7_outputs(3645) <= not(layer6_outputs(1811));
    layer7_outputs(3646) <= not((layer6_outputs(3759)) xor (layer6_outputs(4042)));
    layer7_outputs(3647) <= '0';
    layer7_outputs(3648) <= not(layer6_outputs(3374));
    layer7_outputs(3649) <= not(layer6_outputs(1749));
    layer7_outputs(3650) <= not(layer6_outputs(3886));
    layer7_outputs(3651) <= not(layer6_outputs(4651));
    layer7_outputs(3652) <= (layer6_outputs(3767)) and (layer6_outputs(1907));
    layer7_outputs(3653) <= not(layer6_outputs(2610)) or (layer6_outputs(1382));
    layer7_outputs(3654) <= not((layer6_outputs(4141)) xor (layer6_outputs(3968)));
    layer7_outputs(3655) <= (layer6_outputs(3735)) and not (layer6_outputs(4845));
    layer7_outputs(3656) <= '1';
    layer7_outputs(3657) <= not(layer6_outputs(3044));
    layer7_outputs(3658) <= not(layer6_outputs(4929));
    layer7_outputs(3659) <= not(layer6_outputs(1016));
    layer7_outputs(3660) <= layer6_outputs(4972);
    layer7_outputs(3661) <= layer6_outputs(2259);
    layer7_outputs(3662) <= (layer6_outputs(4260)) and not (layer6_outputs(1513));
    layer7_outputs(3663) <= layer6_outputs(4584);
    layer7_outputs(3664) <= layer6_outputs(4591);
    layer7_outputs(3665) <= layer6_outputs(111);
    layer7_outputs(3666) <= (layer6_outputs(509)) or (layer6_outputs(2516));
    layer7_outputs(3667) <= layer6_outputs(603);
    layer7_outputs(3668) <= not(layer6_outputs(4432)) or (layer6_outputs(4608));
    layer7_outputs(3669) <= (layer6_outputs(1673)) and not (layer6_outputs(3523));
    layer7_outputs(3670) <= not((layer6_outputs(1555)) xor (layer6_outputs(1329)));
    layer7_outputs(3671) <= (layer6_outputs(101)) and not (layer6_outputs(1628));
    layer7_outputs(3672) <= layer6_outputs(2187);
    layer7_outputs(3673) <= layer6_outputs(4833);
    layer7_outputs(3674) <= '0';
    layer7_outputs(3675) <= not(layer6_outputs(5052));
    layer7_outputs(3676) <= not((layer6_outputs(3582)) xor (layer6_outputs(529)));
    layer7_outputs(3677) <= layer6_outputs(4967);
    layer7_outputs(3678) <= not(layer6_outputs(2652));
    layer7_outputs(3679) <= layer6_outputs(1634);
    layer7_outputs(3680) <= layer6_outputs(1583);
    layer7_outputs(3681) <= not(layer6_outputs(3270));
    layer7_outputs(3682) <= not((layer6_outputs(2698)) and (layer6_outputs(1879)));
    layer7_outputs(3683) <= not((layer6_outputs(4065)) and (layer6_outputs(2519)));
    layer7_outputs(3684) <= (layer6_outputs(2768)) or (layer6_outputs(1119));
    layer7_outputs(3685) <= not((layer6_outputs(2133)) and (layer6_outputs(1856)));
    layer7_outputs(3686) <= not(layer6_outputs(1148));
    layer7_outputs(3687) <= layer6_outputs(3584);
    layer7_outputs(3688) <= not(layer6_outputs(3444));
    layer7_outputs(3689) <= layer6_outputs(46);
    layer7_outputs(3690) <= not(layer6_outputs(5056));
    layer7_outputs(3691) <= not((layer6_outputs(605)) or (layer6_outputs(4761)));
    layer7_outputs(3692) <= not(layer6_outputs(3868)) or (layer6_outputs(4517));
    layer7_outputs(3693) <= (layer6_outputs(4577)) and (layer6_outputs(2277));
    layer7_outputs(3694) <= layer6_outputs(2123);
    layer7_outputs(3695) <= (layer6_outputs(468)) and (layer6_outputs(4753));
    layer7_outputs(3696) <= not((layer6_outputs(3141)) xor (layer6_outputs(2550)));
    layer7_outputs(3697) <= not(layer6_outputs(1467)) or (layer6_outputs(1661));
    layer7_outputs(3698) <= (layer6_outputs(3473)) xor (layer6_outputs(2958));
    layer7_outputs(3699) <= (layer6_outputs(1532)) and (layer6_outputs(1855));
    layer7_outputs(3700) <= layer6_outputs(2538);
    layer7_outputs(3701) <= not(layer6_outputs(4266)) or (layer6_outputs(764));
    layer7_outputs(3702) <= not((layer6_outputs(2733)) and (layer6_outputs(1736)));
    layer7_outputs(3703) <= not((layer6_outputs(4148)) and (layer6_outputs(2608)));
    layer7_outputs(3704) <= not((layer6_outputs(1914)) and (layer6_outputs(2753)));
    layer7_outputs(3705) <= (layer6_outputs(391)) xor (layer6_outputs(3195));
    layer7_outputs(3706) <= (layer6_outputs(1750)) and not (layer6_outputs(1764));
    layer7_outputs(3707) <= (layer6_outputs(3882)) xor (layer6_outputs(2786));
    layer7_outputs(3708) <= not(layer6_outputs(279));
    layer7_outputs(3709) <= (layer6_outputs(3398)) xor (layer6_outputs(1469));
    layer7_outputs(3710) <= not(layer6_outputs(1565));
    layer7_outputs(3711) <= not(layer6_outputs(2852));
    layer7_outputs(3712) <= layer6_outputs(1350);
    layer7_outputs(3713) <= not(layer6_outputs(2169));
    layer7_outputs(3714) <= not((layer6_outputs(5113)) xor (layer6_outputs(1373)));
    layer7_outputs(3715) <= '0';
    layer7_outputs(3716) <= not(layer6_outputs(2160)) or (layer6_outputs(1560));
    layer7_outputs(3717) <= not((layer6_outputs(4539)) xor (layer6_outputs(1356)));
    layer7_outputs(3718) <= (layer6_outputs(1211)) and (layer6_outputs(3251));
    layer7_outputs(3719) <= (layer6_outputs(607)) xor (layer6_outputs(2566));
    layer7_outputs(3720) <= (layer6_outputs(3236)) and not (layer6_outputs(1818));
    layer7_outputs(3721) <= not(layer6_outputs(763));
    layer7_outputs(3722) <= layer6_outputs(1261);
    layer7_outputs(3723) <= (layer6_outputs(2743)) and not (layer6_outputs(4969));
    layer7_outputs(3724) <= (layer6_outputs(424)) xor (layer6_outputs(4827));
    layer7_outputs(3725) <= not(layer6_outputs(1413));
    layer7_outputs(3726) <= (layer6_outputs(4559)) and (layer6_outputs(3045));
    layer7_outputs(3727) <= layer6_outputs(5094);
    layer7_outputs(3728) <= not(layer6_outputs(1572));
    layer7_outputs(3729) <= not(layer6_outputs(1144));
    layer7_outputs(3730) <= '0';
    layer7_outputs(3731) <= not(layer6_outputs(590));
    layer7_outputs(3732) <= not(layer6_outputs(3780)) or (layer6_outputs(2420));
    layer7_outputs(3733) <= layer6_outputs(4284);
    layer7_outputs(3734) <= layer6_outputs(4691);
    layer7_outputs(3735) <= not((layer6_outputs(1626)) and (layer6_outputs(3243)));
    layer7_outputs(3736) <= not(layer6_outputs(3960));
    layer7_outputs(3737) <= '1';
    layer7_outputs(3738) <= not(layer6_outputs(4823)) or (layer6_outputs(1134));
    layer7_outputs(3739) <= layer6_outputs(4683);
    layer7_outputs(3740) <= (layer6_outputs(2344)) and (layer6_outputs(3142));
    layer7_outputs(3741) <= '0';
    layer7_outputs(3742) <= (layer6_outputs(2039)) and not (layer6_outputs(2364));
    layer7_outputs(3743) <= (layer6_outputs(3113)) and (layer6_outputs(5087));
    layer7_outputs(3744) <= (layer6_outputs(5091)) and not (layer6_outputs(3454));
    layer7_outputs(3745) <= (layer6_outputs(5079)) and (layer6_outputs(40));
    layer7_outputs(3746) <= layer6_outputs(2976);
    layer7_outputs(3747) <= not(layer6_outputs(2249));
    layer7_outputs(3748) <= (layer6_outputs(691)) and (layer6_outputs(385));
    layer7_outputs(3749) <= not((layer6_outputs(900)) or (layer6_outputs(2509)));
    layer7_outputs(3750) <= (layer6_outputs(3635)) and (layer6_outputs(1942));
    layer7_outputs(3751) <= layer6_outputs(4285);
    layer7_outputs(3752) <= (layer6_outputs(4841)) and not (layer6_outputs(1963));
    layer7_outputs(3753) <= (layer6_outputs(1801)) or (layer6_outputs(1098));
    layer7_outputs(3754) <= not(layer6_outputs(1566)) or (layer6_outputs(104));
    layer7_outputs(3755) <= not(layer6_outputs(874));
    layer7_outputs(3756) <= layer6_outputs(878);
    layer7_outputs(3757) <= not(layer6_outputs(3536));
    layer7_outputs(3758) <= not(layer6_outputs(3832)) or (layer6_outputs(2970));
    layer7_outputs(3759) <= layer6_outputs(1537);
    layer7_outputs(3760) <= layer6_outputs(4268);
    layer7_outputs(3761) <= (layer6_outputs(5006)) and not (layer6_outputs(5112));
    layer7_outputs(3762) <= layer6_outputs(381);
    layer7_outputs(3763) <= layer6_outputs(698);
    layer7_outputs(3764) <= not(layer6_outputs(4295));
    layer7_outputs(3765) <= not(layer6_outputs(1581)) or (layer6_outputs(2255));
    layer7_outputs(3766) <= layer6_outputs(1844);
    layer7_outputs(3767) <= not(layer6_outputs(3669));
    layer7_outputs(3768) <= (layer6_outputs(209)) and (layer6_outputs(2140));
    layer7_outputs(3769) <= not(layer6_outputs(1835));
    layer7_outputs(3770) <= not(layer6_outputs(4802));
    layer7_outputs(3771) <= layer6_outputs(1481);
    layer7_outputs(3772) <= not(layer6_outputs(3815)) or (layer6_outputs(953));
    layer7_outputs(3773) <= layer6_outputs(3782);
    layer7_outputs(3774) <= not(layer6_outputs(5057));
    layer7_outputs(3775) <= not((layer6_outputs(2636)) xor (layer6_outputs(1649)));
    layer7_outputs(3776) <= layer6_outputs(1667);
    layer7_outputs(3777) <= not(layer6_outputs(1204));
    layer7_outputs(3778) <= layer6_outputs(151);
    layer7_outputs(3779) <= not(layer6_outputs(271)) or (layer6_outputs(179));
    layer7_outputs(3780) <= not(layer6_outputs(4234)) or (layer6_outputs(2497));
    layer7_outputs(3781) <= layer6_outputs(2480);
    layer7_outputs(3782) <= not((layer6_outputs(1220)) or (layer6_outputs(1828)));
    layer7_outputs(3783) <= layer6_outputs(168);
    layer7_outputs(3784) <= layer6_outputs(3849);
    layer7_outputs(3785) <= not(layer6_outputs(4236));
    layer7_outputs(3786) <= not((layer6_outputs(1072)) or (layer6_outputs(1217)));
    layer7_outputs(3787) <= (layer6_outputs(2390)) or (layer6_outputs(4851));
    layer7_outputs(3788) <= not(layer6_outputs(4130));
    layer7_outputs(3789) <= not((layer6_outputs(1265)) xor (layer6_outputs(2998)));
    layer7_outputs(3790) <= layer6_outputs(2448);
    layer7_outputs(3791) <= layer6_outputs(3271);
    layer7_outputs(3792) <= not(layer6_outputs(1136));
    layer7_outputs(3793) <= (layer6_outputs(1977)) or (layer6_outputs(571));
    layer7_outputs(3794) <= not(layer6_outputs(3307));
    layer7_outputs(3795) <= not(layer6_outputs(3907));
    layer7_outputs(3796) <= (layer6_outputs(3683)) and not (layer6_outputs(1672));
    layer7_outputs(3797) <= not((layer6_outputs(4068)) xor (layer6_outputs(3727)));
    layer7_outputs(3798) <= not(layer6_outputs(1653));
    layer7_outputs(3799) <= layer6_outputs(513);
    layer7_outputs(3800) <= (layer6_outputs(3540)) and not (layer6_outputs(1348));
    layer7_outputs(3801) <= not((layer6_outputs(2672)) xor (layer6_outputs(2844)));
    layer7_outputs(3802) <= (layer6_outputs(2956)) and not (layer6_outputs(1948));
    layer7_outputs(3803) <= layer6_outputs(5098);
    layer7_outputs(3804) <= layer6_outputs(820);
    layer7_outputs(3805) <= not(layer6_outputs(4195));
    layer7_outputs(3806) <= not(layer6_outputs(1473));
    layer7_outputs(3807) <= not((layer6_outputs(1602)) and (layer6_outputs(2981)));
    layer7_outputs(3808) <= layer6_outputs(3808);
    layer7_outputs(3809) <= (layer6_outputs(2586)) and not (layer6_outputs(2647));
    layer7_outputs(3810) <= not((layer6_outputs(4195)) xor (layer6_outputs(1875)));
    layer7_outputs(3811) <= not(layer6_outputs(4742));
    layer7_outputs(3812) <= not(layer6_outputs(3273));
    layer7_outputs(3813) <= not(layer6_outputs(2837));
    layer7_outputs(3814) <= '1';
    layer7_outputs(3815) <= layer6_outputs(3996);
    layer7_outputs(3816) <= not((layer6_outputs(3948)) or (layer6_outputs(526)));
    layer7_outputs(3817) <= layer6_outputs(971);
    layer7_outputs(3818) <= '0';
    layer7_outputs(3819) <= not(layer6_outputs(3456));
    layer7_outputs(3820) <= not(layer6_outputs(3904));
    layer7_outputs(3821) <= not(layer6_outputs(3919)) or (layer6_outputs(870));
    layer7_outputs(3822) <= (layer6_outputs(1622)) and not (layer6_outputs(612));
    layer7_outputs(3823) <= '1';
    layer7_outputs(3824) <= layer6_outputs(1506);
    layer7_outputs(3825) <= (layer6_outputs(2091)) xor (layer6_outputs(317));
    layer7_outputs(3826) <= layer6_outputs(1796);
    layer7_outputs(3827) <= layer6_outputs(4858);
    layer7_outputs(3828) <= layer6_outputs(3798);
    layer7_outputs(3829) <= not(layer6_outputs(1141));
    layer7_outputs(3830) <= (layer6_outputs(4110)) and (layer6_outputs(891));
    layer7_outputs(3831) <= not(layer6_outputs(2191));
    layer7_outputs(3832) <= not((layer6_outputs(2266)) xor (layer6_outputs(3900)));
    layer7_outputs(3833) <= (layer6_outputs(2128)) and (layer6_outputs(4710));
    layer7_outputs(3834) <= not(layer6_outputs(1265)) or (layer6_outputs(3037));
    layer7_outputs(3835) <= not((layer6_outputs(1208)) xor (layer6_outputs(2866)));
    layer7_outputs(3836) <= not(layer6_outputs(1932));
    layer7_outputs(3837) <= '1';
    layer7_outputs(3838) <= layer6_outputs(1201);
    layer7_outputs(3839) <= (layer6_outputs(4949)) xor (layer6_outputs(2757));
    layer7_outputs(3840) <= not(layer6_outputs(1348));
    layer7_outputs(3841) <= not(layer6_outputs(1046));
    layer7_outputs(3842) <= layer6_outputs(1603);
    layer7_outputs(3843) <= not((layer6_outputs(942)) xor (layer6_outputs(3707)));
    layer7_outputs(3844) <= layer6_outputs(2761);
    layer7_outputs(3845) <= not(layer6_outputs(3757));
    layer7_outputs(3846) <= (layer6_outputs(3465)) and not (layer6_outputs(3603));
    layer7_outputs(3847) <= not(layer6_outputs(395));
    layer7_outputs(3848) <= (layer6_outputs(3589)) and (layer6_outputs(2467));
    layer7_outputs(3849) <= (layer6_outputs(3697)) and (layer6_outputs(489));
    layer7_outputs(3850) <= (layer6_outputs(63)) or (layer6_outputs(1367));
    layer7_outputs(3851) <= not((layer6_outputs(1666)) or (layer6_outputs(1577)));
    layer7_outputs(3852) <= not(layer6_outputs(4267));
    layer7_outputs(3853) <= not((layer6_outputs(4091)) and (layer6_outputs(749)));
    layer7_outputs(3854) <= layer6_outputs(3492);
    layer7_outputs(3855) <= layer6_outputs(3411);
    layer7_outputs(3856) <= not((layer6_outputs(738)) and (layer6_outputs(1701)));
    layer7_outputs(3857) <= layer6_outputs(1358);
    layer7_outputs(3858) <= not(layer6_outputs(1030));
    layer7_outputs(3859) <= layer6_outputs(407);
    layer7_outputs(3860) <= '0';
    layer7_outputs(3861) <= not(layer6_outputs(427));
    layer7_outputs(3862) <= (layer6_outputs(4600)) xor (layer6_outputs(3619));
    layer7_outputs(3863) <= not(layer6_outputs(148));
    layer7_outputs(3864) <= layer6_outputs(1268);
    layer7_outputs(3865) <= (layer6_outputs(1407)) or (layer6_outputs(2288));
    layer7_outputs(3866) <= not(layer6_outputs(2275));
    layer7_outputs(3867) <= not((layer6_outputs(510)) xor (layer6_outputs(4822)));
    layer7_outputs(3868) <= (layer6_outputs(1432)) and not (layer6_outputs(1397));
    layer7_outputs(3869) <= not(layer6_outputs(1210));
    layer7_outputs(3870) <= not((layer6_outputs(2320)) or (layer6_outputs(4519)));
    layer7_outputs(3871) <= layer6_outputs(3658);
    layer7_outputs(3872) <= layer6_outputs(2439);
    layer7_outputs(3873) <= not(layer6_outputs(166));
    layer7_outputs(3874) <= not(layer6_outputs(4573));
    layer7_outputs(3875) <= (layer6_outputs(4074)) xor (layer6_outputs(3157));
    layer7_outputs(3876) <= not((layer6_outputs(3537)) and (layer6_outputs(3088)));
    layer7_outputs(3877) <= not((layer6_outputs(2810)) and (layer6_outputs(3167)));
    layer7_outputs(3878) <= not((layer6_outputs(1693)) xor (layer6_outputs(4639)));
    layer7_outputs(3879) <= (layer6_outputs(4421)) and (layer6_outputs(703));
    layer7_outputs(3880) <= layer6_outputs(2500);
    layer7_outputs(3881) <= layer6_outputs(4564);
    layer7_outputs(3882) <= not(layer6_outputs(2552));
    layer7_outputs(3883) <= layer6_outputs(850);
    layer7_outputs(3884) <= layer6_outputs(105);
    layer7_outputs(3885) <= not((layer6_outputs(1993)) xor (layer6_outputs(615)));
    layer7_outputs(3886) <= (layer6_outputs(5038)) xor (layer6_outputs(1197));
    layer7_outputs(3887) <= layer6_outputs(4686);
    layer7_outputs(3888) <= not((layer6_outputs(1820)) xor (layer6_outputs(4427)));
    layer7_outputs(3889) <= not(layer6_outputs(5098));
    layer7_outputs(3890) <= layer6_outputs(2544);
    layer7_outputs(3891) <= not(layer6_outputs(4506)) or (layer6_outputs(3995));
    layer7_outputs(3892) <= not(layer6_outputs(1267));
    layer7_outputs(3893) <= (layer6_outputs(1280)) and (layer6_outputs(565));
    layer7_outputs(3894) <= not(layer6_outputs(3485)) or (layer6_outputs(4286));
    layer7_outputs(3895) <= not(layer6_outputs(2100));
    layer7_outputs(3896) <= layer6_outputs(542);
    layer7_outputs(3897) <= not(layer6_outputs(3862));
    layer7_outputs(3898) <= '0';
    layer7_outputs(3899) <= layer6_outputs(2245);
    layer7_outputs(3900) <= not((layer6_outputs(4368)) xor (layer6_outputs(4459)));
    layer7_outputs(3901) <= not(layer6_outputs(3955));
    layer7_outputs(3902) <= layer6_outputs(1146);
    layer7_outputs(3903) <= layer6_outputs(1404);
    layer7_outputs(3904) <= layer6_outputs(3546);
    layer7_outputs(3905) <= layer6_outputs(1174);
    layer7_outputs(3906) <= layer6_outputs(3505);
    layer7_outputs(3907) <= not(layer6_outputs(4921));
    layer7_outputs(3908) <= layer6_outputs(282);
    layer7_outputs(3909) <= (layer6_outputs(2129)) xor (layer6_outputs(4808));
    layer7_outputs(3910) <= not((layer6_outputs(3224)) and (layer6_outputs(1948)));
    layer7_outputs(3911) <= (layer6_outputs(4489)) xor (layer6_outputs(1500));
    layer7_outputs(3912) <= not(layer6_outputs(3456)) or (layer6_outputs(1344));
    layer7_outputs(3913) <= not((layer6_outputs(3782)) xor (layer6_outputs(3153)));
    layer7_outputs(3914) <= layer6_outputs(1874);
    layer7_outputs(3915) <= not(layer6_outputs(737));
    layer7_outputs(3916) <= not(layer6_outputs(3466));
    layer7_outputs(3917) <= layer6_outputs(1864);
    layer7_outputs(3918) <= (layer6_outputs(886)) and not (layer6_outputs(1202));
    layer7_outputs(3919) <= (layer6_outputs(4619)) and (layer6_outputs(2169));
    layer7_outputs(3920) <= layer6_outputs(1625);
    layer7_outputs(3921) <= layer6_outputs(4120);
    layer7_outputs(3922) <= not(layer6_outputs(1823));
    layer7_outputs(3923) <= layer6_outputs(2560);
    layer7_outputs(3924) <= layer6_outputs(4898);
    layer7_outputs(3925) <= not(layer6_outputs(3252));
    layer7_outputs(3926) <= not(layer6_outputs(4321));
    layer7_outputs(3927) <= not((layer6_outputs(4122)) xor (layer6_outputs(2706)));
    layer7_outputs(3928) <= (layer6_outputs(4923)) xor (layer6_outputs(185));
    layer7_outputs(3929) <= layer6_outputs(2646);
    layer7_outputs(3930) <= not(layer6_outputs(2038));
    layer7_outputs(3931) <= not((layer6_outputs(5093)) xor (layer6_outputs(1055)));
    layer7_outputs(3932) <= not(layer6_outputs(37));
    layer7_outputs(3933) <= not(layer6_outputs(3248));
    layer7_outputs(3934) <= (layer6_outputs(4123)) and not (layer6_outputs(486));
    layer7_outputs(3935) <= (layer6_outputs(2597)) and not (layer6_outputs(1007));
    layer7_outputs(3936) <= not((layer6_outputs(1178)) and (layer6_outputs(3949)));
    layer7_outputs(3937) <= (layer6_outputs(232)) and (layer6_outputs(1179));
    layer7_outputs(3938) <= not(layer6_outputs(4036));
    layer7_outputs(3939) <= not((layer6_outputs(2945)) xor (layer6_outputs(1568)));
    layer7_outputs(3940) <= (layer6_outputs(2351)) or (layer6_outputs(4874));
    layer7_outputs(3941) <= layer6_outputs(1966);
    layer7_outputs(3942) <= not(layer6_outputs(304));
    layer7_outputs(3943) <= not((layer6_outputs(2188)) and (layer6_outputs(1842)));
    layer7_outputs(3944) <= not(layer6_outputs(766));
    layer7_outputs(3945) <= not((layer6_outputs(1756)) xor (layer6_outputs(3501)));
    layer7_outputs(3946) <= layer6_outputs(1710);
    layer7_outputs(3947) <= not(layer6_outputs(5088));
    layer7_outputs(3948) <= (layer6_outputs(3013)) and not (layer6_outputs(3326));
    layer7_outputs(3949) <= (layer6_outputs(1795)) and not (layer6_outputs(3415));
    layer7_outputs(3950) <= layer6_outputs(3447);
    layer7_outputs(3951) <= (layer6_outputs(4033)) xor (layer6_outputs(2645));
    layer7_outputs(3952) <= layer6_outputs(3890);
    layer7_outputs(3953) <= (layer6_outputs(1047)) and not (layer6_outputs(2128));
    layer7_outputs(3954) <= not((layer6_outputs(3002)) or (layer6_outputs(2210)));
    layer7_outputs(3955) <= not(layer6_outputs(2060));
    layer7_outputs(3956) <= not((layer6_outputs(199)) xor (layer6_outputs(2891)));
    layer7_outputs(3957) <= (layer6_outputs(2677)) and not (layer6_outputs(3225));
    layer7_outputs(3958) <= layer6_outputs(1417);
    layer7_outputs(3959) <= not((layer6_outputs(1936)) and (layer6_outputs(866)));
    layer7_outputs(3960) <= not(layer6_outputs(2491));
    layer7_outputs(3961) <= not(layer6_outputs(5067));
    layer7_outputs(3962) <= layer6_outputs(3846);
    layer7_outputs(3963) <= layer6_outputs(551);
    layer7_outputs(3964) <= not(layer6_outputs(2597));
    layer7_outputs(3965) <= layer6_outputs(3513);
    layer7_outputs(3966) <= (layer6_outputs(1108)) and (layer6_outputs(2448));
    layer7_outputs(3967) <= not(layer6_outputs(4122));
    layer7_outputs(3968) <= (layer6_outputs(483)) and not (layer6_outputs(3767));
    layer7_outputs(3969) <= not(layer6_outputs(1368)) or (layer6_outputs(4269));
    layer7_outputs(3970) <= not(layer6_outputs(2790));
    layer7_outputs(3971) <= not(layer6_outputs(4760));
    layer7_outputs(3972) <= not(layer6_outputs(600)) or (layer6_outputs(2096));
    layer7_outputs(3973) <= not((layer6_outputs(1377)) and (layer6_outputs(1677)));
    layer7_outputs(3974) <= (layer6_outputs(2527)) and (layer6_outputs(547));
    layer7_outputs(3975) <= not(layer6_outputs(1346)) or (layer6_outputs(485));
    layer7_outputs(3976) <= '1';
    layer7_outputs(3977) <= (layer6_outputs(2986)) and not (layer6_outputs(2637));
    layer7_outputs(3978) <= layer6_outputs(4938);
    layer7_outputs(3979) <= layer6_outputs(2252);
    layer7_outputs(3980) <= not(layer6_outputs(4724));
    layer7_outputs(3981) <= layer6_outputs(610);
    layer7_outputs(3982) <= not(layer6_outputs(4822));
    layer7_outputs(3983) <= not(layer6_outputs(1099)) or (layer6_outputs(4023));
    layer7_outputs(3984) <= '1';
    layer7_outputs(3985) <= not((layer6_outputs(750)) or (layer6_outputs(3436)));
    layer7_outputs(3986) <= not((layer6_outputs(3048)) and (layer6_outputs(3212)));
    layer7_outputs(3987) <= (layer6_outputs(3432)) and (layer6_outputs(527));
    layer7_outputs(3988) <= not((layer6_outputs(728)) xor (layer6_outputs(708)));
    layer7_outputs(3989) <= (layer6_outputs(2988)) and not (layer6_outputs(4986));
    layer7_outputs(3990) <= (layer6_outputs(1920)) and not (layer6_outputs(2737));
    layer7_outputs(3991) <= not(layer6_outputs(2));
    layer7_outputs(3992) <= not((layer6_outputs(4684)) or (layer6_outputs(4051)));
    layer7_outputs(3993) <= not((layer6_outputs(2148)) xor (layer6_outputs(3842)));
    layer7_outputs(3994) <= not(layer6_outputs(2973)) or (layer6_outputs(1898));
    layer7_outputs(3995) <= layer6_outputs(2539);
    layer7_outputs(3996) <= not((layer6_outputs(3927)) and (layer6_outputs(4483)));
    layer7_outputs(3997) <= layer6_outputs(590);
    layer7_outputs(3998) <= layer6_outputs(2808);
    layer7_outputs(3999) <= not((layer6_outputs(5104)) xor (layer6_outputs(2778)));
    layer7_outputs(4000) <= (layer6_outputs(4417)) xor (layer6_outputs(454));
    layer7_outputs(4001) <= not(layer6_outputs(3203));
    layer7_outputs(4002) <= layer6_outputs(722);
    layer7_outputs(4003) <= not(layer6_outputs(157));
    layer7_outputs(4004) <= not(layer6_outputs(4370));
    layer7_outputs(4005) <= not(layer6_outputs(4668));
    layer7_outputs(4006) <= (layer6_outputs(1171)) xor (layer6_outputs(3285));
    layer7_outputs(4007) <= not(layer6_outputs(129)) or (layer6_outputs(2729));
    layer7_outputs(4008) <= not(layer6_outputs(3208)) or (layer6_outputs(646));
    layer7_outputs(4009) <= (layer6_outputs(3453)) and not (layer6_outputs(2093));
    layer7_outputs(4010) <= not(layer6_outputs(3175));
    layer7_outputs(4011) <= not(layer6_outputs(4882));
    layer7_outputs(4012) <= layer6_outputs(2395);
    layer7_outputs(4013) <= layer6_outputs(4182);
    layer7_outputs(4014) <= not((layer6_outputs(3842)) and (layer6_outputs(4575)));
    layer7_outputs(4015) <= not((layer6_outputs(990)) or (layer6_outputs(4955)));
    layer7_outputs(4016) <= not(layer6_outputs(1813));
    layer7_outputs(4017) <= '0';
    layer7_outputs(4018) <= layer6_outputs(1863);
    layer7_outputs(4019) <= layer6_outputs(2158);
    layer7_outputs(4020) <= layer6_outputs(116);
    layer7_outputs(4021) <= not(layer6_outputs(1832));
    layer7_outputs(4022) <= layer6_outputs(4798);
    layer7_outputs(4023) <= layer6_outputs(4169);
    layer7_outputs(4024) <= not(layer6_outputs(4454));
    layer7_outputs(4025) <= not(layer6_outputs(2066));
    layer7_outputs(4026) <= (layer6_outputs(2025)) and not (layer6_outputs(4228));
    layer7_outputs(4027) <= (layer6_outputs(4062)) or (layer6_outputs(3014));
    layer7_outputs(4028) <= layer6_outputs(1910);
    layer7_outputs(4029) <= layer6_outputs(3750);
    layer7_outputs(4030) <= not(layer6_outputs(3459));
    layer7_outputs(4031) <= not(layer6_outputs(2987)) or (layer6_outputs(5076));
    layer7_outputs(4032) <= (layer6_outputs(3385)) or (layer6_outputs(1953));
    layer7_outputs(4033) <= layer6_outputs(91);
    layer7_outputs(4034) <= not(layer6_outputs(4138));
    layer7_outputs(4035) <= layer6_outputs(2728);
    layer7_outputs(4036) <= not(layer6_outputs(3093)) or (layer6_outputs(4765));
    layer7_outputs(4037) <= layer6_outputs(332);
    layer7_outputs(4038) <= not(layer6_outputs(4291));
    layer7_outputs(4039) <= not(layer6_outputs(4062));
    layer7_outputs(4040) <= (layer6_outputs(2103)) and (layer6_outputs(5029));
    layer7_outputs(4041) <= not(layer6_outputs(2832));
    layer7_outputs(4042) <= (layer6_outputs(1955)) and (layer6_outputs(3169));
    layer7_outputs(4043) <= (layer6_outputs(907)) and not (layer6_outputs(685));
    layer7_outputs(4044) <= layer6_outputs(81);
    layer7_outputs(4045) <= (layer6_outputs(3313)) and not (layer6_outputs(4281));
    layer7_outputs(4046) <= (layer6_outputs(2836)) or (layer6_outputs(372));
    layer7_outputs(4047) <= not((layer6_outputs(2281)) or (layer6_outputs(3738)));
    layer7_outputs(4048) <= not(layer6_outputs(4433));
    layer7_outputs(4049) <= not(layer6_outputs(275)) or (layer6_outputs(1383));
    layer7_outputs(4050) <= not(layer6_outputs(411)) or (layer6_outputs(2453));
    layer7_outputs(4051) <= layer6_outputs(2826);
    layer7_outputs(4052) <= not((layer6_outputs(1240)) or (layer6_outputs(3498)));
    layer7_outputs(4053) <= not(layer6_outputs(32));
    layer7_outputs(4054) <= (layer6_outputs(3323)) xor (layer6_outputs(2899));
    layer7_outputs(4055) <= not(layer6_outputs(2418)) or (layer6_outputs(5074));
    layer7_outputs(4056) <= not(layer6_outputs(3775));
    layer7_outputs(4057) <= layer6_outputs(945);
    layer7_outputs(4058) <= layer6_outputs(708);
    layer7_outputs(4059) <= not(layer6_outputs(4980)) or (layer6_outputs(3496));
    layer7_outputs(4060) <= not((layer6_outputs(4389)) or (layer6_outputs(3528)));
    layer7_outputs(4061) <= layer6_outputs(871);
    layer7_outputs(4062) <= (layer6_outputs(3477)) and not (layer6_outputs(4493));
    layer7_outputs(4063) <= (layer6_outputs(2144)) xor (layer6_outputs(3617));
    layer7_outputs(4064) <= layer6_outputs(2338);
    layer7_outputs(4065) <= not(layer6_outputs(4013));
    layer7_outputs(4066) <= layer6_outputs(3566);
    layer7_outputs(4067) <= not(layer6_outputs(3367));
    layer7_outputs(4068) <= not(layer6_outputs(3644));
    layer7_outputs(4069) <= not(layer6_outputs(3064)) or (layer6_outputs(4899));
    layer7_outputs(4070) <= layer6_outputs(2848);
    layer7_outputs(4071) <= not(layer6_outputs(1769));
    layer7_outputs(4072) <= not(layer6_outputs(1679));
    layer7_outputs(4073) <= not(layer6_outputs(5108));
    layer7_outputs(4074) <= not(layer6_outputs(913)) or (layer6_outputs(2561));
    layer7_outputs(4075) <= not(layer6_outputs(1179));
    layer7_outputs(4076) <= layer6_outputs(2355);
    layer7_outputs(4077) <= layer6_outputs(789);
    layer7_outputs(4078) <= not(layer6_outputs(549));
    layer7_outputs(4079) <= not((layer6_outputs(1145)) xor (layer6_outputs(1587)));
    layer7_outputs(4080) <= not(layer6_outputs(371)) or (layer6_outputs(1540));
    layer7_outputs(4081) <= (layer6_outputs(931)) and not (layer6_outputs(1678));
    layer7_outputs(4082) <= (layer6_outputs(4109)) xor (layer6_outputs(4046));
    layer7_outputs(4083) <= not((layer6_outputs(4064)) xor (layer6_outputs(3351)));
    layer7_outputs(4084) <= not(layer6_outputs(4836));
    layer7_outputs(4085) <= (layer6_outputs(1195)) and not (layer6_outputs(3264));
    layer7_outputs(4086) <= (layer6_outputs(4354)) xor (layer6_outputs(4058));
    layer7_outputs(4087) <= not((layer6_outputs(1808)) and (layer6_outputs(3811)));
    layer7_outputs(4088) <= (layer6_outputs(4325)) or (layer6_outputs(4450));
    layer7_outputs(4089) <= layer6_outputs(1614);
    layer7_outputs(4090) <= not(layer6_outputs(3555));
    layer7_outputs(4091) <= (layer6_outputs(2195)) or (layer6_outputs(1502));
    layer7_outputs(4092) <= layer6_outputs(384);
    layer7_outputs(4093) <= not(layer6_outputs(4098));
    layer7_outputs(4094) <= layer6_outputs(537);
    layer7_outputs(4095) <= layer6_outputs(420);
    layer7_outputs(4096) <= not((layer6_outputs(1249)) and (layer6_outputs(2139)));
    layer7_outputs(4097) <= layer6_outputs(1523);
    layer7_outputs(4098) <= (layer6_outputs(1716)) or (layer6_outputs(2707));
    layer7_outputs(4099) <= layer6_outputs(4231);
    layer7_outputs(4100) <= layer6_outputs(3124);
    layer7_outputs(4101) <= not(layer6_outputs(242));
    layer7_outputs(4102) <= not((layer6_outputs(2388)) xor (layer6_outputs(4170)));
    layer7_outputs(4103) <= not((layer6_outputs(4976)) or (layer6_outputs(2666)));
    layer7_outputs(4104) <= layer6_outputs(3006);
    layer7_outputs(4105) <= layer6_outputs(244);
    layer7_outputs(4106) <= not((layer6_outputs(2767)) and (layer6_outputs(758)));
    layer7_outputs(4107) <= not((layer6_outputs(84)) or (layer6_outputs(3890)));
    layer7_outputs(4108) <= layer6_outputs(3652);
    layer7_outputs(4109) <= not((layer6_outputs(5040)) or (layer6_outputs(4959)));
    layer7_outputs(4110) <= (layer6_outputs(703)) and not (layer6_outputs(4862));
    layer7_outputs(4111) <= not(layer6_outputs(3358));
    layer7_outputs(4112) <= not((layer6_outputs(26)) or (layer6_outputs(4356)));
    layer7_outputs(4113) <= (layer6_outputs(608)) and not (layer6_outputs(2481));
    layer7_outputs(4114) <= not((layer6_outputs(203)) and (layer6_outputs(3519)));
    layer7_outputs(4115) <= not((layer6_outputs(3947)) and (layer6_outputs(1861)));
    layer7_outputs(4116) <= not(layer6_outputs(3419)) or (layer6_outputs(1207));
    layer7_outputs(4117) <= not((layer6_outputs(4003)) and (layer6_outputs(4799)));
    layer7_outputs(4118) <= not(layer6_outputs(2251));
    layer7_outputs(4119) <= (layer6_outputs(2432)) xor (layer6_outputs(776));
    layer7_outputs(4120) <= layer6_outputs(926);
    layer7_outputs(4121) <= (layer6_outputs(4450)) and not (layer6_outputs(2247));
    layer7_outputs(4122) <= not((layer6_outputs(3508)) or (layer6_outputs(1066)));
    layer7_outputs(4123) <= not(layer6_outputs(345));
    layer7_outputs(4124) <= layer6_outputs(2680);
    layer7_outputs(4125) <= not(layer6_outputs(1991)) or (layer6_outputs(3447));
    layer7_outputs(4126) <= not(layer6_outputs(2789)) or (layer6_outputs(1556));
    layer7_outputs(4127) <= (layer6_outputs(3988)) or (layer6_outputs(2155));
    layer7_outputs(4128) <= not(layer6_outputs(3718)) or (layer6_outputs(734));
    layer7_outputs(4129) <= layer6_outputs(3833);
    layer7_outputs(4130) <= not(layer6_outputs(2531));
    layer7_outputs(4131) <= not((layer6_outputs(2356)) xor (layer6_outputs(1072)));
    layer7_outputs(4132) <= not(layer6_outputs(1292));
    layer7_outputs(4133) <= not(layer6_outputs(510)) or (layer6_outputs(560));
    layer7_outputs(4134) <= not(layer6_outputs(4043));
    layer7_outputs(4135) <= (layer6_outputs(3298)) xor (layer6_outputs(4880));
    layer7_outputs(4136) <= not(layer6_outputs(3470));
    layer7_outputs(4137) <= not(layer6_outputs(4607));
    layer7_outputs(4138) <= not(layer6_outputs(1560));
    layer7_outputs(4139) <= layer6_outputs(3266);
    layer7_outputs(4140) <= layer6_outputs(2454);
    layer7_outputs(4141) <= not((layer6_outputs(598)) or (layer6_outputs(2623)));
    layer7_outputs(4142) <= not((layer6_outputs(98)) or (layer6_outputs(4174)));
    layer7_outputs(4143) <= not(layer6_outputs(2599));
    layer7_outputs(4144) <= not(layer6_outputs(5079));
    layer7_outputs(4145) <= (layer6_outputs(783)) and not (layer6_outputs(1825));
    layer7_outputs(4146) <= not((layer6_outputs(806)) and (layer6_outputs(3868)));
    layer7_outputs(4147) <= not(layer6_outputs(3585));
    layer7_outputs(4148) <= layer6_outputs(13);
    layer7_outputs(4149) <= not(layer6_outputs(1944)) or (layer6_outputs(4936));
    layer7_outputs(4150) <= not(layer6_outputs(3365));
    layer7_outputs(4151) <= '0';
    layer7_outputs(4152) <= (layer6_outputs(1174)) xor (layer6_outputs(1173));
    layer7_outputs(4153) <= not(layer6_outputs(1571));
    layer7_outputs(4154) <= not(layer6_outputs(4342));
    layer7_outputs(4155) <= (layer6_outputs(3701)) xor (layer6_outputs(3743));
    layer7_outputs(4156) <= layer6_outputs(2580);
    layer7_outputs(4157) <= not((layer6_outputs(3369)) and (layer6_outputs(2731)));
    layer7_outputs(4158) <= not((layer6_outputs(2095)) xor (layer6_outputs(1469)));
    layer7_outputs(4159) <= not((layer6_outputs(1700)) xor (layer6_outputs(1979)));
    layer7_outputs(4160) <= not((layer6_outputs(3652)) xor (layer6_outputs(4027)));
    layer7_outputs(4161) <= layer6_outputs(4518);
    layer7_outputs(4162) <= not(layer6_outputs(4129));
    layer7_outputs(4163) <= '0';
    layer7_outputs(4164) <= (layer6_outputs(2983)) and (layer6_outputs(1448));
    layer7_outputs(4165) <= (layer6_outputs(1209)) or (layer6_outputs(281));
    layer7_outputs(4166) <= not(layer6_outputs(771));
    layer7_outputs(4167) <= not((layer6_outputs(4712)) xor (layer6_outputs(4961)));
    layer7_outputs(4168) <= not(layer6_outputs(5062));
    layer7_outputs(4169) <= (layer6_outputs(3747)) and not (layer6_outputs(1464));
    layer7_outputs(4170) <= layer6_outputs(1371);
    layer7_outputs(4171) <= layer6_outputs(804);
    layer7_outputs(4172) <= (layer6_outputs(4272)) and (layer6_outputs(3603));
    layer7_outputs(4173) <= (layer6_outputs(5094)) xor (layer6_outputs(860));
    layer7_outputs(4174) <= not(layer6_outputs(1293)) or (layer6_outputs(1090));
    layer7_outputs(4175) <= (layer6_outputs(1882)) and not (layer6_outputs(2645));
    layer7_outputs(4176) <= not(layer6_outputs(1485));
    layer7_outputs(4177) <= layer6_outputs(2585);
    layer7_outputs(4178) <= not((layer6_outputs(2941)) xor (layer6_outputs(4806)));
    layer7_outputs(4179) <= not(layer6_outputs(3283));
    layer7_outputs(4180) <= not(layer6_outputs(3434)) or (layer6_outputs(1468));
    layer7_outputs(4181) <= layer6_outputs(3618);
    layer7_outputs(4182) <= (layer6_outputs(2709)) and not (layer6_outputs(3715));
    layer7_outputs(4183) <= not((layer6_outputs(2148)) xor (layer6_outputs(4273)));
    layer7_outputs(4184) <= not((layer6_outputs(1183)) xor (layer6_outputs(3416)));
    layer7_outputs(4185) <= not(layer6_outputs(2588));
    layer7_outputs(4186) <= (layer6_outputs(3578)) or (layer6_outputs(1970));
    layer7_outputs(4187) <= not(layer6_outputs(3791)) or (layer6_outputs(1390));
    layer7_outputs(4188) <= '1';
    layer7_outputs(4189) <= (layer6_outputs(575)) xor (layer6_outputs(1086));
    layer7_outputs(4190) <= (layer6_outputs(4106)) and not (layer6_outputs(859));
    layer7_outputs(4191) <= '0';
    layer7_outputs(4192) <= not((layer6_outputs(1552)) xor (layer6_outputs(1408)));
    layer7_outputs(4193) <= not((layer6_outputs(925)) or (layer6_outputs(225)));
    layer7_outputs(4194) <= not(layer6_outputs(102));
    layer7_outputs(4195) <= layer6_outputs(2980);
    layer7_outputs(4196) <= layer6_outputs(2929);
    layer7_outputs(4197) <= layer6_outputs(3691);
    layer7_outputs(4198) <= (layer6_outputs(3400)) or (layer6_outputs(3304));
    layer7_outputs(4199) <= not((layer6_outputs(880)) xor (layer6_outputs(3036)));
    layer7_outputs(4200) <= layer6_outputs(4800);
    layer7_outputs(4201) <= layer6_outputs(1345);
    layer7_outputs(4202) <= not(layer6_outputs(2912));
    layer7_outputs(4203) <= not((layer6_outputs(2607)) or (layer6_outputs(4137)));
    layer7_outputs(4204) <= layer6_outputs(3518);
    layer7_outputs(4205) <= not((layer6_outputs(2547)) and (layer6_outputs(3297)));
    layer7_outputs(4206) <= (layer6_outputs(1204)) or (layer6_outputs(4617));
    layer7_outputs(4207) <= not(layer6_outputs(2494)) or (layer6_outputs(3396));
    layer7_outputs(4208) <= not((layer6_outputs(3987)) or (layer6_outputs(1960)));
    layer7_outputs(4209) <= not(layer6_outputs(5007));
    layer7_outputs(4210) <= not(layer6_outputs(340)) or (layer6_outputs(3670));
    layer7_outputs(4211) <= not(layer6_outputs(4883));
    layer7_outputs(4212) <= not(layer6_outputs(927));
    layer7_outputs(4213) <= not(layer6_outputs(600));
    layer7_outputs(4214) <= (layer6_outputs(1089)) and not (layer6_outputs(837));
    layer7_outputs(4215) <= (layer6_outputs(2796)) and not (layer6_outputs(2918));
    layer7_outputs(4216) <= layer6_outputs(1566);
    layer7_outputs(4217) <= layer6_outputs(3067);
    layer7_outputs(4218) <= not(layer6_outputs(4244)) or (layer6_outputs(3306));
    layer7_outputs(4219) <= layer6_outputs(1241);
    layer7_outputs(4220) <= not(layer6_outputs(4462)) or (layer6_outputs(3986));
    layer7_outputs(4221) <= (layer6_outputs(4373)) xor (layer6_outputs(1134));
    layer7_outputs(4222) <= (layer6_outputs(4204)) and (layer6_outputs(3726));
    layer7_outputs(4223) <= layer6_outputs(1698);
    layer7_outputs(4224) <= not(layer6_outputs(3665));
    layer7_outputs(4225) <= layer6_outputs(2941);
    layer7_outputs(4226) <= not(layer6_outputs(4789));
    layer7_outputs(4227) <= not(layer6_outputs(3894));
    layer7_outputs(4228) <= (layer6_outputs(4601)) and not (layer6_outputs(5037));
    layer7_outputs(4229) <= not(layer6_outputs(4300));
    layer7_outputs(4230) <= (layer6_outputs(4296)) xor (layer6_outputs(4843));
    layer7_outputs(4231) <= layer6_outputs(2725);
    layer7_outputs(4232) <= not((layer6_outputs(2672)) and (layer6_outputs(340)));
    layer7_outputs(4233) <= not(layer6_outputs(2078));
    layer7_outputs(4234) <= (layer6_outputs(2999)) and (layer6_outputs(210));
    layer7_outputs(4235) <= not(layer6_outputs(5045)) or (layer6_outputs(2784));
    layer7_outputs(4236) <= (layer6_outputs(3038)) and not (layer6_outputs(987));
    layer7_outputs(4237) <= (layer6_outputs(4239)) and (layer6_outputs(3079));
    layer7_outputs(4238) <= not((layer6_outputs(526)) or (layer6_outputs(519)));
    layer7_outputs(4239) <= layer6_outputs(3500);
    layer7_outputs(4240) <= (layer6_outputs(3642)) and not (layer6_outputs(2822));
    layer7_outputs(4241) <= not((layer6_outputs(3599)) xor (layer6_outputs(946)));
    layer7_outputs(4242) <= (layer6_outputs(3598)) and not (layer6_outputs(3057));
    layer7_outputs(4243) <= layer6_outputs(813);
    layer7_outputs(4244) <= layer6_outputs(1658);
    layer7_outputs(4245) <= layer6_outputs(2166);
    layer7_outputs(4246) <= (layer6_outputs(1848)) xor (layer6_outputs(817));
    layer7_outputs(4247) <= not(layer6_outputs(4772));
    layer7_outputs(4248) <= not(layer6_outputs(3826));
    layer7_outputs(4249) <= layer6_outputs(2444);
    layer7_outputs(4250) <= not((layer6_outputs(4268)) xor (layer6_outputs(3196)));
    layer7_outputs(4251) <= (layer6_outputs(4242)) and (layer6_outputs(1107));
    layer7_outputs(4252) <= (layer6_outputs(4460)) and not (layer6_outputs(2843));
    layer7_outputs(4253) <= layer6_outputs(1324);
    layer7_outputs(4254) <= layer6_outputs(2057);
    layer7_outputs(4255) <= (layer6_outputs(502)) and not (layer6_outputs(5044));
    layer7_outputs(4256) <= layer6_outputs(2242);
    layer7_outputs(4257) <= layer6_outputs(1849);
    layer7_outputs(4258) <= layer6_outputs(4030);
    layer7_outputs(4259) <= not((layer6_outputs(3784)) or (layer6_outputs(1518)));
    layer7_outputs(4260) <= layer6_outputs(1124);
    layer7_outputs(4261) <= not(layer6_outputs(3476));
    layer7_outputs(4262) <= layer6_outputs(4829);
    layer7_outputs(4263) <= not((layer6_outputs(2973)) and (layer6_outputs(5022)));
    layer7_outputs(4264) <= not(layer6_outputs(899));
    layer7_outputs(4265) <= (layer6_outputs(382)) and not (layer6_outputs(1156));
    layer7_outputs(4266) <= not(layer6_outputs(1459));
    layer7_outputs(4267) <= not((layer6_outputs(2091)) xor (layer6_outputs(4212)));
    layer7_outputs(4268) <= (layer6_outputs(3187)) xor (layer6_outputs(1159));
    layer7_outputs(4269) <= layer6_outputs(3218);
    layer7_outputs(4270) <= not(layer6_outputs(4945));
    layer7_outputs(4271) <= layer6_outputs(3322);
    layer7_outputs(4272) <= layer6_outputs(1447);
    layer7_outputs(4273) <= '0';
    layer7_outputs(4274) <= (layer6_outputs(5066)) or (layer6_outputs(4065));
    layer7_outputs(4275) <= layer6_outputs(3031);
    layer7_outputs(4276) <= layer6_outputs(3846);
    layer7_outputs(4277) <= not(layer6_outputs(3511));
    layer7_outputs(4278) <= not(layer6_outputs(4943));
    layer7_outputs(4279) <= (layer6_outputs(4178)) and not (layer6_outputs(4289));
    layer7_outputs(4280) <= not(layer6_outputs(87));
    layer7_outputs(4281) <= not((layer6_outputs(3065)) xor (layer6_outputs(1477)));
    layer7_outputs(4282) <= '1';
    layer7_outputs(4283) <= not((layer6_outputs(3066)) and (layer6_outputs(1601)));
    layer7_outputs(4284) <= layer6_outputs(390);
    layer7_outputs(4285) <= (layer6_outputs(1336)) or (layer6_outputs(1140));
    layer7_outputs(4286) <= (layer6_outputs(1819)) and not (layer6_outputs(3393));
    layer7_outputs(4287) <= (layer6_outputs(1729)) xor (layer6_outputs(2668));
    layer7_outputs(4288) <= not((layer6_outputs(103)) and (layer6_outputs(4427)));
    layer7_outputs(4289) <= layer6_outputs(2059);
    layer7_outputs(4290) <= layer6_outputs(3678);
    layer7_outputs(4291) <= (layer6_outputs(4767)) and not (layer6_outputs(839));
    layer7_outputs(4292) <= (layer6_outputs(3392)) xor (layer6_outputs(2512));
    layer7_outputs(4293) <= layer6_outputs(400);
    layer7_outputs(4294) <= not((layer6_outputs(3626)) xor (layer6_outputs(688)));
    layer7_outputs(4295) <= (layer6_outputs(1226)) or (layer6_outputs(2307));
    layer7_outputs(4296) <= layer6_outputs(2560);
    layer7_outputs(4297) <= not(layer6_outputs(4699)) or (layer6_outputs(2867));
    layer7_outputs(4298) <= not(layer6_outputs(3775));
    layer7_outputs(4299) <= (layer6_outputs(2630)) xor (layer6_outputs(441));
    layer7_outputs(4300) <= (layer6_outputs(3776)) and (layer6_outputs(1656));
    layer7_outputs(4301) <= (layer6_outputs(4563)) and (layer6_outputs(4004));
    layer7_outputs(4302) <= layer6_outputs(1543);
    layer7_outputs(4303) <= not(layer6_outputs(5053)) or (layer6_outputs(4453));
    layer7_outputs(4304) <= not((layer6_outputs(4815)) xor (layer6_outputs(1915)));
    layer7_outputs(4305) <= not(layer6_outputs(1654));
    layer7_outputs(4306) <= not(layer6_outputs(232)) or (layer6_outputs(2138));
    layer7_outputs(4307) <= not(layer6_outputs(2583));
    layer7_outputs(4308) <= (layer6_outputs(1002)) xor (layer6_outputs(4082));
    layer7_outputs(4309) <= layer6_outputs(4509);
    layer7_outputs(4310) <= not(layer6_outputs(57));
    layer7_outputs(4311) <= not(layer6_outputs(2271));
    layer7_outputs(4312) <= not(layer6_outputs(811)) or (layer6_outputs(448));
    layer7_outputs(4313) <= layer6_outputs(1131);
    layer7_outputs(4314) <= not(layer6_outputs(4596));
    layer7_outputs(4315) <= (layer6_outputs(2760)) xor (layer6_outputs(875));
    layer7_outputs(4316) <= not(layer6_outputs(1983));
    layer7_outputs(4317) <= not(layer6_outputs(3933));
    layer7_outputs(4318) <= not(layer6_outputs(4866));
    layer7_outputs(4319) <= layer6_outputs(2848);
    layer7_outputs(4320) <= layer6_outputs(4481);
    layer7_outputs(4321) <= (layer6_outputs(4813)) and (layer6_outputs(2524));
    layer7_outputs(4322) <= layer6_outputs(988);
    layer7_outputs(4323) <= (layer6_outputs(4693)) xor (layer6_outputs(3891));
    layer7_outputs(4324) <= layer6_outputs(35);
    layer7_outputs(4325) <= layer6_outputs(4723);
    layer7_outputs(4326) <= not((layer6_outputs(2985)) xor (layer6_outputs(3405)));
    layer7_outputs(4327) <= not(layer6_outputs(2793));
    layer7_outputs(4328) <= not(layer6_outputs(1269));
    layer7_outputs(4329) <= (layer6_outputs(3734)) or (layer6_outputs(3992));
    layer7_outputs(4330) <= not(layer6_outputs(2296));
    layer7_outputs(4331) <= not(layer6_outputs(2426));
    layer7_outputs(4332) <= (layer6_outputs(4347)) xor (layer6_outputs(970));
    layer7_outputs(4333) <= layer6_outputs(1900);
    layer7_outputs(4334) <= not(layer6_outputs(651));
    layer7_outputs(4335) <= (layer6_outputs(4879)) and not (layer6_outputs(705));
    layer7_outputs(4336) <= (layer6_outputs(1160)) xor (layer6_outputs(3989));
    layer7_outputs(4337) <= layer6_outputs(4684);
    layer7_outputs(4338) <= not(layer6_outputs(3031)) or (layer6_outputs(2389));
    layer7_outputs(4339) <= (layer6_outputs(3480)) and (layer6_outputs(53));
    layer7_outputs(4340) <= (layer6_outputs(4327)) or (layer6_outputs(4009));
    layer7_outputs(4341) <= not(layer6_outputs(2401)) or (layer6_outputs(88));
    layer7_outputs(4342) <= not(layer6_outputs(1270));
    layer7_outputs(4343) <= not(layer6_outputs(3898));
    layer7_outputs(4344) <= (layer6_outputs(4660)) xor (layer6_outputs(1787));
    layer7_outputs(4345) <= layer6_outputs(5043);
    layer7_outputs(4346) <= (layer6_outputs(3494)) or (layer6_outputs(4237));
    layer7_outputs(4347) <= not((layer6_outputs(2069)) xor (layer6_outputs(4970)));
    layer7_outputs(4348) <= (layer6_outputs(1699)) xor (layer6_outputs(2972));
    layer7_outputs(4349) <= not((layer6_outputs(2100)) xor (layer6_outputs(309)));
    layer7_outputs(4350) <= not((layer6_outputs(2819)) and (layer6_outputs(4598)));
    layer7_outputs(4351) <= layer6_outputs(3275);
    layer7_outputs(4352) <= not((layer6_outputs(2202)) xor (layer6_outputs(1276)));
    layer7_outputs(4353) <= not((layer6_outputs(1133)) xor (layer6_outputs(214)));
    layer7_outputs(4354) <= not(layer6_outputs(3476));
    layer7_outputs(4355) <= not(layer6_outputs(3808));
    layer7_outputs(4356) <= layer6_outputs(1193);
    layer7_outputs(4357) <= layer6_outputs(2892);
    layer7_outputs(4358) <= layer6_outputs(3508);
    layer7_outputs(4359) <= not(layer6_outputs(4903)) or (layer6_outputs(3458));
    layer7_outputs(4360) <= not((layer6_outputs(128)) xor (layer6_outputs(59)));
    layer7_outputs(4361) <= not(layer6_outputs(3847)) or (layer6_outputs(4218));
    layer7_outputs(4362) <= (layer6_outputs(3291)) or (layer6_outputs(4973));
    layer7_outputs(4363) <= not(layer6_outputs(2515));
    layer7_outputs(4364) <= not(layer6_outputs(4477)) or (layer6_outputs(1627));
    layer7_outputs(4365) <= '0';
    layer7_outputs(4366) <= not(layer6_outputs(220));
    layer7_outputs(4367) <= '0';
    layer7_outputs(4368) <= '0';
    layer7_outputs(4369) <= not(layer6_outputs(50));
    layer7_outputs(4370) <= (layer6_outputs(741)) xor (layer6_outputs(3817));
    layer7_outputs(4371) <= not(layer6_outputs(2722));
    layer7_outputs(4372) <= not(layer6_outputs(1853));
    layer7_outputs(4373) <= not((layer6_outputs(405)) xor (layer6_outputs(942)));
    layer7_outputs(4374) <= not(layer6_outputs(2251));
    layer7_outputs(4375) <= layer6_outputs(322);
    layer7_outputs(4376) <= not(layer6_outputs(1042));
    layer7_outputs(4377) <= not(layer6_outputs(434));
    layer7_outputs(4378) <= layer6_outputs(83);
    layer7_outputs(4379) <= not(layer6_outputs(4623));
    layer7_outputs(4380) <= (layer6_outputs(2040)) or (layer6_outputs(248));
    layer7_outputs(4381) <= not(layer6_outputs(2851)) or (layer6_outputs(3800));
    layer7_outputs(4382) <= not(layer6_outputs(1288));
    layer7_outputs(4383) <= layer6_outputs(525);
    layer7_outputs(4384) <= (layer6_outputs(1728)) and not (layer6_outputs(1421));
    layer7_outputs(4385) <= not(layer6_outputs(2036));
    layer7_outputs(4386) <= layer6_outputs(4635);
    layer7_outputs(4387) <= layer6_outputs(1841);
    layer7_outputs(4388) <= '0';
    layer7_outputs(4389) <= not(layer6_outputs(4990));
    layer7_outputs(4390) <= not(layer6_outputs(2051));
    layer7_outputs(4391) <= (layer6_outputs(1542)) and not (layer6_outputs(4435));
    layer7_outputs(4392) <= (layer6_outputs(3845)) and (layer6_outputs(3985));
    layer7_outputs(4393) <= not(layer6_outputs(1858));
    layer7_outputs(4394) <= not((layer6_outputs(1450)) xor (layer6_outputs(1805)));
    layer7_outputs(4395) <= not(layer6_outputs(147));
    layer7_outputs(4396) <= (layer6_outputs(4016)) xor (layer6_outputs(1617));
    layer7_outputs(4397) <= (layer6_outputs(3807)) xor (layer6_outputs(4920));
    layer7_outputs(4398) <= (layer6_outputs(4148)) and not (layer6_outputs(444));
    layer7_outputs(4399) <= (layer6_outputs(4706)) and (layer6_outputs(3287));
    layer7_outputs(4400) <= not(layer6_outputs(3764));
    layer7_outputs(4401) <= (layer6_outputs(1020)) or (layer6_outputs(3020));
    layer7_outputs(4402) <= (layer6_outputs(682)) and not (layer6_outputs(1017));
    layer7_outputs(4403) <= not((layer6_outputs(2769)) and (layer6_outputs(20)));
    layer7_outputs(4404) <= layer6_outputs(2464);
    layer7_outputs(4405) <= not(layer6_outputs(3326));
    layer7_outputs(4406) <= (layer6_outputs(2555)) and not (layer6_outputs(4063));
    layer7_outputs(4407) <= not(layer6_outputs(290));
    layer7_outputs(4408) <= layer6_outputs(516);
    layer7_outputs(4409) <= (layer6_outputs(3448)) and (layer6_outputs(798));
    layer7_outputs(4410) <= not(layer6_outputs(4546));
    layer7_outputs(4411) <= '0';
    layer7_outputs(4412) <= not(layer6_outputs(1562));
    layer7_outputs(4413) <= (layer6_outputs(5025)) and (layer6_outputs(1227));
    layer7_outputs(4414) <= not(layer6_outputs(4385)) or (layer6_outputs(2142));
    layer7_outputs(4415) <= (layer6_outputs(1874)) and not (layer6_outputs(463));
    layer7_outputs(4416) <= not(layer6_outputs(962));
    layer7_outputs(4417) <= not(layer6_outputs(2781));
    layer7_outputs(4418) <= not(layer6_outputs(4779)) or (layer6_outputs(4073));
    layer7_outputs(4419) <= layer6_outputs(363);
    layer7_outputs(4420) <= (layer6_outputs(3602)) and not (layer6_outputs(1487));
    layer7_outputs(4421) <= layer6_outputs(94);
    layer7_outputs(4422) <= (layer6_outputs(4525)) xor (layer6_outputs(1927));
    layer7_outputs(4423) <= (layer6_outputs(1271)) and not (layer6_outputs(3544));
    layer7_outputs(4424) <= (layer6_outputs(629)) or (layer6_outputs(3147));
    layer7_outputs(4425) <= not((layer6_outputs(4936)) xor (layer6_outputs(4773)));
    layer7_outputs(4426) <= not((layer6_outputs(2799)) xor (layer6_outputs(1529)));
    layer7_outputs(4427) <= not(layer6_outputs(1249));
    layer7_outputs(4428) <= not(layer6_outputs(3242)) or (layer6_outputs(3896));
    layer7_outputs(4429) <= layer6_outputs(3980);
    layer7_outputs(4430) <= not((layer6_outputs(1742)) and (layer6_outputs(356)));
    layer7_outputs(4431) <= (layer6_outputs(3369)) and (layer6_outputs(3662));
    layer7_outputs(4432) <= not(layer6_outputs(322)) or (layer6_outputs(1682));
    layer7_outputs(4433) <= not(layer6_outputs(710));
    layer7_outputs(4434) <= layer6_outputs(4719);
    layer7_outputs(4435) <= (layer6_outputs(4681)) xor (layer6_outputs(1410));
    layer7_outputs(4436) <= (layer6_outputs(4290)) xor (layer6_outputs(1506));
    layer7_outputs(4437) <= layer6_outputs(3056);
    layer7_outputs(4438) <= not((layer6_outputs(3850)) xor (layer6_outputs(2341)));
    layer7_outputs(4439) <= (layer6_outputs(3987)) or (layer6_outputs(2841));
    layer7_outputs(4440) <= not(layer6_outputs(3012)) or (layer6_outputs(1165));
    layer7_outputs(4441) <= not(layer6_outputs(2687));
    layer7_outputs(4442) <= not(layer6_outputs(304));
    layer7_outputs(4443) <= (layer6_outputs(4690)) xor (layer6_outputs(871));
    layer7_outputs(4444) <= '0';
    layer7_outputs(4445) <= layer6_outputs(1806);
    layer7_outputs(4446) <= not((layer6_outputs(3255)) xor (layer6_outputs(3137)));
    layer7_outputs(4447) <= not((layer6_outputs(1676)) or (layer6_outputs(2882)));
    layer7_outputs(4448) <= not(layer6_outputs(1745));
    layer7_outputs(4449) <= not(layer6_outputs(3062));
    layer7_outputs(4450) <= layer6_outputs(4209);
    layer7_outputs(4451) <= not(layer6_outputs(1988)) or (layer6_outputs(2844));
    layer7_outputs(4452) <= not(layer6_outputs(1011)) or (layer6_outputs(4308));
    layer7_outputs(4453) <= not(layer6_outputs(928));
    layer7_outputs(4454) <= not(layer6_outputs(3923));
    layer7_outputs(4455) <= (layer6_outputs(58)) xor (layer6_outputs(1628));
    layer7_outputs(4456) <= not(layer6_outputs(1335));
    layer7_outputs(4457) <= not(layer6_outputs(4066));
    layer7_outputs(4458) <= not(layer6_outputs(1075)) or (layer6_outputs(625));
    layer7_outputs(4459) <= not(layer6_outputs(715));
    layer7_outputs(4460) <= (layer6_outputs(1214)) xor (layer6_outputs(743));
    layer7_outputs(4461) <= not(layer6_outputs(892));
    layer7_outputs(4462) <= not((layer6_outputs(1633)) or (layer6_outputs(2003)));
    layer7_outputs(4463) <= (layer6_outputs(1589)) or (layer6_outputs(4424));
    layer7_outputs(4464) <= not(layer6_outputs(611));
    layer7_outputs(4465) <= not((layer6_outputs(2233)) and (layer6_outputs(3330)));
    layer7_outputs(4466) <= layer6_outputs(423);
    layer7_outputs(4467) <= (layer6_outputs(647)) or (layer6_outputs(488));
    layer7_outputs(4468) <= '1';
    layer7_outputs(4469) <= not((layer6_outputs(1766)) xor (layer6_outputs(459)));
    layer7_outputs(4470) <= not(layer6_outputs(3984)) or (layer6_outputs(334));
    layer7_outputs(4471) <= not(layer6_outputs(1228));
    layer7_outputs(4472) <= not((layer6_outputs(453)) and (layer6_outputs(2952)));
    layer7_outputs(4473) <= (layer6_outputs(4957)) xor (layer6_outputs(1637));
    layer7_outputs(4474) <= layer6_outputs(3119);
    layer7_outputs(4475) <= not(layer6_outputs(2306));
    layer7_outputs(4476) <= not(layer6_outputs(4580));
    layer7_outputs(4477) <= (layer6_outputs(1101)) or (layer6_outputs(2173));
    layer7_outputs(4478) <= not(layer6_outputs(3895));
    layer7_outputs(4479) <= not(layer6_outputs(3959));
    layer7_outputs(4480) <= not(layer6_outputs(288));
    layer7_outputs(4481) <= not(layer6_outputs(4887)) or (layer6_outputs(1678));
    layer7_outputs(4482) <= not(layer6_outputs(5012));
    layer7_outputs(4483) <= not(layer6_outputs(874));
    layer7_outputs(4484) <= (layer6_outputs(3250)) xor (layer6_outputs(749));
    layer7_outputs(4485) <= (layer6_outputs(4220)) and (layer6_outputs(2688));
    layer7_outputs(4486) <= layer6_outputs(3150);
    layer7_outputs(4487) <= not(layer6_outputs(2391)) or (layer6_outputs(3135));
    layer7_outputs(4488) <= (layer6_outputs(3857)) or (layer6_outputs(1384));
    layer7_outputs(4489) <= layer6_outputs(4633);
    layer7_outputs(4490) <= layer6_outputs(3899);
    layer7_outputs(4491) <= not(layer6_outputs(2729));
    layer7_outputs(4492) <= not(layer6_outputs(4071));
    layer7_outputs(4493) <= layer6_outputs(1292);
    layer7_outputs(4494) <= not((layer6_outputs(4092)) xor (layer6_outputs(255)));
    layer7_outputs(4495) <= not((layer6_outputs(384)) and (layer6_outputs(4273)));
    layer7_outputs(4496) <= not(layer6_outputs(3024));
    layer7_outputs(4497) <= '0';
    layer7_outputs(4498) <= not(layer6_outputs(3050));
    layer7_outputs(4499) <= layer6_outputs(3491);
    layer7_outputs(4500) <= (layer6_outputs(589)) and not (layer6_outputs(2754));
    layer7_outputs(4501) <= (layer6_outputs(263)) xor (layer6_outputs(1019));
    layer7_outputs(4502) <= not(layer6_outputs(3253));
    layer7_outputs(4503) <= layer6_outputs(3346);
    layer7_outputs(4504) <= (layer6_outputs(2935)) or (layer6_outputs(3709));
    layer7_outputs(4505) <= not(layer6_outputs(3381)) or (layer6_outputs(1951));
    layer7_outputs(4506) <= (layer6_outputs(4923)) and not (layer6_outputs(5102));
    layer7_outputs(4507) <= '0';
    layer7_outputs(4508) <= layer6_outputs(581);
    layer7_outputs(4509) <= layer6_outputs(4956);
    layer7_outputs(4510) <= not((layer6_outputs(2179)) xor (layer6_outputs(3802)));
    layer7_outputs(4511) <= layer6_outputs(2464);
    layer7_outputs(4512) <= (layer6_outputs(455)) or (layer6_outputs(2943));
    layer7_outputs(4513) <= not((layer6_outputs(1326)) xor (layer6_outputs(2953)));
    layer7_outputs(4514) <= not(layer6_outputs(4576)) or (layer6_outputs(2116));
    layer7_outputs(4515) <= layer6_outputs(3288);
    layer7_outputs(4516) <= layer6_outputs(4421);
    layer7_outputs(4517) <= layer6_outputs(3875);
    layer7_outputs(4518) <= layer6_outputs(4977);
    layer7_outputs(4519) <= not(layer6_outputs(2791));
    layer7_outputs(4520) <= not(layer6_outputs(4142));
    layer7_outputs(4521) <= not((layer6_outputs(1534)) or (layer6_outputs(3018)));
    layer7_outputs(4522) <= layer6_outputs(2015);
    layer7_outputs(4523) <= not(layer6_outputs(546));
    layer7_outputs(4524) <= not((layer6_outputs(1937)) or (layer6_outputs(2598)));
    layer7_outputs(4525) <= not(layer6_outputs(802));
    layer7_outputs(4526) <= layer6_outputs(2783);
    layer7_outputs(4527) <= not(layer6_outputs(4935));
    layer7_outputs(4528) <= layer6_outputs(947);
    layer7_outputs(4529) <= layer6_outputs(3715);
    layer7_outputs(4530) <= not(layer6_outputs(2127)) or (layer6_outputs(2308));
    layer7_outputs(4531) <= not((layer6_outputs(4098)) xor (layer6_outputs(1327)));
    layer7_outputs(4532) <= layer6_outputs(2736);
    layer7_outputs(4533) <= layer6_outputs(1852);
    layer7_outputs(4534) <= '1';
    layer7_outputs(4535) <= not(layer6_outputs(3230));
    layer7_outputs(4536) <= not(layer6_outputs(4550));
    layer7_outputs(4537) <= (layer6_outputs(4046)) xor (layer6_outputs(402));
    layer7_outputs(4538) <= not((layer6_outputs(1480)) xor (layer6_outputs(1463)));
    layer7_outputs(4539) <= not((layer6_outputs(263)) xor (layer6_outputs(1578)));
    layer7_outputs(4540) <= not(layer6_outputs(4380));
    layer7_outputs(4541) <= not(layer6_outputs(1067));
    layer7_outputs(4542) <= (layer6_outputs(4310)) or (layer6_outputs(4118));
    layer7_outputs(4543) <= not(layer6_outputs(2910));
    layer7_outputs(4544) <= not((layer6_outputs(4349)) xor (layer6_outputs(1416)));
    layer7_outputs(4545) <= not(layer6_outputs(540));
    layer7_outputs(4546) <= not(layer6_outputs(4817));
    layer7_outputs(4547) <= layer6_outputs(5063);
    layer7_outputs(4548) <= (layer6_outputs(4319)) or (layer6_outputs(1078));
    layer7_outputs(4549) <= (layer6_outputs(1877)) and not (layer6_outputs(1248));
    layer7_outputs(4550) <= layer6_outputs(1088);
    layer7_outputs(4551) <= layer6_outputs(179);
    layer7_outputs(4552) <= not(layer6_outputs(4985));
    layer7_outputs(4553) <= not((layer6_outputs(609)) or (layer6_outputs(2426)));
    layer7_outputs(4554) <= not(layer6_outputs(1558));
    layer7_outputs(4555) <= (layer6_outputs(579)) xor (layer6_outputs(4912));
    layer7_outputs(4556) <= layer6_outputs(873);
    layer7_outputs(4557) <= not((layer6_outputs(4416)) xor (layer6_outputs(163)));
    layer7_outputs(4558) <= not((layer6_outputs(2380)) and (layer6_outputs(222)));
    layer7_outputs(4559) <= layer6_outputs(4191);
    layer7_outputs(4560) <= not(layer6_outputs(4301));
    layer7_outputs(4561) <= (layer6_outputs(3903)) xor (layer6_outputs(2052));
    layer7_outputs(4562) <= (layer6_outputs(535)) and not (layer6_outputs(5106));
    layer7_outputs(4563) <= not(layer6_outputs(2079)) or (layer6_outputs(2161));
    layer7_outputs(4564) <= (layer6_outputs(1720)) or (layer6_outputs(2937));
    layer7_outputs(4565) <= not((layer6_outputs(386)) xor (layer6_outputs(2417)));
    layer7_outputs(4566) <= not(layer6_outputs(451)) or (layer6_outputs(4115));
    layer7_outputs(4567) <= not(layer6_outputs(2290));
    layer7_outputs(4568) <= not((layer6_outputs(93)) xor (layer6_outputs(5021)));
    layer7_outputs(4569) <= not((layer6_outputs(3411)) and (layer6_outputs(4230)));
    layer7_outputs(4570) <= layer6_outputs(4369);
    layer7_outputs(4571) <= not((layer6_outputs(1245)) xor (layer6_outputs(3482)));
    layer7_outputs(4572) <= not(layer6_outputs(1572)) or (layer6_outputs(4892));
    layer7_outputs(4573) <= layer6_outputs(918);
    layer7_outputs(4574) <= layer6_outputs(574);
    layer7_outputs(4575) <= not((layer6_outputs(1936)) xor (layer6_outputs(1525)));
    layer7_outputs(4576) <= layer6_outputs(2000);
    layer7_outputs(4577) <= (layer6_outputs(2748)) and not (layer6_outputs(1549));
    layer7_outputs(4578) <= not(layer6_outputs(3575));
    layer7_outputs(4579) <= layer6_outputs(4314);
    layer7_outputs(4580) <= not(layer6_outputs(1543));
    layer7_outputs(4581) <= (layer6_outputs(1497)) xor (layer6_outputs(1744));
    layer7_outputs(4582) <= not(layer6_outputs(274));
    layer7_outputs(4583) <= layer6_outputs(186);
    layer7_outputs(4584) <= layer6_outputs(3490);
    layer7_outputs(4585) <= (layer6_outputs(852)) and not (layer6_outputs(4665));
    layer7_outputs(4586) <= layer6_outputs(442);
    layer7_outputs(4587) <= layer6_outputs(4186);
    layer7_outputs(4588) <= not(layer6_outputs(2861));
    layer7_outputs(4589) <= not(layer6_outputs(1405)) or (layer6_outputs(1722));
    layer7_outputs(4590) <= (layer6_outputs(2696)) and (layer6_outputs(1389));
    layer7_outputs(4591) <= (layer6_outputs(116)) and (layer6_outputs(1746));
    layer7_outputs(4592) <= not(layer6_outputs(292));
    layer7_outputs(4593) <= not(layer6_outputs(4320)) or (layer6_outputs(806));
    layer7_outputs(4594) <= (layer6_outputs(2431)) xor (layer6_outputs(2561));
    layer7_outputs(4595) <= not((layer6_outputs(1452)) xor (layer6_outputs(729)));
    layer7_outputs(4596) <= not(layer6_outputs(161));
    layer7_outputs(4597) <= layer6_outputs(2625);
    layer7_outputs(4598) <= not(layer6_outputs(8));
    layer7_outputs(4599) <= not(layer6_outputs(2703));
    layer7_outputs(4600) <= layer6_outputs(4807);
    layer7_outputs(4601) <= not((layer6_outputs(3117)) xor (layer6_outputs(1198)));
    layer7_outputs(4602) <= (layer6_outputs(2750)) xor (layer6_outputs(3048));
    layer7_outputs(4603) <= '1';
    layer7_outputs(4604) <= layer6_outputs(5089);
    layer7_outputs(4605) <= not(layer6_outputs(5115)) or (layer6_outputs(2179));
    layer7_outputs(4606) <= not(layer6_outputs(1827));
    layer7_outputs(4607) <= (layer6_outputs(1951)) and (layer6_outputs(4931));
    layer7_outputs(4608) <= not(layer6_outputs(2921));
    layer7_outputs(4609) <= layer6_outputs(4751);
    layer7_outputs(4610) <= layer6_outputs(2117);
    layer7_outputs(4611) <= (layer6_outputs(1005)) and (layer6_outputs(3579));
    layer7_outputs(4612) <= not(layer6_outputs(60));
    layer7_outputs(4613) <= layer6_outputs(1712);
    layer7_outputs(4614) <= layer6_outputs(1521);
    layer7_outputs(4615) <= not(layer6_outputs(4311));
    layer7_outputs(4616) <= not(layer6_outputs(638));
    layer7_outputs(4617) <= not((layer6_outputs(1755)) or (layer6_outputs(1813)));
    layer7_outputs(4618) <= not(layer6_outputs(641));
    layer7_outputs(4619) <= not(layer6_outputs(611));
    layer7_outputs(4620) <= layer6_outputs(298);
    layer7_outputs(4621) <= layer6_outputs(2904);
    layer7_outputs(4622) <= not(layer6_outputs(3646));
    layer7_outputs(4623) <= layer6_outputs(4127);
    layer7_outputs(4624) <= (layer6_outputs(1010)) or (layer6_outputs(3698));
    layer7_outputs(4625) <= (layer6_outputs(2535)) and (layer6_outputs(2707));
    layer7_outputs(4626) <= layer6_outputs(2691);
    layer7_outputs(4627) <= not(layer6_outputs(4438)) or (layer6_outputs(2744));
    layer7_outputs(4628) <= not((layer6_outputs(3481)) or (layer6_outputs(2413)));
    layer7_outputs(4629) <= layer6_outputs(613);
    layer7_outputs(4630) <= not((layer6_outputs(2479)) xor (layer6_outputs(1846)));
    layer7_outputs(4631) <= layer6_outputs(475);
    layer7_outputs(4632) <= layer6_outputs(3058);
    layer7_outputs(4633) <= (layer6_outputs(3223)) xor (layer6_outputs(2341));
    layer7_outputs(4634) <= layer6_outputs(3207);
    layer7_outputs(4635) <= not(layer6_outputs(3658)) or (layer6_outputs(3991));
    layer7_outputs(4636) <= layer6_outputs(752);
    layer7_outputs(4637) <= not((layer6_outputs(4941)) xor (layer6_outputs(2691)));
    layer7_outputs(4638) <= (layer6_outputs(916)) and not (layer6_outputs(1168));
    layer7_outputs(4639) <= layer6_outputs(1274);
    layer7_outputs(4640) <= layer6_outputs(3355);
    layer7_outputs(4641) <= not(layer6_outputs(2705)) or (layer6_outputs(2566));
    layer7_outputs(4642) <= (layer6_outputs(2206)) or (layer6_outputs(2554));
    layer7_outputs(4643) <= (layer6_outputs(3631)) and (layer6_outputs(4544));
    layer7_outputs(4644) <= layer6_outputs(1601);
    layer7_outputs(4645) <= not(layer6_outputs(2366));
    layer7_outputs(4646) <= layer6_outputs(1309);
    layer7_outputs(4647) <= (layer6_outputs(3279)) or (layer6_outputs(1433));
    layer7_outputs(4648) <= layer6_outputs(430);
    layer7_outputs(4649) <= not((layer6_outputs(1471)) xor (layer6_outputs(4504)));
    layer7_outputs(4650) <= not(layer6_outputs(5060));
    layer7_outputs(4651) <= layer6_outputs(4276);
    layer7_outputs(4652) <= layer6_outputs(4494);
    layer7_outputs(4653) <= (layer6_outputs(325)) and not (layer6_outputs(1247));
    layer7_outputs(4654) <= not(layer6_outputs(2595));
    layer7_outputs(4655) <= not(layer6_outputs(4485));
    layer7_outputs(4656) <= (layer6_outputs(2797)) or (layer6_outputs(1437));
    layer7_outputs(4657) <= (layer6_outputs(3819)) or (layer6_outputs(3692));
    layer7_outputs(4658) <= '1';
    layer7_outputs(4659) <= not((layer6_outputs(818)) xor (layer6_outputs(1580)));
    layer7_outputs(4660) <= not(layer6_outputs(4866));
    layer7_outputs(4661) <= not(layer6_outputs(2434));
    layer7_outputs(4662) <= (layer6_outputs(3700)) xor (layer6_outputs(1600));
    layer7_outputs(4663) <= (layer6_outputs(538)) and not (layer6_outputs(673));
    layer7_outputs(4664) <= layer6_outputs(285);
    layer7_outputs(4665) <= not(layer6_outputs(149)) or (layer6_outputs(1772));
    layer7_outputs(4666) <= layer6_outputs(465);
    layer7_outputs(4667) <= not(layer6_outputs(2380));
    layer7_outputs(4668) <= not((layer6_outputs(901)) and (layer6_outputs(4389)));
    layer7_outputs(4669) <= layer6_outputs(3020);
    layer7_outputs(4670) <= layer6_outputs(2990);
    layer7_outputs(4671) <= not((layer6_outputs(705)) and (layer6_outputs(4481)));
    layer7_outputs(4672) <= not((layer6_outputs(446)) or (layer6_outputs(3860)));
    layer7_outputs(4673) <= not((layer6_outputs(387)) or (layer6_outputs(2740)));
    layer7_outputs(4674) <= not(layer6_outputs(1484));
    layer7_outputs(4675) <= (layer6_outputs(2192)) or (layer6_outputs(944));
    layer7_outputs(4676) <= not(layer6_outputs(885));
    layer7_outputs(4677) <= layer6_outputs(1767);
    layer7_outputs(4678) <= (layer6_outputs(4085)) xor (layer6_outputs(5019));
    layer7_outputs(4679) <= (layer6_outputs(370)) and not (layer6_outputs(2045));
    layer7_outputs(4680) <= (layer6_outputs(849)) and (layer6_outputs(3517));
    layer7_outputs(4681) <= not((layer6_outputs(911)) and (layer6_outputs(303)));
    layer7_outputs(4682) <= (layer6_outputs(875)) and not (layer6_outputs(2737));
    layer7_outputs(4683) <= layer6_outputs(543);
    layer7_outputs(4684) <= not(layer6_outputs(15));
    layer7_outputs(4685) <= layer6_outputs(5);
    layer7_outputs(4686) <= not((layer6_outputs(3951)) or (layer6_outputs(4935)));
    layer7_outputs(4687) <= layer6_outputs(4175);
    layer7_outputs(4688) <= not(layer6_outputs(250));
    layer7_outputs(4689) <= layer6_outputs(2331);
    layer7_outputs(4690) <= not(layer6_outputs(294));
    layer7_outputs(4691) <= not(layer6_outputs(677));
    layer7_outputs(4692) <= not((layer6_outputs(2368)) or (layer6_outputs(3721)));
    layer7_outputs(4693) <= layer6_outputs(2523);
    layer7_outputs(4694) <= not(layer6_outputs(1364)) or (layer6_outputs(4627));
    layer7_outputs(4695) <= not(layer6_outputs(243)) or (layer6_outputs(4523));
    layer7_outputs(4696) <= (layer6_outputs(667)) xor (layer6_outputs(1687));
    layer7_outputs(4697) <= not((layer6_outputs(307)) and (layer6_outputs(1899)));
    layer7_outputs(4698) <= layer6_outputs(1517);
    layer7_outputs(4699) <= layer6_outputs(2456);
    layer7_outputs(4700) <= not(layer6_outputs(1624));
    layer7_outputs(4701) <= not(layer6_outputs(4547));
    layer7_outputs(4702) <= not((layer6_outputs(4637)) or (layer6_outputs(1097)));
    layer7_outputs(4703) <= not((layer6_outputs(3758)) and (layer6_outputs(1675)));
    layer7_outputs(4704) <= layer6_outputs(4218);
    layer7_outputs(4705) <= (layer6_outputs(3608)) xor (layer6_outputs(5030));
    layer7_outputs(4706) <= not(layer6_outputs(1717));
    layer7_outputs(4707) <= not(layer6_outputs(3567));
    layer7_outputs(4708) <= layer6_outputs(4174);
    layer7_outputs(4709) <= (layer6_outputs(2604)) xor (layer6_outputs(3526));
    layer7_outputs(4710) <= not((layer6_outputs(1807)) xor (layer6_outputs(2921)));
    layer7_outputs(4711) <= (layer6_outputs(1135)) or (layer6_outputs(4955));
    layer7_outputs(4712) <= not(layer6_outputs(2730));
    layer7_outputs(4713) <= (layer6_outputs(3495)) and (layer6_outputs(26));
    layer7_outputs(4714) <= not(layer6_outputs(5090));
    layer7_outputs(4715) <= (layer6_outputs(172)) or (layer6_outputs(265));
    layer7_outputs(4716) <= layer6_outputs(4147);
    layer7_outputs(4717) <= not(layer6_outputs(2171));
    layer7_outputs(4718) <= not(layer6_outputs(3297));
    layer7_outputs(4719) <= not(layer6_outputs(2532));
    layer7_outputs(4720) <= (layer6_outputs(4578)) and not (layer6_outputs(97));
    layer7_outputs(4721) <= not(layer6_outputs(1126)) or (layer6_outputs(4950));
    layer7_outputs(4722) <= layer6_outputs(3529);
    layer7_outputs(4723) <= not(layer6_outputs(2439));
    layer7_outputs(4724) <= layer6_outputs(3889);
    layer7_outputs(4725) <= not((layer6_outputs(1112)) xor (layer6_outputs(3684)));
    layer7_outputs(4726) <= not((layer6_outputs(3725)) or (layer6_outputs(4425)));
    layer7_outputs(4727) <= not(layer6_outputs(296));
    layer7_outputs(4728) <= '1';
    layer7_outputs(4729) <= (layer6_outputs(3962)) xor (layer6_outputs(3186));
    layer7_outputs(4730) <= layer6_outputs(2951);
    layer7_outputs(4731) <= layer6_outputs(4582);
    layer7_outputs(4732) <= not(layer6_outputs(2242));
    layer7_outputs(4733) <= not((layer6_outputs(2992)) or (layer6_outputs(893)));
    layer7_outputs(4734) <= layer6_outputs(695);
    layer7_outputs(4735) <= not((layer6_outputs(2971)) or (layer6_outputs(954)));
    layer7_outputs(4736) <= not((layer6_outputs(328)) xor (layer6_outputs(2939)));
    layer7_outputs(4737) <= (layer6_outputs(1496)) and not (layer6_outputs(109));
    layer7_outputs(4738) <= not((layer6_outputs(3404)) and (layer6_outputs(2697)));
    layer7_outputs(4739) <= not(layer6_outputs(3634));
    layer7_outputs(4740) <= not((layer6_outputs(450)) xor (layer6_outputs(4423)));
    layer7_outputs(4741) <= not(layer6_outputs(2428)) or (layer6_outputs(890));
    layer7_outputs(4742) <= (layer6_outputs(3274)) or (layer6_outputs(1640));
    layer7_outputs(4743) <= (layer6_outputs(3690)) and (layer6_outputs(1571));
    layer7_outputs(4744) <= (layer6_outputs(2309)) and (layer6_outputs(1191));
    layer7_outputs(4745) <= not(layer6_outputs(2041));
    layer7_outputs(4746) <= layer6_outputs(1546);
    layer7_outputs(4747) <= not(layer6_outputs(449)) or (layer6_outputs(4303));
    layer7_outputs(4748) <= layer6_outputs(4727);
    layer7_outputs(4749) <= (layer6_outputs(3932)) or (layer6_outputs(2250));
    layer7_outputs(4750) <= layer6_outputs(777);
    layer7_outputs(4751) <= layer6_outputs(661);
    layer7_outputs(4752) <= not((layer6_outputs(2763)) and (layer6_outputs(2054)));
    layer7_outputs(4753) <= '1';
    layer7_outputs(4754) <= (layer6_outputs(3821)) xor (layer6_outputs(2748));
    layer7_outputs(4755) <= not((layer6_outputs(1908)) xor (layer6_outputs(4388)));
    layer7_outputs(4756) <= layer6_outputs(1926);
    layer7_outputs(4757) <= (layer6_outputs(1011)) and not (layer6_outputs(4888));
    layer7_outputs(4758) <= not(layer6_outputs(4193));
    layer7_outputs(4759) <= not((layer6_outputs(443)) and (layer6_outputs(4612)));
    layer7_outputs(4760) <= (layer6_outputs(870)) and not (layer6_outputs(1533));
    layer7_outputs(4761) <= (layer6_outputs(2700)) and (layer6_outputs(3727));
    layer7_outputs(4762) <= (layer6_outputs(97)) or (layer6_outputs(3930));
    layer7_outputs(4763) <= '1';
    layer7_outputs(4764) <= not(layer6_outputs(1896)) or (layer6_outputs(1091));
    layer7_outputs(4765) <= (layer6_outputs(2601)) xor (layer6_outputs(3716));
    layer7_outputs(4766) <= not(layer6_outputs(4384));
    layer7_outputs(4767) <= (layer6_outputs(2822)) or (layer6_outputs(2299));
    layer7_outputs(4768) <= not(layer6_outputs(168));
    layer7_outputs(4769) <= not(layer6_outputs(0));
    layer7_outputs(4770) <= layer6_outputs(1975);
    layer7_outputs(4771) <= not(layer6_outputs(1547));
    layer7_outputs(4772) <= not((layer6_outputs(303)) xor (layer6_outputs(3067)));
    layer7_outputs(4773) <= layer6_outputs(4330);
    layer7_outputs(4774) <= layer6_outputs(2942);
    layer7_outputs(4775) <= not((layer6_outputs(2034)) or (layer6_outputs(140)));
    layer7_outputs(4776) <= (layer6_outputs(3979)) xor (layer6_outputs(2340));
    layer7_outputs(4777) <= (layer6_outputs(100)) or (layer6_outputs(3769));
    layer7_outputs(4778) <= (layer6_outputs(4823)) and not (layer6_outputs(923));
    layer7_outputs(4779) <= not(layer6_outputs(3706));
    layer7_outputs(4780) <= not((layer6_outputs(845)) xor (layer6_outputs(3)));
    layer7_outputs(4781) <= not((layer6_outputs(3291)) and (layer6_outputs(3690)));
    layer7_outputs(4782) <= layer6_outputs(3882);
    layer7_outputs(4783) <= layer6_outputs(1528);
    layer7_outputs(4784) <= layer6_outputs(1388);
    layer7_outputs(4785) <= layer6_outputs(3164);
    layer7_outputs(4786) <= not((layer6_outputs(4632)) xor (layer6_outputs(1274)));
    layer7_outputs(4787) <= not(layer6_outputs(1669)) or (layer6_outputs(4184));
    layer7_outputs(4788) <= not((layer6_outputs(642)) or (layer6_outputs(3776)));
    layer7_outputs(4789) <= not(layer6_outputs(4322));
    layer7_outputs(4790) <= not(layer6_outputs(2239));
    layer7_outputs(4791) <= not(layer6_outputs(1535)) or (layer6_outputs(4663));
    layer7_outputs(4792) <= not(layer6_outputs(2379));
    layer7_outputs(4793) <= layer6_outputs(2067);
    layer7_outputs(4794) <= layer6_outputs(4934);
    layer7_outputs(4795) <= (layer6_outputs(1780)) and not (layer6_outputs(4406));
    layer7_outputs(4796) <= not(layer6_outputs(3354));
    layer7_outputs(4797) <= not(layer6_outputs(4814));
    layer7_outputs(4798) <= not(layer6_outputs(3977)) or (layer6_outputs(2446));
    layer7_outputs(4799) <= not((layer6_outputs(2060)) and (layer6_outputs(1616)));
    layer7_outputs(4800) <= not(layer6_outputs(3531));
    layer7_outputs(4801) <= '0';
    layer7_outputs(4802) <= '1';
    layer7_outputs(4803) <= not(layer6_outputs(2785));
    layer7_outputs(4804) <= not(layer6_outputs(752)) or (layer6_outputs(4718));
    layer7_outputs(4805) <= not(layer6_outputs(18));
    layer7_outputs(4806) <= not(layer6_outputs(4476));
    layer7_outputs(4807) <= not((layer6_outputs(3399)) or (layer6_outputs(4577)));
    layer7_outputs(4808) <= (layer6_outputs(346)) and not (layer6_outputs(1260));
    layer7_outputs(4809) <= not(layer6_outputs(2037));
    layer7_outputs(4810) <= layer6_outputs(1384);
    layer7_outputs(4811) <= layer6_outputs(1990);
    layer7_outputs(4812) <= (layer6_outputs(2418)) xor (layer6_outputs(1984));
    layer7_outputs(4813) <= (layer6_outputs(2689)) xor (layer6_outputs(2317));
    layer7_outputs(4814) <= (layer6_outputs(4579)) xor (layer6_outputs(33));
    layer7_outputs(4815) <= not(layer6_outputs(1056));
    layer7_outputs(4816) <= layer6_outputs(365);
    layer7_outputs(4817) <= not(layer6_outputs(1286));
    layer7_outputs(4818) <= not((layer6_outputs(984)) or (layer6_outputs(3773)));
    layer7_outputs(4819) <= not((layer6_outputs(2639)) or (layer6_outputs(4658)));
    layer7_outputs(4820) <= (layer6_outputs(4458)) and (layer6_outputs(2626));
    layer7_outputs(4821) <= (layer6_outputs(78)) xor (layer6_outputs(5008));
    layer7_outputs(4822) <= not((layer6_outputs(410)) and (layer6_outputs(2205)));
    layer7_outputs(4823) <= layer6_outputs(2923);
    layer7_outputs(4824) <= (layer6_outputs(4475)) and not (layer6_outputs(3401));
    layer7_outputs(4825) <= (layer6_outputs(2506)) xor (layer6_outputs(3556));
    layer7_outputs(4826) <= not(layer6_outputs(2103));
    layer7_outputs(4827) <= not((layer6_outputs(3763)) or (layer6_outputs(1997)));
    layer7_outputs(4828) <= not((layer6_outputs(528)) and (layer6_outputs(613)));
    layer7_outputs(4829) <= not(layer6_outputs(3645));
    layer7_outputs(4830) <= not(layer6_outputs(3609));
    layer7_outputs(4831) <= layer6_outputs(3308);
    layer7_outputs(4832) <= not(layer6_outputs(2363)) or (layer6_outputs(1930));
    layer7_outputs(4833) <= layer6_outputs(3182);
    layer7_outputs(4834) <= not((layer6_outputs(289)) and (layer6_outputs(3290)));
    layer7_outputs(4835) <= not((layer6_outputs(1295)) xor (layer6_outputs(3253)));
    layer7_outputs(4836) <= layer6_outputs(4721);
    layer7_outputs(4837) <= not(layer6_outputs(3023)) or (layer6_outputs(1137));
    layer7_outputs(4838) <= not(layer6_outputs(3421));
    layer7_outputs(4839) <= not(layer6_outputs(4352));
    layer7_outputs(4840) <= layer6_outputs(2564);
    layer7_outputs(4841) <= not(layer6_outputs(2612));
    layer7_outputs(4842) <= not(layer6_outputs(3816));
    layer7_outputs(4843) <= not(layer6_outputs(321));
    layer7_outputs(4844) <= (layer6_outputs(4574)) xor (layer6_outputs(4535));
    layer7_outputs(4845) <= (layer6_outputs(1114)) and not (layer6_outputs(6));
    layer7_outputs(4846) <= not(layer6_outputs(3125));
    layer7_outputs(4847) <= not(layer6_outputs(2932)) or (layer6_outputs(1551));
    layer7_outputs(4848) <= not(layer6_outputs(3362)) or (layer6_outputs(2758));
    layer7_outputs(4849) <= (layer6_outputs(1199)) xor (layer6_outputs(940));
    layer7_outputs(4850) <= not(layer6_outputs(1246));
    layer7_outputs(4851) <= not((layer6_outputs(2510)) or (layer6_outputs(1147)));
    layer7_outputs(4852) <= (layer6_outputs(4820)) or (layer6_outputs(3786));
    layer7_outputs(4853) <= not(layer6_outputs(2746));
    layer7_outputs(4854) <= not(layer6_outputs(4945)) or (layer6_outputs(2167));
    layer7_outputs(4855) <= (layer6_outputs(1843)) and not (layer6_outputs(932));
    layer7_outputs(4856) <= layer6_outputs(2402);
    layer7_outputs(4857) <= layer6_outputs(4262);
    layer7_outputs(4858) <= layer6_outputs(3109);
    layer7_outputs(4859) <= (layer6_outputs(1913)) or (layer6_outputs(4278));
    layer7_outputs(4860) <= not(layer6_outputs(687));
    layer7_outputs(4861) <= not(layer6_outputs(2850)) or (layer6_outputs(1733));
    layer7_outputs(4862) <= not(layer6_outputs(3215)) or (layer6_outputs(2798));
    layer7_outputs(4863) <= (layer6_outputs(1872)) and (layer6_outputs(1482));
    layer7_outputs(4864) <= '1';
    layer7_outputs(4865) <= not(layer6_outputs(4833));
    layer7_outputs(4866) <= not(layer6_outputs(991));
    layer7_outputs(4867) <= (layer6_outputs(533)) and not (layer6_outputs(4390));
    layer7_outputs(4868) <= not(layer6_outputs(5057));
    layer7_outputs(4869) <= not(layer6_outputs(2660));
    layer7_outputs(4870) <= not(layer6_outputs(4149));
    layer7_outputs(4871) <= (layer6_outputs(4993)) xor (layer6_outputs(2739));
    layer7_outputs(4872) <= layer6_outputs(40);
    layer7_outputs(4873) <= (layer6_outputs(409)) and not (layer6_outputs(1632));
    layer7_outputs(4874) <= layer6_outputs(4369);
    layer7_outputs(4875) <= not(layer6_outputs(4590));
    layer7_outputs(4876) <= not(layer6_outputs(134));
    layer7_outputs(4877) <= not(layer6_outputs(1642));
    layer7_outputs(4878) <= not((layer6_outputs(2816)) or (layer6_outputs(125)));
    layer7_outputs(4879) <= not(layer6_outputs(1643)) or (layer6_outputs(890));
    layer7_outputs(4880) <= not((layer6_outputs(2577)) or (layer6_outputs(1840)));
    layer7_outputs(4881) <= layer6_outputs(1520);
    layer7_outputs(4882) <= not(layer6_outputs(667));
    layer7_outputs(4883) <= layer6_outputs(825);
    layer7_outputs(4884) <= (layer6_outputs(598)) or (layer6_outputs(2047));
    layer7_outputs(4885) <= not((layer6_outputs(1822)) xor (layer6_outputs(4679)));
    layer7_outputs(4886) <= layer6_outputs(2213);
    layer7_outputs(4887) <= layer6_outputs(1271);
    layer7_outputs(4888) <= not(layer6_outputs(3785)) or (layer6_outputs(3697));
    layer7_outputs(4889) <= not(layer6_outputs(4240));
    layer7_outputs(4890) <= not(layer6_outputs(142)) or (layer6_outputs(4540));
    layer7_outputs(4891) <= '1';
    layer7_outputs(4892) <= (layer6_outputs(1693)) or (layer6_outputs(4610));
    layer7_outputs(4893) <= (layer6_outputs(2416)) and not (layer6_outputs(3151));
    layer7_outputs(4894) <= not(layer6_outputs(3861));
    layer7_outputs(4895) <= layer6_outputs(499);
    layer7_outputs(4896) <= not(layer6_outputs(2978));
    layer7_outputs(4897) <= (layer6_outputs(270)) and not (layer6_outputs(3122));
    layer7_outputs(4898) <= layer6_outputs(2963);
    layer7_outputs(4899) <= not((layer6_outputs(3655)) or (layer6_outputs(1613)));
    layer7_outputs(4900) <= not(layer6_outputs(2679));
    layer7_outputs(4901) <= layer6_outputs(3970);
    layer7_outputs(4902) <= not(layer6_outputs(3212));
    layer7_outputs(4903) <= (layer6_outputs(3762)) xor (layer6_outputs(1762));
    layer7_outputs(4904) <= layer6_outputs(4895);
    layer7_outputs(4905) <= not(layer6_outputs(4694)) or (layer6_outputs(2074));
    layer7_outputs(4906) <= layer6_outputs(3625);
    layer7_outputs(4907) <= not((layer6_outputs(4490)) or (layer6_outputs(3815)));
    layer7_outputs(4908) <= layer6_outputs(4100);
    layer7_outputs(4909) <= '0';
    layer7_outputs(4910) <= layer6_outputs(3149);
    layer7_outputs(4911) <= (layer6_outputs(231)) and not (layer6_outputs(2233));
    layer7_outputs(4912) <= layer6_outputs(3092);
    layer7_outputs(4913) <= layer6_outputs(1158);
    layer7_outputs(4914) <= not((layer6_outputs(4393)) xor (layer6_outputs(3582)));
    layer7_outputs(4915) <= layer6_outputs(3126);
    layer7_outputs(4916) <= not(layer6_outputs(596));
    layer7_outputs(4917) <= layer6_outputs(3160);
    layer7_outputs(4918) <= (layer6_outputs(4475)) xor (layer6_outputs(4511));
    layer7_outputs(4919) <= not(layer6_outputs(205));
    layer7_outputs(4920) <= not(layer6_outputs(2903)) or (layer6_outputs(2625));
    layer7_outputs(4921) <= not((layer6_outputs(2565)) xor (layer6_outputs(3952)));
    layer7_outputs(4922) <= not(layer6_outputs(4030));
    layer7_outputs(4923) <= not((layer6_outputs(474)) or (layer6_outputs(4558)));
    layer7_outputs(4924) <= not((layer6_outputs(3601)) xor (layer6_outputs(3530)));
    layer7_outputs(4925) <= layer6_outputs(662);
    layer7_outputs(4926) <= (layer6_outputs(3311)) or (layer6_outputs(1399));
    layer7_outputs(4927) <= (layer6_outputs(973)) and not (layer6_outputs(2359));
    layer7_outputs(4928) <= not(layer6_outputs(3892));
    layer7_outputs(4929) <= (layer6_outputs(2795)) xor (layer6_outputs(996));
    layer7_outputs(4930) <= not(layer6_outputs(3610)) or (layer6_outputs(61));
    layer7_outputs(4931) <= not(layer6_outputs(3932)) or (layer6_outputs(3205));
    layer7_outputs(4932) <= not(layer6_outputs(1149));
    layer7_outputs(4933) <= not(layer6_outputs(1918));
    layer7_outputs(4934) <= (layer6_outputs(1704)) and not (layer6_outputs(2888));
    layer7_outputs(4935) <= layer6_outputs(2928);
    layer7_outputs(4936) <= layer6_outputs(3466);
    layer7_outputs(4937) <= not(layer6_outputs(1660));
    layer7_outputs(4938) <= layer6_outputs(4668);
    layer7_outputs(4939) <= not((layer6_outputs(4526)) xor (layer6_outputs(4718)));
    layer7_outputs(4940) <= '0';
    layer7_outputs(4941) <= layer6_outputs(1939);
    layer7_outputs(4942) <= not((layer6_outputs(3368)) or (layer6_outputs(606)));
    layer7_outputs(4943) <= (layer6_outputs(3912)) and not (layer6_outputs(3736));
    layer7_outputs(4944) <= layer6_outputs(2991);
    layer7_outputs(4945) <= (layer6_outputs(3880)) xor (layer6_outputs(1547));
    layer7_outputs(4946) <= layer6_outputs(3539);
    layer7_outputs(4947) <= layer6_outputs(13);
    layer7_outputs(4948) <= not(layer6_outputs(2282));
    layer7_outputs(4949) <= not(layer6_outputs(3783));
    layer7_outputs(4950) <= not(layer6_outputs(3879));
    layer7_outputs(4951) <= layer6_outputs(3848);
    layer7_outputs(4952) <= (layer6_outputs(1746)) and (layer6_outputs(939));
    layer7_outputs(4953) <= not((layer6_outputs(2047)) and (layer6_outputs(2042)));
    layer7_outputs(4954) <= (layer6_outputs(1631)) xor (layer6_outputs(2893));
    layer7_outputs(4955) <= layer6_outputs(593);
    layer7_outputs(4956) <= (layer6_outputs(3273)) and not (layer6_outputs(2634));
    layer7_outputs(4957) <= (layer6_outputs(1423)) xor (layer6_outputs(1906));
    layer7_outputs(4958) <= not(layer6_outputs(814));
    layer7_outputs(4959) <= layer6_outputs(4942);
    layer7_outputs(4960) <= not(layer6_outputs(1758));
    layer7_outputs(4961) <= not(layer6_outputs(1049));
    layer7_outputs(4962) <= layer6_outputs(1803);
    layer7_outputs(4963) <= not(layer6_outputs(5102));
    layer7_outputs(4964) <= layer6_outputs(2000);
    layer7_outputs(4965) <= layer6_outputs(4575);
    layer7_outputs(4966) <= not(layer6_outputs(3102));
    layer7_outputs(4967) <= (layer6_outputs(4953)) and not (layer6_outputs(900));
    layer7_outputs(4968) <= layer6_outputs(1231);
    layer7_outputs(4969) <= layer6_outputs(2080);
    layer7_outputs(4970) <= layer6_outputs(2330);
    layer7_outputs(4971) <= not(layer6_outputs(473));
    layer7_outputs(4972) <= layer6_outputs(1446);
    layer7_outputs(4973) <= not(layer6_outputs(2157));
    layer7_outputs(4974) <= not(layer6_outputs(718));
    layer7_outputs(4975) <= '1';
    layer7_outputs(4976) <= (layer6_outputs(1048)) and (layer6_outputs(4917));
    layer7_outputs(4977) <= not(layer6_outputs(4695));
    layer7_outputs(4978) <= (layer6_outputs(4770)) and not (layer6_outputs(857));
    layer7_outputs(4979) <= not(layer6_outputs(27));
    layer7_outputs(4980) <= not(layer6_outputs(2512));
    layer7_outputs(4981) <= not(layer6_outputs(517)) or (layer6_outputs(2487));
    layer7_outputs(4982) <= layer6_outputs(2889);
    layer7_outputs(4983) <= '0';
    layer7_outputs(4984) <= not((layer6_outputs(926)) xor (layer6_outputs(1128)));
    layer7_outputs(4985) <= (layer6_outputs(498)) and not (layer6_outputs(147));
    layer7_outputs(4986) <= '1';
    layer7_outputs(4987) <= layer6_outputs(1101);
    layer7_outputs(4988) <= layer6_outputs(525);
    layer7_outputs(4989) <= not((layer6_outputs(1557)) xor (layer6_outputs(2534)));
    layer7_outputs(4990) <= '1';
    layer7_outputs(4991) <= (layer6_outputs(2145)) and (layer6_outputs(1511));
    layer7_outputs(4992) <= (layer6_outputs(2303)) or (layer6_outputs(4151));
    layer7_outputs(4993) <= not(layer6_outputs(2376));
    layer7_outputs(4994) <= (layer6_outputs(3246)) or (layer6_outputs(3762));
    layer7_outputs(4995) <= not(layer6_outputs(1301));
    layer7_outputs(4996) <= (layer6_outputs(4712)) or (layer6_outputs(2114));
    layer7_outputs(4997) <= not(layer6_outputs(3437)) or (layer6_outputs(3970));
    layer7_outputs(4998) <= not((layer6_outputs(3945)) xor (layer6_outputs(2952)));
    layer7_outputs(4999) <= '1';
    layer7_outputs(5000) <= (layer6_outputs(1423)) or (layer6_outputs(2937));
    layer7_outputs(5001) <= (layer6_outputs(4025)) and not (layer6_outputs(4669));
    layer7_outputs(5002) <= not((layer6_outputs(4410)) xor (layer6_outputs(371)));
    layer7_outputs(5003) <= not(layer6_outputs(4984));
    layer7_outputs(5004) <= not(layer6_outputs(769));
    layer7_outputs(5005) <= (layer6_outputs(741)) and not (layer6_outputs(2136));
    layer7_outputs(5006) <= not(layer6_outputs(2700));
    layer7_outputs(5007) <= layer6_outputs(3679);
    layer7_outputs(5008) <= not((layer6_outputs(2548)) xor (layer6_outputs(1759)));
    layer7_outputs(5009) <= (layer6_outputs(3372)) and not (layer6_outputs(521));
    layer7_outputs(5010) <= layer6_outputs(4214);
    layer7_outputs(5011) <= layer6_outputs(3192);
    layer7_outputs(5012) <= (layer6_outputs(115)) and not (layer6_outputs(4506));
    layer7_outputs(5013) <= (layer6_outputs(3029)) and not (layer6_outputs(4927));
    layer7_outputs(5014) <= (layer6_outputs(4942)) and (layer6_outputs(3377));
    layer7_outputs(5015) <= not((layer6_outputs(4840)) or (layer6_outputs(1316)));
    layer7_outputs(5016) <= (layer6_outputs(3713)) and not (layer6_outputs(2884));
    layer7_outputs(5017) <= not(layer6_outputs(4329));
    layer7_outputs(5018) <= layer6_outputs(956);
    layer7_outputs(5019) <= not(layer6_outputs(4999));
    layer7_outputs(5020) <= layer6_outputs(2070);
    layer7_outputs(5021) <= not(layer6_outputs(934));
    layer7_outputs(5022) <= layer6_outputs(3185);
    layer7_outputs(5023) <= not(layer6_outputs(2253));
    layer7_outputs(5024) <= (layer6_outputs(4453)) xor (layer6_outputs(852));
    layer7_outputs(5025) <= (layer6_outputs(4108)) and not (layer6_outputs(3420));
    layer7_outputs(5026) <= not(layer6_outputs(1434)) or (layer6_outputs(126));
    layer7_outputs(5027) <= not(layer6_outputs(3419));
    layer7_outputs(5028) <= (layer6_outputs(4009)) and not (layer6_outputs(2149));
    layer7_outputs(5029) <= not(layer6_outputs(567));
    layer7_outputs(5030) <= layer6_outputs(5058);
    layer7_outputs(5031) <= layer6_outputs(2421);
    layer7_outputs(5032) <= (layer6_outputs(2868)) or (layer6_outputs(2035));
    layer7_outputs(5033) <= (layer6_outputs(2366)) xor (layer6_outputs(1017));
    layer7_outputs(5034) <= not(layer6_outputs(1831)) or (layer6_outputs(4951));
    layer7_outputs(5035) <= not(layer6_outputs(2325));
    layer7_outputs(5036) <= layer6_outputs(707);
    layer7_outputs(5037) <= not(layer6_outputs(1272)) or (layer6_outputs(4467));
    layer7_outputs(5038) <= (layer6_outputs(3926)) and not (layer6_outputs(2310));
    layer7_outputs(5039) <= not(layer6_outputs(1125));
    layer7_outputs(5040) <= '0';
    layer7_outputs(5041) <= not(layer6_outputs(3418)) or (layer6_outputs(339));
    layer7_outputs(5042) <= not(layer6_outputs(622)) or (layer6_outputs(693));
    layer7_outputs(5043) <= layer6_outputs(1443);
    layer7_outputs(5044) <= not((layer6_outputs(683)) or (layer6_outputs(1050)));
    layer7_outputs(5045) <= layer6_outputs(467);
    layer7_outputs(5046) <= not(layer6_outputs(3953));
    layer7_outputs(5047) <= layer6_outputs(2143);
    layer7_outputs(5048) <= not(layer6_outputs(3175));
    layer7_outputs(5049) <= not((layer6_outputs(1032)) xor (layer6_outputs(3866)));
    layer7_outputs(5050) <= (layer6_outputs(376)) and (layer6_outputs(4207));
    layer7_outputs(5051) <= not((layer6_outputs(1788)) xor (layer6_outputs(4818)));
    layer7_outputs(5052) <= not((layer6_outputs(4772)) xor (layer6_outputs(2593)));
    layer7_outputs(5053) <= not((layer6_outputs(4436)) or (layer6_outputs(155)));
    layer7_outputs(5054) <= not((layer6_outputs(736)) or (layer6_outputs(1868)));
    layer7_outputs(5055) <= (layer6_outputs(1787)) and not (layer6_outputs(317));
    layer7_outputs(5056) <= not(layer6_outputs(4374));
    layer7_outputs(5057) <= (layer6_outputs(1085)) and not (layer6_outputs(2813));
    layer7_outputs(5058) <= layer6_outputs(1924);
    layer7_outputs(5059) <= (layer6_outputs(4648)) and not (layer6_outputs(3094));
    layer7_outputs(5060) <= layer6_outputs(24);
    layer7_outputs(5061) <= not(layer6_outputs(4708));
    layer7_outputs(5062) <= (layer6_outputs(3999)) and not (layer6_outputs(3085));
    layer7_outputs(5063) <= not((layer6_outputs(2202)) and (layer6_outputs(1935)));
    layer7_outputs(5064) <= not(layer6_outputs(10)) or (layer6_outputs(2974));
    layer7_outputs(5065) <= not(layer6_outputs(4952));
    layer7_outputs(5066) <= '0';
    layer7_outputs(5067) <= not((layer6_outputs(2954)) and (layer6_outputs(2820)));
    layer7_outputs(5068) <= (layer6_outputs(680)) and (layer6_outputs(4279));
    layer7_outputs(5069) <= (layer6_outputs(4021)) xor (layer6_outputs(3077));
    layer7_outputs(5070) <= (layer6_outputs(2720)) or (layer6_outputs(4786));
    layer7_outputs(5071) <= layer6_outputs(1625);
    layer7_outputs(5072) <= layer6_outputs(1505);
    layer7_outputs(5073) <= layer6_outputs(1758);
    layer7_outputs(5074) <= (layer6_outputs(2882)) and (layer6_outputs(3836));
    layer7_outputs(5075) <= (layer6_outputs(3134)) or (layer6_outputs(4461));
    layer7_outputs(5076) <= layer6_outputs(1263);
    layer7_outputs(5077) <= (layer6_outputs(435)) xor (layer6_outputs(2662));
    layer7_outputs(5078) <= layer6_outputs(1683);
    layer7_outputs(5079) <= layer6_outputs(4317);
    layer7_outputs(5080) <= layer6_outputs(1441);
    layer7_outputs(5081) <= not(layer6_outputs(3395));
    layer7_outputs(5082) <= layer6_outputs(511);
    layer7_outputs(5083) <= not(layer6_outputs(2203));
    layer7_outputs(5084) <= not((layer6_outputs(771)) and (layer6_outputs(1987)));
    layer7_outputs(5085) <= (layer6_outputs(2582)) and not (layer6_outputs(869));
    layer7_outputs(5086) <= not(layer6_outputs(834));
    layer7_outputs(5087) <= not(layer6_outputs(1147)) or (layer6_outputs(4956));
    layer7_outputs(5088) <= (layer6_outputs(3063)) and not (layer6_outputs(3964));
    layer7_outputs(5089) <= not(layer6_outputs(4208));
    layer7_outputs(5090) <= not((layer6_outputs(3671)) xor (layer6_outputs(985)));
    layer7_outputs(5091) <= (layer6_outputs(1481)) xor (layer6_outputs(4641));
    layer7_outputs(5092) <= not((layer6_outputs(2342)) or (layer6_outputs(3936)));
    layer7_outputs(5093) <= (layer6_outputs(791)) and (layer6_outputs(3744));
    layer7_outputs(5094) <= not((layer6_outputs(309)) or (layer6_outputs(4269)));
    layer7_outputs(5095) <= (layer6_outputs(4087)) xor (layer6_outputs(939));
    layer7_outputs(5096) <= not(layer6_outputs(1420));
    layer7_outputs(5097) <= '0';
    layer7_outputs(5098) <= layer6_outputs(471);
    layer7_outputs(5099) <= not(layer6_outputs(2863)) or (layer6_outputs(2307));
    layer7_outputs(5100) <= not(layer6_outputs(3101));
    layer7_outputs(5101) <= not((layer6_outputs(4356)) or (layer6_outputs(3794)));
    layer7_outputs(5102) <= not((layer6_outputs(2044)) and (layer6_outputs(2473)));
    layer7_outputs(5103) <= not(layer6_outputs(1058)) or (layer6_outputs(3183));
    layer7_outputs(5104) <= layer6_outputs(2887);
    layer7_outputs(5105) <= not(layer6_outputs(2964));
    layer7_outputs(5106) <= not(layer6_outputs(3755));
    layer7_outputs(5107) <= not((layer6_outputs(4080)) xor (layer6_outputs(3711)));
    layer7_outputs(5108) <= (layer6_outputs(5061)) xor (layer6_outputs(4704));
    layer7_outputs(5109) <= layer6_outputs(1942);
    layer7_outputs(5110) <= layer6_outputs(2982);
    layer7_outputs(5111) <= not(layer6_outputs(2292));
    layer7_outputs(5112) <= layer6_outputs(2780);
    layer7_outputs(5113) <= not(layer6_outputs(5033));
    layer7_outputs(5114) <= layer6_outputs(3907);
    layer7_outputs(5115) <= not(layer6_outputs(3293));
    layer7_outputs(5116) <= (layer6_outputs(1290)) or (layer6_outputs(1058));
    layer7_outputs(5117) <= not((layer6_outputs(144)) and (layer6_outputs(989)));
    layer7_outputs(5118) <= layer6_outputs(1667);
    layer7_outputs(5119) <= layer6_outputs(69);
    layer8_outputs(0) <= (layer7_outputs(2963)) and not (layer7_outputs(2875));
    layer8_outputs(1) <= not(layer7_outputs(2835)) or (layer7_outputs(4783));
    layer8_outputs(2) <= (layer7_outputs(2749)) xor (layer7_outputs(4179));
    layer8_outputs(3) <= (layer7_outputs(5110)) and (layer7_outputs(2982));
    layer8_outputs(4) <= not(layer7_outputs(4647));
    layer8_outputs(5) <= (layer7_outputs(2319)) xor (layer7_outputs(2001));
    layer8_outputs(6) <= not(layer7_outputs(1556));
    layer8_outputs(7) <= not(layer7_outputs(2603));
    layer8_outputs(8) <= '1';
    layer8_outputs(9) <= not(layer7_outputs(541));
    layer8_outputs(10) <= not(layer7_outputs(1362)) or (layer7_outputs(3286));
    layer8_outputs(11) <= layer7_outputs(1912);
    layer8_outputs(12) <= layer7_outputs(479);
    layer8_outputs(13) <= not(layer7_outputs(1655)) or (layer7_outputs(776));
    layer8_outputs(14) <= layer7_outputs(2510);
    layer8_outputs(15) <= layer7_outputs(2207);
    layer8_outputs(16) <= layer7_outputs(1061);
    layer8_outputs(17) <= layer7_outputs(1516);
    layer8_outputs(18) <= layer7_outputs(3920);
    layer8_outputs(19) <= not(layer7_outputs(3654));
    layer8_outputs(20) <= (layer7_outputs(776)) and (layer7_outputs(1139));
    layer8_outputs(21) <= (layer7_outputs(2377)) and (layer7_outputs(2549));
    layer8_outputs(22) <= (layer7_outputs(1135)) and not (layer7_outputs(4235));
    layer8_outputs(23) <= not((layer7_outputs(3103)) xor (layer7_outputs(4715)));
    layer8_outputs(24) <= layer7_outputs(3079);
    layer8_outputs(25) <= not(layer7_outputs(702));
    layer8_outputs(26) <= not(layer7_outputs(1058));
    layer8_outputs(27) <= (layer7_outputs(1957)) xor (layer7_outputs(766));
    layer8_outputs(28) <= not(layer7_outputs(769));
    layer8_outputs(29) <= (layer7_outputs(3834)) and not (layer7_outputs(2769));
    layer8_outputs(30) <= not(layer7_outputs(1196));
    layer8_outputs(31) <= not((layer7_outputs(4733)) or (layer7_outputs(1893)));
    layer8_outputs(32) <= not(layer7_outputs(542));
    layer8_outputs(33) <= not((layer7_outputs(1563)) or (layer7_outputs(4981)));
    layer8_outputs(34) <= not(layer7_outputs(2555));
    layer8_outputs(35) <= not(layer7_outputs(2117)) or (layer7_outputs(1688));
    layer8_outputs(36) <= (layer7_outputs(690)) xor (layer7_outputs(2575));
    layer8_outputs(37) <= not(layer7_outputs(43));
    layer8_outputs(38) <= not(layer7_outputs(3800));
    layer8_outputs(39) <= not(layer7_outputs(3612)) or (layer7_outputs(4125));
    layer8_outputs(40) <= (layer7_outputs(1824)) xor (layer7_outputs(2688));
    layer8_outputs(41) <= (layer7_outputs(4092)) xor (layer7_outputs(5029));
    layer8_outputs(42) <= layer7_outputs(792);
    layer8_outputs(43) <= layer7_outputs(4485);
    layer8_outputs(44) <= (layer7_outputs(2777)) and (layer7_outputs(2270));
    layer8_outputs(45) <= not((layer7_outputs(1759)) xor (layer7_outputs(2458)));
    layer8_outputs(46) <= layer7_outputs(8);
    layer8_outputs(47) <= layer7_outputs(2640);
    layer8_outputs(48) <= (layer7_outputs(3486)) xor (layer7_outputs(2601));
    layer8_outputs(49) <= layer7_outputs(4941);
    layer8_outputs(50) <= layer7_outputs(1467);
    layer8_outputs(51) <= layer7_outputs(1683);
    layer8_outputs(52) <= (layer7_outputs(1052)) xor (layer7_outputs(4370));
    layer8_outputs(53) <= not(layer7_outputs(3246)) or (layer7_outputs(1145));
    layer8_outputs(54) <= not(layer7_outputs(4207)) or (layer7_outputs(2407));
    layer8_outputs(55) <= not(layer7_outputs(98)) or (layer7_outputs(481));
    layer8_outputs(56) <= not((layer7_outputs(2577)) or (layer7_outputs(1010)));
    layer8_outputs(57) <= not(layer7_outputs(3365));
    layer8_outputs(58) <= not((layer7_outputs(2970)) xor (layer7_outputs(1101)));
    layer8_outputs(59) <= (layer7_outputs(131)) xor (layer7_outputs(1379));
    layer8_outputs(60) <= (layer7_outputs(4461)) xor (layer7_outputs(3763));
    layer8_outputs(61) <= layer7_outputs(1939);
    layer8_outputs(62) <= not(layer7_outputs(2397));
    layer8_outputs(63) <= (layer7_outputs(4846)) xor (layer7_outputs(2506));
    layer8_outputs(64) <= not((layer7_outputs(1906)) xor (layer7_outputs(4732)));
    layer8_outputs(65) <= '1';
    layer8_outputs(66) <= not(layer7_outputs(1718));
    layer8_outputs(67) <= (layer7_outputs(195)) xor (layer7_outputs(1975));
    layer8_outputs(68) <= layer7_outputs(4748);
    layer8_outputs(69) <= layer7_outputs(1967);
    layer8_outputs(70) <= not(layer7_outputs(4501));
    layer8_outputs(71) <= not(layer7_outputs(2060));
    layer8_outputs(72) <= not(layer7_outputs(726)) or (layer7_outputs(2274));
    layer8_outputs(73) <= not(layer7_outputs(1367));
    layer8_outputs(74) <= (layer7_outputs(2686)) and (layer7_outputs(5093));
    layer8_outputs(75) <= layer7_outputs(988);
    layer8_outputs(76) <= not(layer7_outputs(1315)) or (layer7_outputs(4592));
    layer8_outputs(77) <= (layer7_outputs(4725)) xor (layer7_outputs(2249));
    layer8_outputs(78) <= layer7_outputs(1794);
    layer8_outputs(79) <= layer7_outputs(573);
    layer8_outputs(80) <= not(layer7_outputs(5031)) or (layer7_outputs(429));
    layer8_outputs(81) <= not((layer7_outputs(21)) xor (layer7_outputs(4515)));
    layer8_outputs(82) <= not(layer7_outputs(1289));
    layer8_outputs(83) <= layer7_outputs(2200);
    layer8_outputs(84) <= not(layer7_outputs(4671));
    layer8_outputs(85) <= (layer7_outputs(692)) and (layer7_outputs(424));
    layer8_outputs(86) <= not(layer7_outputs(3617));
    layer8_outputs(87) <= not(layer7_outputs(2408));
    layer8_outputs(88) <= not(layer7_outputs(2760));
    layer8_outputs(89) <= (layer7_outputs(2624)) xor (layer7_outputs(703));
    layer8_outputs(90) <= not((layer7_outputs(446)) xor (layer7_outputs(1015)));
    layer8_outputs(91) <= layer7_outputs(2736);
    layer8_outputs(92) <= (layer7_outputs(1602)) xor (layer7_outputs(1545));
    layer8_outputs(93) <= layer7_outputs(2382);
    layer8_outputs(94) <= not(layer7_outputs(3761));
    layer8_outputs(95) <= (layer7_outputs(2244)) and not (layer7_outputs(4135));
    layer8_outputs(96) <= layer7_outputs(4183);
    layer8_outputs(97) <= layer7_outputs(3942);
    layer8_outputs(98) <= layer7_outputs(3127);
    layer8_outputs(99) <= not((layer7_outputs(3047)) xor (layer7_outputs(3859)));
    layer8_outputs(100) <= not(layer7_outputs(2885));
    layer8_outputs(101) <= not(layer7_outputs(3868));
    layer8_outputs(102) <= not(layer7_outputs(3923));
    layer8_outputs(103) <= '1';
    layer8_outputs(104) <= (layer7_outputs(3479)) and not (layer7_outputs(2062));
    layer8_outputs(105) <= not((layer7_outputs(2626)) xor (layer7_outputs(1554)));
    layer8_outputs(106) <= not((layer7_outputs(4226)) or (layer7_outputs(3857)));
    layer8_outputs(107) <= (layer7_outputs(2479)) and not (layer7_outputs(3996));
    layer8_outputs(108) <= not((layer7_outputs(1978)) or (layer7_outputs(102)));
    layer8_outputs(109) <= (layer7_outputs(437)) or (layer7_outputs(3691));
    layer8_outputs(110) <= not(layer7_outputs(1612));
    layer8_outputs(111) <= not(layer7_outputs(3846)) or (layer7_outputs(591));
    layer8_outputs(112) <= not(layer7_outputs(4369)) or (layer7_outputs(3161));
    layer8_outputs(113) <= layer7_outputs(722);
    layer8_outputs(114) <= layer7_outputs(4232);
    layer8_outputs(115) <= not(layer7_outputs(2688));
    layer8_outputs(116) <= not(layer7_outputs(1051));
    layer8_outputs(117) <= layer7_outputs(2224);
    layer8_outputs(118) <= (layer7_outputs(4816)) xor (layer7_outputs(3347));
    layer8_outputs(119) <= layer7_outputs(2817);
    layer8_outputs(120) <= (layer7_outputs(4787)) xor (layer7_outputs(2384));
    layer8_outputs(121) <= not((layer7_outputs(4296)) xor (layer7_outputs(1488)));
    layer8_outputs(122) <= layer7_outputs(2055);
    layer8_outputs(123) <= (layer7_outputs(1380)) xor (layer7_outputs(218));
    layer8_outputs(124) <= layer7_outputs(1569);
    layer8_outputs(125) <= not(layer7_outputs(302));
    layer8_outputs(126) <= layer7_outputs(1930);
    layer8_outputs(127) <= not((layer7_outputs(773)) xor (layer7_outputs(907)));
    layer8_outputs(128) <= not(layer7_outputs(3990));
    layer8_outputs(129) <= layer7_outputs(2957);
    layer8_outputs(130) <= (layer7_outputs(3879)) and not (layer7_outputs(182));
    layer8_outputs(131) <= (layer7_outputs(2999)) or (layer7_outputs(4616));
    layer8_outputs(132) <= not((layer7_outputs(5069)) xor (layer7_outputs(2583)));
    layer8_outputs(133) <= (layer7_outputs(4400)) and (layer7_outputs(782));
    layer8_outputs(134) <= layer7_outputs(2669);
    layer8_outputs(135) <= (layer7_outputs(4018)) or (layer7_outputs(249));
    layer8_outputs(136) <= layer7_outputs(3046);
    layer8_outputs(137) <= (layer7_outputs(1895)) or (layer7_outputs(2589));
    layer8_outputs(138) <= not(layer7_outputs(3091));
    layer8_outputs(139) <= layer7_outputs(2803);
    layer8_outputs(140) <= layer7_outputs(1405);
    layer8_outputs(141) <= not(layer7_outputs(3231));
    layer8_outputs(142) <= not(layer7_outputs(1008));
    layer8_outputs(143) <= (layer7_outputs(3254)) xor (layer7_outputs(1947));
    layer8_outputs(144) <= layer7_outputs(4819);
    layer8_outputs(145) <= not((layer7_outputs(342)) xor (layer7_outputs(2827)));
    layer8_outputs(146) <= not(layer7_outputs(4979));
    layer8_outputs(147) <= not(layer7_outputs(1152));
    layer8_outputs(148) <= not(layer7_outputs(3084));
    layer8_outputs(149) <= (layer7_outputs(1834)) xor (layer7_outputs(2793));
    layer8_outputs(150) <= not(layer7_outputs(4918));
    layer8_outputs(151) <= not(layer7_outputs(3067)) or (layer7_outputs(4682));
    layer8_outputs(152) <= not(layer7_outputs(1662));
    layer8_outputs(153) <= layer7_outputs(1035);
    layer8_outputs(154) <= (layer7_outputs(1879)) xor (layer7_outputs(1249));
    layer8_outputs(155) <= (layer7_outputs(4611)) xor (layer7_outputs(2756));
    layer8_outputs(156) <= not(layer7_outputs(721)) or (layer7_outputs(4893));
    layer8_outputs(157) <= (layer7_outputs(731)) and not (layer7_outputs(2445));
    layer8_outputs(158) <= not((layer7_outputs(2950)) xor (layer7_outputs(2147)));
    layer8_outputs(159) <= layer7_outputs(4203);
    layer8_outputs(160) <= not(layer7_outputs(4814));
    layer8_outputs(161) <= layer7_outputs(487);
    layer8_outputs(162) <= not((layer7_outputs(453)) and (layer7_outputs(3067)));
    layer8_outputs(163) <= not((layer7_outputs(4455)) xor (layer7_outputs(1542)));
    layer8_outputs(164) <= layer7_outputs(4777);
    layer8_outputs(165) <= layer7_outputs(2397);
    layer8_outputs(166) <= (layer7_outputs(1155)) xor (layer7_outputs(698));
    layer8_outputs(167) <= not(layer7_outputs(3914));
    layer8_outputs(168) <= (layer7_outputs(3238)) and (layer7_outputs(1087));
    layer8_outputs(169) <= (layer7_outputs(3914)) and not (layer7_outputs(975));
    layer8_outputs(170) <= layer7_outputs(4774);
    layer8_outputs(171) <= (layer7_outputs(4033)) or (layer7_outputs(2400));
    layer8_outputs(172) <= not(layer7_outputs(2091));
    layer8_outputs(173) <= (layer7_outputs(4493)) and not (layer7_outputs(2552));
    layer8_outputs(174) <= not((layer7_outputs(1171)) and (layer7_outputs(1570)));
    layer8_outputs(175) <= not((layer7_outputs(1729)) and (layer7_outputs(1511)));
    layer8_outputs(176) <= not(layer7_outputs(3246));
    layer8_outputs(177) <= not((layer7_outputs(3680)) or (layer7_outputs(4634)));
    layer8_outputs(178) <= (layer7_outputs(2310)) xor (layer7_outputs(12));
    layer8_outputs(179) <= not(layer7_outputs(4533)) or (layer7_outputs(1351));
    layer8_outputs(180) <= (layer7_outputs(2178)) xor (layer7_outputs(4040));
    layer8_outputs(181) <= (layer7_outputs(4130)) xor (layer7_outputs(3069));
    layer8_outputs(182) <= not(layer7_outputs(4313));
    layer8_outputs(183) <= '1';
    layer8_outputs(184) <= not(layer7_outputs(1808));
    layer8_outputs(185) <= not(layer7_outputs(2006)) or (layer7_outputs(2566));
    layer8_outputs(186) <= not((layer7_outputs(52)) and (layer7_outputs(1291)));
    layer8_outputs(187) <= layer7_outputs(491);
    layer8_outputs(188) <= layer7_outputs(4734);
    layer8_outputs(189) <= not(layer7_outputs(1217));
    layer8_outputs(190) <= (layer7_outputs(83)) xor (layer7_outputs(2267));
    layer8_outputs(191) <= layer7_outputs(2772);
    layer8_outputs(192) <= (layer7_outputs(1796)) xor (layer7_outputs(455));
    layer8_outputs(193) <= not(layer7_outputs(4212));
    layer8_outputs(194) <= not(layer7_outputs(4664));
    layer8_outputs(195) <= not((layer7_outputs(3245)) xor (layer7_outputs(1002)));
    layer8_outputs(196) <= not((layer7_outputs(2319)) xor (layer7_outputs(3178)));
    layer8_outputs(197) <= layer7_outputs(2649);
    layer8_outputs(198) <= not((layer7_outputs(3338)) xor (layer7_outputs(2062)));
    layer8_outputs(199) <= layer7_outputs(2619);
    layer8_outputs(200) <= not(layer7_outputs(1996));
    layer8_outputs(201) <= not((layer7_outputs(958)) xor (layer7_outputs(3772)));
    layer8_outputs(202) <= not((layer7_outputs(2965)) xor (layer7_outputs(4690)));
    layer8_outputs(203) <= not(layer7_outputs(2766));
    layer8_outputs(204) <= not(layer7_outputs(1587));
    layer8_outputs(205) <= not(layer7_outputs(4088)) or (layer7_outputs(3796));
    layer8_outputs(206) <= (layer7_outputs(4545)) and (layer7_outputs(2546));
    layer8_outputs(207) <= not((layer7_outputs(298)) xor (layer7_outputs(1269)));
    layer8_outputs(208) <= not((layer7_outputs(2971)) xor (layer7_outputs(2626)));
    layer8_outputs(209) <= not((layer7_outputs(1751)) xor (layer7_outputs(143)));
    layer8_outputs(210) <= (layer7_outputs(1262)) and not (layer7_outputs(370));
    layer8_outputs(211) <= not(layer7_outputs(1330));
    layer8_outputs(212) <= (layer7_outputs(2126)) xor (layer7_outputs(575));
    layer8_outputs(213) <= not(layer7_outputs(2629));
    layer8_outputs(214) <= (layer7_outputs(972)) and (layer7_outputs(3080));
    layer8_outputs(215) <= not(layer7_outputs(4067)) or (layer7_outputs(4637));
    layer8_outputs(216) <= layer7_outputs(3542);
    layer8_outputs(217) <= layer7_outputs(4542);
    layer8_outputs(218) <= not((layer7_outputs(1952)) xor (layer7_outputs(833)));
    layer8_outputs(219) <= not((layer7_outputs(344)) xor (layer7_outputs(923)));
    layer8_outputs(220) <= layer7_outputs(4039);
    layer8_outputs(221) <= not(layer7_outputs(196));
    layer8_outputs(222) <= not(layer7_outputs(2091)) or (layer7_outputs(1756));
    layer8_outputs(223) <= layer7_outputs(3064);
    layer8_outputs(224) <= not(layer7_outputs(1072));
    layer8_outputs(225) <= (layer7_outputs(2677)) xor (layer7_outputs(2913));
    layer8_outputs(226) <= not((layer7_outputs(2665)) xor (layer7_outputs(2684)));
    layer8_outputs(227) <= layer7_outputs(460);
    layer8_outputs(228) <= layer7_outputs(2123);
    layer8_outputs(229) <= layer7_outputs(3746);
    layer8_outputs(230) <= (layer7_outputs(4792)) and not (layer7_outputs(4245));
    layer8_outputs(231) <= (layer7_outputs(3017)) xor (layer7_outputs(184));
    layer8_outputs(232) <= layer7_outputs(3705);
    layer8_outputs(233) <= layer7_outputs(3203);
    layer8_outputs(234) <= layer7_outputs(4416);
    layer8_outputs(235) <= not(layer7_outputs(1134));
    layer8_outputs(236) <= layer7_outputs(665);
    layer8_outputs(237) <= (layer7_outputs(3425)) and (layer7_outputs(788));
    layer8_outputs(238) <= not(layer7_outputs(409));
    layer8_outputs(239) <= (layer7_outputs(3263)) xor (layer7_outputs(825));
    layer8_outputs(240) <= not((layer7_outputs(4267)) xor (layer7_outputs(517)));
    layer8_outputs(241) <= not((layer7_outputs(2190)) xor (layer7_outputs(3724)));
    layer8_outputs(242) <= (layer7_outputs(407)) and (layer7_outputs(2728));
    layer8_outputs(243) <= not(layer7_outputs(1850));
    layer8_outputs(244) <= not((layer7_outputs(2789)) xor (layer7_outputs(3667)));
    layer8_outputs(245) <= not(layer7_outputs(4034));
    layer8_outputs(246) <= layer7_outputs(1851);
    layer8_outputs(247) <= not((layer7_outputs(4976)) xor (layer7_outputs(3638)));
    layer8_outputs(248) <= layer7_outputs(928);
    layer8_outputs(249) <= (layer7_outputs(3912)) and not (layer7_outputs(1129));
    layer8_outputs(250) <= (layer7_outputs(1099)) or (layer7_outputs(4196));
    layer8_outputs(251) <= layer7_outputs(1029);
    layer8_outputs(252) <= layer7_outputs(2355);
    layer8_outputs(253) <= (layer7_outputs(3108)) xor (layer7_outputs(4074));
    layer8_outputs(254) <= not(layer7_outputs(1084));
    layer8_outputs(255) <= layer7_outputs(3210);
    layer8_outputs(256) <= (layer7_outputs(2396)) xor (layer7_outputs(3924));
    layer8_outputs(257) <= not((layer7_outputs(2841)) and (layer7_outputs(1382)));
    layer8_outputs(258) <= not(layer7_outputs(4169));
    layer8_outputs(259) <= not(layer7_outputs(662));
    layer8_outputs(260) <= not(layer7_outputs(3148)) or (layer7_outputs(4350));
    layer8_outputs(261) <= not(layer7_outputs(1400));
    layer8_outputs(262) <= not((layer7_outputs(718)) xor (layer7_outputs(2431)));
    layer8_outputs(263) <= not((layer7_outputs(505)) or (layer7_outputs(3416)));
    layer8_outputs(264) <= (layer7_outputs(778)) and not (layer7_outputs(4676));
    layer8_outputs(265) <= (layer7_outputs(2343)) or (layer7_outputs(1753));
    layer8_outputs(266) <= not(layer7_outputs(1674));
    layer8_outputs(267) <= not(layer7_outputs(1198)) or (layer7_outputs(1928));
    layer8_outputs(268) <= not(layer7_outputs(1648));
    layer8_outputs(269) <= not(layer7_outputs(1466)) or (layer7_outputs(4152));
    layer8_outputs(270) <= layer7_outputs(4691);
    layer8_outputs(271) <= not((layer7_outputs(2169)) xor (layer7_outputs(764)));
    layer8_outputs(272) <= not(layer7_outputs(2933));
    layer8_outputs(273) <= not(layer7_outputs(1107));
    layer8_outputs(274) <= not(layer7_outputs(1902));
    layer8_outputs(275) <= not((layer7_outputs(3029)) xor (layer7_outputs(3862)));
    layer8_outputs(276) <= not((layer7_outputs(1876)) and (layer7_outputs(1329)));
    layer8_outputs(277) <= not(layer7_outputs(1984));
    layer8_outputs(278) <= not((layer7_outputs(4829)) xor (layer7_outputs(4398)));
    layer8_outputs(279) <= not(layer7_outputs(4872));
    layer8_outputs(280) <= layer7_outputs(5057);
    layer8_outputs(281) <= not((layer7_outputs(2271)) or (layer7_outputs(1315)));
    layer8_outputs(282) <= not(layer7_outputs(4279));
    layer8_outputs(283) <= not(layer7_outputs(785));
    layer8_outputs(284) <= not((layer7_outputs(5054)) xor (layer7_outputs(4653)));
    layer8_outputs(285) <= (layer7_outputs(2440)) xor (layer7_outputs(5086));
    layer8_outputs(286) <= not((layer7_outputs(3082)) or (layer7_outputs(4111)));
    layer8_outputs(287) <= not(layer7_outputs(1186)) or (layer7_outputs(2443));
    layer8_outputs(288) <= not((layer7_outputs(2943)) and (layer7_outputs(5098)));
    layer8_outputs(289) <= not(layer7_outputs(3730));
    layer8_outputs(290) <= (layer7_outputs(3932)) and (layer7_outputs(1997));
    layer8_outputs(291) <= (layer7_outputs(2817)) and not (layer7_outputs(1309));
    layer8_outputs(292) <= (layer7_outputs(1839)) and not (layer7_outputs(2650));
    layer8_outputs(293) <= layer7_outputs(42);
    layer8_outputs(294) <= layer7_outputs(4774);
    layer8_outputs(295) <= layer7_outputs(4203);
    layer8_outputs(296) <= layer7_outputs(4765);
    layer8_outputs(297) <= not((layer7_outputs(1331)) xor (layer7_outputs(3128)));
    layer8_outputs(298) <= not(layer7_outputs(4952));
    layer8_outputs(299) <= layer7_outputs(4050);
    layer8_outputs(300) <= (layer7_outputs(3411)) xor (layer7_outputs(4205));
    layer8_outputs(301) <= layer7_outputs(1592);
    layer8_outputs(302) <= (layer7_outputs(3781)) or (layer7_outputs(321));
    layer8_outputs(303) <= not((layer7_outputs(2300)) xor (layer7_outputs(2251)));
    layer8_outputs(304) <= not((layer7_outputs(4326)) and (layer7_outputs(2175)));
    layer8_outputs(305) <= layer7_outputs(565);
    layer8_outputs(306) <= layer7_outputs(1509);
    layer8_outputs(307) <= layer7_outputs(3923);
    layer8_outputs(308) <= not((layer7_outputs(1807)) or (layer7_outputs(1031)));
    layer8_outputs(309) <= not(layer7_outputs(2630));
    layer8_outputs(310) <= layer7_outputs(3282);
    layer8_outputs(311) <= not(layer7_outputs(1177));
    layer8_outputs(312) <= (layer7_outputs(3085)) and not (layer7_outputs(4041));
    layer8_outputs(313) <= (layer7_outputs(2646)) xor (layer7_outputs(3668));
    layer8_outputs(314) <= layer7_outputs(821);
    layer8_outputs(315) <= not((layer7_outputs(2130)) xor (layer7_outputs(2063)));
    layer8_outputs(316) <= not((layer7_outputs(4836)) or (layer7_outputs(4468)));
    layer8_outputs(317) <= (layer7_outputs(1546)) xor (layer7_outputs(4433));
    layer8_outputs(318) <= (layer7_outputs(872)) xor (layer7_outputs(1669));
    layer8_outputs(319) <= not(layer7_outputs(3218));
    layer8_outputs(320) <= not((layer7_outputs(619)) xor (layer7_outputs(4718)));
    layer8_outputs(321) <= (layer7_outputs(1319)) and not (layer7_outputs(889));
    layer8_outputs(322) <= layer7_outputs(877);
    layer8_outputs(323) <= not(layer7_outputs(1462));
    layer8_outputs(324) <= not(layer7_outputs(1172));
    layer8_outputs(325) <= layer7_outputs(554);
    layer8_outputs(326) <= (layer7_outputs(1362)) xor (layer7_outputs(4537));
    layer8_outputs(327) <= not(layer7_outputs(2378)) or (layer7_outputs(632));
    layer8_outputs(328) <= (layer7_outputs(2134)) xor (layer7_outputs(2884));
    layer8_outputs(329) <= not(layer7_outputs(1205)) or (layer7_outputs(4966));
    layer8_outputs(330) <= layer7_outputs(3198);
    layer8_outputs(331) <= layer7_outputs(232);
    layer8_outputs(332) <= not(layer7_outputs(2603));
    layer8_outputs(333) <= not(layer7_outputs(658)) or (layer7_outputs(837));
    layer8_outputs(334) <= (layer7_outputs(1468)) xor (layer7_outputs(4201));
    layer8_outputs(335) <= not(layer7_outputs(3757));
    layer8_outputs(336) <= not(layer7_outputs(1690));
    layer8_outputs(337) <= not(layer7_outputs(3877)) or (layer7_outputs(2157));
    layer8_outputs(338) <= not(layer7_outputs(4869));
    layer8_outputs(339) <= not((layer7_outputs(3035)) xor (layer7_outputs(3255)));
    layer8_outputs(340) <= (layer7_outputs(4935)) and (layer7_outputs(1040));
    layer8_outputs(341) <= layer7_outputs(615);
    layer8_outputs(342) <= not((layer7_outputs(3136)) or (layer7_outputs(2018)));
    layer8_outputs(343) <= not(layer7_outputs(168));
    layer8_outputs(344) <= not(layer7_outputs(3288)) or (layer7_outputs(1725));
    layer8_outputs(345) <= not((layer7_outputs(2612)) and (layer7_outputs(2097)));
    layer8_outputs(346) <= layer7_outputs(2246);
    layer8_outputs(347) <= not(layer7_outputs(108));
    layer8_outputs(348) <= layer7_outputs(371);
    layer8_outputs(349) <= layer7_outputs(4832);
    layer8_outputs(350) <= layer7_outputs(3195);
    layer8_outputs(351) <= (layer7_outputs(448)) and (layer7_outputs(642));
    layer8_outputs(352) <= not(layer7_outputs(2949)) or (layer7_outputs(667));
    layer8_outputs(353) <= (layer7_outputs(59)) xor (layer7_outputs(2886));
    layer8_outputs(354) <= not(layer7_outputs(2800));
    layer8_outputs(355) <= layer7_outputs(4076);
    layer8_outputs(356) <= layer7_outputs(3429);
    layer8_outputs(357) <= (layer7_outputs(3080)) xor (layer7_outputs(1654));
    layer8_outputs(358) <= not((layer7_outputs(1689)) xor (layer7_outputs(682)));
    layer8_outputs(359) <= layer7_outputs(2620);
    layer8_outputs(360) <= layer7_outputs(3958);
    layer8_outputs(361) <= not((layer7_outputs(4988)) and (layer7_outputs(907)));
    layer8_outputs(362) <= (layer7_outputs(2184)) xor (layer7_outputs(150));
    layer8_outputs(363) <= (layer7_outputs(2389)) and (layer7_outputs(2692));
    layer8_outputs(364) <= not(layer7_outputs(4144));
    layer8_outputs(365) <= not(layer7_outputs(2931));
    layer8_outputs(366) <= not(layer7_outputs(2898));
    layer8_outputs(367) <= not(layer7_outputs(2402));
    layer8_outputs(368) <= layer7_outputs(1148);
    layer8_outputs(369) <= (layer7_outputs(3550)) xor (layer7_outputs(1905));
    layer8_outputs(370) <= layer7_outputs(3159);
    layer8_outputs(371) <= '1';
    layer8_outputs(372) <= layer7_outputs(3277);
    layer8_outputs(373) <= layer7_outputs(2376);
    layer8_outputs(374) <= not((layer7_outputs(911)) or (layer7_outputs(3869)));
    layer8_outputs(375) <= layer7_outputs(4868);
    layer8_outputs(376) <= not(layer7_outputs(3511)) or (layer7_outputs(1117));
    layer8_outputs(377) <= not((layer7_outputs(3957)) xor (layer7_outputs(3279)));
    layer8_outputs(378) <= not((layer7_outputs(1182)) or (layer7_outputs(3901)));
    layer8_outputs(379) <= layer7_outputs(1132);
    layer8_outputs(380) <= not(layer7_outputs(2815)) or (layer7_outputs(4444));
    layer8_outputs(381) <= not(layer7_outputs(1883));
    layer8_outputs(382) <= not(layer7_outputs(892)) or (layer7_outputs(918));
    layer8_outputs(383) <= not(layer7_outputs(4596)) or (layer7_outputs(1267));
    layer8_outputs(384) <= not(layer7_outputs(2636));
    layer8_outputs(385) <= not(layer7_outputs(4735));
    layer8_outputs(386) <= (layer7_outputs(969)) and not (layer7_outputs(2472));
    layer8_outputs(387) <= layer7_outputs(5064);
    layer8_outputs(388) <= not(layer7_outputs(1877));
    layer8_outputs(389) <= layer7_outputs(619);
    layer8_outputs(390) <= not((layer7_outputs(4250)) and (layer7_outputs(1150)));
    layer8_outputs(391) <= not(layer7_outputs(941)) or (layer7_outputs(1441));
    layer8_outputs(392) <= (layer7_outputs(4518)) or (layer7_outputs(872));
    layer8_outputs(393) <= (layer7_outputs(4303)) xor (layer7_outputs(4287));
    layer8_outputs(394) <= (layer7_outputs(3715)) and (layer7_outputs(4829));
    layer8_outputs(395) <= not(layer7_outputs(755)) or (layer7_outputs(2902));
    layer8_outputs(396) <= (layer7_outputs(3412)) and not (layer7_outputs(4836));
    layer8_outputs(397) <= layer7_outputs(1762);
    layer8_outputs(398) <= not((layer7_outputs(4746)) xor (layer7_outputs(677)));
    layer8_outputs(399) <= layer7_outputs(449);
    layer8_outputs(400) <= not((layer7_outputs(1391)) or (layer7_outputs(3726)));
    layer8_outputs(401) <= not((layer7_outputs(4669)) xor (layer7_outputs(2862)));
    layer8_outputs(402) <= layer7_outputs(4998);
    layer8_outputs(403) <= not((layer7_outputs(876)) or (layer7_outputs(809)));
    layer8_outputs(404) <= (layer7_outputs(1133)) xor (layer7_outputs(4984));
    layer8_outputs(405) <= (layer7_outputs(5018)) or (layer7_outputs(430));
    layer8_outputs(406) <= not(layer7_outputs(2365));
    layer8_outputs(407) <= not(layer7_outputs(165));
    layer8_outputs(408) <= not(layer7_outputs(1234));
    layer8_outputs(409) <= not(layer7_outputs(2089));
    layer8_outputs(410) <= not(layer7_outputs(2088));
    layer8_outputs(411) <= layer7_outputs(563);
    layer8_outputs(412) <= layer7_outputs(5118);
    layer8_outputs(413) <= (layer7_outputs(1826)) xor (layer7_outputs(4372));
    layer8_outputs(414) <= (layer7_outputs(2877)) or (layer7_outputs(1113));
    layer8_outputs(415) <= (layer7_outputs(96)) and not (layer7_outputs(77));
    layer8_outputs(416) <= layer7_outputs(3496);
    layer8_outputs(417) <= (layer7_outputs(4119)) xor (layer7_outputs(4306));
    layer8_outputs(418) <= layer7_outputs(2778);
    layer8_outputs(419) <= not(layer7_outputs(4013));
    layer8_outputs(420) <= layer7_outputs(2672);
    layer8_outputs(421) <= layer7_outputs(4058);
    layer8_outputs(422) <= not((layer7_outputs(2947)) xor (layer7_outputs(3615)));
    layer8_outputs(423) <= layer7_outputs(1838);
    layer8_outputs(424) <= (layer7_outputs(3440)) and (layer7_outputs(3195));
    layer8_outputs(425) <= layer7_outputs(2945);
    layer8_outputs(426) <= layer7_outputs(976);
    layer8_outputs(427) <= (layer7_outputs(2204)) or (layer7_outputs(1994));
    layer8_outputs(428) <= layer7_outputs(1881);
    layer8_outputs(429) <= (layer7_outputs(461)) xor (layer7_outputs(1618));
    layer8_outputs(430) <= layer7_outputs(4633);
    layer8_outputs(431) <= (layer7_outputs(154)) and not (layer7_outputs(2637));
    layer8_outputs(432) <= not(layer7_outputs(3717));
    layer8_outputs(433) <= layer7_outputs(1471);
    layer8_outputs(434) <= layer7_outputs(1791);
    layer8_outputs(435) <= not((layer7_outputs(435)) xor (layer7_outputs(3898)));
    layer8_outputs(436) <= (layer7_outputs(3411)) xor (layer7_outputs(1459));
    layer8_outputs(437) <= layer7_outputs(1728);
    layer8_outputs(438) <= not(layer7_outputs(2255)) or (layer7_outputs(69));
    layer8_outputs(439) <= not(layer7_outputs(141)) or (layer7_outputs(2904));
    layer8_outputs(440) <= layer7_outputs(366);
    layer8_outputs(441) <= (layer7_outputs(2140)) xor (layer7_outputs(1916));
    layer8_outputs(442) <= not((layer7_outputs(4589)) xor (layer7_outputs(5067)));
    layer8_outputs(443) <= not((layer7_outputs(369)) xor (layer7_outputs(244)));
    layer8_outputs(444) <= (layer7_outputs(1432)) and not (layer7_outputs(1639));
    layer8_outputs(445) <= not(layer7_outputs(2258));
    layer8_outputs(446) <= not((layer7_outputs(1089)) or (layer7_outputs(4782)));
    layer8_outputs(447) <= not(layer7_outputs(4740));
    layer8_outputs(448) <= (layer7_outputs(4754)) and (layer7_outputs(4966));
    layer8_outputs(449) <= (layer7_outputs(4665)) and not (layer7_outputs(1212));
    layer8_outputs(450) <= layer7_outputs(1188);
    layer8_outputs(451) <= not((layer7_outputs(3691)) xor (layer7_outputs(50)));
    layer8_outputs(452) <= layer7_outputs(3625);
    layer8_outputs(453) <= (layer7_outputs(4069)) xor (layer7_outputs(4536));
    layer8_outputs(454) <= not((layer7_outputs(1521)) or (layer7_outputs(441)));
    layer8_outputs(455) <= (layer7_outputs(4457)) and not (layer7_outputs(1969));
    layer8_outputs(456) <= layer7_outputs(2592);
    layer8_outputs(457) <= not((layer7_outputs(3669)) xor (layer7_outputs(3013)));
    layer8_outputs(458) <= not(layer7_outputs(1629)) or (layer7_outputs(3840));
    layer8_outputs(459) <= (layer7_outputs(3830)) and (layer7_outputs(4889));
    layer8_outputs(460) <= (layer7_outputs(273)) xor (layer7_outputs(4381));
    layer8_outputs(461) <= not(layer7_outputs(4784)) or (layer7_outputs(3075));
    layer8_outputs(462) <= not(layer7_outputs(4527));
    layer8_outputs(463) <= not(layer7_outputs(2316));
    layer8_outputs(464) <= not(layer7_outputs(4583));
    layer8_outputs(465) <= not((layer7_outputs(1062)) xor (layer7_outputs(4358)));
    layer8_outputs(466) <= not(layer7_outputs(3721));
    layer8_outputs(467) <= not(layer7_outputs(764));
    layer8_outputs(468) <= (layer7_outputs(661)) xor (layer7_outputs(2910));
    layer8_outputs(469) <= layer7_outputs(1563);
    layer8_outputs(470) <= layer7_outputs(2519);
    layer8_outputs(471) <= not(layer7_outputs(1153));
    layer8_outputs(472) <= layer7_outputs(1235);
    layer8_outputs(473) <= not(layer7_outputs(2881));
    layer8_outputs(474) <= layer7_outputs(4214);
    layer8_outputs(475) <= (layer7_outputs(1742)) and not (layer7_outputs(1758));
    layer8_outputs(476) <= layer7_outputs(327);
    layer8_outputs(477) <= not((layer7_outputs(4213)) xor (layer7_outputs(4080)));
    layer8_outputs(478) <= (layer7_outputs(3370)) and not (layer7_outputs(3544));
    layer8_outputs(479) <= '0';
    layer8_outputs(480) <= (layer7_outputs(175)) and (layer7_outputs(1684));
    layer8_outputs(481) <= not((layer7_outputs(4804)) xor (layer7_outputs(40)));
    layer8_outputs(482) <= (layer7_outputs(3553)) xor (layer7_outputs(3799));
    layer8_outputs(483) <= layer7_outputs(4673);
    layer8_outputs(484) <= not(layer7_outputs(2598)) or (layer7_outputs(3878));
    layer8_outputs(485) <= (layer7_outputs(4679)) and not (layer7_outputs(767));
    layer8_outputs(486) <= not((layer7_outputs(388)) xor (layer7_outputs(3149)));
    layer8_outputs(487) <= layer7_outputs(3657);
    layer8_outputs(488) <= (layer7_outputs(959)) and (layer7_outputs(2532));
    layer8_outputs(489) <= layer7_outputs(2919);
    layer8_outputs(490) <= not((layer7_outputs(97)) xor (layer7_outputs(62)));
    layer8_outputs(491) <= layer7_outputs(1782);
    layer8_outputs(492) <= not(layer7_outputs(1082)) or (layer7_outputs(1644));
    layer8_outputs(493) <= (layer7_outputs(385)) xor (layer7_outputs(1492));
    layer8_outputs(494) <= (layer7_outputs(3103)) xor (layer7_outputs(407));
    layer8_outputs(495) <= not(layer7_outputs(4900)) or (layer7_outputs(3640));
    layer8_outputs(496) <= (layer7_outputs(3329)) xor (layer7_outputs(1536));
    layer8_outputs(497) <= layer7_outputs(913);
    layer8_outputs(498) <= not(layer7_outputs(413));
    layer8_outputs(499) <= layer7_outputs(4415);
    layer8_outputs(500) <= (layer7_outputs(4763)) xor (layer7_outputs(5112));
    layer8_outputs(501) <= not(layer7_outputs(1640));
    layer8_outputs(502) <= (layer7_outputs(3910)) xor (layer7_outputs(487));
    layer8_outputs(503) <= layer7_outputs(3952);
    layer8_outputs(504) <= not(layer7_outputs(2212));
    layer8_outputs(505) <= not(layer7_outputs(2362)) or (layer7_outputs(1050));
    layer8_outputs(506) <= not(layer7_outputs(906));
    layer8_outputs(507) <= not((layer7_outputs(4439)) and (layer7_outputs(1899)));
    layer8_outputs(508) <= not(layer7_outputs(2728)) or (layer7_outputs(997));
    layer8_outputs(509) <= not(layer7_outputs(1699));
    layer8_outputs(510) <= not(layer7_outputs(2491)) or (layer7_outputs(1059));
    layer8_outputs(511) <= layer7_outputs(2330);
    layer8_outputs(512) <= layer7_outputs(2864);
    layer8_outputs(513) <= not((layer7_outputs(4090)) xor (layer7_outputs(4060)));
    layer8_outputs(514) <= (layer7_outputs(2121)) and not (layer7_outputs(254));
    layer8_outputs(515) <= layer7_outputs(1041);
    layer8_outputs(516) <= not(layer7_outputs(4833));
    layer8_outputs(517) <= not((layer7_outputs(2980)) xor (layer7_outputs(3997)));
    layer8_outputs(518) <= (layer7_outputs(4066)) xor (layer7_outputs(329));
    layer8_outputs(519) <= not(layer7_outputs(2050)) or (layer7_outputs(4722));
    layer8_outputs(520) <= (layer7_outputs(4328)) and not (layer7_outputs(3427));
    layer8_outputs(521) <= layer7_outputs(4318);
    layer8_outputs(522) <= (layer7_outputs(1673)) and (layer7_outputs(3239));
    layer8_outputs(523) <= layer7_outputs(680);
    layer8_outputs(524) <= not((layer7_outputs(3199)) and (layer7_outputs(4053)));
    layer8_outputs(525) <= not((layer7_outputs(2059)) xor (layer7_outputs(462)));
    layer8_outputs(526) <= not((layer7_outputs(4505)) xor (layer7_outputs(3465)));
    layer8_outputs(527) <= not(layer7_outputs(695));
    layer8_outputs(528) <= not(layer7_outputs(3692)) or (layer7_outputs(2850));
    layer8_outputs(529) <= not((layer7_outputs(2587)) xor (layer7_outputs(4917)));
    layer8_outputs(530) <= layer7_outputs(305);
    layer8_outputs(531) <= layer7_outputs(2145);
    layer8_outputs(532) <= not(layer7_outputs(3251));
    layer8_outputs(533) <= not((layer7_outputs(1613)) or (layer7_outputs(2061)));
    layer8_outputs(534) <= not((layer7_outputs(2425)) xor (layer7_outputs(401)));
    layer8_outputs(535) <= not(layer7_outputs(3819));
    layer8_outputs(536) <= not(layer7_outputs(1438));
    layer8_outputs(537) <= (layer7_outputs(46)) or (layer7_outputs(3135));
    layer8_outputs(538) <= layer7_outputs(2823);
    layer8_outputs(539) <= (layer7_outputs(1497)) xor (layer7_outputs(4067));
    layer8_outputs(540) <= not(layer7_outputs(1741));
    layer8_outputs(541) <= layer7_outputs(4688);
    layer8_outputs(542) <= not((layer7_outputs(1600)) xor (layer7_outputs(1909)));
    layer8_outputs(543) <= layer7_outputs(3652);
    layer8_outputs(544) <= not((layer7_outputs(577)) or (layer7_outputs(4131)));
    layer8_outputs(545) <= (layer7_outputs(2713)) and not (layer7_outputs(3153));
    layer8_outputs(546) <= not(layer7_outputs(3027));
    layer8_outputs(547) <= layer7_outputs(4361);
    layer8_outputs(548) <= not(layer7_outputs(4252)) or (layer7_outputs(2161));
    layer8_outputs(549) <= (layer7_outputs(3694)) or (layer7_outputs(4991));
    layer8_outputs(550) <= not(layer7_outputs(4651));
    layer8_outputs(551) <= not(layer7_outputs(528)) or (layer7_outputs(4059));
    layer8_outputs(552) <= not(layer7_outputs(3560)) or (layer7_outputs(4543));
    layer8_outputs(553) <= not(layer7_outputs(1818));
    layer8_outputs(554) <= (layer7_outputs(1769)) and not (layer7_outputs(560));
    layer8_outputs(555) <= not((layer7_outputs(2210)) xor (layer7_outputs(2692)));
    layer8_outputs(556) <= not(layer7_outputs(428));
    layer8_outputs(557) <= layer7_outputs(3116);
    layer8_outputs(558) <= not(layer7_outputs(1646)) or (layer7_outputs(1572));
    layer8_outputs(559) <= not(layer7_outputs(4877));
    layer8_outputs(560) <= (layer7_outputs(3616)) xor (layer7_outputs(1040));
    layer8_outputs(561) <= not((layer7_outputs(4599)) xor (layer7_outputs(947)));
    layer8_outputs(562) <= layer7_outputs(65);
    layer8_outputs(563) <= not(layer7_outputs(1146));
    layer8_outputs(564) <= not(layer7_outputs(4325));
    layer8_outputs(565) <= layer7_outputs(2722);
    layer8_outputs(566) <= (layer7_outputs(2247)) xor (layer7_outputs(418));
    layer8_outputs(567) <= not(layer7_outputs(3737));
    layer8_outputs(568) <= layer7_outputs(2815);
    layer8_outputs(569) <= not(layer7_outputs(303));
    layer8_outputs(570) <= not(layer7_outputs(1532));
    layer8_outputs(571) <= layer7_outputs(4217);
    layer8_outputs(572) <= layer7_outputs(1539);
    layer8_outputs(573) <= layer7_outputs(1470);
    layer8_outputs(574) <= (layer7_outputs(2244)) and not (layer7_outputs(4779));
    layer8_outputs(575) <= not(layer7_outputs(2336));
    layer8_outputs(576) <= not(layer7_outputs(2186));
    layer8_outputs(577) <= not(layer7_outputs(3057));
    layer8_outputs(578) <= (layer7_outputs(4930)) or (layer7_outputs(4108));
    layer8_outputs(579) <= (layer7_outputs(3917)) and (layer7_outputs(4861));
    layer8_outputs(580) <= (layer7_outputs(174)) and not (layer7_outputs(2449));
    layer8_outputs(581) <= '0';
    layer8_outputs(582) <= layer7_outputs(3566);
    layer8_outputs(583) <= not(layer7_outputs(1212));
    layer8_outputs(584) <= layer7_outputs(3037);
    layer8_outputs(585) <= '0';
    layer8_outputs(586) <= not(layer7_outputs(1531));
    layer8_outputs(587) <= not(layer7_outputs(4489));
    layer8_outputs(588) <= not(layer7_outputs(3530)) or (layer7_outputs(1367));
    layer8_outputs(589) <= layer7_outputs(3476);
    layer8_outputs(590) <= not(layer7_outputs(282));
    layer8_outputs(591) <= not((layer7_outputs(2610)) and (layer7_outputs(4103)));
    layer8_outputs(592) <= not(layer7_outputs(3921));
    layer8_outputs(593) <= (layer7_outputs(338)) xor (layer7_outputs(3223));
    layer8_outputs(594) <= not(layer7_outputs(4685));
    layer8_outputs(595) <= not(layer7_outputs(3896));
    layer8_outputs(596) <= layer7_outputs(1053);
    layer8_outputs(597) <= not(layer7_outputs(1241));
    layer8_outputs(598) <= layer7_outputs(1755);
    layer8_outputs(599) <= not((layer7_outputs(3664)) xor (layer7_outputs(4695)));
    layer8_outputs(600) <= (layer7_outputs(943)) xor (layer7_outputs(734));
    layer8_outputs(601) <= not((layer7_outputs(1564)) xor (layer7_outputs(2609)));
    layer8_outputs(602) <= not(layer7_outputs(4530));
    layer8_outputs(603) <= not(layer7_outputs(3526)) or (layer7_outputs(3298));
    layer8_outputs(604) <= not(layer7_outputs(497)) or (layer7_outputs(4170));
    layer8_outputs(605) <= layer7_outputs(1516);
    layer8_outputs(606) <= not(layer7_outputs(4356));
    layer8_outputs(607) <= not((layer7_outputs(3475)) or (layer7_outputs(3676)));
    layer8_outputs(608) <= (layer7_outputs(4905)) or (layer7_outputs(2907));
    layer8_outputs(609) <= not(layer7_outputs(3813)) or (layer7_outputs(2788));
    layer8_outputs(610) <= layer7_outputs(2702);
    layer8_outputs(611) <= layer7_outputs(1443);
    layer8_outputs(612) <= not((layer7_outputs(2458)) xor (layer7_outputs(2406)));
    layer8_outputs(613) <= layer7_outputs(2484);
    layer8_outputs(614) <= not(layer7_outputs(4333));
    layer8_outputs(615) <= (layer7_outputs(4879)) and (layer7_outputs(318));
    layer8_outputs(616) <= not(layer7_outputs(4392));
    layer8_outputs(617) <= '0';
    layer8_outputs(618) <= layer7_outputs(2689);
    layer8_outputs(619) <= (layer7_outputs(3062)) xor (layer7_outputs(1074));
    layer8_outputs(620) <= layer7_outputs(2519);
    layer8_outputs(621) <= (layer7_outputs(2231)) and not (layer7_outputs(4755));
    layer8_outputs(622) <= not((layer7_outputs(2893)) or (layer7_outputs(270)));
    layer8_outputs(623) <= not(layer7_outputs(2289));
    layer8_outputs(624) <= (layer7_outputs(4236)) and not (layer7_outputs(3750));
    layer8_outputs(625) <= not(layer7_outputs(3498));
    layer8_outputs(626) <= layer7_outputs(4234);
    layer8_outputs(627) <= (layer7_outputs(875)) xor (layer7_outputs(3433));
    layer8_outputs(628) <= layer7_outputs(1691);
    layer8_outputs(629) <= (layer7_outputs(2485)) xor (layer7_outputs(1235));
    layer8_outputs(630) <= (layer7_outputs(4914)) or (layer7_outputs(3325));
    layer8_outputs(631) <= (layer7_outputs(68)) and not (layer7_outputs(2486));
    layer8_outputs(632) <= layer7_outputs(1649);
    layer8_outputs(633) <= (layer7_outputs(416)) and not (layer7_outputs(597));
    layer8_outputs(634) <= layer7_outputs(1445);
    layer8_outputs(635) <= layer7_outputs(3979);
    layer8_outputs(636) <= (layer7_outputs(4789)) xor (layer7_outputs(861));
    layer8_outputs(637) <= (layer7_outputs(1565)) and (layer7_outputs(456));
    layer8_outputs(638) <= not(layer7_outputs(1356));
    layer8_outputs(639) <= not((layer7_outputs(806)) and (layer7_outputs(486)));
    layer8_outputs(640) <= (layer7_outputs(3215)) xor (layer7_outputs(4762));
    layer8_outputs(641) <= layer7_outputs(5111);
    layer8_outputs(642) <= layer7_outputs(4246);
    layer8_outputs(643) <= layer7_outputs(3654);
    layer8_outputs(644) <= not((layer7_outputs(1750)) xor (layer7_outputs(5069)));
    layer8_outputs(645) <= not((layer7_outputs(1507)) or (layer7_outputs(231)));
    layer8_outputs(646) <= not(layer7_outputs(3896));
    layer8_outputs(647) <= layer7_outputs(4928);
    layer8_outputs(648) <= not(layer7_outputs(1454));
    layer8_outputs(649) <= not(layer7_outputs(4700));
    layer8_outputs(650) <= (layer7_outputs(705)) xor (layer7_outputs(627));
    layer8_outputs(651) <= not((layer7_outputs(2572)) xor (layer7_outputs(2648)));
    layer8_outputs(652) <= not(layer7_outputs(1337)) or (layer7_outputs(4993));
    layer8_outputs(653) <= '0';
    layer8_outputs(654) <= not((layer7_outputs(75)) and (layer7_outputs(171)));
    layer8_outputs(655) <= not(layer7_outputs(953));
    layer8_outputs(656) <= (layer7_outputs(2553)) and not (layer7_outputs(1014));
    layer8_outputs(657) <= layer7_outputs(4721);
    layer8_outputs(658) <= layer7_outputs(4555);
    layer8_outputs(659) <= '0';
    layer8_outputs(660) <= not(layer7_outputs(835));
    layer8_outputs(661) <= (layer7_outputs(4822)) and (layer7_outputs(4591));
    layer8_outputs(662) <= not((layer7_outputs(3970)) xor (layer7_outputs(3658)));
    layer8_outputs(663) <= layer7_outputs(908);
    layer8_outputs(664) <= not(layer7_outputs(4550));
    layer8_outputs(665) <= layer7_outputs(1076);
    layer8_outputs(666) <= layer7_outputs(1811);
    layer8_outputs(667) <= layer7_outputs(10);
    layer8_outputs(668) <= not(layer7_outputs(4963));
    layer8_outputs(669) <= not((layer7_outputs(3181)) xor (layer7_outputs(4579)));
    layer8_outputs(670) <= layer7_outputs(366);
    layer8_outputs(671) <= not(layer7_outputs(33)) or (layer7_outputs(637));
    layer8_outputs(672) <= not((layer7_outputs(453)) xor (layer7_outputs(2298)));
    layer8_outputs(673) <= not((layer7_outputs(3627)) xor (layer7_outputs(3084)));
    layer8_outputs(674) <= (layer7_outputs(1926)) or (layer7_outputs(4190));
    layer8_outputs(675) <= not(layer7_outputs(1001));
    layer8_outputs(676) <= '1';
    layer8_outputs(677) <= layer7_outputs(1460);
    layer8_outputs(678) <= not(layer7_outputs(4493));
    layer8_outputs(679) <= (layer7_outputs(3855)) or (layer7_outputs(1353));
    layer8_outputs(680) <= not(layer7_outputs(3992));
    layer8_outputs(681) <= not(layer7_outputs(5080));
    layer8_outputs(682) <= (layer7_outputs(3440)) and (layer7_outputs(1027));
    layer8_outputs(683) <= not(layer7_outputs(2045));
    layer8_outputs(684) <= not((layer7_outputs(100)) xor (layer7_outputs(304)));
    layer8_outputs(685) <= layer7_outputs(119);
    layer8_outputs(686) <= (layer7_outputs(4414)) and not (layer7_outputs(486));
    layer8_outputs(687) <= not(layer7_outputs(451));
    layer8_outputs(688) <= layer7_outputs(2223);
    layer8_outputs(689) <= not(layer7_outputs(3893)) or (layer7_outputs(2675));
    layer8_outputs(690) <= not(layer7_outputs(3557));
    layer8_outputs(691) <= (layer7_outputs(1211)) and (layer7_outputs(3226));
    layer8_outputs(692) <= not(layer7_outputs(2473));
    layer8_outputs(693) <= layer7_outputs(110);
    layer8_outputs(694) <= '0';
    layer8_outputs(695) <= layer7_outputs(2224);
    layer8_outputs(696) <= not(layer7_outputs(1963)) or (layer7_outputs(1406));
    layer8_outputs(697) <= layer7_outputs(64);
    layer8_outputs(698) <= not((layer7_outputs(3438)) xor (layer7_outputs(4835)));
    layer8_outputs(699) <= not((layer7_outputs(4597)) xor (layer7_outputs(2925)));
    layer8_outputs(700) <= layer7_outputs(1126);
    layer8_outputs(701) <= (layer7_outputs(467)) xor (layer7_outputs(3222));
    layer8_outputs(702) <= not(layer7_outputs(3827)) or (layer7_outputs(554));
    layer8_outputs(703) <= not((layer7_outputs(2610)) xor (layer7_outputs(4096)));
    layer8_outputs(704) <= not((layer7_outputs(3850)) xor (layer7_outputs(47)));
    layer8_outputs(705) <= not(layer7_outputs(2740));
    layer8_outputs(706) <= not((layer7_outputs(2087)) xor (layer7_outputs(560)));
    layer8_outputs(707) <= not(layer7_outputs(3889));
    layer8_outputs(708) <= not(layer7_outputs(614)) or (layer7_outputs(3847));
    layer8_outputs(709) <= (layer7_outputs(3650)) xor (layer7_outputs(2604));
    layer8_outputs(710) <= layer7_outputs(4488);
    layer8_outputs(711) <= not(layer7_outputs(3146));
    layer8_outputs(712) <= not(layer7_outputs(506));
    layer8_outputs(713) <= not(layer7_outputs(5027)) or (layer7_outputs(2143));
    layer8_outputs(714) <= (layer7_outputs(4095)) and not (layer7_outputs(4939));
    layer8_outputs(715) <= not(layer7_outputs(4002));
    layer8_outputs(716) <= '1';
    layer8_outputs(717) <= not(layer7_outputs(1228));
    layer8_outputs(718) <= not((layer7_outputs(2346)) and (layer7_outputs(1800)));
    layer8_outputs(719) <= layer7_outputs(4529);
    layer8_outputs(720) <= '0';
    layer8_outputs(721) <= (layer7_outputs(1813)) and not (layer7_outputs(633));
    layer8_outputs(722) <= not(layer7_outputs(107)) or (layer7_outputs(2522));
    layer8_outputs(723) <= not((layer7_outputs(4432)) xor (layer7_outputs(2822)));
    layer8_outputs(724) <= not((layer7_outputs(2666)) xor (layer7_outputs(2588)));
    layer8_outputs(725) <= not(layer7_outputs(1377));
    layer8_outputs(726) <= '1';
    layer8_outputs(727) <= not(layer7_outputs(1190)) or (layer7_outputs(1096));
    layer8_outputs(728) <= layer7_outputs(2999);
    layer8_outputs(729) <= layer7_outputs(4883);
    layer8_outputs(730) <= layer7_outputs(3061);
    layer8_outputs(731) <= not(layer7_outputs(530));
    layer8_outputs(732) <= not(layer7_outputs(3107));
    layer8_outputs(733) <= not((layer7_outputs(4138)) and (layer7_outputs(1682)));
    layer8_outputs(734) <= layer7_outputs(1652);
    layer8_outputs(735) <= layer7_outputs(4094);
    layer8_outputs(736) <= not(layer7_outputs(3241));
    layer8_outputs(737) <= layer7_outputs(689);
    layer8_outputs(738) <= not(layer7_outputs(4969)) or (layer7_outputs(4730));
    layer8_outputs(739) <= (layer7_outputs(4227)) and (layer7_outputs(4870));
    layer8_outputs(740) <= (layer7_outputs(2459)) and not (layer7_outputs(1036));
    layer8_outputs(741) <= not((layer7_outputs(3613)) and (layer7_outputs(2170)));
    layer8_outputs(742) <= not(layer7_outputs(1904));
    layer8_outputs(743) <= not((layer7_outputs(408)) xor (layer7_outputs(475)));
    layer8_outputs(744) <= not(layer7_outputs(3569));
    layer8_outputs(745) <= not(layer7_outputs(4038));
    layer8_outputs(746) <= layer7_outputs(1073);
    layer8_outputs(747) <= '0';
    layer8_outputs(748) <= (layer7_outputs(2716)) and (layer7_outputs(2216));
    layer8_outputs(749) <= layer7_outputs(3991);
    layer8_outputs(750) <= not(layer7_outputs(4657)) or (layer7_outputs(1570));
    layer8_outputs(751) <= layer7_outputs(2843);
    layer8_outputs(752) <= not((layer7_outputs(3429)) and (layer7_outputs(1577)));
    layer8_outputs(753) <= (layer7_outputs(2398)) xor (layer7_outputs(56));
    layer8_outputs(754) <= not(layer7_outputs(708));
    layer8_outputs(755) <= not(layer7_outputs(4470)) or (layer7_outputs(1179));
    layer8_outputs(756) <= (layer7_outputs(3603)) and (layer7_outputs(2695));
    layer8_outputs(757) <= not(layer7_outputs(4525)) or (layer7_outputs(3965));
    layer8_outputs(758) <= not(layer7_outputs(1402));
    layer8_outputs(759) <= not((layer7_outputs(3706)) xor (layer7_outputs(2844)));
    layer8_outputs(760) <= not(layer7_outputs(3237));
    layer8_outputs(761) <= layer7_outputs(4298);
    layer8_outputs(762) <= layer7_outputs(3131);
    layer8_outputs(763) <= not(layer7_outputs(1019));
    layer8_outputs(764) <= not(layer7_outputs(4407)) or (layer7_outputs(95));
    layer8_outputs(765) <= not(layer7_outputs(1931));
    layer8_outputs(766) <= not(layer7_outputs(3770));
    layer8_outputs(767) <= not((layer7_outputs(1100)) xor (layer7_outputs(1022)));
    layer8_outputs(768) <= not(layer7_outputs(2434)) or (layer7_outputs(2500));
    layer8_outputs(769) <= not(layer7_outputs(906));
    layer8_outputs(770) <= layer7_outputs(3299);
    layer8_outputs(771) <= (layer7_outputs(2453)) and (layer7_outputs(90));
    layer8_outputs(772) <= (layer7_outputs(353)) xor (layer7_outputs(2047));
    layer8_outputs(773) <= not((layer7_outputs(2579)) xor (layer7_outputs(908)));
    layer8_outputs(774) <= not((layer7_outputs(2400)) xor (layer7_outputs(3331)));
    layer8_outputs(775) <= not(layer7_outputs(2077));
    layer8_outputs(776) <= not(layer7_outputs(3871));
    layer8_outputs(777) <= not(layer7_outputs(4479));
    layer8_outputs(778) <= layer7_outputs(1862);
    layer8_outputs(779) <= layer7_outputs(2399);
    layer8_outputs(780) <= not((layer7_outputs(1553)) xor (layer7_outputs(4159)));
    layer8_outputs(781) <= (layer7_outputs(580)) and not (layer7_outputs(4797));
    layer8_outputs(782) <= (layer7_outputs(443)) and not (layer7_outputs(4649));
    layer8_outputs(783) <= not((layer7_outputs(568)) xor (layer7_outputs(4512)));
    layer8_outputs(784) <= not((layer7_outputs(3555)) or (layer7_outputs(4852)));
    layer8_outputs(785) <= not((layer7_outputs(4386)) xor (layer7_outputs(3758)));
    layer8_outputs(786) <= not(layer7_outputs(586));
    layer8_outputs(787) <= (layer7_outputs(1708)) xor (layer7_outputs(4639));
    layer8_outputs(788) <= not(layer7_outputs(2307));
    layer8_outputs(789) <= layer7_outputs(824);
    layer8_outputs(790) <= layer7_outputs(4661);
    layer8_outputs(791) <= layer7_outputs(2220);
    layer8_outputs(792) <= not((layer7_outputs(1623)) xor (layer7_outputs(593)));
    layer8_outputs(793) <= not(layer7_outputs(4984));
    layer8_outputs(794) <= (layer7_outputs(1907)) and (layer7_outputs(6));
    layer8_outputs(795) <= (layer7_outputs(1081)) and not (layer7_outputs(3837));
    layer8_outputs(796) <= not(layer7_outputs(3619)) or (layer7_outputs(3334));
    layer8_outputs(797) <= not(layer7_outputs(3904));
    layer8_outputs(798) <= not(layer7_outputs(2581));
    layer8_outputs(799) <= not(layer7_outputs(1424));
    layer8_outputs(800) <= not(layer7_outputs(2699)) or (layer7_outputs(57));
    layer8_outputs(801) <= layer7_outputs(2138);
    layer8_outputs(802) <= layer7_outputs(1420);
    layer8_outputs(803) <= not((layer7_outputs(2850)) or (layer7_outputs(5011)));
    layer8_outputs(804) <= not((layer7_outputs(5042)) or (layer7_outputs(408)));
    layer8_outputs(805) <= not(layer7_outputs(1668)) or (layer7_outputs(1013));
    layer8_outputs(806) <= not(layer7_outputs(170));
    layer8_outputs(807) <= not((layer7_outputs(978)) xor (layer7_outputs(4736)));
    layer8_outputs(808) <= not(layer7_outputs(3477));
    layer8_outputs(809) <= not((layer7_outputs(3718)) xor (layer7_outputs(4409)));
    layer8_outputs(810) <= not(layer7_outputs(1190)) or (layer7_outputs(204));
    layer8_outputs(811) <= layer7_outputs(4453);
    layer8_outputs(812) <= not((layer7_outputs(2555)) xor (layer7_outputs(3834)));
    layer8_outputs(813) <= not(layer7_outputs(1703));
    layer8_outputs(814) <= (layer7_outputs(1882)) and (layer7_outputs(3627));
    layer8_outputs(815) <= not(layer7_outputs(5101));
    layer8_outputs(816) <= not(layer7_outputs(3795));
    layer8_outputs(817) <= (layer7_outputs(3212)) or (layer7_outputs(1703));
    layer8_outputs(818) <= (layer7_outputs(3745)) and (layer7_outputs(909));
    layer8_outputs(819) <= layer7_outputs(4106);
    layer8_outputs(820) <= (layer7_outputs(4902)) and (layer7_outputs(4436));
    layer8_outputs(821) <= not((layer7_outputs(999)) xor (layer7_outputs(3505)));
    layer8_outputs(822) <= (layer7_outputs(3301)) xor (layer7_outputs(4243));
    layer8_outputs(823) <= layer7_outputs(2395);
    layer8_outputs(824) <= not((layer7_outputs(1477)) xor (layer7_outputs(5015)));
    layer8_outputs(825) <= layer7_outputs(887);
    layer8_outputs(826) <= layer7_outputs(3965);
    layer8_outputs(827) <= layer7_outputs(3129);
    layer8_outputs(828) <= not((layer7_outputs(1386)) and (layer7_outputs(4542)));
    layer8_outputs(829) <= layer7_outputs(3777);
    layer8_outputs(830) <= not((layer7_outputs(1677)) or (layer7_outputs(2155)));
    layer8_outputs(831) <= not(layer7_outputs(1770));
    layer8_outputs(832) <= not(layer7_outputs(3299));
    layer8_outputs(833) <= not(layer7_outputs(1633)) or (layer7_outputs(634));
    layer8_outputs(834) <= not(layer7_outputs(4458));
    layer8_outputs(835) <= (layer7_outputs(1943)) and not (layer7_outputs(2357));
    layer8_outputs(836) <= not(layer7_outputs(3529));
    layer8_outputs(837) <= layer7_outputs(4427);
    layer8_outputs(838) <= (layer7_outputs(4584)) or (layer7_outputs(481));
    layer8_outputs(839) <= not(layer7_outputs(2034));
    layer8_outputs(840) <= layer7_outputs(234);
    layer8_outputs(841) <= not(layer7_outputs(2340));
    layer8_outputs(842) <= layer7_outputs(890);
    layer8_outputs(843) <= not(layer7_outputs(4182));
    layer8_outputs(844) <= not(layer7_outputs(1582));
    layer8_outputs(845) <= not(layer7_outputs(1870));
    layer8_outputs(846) <= not(layer7_outputs(227));
    layer8_outputs(847) <= not(layer7_outputs(3963));
    layer8_outputs(848) <= not((layer7_outputs(1665)) and (layer7_outputs(363)));
    layer8_outputs(849) <= not(layer7_outputs(5083));
    layer8_outputs(850) <= (layer7_outputs(2356)) and not (layer7_outputs(4594));
    layer8_outputs(851) <= (layer7_outputs(1517)) xor (layer7_outputs(1798));
    layer8_outputs(852) <= not(layer7_outputs(1067));
    layer8_outputs(853) <= not((layer7_outputs(4840)) xor (layer7_outputs(4022)));
    layer8_outputs(854) <= not((layer7_outputs(4447)) xor (layer7_outputs(4580)));
    layer8_outputs(855) <= not(layer7_outputs(1436));
    layer8_outputs(856) <= not(layer7_outputs(2549));
    layer8_outputs(857) <= not((layer7_outputs(1164)) or (layer7_outputs(2435)));
    layer8_outputs(858) <= not(layer7_outputs(1556));
    layer8_outputs(859) <= not(layer7_outputs(2229)) or (layer7_outputs(4289));
    layer8_outputs(860) <= layer7_outputs(1695);
    layer8_outputs(861) <= layer7_outputs(641);
    layer8_outputs(862) <= layer7_outputs(3789);
    layer8_outputs(863) <= not(layer7_outputs(1343));
    layer8_outputs(864) <= (layer7_outputs(3381)) xor (layer7_outputs(4031));
    layer8_outputs(865) <= layer7_outputs(1851);
    layer8_outputs(866) <= (layer7_outputs(3849)) and not (layer7_outputs(577));
    layer8_outputs(867) <= (layer7_outputs(3099)) xor (layer7_outputs(4383));
    layer8_outputs(868) <= (layer7_outputs(1092)) xor (layer7_outputs(1292));
    layer8_outputs(869) <= layer7_outputs(4939);
    layer8_outputs(870) <= (layer7_outputs(1767)) and not (layer7_outputs(3760));
    layer8_outputs(871) <= not(layer7_outputs(4632)) or (layer7_outputs(1760));
    layer8_outputs(872) <= not(layer7_outputs(4438));
    layer8_outputs(873) <= (layer7_outputs(4046)) and (layer7_outputs(3558));
    layer8_outputs(874) <= layer7_outputs(498);
    layer8_outputs(875) <= not(layer7_outputs(3922)) or (layer7_outputs(1119));
    layer8_outputs(876) <= not(layer7_outputs(124)) or (layer7_outputs(3600));
    layer8_outputs(877) <= layer7_outputs(4381);
    layer8_outputs(878) <= not((layer7_outputs(18)) or (layer7_outputs(3413)));
    layer8_outputs(879) <= not(layer7_outputs(5113));
    layer8_outputs(880) <= not(layer7_outputs(3731));
    layer8_outputs(881) <= not(layer7_outputs(4509));
    layer8_outputs(882) <= not(layer7_outputs(865));
    layer8_outputs(883) <= (layer7_outputs(3431)) xor (layer7_outputs(4977));
    layer8_outputs(884) <= not(layer7_outputs(517));
    layer8_outputs(885) <= not(layer7_outputs(183));
    layer8_outputs(886) <= (layer7_outputs(1737)) and not (layer7_outputs(2668));
    layer8_outputs(887) <= (layer7_outputs(1240)) and not (layer7_outputs(711));
    layer8_outputs(888) <= not(layer7_outputs(630));
    layer8_outputs(889) <= not(layer7_outputs(1346));
    layer8_outputs(890) <= (layer7_outputs(2410)) xor (layer7_outputs(703));
    layer8_outputs(891) <= not((layer7_outputs(2127)) and (layer7_outputs(540)));
    layer8_outputs(892) <= layer7_outputs(3824);
    layer8_outputs(893) <= '1';
    layer8_outputs(894) <= not((layer7_outputs(1323)) and (layer7_outputs(2793)));
    layer8_outputs(895) <= (layer7_outputs(4878)) xor (layer7_outputs(1500));
    layer8_outputs(896) <= (layer7_outputs(2233)) xor (layer7_outputs(1549));
    layer8_outputs(897) <= layer7_outputs(3710);
    layer8_outputs(898) <= not((layer7_outputs(4883)) xor (layer7_outputs(3212)));
    layer8_outputs(899) <= layer7_outputs(2685);
    layer8_outputs(900) <= not(layer7_outputs(670));
    layer8_outputs(901) <= (layer7_outputs(37)) and not (layer7_outputs(3978));
    layer8_outputs(902) <= not((layer7_outputs(3415)) xor (layer7_outputs(3009)));
    layer8_outputs(903) <= not(layer7_outputs(4098));
    layer8_outputs(904) <= layer7_outputs(4927);
    layer8_outputs(905) <= not(layer7_outputs(3989)) or (layer7_outputs(4891));
    layer8_outputs(906) <= (layer7_outputs(4663)) xor (layer7_outputs(4578));
    layer8_outputs(907) <= layer7_outputs(3671);
    layer8_outputs(908) <= not((layer7_outputs(1469)) and (layer7_outputs(4362)));
    layer8_outputs(909) <= not((layer7_outputs(4100)) and (layer7_outputs(307)));
    layer8_outputs(910) <= '0';
    layer8_outputs(911) <= not(layer7_outputs(4747)) or (layer7_outputs(4568));
    layer8_outputs(912) <= not(layer7_outputs(2052));
    layer8_outputs(913) <= not(layer7_outputs(544));
    layer8_outputs(914) <= not(layer7_outputs(719)) or (layer7_outputs(1080));
    layer8_outputs(915) <= not((layer7_outputs(4906)) xor (layer7_outputs(4926)));
    layer8_outputs(916) <= not(layer7_outputs(1819));
    layer8_outputs(917) <= not((layer7_outputs(1285)) and (layer7_outputs(3217)));
    layer8_outputs(918) <= layer7_outputs(3659);
    layer8_outputs(919) <= layer7_outputs(2628);
    layer8_outputs(920) <= (layer7_outputs(180)) and (layer7_outputs(1321));
    layer8_outputs(921) <= not(layer7_outputs(700));
    layer8_outputs(922) <= not(layer7_outputs(1201)) or (layer7_outputs(694));
    layer8_outputs(923) <= layer7_outputs(1485);
    layer8_outputs(924) <= (layer7_outputs(1477)) xor (layer7_outputs(1020));
    layer8_outputs(925) <= layer7_outputs(551);
    layer8_outputs(926) <= layer7_outputs(3588);
    layer8_outputs(927) <= layer7_outputs(1465);
    layer8_outputs(928) <= (layer7_outputs(2582)) and not (layer7_outputs(3267));
    layer8_outputs(929) <= not(layer7_outputs(3981));
    layer8_outputs(930) <= (layer7_outputs(1511)) xor (layer7_outputs(71));
    layer8_outputs(931) <= not(layer7_outputs(1911));
    layer8_outputs(932) <= (layer7_outputs(3336)) and not (layer7_outputs(2403));
    layer8_outputs(933) <= layer7_outputs(3683);
    layer8_outputs(934) <= (layer7_outputs(4529)) xor (layer7_outputs(4346));
    layer8_outputs(935) <= layer7_outputs(1780);
    layer8_outputs(936) <= not(layer7_outputs(2054));
    layer8_outputs(937) <= not(layer7_outputs(2093));
    layer8_outputs(938) <= not(layer7_outputs(1822));
    layer8_outputs(939) <= (layer7_outputs(412)) xor (layer7_outputs(4488));
    layer8_outputs(940) <= not(layer7_outputs(2418));
    layer8_outputs(941) <= layer7_outputs(4354);
    layer8_outputs(942) <= layer7_outputs(4941);
    layer8_outputs(943) <= not(layer7_outputs(583)) or (layer7_outputs(4089));
    layer8_outputs(944) <= '0';
    layer8_outputs(945) <= layer7_outputs(3054);
    layer8_outputs(946) <= layer7_outputs(3665);
    layer8_outputs(947) <= (layer7_outputs(4481)) xor (layer7_outputs(876));
    layer8_outputs(948) <= not(layer7_outputs(1411)) or (layer7_outputs(1551));
    layer8_outputs(949) <= not((layer7_outputs(2307)) or (layer7_outputs(2796)));
    layer8_outputs(950) <= not((layer7_outputs(4540)) or (layer7_outputs(3562)));
    layer8_outputs(951) <= layer7_outputs(3386);
    layer8_outputs(952) <= (layer7_outputs(477)) xor (layer7_outputs(5106));
    layer8_outputs(953) <= (layer7_outputs(664)) xor (layer7_outputs(284));
    layer8_outputs(954) <= (layer7_outputs(4176)) and (layer7_outputs(1882));
    layer8_outputs(955) <= (layer7_outputs(4076)) and not (layer7_outputs(112));
    layer8_outputs(956) <= layer7_outputs(1409);
    layer8_outputs(957) <= (layer7_outputs(1185)) xor (layer7_outputs(2920));
    layer8_outputs(958) <= not((layer7_outputs(1033)) xor (layer7_outputs(3020)));
    layer8_outputs(959) <= not((layer7_outputs(1413)) xor (layer7_outputs(1063)));
    layer8_outputs(960) <= not(layer7_outputs(2448));
    layer8_outputs(961) <= not(layer7_outputs(2707));
    layer8_outputs(962) <= not(layer7_outputs(2103));
    layer8_outputs(963) <= not(layer7_outputs(4897));
    layer8_outputs(964) <= layer7_outputs(4008);
    layer8_outputs(965) <= (layer7_outputs(5089)) xor (layer7_outputs(2463));
    layer8_outputs(966) <= not((layer7_outputs(1177)) xor (layer7_outputs(2287)));
    layer8_outputs(967) <= (layer7_outputs(53)) and (layer7_outputs(1655));
    layer8_outputs(968) <= layer7_outputs(2562);
    layer8_outputs(969) <= layer7_outputs(4109);
    layer8_outputs(970) <= layer7_outputs(2573);
    layer8_outputs(971) <= not(layer7_outputs(3982));
    layer8_outputs(972) <= (layer7_outputs(1858)) or (layer7_outputs(1825));
    layer8_outputs(973) <= not(layer7_outputs(1537));
    layer8_outputs(974) <= not((layer7_outputs(2189)) xor (layer7_outputs(640)));
    layer8_outputs(975) <= not(layer7_outputs(2447)) or (layer7_outputs(3786));
    layer8_outputs(976) <= (layer7_outputs(4841)) and (layer7_outputs(357));
    layer8_outputs(977) <= '0';
    layer8_outputs(978) <= layer7_outputs(3216);
    layer8_outputs(979) <= (layer7_outputs(2836)) xor (layer7_outputs(423));
    layer8_outputs(980) <= not(layer7_outputs(3936));
    layer8_outputs(981) <= not(layer7_outputs(2352)) or (layer7_outputs(5092));
    layer8_outputs(982) <= not(layer7_outputs(3797));
    layer8_outputs(983) <= (layer7_outputs(1709)) and not (layer7_outputs(3376));
    layer8_outputs(984) <= layer7_outputs(2119);
    layer8_outputs(985) <= not(layer7_outputs(4220));
    layer8_outputs(986) <= not(layer7_outputs(4330)) or (layer7_outputs(1502));
    layer8_outputs(987) <= not(layer7_outputs(3204));
    layer8_outputs(988) <= not((layer7_outputs(3504)) or (layer7_outputs(1555)));
    layer8_outputs(989) <= not((layer7_outputs(2930)) xor (layer7_outputs(444)));
    layer8_outputs(990) <= (layer7_outputs(3793)) xor (layer7_outputs(3639));
    layer8_outputs(991) <= layer7_outputs(4908);
    layer8_outputs(992) <= (layer7_outputs(3313)) and (layer7_outputs(4700));
    layer8_outputs(993) <= not(layer7_outputs(744)) or (layer7_outputs(2883));
    layer8_outputs(994) <= not(layer7_outputs(2214));
    layer8_outputs(995) <= (layer7_outputs(3203)) xor (layer7_outputs(1995));
    layer8_outputs(996) <= layer7_outputs(3565);
    layer8_outputs(997) <= not((layer7_outputs(4929)) xor (layer7_outputs(4981)));
    layer8_outputs(998) <= not(layer7_outputs(4997));
    layer8_outputs(999) <= layer7_outputs(590);
    layer8_outputs(1000) <= layer7_outputs(4469);
    layer8_outputs(1001) <= not((layer7_outputs(4132)) and (layer7_outputs(1069)));
    layer8_outputs(1002) <= not(layer7_outputs(4531)) or (layer7_outputs(3868));
    layer8_outputs(1003) <= (layer7_outputs(2411)) and not (layer7_outputs(3866));
    layer8_outputs(1004) <= layer7_outputs(2131);
    layer8_outputs(1005) <= layer7_outputs(521);
    layer8_outputs(1006) <= not((layer7_outputs(3186)) xor (layer7_outputs(4780)));
    layer8_outputs(1007) <= (layer7_outputs(541)) xor (layer7_outputs(2218));
    layer8_outputs(1008) <= not(layer7_outputs(248)) or (layer7_outputs(3937));
    layer8_outputs(1009) <= (layer7_outputs(1982)) xor (layer7_outputs(4124));
    layer8_outputs(1010) <= not(layer7_outputs(4010));
    layer8_outputs(1011) <= not((layer7_outputs(3464)) xor (layer7_outputs(4445)));
    layer8_outputs(1012) <= layer7_outputs(379);
    layer8_outputs(1013) <= layer7_outputs(1574);
    layer8_outputs(1014) <= not(layer7_outputs(4134));
    layer8_outputs(1015) <= (layer7_outputs(3378)) and not (layer7_outputs(618));
    layer8_outputs(1016) <= layer7_outputs(2966);
    layer8_outputs(1017) <= layer7_outputs(5005);
    layer8_outputs(1018) <= not((layer7_outputs(4172)) xor (layer7_outputs(1078)));
    layer8_outputs(1019) <= layer7_outputs(1057);
    layer8_outputs(1020) <= not(layer7_outputs(4121));
    layer8_outputs(1021) <= (layer7_outputs(858)) xor (layer7_outputs(2520));
    layer8_outputs(1022) <= not(layer7_outputs(3177));
    layer8_outputs(1023) <= (layer7_outputs(4113)) and not (layer7_outputs(3825));
    layer8_outputs(1024) <= (layer7_outputs(2112)) or (layer7_outputs(2136));
    layer8_outputs(1025) <= layer7_outputs(239);
    layer8_outputs(1026) <= layer7_outputs(2742);
    layer8_outputs(1027) <= (layer7_outputs(3154)) xor (layer7_outputs(122));
    layer8_outputs(1028) <= layer7_outputs(2755);
    layer8_outputs(1029) <= not((layer7_outputs(1902)) xor (layer7_outputs(375)));
    layer8_outputs(1030) <= layer7_outputs(2694);
    layer8_outputs(1031) <= not((layer7_outputs(4706)) or (layer7_outputs(1245)));
    layer8_outputs(1032) <= not(layer7_outputs(2737));
    layer8_outputs(1033) <= layer7_outputs(2081);
    layer8_outputs(1034) <= layer7_outputs(980);
    layer8_outputs(1035) <= layer7_outputs(3636);
    layer8_outputs(1036) <= (layer7_outputs(5012)) xor (layer7_outputs(1950));
    layer8_outputs(1037) <= (layer7_outputs(2953)) xor (layer7_outputs(4430));
    layer8_outputs(1038) <= layer7_outputs(93);
    layer8_outputs(1039) <= '0';
    layer8_outputs(1040) <= not((layer7_outputs(1581)) xor (layer7_outputs(4270)));
    layer8_outputs(1041) <= (layer7_outputs(1382)) and not (layer7_outputs(4464));
    layer8_outputs(1042) <= not(layer7_outputs(4776));
    layer8_outputs(1043) <= not(layer7_outputs(2679));
    layer8_outputs(1044) <= layer7_outputs(3506);
    layer8_outputs(1045) <= (layer7_outputs(3274)) or (layer7_outputs(4316));
    layer8_outputs(1046) <= layer7_outputs(966);
    layer8_outputs(1047) <= not((layer7_outputs(1711)) xor (layer7_outputs(4560)));
    layer8_outputs(1048) <= '0';
    layer8_outputs(1049) <= layer7_outputs(1192);
    layer8_outputs(1050) <= not((layer7_outputs(2342)) and (layer7_outputs(1710)));
    layer8_outputs(1051) <= not(layer7_outputs(1809));
    layer8_outputs(1052) <= not(layer7_outputs(1202));
    layer8_outputs(1053) <= (layer7_outputs(707)) and (layer7_outputs(4943));
    layer8_outputs(1054) <= (layer7_outputs(3156)) and not (layer7_outputs(715));
    layer8_outputs(1055) <= layer7_outputs(3502);
    layer8_outputs(1056) <= layer7_outputs(4869);
    layer8_outputs(1057) <= not(layer7_outputs(2245));
    layer8_outputs(1058) <= not(layer7_outputs(414));
    layer8_outputs(1059) <= (layer7_outputs(1720)) or (layer7_outputs(182));
    layer8_outputs(1060) <= (layer7_outputs(743)) xor (layer7_outputs(2369));
    layer8_outputs(1061) <= (layer7_outputs(4687)) xor (layer7_outputs(4127));
    layer8_outputs(1062) <= layer7_outputs(2664);
    layer8_outputs(1063) <= not(layer7_outputs(4209));
    layer8_outputs(1064) <= not(layer7_outputs(149));
    layer8_outputs(1065) <= layer7_outputs(4638);
    layer8_outputs(1066) <= layer7_outputs(84);
    layer8_outputs(1067) <= not((layer7_outputs(2536)) or (layer7_outputs(2531)));
    layer8_outputs(1068) <= not(layer7_outputs(2226));
    layer8_outputs(1069) <= not(layer7_outputs(4517));
    layer8_outputs(1070) <= not(layer7_outputs(3147)) or (layer7_outputs(3287));
    layer8_outputs(1071) <= layer7_outputs(1134);
    layer8_outputs(1072) <= not((layer7_outputs(3309)) xor (layer7_outputs(524)));
    layer8_outputs(1073) <= (layer7_outputs(3118)) or (layer7_outputs(480));
    layer8_outputs(1074) <= layer7_outputs(2312);
    layer8_outputs(1075) <= not(layer7_outputs(1723)) or (layer7_outputs(1220));
    layer8_outputs(1076) <= not((layer7_outputs(4258)) xor (layer7_outputs(1917)));
    layer8_outputs(1077) <= layer7_outputs(2308);
    layer8_outputs(1078) <= not(layer7_outputs(3815));
    layer8_outputs(1079) <= layer7_outputs(254);
    layer8_outputs(1080) <= not(layer7_outputs(3332));
    layer8_outputs(1081) <= layer7_outputs(576);
    layer8_outputs(1082) <= '0';
    layer8_outputs(1083) <= layer7_outputs(4079);
    layer8_outputs(1084) <= layer7_outputs(5036);
    layer8_outputs(1085) <= (layer7_outputs(3907)) and not (layer7_outputs(1360));
    layer8_outputs(1086) <= layer7_outputs(3242);
    layer8_outputs(1087) <= layer7_outputs(4826);
    layer8_outputs(1088) <= (layer7_outputs(2643)) and not (layer7_outputs(1741));
    layer8_outputs(1089) <= (layer7_outputs(3330)) xor (layer7_outputs(4543));
    layer8_outputs(1090) <= not(layer7_outputs(3945)) or (layer7_outputs(1272));
    layer8_outputs(1091) <= not(layer7_outputs(1154));
    layer8_outputs(1092) <= not(layer7_outputs(4821));
    layer8_outputs(1093) <= not(layer7_outputs(4556));
    layer8_outputs(1094) <= not((layer7_outputs(4411)) xor (layer7_outputs(4576)));
    layer8_outputs(1095) <= (layer7_outputs(1953)) and not (layer7_outputs(3565));
    layer8_outputs(1096) <= not(layer7_outputs(4265));
    layer8_outputs(1097) <= layer7_outputs(753);
    layer8_outputs(1098) <= not(layer7_outputs(2527));
    layer8_outputs(1099) <= not(layer7_outputs(2156));
    layer8_outputs(1100) <= not(layer7_outputs(818)) or (layer7_outputs(2524));
    layer8_outputs(1101) <= not(layer7_outputs(3998)) or (layer7_outputs(3305));
    layer8_outputs(1102) <= not((layer7_outputs(648)) or (layer7_outputs(2967)));
    layer8_outputs(1103) <= not(layer7_outputs(1933));
    layer8_outputs(1104) <= not((layer7_outputs(4897)) xor (layer7_outputs(4852)));
    layer8_outputs(1105) <= not(layer7_outputs(2176));
    layer8_outputs(1106) <= not(layer7_outputs(4742));
    layer8_outputs(1107) <= not(layer7_outputs(4848)) or (layer7_outputs(4043));
    layer8_outputs(1108) <= not((layer7_outputs(1812)) or (layer7_outputs(2298)));
    layer8_outputs(1109) <= (layer7_outputs(3493)) xor (layer7_outputs(4872));
    layer8_outputs(1110) <= (layer7_outputs(1895)) or (layer7_outputs(4070));
    layer8_outputs(1111) <= layer7_outputs(1537);
    layer8_outputs(1112) <= (layer7_outputs(2121)) and not (layer7_outputs(3063));
    layer8_outputs(1113) <= not(layer7_outputs(1635)) or (layer7_outputs(4659));
    layer8_outputs(1114) <= layer7_outputs(5046);
    layer8_outputs(1115) <= not(layer7_outputs(4652));
    layer8_outputs(1116) <= not((layer7_outputs(1479)) xor (layer7_outputs(2892)));
    layer8_outputs(1117) <= (layer7_outputs(3490)) and not (layer7_outputs(3626));
    layer8_outputs(1118) <= not(layer7_outputs(1161)) or (layer7_outputs(582));
    layer8_outputs(1119) <= not(layer7_outputs(2887)) or (layer7_outputs(4496));
    layer8_outputs(1120) <= layer7_outputs(2055);
    layer8_outputs(1121) <= (layer7_outputs(900)) and not (layer7_outputs(2044));
    layer8_outputs(1122) <= not(layer7_outputs(3658));
    layer8_outputs(1123) <= (layer7_outputs(2997)) xor (layer7_outputs(1653));
    layer8_outputs(1124) <= (layer7_outputs(608)) xor (layer7_outputs(2285));
    layer8_outputs(1125) <= (layer7_outputs(2841)) xor (layer7_outputs(374));
    layer8_outputs(1126) <= (layer7_outputs(997)) xor (layer7_outputs(410));
    layer8_outputs(1127) <= layer7_outputs(237);
    layer8_outputs(1128) <= (layer7_outputs(3954)) xor (layer7_outputs(4042));
    layer8_outputs(1129) <= (layer7_outputs(2765)) xor (layer7_outputs(126));
    layer8_outputs(1130) <= not((layer7_outputs(1491)) xor (layer7_outputs(1831)));
    layer8_outputs(1131) <= layer7_outputs(1930);
    layer8_outputs(1132) <= not(layer7_outputs(1936));
    layer8_outputs(1133) <= not(layer7_outputs(3039));
    layer8_outputs(1134) <= not(layer7_outputs(357));
    layer8_outputs(1135) <= (layer7_outputs(2085)) xor (layer7_outputs(640));
    layer8_outputs(1136) <= not(layer7_outputs(4087));
    layer8_outputs(1137) <= not((layer7_outputs(1418)) xor (layer7_outputs(4147)));
    layer8_outputs(1138) <= not((layer7_outputs(4853)) xor (layer7_outputs(1393)));
    layer8_outputs(1139) <= layer7_outputs(2154);
    layer8_outputs(1140) <= layer7_outputs(3066);
    layer8_outputs(1141) <= layer7_outputs(2710);
    layer8_outputs(1142) <= (layer7_outputs(1972)) or (layer7_outputs(4096));
    layer8_outputs(1143) <= layer7_outputs(2900);
    layer8_outputs(1144) <= (layer7_outputs(2554)) and not (layer7_outputs(2641));
    layer8_outputs(1145) <= layer7_outputs(1250);
    layer8_outputs(1146) <= layer7_outputs(648);
    layer8_outputs(1147) <= (layer7_outputs(1122)) and not (layer7_outputs(4271));
    layer8_outputs(1148) <= not((layer7_outputs(1204)) xor (layer7_outputs(3042)));
    layer8_outputs(1149) <= not(layer7_outputs(3350));
    layer8_outputs(1150) <= layer7_outputs(23);
    layer8_outputs(1151) <= not(layer7_outputs(687));
    layer8_outputs(1152) <= (layer7_outputs(4175)) or (layer7_outputs(1976));
    layer8_outputs(1153) <= not((layer7_outputs(459)) or (layer7_outputs(109)));
    layer8_outputs(1154) <= not((layer7_outputs(3390)) xor (layer7_outputs(2028)));
    layer8_outputs(1155) <= not(layer7_outputs(1515)) or (layer7_outputs(2493));
    layer8_outputs(1156) <= not(layer7_outputs(955)) or (layer7_outputs(3372));
    layer8_outputs(1157) <= not(layer7_outputs(752));
    layer8_outputs(1158) <= not(layer7_outputs(2597));
    layer8_outputs(1159) <= layer7_outputs(2915);
    layer8_outputs(1160) <= not(layer7_outputs(3722));
    layer8_outputs(1161) <= layer7_outputs(927);
    layer8_outputs(1162) <= layer7_outputs(4565);
    layer8_outputs(1163) <= not(layer7_outputs(4924));
    layer8_outputs(1164) <= not((layer7_outputs(4095)) xor (layer7_outputs(3613)));
    layer8_outputs(1165) <= layer7_outputs(5118);
    layer8_outputs(1166) <= not(layer7_outputs(1389));
    layer8_outputs(1167) <= (layer7_outputs(1909)) and (layer7_outputs(1077));
    layer8_outputs(1168) <= layer7_outputs(57);
    layer8_outputs(1169) <= layer7_outputs(1548);
    layer8_outputs(1170) <= layer7_outputs(2945);
    layer8_outputs(1171) <= (layer7_outputs(1385)) and not (layer7_outputs(1306));
    layer8_outputs(1172) <= layer7_outputs(1910);
    layer8_outputs(1173) <= (layer7_outputs(2565)) and (layer7_outputs(5014));
    layer8_outputs(1174) <= not(layer7_outputs(4738)) or (layer7_outputs(4093));
    layer8_outputs(1175) <= (layer7_outputs(2359)) xor (layer7_outputs(299));
    layer8_outputs(1176) <= not((layer7_outputs(2081)) xor (layer7_outputs(5053)));
    layer8_outputs(1177) <= not(layer7_outputs(4914));
    layer8_outputs(1178) <= (layer7_outputs(2021)) and not (layer7_outputs(2451));
    layer8_outputs(1179) <= layer7_outputs(3407);
    layer8_outputs(1180) <= layer7_outputs(4146);
    layer8_outputs(1181) <= (layer7_outputs(4907)) and not (layer7_outputs(1759));
    layer8_outputs(1182) <= layer7_outputs(3261);
    layer8_outputs(1183) <= (layer7_outputs(3656)) xor (layer7_outputs(4029));
    layer8_outputs(1184) <= not((layer7_outputs(2043)) xor (layer7_outputs(728)));
    layer8_outputs(1185) <= not(layer7_outputs(2000));
    layer8_outputs(1186) <= not(layer7_outputs(2593)) or (layer7_outputs(2312));
    layer8_outputs(1187) <= layer7_outputs(1738);
    layer8_outputs(1188) <= not(layer7_outputs(4508));
    layer8_outputs(1189) <= layer7_outputs(4174);
    layer8_outputs(1190) <= (layer7_outputs(2554)) xor (layer7_outputs(2230));
    layer8_outputs(1191) <= (layer7_outputs(403)) or (layer7_outputs(265));
    layer8_outputs(1192) <= layer7_outputs(2995);
    layer8_outputs(1193) <= (layer7_outputs(1519)) or (layer7_outputs(4697));
    layer8_outputs(1194) <= not(layer7_outputs(3961));
    layer8_outputs(1195) <= not(layer7_outputs(2096));
    layer8_outputs(1196) <= (layer7_outputs(2115)) xor (layer7_outputs(3090));
    layer8_outputs(1197) <= layer7_outputs(1693);
    layer8_outputs(1198) <= not((layer7_outputs(3125)) xor (layer7_outputs(3044)));
    layer8_outputs(1199) <= (layer7_outputs(556)) xor (layer7_outputs(1151));
    layer8_outputs(1200) <= layer7_outputs(1431);
    layer8_outputs(1201) <= not(layer7_outputs(3449));
    layer8_outputs(1202) <= (layer7_outputs(3400)) and not (layer7_outputs(727));
    layer8_outputs(1203) <= layer7_outputs(2437);
    layer8_outputs(1204) <= (layer7_outputs(1594)) xor (layer7_outputs(2269));
    layer8_outputs(1205) <= not((layer7_outputs(1327)) xor (layer7_outputs(4908)));
    layer8_outputs(1206) <= not(layer7_outputs(1583));
    layer8_outputs(1207) <= not(layer7_outputs(3019));
    layer8_outputs(1208) <= (layer7_outputs(2303)) and not (layer7_outputs(1476));
    layer8_outputs(1209) <= layer7_outputs(4843);
    layer8_outputs(1210) <= (layer7_outputs(252)) xor (layer7_outputs(2109));
    layer8_outputs(1211) <= '0';
    layer8_outputs(1212) <= layer7_outputs(2205);
    layer8_outputs(1213) <= (layer7_outputs(162)) xor (layer7_outputs(2439));
    layer8_outputs(1214) <= layer7_outputs(1830);
    layer8_outputs(1215) <= not((layer7_outputs(934)) xor (layer7_outputs(3207)));
    layer8_outputs(1216) <= not((layer7_outputs(4822)) xor (layer7_outputs(14)));
    layer8_outputs(1217) <= layer7_outputs(2994);
    layer8_outputs(1218) <= not(layer7_outputs(2257));
    layer8_outputs(1219) <= layer7_outputs(4492);
    layer8_outputs(1220) <= not((layer7_outputs(2242)) xor (layer7_outputs(2503)));
    layer8_outputs(1221) <= (layer7_outputs(2526)) and not (layer7_outputs(4164));
    layer8_outputs(1222) <= (layer7_outputs(1353)) and (layer7_outputs(917));
    layer8_outputs(1223) <= layer7_outputs(4621);
    layer8_outputs(1224) <= (layer7_outputs(2674)) xor (layer7_outputs(2391));
    layer8_outputs(1225) <= not((layer7_outputs(1116)) xor (layer7_outputs(4641)));
    layer8_outputs(1226) <= (layer7_outputs(884)) and not (layer7_outputs(1092));
    layer8_outputs(1227) <= not(layer7_outputs(3698)) or (layer7_outputs(1113));
    layer8_outputs(1228) <= not((layer7_outputs(2310)) xor (layer7_outputs(2915)));
    layer8_outputs(1229) <= (layer7_outputs(3105)) and not (layer7_outputs(757));
    layer8_outputs(1230) <= not(layer7_outputs(4434));
    layer8_outputs(1231) <= '0';
    layer8_outputs(1232) <= layer7_outputs(1617);
    layer8_outputs(1233) <= (layer7_outputs(1213)) and (layer7_outputs(4460));
    layer8_outputs(1234) <= not((layer7_outputs(2234)) xor (layer7_outputs(2801)));
    layer8_outputs(1235) <= (layer7_outputs(2004)) xor (layer7_outputs(4552));
    layer8_outputs(1236) <= not(layer7_outputs(3903));
    layer8_outputs(1237) <= not((layer7_outputs(4582)) xor (layer7_outputs(1642)));
    layer8_outputs(1238) <= '0';
    layer8_outputs(1239) <= layer7_outputs(1164);
    layer8_outputs(1240) <= not(layer7_outputs(2738));
    layer8_outputs(1241) <= not((layer7_outputs(2976)) xor (layer7_outputs(2488)));
    layer8_outputs(1242) <= layer7_outputs(4923);
    layer8_outputs(1243) <= (layer7_outputs(483)) or (layer7_outputs(5026));
    layer8_outputs(1244) <= not(layer7_outputs(111));
    layer8_outputs(1245) <= (layer7_outputs(2180)) xor (layer7_outputs(3881));
    layer8_outputs(1246) <= (layer7_outputs(3884)) xor (layer7_outputs(2061));
    layer8_outputs(1247) <= '1';
    layer8_outputs(1248) <= (layer7_outputs(1338)) and not (layer7_outputs(3409));
    layer8_outputs(1249) <= not(layer7_outputs(2657)) or (layer7_outputs(2854));
    layer8_outputs(1250) <= not((layer7_outputs(3517)) xor (layer7_outputs(1490)));
    layer8_outputs(1251) <= not(layer7_outputs(1336));
    layer8_outputs(1252) <= (layer7_outputs(199)) xor (layer7_outputs(4912));
    layer8_outputs(1253) <= not((layer7_outputs(3127)) xor (layer7_outputs(1136)));
    layer8_outputs(1254) <= (layer7_outputs(1495)) xor (layer7_outputs(3437));
    layer8_outputs(1255) <= not(layer7_outputs(2194));
    layer8_outputs(1256) <= layer7_outputs(3258);
    layer8_outputs(1257) <= layer7_outputs(2513);
    layer8_outputs(1258) <= not((layer7_outputs(2281)) xor (layer7_outputs(3750)));
    layer8_outputs(1259) <= not(layer7_outputs(1434)) or (layer7_outputs(4607));
    layer8_outputs(1260) <= not((layer7_outputs(2819)) and (layer7_outputs(4126)));
    layer8_outputs(1261) <= layer7_outputs(683);
    layer8_outputs(1262) <= not(layer7_outputs(582));
    layer8_outputs(1263) <= layer7_outputs(977);
    layer8_outputs(1264) <= layer7_outputs(3951);
    layer8_outputs(1265) <= not((layer7_outputs(602)) xor (layer7_outputs(536)));
    layer8_outputs(1266) <= not(layer7_outputs(451));
    layer8_outputs(1267) <= (layer7_outputs(2293)) and not (layer7_outputs(4154));
    layer8_outputs(1268) <= not(layer7_outputs(3346));
    layer8_outputs(1269) <= not(layer7_outputs(2275));
    layer8_outputs(1270) <= not(layer7_outputs(4993));
    layer8_outputs(1271) <= not(layer7_outputs(431));
    layer8_outputs(1272) <= not((layer7_outputs(438)) xor (layer7_outputs(2791)));
    layer8_outputs(1273) <= layer7_outputs(1238);
    layer8_outputs(1274) <= (layer7_outputs(3277)) xor (layer7_outputs(762));
    layer8_outputs(1275) <= (layer7_outputs(216)) xor (layer7_outputs(2886));
    layer8_outputs(1276) <= (layer7_outputs(704)) and (layer7_outputs(679));
    layer8_outputs(1277) <= layer7_outputs(2798);
    layer8_outputs(1278) <= not((layer7_outputs(3950)) xor (layer7_outputs(5005)));
    layer8_outputs(1279) <= not(layer7_outputs(3139));
    layer8_outputs(1280) <= (layer7_outputs(330)) or (layer7_outputs(3052));
    layer8_outputs(1281) <= not(layer7_outputs(1499));
    layer8_outputs(1282) <= (layer7_outputs(2718)) xor (layer7_outputs(44));
    layer8_outputs(1283) <= not((layer7_outputs(3421)) xor (layer7_outputs(559)));
    layer8_outputs(1284) <= not(layer7_outputs(103));
    layer8_outputs(1285) <= layer7_outputs(2726);
    layer8_outputs(1286) <= (layer7_outputs(2258)) xor (layer7_outputs(605));
    layer8_outputs(1287) <= not((layer7_outputs(2466)) xor (layer7_outputs(191)));
    layer8_outputs(1288) <= (layer7_outputs(1306)) xor (layer7_outputs(2128));
    layer8_outputs(1289) <= not(layer7_outputs(236));
    layer8_outputs(1290) <= not(layer7_outputs(1816));
    layer8_outputs(1291) <= (layer7_outputs(2917)) xor (layer7_outputs(2476));
    layer8_outputs(1292) <= layer7_outputs(2710);
    layer8_outputs(1293) <= (layer7_outputs(948)) and not (layer7_outputs(889));
    layer8_outputs(1294) <= layer7_outputs(2734);
    layer8_outputs(1295) <= not(layer7_outputs(35));
    layer8_outputs(1296) <= not(layer7_outputs(4990)) or (layer7_outputs(3989));
    layer8_outputs(1297) <= not((layer7_outputs(490)) and (layer7_outputs(710)));
    layer8_outputs(1298) <= not(layer7_outputs(3002));
    layer8_outputs(1299) <= layer7_outputs(4783);
    layer8_outputs(1300) <= layer7_outputs(2691);
    layer8_outputs(1301) <= layer7_outputs(1644);
    layer8_outputs(1302) <= not(layer7_outputs(2873));
    layer8_outputs(1303) <= not(layer7_outputs(3544));
    layer8_outputs(1304) <= (layer7_outputs(1667)) xor (layer7_outputs(2956));
    layer8_outputs(1305) <= (layer7_outputs(4373)) xor (layer7_outputs(3841));
    layer8_outputs(1306) <= not(layer7_outputs(3532));
    layer8_outputs(1307) <= not((layer7_outputs(4197)) xor (layer7_outputs(1375)));
    layer8_outputs(1308) <= (layer7_outputs(562)) and (layer7_outputs(4553));
    layer8_outputs(1309) <= layer7_outputs(3355);
    layer8_outputs(1310) <= not(layer7_outputs(4541));
    layer8_outputs(1311) <= layer7_outputs(2550);
    layer8_outputs(1312) <= layer7_outputs(1392);
    layer8_outputs(1313) <= layer7_outputs(2942);
    layer8_outputs(1314) <= not((layer7_outputs(4867)) or (layer7_outputs(2746)));
    layer8_outputs(1315) <= (layer7_outputs(2655)) xor (layer7_outputs(4870));
    layer8_outputs(1316) <= layer7_outputs(4157);
    layer8_outputs(1317) <= (layer7_outputs(178)) xor (layer7_outputs(3500));
    layer8_outputs(1318) <= (layer7_outputs(1584)) xor (layer7_outputs(653));
    layer8_outputs(1319) <= layer7_outputs(4450);
    layer8_outputs(1320) <= not((layer7_outputs(5025)) xor (layer7_outputs(1411)));
    layer8_outputs(1321) <= layer7_outputs(4201);
    layer8_outputs(1322) <= layer7_outputs(3784);
    layer8_outputs(1323) <= layer7_outputs(2235);
    layer8_outputs(1324) <= not(layer7_outputs(3770));
    layer8_outputs(1325) <= layer7_outputs(2276);
    layer8_outputs(1326) <= (layer7_outputs(2263)) xor (layer7_outputs(1875));
    layer8_outputs(1327) <= layer7_outputs(3104);
    layer8_outputs(1328) <= layer7_outputs(4281);
    layer8_outputs(1329) <= not(layer7_outputs(1257));
    layer8_outputs(1330) <= (layer7_outputs(3719)) xor (layer7_outputs(121));
    layer8_outputs(1331) <= (layer7_outputs(1050)) and (layer7_outputs(3183));
    layer8_outputs(1332) <= not(layer7_outputs(2929));
    layer8_outputs(1333) <= (layer7_outputs(1111)) xor (layer7_outputs(3992));
    layer8_outputs(1334) <= layer7_outputs(3145);
    layer8_outputs(1335) <= not(layer7_outputs(924));
    layer8_outputs(1336) <= layer7_outputs(3783);
    layer8_outputs(1337) <= layer7_outputs(1117);
    layer8_outputs(1338) <= not(layer7_outputs(1789)) or (layer7_outputs(1038));
    layer8_outputs(1339) <= not(layer7_outputs(642));
    layer8_outputs(1340) <= not((layer7_outputs(952)) xor (layer7_outputs(167)));
    layer8_outputs(1341) <= not(layer7_outputs(1416)) or (layer7_outputs(14));
    layer8_outputs(1342) <= layer7_outputs(457);
    layer8_outputs(1343) <= not(layer7_outputs(1062)) or (layer7_outputs(2214));
    layer8_outputs(1344) <= (layer7_outputs(1261)) xor (layer7_outputs(4104));
    layer8_outputs(1345) <= (layer7_outputs(426)) xor (layer7_outputs(3091));
    layer8_outputs(1346) <= not(layer7_outputs(2019));
    layer8_outputs(1347) <= not((layer7_outputs(3739)) and (layer7_outputs(3200)));
    layer8_outputs(1348) <= not(layer7_outputs(2630));
    layer8_outputs(1349) <= (layer7_outputs(4560)) and not (layer7_outputs(3281));
    layer8_outputs(1350) <= '0';
    layer8_outputs(1351) <= not((layer7_outputs(2590)) xor (layer7_outputs(2676)));
    layer8_outputs(1352) <= layer7_outputs(4946);
    layer8_outputs(1353) <= (layer7_outputs(3397)) or (layer7_outputs(406));
    layer8_outputs(1354) <= not(layer7_outputs(750));
    layer8_outputs(1355) <= not(layer7_outputs(3960));
    layer8_outputs(1356) <= not(layer7_outputs(5001)) or (layer7_outputs(2098));
    layer8_outputs(1357) <= layer7_outputs(4896);
    layer8_outputs(1358) <= (layer7_outputs(3614)) and not (layer7_outputs(2852));
    layer8_outputs(1359) <= layer7_outputs(1504);
    layer8_outputs(1360) <= not(layer7_outputs(4581)) or (layer7_outputs(3828));
    layer8_outputs(1361) <= layer7_outputs(2282);
    layer8_outputs(1362) <= layer7_outputs(3366);
    layer8_outputs(1363) <= (layer7_outputs(1354)) xor (layer7_outputs(3406));
    layer8_outputs(1364) <= layer7_outputs(1637);
    layer8_outputs(1365) <= (layer7_outputs(4199)) and not (layer7_outputs(1157));
    layer8_outputs(1366) <= not(layer7_outputs(3034));
    layer8_outputs(1367) <= not((layer7_outputs(293)) or (layer7_outputs(1313)));
    layer8_outputs(1368) <= layer7_outputs(933);
    layer8_outputs(1369) <= layer7_outputs(529);
    layer8_outputs(1370) <= not((layer7_outputs(207)) and (layer7_outputs(3861)));
    layer8_outputs(1371) <= not((layer7_outputs(2721)) xor (layer7_outputs(671)));
    layer8_outputs(1372) <= layer7_outputs(1408);
    layer8_outputs(1373) <= not((layer7_outputs(4628)) xor (layer7_outputs(4223)));
    layer8_outputs(1374) <= layer7_outputs(4460);
    layer8_outputs(1375) <= (layer7_outputs(1304)) xor (layer7_outputs(2305));
    layer8_outputs(1376) <= not(layer7_outputs(3008));
    layer8_outputs(1377) <= not(layer7_outputs(337)) or (layer7_outputs(934));
    layer8_outputs(1378) <= not(layer7_outputs(938));
    layer8_outputs(1379) <= not((layer7_outputs(169)) and (layer7_outputs(4068)));
    layer8_outputs(1380) <= not(layer7_outputs(3875)) or (layer7_outputs(1754));
    layer8_outputs(1381) <= layer7_outputs(1390);
    layer8_outputs(1382) <= (layer7_outputs(820)) and not (layer7_outputs(3018));
    layer8_outputs(1383) <= (layer7_outputs(1011)) xor (layer7_outputs(521));
    layer8_outputs(1384) <= not(layer7_outputs(2127));
    layer8_outputs(1385) <= not(layer7_outputs(3406));
    layer8_outputs(1386) <= (layer7_outputs(130)) and (layer7_outputs(397));
    layer8_outputs(1387) <= not(layer7_outputs(196)) or (layer7_outputs(2208));
    layer8_outputs(1388) <= not(layer7_outputs(158));
    layer8_outputs(1389) <= (layer7_outputs(170)) and not (layer7_outputs(1713));
    layer8_outputs(1390) <= not(layer7_outputs(1996));
    layer8_outputs(1391) <= not(layer7_outputs(1843));
    layer8_outputs(1392) <= not(layer7_outputs(2082));
    layer8_outputs(1393) <= not(layer7_outputs(307));
    layer8_outputs(1394) <= (layer7_outputs(3513)) xor (layer7_outputs(3065));
    layer8_outputs(1395) <= not(layer7_outputs(4837));
    layer8_outputs(1396) <= not(layer7_outputs(2225));
    layer8_outputs(1397) <= (layer7_outputs(363)) xor (layer7_outputs(3641));
    layer8_outputs(1398) <= not(layer7_outputs(4798));
    layer8_outputs(1399) <= (layer7_outputs(2428)) and not (layer7_outputs(620));
    layer8_outputs(1400) <= not((layer7_outputs(274)) and (layer7_outputs(564)));
    layer8_outputs(1401) <= layer7_outputs(5051);
    layer8_outputs(1402) <= not(layer7_outputs(1879));
    layer8_outputs(1403) <= layer7_outputs(1464);
    layer8_outputs(1404) <= not(layer7_outputs(135));
    layer8_outputs(1405) <= layer7_outputs(2632);
    layer8_outputs(1406) <= layer7_outputs(1605);
    layer8_outputs(1407) <= not((layer7_outputs(939)) xor (layer7_outputs(2280)));
    layer8_outputs(1408) <= layer7_outputs(4686);
    layer8_outputs(1409) <= (layer7_outputs(1532)) and not (layer7_outputs(226));
    layer8_outputs(1410) <= layer7_outputs(4826);
    layer8_outputs(1411) <= not((layer7_outputs(1472)) or (layer7_outputs(2442)));
    layer8_outputs(1412) <= (layer7_outputs(1248)) xor (layer7_outputs(3736));
    layer8_outputs(1413) <= not((layer7_outputs(4274)) or (layer7_outputs(2747)));
    layer8_outputs(1414) <= not(layer7_outputs(348));
    layer8_outputs(1415) <= not(layer7_outputs(340));
    layer8_outputs(1416) <= not(layer7_outputs(3418));
    layer8_outputs(1417) <= layer7_outputs(1371);
    layer8_outputs(1418) <= not(layer7_outputs(4950)) or (layer7_outputs(5072));
    layer8_outputs(1419) <= not((layer7_outputs(2670)) xor (layer7_outputs(1710)));
    layer8_outputs(1420) <= (layer7_outputs(4521)) and not (layer7_outputs(1167));
    layer8_outputs(1421) <= not(layer7_outputs(3535));
    layer8_outputs(1422) <= not(layer7_outputs(1123));
    layer8_outputs(1423) <= layer7_outputs(2251);
    layer8_outputs(1424) <= layer7_outputs(515);
    layer8_outputs(1425) <= not(layer7_outputs(4242));
    layer8_outputs(1426) <= layer7_outputs(880);
    layer8_outputs(1427) <= not(layer7_outputs(1590));
    layer8_outputs(1428) <= layer7_outputs(4291);
    layer8_outputs(1429) <= (layer7_outputs(3713)) and not (layer7_outputs(80));
    layer8_outputs(1430) <= not(layer7_outputs(4528));
    layer8_outputs(1431) <= not((layer7_outputs(339)) xor (layer7_outputs(3967)));
    layer8_outputs(1432) <= layer7_outputs(432);
    layer8_outputs(1433) <= not((layer7_outputs(3163)) xor (layer7_outputs(3131)));
    layer8_outputs(1434) <= not((layer7_outputs(2108)) xor (layer7_outputs(161)));
    layer8_outputs(1435) <= layer7_outputs(3225);
    layer8_outputs(1436) <= not((layer7_outputs(805)) xor (layer7_outputs(4213)));
    layer8_outputs(1437) <= (layer7_outputs(2444)) xor (layer7_outputs(3532));
    layer8_outputs(1438) <= not(layer7_outputs(3643));
    layer8_outputs(1439) <= layer7_outputs(1708);
    layer8_outputs(1440) <= layer7_outputs(3918);
    layer8_outputs(1441) <= not(layer7_outputs(1676));
    layer8_outputs(1442) <= (layer7_outputs(2690)) and not (layer7_outputs(322));
    layer8_outputs(1443) <= (layer7_outputs(1275)) and not (layer7_outputs(3430));
    layer8_outputs(1444) <= layer7_outputs(1712);
    layer8_outputs(1445) <= not(layer7_outputs(4842)) or (layer7_outputs(292));
    layer8_outputs(1446) <= not(layer7_outputs(2906));
    layer8_outputs(1447) <= not(layer7_outputs(163));
    layer8_outputs(1448) <= layer7_outputs(419);
    layer8_outputs(1449) <= not(layer7_outputs(2006)) or (layer7_outputs(2781));
    layer8_outputs(1450) <= (layer7_outputs(4953)) xor (layer7_outputs(719));
    layer8_outputs(1451) <= (layer7_outputs(1967)) and not (layer7_outputs(3945));
    layer8_outputs(1452) <= not(layer7_outputs(3646));
    layer8_outputs(1453) <= (layer7_outputs(4210)) xor (layer7_outputs(1518));
    layer8_outputs(1454) <= not(layer7_outputs(5056));
    layer8_outputs(1455) <= not(layer7_outputs(4283)) or (layer7_outputs(2177));
    layer8_outputs(1456) <= layer7_outputs(3968);
    layer8_outputs(1457) <= not((layer7_outputs(2435)) xor (layer7_outputs(128)));
    layer8_outputs(1458) <= layer7_outputs(1243);
    layer8_outputs(1459) <= not((layer7_outputs(3539)) xor (layer7_outputs(3023)));
    layer8_outputs(1460) <= not(layer7_outputs(3711));
    layer8_outputs(1461) <= not(layer7_outputs(720));
    layer8_outputs(1462) <= (layer7_outputs(4487)) xor (layer7_outputs(4602));
    layer8_outputs(1463) <= not(layer7_outputs(2843)) or (layer7_outputs(3423));
    layer8_outputs(1464) <= layer7_outputs(2764);
    layer8_outputs(1465) <= not(layer7_outputs(4107));
    layer8_outputs(1466) <= (layer7_outputs(900)) and (layer7_outputs(243));
    layer8_outputs(1467) <= not(layer7_outputs(4711));
    layer8_outputs(1468) <= not(layer7_outputs(4501));
    layer8_outputs(1469) <= not(layer7_outputs(519));
    layer8_outputs(1470) <= not((layer7_outputs(452)) xor (layer7_outputs(139)));
    layer8_outputs(1471) <= layer7_outputs(1545);
    layer8_outputs(1472) <= not(layer7_outputs(330));
    layer8_outputs(1473) <= not((layer7_outputs(2908)) and (layer7_outputs(3975)));
    layer8_outputs(1474) <= layer7_outputs(4238);
    layer8_outputs(1475) <= layer7_outputs(4944);
    layer8_outputs(1476) <= not(layer7_outputs(3186));
    layer8_outputs(1477) <= not((layer7_outputs(1108)) xor (layer7_outputs(1039)));
    layer8_outputs(1478) <= (layer7_outputs(310)) xor (layer7_outputs(262));
    layer8_outputs(1479) <= not(layer7_outputs(1596));
    layer8_outputs(1480) <= layer7_outputs(4613);
    layer8_outputs(1481) <= (layer7_outputs(2227)) xor (layer7_outputs(2420));
    layer8_outputs(1482) <= not((layer7_outputs(4080)) xor (layer7_outputs(4300)));
    layer8_outputs(1483) <= not((layer7_outputs(235)) xor (layer7_outputs(2763)));
    layer8_outputs(1484) <= not(layer7_outputs(1355));
    layer8_outputs(1485) <= layer7_outputs(332);
    layer8_outputs(1486) <= not(layer7_outputs(2419));
    layer8_outputs(1487) <= (layer7_outputs(2329)) and (layer7_outputs(4399));
    layer8_outputs(1488) <= not((layer7_outputs(4370)) or (layer7_outputs(2007)));
    layer8_outputs(1489) <= not(layer7_outputs(1701));
    layer8_outputs(1490) <= not(layer7_outputs(4359));
    layer8_outputs(1491) <= not(layer7_outputs(1455));
    layer8_outputs(1492) <= layer7_outputs(66);
    layer8_outputs(1493) <= not((layer7_outputs(3620)) xor (layer7_outputs(2340)));
    layer8_outputs(1494) <= not(layer7_outputs(4043));
    layer8_outputs(1495) <= layer7_outputs(1204);
    layer8_outputs(1496) <= (layer7_outputs(3911)) and not (layer7_outputs(3319));
    layer8_outputs(1497) <= not(layer7_outputs(4689));
    layer8_outputs(1498) <= not((layer7_outputs(944)) xor (layer7_outputs(295)));
    layer8_outputs(1499) <= '0';
    layer8_outputs(1500) <= (layer7_outputs(4949)) or (layer7_outputs(2149));
    layer8_outputs(1501) <= layer7_outputs(4772);
    layer8_outputs(1502) <= not(layer7_outputs(1102)) or (layer7_outputs(4971));
    layer8_outputs(1503) <= not(layer7_outputs(1079));
    layer8_outputs(1504) <= not(layer7_outputs(936)) or (layer7_outputs(2217));
    layer8_outputs(1505) <= (layer7_outputs(234)) xor (layer7_outputs(1159));
    layer8_outputs(1506) <= not(layer7_outputs(3690));
    layer8_outputs(1507) <= not(layer7_outputs(3719));
    layer8_outputs(1508) <= (layer7_outputs(594)) xor (layer7_outputs(4880));
    layer8_outputs(1509) <= not(layer7_outputs(3457));
    layer8_outputs(1510) <= not((layer7_outputs(3494)) xor (layer7_outputs(3398)));
    layer8_outputs(1511) <= not(layer7_outputs(4037));
    layer8_outputs(1512) <= not(layer7_outputs(3751));
    layer8_outputs(1513) <= not((layer7_outputs(3935)) or (layer7_outputs(4625)));
    layer8_outputs(1514) <= layer7_outputs(2615);
    layer8_outputs(1515) <= (layer7_outputs(2941)) xor (layer7_outputs(1686));
    layer8_outputs(1516) <= not(layer7_outputs(3583));
    layer8_outputs(1517) <= not((layer7_outputs(2847)) xor (layer7_outputs(1231)));
    layer8_outputs(1518) <= layer7_outputs(2040);
    layer8_outputs(1519) <= (layer7_outputs(945)) or (layer7_outputs(1035));
    layer8_outputs(1520) <= not((layer7_outputs(3959)) and (layer7_outputs(75)));
    layer8_outputs(1521) <= (layer7_outputs(3713)) xor (layer7_outputs(4990));
    layer8_outputs(1522) <= (layer7_outputs(3110)) and (layer7_outputs(841));
    layer8_outputs(1523) <= (layer7_outputs(4178)) and (layer7_outputs(1966));
    layer8_outputs(1524) <= not(layer7_outputs(2867));
    layer8_outputs(1525) <= not((layer7_outputs(674)) xor (layer7_outputs(4650)));
    layer8_outputs(1526) <= layer7_outputs(280);
    layer8_outputs(1527) <= not((layer7_outputs(4024)) xor (layer7_outputs(4010)));
    layer8_outputs(1528) <= not(layer7_outputs(5023)) or (layer7_outputs(3712));
    layer8_outputs(1529) <= not((layer7_outputs(1490)) or (layer7_outputs(2833)));
    layer8_outputs(1530) <= (layer7_outputs(1214)) and not (layer7_outputs(2461));
    layer8_outputs(1531) <= (layer7_outputs(4104)) xor (layer7_outputs(4656));
    layer8_outputs(1532) <= layer7_outputs(354);
    layer8_outputs(1533) <= not((layer7_outputs(2181)) or (layer7_outputs(2535)));
    layer8_outputs(1534) <= not(layer7_outputs(4117));
    layer8_outputs(1535) <= layer7_outputs(3106);
    layer8_outputs(1536) <= not((layer7_outputs(781)) xor (layer7_outputs(4904)));
    layer8_outputs(1537) <= not(layer7_outputs(4057));
    layer8_outputs(1538) <= not(layer7_outputs(964));
    layer8_outputs(1539) <= layer7_outputs(32);
    layer8_outputs(1540) <= layer7_outputs(3913);
    layer8_outputs(1541) <= not(layer7_outputs(3568)) or (layer7_outputs(1662));
    layer8_outputs(1542) <= not((layer7_outputs(3972)) and (layer7_outputs(1335)));
    layer8_outputs(1543) <= not(layer7_outputs(5045)) or (layer7_outputs(3155));
    layer8_outputs(1544) <= (layer7_outputs(4086)) xor (layer7_outputs(1627));
    layer8_outputs(1545) <= (layer7_outputs(2848)) and not (layer7_outputs(4153));
    layer8_outputs(1546) <= not(layer7_outputs(3167));
    layer8_outputs(1547) <= layer7_outputs(675);
    layer8_outputs(1548) <= not((layer7_outputs(4622)) xor (layer7_outputs(2968)));
    layer8_outputs(1549) <= not(layer7_outputs(4254));
    layer8_outputs(1550) <= (layer7_outputs(1631)) or (layer7_outputs(3400));
    layer8_outputs(1551) <= not(layer7_outputs(4956));
    layer8_outputs(1552) <= not(layer7_outputs(2782)) or (layer7_outputs(586));
    layer8_outputs(1553) <= layer7_outputs(2565);
    layer8_outputs(1554) <= layer7_outputs(4422);
    layer8_outputs(1555) <= not((layer7_outputs(1964)) xor (layer7_outputs(392)));
    layer8_outputs(1556) <= not((layer7_outputs(699)) xor (layer7_outputs(3477)));
    layer8_outputs(1557) <= not(layer7_outputs(2599));
    layer8_outputs(1558) <= (layer7_outputs(4579)) and (layer7_outputs(1697));
    layer8_outputs(1559) <= not(layer7_outputs(3150));
    layer8_outputs(1560) <= not((layer7_outputs(3292)) xor (layer7_outputs(3053)));
    layer8_outputs(1561) <= layer7_outputs(998);
    layer8_outputs(1562) <= (layer7_outputs(3443)) xor (layer7_outputs(4241));
    layer8_outputs(1563) <= '1';
    layer8_outputs(1564) <= not((layer7_outputs(792)) xor (layer7_outputs(624)));
    layer8_outputs(1565) <= layer7_outputs(2711);
    layer8_outputs(1566) <= (layer7_outputs(3684)) and not (layer7_outputs(1589));
    layer8_outputs(1567) <= layer7_outputs(4636);
    layer8_outputs(1568) <= not(layer7_outputs(2872));
    layer8_outputs(1569) <= not(layer7_outputs(485));
    layer8_outputs(1570) <= (layer7_outputs(4960)) xor (layer7_outputs(151));
    layer8_outputs(1571) <= not(layer7_outputs(3763)) or (layer7_outputs(3071));
    layer8_outputs(1572) <= layer7_outputs(3236);
    layer8_outputs(1573) <= not((layer7_outputs(1887)) xor (layer7_outputs(3591)));
    layer8_outputs(1574) <= (layer7_outputs(3353)) xor (layer7_outputs(3160));
    layer8_outputs(1575) <= layer7_outputs(4198);
    layer8_outputs(1576) <= not(layer7_outputs(2039)) or (layer7_outputs(4000));
    layer8_outputs(1577) <= not(layer7_outputs(2421)) or (layer7_outputs(2443));
    layer8_outputs(1578) <= (layer7_outputs(2835)) xor (layer7_outputs(4848));
    layer8_outputs(1579) <= not(layer7_outputs(1004)) or (layer7_outputs(4282));
    layer8_outputs(1580) <= not(layer7_outputs(2522));
    layer8_outputs(1581) <= (layer7_outputs(3876)) and not (layer7_outputs(1144));
    layer8_outputs(1582) <= not((layer7_outputs(4393)) xor (layer7_outputs(3908)));
    layer8_outputs(1583) <= layer7_outputs(822);
    layer8_outputs(1584) <= layer7_outputs(181);
    layer8_outputs(1585) <= (layer7_outputs(2284)) xor (layer7_outputs(3700));
    layer8_outputs(1586) <= not(layer7_outputs(17));
    layer8_outputs(1587) <= layer7_outputs(3807);
    layer8_outputs(1588) <= layer7_outputs(4571);
    layer8_outputs(1589) <= not((layer7_outputs(2420)) or (layer7_outputs(1858)));
    layer8_outputs(1590) <= not((layer7_outputs(5059)) xor (layer7_outputs(165)));
    layer8_outputs(1591) <= not(layer7_outputs(1634));
    layer8_outputs(1592) <= not(layer7_outputs(3966));
    layer8_outputs(1593) <= (layer7_outputs(3276)) xor (layer7_outputs(3622));
    layer8_outputs(1594) <= not((layer7_outputs(3237)) xor (layer7_outputs(1033)));
    layer8_outputs(1595) <= not(layer7_outputs(3425));
    layer8_outputs(1596) <= (layer7_outputs(3716)) xor (layer7_outputs(4561));
    layer8_outputs(1597) <= not(layer7_outputs(2954));
    layer8_outputs(1598) <= layer7_outputs(4458);
    layer8_outputs(1599) <= not((layer7_outputs(2408)) xor (layer7_outputs(3341)));
    layer8_outputs(1600) <= not(layer7_outputs(3846));
    layer8_outputs(1601) <= not(layer7_outputs(963)) or (layer7_outputs(1030));
    layer8_outputs(1602) <= not(layer7_outputs(1398));
    layer8_outputs(1603) <= not(layer7_outputs(765));
    layer8_outputs(1604) <= not(layer7_outputs(2221));
    layer8_outputs(1605) <= (layer7_outputs(958)) xor (layer7_outputs(4952));
    layer8_outputs(1606) <= '1';
    layer8_outputs(1607) <= (layer7_outputs(4562)) and (layer7_outputs(882));
    layer8_outputs(1608) <= (layer7_outputs(3302)) and not (layer7_outputs(1669));
    layer8_outputs(1609) <= not((layer7_outputs(3771)) xor (layer7_outputs(2228)));
    layer8_outputs(1610) <= (layer7_outputs(4855)) and not (layer7_outputs(2695));
    layer8_outputs(1611) <= layer7_outputs(2107);
    layer8_outputs(1612) <= (layer7_outputs(3524)) xor (layer7_outputs(2505));
    layer8_outputs(1613) <= not(layer7_outputs(171));
    layer8_outputs(1614) <= not(layer7_outputs(1987));
    layer8_outputs(1615) <= layer7_outputs(469);
    layer8_outputs(1616) <= layer7_outputs(3164);
    layer8_outputs(1617) <= (layer7_outputs(546)) xor (layer7_outputs(2876));
    layer8_outputs(1618) <= not(layer7_outputs(1971));
    layer8_outputs(1619) <= layer7_outputs(535);
    layer8_outputs(1620) <= (layer7_outputs(2750)) or (layer7_outputs(1730));
    layer8_outputs(1621) <= layer7_outputs(372);
    layer8_outputs(1622) <= not((layer7_outputs(4463)) xor (layer7_outputs(1736)));
    layer8_outputs(1623) <= not(layer7_outputs(4672));
    layer8_outputs(1624) <= layer7_outputs(2068);
    layer8_outputs(1625) <= not(layer7_outputs(2075));
    layer8_outputs(1626) <= not(layer7_outputs(3723));
    layer8_outputs(1627) <= not(layer7_outputs(730));
    layer8_outputs(1628) <= not(layer7_outputs(4523));
    layer8_outputs(1629) <= not(layer7_outputs(3401));
    layer8_outputs(1630) <= layer7_outputs(38);
    layer8_outputs(1631) <= layer7_outputs(4001);
    layer8_outputs(1632) <= not(layer7_outputs(1160)) or (layer7_outputs(93));
    layer8_outputs(1633) <= layer7_outputs(187);
    layer8_outputs(1634) <= not((layer7_outputs(1286)) xor (layer7_outputs(1661)));
    layer8_outputs(1635) <= not(layer7_outputs(3468));
    layer8_outputs(1636) <= (layer7_outputs(3059)) and not (layer7_outputs(60));
    layer8_outputs(1637) <= layer7_outputs(2538);
    layer8_outputs(1638) <= (layer7_outputs(2267)) or (layer7_outputs(1207));
    layer8_outputs(1639) <= (layer7_outputs(952)) or (layer7_outputs(4077));
    layer8_outputs(1640) <= layer7_outputs(669);
    layer8_outputs(1641) <= (layer7_outputs(3227)) and (layer7_outputs(5034));
    layer8_outputs(1642) <= (layer7_outputs(1481)) xor (layer7_outputs(2361));
    layer8_outputs(1643) <= (layer7_outputs(2027)) or (layer7_outputs(4967));
    layer8_outputs(1644) <= layer7_outputs(2453);
    layer8_outputs(1645) <= not(layer7_outputs(3112));
    layer8_outputs(1646) <= layer7_outputs(4785);
    layer8_outputs(1647) <= layer7_outputs(2752);
    layer8_outputs(1648) <= (layer7_outputs(218)) xor (layer7_outputs(4409));
    layer8_outputs(1649) <= '1';
    layer8_outputs(1650) <= not(layer7_outputs(1999)) or (layer7_outputs(3508));
    layer8_outputs(1651) <= not(layer7_outputs(780)) or (layer7_outputs(1163));
    layer8_outputs(1652) <= (layer7_outputs(4623)) xor (layer7_outputs(1448));
    layer8_outputs(1653) <= not(layer7_outputs(5078)) or (layer7_outputs(3955));
    layer8_outputs(1654) <= not(layer7_outputs(3909));
    layer8_outputs(1655) <= not(layer7_outputs(1760));
    layer8_outputs(1656) <= layer7_outputs(3197);
    layer8_outputs(1657) <= not((layer7_outputs(2561)) and (layer7_outputs(2851)));
    layer8_outputs(1658) <= not(layer7_outputs(4933));
    layer8_outputs(1659) <= not(layer7_outputs(709));
    layer8_outputs(1660) <= (layer7_outputs(2460)) or (layer7_outputs(612));
    layer8_outputs(1661) <= not((layer7_outputs(260)) and (layer7_outputs(3458)));
    layer8_outputs(1662) <= not(layer7_outputs(2294)) or (layer7_outputs(1185));
    layer8_outputs(1663) <= not(layer7_outputs(2802));
    layer8_outputs(1664) <= (layer7_outputs(2657)) xor (layer7_outputs(4344));
    layer8_outputs(1665) <= not((layer7_outputs(2374)) xor (layer7_outputs(4797)));
    layer8_outputs(1666) <= (layer7_outputs(3322)) or (layer7_outputs(1410));
    layer8_outputs(1667) <= layer7_outputs(847);
    layer8_outputs(1668) <= not(layer7_outputs(3689));
    layer8_outputs(1669) <= not(layer7_outputs(1726));
    layer8_outputs(1670) <= layer7_outputs(4059);
    layer8_outputs(1671) <= not((layer7_outputs(3481)) or (layer7_outputs(359)));
    layer8_outputs(1672) <= (layer7_outputs(3692)) and not (layer7_outputs(1755));
    layer8_outputs(1673) <= (layer7_outputs(4013)) and (layer7_outputs(2489));
    layer8_outputs(1674) <= not(layer7_outputs(145));
    layer8_outputs(1675) <= not((layer7_outputs(585)) xor (layer7_outputs(524)));
    layer8_outputs(1676) <= (layer7_outputs(1872)) or (layer7_outputs(2314));
    layer8_outputs(1677) <= (layer7_outputs(2951)) and (layer7_outputs(3335));
    layer8_outputs(1678) <= (layer7_outputs(4776)) and not (layer7_outputs(95));
    layer8_outputs(1679) <= (layer7_outputs(574)) xor (layer7_outputs(2545));
    layer8_outputs(1680) <= not(layer7_outputs(2776)) or (layer7_outputs(2058));
    layer8_outputs(1681) <= not((layer7_outputs(2722)) or (layer7_outputs(2097)));
    layer8_outputs(1682) <= not((layer7_outputs(2162)) xor (layer7_outputs(3071)));
    layer8_outputs(1683) <= not(layer7_outputs(3598));
    layer8_outputs(1684) <= not(layer7_outputs(1233)) or (layer7_outputs(1950));
    layer8_outputs(1685) <= '1';
    layer8_outputs(1686) <= layer7_outputs(4459);
    layer8_outputs(1687) <= '0';
    layer8_outputs(1688) <= layer7_outputs(1301);
    layer8_outputs(1689) <= not(layer7_outputs(3785));
    layer8_outputs(1690) <= not(layer7_outputs(3855));
    layer8_outputs(1691) <= not((layer7_outputs(1958)) or (layer7_outputs(505)));
    layer8_outputs(1692) <= not((layer7_outputs(211)) xor (layer7_outputs(3182)));
    layer8_outputs(1693) <= (layer7_outputs(2704)) xor (layer7_outputs(914));
    layer8_outputs(1694) <= layer7_outputs(1446);
    layer8_outputs(1695) <= (layer7_outputs(1561)) and not (layer7_outputs(2771));
    layer8_outputs(1696) <= (layer7_outputs(227)) xor (layer7_outputs(1279));
    layer8_outputs(1697) <= not(layer7_outputs(3817));
    layer8_outputs(1698) <= not(layer7_outputs(3258));
    layer8_outputs(1699) <= not((layer7_outputs(732)) xor (layer7_outputs(4638)));
    layer8_outputs(1700) <= layer7_outputs(81);
    layer8_outputs(1701) <= not(layer7_outputs(1304)) or (layer7_outputs(1107));
    layer8_outputs(1702) <= not(layer7_outputs(1316));
    layer8_outputs(1703) <= not(layer7_outputs(3420)) or (layer7_outputs(3152));
    layer8_outputs(1704) <= layer7_outputs(3069);
    layer8_outputs(1705) <= not((layer7_outputs(566)) xor (layer7_outputs(3173)));
    layer8_outputs(1706) <= layer7_outputs(445);
    layer8_outputs(1707) <= (layer7_outputs(4901)) xor (layer7_outputs(5020));
    layer8_outputs(1708) <= not(layer7_outputs(2857));
    layer8_outputs(1709) <= not((layer7_outputs(3022)) xor (layer7_outputs(525)));
    layer8_outputs(1710) <= not(layer7_outputs(2820)) or (layer7_outputs(2958));
    layer8_outputs(1711) <= not((layer7_outputs(3995)) and (layer7_outputs(539)));
    layer8_outputs(1712) <= not(layer7_outputs(4770));
    layer8_outputs(1713) <= layer7_outputs(2952);
    layer8_outputs(1714) <= (layer7_outputs(750)) or (layer7_outputs(3404));
    layer8_outputs(1715) <= '0';
    layer8_outputs(1716) <= not(layer7_outputs(302));
    layer8_outputs(1717) <= layer7_outputs(104);
    layer8_outputs(1718) <= not((layer7_outputs(725)) xor (layer7_outputs(888)));
    layer8_outputs(1719) <= (layer7_outputs(2129)) and not (layer7_outputs(3899));
    layer8_outputs(1720) <= layer7_outputs(1347);
    layer8_outputs(1721) <= not(layer7_outputs(3894));
    layer8_outputs(1722) <= (layer7_outputs(882)) xor (layer7_outputs(1536));
    layer8_outputs(1723) <= not((layer7_outputs(2235)) xor (layer7_outputs(2110)));
    layer8_outputs(1724) <= not(layer7_outputs(2180));
    layer8_outputs(1725) <= not(layer7_outputs(1927));
    layer8_outputs(1726) <= (layer7_outputs(1206)) and not (layer7_outputs(1388));
    layer8_outputs(1727) <= not((layer7_outputs(2700)) xor (layer7_outputs(3645)));
    layer8_outputs(1728) <= not(layer7_outputs(4202)) or (layer7_outputs(4195));
    layer8_outputs(1729) <= not(layer7_outputs(3495));
    layer8_outputs(1730) <= layer7_outputs(5);
    layer8_outputs(1731) <= not((layer7_outputs(4884)) xor (layer7_outputs(21)));
    layer8_outputs(1732) <= layer7_outputs(88);
    layer8_outputs(1733) <= layer7_outputs(1373);
    layer8_outputs(1734) <= '0';
    layer8_outputs(1735) <= layer7_outputs(2350);
    layer8_outputs(1736) <= layer7_outputs(2110);
    layer8_outputs(1737) <= (layer7_outputs(2531)) or (layer7_outputs(425));
    layer8_outputs(1738) <= not(layer7_outputs(2755));
    layer8_outputs(1739) <= not((layer7_outputs(714)) or (layer7_outputs(2718)));
    layer8_outputs(1740) <= not((layer7_outputs(390)) or (layer7_outputs(1590)));
    layer8_outputs(1741) <= (layer7_outputs(3903)) xor (layer7_outputs(3470));
    layer8_outputs(1742) <= not(layer7_outputs(2099)) or (layer7_outputs(147));
    layer8_outputs(1743) <= not(layer7_outputs(183));
    layer8_outputs(1744) <= layer7_outputs(2558);
    layer8_outputs(1745) <= (layer7_outputs(3428)) xor (layer7_outputs(2257));
    layer8_outputs(1746) <= not(layer7_outputs(1104)) or (layer7_outputs(974));
    layer8_outputs(1747) <= (layer7_outputs(442)) and not (layer7_outputs(3699));
    layer8_outputs(1748) <= layer7_outputs(1384);
    layer8_outputs(1749) <= not(layer7_outputs(4231));
    layer8_outputs(1750) <= not(layer7_outputs(1699));
    layer8_outputs(1751) <= layer7_outputs(1435);
    layer8_outputs(1752) <= layer7_outputs(2611);
    layer8_outputs(1753) <= not((layer7_outputs(3)) xor (layer7_outputs(4443)));
    layer8_outputs(1754) <= not(layer7_outputs(3188)) or (layer7_outputs(2477));
    layer8_outputs(1755) <= not((layer7_outputs(362)) and (layer7_outputs(326)));
    layer8_outputs(1756) <= layer7_outputs(4846);
    layer8_outputs(1757) <= not((layer7_outputs(1972)) xor (layer7_outputs(445)));
    layer8_outputs(1758) <= layer7_outputs(1863);
    layer8_outputs(1759) <= not((layer7_outputs(3519)) xor (layer7_outputs(173)));
    layer8_outputs(1760) <= not((layer7_outputs(5104)) and (layer7_outputs(613)));
    layer8_outputs(1761) <= layer7_outputs(885);
    layer8_outputs(1762) <= layer7_outputs(782);
    layer8_outputs(1763) <= (layer7_outputs(4351)) and not (layer7_outputs(2248));
    layer8_outputs(1764) <= not(layer7_outputs(2131));
    layer8_outputs(1765) <= not(layer7_outputs(2192));
    layer8_outputs(1766) <= not((layer7_outputs(3791)) and (layer7_outputs(1450)));
    layer8_outputs(1767) <= (layer7_outputs(4752)) and not (layer7_outputs(1534));
    layer8_outputs(1768) <= layer7_outputs(4819);
    layer8_outputs(1769) <= layer7_outputs(2894);
    layer8_outputs(1770) <= not((layer7_outputs(2620)) and (layer7_outputs(3371)));
    layer8_outputs(1771) <= (layer7_outputs(2613)) xor (layer7_outputs(4170));
    layer8_outputs(1772) <= (layer7_outputs(3369)) and not (layer7_outputs(1351));
    layer8_outputs(1773) <= not(layer7_outputs(4885));
    layer8_outputs(1774) <= not(layer7_outputs(4051));
    layer8_outputs(1775) <= not(layer7_outputs(1296));
    layer8_outputs(1776) <= not(layer7_outputs(1158));
    layer8_outputs(1777) <= not(layer7_outputs(1425)) or (layer7_outputs(1832));
    layer8_outputs(1778) <= not(layer7_outputs(3151));
    layer8_outputs(1779) <= layer7_outputs(4454);
    layer8_outputs(1780) <= not(layer7_outputs(2326));
    layer8_outputs(1781) <= (layer7_outputs(4697)) or (layer7_outputs(4761));
    layer8_outputs(1782) <= not((layer7_outputs(2370)) and (layer7_outputs(523)));
    layer8_outputs(1783) <= layer7_outputs(4550);
    layer8_outputs(1784) <= not(layer7_outputs(4151));
    layer8_outputs(1785) <= layer7_outputs(4212);
    layer8_outputs(1786) <= (layer7_outputs(2065)) or (layer7_outputs(3308));
    layer8_outputs(1787) <= not((layer7_outputs(5117)) xor (layer7_outputs(41)));
    layer8_outputs(1788) <= not(layer7_outputs(3563));
    layer8_outputs(1789) <= not((layer7_outputs(3788)) and (layer7_outputs(726)));
    layer8_outputs(1790) <= not((layer7_outputs(4322)) and (layer7_outputs(4194)));
    layer8_outputs(1791) <= not(layer7_outputs(4934));
    layer8_outputs(1792) <= not(layer7_outputs(2523));
    layer8_outputs(1793) <= layer7_outputs(2871);
    layer8_outputs(1794) <= not(layer7_outputs(1801)) or (layer7_outputs(768));
    layer8_outputs(1795) <= not(layer7_outputs(2639));
    layer8_outputs(1796) <= not((layer7_outputs(1399)) xor (layer7_outputs(2969)));
    layer8_outputs(1797) <= not(layer7_outputs(2762));
    layer8_outputs(1798) <= (layer7_outputs(2438)) xor (layer7_outputs(1203));
    layer8_outputs(1799) <= (layer7_outputs(3322)) xor (layer7_outputs(1361));
    layer8_outputs(1800) <= not((layer7_outputs(3062)) and (layer7_outputs(1744)));
    layer8_outputs(1801) <= layer7_outputs(4936);
    layer8_outputs(1802) <= layer7_outputs(866);
    layer8_outputs(1803) <= layer7_outputs(5072);
    layer8_outputs(1804) <= (layer7_outputs(152)) xor (layer7_outputs(436));
    layer8_outputs(1805) <= layer7_outputs(4611);
    layer8_outputs(1806) <= (layer7_outputs(1620)) xor (layer7_outputs(3762));
    layer8_outputs(1807) <= layer7_outputs(1309);
    layer8_outputs(1808) <= not(layer7_outputs(1176));
    layer8_outputs(1809) <= not((layer7_outputs(2908)) xor (layer7_outputs(3135)));
    layer8_outputs(1810) <= (layer7_outputs(1934)) or (layer7_outputs(198));
    layer8_outputs(1811) <= not((layer7_outputs(4482)) and (layer7_outputs(810)));
    layer8_outputs(1812) <= (layer7_outputs(2889)) or (layer7_outputs(3145));
    layer8_outputs(1813) <= layer7_outputs(2394);
    layer8_outputs(1814) <= layer7_outputs(1612);
    layer8_outputs(1815) <= not(layer7_outputs(4408));
    layer8_outputs(1816) <= not(layer7_outputs(2967));
    layer8_outputs(1817) <= (layer7_outputs(2021)) xor (layer7_outputs(659));
    layer8_outputs(1818) <= not(layer7_outputs(383));
    layer8_outputs(1819) <= not((layer7_outputs(3533)) xor (layer7_outputs(4541)));
    layer8_outputs(1820) <= not((layer7_outputs(89)) xor (layer7_outputs(2385)));
    layer8_outputs(1821) <= not(layer7_outputs(865));
    layer8_outputs(1822) <= (layer7_outputs(2936)) and not (layer7_outputs(4515));
    layer8_outputs(1823) <= (layer7_outputs(1431)) and not (layer7_outputs(310));
    layer8_outputs(1824) <= layer7_outputs(99);
    layer8_outputs(1825) <= not((layer7_outputs(3839)) xor (layer7_outputs(3742)));
    layer8_outputs(1826) <= layer7_outputs(721);
    layer8_outputs(1827) <= layer7_outputs(444);
    layer8_outputs(1828) <= layer7_outputs(1025);
    layer8_outputs(1829) <= not((layer7_outputs(2498)) xor (layer7_outputs(3077)));
    layer8_outputs(1830) <= not(layer7_outputs(1486));
    layer8_outputs(1831) <= not((layer7_outputs(4546)) and (layer7_outputs(5054)));
    layer8_outputs(1832) <= (layer7_outputs(813)) and not (layer7_outputs(1877));
    layer8_outputs(1833) <= '1';
    layer8_outputs(1834) <= (layer7_outputs(3012)) and not (layer7_outputs(3693));
    layer8_outputs(1835) <= (layer7_outputs(3006)) or (layer7_outputs(117));
    layer8_outputs(1836) <= not((layer7_outputs(2384)) or (layer7_outputs(4285)));
    layer8_outputs(1837) <= not(layer7_outputs(4129));
    layer8_outputs(1838) <= not((layer7_outputs(2712)) xor (layer7_outputs(4677)));
    layer8_outputs(1839) <= layer7_outputs(1691);
    layer8_outputs(1840) <= not(layer7_outputs(1530));
    layer8_outputs(1841) <= not(layer7_outputs(1219));
    layer8_outputs(1842) <= not((layer7_outputs(5020)) and (layer7_outputs(2656)));
    layer8_outputs(1843) <= not((layer7_outputs(3860)) xor (layer7_outputs(4078)));
    layer8_outputs(1844) <= not(layer7_outputs(1831));
    layer8_outputs(1845) <= not((layer7_outputs(3485)) xor (layer7_outputs(3180)));
    layer8_outputs(1846) <= not(layer7_outputs(2678));
    layer8_outputs(1847) <= '0';
    layer8_outputs(1848) <= layer7_outputs(3696);
    layer8_outputs(1849) <= (layer7_outputs(1436)) or (layer7_outputs(2534));
    layer8_outputs(1850) <= (layer7_outputs(4629)) and (layer7_outputs(76));
    layer8_outputs(1851) <= not((layer7_outputs(3055)) xor (layer7_outputs(4809)));
    layer8_outputs(1852) <= not(layer7_outputs(3841));
    layer8_outputs(1853) <= not((layer7_outputs(1303)) and (layer7_outputs(118)));
    layer8_outputs(1854) <= not(layer7_outputs(3273));
    layer8_outputs(1855) <= (layer7_outputs(1100)) xor (layer7_outputs(374));
    layer8_outputs(1856) <= (layer7_outputs(3624)) or (layer7_outputs(3549));
    layer8_outputs(1857) <= (layer7_outputs(2751)) xor (layer7_outputs(142));
    layer8_outputs(1858) <= layer7_outputs(5087);
    layer8_outputs(1859) <= not((layer7_outputs(5093)) or (layer7_outputs(3268)));
    layer8_outputs(1860) <= not(layer7_outputs(966));
    layer8_outputs(1861) <= not(layer7_outputs(1740));
    layer8_outputs(1862) <= layer7_outputs(2350);
    layer8_outputs(1863) <= layer7_outputs(3057);
    layer8_outputs(1864) <= (layer7_outputs(337)) xor (layer7_outputs(1829));
    layer8_outputs(1865) <= layer7_outputs(3291);
    layer8_outputs(1866) <= not(layer7_outputs(1704)) or (layer7_outputs(2717));
    layer8_outputs(1867) <= not((layer7_outputs(2203)) or (layer7_outputs(4631)));
    layer8_outputs(1868) <= not((layer7_outputs(2604)) or (layer7_outputs(3579)));
    layer8_outputs(1869) <= not(layer7_outputs(3041));
    layer8_outputs(1870) <= layer7_outputs(4779);
    layer8_outputs(1871) <= layer7_outputs(373);
    layer8_outputs(1872) <= layer7_outputs(300);
    layer8_outputs(1873) <= not(layer7_outputs(2208)) or (layer7_outputs(4466));
    layer8_outputs(1874) <= not(layer7_outputs(2567)) or (layer7_outputs(3668));
    layer8_outputs(1875) <= not((layer7_outputs(4522)) xor (layer7_outputs(793)));
    layer8_outputs(1876) <= (layer7_outputs(4030)) xor (layer7_outputs(927));
    layer8_outputs(1877) <= not(layer7_outputs(1461));
    layer8_outputs(1878) <= layer7_outputs(967);
    layer8_outputs(1879) <= not(layer7_outputs(2942));
    layer8_outputs(1880) <= not(layer7_outputs(1252));
    layer8_outputs(1881) <= not((layer7_outputs(3367)) xor (layer7_outputs(4294)));
    layer8_outputs(1882) <= not(layer7_outputs(3221));
    layer8_outputs(1883) <= (layer7_outputs(4442)) and not (layer7_outputs(570));
    layer8_outputs(1884) <= (layer7_outputs(1965)) or (layer7_outputs(208));
    layer8_outputs(1885) <= layer7_outputs(2221);
    layer8_outputs(1886) <= (layer7_outputs(967)) xor (layer7_outputs(3752));
    layer8_outputs(1887) <= (layer7_outputs(4831)) and (layer7_outputs(4270));
    layer8_outputs(1888) <= layer7_outputs(2528);
    layer8_outputs(1889) <= not(layer7_outputs(4641));
    layer8_outputs(1890) <= not(layer7_outputs(3835)) or (layer7_outputs(1349));
    layer8_outputs(1891) <= layer7_outputs(1400);
    layer8_outputs(1892) <= not(layer7_outputs(2465));
    layer8_outputs(1893) <= not((layer7_outputs(1444)) xor (layer7_outputs(4823)));
    layer8_outputs(1894) <= not(layer7_outputs(3902));
    layer8_outputs(1895) <= not(layer7_outputs(2358));
    layer8_outputs(1896) <= (layer7_outputs(2159)) and not (layer7_outputs(4110));
    layer8_outputs(1897) <= not((layer7_outputs(2899)) or (layer7_outputs(3239)));
    layer8_outputs(1898) <= not(layer7_outputs(4805));
    layer8_outputs(1899) <= not((layer7_outputs(4863)) xor (layer7_outputs(1332)));
    layer8_outputs(1900) <= layer7_outputs(1131);
    layer8_outputs(1901) <= layer7_outputs(503);
    layer8_outputs(1902) <= (layer7_outputs(1207)) and (layer7_outputs(3678));
    layer8_outputs(1903) <= (layer7_outputs(4648)) xor (layer7_outputs(4188));
    layer8_outputs(1904) <= not(layer7_outputs(4061));
    layer8_outputs(1905) <= not((layer7_outputs(4042)) xor (layer7_outputs(240)));
    layer8_outputs(1906) <= (layer7_outputs(1871)) or (layer7_outputs(1342));
    layer8_outputs(1907) <= not(layer7_outputs(2998));
    layer8_outputs(1908) <= not((layer7_outputs(4264)) xor (layer7_outputs(384)));
    layer8_outputs(1909) <= not(layer7_outputs(2300));
    layer8_outputs(1910) <= not(layer7_outputs(1317)) or (layer7_outputs(1284));
    layer8_outputs(1911) <= layer7_outputs(4211);
    layer8_outputs(1912) <= not((layer7_outputs(1929)) and (layer7_outputs(3702)));
    layer8_outputs(1913) <= not(layer7_outputs(1788));
    layer8_outputs(1914) <= not(layer7_outputs(125));
    layer8_outputs(1915) <= not(layer7_outputs(3572));
    layer8_outputs(1916) <= layer7_outputs(4105);
    layer8_outputs(1917) <= layer7_outputs(3327);
    layer8_outputs(1918) <= layer7_outputs(2551);
    layer8_outputs(1919) <= not(layer7_outputs(272));
    layer8_outputs(1920) <= (layer7_outputs(5087)) and not (layer7_outputs(3753));
    layer8_outputs(1921) <= layer7_outputs(4613);
    layer8_outputs(1922) <= (layer7_outputs(1478)) and not (layer7_outputs(2404));
    layer8_outputs(1923) <= not(layer7_outputs(1597));
    layer8_outputs(1924) <= (layer7_outputs(4904)) xor (layer7_outputs(4853));
    layer8_outputs(1925) <= not((layer7_outputs(2355)) xor (layer7_outputs(100)));
    layer8_outputs(1926) <= not(layer7_outputs(54)) or (layer7_outputs(570));
    layer8_outputs(1927) <= layer7_outputs(3503);
    layer8_outputs(1928) <= not(layer7_outputs(1303));
    layer8_outputs(1929) <= not(layer7_outputs(1509));
    layer8_outputs(1930) <= not(layer7_outputs(657)) or (layer7_outputs(1424));
    layer8_outputs(1931) <= layer7_outputs(3153);
    layer8_outputs(1932) <= not(layer7_outputs(4709)) or (layer7_outputs(412));
    layer8_outputs(1933) <= not((layer7_outputs(3788)) xor (layer7_outputs(1591)));
    layer8_outputs(1934) <= (layer7_outputs(3381)) xor (layer7_outputs(2318));
    layer8_outputs(1935) <= (layer7_outputs(903)) and not (layer7_outputs(4091));
    layer8_outputs(1936) <= (layer7_outputs(3169)) xor (layer7_outputs(2680));
    layer8_outputs(1937) <= not((layer7_outputs(784)) or (layer7_outputs(2869)));
    layer8_outputs(1938) <= not(layer7_outputs(452));
    layer8_outputs(1939) <= not((layer7_outputs(492)) xor (layer7_outputs(5046)));
    layer8_outputs(1940) <= layer7_outputs(174);
    layer8_outputs(1941) <= not((layer7_outputs(4171)) xor (layer7_outputs(2354)));
    layer8_outputs(1942) <= layer7_outputs(4152);
    layer8_outputs(1943) <= (layer7_outputs(1375)) or (layer7_outputs(3248));
    layer8_outputs(1944) <= layer7_outputs(4649);
    layer8_outputs(1945) <= not(layer7_outputs(1862));
    layer8_outputs(1946) <= (layer7_outputs(4028)) xor (layer7_outputs(2187));
    layer8_outputs(1947) <= not(layer7_outputs(2080));
    layer8_outputs(1948) <= not(layer7_outputs(2911));
    layer8_outputs(1949) <= layer7_outputs(1209);
    layer8_outputs(1950) <= not(layer7_outputs(4199));
    layer8_outputs(1951) <= not(layer7_outputs(1986));
    layer8_outputs(1952) <= (layer7_outputs(2932)) and not (layer7_outputs(4983));
    layer8_outputs(1953) <= (layer7_outputs(1459)) xor (layer7_outputs(4089));
    layer8_outputs(1954) <= (layer7_outputs(579)) and not (layer7_outputs(1645));
    layer8_outputs(1955) <= not(layer7_outputs(4122));
    layer8_outputs(1956) <= not(layer7_outputs(79));
    layer8_outputs(1957) <= not((layer7_outputs(1628)) or (layer7_outputs(358)));
    layer8_outputs(1958) <= layer7_outputs(2297);
    layer8_outputs(1959) <= (layer7_outputs(1822)) and not (layer7_outputs(2275));
    layer8_outputs(1960) <= layer7_outputs(1197);
    layer8_outputs(1961) <= not(layer7_outputs(4193));
    layer8_outputs(1962) <= not(layer7_outputs(3004));
    layer8_outputs(1963) <= not(layer7_outputs(4248));
    layer8_outputs(1964) <= not((layer7_outputs(417)) xor (layer7_outputs(4451)));
    layer8_outputs(1965) <= (layer7_outputs(935)) and not (layer7_outputs(4160));
    layer8_outputs(1966) <= layer7_outputs(886);
    layer8_outputs(1967) <= (layer7_outputs(1792)) xor (layer7_outputs(1896));
    layer8_outputs(1968) <= not(layer7_outputs(2511));
    layer8_outputs(1969) <= not(layer7_outputs(1733));
    layer8_outputs(1970) <= not(layer7_outputs(399));
    layer8_outputs(1971) <= layer7_outputs(279);
    layer8_outputs(1972) <= not(layer7_outputs(464));
    layer8_outputs(1973) <= not(layer7_outputs(3649));
    layer8_outputs(1974) <= not((layer7_outputs(4652)) xor (layer7_outputs(2659)));
    layer8_outputs(1975) <= (layer7_outputs(2424)) xor (layer7_outputs(1683));
    layer8_outputs(1976) <= '1';
    layer8_outputs(1977) <= layer7_outputs(852);
    layer8_outputs(1978) <= layer7_outputs(2981);
    layer8_outputs(1979) <= not((layer7_outputs(973)) xor (layer7_outputs(3513)));
    layer8_outputs(1980) <= layer7_outputs(1795);
    layer8_outputs(1981) <= not((layer7_outputs(1664)) or (layer7_outputs(231)));
    layer8_outputs(1982) <= layer7_outputs(615);
    layer8_outputs(1983) <= layer7_outputs(1358);
    layer8_outputs(1984) <= not((layer7_outputs(3297)) or (layer7_outputs(4538)));
    layer8_outputs(1985) <= not((layer7_outputs(300)) and (layer7_outputs(1012)));
    layer8_outputs(1986) <= not(layer7_outputs(4721));
    layer8_outputs(1987) <= not(layer7_outputs(4937));
    layer8_outputs(1988) <= (layer7_outputs(4049)) or (layer7_outputs(335));
    layer8_outputs(1989) <= not(layer7_outputs(4714));
    layer8_outputs(1990) <= not((layer7_outputs(2568)) and (layer7_outputs(129)));
    layer8_outputs(1991) <= layer7_outputs(1766);
    layer8_outputs(1992) <= not(layer7_outputs(3339));
    layer8_outputs(1993) <= (layer7_outputs(3507)) xor (layer7_outputs(4196));
    layer8_outputs(1994) <= not(layer7_outputs(3491)) or (layer7_outputs(3926));
    layer8_outputs(1995) <= not(layer7_outputs(3640));
    layer8_outputs(1996) <= not(layer7_outputs(1917));
    layer8_outputs(1997) <= not(layer7_outputs(3817));
    layer8_outputs(1998) <= not(layer7_outputs(3973));
    layer8_outputs(1999) <= layer7_outputs(4396);
    layer8_outputs(2000) <= not((layer7_outputs(4696)) xor (layer7_outputs(313)));
    layer8_outputs(2001) <= not(layer7_outputs(352));
    layer8_outputs(2002) <= layer7_outputs(1566);
    layer8_outputs(2003) <= not((layer7_outputs(3895)) xor (layer7_outputs(3384)));
    layer8_outputs(2004) <= (layer7_outputs(2144)) xor (layer7_outputs(3271));
    layer8_outputs(2005) <= not(layer7_outputs(1346));
    layer8_outputs(2006) <= layer7_outputs(2923);
    layer8_outputs(2007) <= not((layer7_outputs(3885)) or (layer7_outputs(3206)));
    layer8_outputs(2008) <= not((layer7_outputs(990)) xor (layer7_outputs(4647)));
    layer8_outputs(2009) <= (layer7_outputs(22)) and not (layer7_outputs(2212));
    layer8_outputs(2010) <= not(layer7_outputs(2707));
    layer8_outputs(2011) <= layer7_outputs(3073);
    layer8_outputs(2012) <= layer7_outputs(3941);
    layer8_outputs(2013) <= not(layer7_outputs(1885));
    layer8_outputs(2014) <= not((layer7_outputs(3782)) xor (layer7_outputs(309)));
    layer8_outputs(2015) <= (layer7_outputs(113)) xor (layer7_outputs(2112));
    layer8_outputs(2016) <= layer7_outputs(4102);
    layer8_outputs(2017) <= not(layer7_outputs(219));
    layer8_outputs(2018) <= (layer7_outputs(2036)) and (layer7_outputs(2387));
    layer8_outputs(2019) <= (layer7_outputs(1593)) and not (layer7_outputs(4295));
    layer8_outputs(2020) <= '0';
    layer8_outputs(2021) <= not((layer7_outputs(1012)) xor (layer7_outputs(3232)));
    layer8_outputs(2022) <= layer7_outputs(3939);
    layer8_outputs(2023) <= layer7_outputs(322);
    layer8_outputs(2024) <= layer7_outputs(2605);
    layer8_outputs(2025) <= not(layer7_outputs(510)) or (layer7_outputs(1086));
    layer8_outputs(2026) <= (layer7_outputs(1379)) xor (layer7_outputs(508));
    layer8_outputs(2027) <= layer7_outputs(3800);
    layer8_outputs(2028) <= not(layer7_outputs(438));
    layer8_outputs(2029) <= layer7_outputs(1019);
    layer8_outputs(2030) <= not((layer7_outputs(401)) and (layer7_outputs(3360)));
    layer8_outputs(2031) <= not(layer7_outputs(3020));
    layer8_outputs(2032) <= not((layer7_outputs(1611)) and (layer7_outputs(3618)));
    layer8_outputs(2033) <= not(layer7_outputs(259)) or (layer7_outputs(4842));
    layer8_outputs(2034) <= (layer7_outputs(1664)) xor (layer7_outputs(3254));
    layer8_outputs(2035) <= not((layer7_outputs(4288)) xor (layer7_outputs(1287)));
    layer8_outputs(2036) <= not(layer7_outputs(2118));
    layer8_outputs(2037) <= not(layer7_outputs(3375));
    layer8_outputs(2038) <= not(layer7_outputs(4795));
    layer8_outputs(2039) <= not(layer7_outputs(1646));
    layer8_outputs(2040) <= not(layer7_outputs(3595));
    layer8_outputs(2041) <= not(layer7_outputs(1505));
    layer8_outputs(2042) <= not(layer7_outputs(669));
    layer8_outputs(2043) <= (layer7_outputs(3133)) and not (layer7_outputs(1441));
    layer8_outputs(2044) <= not(layer7_outputs(2903));
    layer8_outputs(2045) <= not((layer7_outputs(4367)) xor (layer7_outputs(891)));
    layer8_outputs(2046) <= layer7_outputs(4670);
    layer8_outputs(2047) <= '1';
    layer8_outputs(2048) <= not(layer7_outputs(3471));
    layer8_outputs(2049) <= layer7_outputs(1438);
    layer8_outputs(2050) <= not(layer7_outputs(3768));
    layer8_outputs(2051) <= (layer7_outputs(2395)) and not (layer7_outputs(1449));
    layer8_outputs(2052) <= not(layer7_outputs(250));
    layer8_outputs(2053) <= not(layer7_outputs(23)) or (layer7_outputs(4773));
    layer8_outputs(2054) <= (layer7_outputs(668)) or (layer7_outputs(1266));
    layer8_outputs(2055) <= not(layer7_outputs(2405));
    layer8_outputs(2056) <= (layer7_outputs(1880)) and not (layer7_outputs(3032));
    layer8_outputs(2057) <= layer7_outputs(5000);
    layer8_outputs(2058) <= not((layer7_outputs(4584)) xor (layer7_outputs(5039)));
    layer8_outputs(2059) <= not(layer7_outputs(4414));
    layer8_outputs(2060) <= not(layer7_outputs(811));
    layer8_outputs(2061) <= layer7_outputs(2145);
    layer8_outputs(2062) <= (layer7_outputs(3805)) xor (layer7_outputs(1526));
    layer8_outputs(2063) <= not((layer7_outputs(1300)) xor (layer7_outputs(399)));
    layer8_outputs(2064) <= layer7_outputs(2069);
    layer8_outputs(2065) <= (layer7_outputs(3191)) xor (layer7_outputs(3708));
    layer8_outputs(2066) <= (layer7_outputs(1374)) xor (layer7_outputs(78));
    layer8_outputs(2067) <= not(layer7_outputs(4390));
    layer8_outputs(2068) <= not(layer7_outputs(4843));
    layer8_outputs(2069) <= layer7_outputs(4277);
    layer8_outputs(2070) <= not((layer7_outputs(4651)) or (layer7_outputs(2552)));
    layer8_outputs(2071) <= not((layer7_outputs(552)) and (layer7_outputs(4486)));
    layer8_outputs(2072) <= layer7_outputs(4849);
    layer8_outputs(2073) <= not(layer7_outputs(494));
    layer8_outputs(2074) <= not(layer7_outputs(4216));
    layer8_outputs(2075) <= not((layer7_outputs(795)) or (layer7_outputs(3457)));
    layer8_outputs(2076) <= layer7_outputs(411);
    layer8_outputs(2077) <= not((layer7_outputs(2866)) xor (layer7_outputs(4773)));
    layer8_outputs(2078) <= layer7_outputs(1557);
    layer8_outputs(2079) <= (layer7_outputs(4497)) xor (layer7_outputs(3660));
    layer8_outputs(2080) <= not(layer7_outputs(3346));
    layer8_outputs(2081) <= layer7_outputs(3343);
    layer8_outputs(2082) <= not(layer7_outputs(3086));
    layer8_outputs(2083) <= not((layer7_outputs(5097)) and (layer7_outputs(4066)));
    layer8_outputs(2084) <= not(layer7_outputs(4544));
    layer8_outputs(2085) <= not((layer7_outputs(4482)) xor (layer7_outputs(3403)));
    layer8_outputs(2086) <= not((layer7_outputs(4420)) or (layer7_outputs(665)));
    layer8_outputs(2087) <= (layer7_outputs(523)) xor (layer7_outputs(205));
    layer8_outputs(2088) <= not((layer7_outputs(4668)) xor (layer7_outputs(1777)));
    layer8_outputs(2089) <= not(layer7_outputs(880)) or (layer7_outputs(1942));
    layer8_outputs(2090) <= not(layer7_outputs(4219));
    layer8_outputs(2091) <= (layer7_outputs(3174)) and (layer7_outputs(4601));
    layer8_outputs(2092) <= layer7_outputs(2249);
    layer8_outputs(2093) <= (layer7_outputs(20)) and not (layer7_outputs(4183));
    layer8_outputs(2094) <= not((layer7_outputs(380)) xor (layer7_outputs(5019)));
    layer8_outputs(2095) <= layer7_outputs(3621);
    layer8_outputs(2096) <= not(layer7_outputs(4169));
    layer8_outputs(2097) <= not((layer7_outputs(4669)) xor (layer7_outputs(4266)));
    layer8_outputs(2098) <= (layer7_outputs(4327)) and not (layer7_outputs(1776));
    layer8_outputs(2099) <= not(layer7_outputs(2261)) or (layer7_outputs(2576));
    layer8_outputs(2100) <= layer7_outputs(507);
    layer8_outputs(2101) <= not(layer7_outputs(3360));
    layer8_outputs(2102) <= not((layer7_outputs(844)) xor (layer7_outputs(846)));
    layer8_outputs(2103) <= not(layer7_outputs(2336));
    layer8_outputs(2104) <= layer7_outputs(4945);
    layer8_outputs(2105) <= not(layer7_outputs(2358)) or (layer7_outputs(681));
    layer8_outputs(2106) <= not((layer7_outputs(3848)) and (layer7_outputs(1203)));
    layer8_outputs(2107) <= not(layer7_outputs(1620));
    layer8_outputs(2108) <= (layer7_outputs(146)) and (layer7_outputs(1016));
    layer8_outputs(2109) <= not(layer7_outputs(4575)) or (layer7_outputs(4113));
    layer8_outputs(2110) <= (layer7_outputs(2041)) and not (layer7_outputs(4180));
    layer8_outputs(2111) <= not(layer7_outputs(2405));
    layer8_outputs(2112) <= (layer7_outputs(55)) xor (layer7_outputs(3610));
    layer8_outputs(2113) <= (layer7_outputs(4947)) and (layer7_outputs(4315));
    layer8_outputs(2114) <= not(layer7_outputs(4932)) or (layer7_outputs(308));
    layer8_outputs(2115) <= (layer7_outputs(3257)) or (layer7_outputs(3806));
    layer8_outputs(2116) <= layer7_outputs(4895);
    layer8_outputs(2117) <= not((layer7_outputs(837)) xor (layer7_outputs(287)));
    layer8_outputs(2118) <= not(layer7_outputs(4402));
    layer8_outputs(2119) <= layer7_outputs(3132);
    layer8_outputs(2120) <= (layer7_outputs(808)) xor (layer7_outputs(4895));
    layer8_outputs(2121) <= layer7_outputs(4376);
    layer8_outputs(2122) <= (layer7_outputs(5024)) xor (layer7_outputs(2901));
    layer8_outputs(2123) <= (layer7_outputs(1932)) xor (layer7_outputs(3732));
    layer8_outputs(2124) <= not(layer7_outputs(2903));
    layer8_outputs(2125) <= not((layer7_outputs(3865)) xor (layer7_outputs(4333)));
    layer8_outputs(2126) <= layer7_outputs(3332);
    layer8_outputs(2127) <= (layer7_outputs(1365)) or (layer7_outputs(241));
    layer8_outputs(2128) <= layer7_outputs(4833);
    layer8_outputs(2129) <= (layer7_outputs(4963)) and not (layer7_outputs(428));
    layer8_outputs(2130) <= layer7_outputs(4956);
    layer8_outputs(2131) <= layer7_outputs(3226);
    layer8_outputs(2132) <= layer7_outputs(288);
    layer8_outputs(2133) <= not((layer7_outputs(397)) xor (layer7_outputs(4804)));
    layer8_outputs(2134) <= not((layer7_outputs(1836)) and (layer7_outputs(3143)));
    layer8_outputs(2135) <= layer7_outputs(945);
    layer8_outputs(2136) <= not((layer7_outputs(1656)) and (layer7_outputs(3766)));
    layer8_outputs(2137) <= not(layer7_outputs(2429));
    layer8_outputs(2138) <= not(layer7_outputs(700));
    layer8_outputs(2139) <= not(layer7_outputs(4959)) or (layer7_outputs(1817));
    layer8_outputs(2140) <= layer7_outputs(2376);
    layer8_outputs(2141) <= not(layer7_outputs(4859));
    layer8_outputs(2142) <= (layer7_outputs(3629)) xor (layer7_outputs(3491));
    layer8_outputs(2143) <= not(layer7_outputs(691)) or (layer7_outputs(242));
    layer8_outputs(2144) <= (layer7_outputs(1647)) xor (layer7_outputs(777));
    layer8_outputs(2145) <= not(layer7_outputs(2051));
    layer8_outputs(2146) <= (layer7_outputs(4271)) xor (layer7_outputs(1042));
    layer8_outputs(2147) <= not((layer7_outputs(1891)) or (layer7_outputs(3937)));
    layer8_outputs(2148) <= not((layer7_outputs(3806)) and (layer7_outputs(3618)));
    layer8_outputs(2149) <= (layer7_outputs(638)) xor (layer7_outputs(3999));
    layer8_outputs(2150) <= not(layer7_outputs(4660));
    layer8_outputs(2151) <= not(layer7_outputs(213));
    layer8_outputs(2152) <= (layer7_outputs(1199)) xor (layer7_outputs(36));
    layer8_outputs(2153) <= not(layer7_outputs(512));
    layer8_outputs(2154) <= not(layer7_outputs(49));
    layer8_outputs(2155) <= not((layer7_outputs(3663)) xor (layer7_outputs(1889)));
    layer8_outputs(2156) <= layer7_outputs(2984);
    layer8_outputs(2157) <= not(layer7_outputs(4132));
    layer8_outputs(2158) <= (layer7_outputs(211)) xor (layer7_outputs(91));
    layer8_outputs(2159) <= not(layer7_outputs(4316));
    layer8_outputs(2160) <= not((layer7_outputs(415)) xor (layer7_outputs(1785)));
    layer8_outputs(2161) <= (layer7_outputs(2280)) and not (layer7_outputs(1815));
    layer8_outputs(2162) <= not((layer7_outputs(3830)) and (layer7_outputs(2253)));
    layer8_outputs(2163) <= (layer7_outputs(1521)) xor (layer7_outputs(993));
    layer8_outputs(2164) <= (layer7_outputs(2989)) xor (layer7_outputs(2187));
    layer8_outputs(2165) <= not((layer7_outputs(3096)) xor (layer7_outputs(4128)));
    layer8_outputs(2166) <= '0';
    layer8_outputs(2167) <= layer7_outputs(2949);
    layer8_outputs(2168) <= not(layer7_outputs(1175));
    layer8_outputs(2169) <= layer7_outputs(3395);
    layer8_outputs(2170) <= not((layer7_outputs(831)) xor (layer7_outputs(1183)));
    layer8_outputs(2171) <= (layer7_outputs(4211)) and not (layer7_outputs(3577));
    layer8_outputs(2172) <= layer7_outputs(4495);
    layer8_outputs(2173) <= not((layer7_outputs(40)) xor (layer7_outputs(3296)));
    layer8_outputs(2174) <= (layer7_outputs(3033)) and not (layer7_outputs(4242));
    layer8_outputs(2175) <= (layer7_outputs(1151)) and not (layer7_outputs(4778));
    layer8_outputs(2176) <= not(layer7_outputs(4841)) or (layer7_outputs(1333));
    layer8_outputs(2177) <= layer7_outputs(1273);
    layer8_outputs(2178) <= layer7_outputs(3019);
    layer8_outputs(2179) <= not(layer7_outputs(3768)) or (layer7_outputs(94));
    layer8_outputs(2180) <= layer7_outputs(82);
    layer8_outputs(2181) <= layer7_outputs(1402);
    layer8_outputs(2182) <= not(layer7_outputs(3376));
    layer8_outputs(2183) <= layer7_outputs(1565);
    layer8_outputs(2184) <= layer7_outputs(697);
    layer8_outputs(2185) <= not(layer7_outputs(2490));
    layer8_outputs(2186) <= (layer7_outputs(2082)) xor (layer7_outputs(926));
    layer8_outputs(2187) <= '0';
    layer8_outputs(2188) <= layer7_outputs(2073);
    layer8_outputs(2189) <= (layer7_outputs(288)) xor (layer7_outputs(2725));
    layer8_outputs(2190) <= (layer7_outputs(4796)) xor (layer7_outputs(741));
    layer8_outputs(2191) <= (layer7_outputs(501)) xor (layer7_outputs(1530));
    layer8_outputs(2192) <= layer7_outputs(3540);
    layer8_outputs(2193) <= layer7_outputs(1873);
    layer8_outputs(2194) <= (layer7_outputs(2521)) and not (layer7_outputs(3090));
    layer8_outputs(2195) <= not((layer7_outputs(3624)) xor (layer7_outputs(2987)));
    layer8_outputs(2196) <= layer7_outputs(2448);
    layer8_outputs(2197) <= not(layer7_outputs(1039));
    layer8_outputs(2198) <= (layer7_outputs(4176)) or (layer7_outputs(3538));
    layer8_outputs(2199) <= not(layer7_outputs(2185));
    layer8_outputs(2200) <= layer7_outputs(1462);
    layer8_outputs(2201) <= not((layer7_outputs(4907)) xor (layer7_outputs(895)));
    layer8_outputs(2202) <= layer7_outputs(4544);
    layer8_outputs(2203) <= (layer7_outputs(592)) or (layer7_outputs(2698));
    layer8_outputs(2204) <= not((layer7_outputs(915)) or (layer7_outputs(2481)));
    layer8_outputs(2205) <= not(layer7_outputs(24));
    layer8_outputs(2206) <= not(layer7_outputs(1426));
    layer8_outputs(2207) <= (layer7_outputs(4332)) and (layer7_outputs(3375));
    layer8_outputs(2208) <= layer7_outputs(624);
    layer8_outputs(2209) <= (layer7_outputs(1674)) xor (layer7_outputs(1071));
    layer8_outputs(2210) <= not(layer7_outputs(4038));
    layer8_outputs(2211) <= layer7_outputs(2955);
    layer8_outputs(2212) <= layer7_outputs(490);
    layer8_outputs(2213) <= layer7_outputs(3559);
    layer8_outputs(2214) <= layer7_outputs(1342);
    layer8_outputs(2215) <= (layer7_outputs(3780)) and not (layer7_outputs(2660));
    layer8_outputs(2216) <= (layer7_outputs(4490)) or (layer7_outputs(1103));
    layer8_outputs(2217) <= (layer7_outputs(4643)) xor (layer7_outputs(2830));
    layer8_outputs(2218) <= (layer7_outputs(0)) xor (layer7_outputs(4151));
    layer8_outputs(2219) <= (layer7_outputs(3112)) and not (layer7_outputs(720));
    layer8_outputs(2220) <= (layer7_outputs(1595)) xor (layer7_outputs(538));
    layer8_outputs(2221) <= layer7_outputs(2427);
    layer8_outputs(2222) <= (layer7_outputs(3631)) xor (layer7_outputs(4921));
    layer8_outputs(2223) <= (layer7_outputs(2540)) and (layer7_outputs(1722));
    layer8_outputs(2224) <= (layer7_outputs(4559)) and not (layer7_outputs(883));
    layer8_outputs(2225) <= not(layer7_outputs(2467));
    layer8_outputs(2226) <= not((layer7_outputs(1774)) xor (layer7_outputs(4305)));
    layer8_outputs(2227) <= (layer7_outputs(2233)) xor (layer7_outputs(3104));
    layer8_outputs(2228) <= layer7_outputs(4224);
    layer8_outputs(2229) <= (layer7_outputs(866)) and not (layer7_outputs(4400));
    layer8_outputs(2230) <= not(layer7_outputs(1439));
    layer8_outputs(2231) <= layer7_outputs(3382);
    layer8_outputs(2232) <= layer7_outputs(3309);
    layer8_outputs(2233) <= (layer7_outputs(1089)) or (layer7_outputs(834));
    layer8_outputs(2234) <= (layer7_outputs(3304)) and (layer7_outputs(1245));
    layer8_outputs(2235) <= '1';
    layer8_outputs(2236) <= not(layer7_outputs(1258));
    layer8_outputs(2237) <= layer7_outputs(4624);
    layer8_outputs(2238) <= layer7_outputs(478);
    layer8_outputs(2239) <= layer7_outputs(652);
    layer8_outputs(2240) <= layer7_outputs(3021);
    layer8_outputs(2241) <= not(layer7_outputs(4133));
    layer8_outputs(2242) <= (layer7_outputs(653)) and (layer7_outputs(489));
    layer8_outputs(2243) <= layer7_outputs(3265);
    layer8_outputs(2244) <= not(layer7_outputs(1813));
    layer8_outputs(2245) <= not(layer7_outputs(3408));
    layer8_outputs(2246) <= not((layer7_outputs(422)) xor (layer7_outputs(903)));
    layer8_outputs(2247) <= (layer7_outputs(3755)) and not (layer7_outputs(4808));
    layer8_outputs(2248) <= not(layer7_outputs(1155));
    layer8_outputs(2249) <= not((layer7_outputs(45)) xor (layer7_outputs(2944)));
    layer8_outputs(2250) <= not(layer7_outputs(3667));
    layer8_outputs(2251) <= layer7_outputs(1254);
    layer8_outputs(2252) <= layer7_outputs(2785);
    layer8_outputs(2253) <= (layer7_outputs(5019)) xor (layer7_outputs(751));
    layer8_outputs(2254) <= layer7_outputs(3690);
    layer8_outputs(2255) <= layer7_outputs(2794);
    layer8_outputs(2256) <= layer7_outputs(2391);
    layer8_outputs(2257) <= layer7_outputs(664);
    layer8_outputs(2258) <= (layer7_outputs(1216)) xor (layer7_outputs(919));
    layer8_outputs(2259) <= (layer7_outputs(3021)) and not (layer7_outputs(3930));
    layer8_outputs(2260) <= layer7_outputs(4051);
    layer8_outputs(2261) <= not((layer7_outputs(2440)) or (layer7_outputs(4003)));
    layer8_outputs(2262) <= (layer7_outputs(472)) xor (layer7_outputs(2741));
    layer8_outputs(2263) <= not(layer7_outputs(3424));
    layer8_outputs(2264) <= (layer7_outputs(4005)) xor (layer7_outputs(455));
    layer8_outputs(2265) <= layer7_outputs(1640);
    layer8_outputs(2266) <= (layer7_outputs(64)) xor (layer7_outputs(3190));
    layer8_outputs(2267) <= not((layer7_outputs(3522)) xor (layer7_outputs(3805)));
    layer8_outputs(2268) <= layer7_outputs(4336);
    layer8_outputs(2269) <= not((layer7_outputs(3221)) and (layer7_outputs(2977)));
    layer8_outputs(2270) <= not(layer7_outputs(4665));
    layer8_outputs(2271) <= not(layer7_outputs(561));
    layer8_outputs(2272) <= layer7_outputs(4158);
    layer8_outputs(2273) <= not(layer7_outputs(1997));
    layer8_outputs(2274) <= not(layer7_outputs(1800));
    layer8_outputs(2275) <= layer7_outputs(3720);
    layer8_outputs(2276) <= not((layer7_outputs(4368)) xor (layer7_outputs(957)));
    layer8_outputs(2277) <= not(layer7_outputs(207)) or (layer7_outputs(4858));
    layer8_outputs(2278) <= not((layer7_outputs(4875)) xor (layer7_outputs(1888)));
    layer8_outputs(2279) <= not(layer7_outputs(4164));
    layer8_outputs(2280) <= layer7_outputs(2154);
    layer8_outputs(2281) <= layer7_outputs(2558);
    layer8_outputs(2282) <= not((layer7_outputs(4476)) and (layer7_outputs(2529)));
    layer8_outputs(2283) <= (layer7_outputs(4722)) xor (layer7_outputs(2029));
    layer8_outputs(2284) <= not(layer7_outputs(579));
    layer8_outputs(2285) <= (layer7_outputs(1137)) xor (layer7_outputs(4298));
    layer8_outputs(2286) <= (layer7_outputs(3971)) and (layer7_outputs(4352));
    layer8_outputs(2287) <= (layer7_outputs(3916)) or (layer7_outputs(4709));
    layer8_outputs(2288) <= not(layer7_outputs(1717)) or (layer7_outputs(4658));
    layer8_outputs(2289) <= not(layer7_outputs(1));
    layer8_outputs(2290) <= layer7_outputs(2993);
    layer8_outputs(2291) <= (layer7_outputs(3808)) and (layer7_outputs(4968));
    layer8_outputs(2292) <= not(layer7_outputs(4615));
    layer8_outputs(2293) <= not((layer7_outputs(772)) and (layer7_outputs(3883)));
    layer8_outputs(2294) <= layer7_outputs(2779);
    layer8_outputs(2295) <= not(layer7_outputs(4704));
    layer8_outputs(2296) <= layer7_outputs(2686);
    layer8_outputs(2297) <= not(layer7_outputs(1333));
    layer8_outputs(2298) <= not(layer7_outputs(5056));
    layer8_outputs(2299) <= not(layer7_outputs(510)) or (layer7_outputs(1619));
    layer8_outputs(2300) <= layer7_outputs(2132);
    layer8_outputs(2301) <= not(layer7_outputs(128)) or (layer7_outputs(5033));
    layer8_outputs(2302) <= (layer7_outputs(3984)) and not (layer7_outputs(3777));
    layer8_outputs(2303) <= not((layer7_outputs(283)) xor (layer7_outputs(1623)));
    layer8_outputs(2304) <= layer7_outputs(2724);
    layer8_outputs(2305) <= not(layer7_outputs(3463));
    layer8_outputs(2306) <= layer7_outputs(2333);
    layer8_outputs(2307) <= not((layer7_outputs(749)) xor (layer7_outputs(2523)));
    layer8_outputs(2308) <= not((layer7_outputs(1491)) xor (layer7_outputs(2515)));
    layer8_outputs(2309) <= not((layer7_outputs(835)) and (layer7_outputs(597)));
    layer8_outputs(2310) <= not(layer7_outputs(4165));
    layer8_outputs(2311) <= not((layer7_outputs(2320)) or (layer7_outputs(1768)));
    layer8_outputs(2312) <= not(layer7_outputs(479));
    layer8_outputs(2313) <= (layer7_outputs(2499)) and not (layer7_outputs(3262));
    layer8_outputs(2314) <= not((layer7_outputs(1472)) or (layer7_outputs(1666)));
    layer8_outputs(2315) <= not(layer7_outputs(276));
    layer8_outputs(2316) <= not(layer7_outputs(1091));
    layer8_outputs(2317) <= layer7_outputs(3933);
    layer8_outputs(2318) <= not(layer7_outputs(3083)) or (layer7_outputs(1310));
    layer8_outputs(2319) <= not((layer7_outputs(4345)) xor (layer7_outputs(85)));
    layer8_outputs(2320) <= (layer7_outputs(1188)) or (layer7_outputs(559));
    layer8_outputs(2321) <= (layer7_outputs(3288)) and not (layer7_outputs(2775));
    layer8_outputs(2322) <= layer7_outputs(4103);
    layer8_outputs(2323) <= (layer7_outputs(2164)) and not (layer7_outputs(4358));
    layer8_outputs(2324) <= (layer7_outputs(3293)) or (layer7_outputs(2861));
    layer8_outputs(2325) <= layer7_outputs(954);
    layer8_outputs(2326) <= layer7_outputs(5114);
    layer8_outputs(2327) <= not(layer7_outputs(2381)) or (layer7_outputs(201));
    layer8_outputs(2328) <= not((layer7_outputs(1956)) xor (layer7_outputs(4514)));
    layer8_outputs(2329) <= (layer7_outputs(2056)) xor (layer7_outputs(4558));
    layer8_outputs(2330) <= not((layer7_outputs(2274)) and (layer7_outputs(2745)));
    layer8_outputs(2331) <= (layer7_outputs(1942)) and not (layer7_outputs(406));
    layer8_outputs(2332) <= (layer7_outputs(1730)) or (layer7_outputs(3399));
    layer8_outputs(2333) <= (layer7_outputs(2247)) and not (layer7_outputs(2613));
    layer8_outputs(2334) <= not(layer7_outputs(771));
    layer8_outputs(2335) <= not(layer7_outputs(2416));
    layer8_outputs(2336) <= (layer7_outputs(5053)) and not (layer7_outputs(382));
    layer8_outputs(2337) <= layer7_outputs(3189);
    layer8_outputs(2338) <= (layer7_outputs(2452)) and (layer7_outputs(1901));
    layer8_outputs(2339) <= layer7_outputs(2125);
    layer8_outputs(2340) <= (layer7_outputs(98)) xor (layer7_outputs(4234));
    layer8_outputs(2341) <= not((layer7_outputs(4054)) or (layer7_outputs(2996)));
    layer8_outputs(2342) <= layer7_outputs(1223);
    layer8_outputs(2343) <= layer7_outputs(4634);
    layer8_outputs(2344) <= layer7_outputs(394);
    layer8_outputs(2345) <= (layer7_outputs(349)) xor (layer7_outputs(2185));
    layer8_outputs(2346) <= not(layer7_outputs(1948));
    layer8_outputs(2347) <= not(layer7_outputs(1282)) or (layer7_outputs(4027));
    layer8_outputs(2348) <= not((layer7_outputs(4268)) xor (layer7_outputs(2179)));
    layer8_outputs(2349) <= not((layer7_outputs(1713)) xor (layer7_outputs(4739)));
    layer8_outputs(2350) <= (layer7_outputs(3482)) and (layer7_outputs(4815));
    layer8_outputs(2351) <= not((layer7_outputs(4713)) xor (layer7_outputs(1659)));
    layer8_outputs(2352) <= not(layer7_outputs(4364));
    layer8_outputs(2353) <= not(layer7_outputs(941));
    layer8_outputs(2354) <= layer7_outputs(2418);
    layer8_outputs(2355) <= not((layer7_outputs(3206)) or (layer7_outputs(1848)));
    layer8_outputs(2356) <= not(layer7_outputs(3148));
    layer8_outputs(2357) <= (layer7_outputs(76)) and not (layer7_outputs(181));
    layer8_outputs(2358) <= layer7_outputs(4341);
    layer8_outputs(2359) <= layer7_outputs(626);
    layer8_outputs(2360) <= (layer7_outputs(2313)) and not (layer7_outputs(954));
    layer8_outputs(2361) <= not((layer7_outputs(4737)) or (layer7_outputs(2537)));
    layer8_outputs(2362) <= not(layer7_outputs(3251));
    layer8_outputs(2363) <= (layer7_outputs(4338)) and (layer7_outputs(1538));
    layer8_outputs(2364) <= not(layer7_outputs(4166));
    layer8_outputs(2365) <= not(layer7_outputs(1577));
    layer8_outputs(2366) <= layer7_outputs(5076);
    layer8_outputs(2367) <= not(layer7_outputs(2321));
    layer8_outputs(2368) <= layer7_outputs(2044);
    layer8_outputs(2369) <= not(layer7_outputs(737));
    layer8_outputs(2370) <= layer7_outputs(3574);
    layer8_outputs(2371) <= layer7_outputs(1194);
    layer8_outputs(2372) <= layer7_outputs(2780);
    layer8_outputs(2373) <= (layer7_outputs(2990)) xor (layer7_outputs(3124));
    layer8_outputs(2374) <= layer7_outputs(4063);
    layer8_outputs(2375) <= not(layer7_outputs(1081));
    layer8_outputs(2376) <= (layer7_outputs(544)) or (layer7_outputs(1832));
    layer8_outputs(2377) <= not((layer7_outputs(701)) and (layer7_outputs(1095)));
    layer8_outputs(2378) <= not(layer7_outputs(135)) or (layer7_outputs(2964));
    layer8_outputs(2379) <= layer7_outputs(2411);
    layer8_outputs(2380) <= '1';
    layer8_outputs(2381) <= not(layer7_outputs(4198));
    layer8_outputs(2382) <= (layer7_outputs(316)) and (layer7_outputs(4399));
    layer8_outputs(2383) <= not(layer7_outputs(4008));
    layer8_outputs(2384) <= not((layer7_outputs(2577)) xor (layer7_outputs(214)));
    layer8_outputs(2385) <= layer7_outputs(4477);
    layer8_outputs(2386) <= (layer7_outputs(4253)) and not (layer7_outputs(3516));
    layer8_outputs(2387) <= not(layer7_outputs(519));
    layer8_outputs(2388) <= (layer7_outputs(5099)) or (layer7_outputs(1427));
    layer8_outputs(2389) <= not(layer7_outputs(3278));
    layer8_outputs(2390) <= layer7_outputs(1144);
    layer8_outputs(2391) <= not(layer7_outputs(2020));
    layer8_outputs(2392) <= (layer7_outputs(2537)) and not (layer7_outputs(2543));
    layer8_outputs(2393) <= not(layer7_outputs(4552));
    layer8_outputs(2394) <= not(layer7_outputs(2232));
    layer8_outputs(2395) <= not(layer7_outputs(3285));
    layer8_outputs(2396) <= not((layer7_outputs(124)) and (layer7_outputs(4708)));
    layer8_outputs(2397) <= (layer7_outputs(4964)) xor (layer7_outputs(2113));
    layer8_outputs(2398) <= (layer7_outputs(4536)) or (layer7_outputs(116));
    layer8_outputs(2399) <= (layer7_outputs(3942)) and not (layer7_outputs(712));
    layer8_outputs(2400) <= layer7_outputs(680);
    layer8_outputs(2401) <= not((layer7_outputs(763)) xor (layer7_outputs(3070)));
    layer8_outputs(2402) <= layer7_outputs(1499);
    layer8_outputs(2403) <= not((layer7_outputs(2446)) xor (layer7_outputs(3598)));
    layer8_outputs(2404) <= not(layer7_outputs(1598)) or (layer7_outputs(3455));
    layer8_outputs(2405) <= not((layer7_outputs(4572)) xor (layer7_outputs(2717)));
    layer8_outputs(2406) <= not((layer7_outputs(3188)) xor (layer7_outputs(2504)));
    layer8_outputs(2407) <= not(layer7_outputs(1651));
    layer8_outputs(2408) <= not(layer7_outputs(4758));
    layer8_outputs(2409) <= not((layer7_outputs(1775)) xor (layer7_outputs(1292)));
    layer8_outputs(2410) <= (layer7_outputs(2090)) and (layer7_outputs(4702));
    layer8_outputs(2411) <= layer7_outputs(3144);
    layer8_outputs(2412) <= layer7_outputs(2904);
    layer8_outputs(2413) <= layer7_outputs(2226);
    layer8_outputs(2414) <= not(layer7_outputs(4714));
    layer8_outputs(2415) <= layer7_outputs(157);
    layer8_outputs(2416) <= layer7_outputs(2740);
    layer8_outputs(2417) <= not(layer7_outputs(4980)) or (layer7_outputs(3767));
    layer8_outputs(2418) <= not(layer7_outputs(1672)) or (layer7_outputs(775));
    layer8_outputs(2419) <= (layer7_outputs(2030)) xor (layer7_outputs(4903));
    layer8_outputs(2420) <= layer7_outputs(1416);
    layer8_outputs(2421) <= not((layer7_outputs(2813)) xor (layer7_outputs(2885)));
    layer8_outputs(2422) <= not((layer7_outputs(3744)) xor (layer7_outputs(3147)));
    layer8_outputs(2423) <= (layer7_outputs(3988)) xor (layer7_outputs(304));
    layer8_outputs(2424) <= not((layer7_outputs(3105)) xor (layer7_outputs(3466)));
    layer8_outputs(2425) <= not(layer7_outputs(2054));
    layer8_outputs(2426) <= layer7_outputs(2568);
    layer8_outputs(2427) <= not((layer7_outputs(5066)) or (layer7_outputs(4426)));
    layer8_outputs(2428) <= not(layer7_outputs(1939));
    layer8_outputs(2429) <= not(layer7_outputs(1074));
    layer8_outputs(2430) <= not(layer7_outputs(4186));
    layer8_outputs(2431) <= (layer7_outputs(3879)) xor (layer7_outputs(2926));
    layer8_outputs(2432) <= (layer7_outputs(2991)) or (layer7_outputs(3891));
    layer8_outputs(2433) <= not(layer7_outputs(2374));
    layer8_outputs(2434) <= (layer7_outputs(4236)) and not (layer7_outputs(656));
    layer8_outputs(2435) <= not(layer7_outputs(2853)) or (layer7_outputs(1845));
    layer8_outputs(2436) <= layer7_outputs(2476);
    layer8_outputs(2437) <= layer7_outputs(78);
    layer8_outputs(2438) <= not((layer7_outputs(3738)) xor (layer7_outputs(1357)));
    layer8_outputs(2439) <= (layer7_outputs(1000)) or (layer7_outputs(905));
    layer8_outputs(2440) <= (layer7_outputs(1806)) and not (layer7_outputs(4684));
    layer8_outputs(2441) <= not((layer7_outputs(1381)) xor (layer7_outputs(2174)));
    layer8_outputs(2442) <= (layer7_outputs(3695)) and not (layer7_outputs(150));
    layer8_outputs(2443) <= not(layer7_outputs(2685));
    layer8_outputs(2444) <= layer7_outputs(4131);
    layer8_outputs(2445) <= not((layer7_outputs(3078)) xor (layer7_outputs(3671)));
    layer8_outputs(2446) <= not(layer7_outputs(850));
    layer8_outputs(2447) <= not(layer7_outputs(4945));
    layer8_outputs(2448) <= not((layer7_outputs(2401)) and (layer7_outputs(2345)));
    layer8_outputs(2449) <= layer7_outputs(4190);
    layer8_outputs(2450) <= not(layer7_outputs(4838));
    layer8_outputs(2451) <= (layer7_outputs(3214)) xor (layer7_outputs(3371));
    layer8_outputs(2452) <= not(layer7_outputs(2151));
    layer8_outputs(2453) <= not((layer7_outputs(3858)) xor (layer7_outputs(3863)));
    layer8_outputs(2454) <= (layer7_outputs(814)) xor (layer7_outputs(1056));
    layer8_outputs(2455) <= (layer7_outputs(540)) and not (layer7_outputs(1423));
    layer8_outputs(2456) <= '1';
    layer8_outputs(2457) <= layer7_outputs(230);
    layer8_outputs(2458) <= (layer7_outputs(1621)) xor (layer7_outputs(1085));
    layer8_outputs(2459) <= layer7_outputs(3341);
    layer8_outputs(2460) <= layer7_outputs(684);
    layer8_outputs(2461) <= not((layer7_outputs(3327)) and (layer7_outputs(2727)));
    layer8_outputs(2462) <= (layer7_outputs(742)) xor (layer7_outputs(3443));
    layer8_outputs(2463) <= (layer7_outputs(3498)) xor (layer7_outputs(2190));
    layer8_outputs(2464) <= not(layer7_outputs(2206)) or (layer7_outputs(2305));
    layer8_outputs(2465) <= not(layer7_outputs(3790)) or (layer7_outputs(2868));
    layer8_outputs(2466) <= not(layer7_outputs(389));
    layer8_outputs(2467) <= layer7_outputs(4682);
    layer8_outputs(2468) <= not((layer7_outputs(2328)) or (layer7_outputs(2071)));
    layer8_outputs(2469) <= layer7_outputs(3106);
    layer8_outputs(2470) <= layer7_outputs(2158);
    layer8_outputs(2471) <= layer7_outputs(3747);
    layer8_outputs(2472) <= layer7_outputs(4214);
    layer8_outputs(2473) <= not((layer7_outputs(609)) or (layer7_outputs(3454)));
    layer8_outputs(2474) <= (layer7_outputs(4594)) and (layer7_outputs(1352));
    layer8_outputs(2475) <= layer7_outputs(4879);
    layer8_outputs(2476) <= layer7_outputs(3472);
    layer8_outputs(2477) <= (layer7_outputs(3687)) and not (layer7_outputs(2193));
    layer8_outputs(2478) <= not(layer7_outputs(4073)) or (layer7_outputs(922));
    layer8_outputs(2479) <= not((layer7_outputs(4705)) xor (layer7_outputs(843)));
    layer8_outputs(2480) <= not((layer7_outputs(4672)) and (layer7_outputs(804)));
    layer8_outputs(2481) <= (layer7_outputs(1855)) xor (layer7_outputs(4473));
    layer8_outputs(2482) <= (layer7_outputs(569)) or (layer7_outputs(3888));
    layer8_outputs(2483) <= (layer7_outputs(1084)) and not (layer7_outputs(3587));
    layer8_outputs(2484) <= not(layer7_outputs(114));
    layer8_outputs(2485) <= (layer7_outputs(144)) xor (layer7_outputs(3665));
    layer8_outputs(2486) <= layer7_outputs(3264);
    layer8_outputs(2487) <= layer7_outputs(1378);
    layer8_outputs(2488) <= '1';
    layer8_outputs(2489) <= not((layer7_outputs(2878)) or (layer7_outputs(864)));
    layer8_outputs(2490) <= not(layer7_outputs(2148));
    layer8_outputs(2491) <= (layer7_outputs(2731)) xor (layer7_outputs(4301));
    layer8_outputs(2492) <= not(layer7_outputs(735));
    layer8_outputs(2493) <= layer7_outputs(3036);
    layer8_outputs(2494) <= (layer7_outputs(294)) xor (layer7_outputs(688));
    layer8_outputs(2495) <= not((layer7_outputs(482)) and (layer7_outputs(2334)));
    layer8_outputs(2496) <= not(layer7_outputs(3716));
    layer8_outputs(2497) <= (layer7_outputs(3347)) and not (layer7_outputs(2444));
    layer8_outputs(2498) <= not((layer7_outputs(4116)) or (layer7_outputs(3474)));
    layer8_outputs(2499) <= not(layer7_outputs(4484)) or (layer7_outputs(2));
    layer8_outputs(2500) <= not(layer7_outputs(4027)) or (layer7_outputs(4269));
    layer8_outputs(2501) <= layer7_outputs(3268);
    layer8_outputs(2502) <= not(layer7_outputs(3129));
    layer8_outputs(2503) <= not(layer7_outputs(2125));
    layer8_outputs(2504) <= not((layer7_outputs(4204)) or (layer7_outputs(4947)));
    layer8_outputs(2505) <= layer7_outputs(2580);
    layer8_outputs(2506) <= (layer7_outputs(4385)) and not (layer7_outputs(761));
    layer8_outputs(2507) <= layer7_outputs(4710);
    layer8_outputs(2508) <= not(layer7_outputs(3367)) or (layer7_outputs(3978));
    layer8_outputs(2509) <= layer7_outputs(4243);
    layer8_outputs(2510) <= not((layer7_outputs(3648)) and (layer7_outputs(1125)));
    layer8_outputs(2511) <= layer7_outputs(4818);
    layer8_outputs(2512) <= (layer7_outputs(172)) xor (layer7_outputs(989));
    layer8_outputs(2513) <= layer7_outputs(1622);
    layer8_outputs(2514) <= (layer7_outputs(275)) and not (layer7_outputs(256));
    layer8_outputs(2515) <= not(layer7_outputs(1880)) or (layer7_outputs(3010));
    layer8_outputs(2516) <= (layer7_outputs(459)) xor (layer7_outputs(3880));
    layer8_outputs(2517) <= not((layer7_outputs(4626)) xor (layer7_outputs(946)));
    layer8_outputs(2518) <= not(layer7_outputs(1319));
    layer8_outputs(2519) <= layer7_outputs(960);
    layer8_outputs(2520) <= not((layer7_outputs(1954)) and (layer7_outputs(4071)));
    layer8_outputs(2521) <= not(layer7_outputs(3158));
    layer8_outputs(2522) <= layer7_outputs(1046);
    layer8_outputs(2523) <= (layer7_outputs(133)) xor (layer7_outputs(634));
    layer8_outputs(2524) <= (layer7_outputs(267)) and not (layer7_outputs(278));
    layer8_outputs(2525) <= not(layer7_outputs(77));
    layer8_outputs(2526) <= (layer7_outputs(991)) and not (layer7_outputs(3567));
    layer8_outputs(2527) <= not((layer7_outputs(522)) xor (layer7_outputs(3931)));
    layer8_outputs(2528) <= (layer7_outputs(1352)) and not (layer7_outputs(3961));
    layer8_outputs(2529) <= (layer7_outputs(5016)) and (layer7_outputs(724));
    layer8_outputs(2530) <= not(layer7_outputs(3995));
    layer8_outputs(2531) <= not((layer7_outputs(193)) xor (layer7_outputs(1288)));
    layer8_outputs(2532) <= not((layer7_outputs(4384)) or (layer7_outputs(3919)));
    layer8_outputs(2533) <= layer7_outputs(3414);
    layer8_outputs(2534) <= (layer7_outputs(3676)) and not (layer7_outputs(4510));
    layer8_outputs(2535) <= (layer7_outputs(1480)) xor (layer7_outputs(1650));
    layer8_outputs(2536) <= not(layer7_outputs(557));
    layer8_outputs(2537) <= (layer7_outputs(2713)) xor (layer7_outputs(229));
    layer8_outputs(2538) <= not(layer7_outputs(5018)) or (layer7_outputs(1372));
    layer8_outputs(2539) <= not(layer7_outputs(4182));
    layer8_outputs(2540) <= '1';
    layer8_outputs(2541) <= (layer7_outputs(3789)) and (layer7_outputs(4343));
    layer8_outputs(2542) <= not(layer7_outputs(1335));
    layer8_outputs(2543) <= not(layer7_outputs(5084));
    layer8_outputs(2544) <= layer7_outputs(3559);
    layer8_outputs(2545) <= (layer7_outputs(5010)) xor (layer7_outputs(4127));
    layer8_outputs(2546) <= layer7_outputs(4840);
    layer8_outputs(2547) <= not(layer7_outputs(2780));
    layer8_outputs(2548) <= not(layer7_outputs(4267)) or (layer7_outputs(2014));
    layer8_outputs(2549) <= not((layer7_outputs(2118)) and (layer7_outputs(2790)));
    layer8_outputs(2550) <= layer7_outputs(3487);
    layer8_outputs(2551) <= not((layer7_outputs(3388)) xor (layer7_outputs(2331)));
    layer8_outputs(2552) <= not(layer7_outputs(4587)) or (layer7_outputs(1225));
    layer8_outputs(2553) <= not(layer7_outputs(3895));
    layer8_outputs(2554) <= not(layer7_outputs(1439)) or (layer7_outputs(2933));
    layer8_outputs(2555) <= not((layer7_outputs(1638)) xor (layer7_outputs(2056)));
    layer8_outputs(2556) <= not(layer7_outputs(734)) or (layer7_outputs(1196));
    layer8_outputs(2557) <= not((layer7_outputs(2010)) xor (layer7_outputs(4513)));
    layer8_outputs(2558) <= (layer7_outputs(3792)) xor (layer7_outputs(4440));
    layer8_outputs(2559) <= (layer7_outputs(788)) xor (layer7_outputs(3956));
    layer8_outputs(2560) <= layer7_outputs(863);
    layer8_outputs(2561) <= layer7_outputs(3701);
    layer8_outputs(2562) <= (layer7_outputs(4365)) xor (layer7_outputs(16));
    layer8_outputs(2563) <= layer7_outputs(3645);
    layer8_outputs(2564) <= not((layer7_outputs(4703)) xor (layer7_outputs(2101)));
    layer8_outputs(2565) <= not(layer7_outputs(4757));
    layer8_outputs(2566) <= (layer7_outputs(2810)) xor (layer7_outputs(4612));
    layer8_outputs(2567) <= not(layer7_outputs(2067));
    layer8_outputs(2568) <= not(layer7_outputs(2831));
    layer8_outputs(2569) <= layer7_outputs(5088);
    layer8_outputs(2570) <= not(layer7_outputs(217));
    layer8_outputs(2571) <= not((layer7_outputs(2066)) xor (layer7_outputs(3056)));
    layer8_outputs(2572) <= (layer7_outputs(1863)) and not (layer7_outputs(5084));
    layer8_outputs(2573) <= not(layer7_outputs(2526));
    layer8_outputs(2574) <= layer7_outputs(4033);
    layer8_outputs(2575) <= not(layer7_outputs(3199));
    layer8_outputs(2576) <= layer7_outputs(1343);
    layer8_outputs(2577) <= not(layer7_outputs(581)) or (layer7_outputs(4275));
    layer8_outputs(2578) <= not(layer7_outputs(534));
    layer8_outputs(2579) <= (layer7_outputs(4041)) xor (layer7_outputs(1733));
    layer8_outputs(2580) <= layer7_outputs(3200);
    layer8_outputs(2581) <= (layer7_outputs(547)) xor (layer7_outputs(2203));
    layer8_outputs(2582) <= layer7_outputs(4039);
    layer8_outputs(2583) <= not(layer7_outputs(917));
    layer8_outputs(2584) <= not((layer7_outputs(1748)) and (layer7_outputs(2584)));
    layer8_outputs(2585) <= not(layer7_outputs(3590));
    layer8_outputs(2586) <= not(layer7_outputs(1085)) or (layer7_outputs(2018));
    layer8_outputs(2587) <= not(layer7_outputs(1394));
    layer8_outputs(2588) <= not(layer7_outputs(808));
    layer8_outputs(2589) <= not((layer7_outputs(2334)) and (layer7_outputs(2509)));
    layer8_outputs(2590) <= not(layer7_outputs(3305));
    layer8_outputs(2591) <= not((layer7_outputs(821)) and (layer7_outputs(4187)));
    layer8_outputs(2592) <= (layer7_outputs(4745)) and (layer7_outputs(987));
    layer8_outputs(2593) <= not(layer7_outputs(3614));
    layer8_outputs(2594) <= not((layer7_outputs(4321)) or (layer7_outputs(2246)));
    layer8_outputs(2595) <= layer7_outputs(2623);
    layer8_outputs(2596) <= not(layer7_outputs(5));
    layer8_outputs(2597) <= not(layer7_outputs(4949)) or (layer7_outputs(3399));
    layer8_outputs(2598) <= not(layer7_outputs(3936)) or (layer7_outputs(985));
    layer8_outputs(2599) <= layer7_outputs(1503);
    layer8_outputs(2600) <= (layer7_outputs(3694)) or (layer7_outputs(1120));
    layer8_outputs(2601) <= layer7_outputs(716);
    layer8_outputs(2602) <= (layer7_outputs(3725)) xor (layer7_outputs(1034));
    layer8_outputs(2603) <= not(layer7_outputs(1985));
    layer8_outputs(2604) <= layer7_outputs(2277);
    layer8_outputs(2605) <= not((layer7_outputs(3230)) and (layer7_outputs(192)));
    layer8_outputs(2606) <= not(layer7_outputs(1968));
    layer8_outputs(2607) <= layer7_outputs(1230);
    layer8_outputs(2608) <= not(layer7_outputs(2063));
    layer8_outputs(2609) <= (layer7_outputs(663)) and not (layer7_outputs(3518));
    layer8_outputs(2610) <= (layer7_outputs(1839)) and (layer7_outputs(2594));
    layer8_outputs(2611) <= layer7_outputs(1973);
    layer8_outputs(2612) <= not(layer7_outputs(2067));
    layer8_outputs(2613) <= layer7_outputs(336);
    layer8_outputs(2614) <= not((layer7_outputs(5007)) or (layer7_outputs(4145)));
    layer8_outputs(2615) <= not(layer7_outputs(3162));
    layer8_outputs(2616) <= not((layer7_outputs(3704)) xor (layer7_outputs(2731)));
    layer8_outputs(2617) <= (layer7_outputs(3576)) and (layer7_outputs(4835));
    layer8_outputs(2618) <= not(layer7_outputs(1474));
    layer8_outputs(2619) <= (layer7_outputs(345)) xor (layer7_outputs(3316));
    layer8_outputs(2620) <= layer7_outputs(1172);
    layer8_outputs(2621) <= not(layer7_outputs(3629));
    layer8_outputs(2622) <= not((layer7_outputs(4389)) or (layer7_outputs(142)));
    layer8_outputs(2623) <= not(layer7_outputs(3688));
    layer8_outputs(2624) <= not((layer7_outputs(2645)) and (layer7_outputs(5113)));
    layer8_outputs(2625) <= not(layer7_outputs(2542));
    layer8_outputs(2626) <= not((layer7_outputs(3601)) xor (layer7_outputs(4653)));
    layer8_outputs(2627) <= not(layer7_outputs(8));
    layer8_outputs(2628) <= not(layer7_outputs(1543)) or (layer7_outputs(3349));
    layer8_outputs(2629) <= not(layer7_outputs(368));
    layer8_outputs(2630) <= not((layer7_outputs(2725)) xor (layer7_outputs(1604)));
    layer8_outputs(2631) <= not(layer7_outputs(279));
    layer8_outputs(2632) <= (layer7_outputs(5075)) xor (layer7_outputs(1991));
    layer8_outputs(2633) <= not(layer7_outputs(2512)) or (layer7_outputs(225));
    layer8_outputs(2634) <= not(layer7_outputs(4903));
    layer8_outputs(2635) <= not(layer7_outputs(1632)) or (layer7_outputs(442));
    layer8_outputs(2636) <= not(layer7_outputs(1021)) or (layer7_outputs(1786));
    layer8_outputs(2637) <= (layer7_outputs(1136)) and not (layer7_outputs(449));
    layer8_outputs(2638) <= not(layer7_outputs(657));
    layer8_outputs(2639) <= layer7_outputs(3729);
    layer8_outputs(2640) <= layer7_outputs(3582);
    layer8_outputs(2641) <= (layer7_outputs(2638)) and (layer7_outputs(978));
    layer8_outputs(2642) <= not((layer7_outputs(1815)) and (layer7_outputs(1017)));
    layer8_outputs(2643) <= not((layer7_outputs(4115)) and (layer7_outputs(2634)));
    layer8_outputs(2644) <= layer7_outputs(5108);
    layer8_outputs(2645) <= layer7_outputs(1010);
    layer8_outputs(2646) <= not(layer7_outputs(3193));
    layer8_outputs(2647) <= not((layer7_outputs(632)) xor (layer7_outputs(3378)));
    layer8_outputs(2648) <= not(layer7_outputs(475));
    layer8_outputs(2649) <= not(layer7_outputs(4815));
    layer8_outputs(2650) <= layer7_outputs(4478);
    layer8_outputs(2651) <= not((layer7_outputs(2939)) xor (layer7_outputs(1533)));
    layer8_outputs(2652) <= not(layer7_outputs(1729));
    layer8_outputs(2653) <= (layer7_outputs(1426)) xor (layer7_outputs(3905));
    layer8_outputs(2654) <= (layer7_outputs(4523)) and not (layer7_outputs(2367));
    layer8_outputs(2655) <= (layer7_outputs(1632)) and not (layer7_outputs(3725));
    layer8_outputs(2656) <= layer7_outputs(2785);
    layer8_outputs(2657) <= layer7_outputs(3982);
    layer8_outputs(2658) <= layer7_outputs(3256);
    layer8_outputs(2659) <= layer7_outputs(4619);
    layer8_outputs(2660) <= (layer7_outputs(1294)) xor (layer7_outputs(4060));
    layer8_outputs(2661) <= (layer7_outputs(633)) and (layer7_outputs(2048));
    layer8_outputs(2662) <= (layer7_outputs(3682)) xor (layer7_outputs(3783));
    layer8_outputs(2663) <= not(layer7_outputs(5001));
    layer8_outputs(2664) <= '1';
    layer8_outputs(2665) <= not((layer7_outputs(3181)) and (layer7_outputs(2525)));
    layer8_outputs(2666) <= layer7_outputs(2965);
    layer8_outputs(2667) <= not(layer7_outputs(2116));
    layer8_outputs(2668) <= (layer7_outputs(666)) and (layer7_outputs(1749));
    layer8_outputs(2669) <= (layer7_outputs(1488)) xor (layer7_outputs(1595));
    layer8_outputs(2670) <= (layer7_outputs(2697)) and not (layer7_outputs(4782));
    layer8_outputs(2671) <= '1';
    layer8_outputs(2672) <= (layer7_outputs(4353)) xor (layer7_outputs(3772));
    layer8_outputs(2673) <= not(layer7_outputs(99));
    layer8_outputs(2674) <= (layer7_outputs(2758)) and not (layer7_outputs(3577));
    layer8_outputs(2675) <= not((layer7_outputs(3116)) or (layer7_outputs(3661)));
    layer8_outputs(2676) <= (layer7_outputs(3046)) xor (layer7_outputs(3528));
    layer8_outputs(2677) <= (layer7_outputs(3631)) and not (layer7_outputs(3351));
    layer8_outputs(2678) <= not((layer7_outputs(4174)) and (layer7_outputs(1781)));
    layer8_outputs(2679) <= not(layer7_outputs(3301));
    layer8_outputs(2680) <= layer7_outputs(3123);
    layer8_outputs(2681) <= not((layer7_outputs(3969)) or (layer7_outputs(1872)));
    layer8_outputs(2682) <= not(layer7_outputs(4675));
    layer8_outputs(2683) <= (layer7_outputs(3085)) xor (layer7_outputs(970));
    layer8_outputs(2684) <= layer7_outputs(816);
    layer8_outputs(2685) <= not((layer7_outputs(601)) and (layer7_outputs(4248)));
    layer8_outputs(2686) <= not((layer7_outputs(393)) xor (layer7_outputs(4530)));
    layer8_outputs(2687) <= not((layer7_outputs(2564)) or (layer7_outputs(1946)));
    layer8_outputs(2688) <= not(layer7_outputs(3653));
    layer8_outputs(2689) <= not((layer7_outputs(2124)) xor (layer7_outputs(3946)));
    layer8_outputs(2690) <= layer7_outputs(1510);
    layer8_outputs(2691) <= layer7_outputs(1720);
    layer8_outputs(2692) <= layer7_outputs(4591);
    layer8_outputs(2693) <= not(layer7_outputs(4448));
    layer8_outputs(2694) <= layer7_outputs(1);
    layer8_outputs(2695) <= layer7_outputs(245);
    layer8_outputs(2696) <= not(layer7_outputs(1447)) or (layer7_outputs(584));
    layer8_outputs(2697) <= (layer7_outputs(2825)) and not (layer7_outputs(5016));
    layer8_outputs(2698) <= not(layer7_outputs(3300));
    layer8_outputs(2699) <= not((layer7_outputs(701)) and (layer7_outputs(4535)));
    layer8_outputs(2700) <= layer7_outputs(1606);
    layer8_outputs(2701) <= not(layer7_outputs(2774));
    layer8_outputs(2702) <= not((layer7_outputs(3324)) and (layer7_outputs(2215)));
    layer8_outputs(2703) <= not((layer7_outputs(1246)) xor (layer7_outputs(3609)));
    layer8_outputs(2704) <= not((layer7_outputs(3545)) xor (layer7_outputs(1978)));
    layer8_outputs(2705) <= layer7_outputs(3342);
    layer8_outputs(2706) <= not(layer7_outputs(1268));
    layer8_outputs(2707) <= '0';
    layer8_outputs(2708) <= not((layer7_outputs(3845)) or (layer7_outputs(4466)));
    layer8_outputs(2709) <= layer7_outputs(3130);
    layer8_outputs(2710) <= not((layer7_outputs(1523)) xor (layer7_outputs(1255)));
    layer8_outputs(2711) <= layer7_outputs(1254);
    layer8_outputs(2712) <= not((layer7_outputs(2422)) or (layer7_outputs(3944)));
    layer8_outputs(2713) <= not((layer7_outputs(2708)) xor (layer7_outputs(3430)));
    layer8_outputs(2714) <= layer7_outputs(4629);
    layer8_outputs(2715) <= layer7_outputs(2653);
    layer8_outputs(2716) <= (layer7_outputs(2431)) xor (layer7_outputs(3844));
    layer8_outputs(2717) <= not(layer7_outputs(2480));
    layer8_outputs(2718) <= not(layer7_outputs(3088));
    layer8_outputs(2719) <= not(layer7_outputs(362));
    layer8_outputs(2720) <= (layer7_outputs(3337)) xor (layer7_outputs(1810));
    layer8_outputs(2721) <= layer7_outputs(956);
    layer8_outputs(2722) <= not(layer7_outputs(2032));
    layer8_outputs(2723) <= not(layer7_outputs(1894));
    layer8_outputs(2724) <= not((layer7_outputs(1724)) xor (layer7_outputs(3036)));
    layer8_outputs(2725) <= not(layer7_outputs(4016));
    layer8_outputs(2726) <= not((layer7_outputs(558)) xor (layer7_outputs(2088)));
    layer8_outputs(2727) <= not((layer7_outputs(1082)) xor (layer7_outputs(1372)));
    layer8_outputs(2728) <= not(layer7_outputs(2335));
    layer8_outputs(2729) <= (layer7_outputs(3383)) xor (layer7_outputs(2456));
    layer8_outputs(2730) <= (layer7_outputs(251)) or (layer7_outputs(1371));
    layer8_outputs(2731) <= not((layer7_outputs(4519)) xor (layer7_outputs(3551)));
    layer8_outputs(2732) <= '1';
    layer8_outputs(2733) <= layer7_outputs(4906);
    layer8_outputs(2734) <= not((layer7_outputs(203)) or (layer7_outputs(996)));
    layer8_outputs(2735) <= not(layer7_outputs(3687));
    layer8_outputs(2736) <= not(layer7_outputs(61));
    layer8_outputs(2737) <= not((layer7_outputs(1349)) xor (layer7_outputs(2900)));
    layer8_outputs(2738) <= not(layer7_outputs(2591));
    layer8_outputs(2739) <= not(layer7_outputs(1734));
    layer8_outputs(2740) <= not((layer7_outputs(387)) xor (layer7_outputs(4847)));
    layer8_outputs(2741) <= (layer7_outputs(4881)) xor (layer7_outputs(2492));
    layer8_outputs(2742) <= (layer7_outputs(1322)) and not (layer7_outputs(2239));
    layer8_outputs(2743) <= '0';
    layer8_outputs(2744) <= layer7_outputs(2050);
    layer8_outputs(2745) <= not(layer7_outputs(2469)) or (layer7_outputs(4757));
    layer8_outputs(2746) <= layer7_outputs(2071);
    layer8_outputs(2747) <= layer7_outputs(1923);
    layer8_outputs(2748) <= not(layer7_outputs(2252)) or (layer7_outputs(3143));
    layer8_outputs(2749) <= not(layer7_outputs(2584));
    layer8_outputs(2750) <= layer7_outputs(854);
    layer8_outputs(2751) <= not(layer7_outputs(2123));
    layer8_outputs(2752) <= (layer7_outputs(3727)) xor (layer7_outputs(497));
    layer8_outputs(2753) <= not(layer7_outputs(1566));
    layer8_outputs(2754) <= (layer7_outputs(4850)) xor (layer7_outputs(4928));
    layer8_outputs(2755) <= not((layer7_outputs(4728)) xor (layer7_outputs(963)));
    layer8_outputs(2756) <= layer7_outputs(4436);
    layer8_outputs(2757) <= not(layer7_outputs(4484));
    layer8_outputs(2758) <= not(layer7_outputs(439));
    layer8_outputs(2759) <= layer7_outputs(2539);
    layer8_outputs(2760) <= layer7_outputs(1803);
    layer8_outputs(2761) <= not(layer7_outputs(3219));
    layer8_outputs(2762) <= (layer7_outputs(3451)) xor (layer7_outputs(5071));
    layer8_outputs(2763) <= not((layer7_outputs(1850)) xor (layer7_outputs(4276)));
    layer8_outputs(2764) <= (layer7_outputs(4670)) and (layer7_outputs(3374));
    layer8_outputs(2765) <= not(layer7_outputs(448)) or (layer7_outputs(4660));
    layer8_outputs(2766) <= (layer7_outputs(92)) or (layer7_outputs(1422));
    layer8_outputs(2767) <= not(layer7_outputs(4982)) or (layer7_outputs(4582));
    layer8_outputs(2768) <= not(layer7_outputs(4570));
    layer8_outputs(2769) <= layer7_outputs(2653);
    layer8_outputs(2770) <= not((layer7_outputs(4788)) xor (layer7_outputs(3178)));
    layer8_outputs(2771) <= not((layer7_outputs(715)) xor (layer7_outputs(3285)));
    layer8_outputs(2772) <= not((layer7_outputs(351)) xor (layer7_outputs(3630)));
    layer8_outputs(2773) <= (layer7_outputs(3767)) xor (layer7_outputs(2141));
    layer8_outputs(2774) <= (layer7_outputs(4718)) xor (layer7_outputs(309));
    layer8_outputs(2775) <= not((layer7_outputs(1178)) xor (layer7_outputs(3697)));
    layer8_outputs(2776) <= layer7_outputs(4403);
    layer8_outputs(2777) <= not(layer7_outputs(961));
    layer8_outputs(2778) <= not(layer7_outputs(2468));
    layer8_outputs(2779) <= layer7_outputs(410);
    layer8_outputs(2780) <= (layer7_outputs(3066)) or (layer7_outputs(2824));
    layer8_outputs(2781) <= layer7_outputs(268);
    layer8_outputs(2782) <= layer7_outputs(2412);
    layer8_outputs(2783) <= not(layer7_outputs(1875));
    layer8_outputs(2784) <= (layer7_outputs(723)) xor (layer7_outputs(1582));
    layer8_outputs(2785) <= not((layer7_outputs(2521)) xor (layer7_outputs(4617)));
    layer8_outputs(2786) <= layer7_outputs(3056);
    layer8_outputs(2787) <= layer7_outputs(1070);
    layer8_outputs(2788) <= not(layer7_outputs(2687)) or (layer7_outputs(2090));
    layer8_outputs(2789) <= (layer7_outputs(868)) and not (layer7_outputs(699));
    layer8_outputs(2790) <= not((layer7_outputs(4011)) xor (layer7_outputs(2544)));
    layer8_outputs(2791) <= layer7_outputs(2368);
    layer8_outputs(2792) <= (layer7_outputs(5010)) xor (layer7_outputs(340));
    layer8_outputs(2793) <= not((layer7_outputs(3228)) xor (layer7_outputs(4295)));
    layer8_outputs(2794) <= layer7_outputs(1578);
    layer8_outputs(2795) <= not(layer7_outputs(571));
    layer8_outputs(2796) <= layer7_outputs(4512);
    layer8_outputs(2797) <= not((layer7_outputs(1437)) xor (layer7_outputs(3891)));
    layer8_outputs(2798) <= layer7_outputs(1779);
    layer8_outputs(2799) <= layer7_outputs(2821);
    layer8_outputs(2800) <= not(layer7_outputs(4291));
    layer8_outputs(2801) <= not((layer7_outputs(5017)) xor (layer7_outputs(4339)));
    layer8_outputs(2802) <= not((layer7_outputs(2796)) xor (layer7_outputs(2483)));
    layer8_outputs(2803) <= (layer7_outputs(2360)) and not (layer7_outputs(74));
    layer8_outputs(2804) <= not((layer7_outputs(2897)) xor (layer7_outputs(2667)));
    layer8_outputs(2805) <= layer7_outputs(3167);
    layer8_outputs(2806) <= not((layer7_outputs(4368)) xor (layer7_outputs(4970)));
    layer8_outputs(2807) <= not(layer7_outputs(2028));
    layer8_outputs(2808) <= (layer7_outputs(1445)) xor (layer7_outputs(4522));
    layer8_outputs(2809) <= (layer7_outputs(2826)) and not (layer7_outputs(2478));
    layer8_outputs(2810) <= layer7_outputs(430);
    layer8_outputs(2811) <= not(layer7_outputs(4803)) or (layer7_outputs(904));
    layer8_outputs(2812) <= (layer7_outputs(1293)) and (layer7_outputs(3256));
    layer8_outputs(2813) <= not(layer7_outputs(3354));
    layer8_outputs(2814) <= layer7_outputs(1453);
    layer8_outputs(2815) <= not(layer7_outputs(3515));
    layer8_outputs(2816) <= layer7_outputs(1515);
    layer8_outputs(2817) <= not((layer7_outputs(4403)) xor (layer7_outputs(1054)));
    layer8_outputs(2818) <= layer7_outputs(301);
    layer8_outputs(2819) <= not((layer7_outputs(654)) xor (layer7_outputs(3481)));
    layer8_outputs(2820) <= (layer7_outputs(4890)) and not (layer7_outputs(3911));
    layer8_outputs(2821) <= not(layer7_outputs(3801)) or (layer7_outputs(1559));
    layer8_outputs(2822) <= not(layer7_outputs(3487));
    layer8_outputs(2823) <= layer7_outputs(70);
    layer8_outputs(2824) <= layer7_outputs(483);
    layer8_outputs(2825) <= layer7_outputs(2709);
    layer8_outputs(2826) <= (layer7_outputs(1615)) xor (layer7_outputs(1888));
    layer8_outputs(2827) <= layer7_outputs(4348);
    layer8_outputs(2828) <= not(layer7_outputs(3915));
    layer8_outputs(2829) <= not(layer7_outputs(3489));
    layer8_outputs(2830) <= not(layer7_outputs(4954)) or (layer7_outputs(4748));
    layer8_outputs(2831) <= not((layer7_outputs(4230)) and (layer7_outputs(1434)));
    layer8_outputs(2832) <= layer7_outputs(4528);
    layer8_outputs(2833) <= layer7_outputs(1893);
    layer8_outputs(2834) <= (layer7_outputs(4678)) xor (layer7_outputs(4061));
    layer8_outputs(2835) <= layer7_outputs(4692);
    layer8_outputs(2836) <= not((layer7_outputs(787)) and (layer7_outputs(4866)));
    layer8_outputs(2837) <= not(layer7_outputs(2906));
    layer8_outputs(2838) <= layer7_outputs(802);
    layer8_outputs(2839) <= not((layer7_outputs(3321)) xor (layer7_outputs(319)));
    layer8_outputs(2840) <= not(layer7_outputs(4622));
    layer8_outputs(2841) <= (layer7_outputs(2879)) xor (layer7_outputs(2922));
    layer8_outputs(2842) <= (layer7_outputs(1970)) xor (layer7_outputs(2472));
    layer8_outputs(2843) <= not(layer7_outputs(1671)) or (layer7_outputs(2465));
    layer8_outputs(2844) <= (layer7_outputs(2927)) xor (layer7_outputs(1075));
    layer8_outputs(2845) <= not((layer7_outputs(4737)) xor (layer7_outputs(4426)));
    layer8_outputs(2846) <= layer7_outputs(169);
    layer8_outputs(2847) <= not((layer7_outputs(1458)) or (layer7_outputs(3526)));
    layer8_outputs(2848) <= not((layer7_outputs(728)) and (layer7_outputs(5082)));
    layer8_outputs(2849) <= not(layer7_outputs(815));
    layer8_outputs(2850) <= (layer7_outputs(3611)) xor (layer7_outputs(3615));
    layer8_outputs(2851) <= (layer7_outputs(1274)) xor (layer7_outputs(1840));
    layer8_outputs(2852) <= '1';
    layer8_outputs(2853) <= not(layer7_outputs(1181));
    layer8_outputs(2854) <= not((layer7_outputs(1952)) or (layer7_outputs(3225)));
    layer8_outputs(2855) <= layer7_outputs(2096);
    layer8_outputs(2856) <= (layer7_outputs(1908)) and not (layer7_outputs(3880));
    layer8_outputs(2857) <= layer7_outputs(4926);
    layer8_outputs(2858) <= not((layer7_outputs(1336)) xor (layer7_outputs(2979)));
    layer8_outputs(2859) <= layer7_outputs(4411);
    layer8_outputs(2860) <= (layer7_outputs(4380)) and not (layer7_outputs(3353));
    layer8_outputs(2861) <= (layer7_outputs(4593)) xor (layer7_outputs(188));
    layer8_outputs(2862) <= not(layer7_outputs(314));
    layer8_outputs(2863) <= (layer7_outputs(1824)) and not (layer7_outputs(886));
    layer8_outputs(2864) <= (layer7_outputs(1981)) xor (layer7_outputs(4516));
    layer8_outputs(2865) <= (layer7_outputs(3286)) xor (layer7_outputs(3674));
    layer8_outputs(2866) <= layer7_outputs(3824);
    layer8_outputs(2867) <= not(layer7_outputs(2893));
    layer8_outputs(2868) <= (layer7_outputs(48)) xor (layer7_outputs(951));
    layer8_outputs(2869) <= layer7_outputs(1206);
    layer8_outputs(2870) <= not((layer7_outputs(3741)) xor (layer7_outputs(5071)));
    layer8_outputs(2871) <= not((layer7_outputs(4752)) xor (layer7_outputs(4434)));
    layer8_outputs(2872) <= layer7_outputs(2493);
    layer8_outputs(2873) <= not(layer7_outputs(1981));
    layer8_outputs(2874) <= layer7_outputs(180);
    layer8_outputs(2875) <= not((layer7_outputs(2015)) xor (layer7_outputs(4350)));
    layer8_outputs(2876) <= not(layer7_outputs(1449));
    layer8_outputs(2877) <= not(layer7_outputs(4082));
    layer8_outputs(2878) <= not((layer7_outputs(2078)) xor (layer7_outputs(686)));
    layer8_outputs(2879) <= not(layer7_outputs(2910));
    layer8_outputs(2880) <= not(layer7_outputs(61));
    layer8_outputs(2881) <= not(layer7_outputs(1546)) or (layer7_outputs(233));
    layer8_outputs(2882) <= (layer7_outputs(5047)) or (layer7_outputs(2768));
    layer8_outputs(2883) <= (layer7_outputs(5002)) xor (layer7_outputs(4888));
    layer8_outputs(2884) <= not(layer7_outputs(3383));
    layer8_outputs(2885) <= (layer7_outputs(2836)) xor (layer7_outputs(2596));
    layer8_outputs(2886) <= not(layer7_outputs(4556));
    layer8_outputs(2887) <= not(layer7_outputs(4942));
    layer8_outputs(2888) <= layer7_outputs(4345);
    layer8_outputs(2889) <= layer7_outputs(3426);
    layer8_outputs(2890) <= (layer7_outputs(1624)) and (layer7_outputs(1348));
    layer8_outputs(2891) <= layer7_outputs(1602);
    layer8_outputs(2892) <= (layer7_outputs(4387)) xor (layer7_outputs(2615));
    layer8_outputs(2893) <= not(layer7_outputs(4184));
    layer8_outputs(2894) <= (layer7_outputs(3723)) xor (layer7_outputs(4668));
    layer8_outputs(2895) <= (layer7_outputs(995)) xor (layer7_outputs(1579));
    layer8_outputs(2896) <= not((layer7_outputs(4366)) xor (layer7_outputs(1470)));
    layer8_outputs(2897) <= layer7_outputs(2747);
    layer8_outputs(2898) <= layer7_outputs(1308);
    layer8_outputs(2899) <= not(layer7_outputs(2939));
    layer8_outputs(2900) <= not(layer7_outputs(2673)) or (layer7_outputs(1266));
    layer8_outputs(2901) <= layer7_outputs(2854);
    layer8_outputs(2902) <= not((layer7_outputs(4178)) xor (layer7_outputs(2752)));
    layer8_outputs(2903) <= '0';
    layer8_outputs(2904) <= not((layer7_outputs(3451)) or (layer7_outputs(576)));
    layer8_outputs(2905) <= (layer7_outputs(4798)) xor (layer7_outputs(4413));
    layer8_outputs(2906) <= not(layer7_outputs(4695)) or (layer7_outputs(258));
    layer8_outputs(2907) <= not(layer7_outputs(1046)) or (layer7_outputs(643));
    layer8_outputs(2908) <= (layer7_outputs(4423)) and (layer7_outputs(2192));
    layer8_outputs(2909) <= not(layer7_outputs(2288)) or (layer7_outputs(3555));
    layer8_outputs(2910) <= (layer7_outputs(1986)) and (layer7_outputs(1567));
    layer8_outputs(2911) <= not(layer7_outputs(4302));
    layer8_outputs(2912) <= not((layer7_outputs(437)) xor (layer7_outputs(3052)));
    layer8_outputs(2913) <= not((layer7_outputs(3102)) xor (layer7_outputs(2352)));
    layer8_outputs(2914) <= not(layer7_outputs(1253));
    layer8_outputs(2915) <= (layer7_outputs(594)) or (layer7_outputs(4973));
    layer8_outputs(2916) <= layer7_outputs(2632);
    layer8_outputs(2917) <= layer7_outputs(2975);
    layer8_outputs(2918) <= layer7_outputs(1571);
    layer8_outputs(2919) <= layer7_outputs(3680);
    layer8_outputs(2920) <= not(layer7_outputs(1463));
    layer8_outputs(2921) <= (layer7_outputs(2832)) and not (layer7_outputs(1744));
    layer8_outputs(2922) <= not((layer7_outputs(3141)) or (layer7_outputs(3416)));
    layer8_outputs(2923) <= not((layer7_outputs(3743)) xor (layer7_outputs(2937)));
    layer8_outputs(2924) <= layer7_outputs(3274);
    layer8_outputs(2925) <= not(layer7_outputs(4614)) or (layer7_outputs(4824));
    layer8_outputs(2926) <= (layer7_outputs(1243)) xor (layer7_outputs(2048));
    layer8_outputs(2927) <= (layer7_outputs(4729)) xor (layer7_outputs(2155));
    layer8_outputs(2928) <= not(layer7_outputs(2578));
    layer8_outputs(2929) <= layer7_outputs(4988);
    layer8_outputs(2930) <= '1';
    layer8_outputs(2931) <= not((layer7_outputs(1865)) xor (layer7_outputs(1805)));
    layer8_outputs(2932) <= (layer7_outputs(222)) xor (layer7_outputs(2849));
    layer8_outputs(2933) <= (layer7_outputs(1706)) xor (layer7_outputs(2348));
    layer8_outputs(2934) <= (layer7_outputs(1300)) and not (layer7_outputs(830));
    layer8_outputs(2935) <= (layer7_outputs(4813)) and not (layer7_outputs(2807));
    layer8_outputs(2936) <= (layer7_outputs(2961)) and not (layer7_outputs(803));
    layer8_outputs(2937) <= (layer7_outputs(2475)) and not (layer7_outputs(3215));
    layer8_outputs(2938) <= not(layer7_outputs(140));
    layer8_outputs(2939) <= (layer7_outputs(1568)) and not (layer7_outputs(2278));
    layer8_outputs(2940) <= not((layer7_outputs(1749)) or (layer7_outputs(480)));
    layer8_outputs(2941) <= (layer7_outputs(2283)) or (layer7_outputs(2087));
    layer8_outputs(2942) <= layer7_outputs(2370);
    layer8_outputs(2943) <= not(layer7_outputs(987)) or (layer7_outputs(4834));
    layer8_outputs(2944) <= not(layer7_outputs(646));
    layer8_outputs(2945) <= layer7_outputs(3345);
    layer8_outputs(2946) <= (layer7_outputs(893)) xor (layer7_outputs(4215));
    layer8_outputs(2947) <= (layer7_outputs(3711)) xor (layer7_outputs(2086));
    layer8_outputs(2948) <= not(layer7_outputs(2879));
    layer8_outputs(2949) <= (layer7_outputs(115)) or (layer7_outputs(4913));
    layer8_outputs(2950) <= not(layer7_outputs(3904));
    layer8_outputs(2951) <= (layer7_outputs(1370)) xor (layer7_outputs(599));
    layer8_outputs(2952) <= (layer7_outputs(1598)) xor (layer7_outputs(3831));
    layer8_outputs(2953) <= layer7_outputs(4442);
    layer8_outputs(2954) <= layer7_outputs(769);
    layer8_outputs(2955) <= layer7_outputs(1597);
    layer8_outputs(2956) <= (layer7_outputs(224)) and (layer7_outputs(2627));
    layer8_outputs(2957) <= not((layer7_outputs(3644)) or (layer7_outputs(3929)));
    layer8_outputs(2958) <= (layer7_outputs(834)) xor (layer7_outputs(690));
    layer8_outputs(2959) <= not((layer7_outputs(2655)) xor (layer7_outputs(1079)));
    layer8_outputs(2960) <= (layer7_outputs(4144)) and (layer7_outputs(1761));
    layer8_outputs(2961) <= (layer7_outputs(2424)) xor (layer7_outputs(3396));
    layer8_outputs(2962) <= layer7_outputs(4574);
    layer8_outputs(2963) <= layer7_outputs(4618);
    layer8_outputs(2964) <= not(layer7_outputs(2508));
    layer8_outputs(2965) <= not(layer7_outputs(1044));
    layer8_outputs(2966) <= layer7_outputs(4110);
    layer8_outputs(2967) <= not(layer7_outputs(4707));
    layer8_outputs(2968) <= not(layer7_outputs(4688));
    layer8_outputs(2969) <= layer7_outputs(1028);
    layer8_outputs(2970) <= not(layer7_outputs(2890));
    layer8_outputs(2971) <= not((layer7_outputs(951)) and (layer7_outputs(378)));
    layer8_outputs(2972) <= not((layer7_outputs(4007)) and (layer7_outputs(3350)));
    layer8_outputs(2973) <= not((layer7_outputs(4749)) xor (layer7_outputs(229)));
    layer8_outputs(2974) <= not(layer7_outputs(4747)) or (layer7_outputs(3081));
    layer8_outputs(2975) <= not((layer7_outputs(2829)) or (layer7_outputs(2353)));
    layer8_outputs(2976) <= not((layer7_outputs(4380)) and (layer7_outputs(2828)));
    layer8_outputs(2977) <= (layer7_outputs(841)) and not (layer7_outputs(3821));
    layer8_outputs(2978) <= '0';
    layer8_outputs(2979) <= not(layer7_outputs(3604)) or (layer7_outputs(2291));
    layer8_outputs(2980) <= not((layer7_outputs(4763)) xor (layer7_outputs(4517)));
    layer8_outputs(2981) <= not((layer7_outputs(3307)) xor (layer7_outputs(2016)));
    layer8_outputs(2982) <= (layer7_outputs(2015)) xor (layer7_outputs(194));
    layer8_outputs(2983) <= not(layer7_outputs(2240));
    layer8_outputs(2984) <= (layer7_outputs(3219)) xor (layer7_outputs(4255));
    layer8_outputs(2985) <= layer7_outputs(1115);
    layer8_outputs(2986) <= not(layer7_outputs(4976)) or (layer7_outputs(3392));
    layer8_outputs(2987) <= layer7_outputs(3997);
    layer8_outputs(2988) <= (layer7_outputs(2047)) xor (layer7_outputs(4708));
    layer8_outputs(2989) <= not(layer7_outputs(2838));
    layer8_outputs(2990) <= (layer7_outputs(4233)) xor (layer7_outputs(2494));
    layer8_outputs(2991) <= (layer7_outputs(51)) xor (layer7_outputs(3685));
    layer8_outputs(2992) <= (layer7_outputs(2149)) xor (layer7_outputs(627));
    layer8_outputs(2993) <= not((layer7_outputs(4955)) and (layer7_outputs(2548)));
    layer8_outputs(2994) <= (layer7_outputs(2079)) and not (layer7_outputs(1044));
    layer8_outputs(2995) <= layer7_outputs(2076);
    layer8_outputs(2996) <= not((layer7_outputs(358)) or (layer7_outputs(3488)));
    layer8_outputs(2997) <= not(layer7_outputs(4818)) or (layer7_outputs(1283));
    layer8_outputs(2998) <= not(layer7_outputs(164));
    layer8_outputs(2999) <= layer7_outputs(4320);
    layer8_outputs(3000) <= not(layer7_outputs(781)) or (layer7_outputs(4331));
    layer8_outputs(3001) <= layer7_outputs(3402);
    layer8_outputs(3002) <= (layer7_outputs(2986)) xor (layer7_outputs(484));
    layer8_outputs(3003) <= not(layer7_outputs(1055));
    layer8_outputs(3004) <= layer7_outputs(2156);
    layer8_outputs(3005) <= (layer7_outputs(1761)) xor (layer7_outputs(2714));
    layer8_outputs(3006) <= (layer7_outputs(1183)) and (layer7_outputs(3863));
    layer8_outputs(3007) <= not(layer7_outputs(811));
    layer8_outputs(3008) <= not((layer7_outputs(3672)) xor (layer7_outputs(328)));
    layer8_outputs(3009) <= (layer7_outputs(2322)) xor (layer7_outputs(286));
    layer8_outputs(3010) <= layer7_outputs(4516);
    layer8_outputs(3011) <= (layer7_outputs(3967)) xor (layer7_outputs(5115));
    layer8_outputs(3012) <= layer7_outputs(3130);
    layer8_outputs(3013) <= layer7_outputs(3520);
    layer8_outputs(3014) <= not((layer7_outputs(3960)) xor (layer7_outputs(4507)));
    layer8_outputs(3015) <= (layer7_outputs(4887)) or (layer7_outputs(1739));
    layer8_outputs(3016) <= not((layer7_outputs(1149)) and (layer7_outputs(395)));
    layer8_outputs(3017) <= not(layer7_outputs(398));
    layer8_outputs(3018) <= not(layer7_outputs(1694));
    layer8_outputs(3019) <= not(layer7_outputs(3247));
    layer8_outputs(3020) <= layer7_outputs(1918);
    layer8_outputs(3021) <= (layer7_outputs(789)) xor (layer7_outputs(1297));
    layer8_outputs(3022) <= layer7_outputs(3397);
    layer8_outputs(3023) <= layer7_outputs(228);
    layer8_outputs(3024) <= not(layer7_outputs(1440)) or (layer7_outputs(3445));
    layer8_outputs(3025) <= layer7_outputs(2260);
    layer8_outputs(3026) <= (layer7_outputs(4467)) or (layer7_outputs(2202));
    layer8_outputs(3027) <= (layer7_outputs(3351)) xor (layer7_outputs(4188));
    layer8_outputs(3028) <= layer7_outputs(4045);
    layer8_outputs(3029) <= not(layer7_outputs(3589)) or (layer7_outputs(3393));
    layer8_outputs(3030) <= layer7_outputs(1756);
    layer8_outputs(3031) <= not(layer7_outputs(9)) or (layer7_outputs(4503));
    layer8_outputs(3032) <= not(layer7_outputs(4483)) or (layer7_outputs(3785));
    layer8_outputs(3033) <= '0';
    layer8_outputs(3034) <= not((layer7_outputs(331)) xor (layer7_outputs(2478)));
    layer8_outputs(3035) <= not((layer7_outputs(2978)) xor (layer7_outputs(3033)));
    layer8_outputs(3036) <= layer7_outputs(29);
    layer8_outputs(3037) <= not(layer7_outputs(1838));
    layer8_outputs(3038) <= layer7_outputs(2211);
    layer8_outputs(3039) <= layer7_outputs(2825);
    layer8_outputs(3040) <= not(layer7_outputs(3048));
    layer8_outputs(3041) <= not(layer7_outputs(2218));
    layer8_outputs(3042) <= not(layer7_outputs(2490));
    layer8_outputs(3043) <= not((layer7_outputs(1098)) xor (layer7_outputs(706)));
    layer8_outputs(3044) <= not((layer7_outputs(2132)) or (layer7_outputs(4355)));
    layer8_outputs(3045) <= not(layer7_outputs(2262));
    layer8_outputs(3046) <= (layer7_outputs(2574)) and not (layer7_outputs(1230));
    layer8_outputs(3047) <= not(layer7_outputs(2353)) or (layer7_outputs(706));
    layer8_outputs(3048) <= not((layer7_outputs(4731)) xor (layer7_outputs(3543)));
    layer8_outputs(3049) <= not(layer7_outputs(4012));
    layer8_outputs(3050) <= not(layer7_outputs(4435));
    layer8_outputs(3051) <= layer7_outputs(4206);
    layer8_outputs(3052) <= layer7_outputs(4938);
    layer8_outputs(3053) <= layer7_outputs(2171);
    layer8_outputs(3054) <= layer7_outputs(3781);
    layer8_outputs(3055) <= (layer7_outputs(2790)) and (layer7_outputs(2762));
    layer8_outputs(3056) <= not(layer7_outputs(3568));
    layer8_outputs(3057) <= (layer7_outputs(1914)) xor (layer7_outputs(4547));
    layer8_outputs(3058) <= (layer7_outputs(2171)) and (layer7_outputs(3681));
    layer8_outputs(3059) <= not(layer7_outputs(2000));
    layer8_outputs(3060) <= not((layer7_outputs(283)) and (layer7_outputs(1892)));
    layer8_outputs(3061) <= not(layer7_outputs(1455));
    layer8_outputs(3062) <= (layer7_outputs(3921)) and (layer7_outputs(3280));
    layer8_outputs(3063) <= layer7_outputs(270);
    layer8_outputs(3064) <= layer7_outputs(3606);
    layer8_outputs(3065) <= not((layer7_outputs(824)) or (layer7_outputs(2074)));
    layer8_outputs(3066) <= not(layer7_outputs(2636)) or (layer7_outputs(2895));
    layer8_outputs(3067) <= layer7_outputs(2696);
    layer8_outputs(3068) <= not(layer7_outputs(1350)) or (layer7_outputs(1097));
    layer8_outputs(3069) <= not(layer7_outputs(2727)) or (layer7_outputs(5091));
    layer8_outputs(3070) <= not(layer7_outputs(1249));
    layer8_outputs(3071) <= not((layer7_outputs(895)) xor (layer7_outputs(3072)));
    layer8_outputs(3072) <= not(layer7_outputs(4562));
    layer8_outputs(3073) <= not(layer7_outputs(3673)) or (layer7_outputs(1093));
    layer8_outputs(3074) <= not(layer7_outputs(1225));
    layer8_outputs(3075) <= not((layer7_outputs(454)) xor (layer7_outputs(278)));
    layer8_outputs(3076) <= not((layer7_outputs(2407)) xor (layer7_outputs(3703)));
    layer8_outputs(3077) <= not(layer7_outputs(826));
    layer8_outputs(3078) <= (layer7_outputs(4394)) or (layer7_outputs(2106));
    layer8_outputs(3079) <= (layer7_outputs(4871)) or (layer7_outputs(4655));
    layer8_outputs(3080) <= (layer7_outputs(4251)) or (layer7_outputs(3707));
    layer8_outputs(3081) <= not(layer7_outputs(4874));
    layer8_outputs(3082) <= (layer7_outputs(655)) or (layer7_outputs(817));
    layer8_outputs(3083) <= not(layer7_outputs(3697));
    layer8_outputs(3084) <= layer7_outputs(3410);
    layer8_outputs(3085) <= layer7_outputs(1721);
    layer8_outputs(3086) <= not(layer7_outputs(1051));
    layer8_outputs(3087) <= not(layer7_outputs(2052));
    layer8_outputs(3088) <= layer7_outputs(765);
    layer8_outputs(3089) <= layer7_outputs(2642);
    layer8_outputs(3090) <= not((layer7_outputs(2767)) xor (layer7_outputs(104)));
    layer8_outputs(3091) <= layer7_outputs(2932);
    layer8_outputs(3092) <= (layer7_outputs(1131)) or (layer7_outputs(3306));
    layer8_outputs(3093) <= not(layer7_outputs(2956));
    layer8_outputs(3094) <= (layer7_outputs(457)) xor (layer7_outputs(2948));
    layer8_outputs(3095) <= not(layer7_outputs(4518)) or (layer7_outputs(113));
    layer8_outputs(3096) <= (layer7_outputs(3908)) and not (layer7_outputs(1408));
    layer8_outputs(3097) <= not(layer7_outputs(101));
    layer8_outputs(3098) <= not((layer7_outputs(3758)) xor (layer7_outputs(2496)));
    layer8_outputs(3099) <= not(layer7_outputs(4261));
    layer8_outputs(3100) <= not(layer7_outputs(4806));
    layer8_outputs(3101) <= not((layer7_outputs(3190)) xor (layer7_outputs(689)));
    layer8_outputs(3102) <= layer7_outputs(250);
    layer8_outputs(3103) <= not(layer7_outputs(2302));
    layer8_outputs(3104) <= (layer7_outputs(4166)) xor (layer7_outputs(1156));
    layer8_outputs(3105) <= not(layer7_outputs(4655)) or (layer7_outputs(3214));
    layer8_outputs(3106) <= not(layer7_outputs(1764));
    layer8_outputs(3107) <= layer7_outputs(2909);
    layer8_outputs(3108) <= layer7_outputs(2354);
    layer8_outputs(3109) <= not((layer7_outputs(1541)) xor (layer7_outputs(2873)));
    layer8_outputs(3110) <= not(layer7_outputs(4216));
    layer8_outputs(3111) <= layer7_outputs(3661);
    layer8_outputs(3112) <= layer7_outputs(3864);
    layer8_outputs(3113) <= not(layer7_outputs(4427));
    layer8_outputs(3114) <= layer7_outputs(4924);
    layer8_outputs(3115) <= (layer7_outputs(773)) or (layer7_outputs(4635));
    layer8_outputs(3116) <= (layer7_outputs(4620)) xor (layer7_outputs(4489));
    layer8_outputs(3117) <= not(layer7_outputs(983));
    layer8_outputs(3118) <= not(layer7_outputs(3073));
    layer8_outputs(3119) <= not(layer7_outputs(1953)) or (layer7_outputs(729));
    layer8_outputs(3120) <= not((layer7_outputs(4768)) or (layer7_outputs(2166)));
    layer8_outputs(3121) <= not(layer7_outputs(2513));
    layer8_outputs(3122) <= (layer7_outputs(4972)) and not (layer7_outputs(2157));
    layer8_outputs(3123) <= (layer7_outputs(1484)) and not (layer7_outputs(1785));
    layer8_outputs(3124) <= not(layer7_outputs(432));
    layer8_outputs(3125) <= not(layer7_outputs(2940));
    layer8_outputs(3126) <= not(layer7_outputs(1870));
    layer8_outputs(3127) <= layer7_outputs(4202);
    layer8_outputs(3128) <= layer7_outputs(336);
    layer8_outputs(3129) <= not((layer7_outputs(3432)) xor (layer7_outputs(2264)));
    layer8_outputs(3130) <= not(layer7_outputs(2952)) or (layer7_outputs(514));
    layer8_outputs(3131) <= (layer7_outputs(3549)) xor (layer7_outputs(478));
    layer8_outputs(3132) <= layer7_outputs(4554);
    layer8_outputs(3133) <= (layer7_outputs(3862)) xor (layer7_outputs(1768));
    layer8_outputs(3134) <= not((layer7_outputs(797)) xor (layer7_outputs(2184)));
    layer8_outputs(3135) <= not(layer7_outputs(3581));
    layer8_outputs(3136) <= layer7_outputs(4547);
    layer8_outputs(3137) <= not(layer7_outputs(2283));
    layer8_outputs(3138) <= (layer7_outputs(3628)) and not (layer7_outputs(1407));
    layer8_outputs(3139) <= layer7_outputs(1898);
    layer8_outputs(3140) <= layer7_outputs(3266);
    layer8_outputs(3141) <= layer7_outputs(4311);
    layer8_outputs(3142) <= not((layer7_outputs(4081)) and (layer7_outputs(1954)));
    layer8_outputs(3143) <= layer7_outputs(2276);
    layer8_outputs(3144) <= not(layer7_outputs(3575));
    layer8_outputs(3145) <= layer7_outputs(4575);
    layer8_outputs(3146) <= layer7_outputs(3097);
    layer8_outputs(3147) <= not(layer7_outputs(4022));
    layer8_outputs(3148) <= (layer7_outputs(3508)) and not (layer7_outputs(1553));
    layer8_outputs(3149) <= layer7_outputs(2069);
    layer8_outputs(3150) <= not(layer7_outputs(1043));
    layer8_outputs(3151) <= layer7_outputs(2434);
    layer8_outputs(3152) <= (layer7_outputs(830)) xor (layer7_outputs(4861));
    layer8_outputs(3153) <= (layer7_outputs(4977)) and not (layer7_outputs(1064));
    layer8_outputs(3154) <= layer7_outputs(2954);
    layer8_outputs(3155) <= not(layer7_outputs(4957));
    layer8_outputs(3156) <= (layer7_outputs(1412)) xor (layer7_outputs(312));
    layer8_outputs(3157) <= (layer7_outputs(3926)) or (layer7_outputs(3016));
    layer8_outputs(3158) <= layer7_outputs(2980);
    layer8_outputs(3159) <= (layer7_outputs(1364)) xor (layer7_outputs(877));
    layer8_outputs(3160) <= layer7_outputs(1833);
    layer8_outputs(3161) <= not((layer7_outputs(4507)) or (layer7_outputs(198)));
    layer8_outputs(3162) <= not((layer7_outputs(4630)) xor (layer7_outputs(1524)));
    layer8_outputs(3163) <= not(layer7_outputs(3736));
    layer8_outputs(3164) <= not((layer7_outputs(4944)) or (layer7_outputs(2898)));
    layer8_outputs(3165) <= (layer7_outputs(3782)) xor (layer7_outputs(2972));
    layer8_outputs(3166) <= not(layer7_outputs(2078));
    layer8_outputs(3167) <= layer7_outputs(1130);
    layer8_outputs(3168) <= not((layer7_outputs(4610)) xor (layer7_outputs(465)));
    layer8_outputs(3169) <= not(layer7_outputs(3502));
    layer8_outputs(3170) <= (layer7_outputs(2318)) xor (layer7_outputs(4717));
    layer8_outputs(3171) <= (layer7_outputs(1764)) and not (layer7_outputs(2684));
    layer8_outputs(3172) <= layer7_outputs(868);
    layer8_outputs(3173) <= (layer7_outputs(2905)) or (layer7_outputs(3245));
    layer8_outputs(3174) <= layer7_outputs(888);
    layer8_outputs(3175) <= not(layer7_outputs(3003)) or (layer7_outputs(3514));
    layer8_outputs(3176) <= (layer7_outputs(1603)) and not (layer7_outputs(1405));
    layer8_outputs(3177) <= not(layer7_outputs(4116)) or (layer7_outputs(1569));
    layer8_outputs(3178) <= layer7_outputs(3980);
    layer8_outputs(3179) <= not((layer7_outputs(3026)) xor (layer7_outputs(5074)));
    layer8_outputs(3180) <= layer7_outputs(4222);
    layer8_outputs(3181) <= not(layer7_outputs(2887));
    layer8_outputs(3182) <= layer7_outputs(1067);
    layer8_outputs(3183) <= layer7_outputs(4744);
    layer8_outputs(3184) <= not(layer7_outputs(4481));
    layer8_outputs(3185) <= not(layer7_outputs(296));
    layer8_outputs(3186) <= layer7_outputs(1179);
    layer8_outputs(3187) <= layer7_outputs(568);
    layer8_outputs(3188) <= layer7_outputs(1522);
    layer8_outputs(3189) <= not(layer7_outputs(2525)) or (layer7_outputs(2634));
    layer8_outputs(3190) <= not((layer7_outputs(4099)) and (layer7_outputs(4817)));
    layer8_outputs(3191) <= not(layer7_outputs(1430));
    layer8_outputs(3192) <= layer7_outputs(2430);
    layer8_outputs(3193) <= not(layer7_outputs(982));
    layer8_outputs(3194) <= not((layer7_outputs(2101)) xor (layer7_outputs(189)));
    layer8_outputs(3195) <= (layer7_outputs(667)) and not (layer7_outputs(1547));
    layer8_outputs(3196) <= (layer7_outputs(3061)) or (layer7_outputs(1415));
    layer8_outputs(3197) <= layer7_outputs(686);
    layer8_outputs(3198) <= layer7_outputs(1855);
    layer8_outputs(3199) <= layer7_outputs(3247);
    layer8_outputs(3200) <= not(layer7_outputs(1809));
    layer8_outputs(3201) <= (layer7_outputs(2983)) or (layer7_outputs(1845));
    layer8_outputs(3202) <= not(layer7_outputs(3931));
    layer8_outputs(3203) <= layer7_outputs(4102);
    layer8_outputs(3204) <= not(layer7_outputs(2756));
    layer8_outputs(3205) <= not(layer7_outputs(2422));
    layer8_outputs(3206) <= not((layer7_outputs(3424)) xor (layer7_outputs(3079)));
    layer8_outputs(3207) <= '1';
    layer8_outputs(3208) <= (layer7_outputs(4335)) xor (layer7_outputs(1580));
    layer8_outputs(3209) <= not(layer7_outputs(460));
    layer8_outputs(3210) <= not(layer7_outputs(441)) or (layer7_outputs(4623));
    layer8_outputs(3211) <= layer7_outputs(313);
    layer8_outputs(3212) <= not(layer7_outputs(2306));
    layer8_outputs(3213) <= (layer7_outputs(5070)) xor (layer7_outputs(1143));
    layer8_outputs(3214) <= not(layer7_outputs(1586));
    layer8_outputs(3215) <= (layer7_outputs(4070)) xor (layer7_outputs(1496));
    layer8_outputs(3216) <= (layer7_outputs(2004)) xor (layer7_outputs(4982));
    layer8_outputs(3217) <= (layer7_outputs(1038)) xor (layer7_outputs(177));
    layer8_outputs(3218) <= not(layer7_outputs(4252));
    layer8_outputs(3219) <= (layer7_outputs(2753)) and not (layer7_outputs(4301));
    layer8_outputs(3220) <= (layer7_outputs(3323)) or (layer7_outputs(3032));
    layer8_outputs(3221) <= not((layer7_outputs(4948)) xor (layer7_outputs(4374)));
    layer8_outputs(3222) <= not((layer7_outputs(1192)) xor (layer7_outputs(2856)));
    layer8_outputs(3223) <= (layer7_outputs(4307)) xor (layer7_outputs(2924));
    layer8_outputs(3224) <= not((layer7_outputs(4461)) or (layer7_outputs(3213)));
    layer8_outputs(3225) <= layer7_outputs(4037);
    layer8_outputs(3226) <= layer7_outputs(3417);
    layer8_outputs(3227) <= layer7_outputs(2117);
    layer8_outputs(3228) <= layer7_outputs(2974);
    layer8_outputs(3229) <= not(layer7_outputs(2683));
    layer8_outputs(3230) <= layer7_outputs(2076);
    layer8_outputs(3231) <= not((layer7_outputs(2536)) xor (layer7_outputs(3593)));
    layer8_outputs(3232) <= not(layer7_outputs(3775));
    layer8_outputs(3233) <= not(layer7_outputs(473));
    layer8_outputs(3234) <= layer7_outputs(2332);
    layer8_outputs(3235) <= not(layer7_outputs(5004)) or (layer7_outputs(942));
    layer8_outputs(3236) <= (layer7_outputs(1678)) xor (layer7_outputs(2870));
    layer8_outputs(3237) <= (layer7_outputs(4827)) and (layer7_outputs(844));
    layer8_outputs(3238) <= not((layer7_outputs(1000)) or (layer7_outputs(255)));
    layer8_outputs(3239) <= not(layer7_outputs(744));
    layer8_outputs(3240) <= not(layer7_outputs(896));
    layer8_outputs(3241) <= not(layer7_outputs(3580));
    layer8_outputs(3242) <= not(layer7_outputs(3139));
    layer8_outputs(3243) <= (layer7_outputs(141)) and (layer7_outputs(2647));
    layer8_outputs(3244) <= not(layer7_outputs(3605));
    layer8_outputs(3245) <= layer7_outputs(3867);
    layer8_outputs(3246) <= layer7_outputs(2533);
    layer8_outputs(3247) <= not(layer7_outputs(3836));
    layer8_outputs(3248) <= (layer7_outputs(2252)) xor (layer7_outputs(2869));
    layer8_outputs(3249) <= (layer7_outputs(2445)) xor (layer7_outputs(1083));
    layer8_outputs(3250) <= (layer7_outputs(2907)) and not (layer7_outputs(2146));
    layer8_outputs(3251) <= not((layer7_outputs(1340)) xor (layer7_outputs(2162)));
    layer8_outputs(3252) <= not(layer7_outputs(2012));
    layer8_outputs(3253) <= (layer7_outputs(72)) xor (layer7_outputs(2820));
    layer8_outputs(3254) <= layer7_outputs(2025);
    layer8_outputs(3255) <= (layer7_outputs(3648)) and not (layer7_outputs(2930));
    layer8_outputs(3256) <= layer7_outputs(447);
    layer8_outputs(3257) <= (layer7_outputs(3955)) and not (layer7_outputs(4303));
    layer8_outputs(3258) <= not((layer7_outputs(3756)) and (layer7_outputs(4698)));
    layer8_outputs(3259) <= not((layer7_outputs(4185)) and (layer7_outputs(4608)));
    layer8_outputs(3260) <= not((layer7_outputs(685)) and (layer7_outputs(4755)));
    layer8_outputs(3261) <= not((layer7_outputs(2502)) xor (layer7_outputs(297)));
    layer8_outputs(3262) <= not(layer7_outputs(2929));
    layer8_outputs(3263) <= layer7_outputs(968);
    layer8_outputs(3264) <= not(layer7_outputs(1237));
    layer8_outputs(3265) <= (layer7_outputs(3122)) xor (layer7_outputs(1126));
    layer8_outputs(3266) <= layer7_outputs(3166);
    layer8_outputs(3267) <= not((layer7_outputs(1118)) xor (layer7_outputs(649)));
    layer8_outputs(3268) <= not(layer7_outputs(4810));
    layer8_outputs(3269) <= (layer7_outputs(1964)) xor (layer7_outputs(350));
    layer8_outputs(3270) <= (layer7_outputs(2385)) xor (layer7_outputs(580));
    layer8_outputs(3271) <= not(layer7_outputs(160));
    layer8_outputs(3272) <= not(layer7_outputs(2979)) or (layer7_outputs(3847));
    layer8_outputs(3273) <= (layer7_outputs(4319)) and not (layer7_outputs(4951));
    layer8_outputs(3274) <= not((layer7_outputs(2086)) xor (layer7_outputs(1141)));
    layer8_outputs(3275) <= not(layer7_outputs(1677));
    layer8_outputs(3276) <= not(layer7_outputs(3232)) or (layer7_outputs(1189));
    layer8_outputs(3277) <= not((layer7_outputs(3673)) xor (layer7_outputs(5085)));
    layer8_outputs(3278) <= not(layer7_outputs(1395));
    layer8_outputs(3279) <= not(layer7_outputs(730));
    layer8_outputs(3280) <= not(layer7_outputs(1420));
    layer8_outputs(3281) <= not(layer7_outputs(1639));
    layer8_outputs(3282) <= not((layer7_outputs(4871)) xor (layer7_outputs(747)));
    layer8_outputs(3283) <= not(layer7_outputs(3829)) or (layer7_outputs(2272));
    layer8_outputs(3284) <= layer7_outputs(464);
    layer8_outputs(3285) <= not(layer7_outputs(1110)) or (layer7_outputs(911));
    layer8_outputs(3286) <= layer7_outputs(670);
    layer8_outputs(3287) <= (layer7_outputs(1873)) and not (layer7_outputs(1852));
    layer8_outputs(3288) <= not(layer7_outputs(1864)) or (layer7_outputs(1080));
    layer8_outputs(3289) <= (layer7_outputs(4004)) xor (layer7_outputs(311));
    layer8_outputs(3290) <= not(layer7_outputs(2923));
    layer8_outputs(3291) <= not(layer7_outputs(1101));
    layer8_outputs(3292) <= layer7_outputs(3205);
    layer8_outputs(3293) <= (layer7_outputs(2454)) and (layer7_outputs(4554));
    layer8_outputs(3294) <= not(layer7_outputs(166));
    layer8_outputs(3295) <= (layer7_outputs(2819)) or (layer7_outputs(1929));
    layer8_outputs(3296) <= not((layer7_outputs(1274)) xor (layer7_outputs(3677)));
    layer8_outputs(3297) <= not(layer7_outputs(1478));
    layer8_outputs(3298) <= layer7_outputs(2462);
    layer8_outputs(3299) <= layer7_outputs(3407);
    layer8_outputs(3300) <= not(layer7_outputs(3478)) or (layer7_outputs(4064));
    layer8_outputs(3301) <= (layer7_outputs(3977)) and not (layer7_outputs(1251));
    layer8_outputs(3302) <= layer7_outputs(5033);
    layer8_outputs(3303) <= layer7_outputs(2243);
    layer8_outputs(3304) <= layer7_outputs(1105);
    layer8_outputs(3305) <= (layer7_outputs(4139)) xor (layer7_outputs(2813));
    layer8_outputs(3306) <= not((layer7_outputs(4020)) xor (layer7_outputs(4531)));
    layer8_outputs(3307) <= not(layer7_outputs(2842));
    layer8_outputs(3308) <= layer7_outputs(4129);
    layer8_outputs(3309) <= not(layer7_outputs(831));
    layer8_outputs(3310) <= not(layer7_outputs(3893));
    layer8_outputs(3311) <= (layer7_outputs(796)) and (layer7_outputs(2575));
    layer8_outputs(3312) <= (layer7_outputs(965)) and (layer7_outputs(4205));
    layer8_outputs(3313) <= (layer7_outputs(116)) xor (layer7_outputs(618));
    layer8_outputs(3314) <= not((layer7_outputs(3530)) xor (layer7_outputs(2135)));
    layer8_outputs(3315) <= not(layer7_outputs(2114));
    layer8_outputs(3316) <= not((layer7_outputs(4029)) xor (layer7_outputs(4373)));
    layer8_outputs(3317) <= (layer7_outputs(3369)) xor (layer7_outputs(4513));
    layer8_outputs(3318) <= not(layer7_outputs(1276)) or (layer7_outputs(4743));
    layer8_outputs(3319) <= layer7_outputs(4667);
    layer8_outputs(3320) <= not(layer7_outputs(3076)) or (layer7_outputs(2644));
    layer8_outputs(3321) <= (layer7_outputs(4221)) xor (layer7_outputs(4192));
    layer8_outputs(3322) <= layer7_outputs(2293);
    layer8_outputs(3323) <= layer7_outputs(2288);
    layer8_outputs(3324) <= not(layer7_outputs(1956));
    layer8_outputs(3325) <= not((layer7_outputs(1417)) and (layer7_outputs(4711)));
    layer8_outputs(3326) <= (layer7_outputs(4951)) and not (layer7_outputs(961));
    layer8_outputs(3327) <= layer7_outputs(1383);
    layer8_outputs(3328) <= not(layer7_outputs(4078));
    layer8_outputs(3329) <= (layer7_outputs(644)) and (layer7_outputs(2466));
    layer8_outputs(3330) <= not((layer7_outputs(471)) xor (layer7_outputs(2530)));
    layer8_outputs(3331) <= layer7_outputs(386);
    layer8_outputs(3332) <= layer7_outputs(3537);
    layer8_outputs(3333) <= (layer7_outputs(2970)) xor (layer7_outputs(3151));
    layer8_outputs(3334) <= (layer7_outputs(1216)) xor (layer7_outputs(4606));
    layer8_outputs(3335) <= not(layer7_outputs(2732));
    layer8_outputs(3336) <= not(layer7_outputs(1421));
    layer8_outputs(3337) <= (layer7_outputs(3291)) xor (layer7_outputs(3224));
    layer8_outputs(3338) <= (layer7_outputs(3753)) xor (layer7_outputs(4824));
    layer8_outputs(3339) <= not(layer7_outputs(1487)) or (layer7_outputs(2451));
    layer8_outputs(3340) <= not((layer7_outputs(3244)) or (layer7_outputs(3964)));
    layer8_outputs(3341) <= layer7_outputs(1818);
    layer8_outputs(3342) <= not(layer7_outputs(3252));
    layer8_outputs(3343) <= (layer7_outputs(212)) and not (layer7_outputs(2721));
    layer8_outputs(3344) <= (layer7_outputs(3871)) xor (layer7_outputs(893));
    layer8_outputs(3345) <= (layer7_outputs(54)) xor (layer7_outputs(2749));
    layer8_outputs(3346) <= not(layer7_outputs(4539));
    layer8_outputs(3347) <= layer7_outputs(2857);
    layer8_outputs(3348) <= not(layer7_outputs(4912));
    layer8_outputs(3349) <= not(layer7_outputs(5013));
    layer8_outputs(3350) <= not(layer7_outputs(3109));
    layer8_outputs(3351) <= (layer7_outputs(3444)) and not (layer7_outputs(3924));
    layer8_outputs(3352) <= not(layer7_outputs(3329)) or (layer7_outputs(1897));
    layer8_outputs(3353) <= (layer7_outputs(156)) and (layer7_outputs(1301));
    layer8_outputs(3354) <= layer7_outputs(899);
    layer8_outputs(3355) <= layer7_outputs(1668);
    layer8_outputs(3356) <= not(layer7_outputs(2438));
    layer8_outputs(3357) <= not(layer7_outputs(4101)) or (layer7_outputs(902));
    layer8_outputs(3358) <= layer7_outputs(1609);
    layer8_outputs(3359) <= not(layer7_outputs(3608)) or (layer7_outputs(209));
    layer8_outputs(3360) <= (layer7_outputs(4395)) and not (layer7_outputs(4115));
    layer8_outputs(3361) <= layer7_outputs(928);
    layer8_outputs(3362) <= layer7_outputs(1618);
    layer8_outputs(3363) <= (layer7_outputs(4161)) xor (layer7_outputs(1211));
    layer8_outputs(3364) <= not((layer7_outputs(392)) xor (layer7_outputs(26)));
    layer8_outputs(3365) <= not((layer7_outputs(2888)) or (layer7_outputs(4294)));
    layer8_outputs(3366) <= not((layer7_outputs(1394)) or (layer7_outputs(3535)));
    layer8_outputs(3367) <= layer7_outputs(4130);
    layer8_outputs(3368) <= layer7_outputs(641);
    layer8_outputs(3369) <= (layer7_outputs(488)) and not (layer7_outputs(215));
    layer8_outputs(3370) <= (layer7_outputs(1854)) xor (layer7_outputs(2601));
    layer8_outputs(3371) <= not(layer7_outputs(224));
    layer8_outputs(3372) <= not(layer7_outputs(2172));
    layer8_outputs(3373) <= not((layer7_outputs(762)) xor (layer7_outputs(607)));
    layer8_outputs(3374) <= not((layer7_outputs(2473)) xor (layer7_outputs(3545)));
    layer8_outputs(3375) <= layer7_outputs(5095);
    layer8_outputs(3376) <= layer7_outputs(1323);
    layer8_outputs(3377) <= layer7_outputs(1332);
    layer8_outputs(3378) <= not((layer7_outputs(1531)) or (layer7_outputs(2716)));
    layer8_outputs(3379) <= (layer7_outputs(3111)) xor (layer7_outputs(2253));
    layer8_outputs(3380) <= (layer7_outputs(1629)) and (layer7_outputs(4954));
    layer8_outputs(3381) <= not(layer7_outputs(66));
    layer8_outputs(3382) <= not(layer7_outputs(1561));
    layer8_outputs(3383) <= (layer7_outputs(3261)) and (layer7_outputs(3861));
    layer8_outputs(3384) <= '1';
    layer8_outputs(3385) <= (layer7_outputs(3583)) or (layer7_outputs(2165));
    layer8_outputs(3386) <= (layer7_outputs(832)) or (layer7_outputs(1231));
    layer8_outputs(3387) <= not((layer7_outputs(3632)) or (layer7_outputs(2892)));
    layer8_outputs(3388) <= not((layer7_outputs(2064)) and (layer7_outputs(88)));
    layer8_outputs(3389) <= not(layer7_outputs(1933)) or (layer7_outputs(418));
    layer8_outputs(3390) <= not((layer7_outputs(1528)) xor (layer7_outputs(1584)));
    layer8_outputs(3391) <= layer7_outputs(3359);
    layer8_outputs(3392) <= (layer7_outputs(4471)) and not (layer7_outputs(4662));
    layer8_outputs(3393) <= layer7_outputs(988);
    layer8_outputs(3394) <= layer7_outputs(2410);
    layer8_outputs(3395) <= not(layer7_outputs(4893)) or (layer7_outputs(1422));
    layer8_outputs(3396) <= layer7_outputs(3295);
    layer8_outputs(3397) <= (layer7_outputs(1575)) and not (layer7_outputs(2683));
    layer8_outputs(3398) <= layer7_outputs(550);
    layer8_outputs(3399) <= (layer7_outputs(2005)) xor (layer7_outputs(2188));
    layer8_outputs(3400) <= (layer7_outputs(2563)) and not (layer7_outputs(194));
    layer8_outputs(3401) <= not((layer7_outputs(4404)) xor (layer7_outputs(3086)));
    layer8_outputs(3402) <= not(layer7_outputs(2023));
    layer8_outputs(3403) <= not(layer7_outputs(3683));
    layer8_outputs(3404) <= (layer7_outputs(1006)) and (layer7_outputs(4910));
    layer8_outputs(3405) <= (layer7_outputs(1280)) and (layer7_outputs(3953));
    layer8_outputs(3406) <= not(layer7_outputs(1608));
    layer8_outputs(3407) <= not(layer7_outputs(13));
    layer8_outputs(3408) <= not((layer7_outputs(1694)) and (layer7_outputs(4470)));
    layer8_outputs(3409) <= not(layer7_outputs(4813));
    layer8_outputs(3410) <= (layer7_outputs(2271)) and not (layer7_outputs(2567));
    layer8_outputs(3411) <= (layer7_outputs(870)) and (layer7_outputs(4600));
    layer8_outputs(3412) <= not((layer7_outputs(5040)) xor (layer7_outputs(2016)));
    layer8_outputs(3413) <= not(layer7_outputs(323));
    layer8_outputs(3414) <= (layer7_outputs(2674)) xor (layer7_outputs(651));
    layer8_outputs(3415) <= not(layer7_outputs(2272));
    layer8_outputs(3416) <= not(layer7_outputs(3816));
    layer8_outputs(3417) <= layer7_outputs(4793);
    layer8_outputs(3418) <= layer7_outputs(70);
    layer8_outputs(3419) <= (layer7_outputs(2140)) or (layer7_outputs(1816));
    layer8_outputs(3420) <= not(layer7_outputs(3754));
    layer8_outputs(3421) <= not(layer7_outputs(2135));
    layer8_outputs(3422) <= layer7_outputs(4771);
    layer8_outputs(3423) <= not((layer7_outputs(112)) xor (layer7_outputs(1181)));
    layer8_outputs(3424) <= layer7_outputs(3561);
    layer8_outputs(3425) <= not(layer7_outputs(2392));
    layer8_outputs(3426) <= layer7_outputs(3662);
    layer8_outputs(3427) <= (layer7_outputs(1928)) xor (layer7_outputs(2878));
    layer8_outputs(3428) <= layer7_outputs(4177);
    layer8_outputs(3429) <= (layer7_outputs(4573)) xor (layer7_outputs(2250));
    layer8_outputs(3430) <= not((layer7_outputs(5027)) and (layer7_outputs(4498)));
    layer8_outputs(3431) <= layer7_outputs(1227);
    layer8_outputs(3432) <= layer7_outputs(4299);
    layer8_outputs(3433) <= not(layer7_outputs(5101));
    layer8_outputs(3434) <= not((layer7_outputs(2232)) xor (layer7_outputs(2745)));
    layer8_outputs(3435) <= layer7_outputs(1649);
    layer8_outputs(3436) <= not(layer7_outputs(2158));
    layer8_outputs(3437) <= not(layer7_outputs(2122));
    layer8_outputs(3438) <= not(layer7_outputs(1378));
    layer8_outputs(3439) <= (layer7_outputs(2736)) and not (layer7_outputs(3794));
    layer8_outputs(3440) <= layer7_outputs(3592);
    layer8_outputs(3441) <= not(layer7_outputs(2988));
    layer8_outputs(3442) <= not(layer7_outputs(1672)) or (layer7_outputs(4314));
    layer8_outputs(3443) <= not(layer7_outputs(4671));
    layer8_outputs(3444) <= layer7_outputs(4019);
    layer8_outputs(3445) <= not((layer7_outputs(1496)) xor (layer7_outputs(1626)));
    layer8_outputs(3446) <= layer7_outputs(1633);
    layer8_outputs(3447) <= not((layer7_outputs(2807)) and (layer7_outputs(2150)));
    layer8_outputs(3448) <= (layer7_outputs(1856)) xor (layer7_outputs(572));
    layer8_outputs(3449) <= not(layer7_outputs(4785));
    layer8_outputs(3450) <= (layer7_outputs(3304)) xor (layer7_outputs(3826));
    layer8_outputs(3451) <= layer7_outputs(944);
    layer8_outputs(3452) <= (layer7_outputs(1318)) or (layer7_outputs(2951));
    layer8_outputs(3453) <= (layer7_outputs(3579)) xor (layer7_outputs(3620));
    layer8_outputs(3454) <= layer7_outputs(1520);
    layer8_outputs(3455) <= not(layer7_outputs(4257));
    layer8_outputs(3456) <= (layer7_outputs(671)) xor (layer7_outputs(4079));
    layer8_outputs(3457) <= not((layer7_outputs(5015)) or (layer7_outputs(2143)));
    layer8_outputs(3458) <= '1';
    layer8_outputs(3459) <= layer7_outputs(1599);
    layer8_outputs(3460) <= not(layer7_outputs(1604));
    layer8_outputs(3461) <= not((layer7_outputs(666)) or (layer7_outputs(1534)));
    layer8_outputs(3462) <= (layer7_outputs(2363)) or (layer7_outputs(3842));
    layer8_outputs(3463) <= not((layer7_outputs(4511)) and (layer7_outputs(3612)));
    layer8_outputs(3464) <= not(layer7_outputs(935));
    layer8_outputs(3465) <= not(layer7_outputs(4572));
    layer8_outputs(3466) <= not((layer7_outputs(3158)) and (layer7_outputs(4282)));
    layer8_outputs(3467) <= not(layer7_outputs(405)) or (layer7_outputs(2104));
    layer8_outputs(3468) <= (layer7_outputs(2469)) xor (layer7_outputs(1034));
    layer8_outputs(3469) <= not(layer7_outputs(3194));
    layer8_outputs(3470) <= not((layer7_outputs(4989)) xor (layer7_outputs(739)));
    layer8_outputs(3471) <= not((layer7_outputs(953)) xor (layer7_outputs(59)));
    layer8_outputs(3472) <= layer7_outputs(2798);
    layer8_outputs(3473) <= not((layer7_outputs(3156)) xor (layer7_outputs(1366)));
    layer8_outputs(3474) <= (layer7_outputs(1663)) xor (layer7_outputs(2142));
    layer8_outputs(3475) <= (layer7_outputs(4382)) and not (layer7_outputs(3049));
    layer8_outputs(3476) <= (layer7_outputs(2460)) xor (layer7_outputs(4384));
    layer8_outputs(3477) <= not(layer7_outputs(2812));
    layer8_outputs(3478) <= not(layer7_outputs(985)) or (layer7_outputs(842));
    layer8_outputs(3479) <= not(layer7_outputs(327));
    layer8_outputs(3480) <= (layer7_outputs(1109)) xor (layer7_outputs(36));
    layer8_outputs(3481) <= not(layer7_outputs(2297));
    layer8_outputs(3482) <= layer7_outputs(3138);
    layer8_outputs(3483) <= not(layer7_outputs(4533));
    layer8_outputs(3484) <= not(layer7_outputs(4021));
    layer8_outputs(3485) <= not(layer7_outputs(3900)) or (layer7_outputs(3366));
    layer8_outputs(3486) <= not(layer7_outputs(3628)) or (layer7_outputs(2997));
    layer8_outputs(3487) <= not((layer7_outputs(4023)) xor (layer7_outputs(7)));
    layer8_outputs(3488) <= not(layer7_outputs(19)) or (layer7_outputs(3325));
    layer8_outputs(3489) <= not(layer7_outputs(2960));
    layer8_outputs(3490) <= layer7_outputs(3157);
    layer8_outputs(3491) <= not(layer7_outputs(5109)) or (layer7_outputs(3209));
    layer8_outputs(3492) <= '0';
    layer8_outputs(3493) <= not(layer7_outputs(4588));
    layer8_outputs(3494) <= layer7_outputs(3336);
    layer8_outputs(3495) <= (layer7_outputs(404)) and not (layer7_outputs(863));
    layer8_outputs(3496) <= not(layer7_outputs(1066));
    layer8_outputs(3497) <= not((layer7_outputs(3101)) xor (layer7_outputs(647)));
    layer8_outputs(3498) <= not((layer7_outputs(2412)) xor (layer7_outputs(3452)));
    layer8_outputs(3499) <= layer7_outputs(3003);
    layer8_outputs(3500) <= not(layer7_outputs(589)) or (layer7_outputs(163));
    layer8_outputs(3501) <= (layer7_outputs(3210)) and (layer7_outputs(3633));
    layer8_outputs(3502) <= layer7_outputs(1068);
    layer8_outputs(3503) <= not((layer7_outputs(384)) xor (layer7_outputs(5038)));
    layer8_outputs(3504) <= (layer7_outputs(39)) xor (layer7_outputs(3765));
    layer8_outputs(3505) <= not(layer7_outputs(420));
    layer8_outputs(3506) <= not(layer7_outputs(1725));
    layer8_outputs(3507) <= layer7_outputs(1275);
    layer8_outputs(3508) <= not(layer7_outputs(1989));
    layer8_outputs(3509) <= not(layer7_outputs(3303));
    layer8_outputs(3510) <= (layer7_outputs(4260)) or (layer7_outputs(3002));
    layer8_outputs(3511) <= (layer7_outputs(179)) and not (layer7_outputs(317));
    layer8_outputs(3512) <= layer7_outputs(4147);
    layer8_outputs(3513) <= not(layer7_outputs(1793));
    layer8_outputs(3514) <= (layer7_outputs(1095)) and not (layer7_outputs(3077));
    layer8_outputs(3515) <= not(layer7_outputs(1657));
    layer8_outputs(3516) <= layer7_outputs(4911);
    layer8_outputs(3517) <= not(layer7_outputs(4372));
    layer8_outputs(3518) <= not(layer7_outputs(242));
    layer8_outputs(3519) <= not((layer7_outputs(3751)) and (layer7_outputs(3500)));
    layer8_outputs(3520) <= layer7_outputs(1647);
    layer8_outputs(3521) <= not(layer7_outputs(3294));
    layer8_outputs(3522) <= (layer7_outputs(269)) xor (layer7_outputs(3928));
    layer8_outputs(3523) <= layer7_outputs(3584);
    layer8_outputs(3524) <= not(layer7_outputs(4866)) or (layer7_outputs(838));
    layer8_outputs(3525) <= not(layer7_outputs(733));
    layer8_outputs(3526) <= layer7_outputs(3659);
    layer8_outputs(3527) <= layer7_outputs(4048);
    layer8_outputs(3528) <= layer7_outputs(5025);
    layer8_outputs(3529) <= layer7_outputs(1218);
    layer8_outputs(3530) <= (layer7_outputs(4619)) xor (layer7_outputs(879));
    layer8_outputs(3531) <= (layer7_outputs(3339)) or (layer7_outputs(2821));
    layer8_outputs(3532) <= not(layer7_outputs(4683));
    layer8_outputs(3533) <= not(layer7_outputs(2759));
    layer8_outputs(3534) <= (layer7_outputs(3095)) xor (layer7_outputs(5098));
    layer8_outputs(3535) <= not(layer7_outputs(5115));
    layer8_outputs(3536) <= not(layer7_outputs(3747));
    layer8_outputs(3537) <= not(layer7_outputs(3534)) or (layer7_outputs(2739));
    layer8_outputs(3538) <= '0';
    layer8_outputs(3539) <= not(layer7_outputs(2704));
    layer8_outputs(3540) <= (layer7_outputs(4628)) xor (layer7_outputs(3634));
    layer8_outputs(3541) <= not((layer7_outputs(957)) and (layer7_outputs(1160)));
    layer8_outputs(3542) <= layer7_outputs(983);
    layer8_outputs(3543) <= layer7_outputs(2325);
    layer8_outputs(3544) <= (layer7_outputs(828)) and not (layer7_outputs(2507));
    layer8_outputs(3545) <= (layer7_outputs(3562)) and (layer7_outputs(2497));
    layer8_outputs(3546) <= (layer7_outputs(1270)) xor (layer7_outputs(881));
    layer8_outputs(3547) <= (layer7_outputs(3647)) or (layer7_outputs(273));
    layer8_outputs(3548) <= layer7_outputs(1921);
    layer8_outputs(3549) <= not(layer7_outputs(4375));
    layer8_outputs(3550) <= not(layer7_outputs(3318));
    layer8_outputs(3551) <= layer7_outputs(1457);
    layer8_outputs(3552) <= not((layer7_outputs(3420)) xor (layer7_outputs(431)));
    layer8_outputs(3553) <= not(layer7_outputs(2808));
    layer8_outputs(3554) <= not(layer7_outputs(2093)) or (layer7_outputs(1637));
    layer8_outputs(3555) <= layer7_outputs(3859);
    layer8_outputs(3556) <= (layer7_outputs(1020)) or (layer7_outputs(2106));
    layer8_outputs(3557) <= not((layer7_outputs(4419)) xor (layer7_outputs(2635)));
    layer8_outputs(3558) <= not(layer7_outputs(4376)) or (layer7_outputs(2295));
    layer8_outputs(3559) <= (layer7_outputs(1258)) xor (layer7_outputs(2264));
    layer8_outputs(3560) <= (layer7_outputs(2701)) and not (layer7_outputs(3240));
    layer8_outputs(3561) <= (layer7_outputs(201)) xor (layer7_outputs(631));
    layer8_outputs(3562) <= not(layer7_outputs(3506));
    layer8_outputs(3563) <= layer7_outputs(4727);
    layer8_outputs(3564) <= (layer7_outputs(4020)) and (layer7_outputs(1409));
    layer8_outputs(3565) <= (layer7_outputs(2669)) and not (layer7_outputs(4259));
    layer8_outputs(3566) <= not(layer7_outputs(1923)) or (layer7_outputs(4646));
    layer8_outputs(3567) <= not(layer7_outputs(4049));
    layer8_outputs(3568) <= not((layer7_outputs(1951)) xor (layer7_outputs(3748)));
    layer8_outputs(3569) <= not(layer7_outputs(2170));
    layer8_outputs(3570) <= layer7_outputs(106);
    layer8_outputs(3571) <= layer7_outputs(1399);
    layer8_outputs(3572) <= not((layer7_outputs(607)) xor (layer7_outputs(3362)));
    layer8_outputs(3573) <= layer7_outputs(5066);
    layer8_outputs(3574) <= (layer7_outputs(4429)) xor (layer7_outputs(4229));
    layer8_outputs(3575) <= layer7_outputs(2678);
    layer8_outputs(3576) <= layer7_outputs(2504);
    layer8_outputs(3577) <= (layer7_outputs(91)) and not (layer7_outputs(4559));
    layer8_outputs(3578) <= not((layer7_outputs(49)) and (layer7_outputs(4209)));
    layer8_outputs(3579) <= not((layer7_outputs(2880)) or (layer7_outputs(3712)));
    layer8_outputs(3580) <= layer7_outputs(4760);
    layer8_outputs(3581) <= not(layer7_outputs(2209));
    layer8_outputs(3582) <= (layer7_outputs(3792)) and (layer7_outputs(4134));
    layer8_outputs(3583) <= layer7_outputs(1790);
    layer8_outputs(3584) <= not((layer7_outputs(596)) or (layer7_outputs(4616)));
    layer8_outputs(3585) <= not(layer7_outputs(3179));
    layer8_outputs(3586) <= not((layer7_outputs(1837)) and (layer7_outputs(1264)));
    layer8_outputs(3587) <= not(layer7_outputs(188));
    layer8_outputs(3588) <= layer7_outputs(4025);
    layer8_outputs(3589) <= layer7_outputs(1700);
    layer8_outputs(3590) <= not(layer7_outputs(387)) or (layer7_outputs(1731));
    layer8_outputs(3591) <= not(layer7_outputs(3934));
    layer8_outputs(3592) <= not(layer7_outputs(2311)) or (layer7_outputs(308));
    layer8_outputs(3593) <= '1';
    layer8_outputs(3594) <= not((layer7_outputs(4274)) xor (layer7_outputs(6)));
    layer8_outputs(3595) <= not((layer7_outputs(320)) xor (layer7_outputs(2514)));
    layer8_outputs(3596) <= not(layer7_outputs(314));
    layer8_outputs(3597) <= not(layer7_outputs(4155));
    layer8_outputs(3598) <= (layer7_outputs(3358)) and not (layer7_outputs(1403));
    layer8_outputs(3599) <= (layer7_outputs(347)) xor (layer7_outputs(749));
    layer8_outputs(3600) <= not(layer7_outputs(3558));
    layer8_outputs(3601) <= layer7_outputs(2920);
    layer8_outputs(3602) <= layer7_outputs(3572);
    layer8_outputs(3603) <= (layer7_outputs(271)) and not (layer7_outputs(4117));
    layer8_outputs(3604) <= (layer7_outputs(1606)) and not (layer7_outputs(2026));
    layer8_outputs(3605) <= not(layer7_outputs(3641)) or (layer7_outputs(468));
    layer8_outputs(3606) <= not((layer7_outputs(965)) xor (layer7_outputs(2516)));
    layer8_outputs(3607) <= not(layer7_outputs(2748));
    layer8_outputs(3608) <= (layer7_outputs(4935)) and not (layer7_outputs(1262));
    layer8_outputs(3609) <= (layer7_outputs(1581)) and not (layer7_outputs(1045));
    layer8_outputs(3610) <= not(layer7_outputs(4916));
    layer8_outputs(3611) <= (layer7_outputs(3646)) or (layer7_outputs(2744));
    layer8_outputs(3612) <= not((layer7_outputs(58)) or (layer7_outputs(3816)));
    layer8_outputs(3613) <= layer7_outputs(1513);
    layer8_outputs(3614) <= '0';
    layer8_outputs(3615) <= (layer7_outputs(276)) or (layer7_outputs(3374));
    layer8_outputs(3616) <= not(layer7_outputs(1641));
    layer8_outputs(3617) <= not(layer7_outputs(2046)) or (layer7_outputs(4992));
    layer8_outputs(3618) <= layer7_outputs(215);
    layer8_outputs(3619) <= (layer7_outputs(2441)) or (layer7_outputs(3082));
    layer8_outputs(3620) <= (layer7_outputs(1681)) and not (layer7_outputs(2164));
    layer8_outputs(3621) <= not(layer7_outputs(425));
    layer8_outputs(3622) <= not(layer7_outputs(791));
    layer8_outputs(3623) <= (layer7_outputs(1334)) xor (layer7_outputs(277));
    layer8_outputs(3624) <= layer7_outputs(2240);
    layer8_outputs(3625) <= not(layer7_outputs(4577)) or (layer7_outputs(3415));
    layer8_outputs(3626) <= layer7_outputs(3393);
    layer8_outputs(3627) <= not(layer7_outputs(2199));
    layer8_outputs(3628) <= layer7_outputs(4410);
    layer8_outputs(3629) <= not((layer7_outputs(400)) xor (layer7_outputs(950)));
    layer8_outputs(3630) <= not(layer7_outputs(144));
    layer8_outputs(3631) <= (layer7_outputs(1318)) and not (layer7_outputs(4006));
    layer8_outputs(3632) <= not(layer7_outputs(3295));
    layer8_outputs(3633) <= not(layer7_outputs(2066)) or (layer7_outputs(3877));
    layer8_outputs(3634) <= (layer7_outputs(3119)) xor (layer7_outputs(839));
    layer8_outputs(3635) <= not((layer7_outputs(2484)) xor (layer7_outputs(3675)));
    layer8_outputs(3636) <= not((layer7_outputs(351)) and (layer7_outputs(349)));
    layer8_outputs(3637) <= not(layer7_outputs(1784));
    layer8_outputs(3638) <= not(layer7_outputs(534)) or (layer7_outputs(759));
    layer8_outputs(3639) <= layer7_outputs(1825);
    layer8_outputs(3640) <= layer7_outputs(707);
    layer8_outputs(3641) <= layer7_outputs(1153);
    layer8_outputs(3642) <= layer7_outputs(3580);
    layer8_outputs(3643) <= not((layer7_outputs(4072)) xor (layer7_outputs(2486)));
    layer8_outputs(3644) <= layer7_outputs(2265);
    layer8_outputs(3645) <= (layer7_outputs(3636)) xor (layer7_outputs(4314));
    layer8_outputs(3646) <= not(layer7_outputs(474));
    layer8_outputs(3647) <= not(layer7_outputs(2313));
    layer8_outputs(3648) <= not(layer7_outputs(2679));
    layer8_outputs(3649) <= layer7_outputs(4231);
    layer8_outputs(3650) <= (layer7_outputs(4262)) xor (layer7_outputs(422));
    layer8_outputs(3651) <= (layer7_outputs(4194)) and not (layer7_outputs(3161));
    layer8_outputs(3652) <= (layer7_outputs(1239)) xor (layer7_outputs(3342));
    layer8_outputs(3653) <= layer7_outputs(2450);
    layer8_outputs(3654) <= not(layer7_outputs(3540));
    layer8_outputs(3655) <= not(layer7_outputs(1783));
    layer8_outputs(3656) <= (layer7_outputs(320)) and not (layer7_outputs(5055));
    layer8_outputs(3657) <= layer7_outputs(2984);
    layer8_outputs(3658) <= not(layer7_outputs(1453));
    layer8_outputs(3659) <= layer7_outputs(4657);
    layer8_outputs(3660) <= not(layer7_outputs(3994));
    layer8_outputs(3661) <= (layer7_outputs(936)) and not (layer7_outputs(2708));
    layer8_outputs(3662) <= not(layer7_outputs(2262));
    layer8_outputs(3663) <= not((layer7_outputs(5085)) xor (layer7_outputs(2735)));
    layer8_outputs(3664) <= not((layer7_outputs(4702)) or (layer7_outputs(2138)));
    layer8_outputs(3665) <= not(layer7_outputs(3749)) or (layer7_outputs(1636));
    layer8_outputs(3666) <= not((layer7_outputs(1732)) xor (layer7_outputs(1860)));
    layer8_outputs(3667) <= not(layer7_outputs(4230)) or (layer7_outputs(2541));
    layer8_outputs(3668) <= not(layer7_outputs(4245));
    layer8_outputs(3669) <= (layer7_outputs(122)) xor (layer7_outputs(3993));
    layer8_outputs(3670) <= layer7_outputs(416);
    layer8_outputs(3671) <= not(layer7_outputs(998)) or (layer7_outputs(4476));
    layer8_outputs(3672) <= not((layer7_outputs(3688)) or (layer7_outputs(3726)));
    layer8_outputs(3673) <= layer7_outputs(1234);
    layer8_outputs(3674) <= not((layer7_outputs(3706)) or (layer7_outputs(1237)));
    layer8_outputs(3675) <= not(layer7_outputs(326));
    layer8_outputs(3676) <= not(layer7_outputs(5079));
    layer8_outputs(3677) <= layer7_outputs(3240);
    layer8_outputs(3678) <= layer7_outputs(2860);
    layer8_outputs(3679) <= layer7_outputs(447);
    layer8_outputs(3680) <= not(layer7_outputs(982));
    layer8_outputs(3681) <= (layer7_outputs(3390)) xor (layer7_outputs(1941));
    layer8_outputs(3682) <= not(layer7_outputs(800)) or (layer7_outputs(3709));
    layer8_outputs(3683) <= layer7_outputs(1985);
    layer8_outputs(3684) <= layer7_outputs(360);
    layer8_outputs(3685) <= (layer7_outputs(2985)) xor (layer7_outputs(3625));
    layer8_outputs(3686) <= not((layer7_outputs(644)) and (layer7_outputs(3315)));
    layer8_outputs(3687) <= not(layer7_outputs(3599));
    layer8_outputs(3688) <= (layer7_outputs(161)) and (layer7_outputs(2676));
    layer8_outputs(3689) <= (layer7_outputs(1842)) and not (layer7_outputs(2925));
    layer8_outputs(3690) <= not(layer7_outputs(3686));
    layer8_outputs(3691) <= not(layer7_outputs(1562));
    layer8_outputs(3692) <= (layer7_outputs(4416)) xor (layer7_outputs(1397));
    layer8_outputs(3693) <= not(layer7_outputs(807));
    layer8_outputs(3694) <= (layer7_outputs(1269)) xor (layer7_outputs(2));
    layer8_outputs(3695) <= not((layer7_outputs(3379)) xor (layer7_outputs(4227)));
    layer8_outputs(3696) <= (layer7_outputs(3266)) and (layer7_outputs(4306));
    layer8_outputs(3697) <= not(layer7_outputs(4296));
    layer8_outputs(3698) <= layer7_outputs(1519);
    layer8_outputs(3699) <= (layer7_outputs(1540)) xor (layer7_outputs(2425));
    layer8_outputs(3700) <= not((layer7_outputs(4743)) and (layer7_outputs(1146)));
    layer8_outputs(3701) <= not(layer7_outputs(1867));
    layer8_outputs(3702) <= not(layer7_outputs(4114));
    layer8_outputs(3703) <= not(layer7_outputs(1464));
    layer8_outputs(3704) <= not(layer7_outputs(4764));
    layer8_outputs(3705) <= not(layer7_outputs(2317));
    layer8_outputs(3706) <= not((layer7_outputs(398)) or (layer7_outputs(1529)));
    layer8_outputs(3707) <= layer7_outputs(4635);
    layer8_outputs(3708) <= layer7_outputs(4958);
    layer8_outputs(3709) <= not(layer7_outputs(1528));
    layer8_outputs(3710) <= not(layer7_outputs(82)) or (layer7_outputs(2696));
    layer8_outputs(3711) <= not(layer7_outputs(1678));
    layer8_outputs(3712) <= layer7_outputs(470);
    layer8_outputs(3713) <= not((layer7_outputs(3854)) and (layer7_outputs(3134)));
    layer8_outputs(3714) <= (layer7_outputs(332)) or (layer7_outputs(2880));
    layer8_outputs(3715) <= (layer7_outputs(543)) xor (layer7_outputs(4919));
    layer8_outputs(3716) <= not((layer7_outputs(4985)) xor (layer7_outputs(375)));
    layer8_outputs(3717) <= not((layer7_outputs(2733)) xor (layer7_outputs(4767)));
    layer8_outputs(3718) <= (layer7_outputs(4308)) or (layer7_outputs(4309));
    layer8_outputs(3719) <= (layer7_outputs(3027)) and (layer7_outputs(2670));
    layer8_outputs(3720) <= '1';
    layer8_outputs(3721) <= (layer7_outputs(3)) and not (layer7_outputs(3602));
    layer8_outputs(3722) <= not(layer7_outputs(4162));
    layer8_outputs(3723) <= not((layer7_outputs(4891)) and (layer7_outputs(2379)));
    layer8_outputs(3724) <= (layer7_outputs(4595)) xor (layer7_outputs(2629));
    layer8_outputs(3725) <= not(layer7_outputs(1814));
    layer8_outputs(3726) <= layer7_outputs(3271);
    layer8_outputs(3727) <= not((layer7_outputs(5034)) or (layer7_outputs(371)));
    layer8_outputs(3728) <= (layer7_outputs(922)) or (layer7_outputs(2533));
    layer8_outputs(3729) <= not(layer7_outputs(3851));
    layer8_outputs(3730) <= (layer7_outputs(2346)) or (layer7_outputs(3267));
    layer8_outputs(3731) <= layer7_outputs(4357);
    layer8_outputs(3732) <= not(layer7_outputs(4961));
    layer8_outputs(3733) <= not(layer7_outputs(3872));
    layer8_outputs(3734) <= not(layer7_outputs(740));
    layer8_outputs(3735) <= layer7_outputs(3208);
    layer8_outputs(3736) <= (layer7_outputs(5061)) xor (layer7_outputs(1458));
    layer8_outputs(3737) <= layer7_outputs(1222);
    layer8_outputs(3738) <= not(layer7_outputs(4437));
    layer8_outputs(3739) <= not(layer7_outputs(3045));
    layer8_outputs(3740) <= layer7_outputs(3731);
    layer8_outputs(3741) <= not((layer7_outputs(1745)) xor (layer7_outputs(2855)));
    layer8_outputs(3742) <= not(layer7_outputs(94));
    layer8_outputs(3743) <= (layer7_outputs(592)) xor (layer7_outputs(2875));
    layer8_outputs(3744) <= not(layer7_outputs(4735)) or (layer7_outputs(3790));
    layer8_outputs(3745) <= layer7_outputs(2741);
    layer8_outputs(3746) <= not((layer7_outputs(4275)) xor (layer7_outputs(4289)));
    layer8_outputs(3747) <= not((layer7_outputs(4667)) xor (layer7_outputs(616)));
    layer8_outputs(3748) <= layer7_outputs(4123);
    layer8_outputs(3749) <= not(layer7_outputs(2477));
    layer8_outputs(3750) <= not(layer7_outputs(3571));
    layer8_outputs(3751) <= not(layer7_outputs(774)) or (layer7_outputs(5061));
    layer8_outputs(3752) <= not(layer7_outputs(1295));
    layer8_outputs(3753) <= not((layer7_outputs(4165)) or (layer7_outputs(2777)));
    layer8_outputs(3754) <= not(layer7_outputs(2539));
    layer8_outputs(3755) <= not((layer7_outputs(67)) and (layer7_outputs(4173)));
    layer8_outputs(3756) <= not((layer7_outputs(2324)) xor (layer7_outputs(4377)));
    layer8_outputs(3757) <= layer7_outputs(1904);
    layer8_outputs(3758) <= not((layer7_outputs(2596)) or (layer7_outputs(2191)));
    layer8_outputs(3759) <= layer7_outputs(2254);
    layer8_outputs(3760) <= layer7_outputs(1369);
    layer8_outputs(3761) <= (layer7_outputs(344)) and not (layer7_outputs(1807));
    layer8_outputs(3762) <= not(layer7_outputs(1823));
    layer8_outputs(3763) <= (layer7_outputs(4150)) xor (layer7_outputs(2806));
    layer8_outputs(3764) <= not((layer7_outputs(1871)) xor (layer7_outputs(4181)));
    layer8_outputs(3765) <= (layer7_outputs(4659)) and not (layer7_outputs(4514));
    layer8_outputs(3766) <= layer7_outputs(3878);
    layer8_outputs(3767) <= not((layer7_outputs(3958)) xor (layer7_outputs(2482)));
    layer8_outputs(3768) <= (layer7_outputs(3303)) or (layer7_outputs(539));
    layer8_outputs(3769) <= not(layer7_outputs(1648));
    layer8_outputs(3770) <= layer7_outputs(2551);
    layer8_outputs(3771) <= (layer7_outputs(5079)) and (layer7_outputs(4472));
    layer8_outputs(3772) <= not(layer7_outputs(323));
    layer8_outputs(3773) <= not(layer7_outputs(5099)) or (layer7_outputs(4946));
    layer8_outputs(3774) <= not(layer7_outputs(3024)) or (layer7_outputs(3947));
    layer8_outputs(3775) <= (layer7_outputs(2013)) and not (layer7_outputs(435));
    layer8_outputs(3776) <= layer7_outputs(221);
    layer8_outputs(3777) <= (layer7_outputs(5119)) xor (layer7_outputs(2698));
    layer8_outputs(3778) <= (layer7_outputs(1747)) xor (layer7_outputs(1886));
    layer8_outputs(3779) <= not(layer7_outputs(628)) or (layer7_outputs(2753));
    layer8_outputs(3780) <= layer7_outputs(2848);
    layer8_outputs(3781) <= (layer7_outputs(2161)) and not (layer7_outputs(2617));
    layer8_outputs(3782) <= layer7_outputs(1690);
    layer8_outputs(3783) <= not(layer7_outputs(825));
    layer8_outputs(3784) <= not((layer7_outputs(3738)) xor (layer7_outputs(2080)));
    layer8_outputs(3785) <= layer7_outputs(3682);
    layer8_outputs(3786) <= layer7_outputs(548);
    layer8_outputs(3787) <= not((layer7_outputs(1828)) or (layer7_outputs(2392)));
    layer8_outputs(3788) <= layer7_outputs(4193);
    layer8_outputs(3789) <= not((layer7_outputs(2818)) and (layer7_outputs(4968)));
    layer8_outputs(3790) <= (layer7_outputs(72)) or (layer7_outputs(4148));
    layer8_outputs(3791) <= layer7_outputs(4896);
    layer8_outputs(3792) <= (layer7_outputs(3910)) and not (layer7_outputs(1494));
    layer8_outputs(3793) <= layer7_outputs(3037);
    layer8_outputs(3794) <= not(layer7_outputs(1680));
    layer8_outputs(3795) <= not(layer7_outputs(2075));
    layer8_outputs(3796) <= (layer7_outputs(3182)) xor (layer7_outputs(1247));
    layer8_outputs(3797) <= not((layer7_outputs(2642)) xor (layer7_outputs(138)));
    layer8_outputs(3798) <= layer7_outputs(492);
    layer8_outputs(3799) <= (layer7_outputs(2840)) xor (layer7_outputs(2216));
    layer8_outputs(3800) <= not(layer7_outputs(2386));
    layer8_outputs(3801) <= layer7_outputs(3541);
    layer8_outputs(3802) <= '0';
    layer8_outputs(3803) <= (layer7_outputs(1793)) or (layer7_outputs(3113));
    layer8_outputs(3804) <= not(layer7_outputs(1294));
    layer8_outputs(3805) <= (layer7_outputs(2278)) xor (layer7_outputs(2783));
    layer8_outputs(3806) <= not(layer7_outputs(2556));
    layer8_outputs(3807) <= layer7_outputs(4007);
    layer8_outputs(3808) <= not(layer7_outputs(2383)) or (layer7_outputs(4595));
    layer8_outputs(3809) <= (layer7_outputs(2335)) xor (layer7_outputs(1281));
    layer8_outputs(3810) <= not(layer7_outputs(1998)) or (layer7_outputs(4305));
    layer8_outputs(3811) <= not(layer7_outputs(733));
    layer8_outputs(3812) <= not(layer7_outputs(4973));
    layer8_outputs(3813) <= not((layer7_outputs(2922)) xor (layer7_outputs(3546)));
    layer8_outputs(3814) <= layer7_outputs(377);
    layer8_outputs(3815) <= (layer7_outputs(4936)) and not (layer7_outputs(3185));
    layer8_outputs(3816) <= layer7_outputs(43);
    layer8_outputs(3817) <= (layer7_outputs(1380)) xor (layer7_outputs(3260));
    layer8_outputs(3818) <= '0';
    layer8_outputs(3819) <= not(layer7_outputs(768)) or (layer7_outputs(4287));
    layer8_outputs(3820) <= (layer7_outputs(3515)) and (layer7_outputs(1941));
    layer8_outputs(3821) <= layer7_outputs(2070);
    layer8_outputs(3822) <= (layer7_outputs(1737)) xor (layer7_outputs(293));
    layer8_outputs(3823) <= layer7_outputs(3927);
    layer8_outputs(3824) <= (layer7_outputs(502)) xor (layer7_outputs(5031));
    layer8_outputs(3825) <= (layer7_outputs(2236)) and not (layer7_outputs(4527));
    layer8_outputs(3826) <= not((layer7_outputs(520)) xor (layer7_outputs(596)));
    layer8_outputs(3827) <= (layer7_outputs(3928)) xor (layer7_outputs(526));
    layer8_outputs(3828) <= (layer7_outputs(2035)) and (layer7_outputs(878));
    layer8_outputs(3829) <= layer7_outputs(3537);
    layer8_outputs(3830) <= (layer7_outputs(4985)) xor (layer7_outputs(571));
    layer8_outputs(3831) <= not(layer7_outputs(4261));
    layer8_outputs(3832) <= layer7_outputs(4580);
    layer8_outputs(3833) <= (layer7_outputs(317)) and (layer7_outputs(3894));
    layer8_outputs(3834) <= layer7_outputs(4740);
    layer8_outputs(3835) <= not(layer7_outputs(4837));
    layer8_outputs(3836) <= layer7_outputs(3885);
    layer8_outputs(3837) <= not(layer7_outputs(2137)) or (layer7_outputs(3055));
    layer8_outputs(3838) <= not((layer7_outputs(4746)) xor (layer7_outputs(1949)));
    layer8_outputs(3839) <= not(layer7_outputs(1876)) or (layer7_outputs(848));
    layer8_outputs(3840) <= not(layer7_outputs(2225));
    layer8_outputs(3841) <= not((layer7_outputs(3035)) xor (layer7_outputs(3582)));
    layer8_outputs(3842) <= (layer7_outputs(2150)) or (layer7_outputs(5017));
    layer8_outputs(3843) <= (layer7_outputs(704)) xor (layer7_outputs(1178));
    layer8_outputs(3844) <= (layer7_outputs(253)) and not (layer7_outputs(3048));
    layer8_outputs(3845) <= not(layer7_outputs(3042)) or (layer7_outputs(2693));
    layer8_outputs(3846) <= not(layer7_outputs(2237));
    layer8_outputs(3847) <= (layer7_outputs(3503)) and not (layer7_outputs(968));
    layer8_outputs(3848) <= layer7_outputs(4692);
    layer8_outputs(3849) <= (layer7_outputs(4240)) and not (layer7_outputs(3387));
    layer8_outputs(3850) <= layer7_outputs(2342);
    layer8_outputs(3851) <= layer7_outputs(204);
    layer8_outputs(3852) <= not(layer7_outputs(210));
    layer8_outputs(3853) <= layer7_outputs(501);
    layer8_outputs(3854) <= not(layer7_outputs(3496)) or (layer7_outputs(4179));
    layer8_outputs(3855) <= not((layer7_outputs(3471)) or (layer7_outputs(4838)));
    layer8_outputs(3856) <= layer7_outputs(1267);
    layer8_outputs(3857) <= not(layer7_outputs(552));
    layer8_outputs(3858) <= not(layer7_outputs(3840));
    layer8_outputs(3859) <= layer7_outputs(79);
    layer8_outputs(3860) <= not((layer7_outputs(2302)) xor (layer7_outputs(4083)));
    layer8_outputs(3861) <= (layer7_outputs(1867)) xor (layer7_outputs(3497));
    layer8_outputs(3862) <= not(layer7_outputs(1397));
    layer8_outputs(3863) <= layer7_outputs(2077);
    layer8_outputs(3864) <= (layer7_outputs(4880)) and (layer7_outputs(4999));
    layer8_outputs(3865) <= layer7_outputs(1147);
    layer8_outputs(3866) <= (layer7_outputs(2474)) or (layer7_outputs(2409));
    layer8_outputs(3867) <= (layer7_outputs(3686)) xor (layer7_outputs(1670));
    layer8_outputs(3868) <= not(layer7_outputs(708));
    layer8_outputs(3869) <= layer7_outputs(1788);
    layer8_outputs(3870) <= not(layer7_outputs(1238)) or (layer7_outputs(3769));
    layer8_outputs(3871) <= not((layer7_outputs(1962)) xor (layer7_outputs(3045)));
    layer8_outputs(3872) <= not(layer7_outputs(2194));
    layer8_outputs(3873) <= (layer7_outputs(549)) and (layer7_outputs(1731));
    layer8_outputs(3874) <= layer7_outputs(4620);
    layer8_outputs(3875) <= (layer7_outputs(3866)) and not (layer7_outputs(4607));
    layer8_outputs(3876) <= not((layer7_outputs(296)) xor (layer7_outputs(4909)));
    layer8_outputs(3877) <= not(layer7_outputs(4389));
    layer8_outputs(3878) <= layer7_outputs(1220);
    layer8_outputs(3879) <= not((layer7_outputs(948)) xor (layer7_outputs(87)));
    layer8_outputs(3880) <= not(layer7_outputs(3749));
    layer8_outputs(3881) <= (layer7_outputs(1482)) xor (layer7_outputs(1885));
    layer8_outputs(3882) <= not((layer7_outputs(1419)) and (layer7_outputs(4159)));
    layer8_outputs(3883) <= layer7_outputs(1476);
    layer8_outputs(3884) <= not((layer7_outputs(1009)) or (layer7_outputs(3875)));
    layer8_outputs(3885) <= layer7_outputs(3547);
    layer8_outputs(3886) <= not((layer7_outputs(4308)) xor (layer7_outputs(4704)));
    layer8_outputs(3887) <= (layer7_outputs(2928)) xor (layer7_outputs(2014));
    layer8_outputs(3888) <= (layer7_outputs(3453)) xor (layer7_outputs(2265));
    layer8_outputs(3889) <= not((layer7_outputs(4349)) xor (layer7_outputs(2644)));
    layer8_outputs(3890) <= not(layer7_outputs(3974));
    layer8_outputs(3891) <= (layer7_outputs(2446)) xor (layer7_outputs(3759));
    layer8_outputs(3892) <= layer7_outputs(3335);
    layer8_outputs(3893) <= not((layer7_outputs(819)) xor (layer7_outputs(727)));
    layer8_outputs(3894) <= not((layer7_outputs(949)) and (layer7_outputs(4805)));
    layer8_outputs(3895) <= (layer7_outputs(491)) xor (layer7_outputs(4371));
    layer8_outputs(3896) <= (layer7_outputs(2868)) xor (layer7_outputs(3801));
    layer8_outputs(3897) <= (layer7_outputs(741)) and (layer7_outputs(2447));
    layer8_outputs(3898) <= layer7_outputs(2643);
    layer8_outputs(3899) <= (layer7_outputs(1256)) and (layer7_outputs(5014));
    layer8_outputs(3900) <= not((layer7_outputs(101)) xor (layer7_outputs(574)));
    layer8_outputs(3901) <= not(layer7_outputs(4369));
    layer8_outputs(3902) <= layer7_outputs(1780);
    layer8_outputs(3903) <= layer7_outputs(3739);
    layer8_outputs(3904) <= not(layer7_outputs(859));
    layer8_outputs(3905) <= (layer7_outputs(514)) or (layer7_outputs(1795));
    layer8_outputs(3906) <= layer7_outputs(1508);
    layer8_outputs(3907) <= layer7_outputs(4415);
    layer8_outputs(3908) <= not(layer7_outputs(4971));
    layer8_outputs(3909) <= not(layer7_outputs(3901));
    layer8_outputs(3910) <= (layer7_outputs(2534)) or (layer7_outputs(3563));
    layer8_outputs(3911) <= layer7_outputs(4539);
    layer8_outputs(3912) <= layer7_outputs(4901);
    layer8_outputs(3913) <= not(layer7_outputs(2038));
    layer8_outputs(3914) <= (layer7_outputs(3422)) and (layer7_outputs(364));
    layer8_outputs(3915) <= layer7_outputs(2839);
    layer8_outputs(3916) <= not(layer7_outputs(4404));
    layer8_outputs(3917) <= not(layer7_outputs(1608)) or (layer7_outputs(3417));
    layer8_outputs(3918) <= (layer7_outputs(5073)) or (layer7_outputs(2042));
    layer8_outputs(3919) <= (layer7_outputs(5000)) and not (layer7_outputs(3734));
    layer8_outputs(3920) <= layer7_outputs(3354);
    layer8_outputs(3921) <= (layer7_outputs(3312)) and not (layer7_outputs(2935));
    layer8_outputs(3922) <= not((layer7_outputs(3915)) xor (layer7_outputs(5074)));
    layer8_outputs(3923) <= not(layer7_outputs(4693)) or (layer7_outputs(2934));
    layer8_outputs(3924) <= not(layer7_outputs(1007));
    layer8_outputs(3925) <= layer7_outputs(971);
    layer8_outputs(3926) <= layer7_outputs(413);
    layer8_outputs(3927) <= (layer7_outputs(1140)) and not (layer7_outputs(1958));
    layer8_outputs(3928) <= (layer7_outputs(3461)) xor (layer7_outputs(1979));
    layer8_outputs(3929) <= not(layer7_outputs(2009));
    layer8_outputs(3930) <= layer7_outputs(4257);
    layer8_outputs(3931) <= not(layer7_outputs(902));
    layer8_outputs(3932) <= (layer7_outputs(2579)) and (layer7_outputs(1752));
    layer8_outputs(3933) <= layer7_outputs(2020);
    layer8_outputs(3934) <= (layer7_outputs(2459)) and not (layer7_outputs(4235));
    layer8_outputs(3935) <= not(layer7_outputs(2487));
    layer8_outputs(3936) <= not(layer7_outputs(3821));
    layer8_outputs(3937) <= not(layer7_outputs(5048));
    layer8_outputs(3938) <= not(layer7_outputs(971));
    layer8_outputs(3939) <= layer7_outputs(4118);
    layer8_outputs(3940) <= not(layer7_outputs(1024)) or (layer7_outputs(2023));
    layer8_outputs(3941) <= layer7_outputs(3233);
    layer8_outputs(3942) <= layer7_outputs(2931);
    layer8_outputs(3943) <= layer7_outputs(2774);
    layer8_outputs(3944) <= not(layer7_outputs(355));
    layer8_outputs(3945) <= (layer7_outputs(4898)) xor (layer7_outputs(1241));
    layer8_outputs(3946) <= not((layer7_outputs(600)) and (layer7_outputs(3386)));
    layer8_outputs(3947) <= (layer7_outputs(4684)) xor (layer7_outputs(1374));
    layer8_outputs(3948) <= (layer7_outputs(2009)) and not (layer7_outputs(3701));
    layer8_outputs(3949) <= not(layer7_outputs(1410));
    layer8_outputs(3950) <= (layer7_outputs(1653)) or (layer7_outputs(2706));
    layer8_outputs(3951) <= not(layer7_outputs(3677));
    layer8_outputs(3952) <= (layer7_outputs(4640)) and (layer7_outputs(1302));
    layer8_outputs(3953) <= not(layer7_outputs(4639)) or (layer7_outputs(791));
    layer8_outputs(3954) <= not((layer7_outputs(4601)) xor (layer7_outputs(423)));
    layer8_outputs(3955) <= not(layer7_outputs(2102));
    layer8_outputs(3956) <= not(layer7_outputs(3531)) or (layer7_outputs(3058));
    layer8_outputs(3957) <= (layer7_outputs(3164)) and not (layer7_outputs(1599));
    layer8_outputs(3958) <= layer7_outputs(2754);
    layer8_outputs(3959) <= layer7_outputs(3373);
    layer8_outputs(3960) <= not(layer7_outputs(3933));
    layer8_outputs(3961) <= not(layer7_outputs(4237));
    layer8_outputs(3962) <= layer7_outputs(3175);
    layer8_outputs(3963) <= not(layer7_outputs(3890));
    layer8_outputs(3964) <= layer7_outputs(1945);
    layer8_outputs(3965) <= (layer7_outputs(3497)) and not (layer7_outputs(2837));
    layer8_outputs(3966) <= layer7_outputs(3826);
    layer8_outputs(3967) <= layer7_outputs(3484);
    layer8_outputs(3968) <= not(layer7_outputs(33));
    layer8_outputs(3969) <= (layer7_outputs(1861)) xor (layer7_outputs(3152));
    layer8_outputs(3970) <= not((layer7_outputs(504)) xor (layer7_outputs(4778)));
    layer8_outputs(3971) <= layer7_outputs(1363);
    layer8_outputs(3972) <= layer7_outputs(2294);
    layer8_outputs(3973) <= not(layer7_outputs(239)) or (layer7_outputs(4406));
    layer8_outputs(3974) <= not(layer7_outputs(3561));
    layer8_outputs(3975) <= layer7_outputs(4902);
    layer8_outputs(3976) <= (layer7_outputs(4934)) and not (layer7_outputs(4519));
    layer8_outputs(3977) <= (layer7_outputs(1182)) and not (layer7_outputs(1110));
    layer8_outputs(3978) <= layer7_outputs(4794);
    layer8_outputs(3979) <= not(layer7_outputs(2608));
    layer8_outputs(3980) <= not(layer7_outputs(1312)) or (layer7_outputs(1387));
    layer8_outputs(3981) <= (layer7_outputs(3940)) or (layer7_outputs(1331));
    layer8_outputs(3982) <= not((layer7_outputs(1045)) xor (layer7_outputs(1748)));
    layer8_outputs(3983) <= (layer7_outputs(385)) and not (layer7_outputs(1429));
    layer8_outputs(3984) <= not(layer7_outputs(3722));
    layer8_outputs(3985) <= layer7_outputs(4876);
    layer8_outputs(3986) <= layer7_outputs(1679);
    layer8_outputs(3987) <= not((layer7_outputs(504)) or (layer7_outputs(901)));
    layer8_outputs(3988) <= not(layer7_outputs(4713));
    layer8_outputs(3989) <= (layer7_outputs(5004)) and not (layer7_outputs(191));
    layer8_outputs(3990) <= not(layer7_outputs(3241)) or (layer7_outputs(1468));
    layer8_outputs(3991) <= not((layer7_outputs(4083)) xor (layer7_outputs(4325)));
    layer8_outputs(3992) <= not(layer7_outputs(3823));
    layer8_outputs(3993) <= not(layer7_outputs(4390)) or (layer7_outputs(851));
    layer8_outputs(3994) <= layer7_outputs(1934);
    layer8_outputs(3995) <= (layer7_outputs(2557)) xor (layer7_outputs(3211));
    layer8_outputs(3996) <= not(layer7_outputs(3075));
    layer8_outputs(3997) <= not(layer7_outputs(2152));
    layer8_outputs(3998) <= not(layer7_outputs(4478));
    layer8_outputs(3999) <= layer7_outputs(4124);
    layer8_outputs(4000) <= not((layer7_outputs(1572)) xor (layer7_outputs(2166)));
    layer8_outputs(4001) <= not(layer7_outputs(484));
    layer8_outputs(4002) <= not(layer7_outputs(2797));
    layer8_outputs(4003) <= (layer7_outputs(1088)) and not (layer7_outputs(2520));
    layer8_outputs(4004) <= (layer7_outputs(4015)) xor (layer7_outputs(4065));
    layer8_outputs(4005) <= (layer7_outputs(685)) xor (layer7_outputs(315));
    layer8_outputs(4006) <= layer7_outputs(3252);
    layer8_outputs(4007) <= (layer7_outputs(403)) and not (layer7_outputs(1884));
    layer8_outputs(4008) <= (layer7_outputs(2709)) and (layer7_outputs(4121));
    layer8_outputs(4009) <= layer7_outputs(2167);
    layer8_outputs(4010) <= (layer7_outputs(1508)) and not (layer7_outputs(647));
    layer8_outputs(4011) <= (layer7_outputs(4146)) and not (layer7_outputs(240));
    layer8_outputs(4012) <= not(layer7_outputs(3025)) or (layer7_outputs(2279));
    layer8_outputs(4013) <= (layer7_outputs(3319)) xor (layer7_outputs(2651));
    layer8_outputs(4014) <= (layer7_outputs(4715)) and (layer7_outputs(1393));
    layer8_outputs(4015) <= not(layer7_outputs(2772));
    layer8_outputs(4016) <= not(layer7_outputs(756));
    layer8_outputs(4017) <= not((layer7_outputs(2483)) xor (layer7_outputs(4387)));
    layer8_outputs(4018) <= layer7_outputs(622);
    layer8_outputs(4019) <= not((layer7_outputs(2800)) xor (layer7_outputs(5106)));
    layer8_outputs(4020) <= not(layer7_outputs(617)) or (layer7_outputs(5013));
    layer8_outputs(4021) <= layer7_outputs(1938);
    layer8_outputs(4022) <= (layer7_outputs(2348)) xor (layer7_outputs(1322));
    layer8_outputs(4023) <= not((layer7_outputs(1329)) and (layer7_outputs(2186)));
    layer8_outputs(4024) <= not(layer7_outputs(4756));
    layer8_outputs(4025) <= layer7_outputs(339);
    layer8_outputs(4026) <= (layer7_outputs(1401)) or (layer7_outputs(636));
    layer8_outputs(4027) <= layer7_outputs(5116);
    layer8_outputs(4028) <= not((layer7_outputs(4272)) or (layer7_outputs(4081)));
    layer8_outputs(4029) <= not(layer7_outputs(1435));
    layer8_outputs(4030) <= layer7_outputs(289);
    layer8_outputs(4031) <= (layer7_outputs(1094)) and not (layer7_outputs(1679));
    layer8_outputs(4032) <= layer7_outputs(1248);
    layer8_outputs(4033) <= layer7_outputs(3174);
    layer8_outputs(4034) <= not(layer7_outputs(3585));
    layer8_outputs(4035) <= not(layer7_outputs(3799)) or (layer7_outputs(2592));
    layer8_outputs(4036) <= layer7_outputs(3249);
    layer8_outputs(4037) <= not((layer7_outputs(3314)) xor (layer7_outputs(940)));
    layer8_outputs(4038) <= not(layer7_outputs(3439)) or (layer7_outputs(1063));
    layer8_outputs(4039) <= layer7_outputs(1494);
    layer8_outputs(4040) <= layer7_outputs(3308);
    layer8_outputs(4041) <= (layer7_outputs(775)) and not (layer7_outputs(3812));
    layer8_outputs(4042) <= not(layer7_outputs(2068));
    layer8_outputs(4043) <= not(layer7_outputs(1634));
    layer8_outputs(4044) <= (layer7_outputs(4106)) xor (layer7_outputs(3664));
    layer8_outputs(4045) <= (layer7_outputs(1903)) xor (layer7_outputs(3827));
    layer8_outputs(4046) <= not(layer7_outputs(2598));
    layer8_outputs(4047) <= (layer7_outputs(1641)) and (layer7_outputs(2889));
    layer8_outputs(4048) <= not((layer7_outputs(600)) xor (layer7_outputs(3590)));
    layer8_outputs(4049) <= layer7_outputs(5043);
    layer8_outputs(4050) <= not((layer7_outputs(2242)) xor (layer7_outputs(1493)));
    layer8_outputs(4051) <= layer7_outputs(2608);
    layer8_outputs(4052) <= not((layer7_outputs(4477)) xor (layer7_outputs(4694)));
    layer8_outputs(4053) <= (layer7_outputs(3531)) and not (layer7_outputs(1659));
    layer8_outputs(4054) <= (layer7_outputs(3611)) and (layer7_outputs(2858));
    layer8_outputs(4055) <= not(layer7_outputs(489));
    layer8_outputs(4056) <= not(layer7_outputs(595));
    layer8_outputs(4057) <= not(layer7_outputs(2914)) or (layer7_outputs(1330));
    layer8_outputs(4058) <= not(layer7_outputs(176));
    layer8_outputs(4059) <= not(layer7_outputs(802));
    layer8_outputs(4060) <= not(layer7_outputs(4413)) or (layer7_outputs(1881));
    layer8_outputs(4061) <= not((layer7_outputs(2595)) xor (layer7_outputs(3775)));
    layer8_outputs(4062) <= not(layer7_outputs(2909));
    layer8_outputs(4063) <= not(layer7_outputs(4525));
    layer8_outputs(4064) <= layer7_outputs(2213);
    layer8_outputs(4065) <= not((layer7_outputs(879)) xor (layer7_outputs(655)));
    layer8_outputs(4066) <= not(layer7_outputs(3756));
    layer8_outputs(4067) <= not((layer7_outputs(543)) and (layer7_outputs(2107)));
    layer8_outputs(4068) <= not((layer7_outputs(4950)) xor (layer7_outputs(960)));
    layer8_outputs(4069) <= layer7_outputs(341);
    layer8_outputs(4070) <= layer7_outputs(1295);
    layer8_outputs(4071) <= layer7_outputs(2327);
    layer8_outputs(4072) <= (layer7_outputs(912)) xor (layer7_outputs(2962));
    layer8_outputs(4073) <= not((layer7_outputs(3990)) and (layer7_outputs(35)));
    layer8_outputs(4074) <= not((layer7_outputs(806)) and (layer7_outputs(4215)));
    layer8_outputs(4075) <= not(layer7_outputs(931)) or (layer7_outputs(1385));
    layer8_outputs(4076) <= not((layer7_outputs(4317)) xor (layer7_outputs(2181)));
    layer8_outputs(4077) <= layer7_outputs(617);
    layer8_outputs(4078) <= not(layer7_outputs(1709));
    layer8_outputs(4079) <= layer7_outputs(1228);
    layer8_outputs(4080) <= not((layer7_outputs(2223)) and (layer7_outputs(4058)));
    layer8_outputs(4081) <= not(layer7_outputs(3887));
    layer8_outputs(4082) <= not(layer7_outputs(774));
    layer8_outputs(4083) <= layer7_outputs(3754);
    layer8_outputs(4084) <= not((layer7_outputs(1890)) xor (layer7_outputs(3333)));
    layer8_outputs(4085) <= not((layer7_outputs(4817)) and (layer7_outputs(1905)));
    layer8_outputs(4086) <= not(layer7_outputs(3718));
    layer8_outputs(4087) <= not(layer7_outputs(4328)) or (layer7_outputs(638));
    layer8_outputs(4088) <= layer7_outputs(1098);
    layer8_outputs(4089) <= layer7_outputs(4662);
    layer8_outputs(4090) <= not((layer7_outputs(2119)) xor (layer7_outputs(1354)));
    layer8_outputs(4091) <= not(layer7_outputs(2993));
    layer8_outputs(4092) <= not(layer7_outputs(1442));
    layer8_outputs(4093) <= layer7_outputs(2668);
    layer8_outputs(4094) <= layer7_outputs(2996);
    layer8_outputs(4095) <= (layer7_outputs(4490)) xor (layer7_outputs(770));
    layer8_outputs(4096) <= not(layer7_outputs(918));
    layer8_outputs(4097) <= not(layer7_outputs(1270));
    layer8_outputs(4098) <= layer7_outputs(3038);
    layer8_outputs(4099) <= layer7_outputs(1217);
    layer8_outputs(4100) <= layer7_outputs(2402);
    layer8_outputs(4101) <= not((layer7_outputs(2238)) xor (layer7_outputs(1626)));
    layer8_outputs(4102) <= not((layer7_outputs(4720)) xor (layer7_outputs(496)));
    layer8_outputs(4103) <= not(layer7_outputs(1617));
    layer8_outputs(4104) <= not((layer7_outputs(3675)) xor (layer7_outputs(3870)));
    layer8_outputs(4105) <= not((layer7_outputs(2027)) or (layer7_outputs(2072)));
    layer8_outputs(4106) <= layer7_outputs(2126);
    layer8_outputs(4107) <= not(layer7_outputs(850));
    layer8_outputs(4108) <= not(layer7_outputs(1642));
    layer8_outputs(4109) <= not(layer7_outputs(3307));
    layer8_outputs(4110) <= not(layer7_outputs(4446));
    layer8_outputs(4111) <= (layer7_outputs(2681)) and not (layer7_outputs(3315));
    layer8_outputs(4112) <= (layer7_outputs(3643)) and not (layer7_outputs(136));
    layer8_outputs(4113) <= not(layer7_outputs(2863));
    layer8_outputs(4114) <= not((layer7_outputs(138)) xor (layer7_outputs(2779)));
    layer8_outputs(4115) <= (layer7_outputs(1473)) xor (layer7_outputs(5114));
    layer8_outputs(4116) <= not((layer7_outputs(2349)) xor (layer7_outputs(476)));
    layer8_outputs(4117) <= (layer7_outputs(4357)) and not (layer7_outputs(4034));
    layer8_outputs(4118) <= not(layer7_outputs(2200));
    layer8_outputs(4119) <= layer7_outputs(4352);
    layer8_outputs(4120) <= not(layer7_outputs(328));
    layer8_outputs(4121) <= layer7_outputs(4225);
    layer8_outputs(4122) <= layer7_outputs(3897);
    layer8_outputs(4123) <= '0';
    layer8_outputs(4124) <= not(layer7_outputs(815));
    layer8_outputs(4125) <= (layer7_outputs(2703)) or (layer7_outputs(1796));
    layer8_outputs(4126) <= (layer7_outputs(4356)) and not (layer7_outputs(3985));
    layer8_outputs(4127) <= layer7_outputs(2515);
    layer8_outputs(4128) <= not(layer7_outputs(1752));
    layer8_outputs(4129) <= layer7_outputs(3949);
    layer8_outputs(4130) <= not(layer7_outputs(4576));
    layer8_outputs(4131) <= not(layer7_outputs(1433)) or (layer7_outputs(1073));
    layer8_outputs(4132) <= layer7_outputs(869);
    layer8_outputs(4133) <= (layer7_outputs(1571)) or (layer7_outputs(4685));
    layer8_outputs(4134) <= (layer7_outputs(625)) xor (layer7_outputs(3438));
    layer8_outputs(4135) <= not(layer7_outputs(3280)) or (layer7_outputs(3175));
    layer8_outputs(4136) <= layer7_outputs(1906);
    layer8_outputs(4137) <= not(layer7_outputs(4321));
    layer8_outputs(4138) <= layer7_outputs(5080);
    layer8_outputs(4139) <= not(layer7_outputs(1414));
    layer8_outputs(4140) <= (layer7_outputs(1023)) and (layer7_outputs(2241));
    layer8_outputs(4141) <= not((layer7_outputs(3005)) or (layer7_outputs(1481)));
    layer8_outputs(4142) <= layer7_outputs(4072);
    layer8_outputs(4143) <= not(layer7_outputs(140));
    layer8_outputs(4144) <= not(layer7_outputs(4286));
    layer8_outputs(4145) <= not((layer7_outputs(2182)) xor (layer7_outputs(2254)));
    layer8_outputs(4146) <= not(layer7_outputs(499)) or (layer7_outputs(857));
    layer8_outputs(4147) <= layer7_outputs(4588);
    layer8_outputs(4148) <= not(layer7_outputs(4286)) or (layer7_outputs(798));
    layer8_outputs(4149) <= layer7_outputs(2414);
    layer8_outputs(4150) <= not(layer7_outputs(247));
    layer8_outputs(4151) <= layer7_outputs(2241);
    layer8_outputs(4152) <= not((layer7_outputs(1359)) xor (layer7_outputs(440)));
    layer8_outputs(4153) <= not(layer7_outputs(3760));
    layer8_outputs(4154) <= layer7_outputs(2806);
    layer8_outputs(4155) <= (layer7_outputs(4012)) and (layer7_outputs(1611));
    layer8_outputs(4156) <= not((layer7_outputs(4462)) xor (layer7_outputs(1442)));
    layer8_outputs(4157) <= layer7_outputs(3154);
    layer8_outputs(4158) <= (layer7_outputs(3089)) and (layer7_outputs(2978));
    layer8_outputs(4159) <= not(layer7_outputs(1992));
    layer8_outputs(4160) <= not((layer7_outputs(63)) xor (layer7_outputs(2712)));
    layer8_outputs(4161) <= not((layer7_outputs(3379)) xor (layer7_outputs(2380)));
    layer8_outputs(4162) <= '0';
    layer8_outputs(4163) <= layer7_outputs(1355);
    layer8_outputs(4164) <= not(layer7_outputs(2761)) or (layer7_outputs(4587));
    layer8_outputs(4165) <= not(layer7_outputs(2176));
    layer8_outputs(4166) <= not(layer7_outputs(4524));
    layer8_outputs(4167) <= not(layer7_outputs(4141));
    layer8_outputs(4168) <= layer7_outputs(162);
    layer8_outputs(4169) <= not((layer7_outputs(1345)) and (layer7_outputs(2791)));
    layer8_outputs(4170) <= layer7_outputs(1061);
    layer8_outputs(4171) <= layer7_outputs(3068);
    layer8_outputs(4172) <= '1';
    layer8_outputs(4173) <= not((layer7_outputs(3964)) and (layer7_outputs(695)));
    layer8_outputs(4174) <= (layer7_outputs(3281)) and (layer7_outputs(4112));
    layer8_outputs(4175) <= not(layer7_outputs(3969)) or (layer7_outputs(3031));
    layer8_outputs(4176) <= not((layer7_outputs(4703)) xor (layer7_outputs(4330)));
    layer8_outputs(4177) <= not((layer7_outputs(3796)) and (layer7_outputs(3083)));
    layer8_outputs(4178) <= not(layer7_outputs(3207));
    layer8_outputs(4179) <= (layer7_outputs(758)) and not (layer7_outputs(1443));
    layer8_outputs(4180) <= layer7_outputs(151);
    layer8_outputs(4181) <= not(layer7_outputs(4725));
    layer8_outputs(4182) <= not(layer7_outputs(5041));
    layer8_outputs(4183) <= not(layer7_outputs(166));
    layer8_outputs(4184) <= not(layer7_outputs(2694));
    layer8_outputs(4185) <= not(layer7_outputs(4878)) or (layer7_outputs(4364));
    layer8_outputs(4186) <= layer7_outputs(901);
    layer8_outputs(4187) <= not(layer7_outputs(976));
    layer8_outputs(4188) <= not(layer7_outputs(5051));
    layer8_outputs(4189) <= not((layer7_outputs(1808)) xor (layer7_outputs(820)));
    layer8_outputs(4190) <= layer7_outputs(1957);
    layer8_outputs(4191) <= not((layer7_outputs(343)) or (layer7_outputs(118)));
    layer8_outputs(4192) <= (layer7_outputs(3001)) and (layer7_outputs(2863));
    layer8_outputs(4193) <= (layer7_outputs(2347)) xor (layer7_outputs(4));
    layer8_outputs(4194) <= not(layer7_outputs(803)) or (layer7_outputs(1727));
    layer8_outputs(4195) <= not(layer7_outputs(813));
    layer8_outputs(4196) <= not(layer7_outputs(4386)) or (layer7_outputs(3357));
    layer8_outputs(4197) <= (layer7_outputs(2169)) and not (layer7_outputs(1743));
    layer8_outputs(4198) <= not((layer7_outputs(4192)) xor (layer7_outputs(783)));
    layer8_outputs(4199) <= not((layer7_outputs(4418)) and (layer7_outputs(2964)));
    layer8_outputs(4200) <= layer7_outputs(1753);
    layer8_outputs(4201) <= (layer7_outputs(3321)) xor (layer7_outputs(4675));
    layer8_outputs(4202) <= (layer7_outputs(1998)) and (layer7_outputs(3569));
    layer8_outputs(4203) <= (layer7_outputs(2432)) and not (layer7_outputs(4730));
    layer8_outputs(4204) <= (layer7_outputs(2255)) and not (layer7_outputs(1001));
    layer8_outputs(4205) <= layer7_outputs(2195);
    layer8_outputs(4206) <= (layer7_outputs(1704)) and not (layer7_outputs(4133));
    layer8_outputs(4207) <= '1';
    layer8_outputs(4208) <= not((layer7_outputs(4994)) or (layer7_outputs(2705)));
    layer8_outputs(4209) <= not(layer7_outputs(4578));
    layer8_outputs(4210) <= not(layer7_outputs(1513));
    layer8_outputs(4211) <= (layer7_outputs(2301)) xor (layer7_outputs(5059));
    layer8_outputs(4212) <= not((layer7_outputs(3998)) xor (layer7_outputs(4979)));
    layer8_outputs(4213) <= layer7_outputs(4823);
    layer8_outputs(4214) <= not(layer7_outputs(3455));
    layer8_outputs(4215) <= layer7_outputs(148);
    layer8_outputs(4216) <= not((layer7_outputs(1869)) xor (layer7_outputs(621)));
    layer8_outputs(4217) <= not(layer7_outputs(1596));
    layer8_outputs(4218) <= (layer7_outputs(2689)) xor (layer7_outputs(3604));
    layer8_outputs(4219) <= (layer7_outputs(1758)) and not (layer7_outputs(1005));
    layer8_outputs(4220) <= (layer7_outputs(3344)) xor (layer7_outputs(3986));
    layer8_outputs(4221) <= not(layer7_outputs(243));
    layer8_outputs(4222) <= not((layer7_outputs(3804)) xor (layer7_outputs(3930)));
    layer8_outputs(4223) <= not(layer7_outputs(4806));
    layer8_outputs(4224) <= not((layer7_outputs(661)) xor (layer7_outputs(1128)));
    layer8_outputs(4225) <= (layer7_outputs(1265)) xor (layer7_outputs(2270));
    layer8_outputs(4226) <= layer7_outputs(345);
    layer8_outputs(4227) <= not(layer7_outputs(522));
    layer8_outputs(4228) <= not((layer7_outputs(874)) xor (layer7_outputs(1787)));
    layer8_outputs(4229) <= not((layer7_outputs(4149)) xor (layer7_outputs(5077)));
    layer8_outputs(4230) <= not(layer7_outputs(3365)) or (layer7_outputs(1384));
    layer8_outputs(4231) <= not(layer7_outputs(891));
    layer8_outputs(4232) <= not((layer7_outputs(4360)) xor (layer7_outputs(4336)));
    layer8_outputs(4233) <= not(layer7_outputs(3787));
    layer8_outputs(4234) <= not(layer7_outputs(2159));
    layer8_outputs(4235) <= (layer7_outputs(4410)) or (layer7_outputs(3218));
    layer8_outputs(4236) <= (layer7_outputs(3007)) and not (layer7_outputs(2652));
    layer8_outputs(4237) <= not((layer7_outputs(2553)) or (layer7_outputs(1754)));
    layer8_outputs(4238) <= layer7_outputs(565);
    layer8_outputs(4239) <= (layer7_outputs(2426)) and (layer7_outputs(2178));
    layer8_outputs(4240) <= not(layer7_outputs(532));
    layer8_outputs(4241) <= layer7_outputs(1314);
    layer8_outputs(4242) <= not((layer7_outputs(790)) xor (layer7_outputs(1387)));
    layer8_outputs(4243) <= layer7_outputs(4690);
    layer8_outputs(4244) <= not(layer7_outputs(5044));
    layer8_outputs(4245) <= not((layer7_outputs(2517)) and (layer7_outputs(1601)));
    layer8_outputs(4246) <= layer7_outputs(1272);
    layer8_outputs(4247) <= not(layer7_outputs(2902));
    layer8_outputs(4248) <= (layer7_outputs(4892)) and not (layer7_outputs(4787));
    layer8_outputs(4249) <= not(layer7_outputs(4401));
    layer8_outputs(4250) <= not((layer7_outputs(305)) xor (layer7_outputs(3651)));
    layer8_outputs(4251) <= not(layer7_outputs(2147)) or (layer7_outputs(4499));
    layer8_outputs(4252) <= not((layer7_outputs(839)) and (layer7_outputs(2986)));
    layer8_outputs(4253) <= not((layer7_outputs(260)) xor (layer7_outputs(1337)));
    layer8_outputs(4254) <= not((layer7_outputs(4262)) xor (layer7_outputs(454)));
    layer8_outputs(4255) <= not(layer7_outputs(3228));
    layer8_outputs(4256) <= not(layer7_outputs(111));
    layer8_outputs(4257) <= not((layer7_outputs(3798)) xor (layer7_outputs(2795)));
    layer8_outputs(4258) <= (layer7_outputs(499)) xor (layer7_outputs(359));
    layer8_outputs(4259) <= (layer7_outputs(1338)) and not (layer7_outputs(4800));
    layer8_outputs(4260) <= not((layer7_outputs(2811)) xor (layer7_outputs(1065)));
    layer8_outputs(4261) <= not(layer7_outputs(583));
    layer8_outputs(4262) <= (layer7_outputs(4674)) or (layer7_outputs(3107));
    layer8_outputs(4263) <= not(layer7_outputs(4862)) or (layer7_outputs(3553));
    layer8_outputs(4264) <= not(layer7_outputs(3864));
    layer8_outputs(4265) <= layer7_outputs(9);
    layer8_outputs(4266) <= not(layer7_outputs(3941));
    layer8_outputs(4267) <= not(layer7_outputs(4506));
    layer8_outputs(4268) <= (layer7_outputs(4917)) and (layer7_outputs(2548));
    layer8_outputs(4269) <= layer7_outputs(578);
    layer8_outputs(4270) <= (layer7_outputs(1242)) xor (layer7_outputs(3999));
    layer8_outputs(4271) <= (layer7_outputs(672)) xor (layer7_outputs(3642));
    layer8_outputs(4272) <= not(layer7_outputs(4118));
    layer8_outputs(4273) <= not(layer7_outputs(551));
    layer8_outputs(4274) <= layer7_outputs(4026);
    layer8_outputs(4275) <= not(layer7_outputs(2259));
    layer8_outputs(4276) <= layer7_outputs(4810);
    layer8_outputs(4277) <= layer7_outputs(4535);
    layer8_outputs(4278) <= not((layer7_outputs(1173)) xor (layer7_outputs(177)));
    layer8_outputs(4279) <= (layer7_outputs(5062)) xor (layer7_outputs(940));
    layer8_outputs(4280) <= layer7_outputs(360);
    layer8_outputs(4281) <= not((layer7_outputs(646)) xor (layer7_outputs(887)));
    layer8_outputs(4282) <= not(layer7_outputs(4498));
    layer8_outputs(4283) <= not(layer7_outputs(4767));
    layer8_outputs(4284) <= not((layer7_outputs(3854)) or (layer7_outputs(3850)));
    layer8_outputs(4285) <= '1';
    layer8_outputs(4286) <= (layer7_outputs(3564)) and not (layer7_outputs(4001));
    layer8_outputs(4287) <= not(layer7_outputs(3120)) or (layer7_outputs(629));
    layer8_outputs(4288) <= layer7_outputs(3635);
    layer8_outputs(4289) <= layer7_outputs(2560);
    layer8_outputs(4290) <= not(layer7_outputs(4378)) or (layer7_outputs(2074));
    layer8_outputs(4291) <= not(layer7_outputs(793));
    layer8_outputs(4292) <= (layer7_outputs(1483)) and not (layer7_outputs(3829));
    layer8_outputs(4293) <= not(layer7_outputs(4674));
    layer8_outputs(4294) <= (layer7_outputs(3740)) and not (layer7_outputs(2436));
    layer8_outputs(4295) <= layer7_outputs(275);
    layer8_outputs(4296) <= (layer7_outputs(1687)) xor (layer7_outputs(4107));
    layer8_outputs(4297) <= layer7_outputs(3757);
    layer8_outputs(4298) <= (layer7_outputs(1897)) and (layer7_outputs(2714));
    layer8_outputs(4299) <= layer7_outputs(4845);
    layer8_outputs(4300) <= layer7_outputs(1874);
    layer8_outputs(4301) <= layer7_outputs(3809);
    layer8_outputs(4302) <= (layer7_outputs(705)) xor (layer7_outputs(1271));
    layer8_outputs(4303) <= not(layer7_outputs(1370));
    layer8_outputs(4304) <= not((layer7_outputs(3542)) and (layer7_outputs(528)));
    layer8_outputs(4305) <= not((layer7_outputs(1404)) or (layer7_outputs(4463)));
    layer8_outputs(4306) <= not(layer7_outputs(1055)) or (layer7_outputs(759));
    layer8_outputs(4307) <= layer7_outputs(2498);
    layer8_outputs(4308) <= not(layer7_outputs(2872));
    layer8_outputs(4309) <= not(layer7_outputs(2982));
    layer8_outputs(4310) <= not(layer7_outputs(3462)) or (layer7_outputs(1115));
    layer8_outputs(4311) <= (layer7_outputs(3363)) xor (layer7_outputs(2517));
    layer8_outputs(4312) <= not((layer7_outputs(2767)) xor (layer7_outputs(1377)));
    layer8_outputs(4313) <= not(layer7_outputs(3600));
    layer8_outputs(4314) <= not(layer7_outputs(3632));
    layer8_outputs(4315) <= not(layer7_outputs(3693));
    layer8_outputs(4316) <= layer7_outputs(4184);
    layer8_outputs(4317) <= not((layer7_outputs(3917)) xor (layer7_outputs(914)));
    layer8_outputs(4318) <= not(layer7_outputs(867));
    layer8_outputs(4319) <= not(layer7_outputs(3892));
    layer8_outputs(4320) <= (layer7_outputs(4068)) xor (layer7_outputs(913));
    layer8_outputs(4321) <= not(layer7_outputs(836)) or (layer7_outputs(2706));
    layer8_outputs(4322) <= not((layer7_outputs(4551)) xor (layer7_outputs(4511)));
    layer8_outputs(4323) <= layer7_outputs(2770);
    layer8_outputs(4324) <= (layer7_outputs(38)) xor (layer7_outputs(3187));
    layer8_outputs(4325) <= not(layer7_outputs(710));
    layer8_outputs(4326) <= not((layer7_outputs(1955)) and (layer7_outputs(3987)));
    layer8_outputs(4327) <= not(layer7_outputs(5008));
    layer8_outputs(4328) <= layer7_outputs(2992);
    layer8_outputs(4329) <= not(layer7_outputs(187)) or (layer7_outputs(1746));
    layer8_outputs(4330) <= (layer7_outputs(919)) xor (layer7_outputs(4831));
    layer8_outputs(4331) <= not(layer7_outputs(2969));
    layer8_outputs(4332) <= not(layer7_outputs(3166)) or (layer7_outputs(4189));
    layer8_outputs(4333) <= not(layer7_outputs(4320));
    layer8_outputs(4334) <= layer7_outputs(2238);
    layer8_outputs(4335) <= (layer7_outputs(3435)) xor (layer7_outputs(3168));
    layer8_outputs(4336) <= not((layer7_outputs(3326)) or (layer7_outputs(3929)));
    layer8_outputs(4337) <= not(layer7_outputs(2311));
    layer8_outputs(4338) <= layer7_outputs(4053);
    layer8_outputs(4339) <= layer7_outputs(4666);
    layer8_outputs(4340) <= not(layer7_outputs(212));
    layer8_outputs(4341) <= (layer7_outputs(789)) or (layer7_outputs(3514));
    layer8_outputs(4342) <= not((layer7_outputs(3968)) and (layer7_outputs(3714)));
    layer8_outputs(4343) <= not((layer7_outputs(4753)) xor (layer7_outputs(2299)));
    layer8_outputs(4344) <= '0';
    layer8_outputs(4345) <= layer7_outputs(3404);
    layer8_outputs(4346) <= layer7_outputs(3216);
    layer8_outputs(4347) <= not(layer7_outputs(233));
    layer8_outputs(4348) <= layer7_outputs(2581);
    layer8_outputs(4349) <= layer7_outputs(3619);
    layer8_outputs(4350) <= not((layer7_outputs(3727)) and (layer7_outputs(4143)));
    layer8_outputs(4351) <= layer7_outputs(3011);
    layer8_outputs(4352) <= layer7_outputs(3482);
    layer8_outputs(4353) <= not(layer7_outputs(3463));
    layer8_outputs(4354) <= not(layer7_outputs(4593));
    layer8_outputs(4355) <= not((layer7_outputs(4726)) or (layer7_outputs(3401)));
    layer8_outputs(4356) <= not(layer7_outputs(3014));
    layer8_outputs(4357) <= not((layer7_outputs(1751)) xor (layer7_outputs(1527)));
    layer8_outputs(4358) <= not((layer7_outputs(845)) xor (layer7_outputs(3521)));
    layer8_outputs(4359) <= not((layer7_outputs(11)) xor (layer7_outputs(1789)));
    layer8_outputs(4360) <= not(layer7_outputs(4564));
    layer8_outputs(4361) <= layer7_outputs(2429);
    layer8_outputs(4362) <= not(layer7_outputs(1702));
    layer8_outputs(4363) <= not(layer7_outputs(206));
    layer8_outputs(4364) <= layer7_outputs(1041);
    layer8_outputs(4365) <= not((layer7_outputs(2583)) or (layer7_outputs(2527)));
    layer8_outputs(4366) <= (layer7_outputs(2033)) and not (layer7_outputs(3318));
    layer8_outputs(4367) <= not(layer7_outputs(2890));
    layer8_outputs(4368) <= layer7_outputs(325);
    layer8_outputs(4369) <= not(layer7_outputs(3114));
    layer8_outputs(4370) <= not(layer7_outputs(4526));
    layer8_outputs(4371) <= not(layer7_outputs(2487));
    layer8_outputs(4372) <= not(layer7_outputs(2479));
    layer8_outputs(4373) <= (layer7_outputs(650)) and not (layer7_outputs(1480));
    layer8_outputs(4374) <= (layer7_outputs(1448)) or (layer7_outputs(1341));
    layer8_outputs(4375) <= not(layer7_outputs(154)) or (layer7_outputs(1493));
    layer8_outputs(4376) <= not((layer7_outputs(2182)) xor (layer7_outputs(674)));
    layer8_outputs(4377) <= not(layer7_outputs(1293));
    layer8_outputs(4378) <= not(layer7_outputs(4140)) or (layer7_outputs(388));
    layer8_outputs(4379) <= not((layer7_outputs(3899)) xor (layer7_outputs(147)));
    layer8_outputs(4380) <= layer7_outputs(3264);
    layer8_outputs(4381) <= layer7_outputs(2560);
    layer8_outputs(4382) <= (layer7_outputs(3743)) xor (layer7_outputs(675));
    layer8_outputs(4383) <= (layer7_outputs(5103)) or (layer7_outputs(3298));
    layer8_outputs(4384) <= (layer7_outputs(4508)) or (layer7_outputs(2256));
    layer8_outputs(4385) <= not((layer7_outputs(1088)) and (layer7_outputs(636)));
    layer8_outputs(4386) <= not(layer7_outputs(1279));
    layer8_outputs(4387) <= not((layer7_outputs(4609)) xor (layer7_outputs(2041)));
    layer8_outputs(4388) <= not(layer7_outputs(3249));
    layer8_outputs(4389) <= not((layer7_outputs(2866)) or (layer7_outputs(415)));
    layer8_outputs(4390) <= layer7_outputs(3946);
    layer8_outputs(4391) <= not(layer7_outputs(2038));
    layer8_outputs(4392) <= not((layer7_outputs(3856)) xor (layer7_outputs(605)));
    layer8_outputs(4393) <= layer7_outputs(3798);
    layer8_outputs(4394) <= (layer7_outputs(5076)) xor (layer7_outputs(1783));
    layer8_outputs(4395) <= layer7_outputs(1944);
    layer8_outputs(4396) <= '1';
    layer8_outputs(4397) <= layer7_outputs(3626);
    layer8_outputs(4398) <= (layer7_outputs(2309)) and (layer7_outputs(4279));
    layer8_outputs(4399) <= not(layer7_outputs(1779));
    layer8_outputs(4400) <= layer7_outputs(232);
    layer8_outputs(4401) <= layer7_outputs(5065);
    layer8_outputs(4402) <= not(layer7_outputs(2955));
    layer8_outputs(4403) <= (layer7_outputs(1865)) xor (layer7_outputs(3270));
    layer8_outputs(4404) <= not((layer7_outputs(3125)) or (layer7_outputs(2454)));
    layer8_outputs(4405) <= not(layer7_outputs(1722)) or (layer7_outputs(4359));
    layer8_outputs(4406) <= not(layer7_outputs(3449));
    layer8_outputs(4407) <= not(layer7_outputs(1004));
    layer8_outputs(4408) <= layer7_outputs(238);
    layer8_outputs(4409) <= not(layer7_outputs(5021)) or (layer7_outputs(10));
    layer8_outputs(4410) <= layer7_outputs(1915);
    layer8_outputs(4411) <= layer7_outputs(4397);
    layer8_outputs(4412) <= not((layer7_outputs(1962)) and (layer7_outputs(1138)));
    layer8_outputs(4413) <= not(layer7_outputs(325)) or (layer7_outputs(2199));
    layer8_outputs(4414) <= not(layer7_outputs(2663));
    layer8_outputs(4415) <= layer7_outputs(3793);
    layer8_outputs(4416) <= layer7_outputs(3717);
    layer8_outputs(4417) <= layer7_outputs(294);
    layer8_outputs(4418) <= not((layer7_outputs(80)) xor (layer7_outputs(4112)));
    layer8_outputs(4419) <= not(layer7_outputs(3595));
    layer8_outputs(4420) <= (layer7_outputs(396)) or (layer7_outputs(1645));
    layer8_outputs(4421) <= layer7_outputs(3883);
    layer8_outputs(4422) <= (layer7_outputs(3776)) and (layer7_outputs(3707));
    layer8_outputs(4423) <= not((layer7_outputs(3410)) or (layer7_outputs(3047)));
    layer8_outputs(4424) <= not(layer7_outputs(3377));
    layer8_outputs(4425) <= (layer7_outputs(3728)) and not (layer7_outputs(3685));
    layer8_outputs(4426) <= not(layer7_outputs(3981));
    layer8_outputs(4427) <= (layer7_outputs(955)) xor (layer7_outputs(4789));
    layer8_outputs(4428) <= not(layer7_outputs(1221));
    layer8_outputs(4429) <= layer7_outputs(4851);
    layer8_outputs(4430) <= not(layer7_outputs(1840));
    layer8_outputs(4431) <= not((layer7_outputs(2687)) xor (layer7_outputs(1643)));
    layer8_outputs(4432) <= not((layer7_outputs(567)) xor (layer7_outputs(4464)));
    layer8_outputs(4433) <= not(layer7_outputs(1861));
    layer8_outputs(4434) <= not(layer7_outputs(3818));
    layer8_outputs(4435) <= not(layer7_outputs(1899));
    layer8_outputs(4436) <= layer7_outputs(3162);
    layer8_outputs(4437) <= (layer7_outputs(527)) xor (layer7_outputs(3467));
    layer8_outputs(4438) <= not((layer7_outputs(3275)) or (layer7_outputs(3876)));
    layer8_outputs(4439) <= not((layer7_outputs(4221)) xor (layer7_outputs(3825)));
    layer8_outputs(4440) <= layer7_outputs(160);
    layer8_outputs(4441) <= not((layer7_outputs(3651)) xor (layer7_outputs(3364)));
    layer8_outputs(4442) <= (layer7_outputs(2665)) xor (layer7_outputs(129));
    layer8_outputs(4443) <= not((layer7_outputs(4167)) and (layer7_outputs(290)));
    layer8_outputs(4444) <= (layer7_outputs(2746)) xor (layer7_outputs(2292));
    layer8_outputs(4445) <= not(layer7_outputs(4363));
    layer8_outputs(4446) <= not((layer7_outputs(2607)) xor (layer7_outputs(3724)));
    layer8_outputs(4447) <= layer7_outputs(2760);
    layer8_outputs(4448) <= not(layer7_outputs(2711));
    layer8_outputs(4449) <= (layer7_outputs(2671)) xor (layer7_outputs(1296));
    layer8_outputs(4450) <= (layer7_outputs(722)) xor (layer7_outputs(421));
    layer8_outputs(4451) <= not(layer7_outputs(4566));
    layer8_outputs(4452) <= layer7_outputs(2282);
    layer8_outputs(4453) <= not((layer7_outputs(4567)) and (layer7_outputs(5119)));
    layer8_outputs(4454) <= not((layer7_outputs(5009)) and (layer7_outputs(4732)));
    layer8_outputs(4455) <= not(layer7_outputs(613)) or (layer7_outputs(4573));
    layer8_outputs(4456) <= (layer7_outputs(1856)) xor (layer7_outputs(3810));
    layer8_outputs(4457) <= not(layer7_outputs(3881)) or (layer7_outputs(3597));
    layer8_outputs(4458) <= layer7_outputs(4781);
    layer8_outputs(4459) <= not((layer7_outputs(1910)) xor (layer7_outputs(3519)));
    layer8_outputs(4460) <= not((layer7_outputs(3446)) xor (layer7_outputs(1925)));
    layer8_outputs(4461) <= not(layer7_outputs(1395));
    layer8_outputs(4462) <= not((layer7_outputs(3529)) xor (layer7_outputs(4631)));
    layer8_outputs(4463) <= layer7_outputs(3602);
    layer8_outputs(4464) <= layer7_outputs(3013);
    layer8_outputs(4465) <= not(layer7_outputs(329));
    layer8_outputs(4466) <= not(layer7_outputs(3795));
    layer8_outputs(4467) <= not(layer7_outputs(1718));
    layer8_outputs(4468) <= not(layer7_outputs(742));
    layer8_outputs(4469) <= (layer7_outputs(4962)) and not (layer7_outputs(2599));
    layer8_outputs(4470) <= layer7_outputs(2759);
    layer8_outputs(4471) <= (layer7_outputs(2286)) xor (layer7_outputs(3813));
    layer8_outputs(4472) <= (layer7_outputs(688)) xor (layer7_outputs(3109));
    layer8_outputs(4473) <= not(layer7_outputs(2623));
    layer8_outputs(4474) <= not(layer7_outputs(1180));
    layer8_outputs(4475) <= not((layer7_outputs(4313)) or (layer7_outputs(2563)));
    layer8_outputs(4476) <= layer7_outputs(5022);
    layer8_outputs(4477) <= (layer7_outputs(4140)) xor (layer7_outputs(840));
    layer8_outputs(4478) <= layer7_outputs(4329);
    layer8_outputs(4479) <= '0';
    layer8_outputs(4480) <= not((layer7_outputs(5035)) xor (layer7_outputs(3735)));
    layer8_outputs(4481) <= (layer7_outputs(259)) and (layer7_outputs(2153));
    layer8_outputs(4482) <= layer7_outputs(3512);
    layer8_outputs(4483) <= '1';
    layer8_outputs(4484) <= layer7_outputs(1226);
    layer8_outputs(4485) <= '1';
    layer8_outputs(4486) <= not(layer7_outputs(4888)) or (layer7_outputs(4719));
    layer8_outputs(4487) <= not(layer7_outputs(3975));
    layer8_outputs(4488) <= not((layer7_outputs(2891)) or (layer7_outputs(3123)));
    layer8_outputs(4489) <= (layer7_outputs(2151)) xor (layer7_outputs(3269));
    layer8_outputs(4490) <= not(layer7_outputs(3095));
    layer8_outputs(4491) <= (layer7_outputs(4526)) and not (layer7_outputs(2373));
    layer8_outputs(4492) <= layer7_outputs(693);
    layer8_outputs(4493) <= not((layer7_outputs(4707)) xor (layer7_outputs(4942)));
    layer8_outputs(4494) <= layer7_outputs(2975);
    layer8_outputs(4495) <= not(layer7_outputs(333));
    layer8_outputs(4496) <= (layer7_outputs(1740)) and not (layer7_outputs(2574));
    layer8_outputs(4497) <= (layer7_outputs(1280)) xor (layer7_outputs(3466));
    layer8_outputs(4498) <= not(layer7_outputs(1047));
    layer8_outputs(4499) <= (layer7_outputs(2586)) and not (layer7_outputs(3780));
    layer8_outputs(4500) <= layer7_outputs(4195);
    layer8_outputs(4501) <= not(layer7_outputs(3368));
    layer8_outputs(4502) <= layer7_outputs(3681);
    layer8_outputs(4503) <= not(layer7_outputs(3483));
    layer8_outputs(4504) <= layer7_outputs(291);
    layer8_outputs(4505) <= (layer7_outputs(548)) xor (layer7_outputs(1834));
    layer8_outputs(4506) <= (layer7_outputs(1507)) and not (layer7_outputs(1514));
    layer8_outputs(4507) <= (layer7_outputs(1868)) xor (layer7_outputs(4128));
    layer8_outputs(4508) <= layer7_outputs(2195);
    layer8_outputs(4509) <= not((layer7_outputs(1600)) xor (layer7_outputs(4003)));
    layer8_outputs(4510) <= not(layer7_outputs(2972)) or (layer7_outputs(1026));
    layer8_outputs(4511) <= not(layer7_outputs(1806));
    layer8_outputs(4512) <= not(layer7_outputs(3962));
    layer8_outputs(4513) <= (layer7_outputs(4645)) xor (layer7_outputs(1506));
    layer8_outputs(4514) <= not(layer7_outputs(1529));
    layer8_outputs(4515) <= not(layer7_outputs(838));
    layer8_outputs(4516) <= not(layer7_outputs(1469));
    layer8_outputs(4517) <= layer7_outputs(157);
    layer8_outputs(4518) <= (layer7_outputs(1276)) and not (layer7_outputs(2403));
    layer8_outputs(4519) <= not(layer7_outputs(5083));
    layer8_outputs(4520) <= (layer7_outputs(4534)) xor (layer7_outputs(2409));
    layer8_outputs(4521) <= layer7_outputs(236);
    layer8_outputs(4522) <= not((layer7_outputs(3663)) or (layer7_outputs(1976)));
    layer8_outputs(4523) <= (layer7_outputs(4648)) xor (layer7_outputs(3255));
    layer8_outputs(4524) <= not(layer7_outputs(426));
    layer8_outputs(4525) <= not(layer7_outputs(1383));
    layer8_outputs(4526) <= (layer7_outputs(4705)) or (layer7_outputs(2994));
    layer8_outputs(4527) <= not(layer7_outputs(4082)) or (layer7_outputs(3434));
    layer8_outputs(4528) <= layer7_outputs(105);
    layer8_outputs(4529) <= (layer7_outputs(495)) and not (layer7_outputs(5021));
    layer8_outputs(4530) <= layer7_outputs(4830);
    layer8_outputs(4531) <= layer7_outputs(1684);
    layer8_outputs(4532) <= layer7_outputs(2414);
    layer8_outputs(4533) <= (layer7_outputs(5048)) xor (layer7_outputs(2542));
    layer8_outputs(4534) <= layer7_outputs(2538);
    layer8_outputs(4535) <= layer7_outputs(1170);
    layer8_outputs(4536) <= not(layer7_outputs(620));
    layer8_outputs(4537) <= layer7_outputs(4656);
    layer8_outputs(4538) <= '1';
    layer8_outputs(4539) <= not((layer7_outputs(4661)) xor (layer7_outputs(3235)));
    layer8_outputs(4540) <= not((layer7_outputs(1591)) xor (layer7_outputs(1638)));
    layer8_outputs(4541) <= not(layer7_outputs(2589));
    layer8_outputs(4542) <= (layer7_outputs(740)) and not (layer7_outputs(2329));
    layer8_outputs(4543) <= (layer7_outputs(1878)) or (layer7_outputs(2805));
    layer8_outputs(4544) <= (layer7_outputs(2173)) xor (layer7_outputs(745));
    layer8_outputs(4545) <= (layer7_outputs(282)) and not (layer7_outputs(4644));
    layer8_outputs(4546) <= not(layer7_outputs(5073));
    layer8_outputs(4547) <= not((layer7_outputs(4074)) or (layer7_outputs(108)));
    layer8_outputs(4548) <= (layer7_outputs(4491)) and not (layer7_outputs(1894));
    layer8_outputs(4549) <= not((layer7_outputs(3657)) xor (layer7_outputs(3272)));
    layer8_outputs(4550) <= not(layer7_outputs(1467)) or (layer7_outputs(2733));
    layer8_outputs(4551) <= not(layer7_outputs(2944)) or (layer7_outputs(3802));
    layer8_outputs(4552) <= not((layer7_outputs(1506)) xor (layer7_outputs(4407)));
    layer8_outputs(4553) <= not(layer7_outputs(3146)) or (layer7_outputs(1175));
    layer8_outputs(4554) <= not(layer7_outputs(595));
    layer8_outputs(4555) <= not(layer7_outputs(1918));
    layer8_outputs(4556) <= not(layer7_outputs(3278));
    layer8_outputs(4557) <= layer7_outputs(4854);
    layer8_outputs(4558) <= (layer7_outputs(4664)) or (layer7_outputs(4663));
    layer8_outputs(4559) <= (layer7_outputs(712)) or (layer7_outputs(3229));
    layer8_outputs(4560) <= not((layer7_outputs(4014)) xor (layer7_outputs(5065)));
    layer8_outputs(4561) <= layer7_outputs(3833);
    layer8_outputs(4562) <= not(layer7_outputs(3395));
    layer8_outputs(4563) <= not(layer7_outputs(1819));
    layer8_outputs(4564) <= (layer7_outputs(5063)) xor (layer7_outputs(4086));
    layer8_outputs(4565) <= not(layer7_outputs(303));
    layer8_outputs(4566) <= (layer7_outputs(2303)) or (layer7_outputs(4742));
    layer8_outputs(4567) <= (layer7_outputs(1916)) and not (layer7_outputs(1721));
    layer8_outputs(4568) <= not((layer7_outputs(2351)) and (layer7_outputs(691)));
    layer8_outputs(4569) <= not(layer7_outputs(4256));
    layer8_outputs(4570) <= not(layer7_outputs(2832)) or (layer7_outputs(4186));
    layer8_outputs(4571) <= '1';
    layer8_outputs(4572) <= not((layer7_outputs(4905)) and (layer7_outputs(2197)));
    layer8_outputs(4573) <= not(layer7_outputs(5024));
    layer8_outputs(4574) <= not(layer7_outputs(3229)) or (layer7_outputs(899));
    layer8_outputs(4575) <= not((layer7_outputs(4612)) xor (layer7_outputs(1285)));
    layer8_outputs(4576) <= not(layer7_outputs(2120)) or (layer7_outputs(852));
    layer8_outputs(4577) <= (layer7_outputs(2896)) xor (layer7_outputs(4816));
    layer8_outputs(4578) <= not(layer7_outputs(1016)) or (layer7_outputs(83));
    layer8_outputs(4579) <= not(layer7_outputs(3242));
    layer8_outputs(4580) <= not((layer7_outputs(102)) or (layer7_outputs(2591)));
    layer8_outputs(4581) <= (layer7_outputs(2109)) and not (layer7_outputs(3744));
    layer8_outputs(4582) <= layer7_outputs(4047);
    layer8_outputs(4583) <= not(layer7_outputs(2921));
    layer8_outputs(4584) <= layer7_outputs(4431);
    layer8_outputs(4585) <= layer7_outputs(683);
    layer8_outputs(4586) <= (layer7_outputs(4569)) xor (layer7_outputs(3040));
    layer8_outputs(4587) <= layer7_outputs(1008);
    layer8_outputs(4588) <= not(layer7_outputs(4019)) or (layer7_outputs(1233));
    layer8_outputs(4589) <= '0';
    layer8_outputs(4590) <= not((layer7_outputs(3352)) and (layer7_outputs(2792)));
    layer8_outputs(4591) <= (layer7_outputs(610)) and (layer7_outputs(3442));
    layer8_outputs(4592) <= layer7_outputs(5038);
    layer8_outputs(4593) <= not(layer7_outputs(745));
    layer8_outputs(4594) <= layer7_outputs(4437);
    layer8_outputs(4595) <= not(layer7_outputs(1290));
    layer8_outputs(4596) <= (layer7_outputs(3769)) and not (layer7_outputs(209));
    layer8_outputs(4597) <= (layer7_outputs(3608)) xor (layer7_outputs(3220));
    layer8_outputs(4598) <= not((layer7_outputs(1628)) xor (layer7_outputs(3275)));
    layer8_outputs(4599) <= not(layer7_outputs(159));
    layer8_outputs(4600) <= (layer7_outputs(4312)) xor (layer7_outputs(3490));
    layer8_outputs(4601) <= not(layer7_outputs(4500));
    layer8_outputs(4602) <= not((layer7_outputs(1552)) xor (layer7_outputs(4997)));
    layer8_outputs(4603) <= (layer7_outputs(3394)) and (layer7_outputs(4938));
    layer8_outputs(4604) <= layer7_outputs(228);
    layer8_outputs(4605) <= layer7_outputs(249);
    layer8_outputs(4606) <= layer7_outputs(3916);
    layer8_outputs(4607) <= not(layer7_outputs(1766));
    layer8_outputs(4608) <= not((layer7_outputs(684)) or (layer7_outputs(4453)));
    layer8_outputs(4609) <= not(layer7_outputs(1421));
    layer8_outputs(4610) <= (layer7_outputs(4341)) xor (layer7_outputs(2654));
    layer8_outputs(4611) <= layer7_outputs(1605);
    layer8_outputs(4612) <= layer7_outputs(4273);
    layer8_outputs(4613) <= layer7_outputs(4097);
    layer8_outputs(4614) <= not((layer7_outputs(2361)) or (layer7_outputs(469)));
    layer8_outputs(4615) <= not(layer7_outputs(4532));
    layer8_outputs(4616) <= (layer7_outputs(4859)) xor (layer7_outputs(4105));
    layer8_outputs(4617) <= not((layer7_outputs(1097)) and (layer7_outputs(4754)));
    layer8_outputs(4618) <= (layer7_outputs(840)) xor (layer7_outputs(2463));
    layer8_outputs(4619) <= (layer7_outputs(4077)) xor (layer7_outputs(535));
    layer8_outputs(4620) <= (layer7_outputs(4281)) xor (layer7_outputs(692));
    layer8_outputs(4621) <= (layer7_outputs(4241)) xor (layer7_outputs(3051));
    layer8_outputs(4622) <= not(layer7_outputs(324));
    layer8_outputs(4623) <= not(layer7_outputs(4310));
    layer8_outputs(4624) <= (layer7_outputs(2389)) xor (layer7_outputs(3348));
    layer8_outputs(4625) <= layer7_outputs(1486);
    layer8_outputs(4626) <= (layer7_outputs(3217)) xor (layer7_outputs(3586));
    layer8_outputs(4627) <= layer7_outputs(2133);
    layer8_outputs(4628) <= layer7_outputs(1359);
    layer8_outputs(4629) <= (layer7_outputs(3538)) and not (layer7_outputs(1578));
    layer8_outputs(4630) <= layer7_outputs(2228);
    layer8_outputs(4631) <= not((layer7_outputs(4970)) xor (layer7_outputs(3809)));
    layer8_outputs(4632) <= layer7_outputs(2935);
    layer8_outputs(4633) <= not((layer7_outputs(1002)) and (layer7_outputs(1794)));
    layer8_outputs(4634) <= (layer7_outputs(2079)) xor (layer7_outputs(4654));
    layer8_outputs(4635) <= (layer7_outputs(4090)) xor (layer7_outputs(2628));
    layer8_outputs(4636) <= not((layer7_outputs(5028)) xor (layer7_outputs(266)));
    layer8_outputs(4637) <= not(layer7_outputs(3585));
    layer8_outputs(4638) <= not(layer7_outputs(4047));
    layer8_outputs(4639) <= layer7_outputs(1226);
    layer8_outputs(4640) <= not((layer7_outputs(4428)) xor (layer7_outputs(2776)));
    layer8_outputs(4641) <= not((layer7_outputs(167)) xor (layer7_outputs(4766)));
    layer8_outputs(4642) <= not(layer7_outputs(2051));
    layer8_outputs(4643) <= not((layer7_outputs(1167)) xor (layer7_outputs(7)));
    layer8_outputs(4644) <= not(layer7_outputs(2116));
    layer8_outputs(4645) <= not(layer7_outputs(713));
    layer8_outputs(4646) <= not(layer7_outputs(2437));
    layer8_outputs(4647) <= not((layer7_outputs(370)) xor (layer7_outputs(1307)));
    layer8_outputs(4648) <= (layer7_outputs(4311)) xor (layer7_outputs(639));
    layer8_outputs(4649) <= not(layer7_outputs(4299));
    layer8_outputs(4650) <= not((layer7_outputs(1143)) or (layer7_outputs(3170)));
    layer8_outputs(4651) <= layer7_outputs(4965);
    layer8_outputs(4652) <= not(layer7_outputs(1121));
    layer8_outputs(4653) <= (layer7_outputs(1162)) xor (layer7_outputs(3536));
    layer8_outputs(4654) <= not(layer7_outputs(4343));
    layer8_outputs(4655) <= (layer7_outputs(904)) xor (layer7_outputs(4847));
    layer8_outputs(4656) <= layer7_outputs(3094);
    layer8_outputs(4657) <= (layer7_outputs(533)) xor (layer7_outputs(1414));
    layer8_outputs(4658) <= (layer7_outputs(2133)) xor (layer7_outputs(2144));
    layer8_outputs(4659) <= layer7_outputs(5116);
    layer8_outputs(4660) <= not(layer7_outputs(2122)) or (layer7_outputs(4764));
    layer8_outputs(4661) <= not((layer7_outputs(1252)) xor (layer7_outputs(178)));
    layer8_outputs(4662) <= not(layer7_outputs(3852));
    layer8_outputs(4663) <= '1';
    layer8_outputs(4664) <= not(layer7_outputs(4344)) or (layer7_outputs(315));
    layer8_outputs(4665) <= layer7_outputs(1373);
    layer8_outputs(4666) <= (layer7_outputs(18)) or (layer7_outputs(1551));
    layer8_outputs(4667) <= not(layer7_outputs(2580));
    layer8_outputs(4668) <= not((layer7_outputs(923)) xor (layer7_outputs(1847)));
    layer8_outputs(4669) <= not((layer7_outputs(801)) xor (layer7_outputs(3488)));
    layer8_outputs(4670) <= layer7_outputs(564);
    layer8_outputs(4671) <= not((layer7_outputs(2481)) xor (layer7_outputs(1250)));
    layer8_outputs(4672) <= (layer7_outputs(2611)) and (layer7_outputs(120));
    layer8_outputs(4673) <= not(layer7_outputs(3227));
    layer8_outputs(4674) <= (layer7_outputs(380)) xor (layer7_outputs(372));
    layer8_outputs(4675) <= (layer7_outputs(1198)) and not (layer7_outputs(2003));
    layer8_outputs(4676) <= not(layer7_outputs(219));
    layer8_outputs(4677) <= layer7_outputs(1549);
    layer8_outputs(4678) <= not((layer7_outputs(2495)) xor (layer7_outputs(4898)));
    layer8_outputs(4679) <= layer7_outputs(4830);
    layer8_outputs(4680) <= not((layer7_outputs(2139)) and (layer7_outputs(4363)));
    layer8_outputs(4681) <= layer7_outputs(3120);
    layer8_outputs(4682) <= not((layer7_outputs(994)) and (layer7_outputs(3173)));
    layer8_outputs(4683) <= (layer7_outputs(4355)) and (layer7_outputs(937));
    layer8_outputs(4684) <= layer7_outputs(1091);
    layer8_outputs(4685) <= (layer7_outputs(4156)) or (layer7_outputs(4828));
    layer8_outputs(4686) <= layer7_outputs(352);
    layer8_outputs(4687) <= not((layer7_outputs(3180)) or (layer7_outputs(4603)));
    layer8_outputs(4688) <= layer7_outputs(3596);
    layer8_outputs(4689) <= layer7_outputs(1413);
    layer8_outputs(4690) <= layer7_outputs(3223);
    layer8_outputs(4691) <= not(layer7_outputs(2816));
    layer8_outputs(4692) <= (layer7_outputs(1523)) xor (layer7_outputs(2758));
    layer8_outputs(4693) <= layer7_outputs(2309);
    layer8_outputs(4694) <= (layer7_outputs(3257)) xor (layer7_outputs(434));
    layer8_outputs(4695) <= not(layer7_outputs(4794)) or (layer7_outputs(3977));
    layer8_outputs(4696) <= (layer7_outputs(4443)) xor (layer7_outputs(1014));
    layer8_outputs(4697) <= layer7_outputs(318);
    layer8_outputs(4698) <= (layer7_outputs(5049)) xor (layer7_outputs(2461));
    layer8_outputs(4699) <= not((layer7_outputs(660)) xor (layer7_outputs(3843)));
    layer8_outputs(4700) <= not((layer7_outputs(1781)) xor (layer7_outputs(3213)));
    layer8_outputs(4701) <= layer7_outputs(1900);
    layer8_outputs(4702) <= (layer7_outputs(920)) xor (layer7_outputs(223));
    layer8_outputs(4703) <= layer7_outputs(714);
    layer8_outputs(4704) <= (layer7_outputs(3872)) and (layer7_outputs(3070));
    layer8_outputs(4705) <= not(layer7_outputs(556));
    layer8_outputs(4706) <= layer7_outputs(5081);
    layer8_outputs(4707) <= (layer7_outputs(3852)) and not (layer7_outputs(518));
    layer8_outputs(4708) <= not((layer7_outputs(1388)) and (layer7_outputs(3348)));
    layer8_outputs(4709) <= layer7_outputs(4969);
    layer8_outputs(4710) <= not(layer7_outputs(851));
    layer8_outputs(4711) <= layer7_outputs(1328);
    layer8_outputs(4712) <= (layer7_outputs(2633)) and not (layer7_outputs(3495));
    layer8_outputs(4713) <= (layer7_outputs(4860)) xor (layer7_outputs(1913));
    layer8_outputs(4714) <= (layer7_outputs(381)) or (layer7_outputs(4925));
    layer8_outputs(4715) <= not(layer7_outputs(3702)) or (layer7_outputs(1148));
    layer8_outputs(4716) <= '1';
    layer8_outputs(4717) <= not(layer7_outputs(845));
    layer8_outputs(4718) <= not(layer7_outputs(2415));
    layer8_outputs(4719) <= (layer7_outputs(4563)) xor (layer7_outputs(2658));
    layer8_outputs(4720) <= not((layer7_outputs(930)) xor (layer7_outputs(354)));
    layer8_outputs(4721) <= (layer7_outputs(3988)) and (layer7_outputs(186));
    layer8_outputs(4722) <= (layer7_outputs(1328)) and (layer7_outputs(4974));
    layer8_outputs(4723) <= layer7_outputs(2703);
    layer8_outputs(4724) <= layer7_outputs(603);
    layer8_outputs(4725) <= not((layer7_outputs(2364)) xor (layer7_outputs(1229)));
    layer8_outputs(4726) <= not(layer7_outputs(1350));
    layer8_outputs(4727) <= not((layer7_outputs(3155)) xor (layer7_outputs(4487)));
    layer8_outputs(4728) <= not(layer7_outputs(2083)) or (layer7_outputs(29));
    layer8_outputs(4729) <= (layer7_outputs(4728)) or (layer7_outputs(1157));
    layer8_outputs(4730) <= not(layer7_outputs(3774));
    layer8_outputs(4731) <= (layer7_outputs(3391)) and (layer7_outputs(2824));
    layer8_outputs(4732) <= not(layer7_outputs(3283));
    layer8_outputs(4733) <= layer7_outputs(3839);
    layer8_outputs(4734) <= not((layer7_outputs(158)) xor (layer7_outputs(2600)));
    layer8_outputs(4735) <= not(layer7_outputs(4018));
    layer8_outputs(4736) <= not(layer7_outputs(3547));
    layer8_outputs(4737) <= not((layer7_outputs(4122)) and (layer7_outputs(2368)));
    layer8_outputs(4738) <= not((layer7_outputs(3427)) xor (layer7_outputs(4596)));
    layer8_outputs(4739) <= layer7_outputs(2471);
    layer8_outputs(4740) <= layer7_outputs(3382);
    layer8_outputs(4741) <= layer7_outputs(1777);
    layer8_outputs(4742) <= not(layer7_outputs(1418));
    layer8_outputs(4743) <= (layer7_outputs(509)) xor (layer7_outputs(3121));
    layer8_outputs(4744) <= layer7_outputs(2441);
    layer8_outputs(4745) <= not(layer7_outputs(4802)) or (layer7_outputs(1174));
    layer8_outputs(4746) <= not(layer7_outputs(2084));
    layer8_outputs(4747) <= not(layer7_outputs(0)) or (layer7_outputs(5117));
    layer8_outputs(4748) <= layer7_outputs(3114);
    layer8_outputs(4749) <= not(layer7_outputs(4475));
    layer8_outputs(4750) <= not(layer7_outputs(3705));
    layer8_outputs(4751) <= not(layer7_outputs(4452));
    layer8_outputs(4752) <= not(layer7_outputs(3802));
    layer8_outputs(4753) <= layer7_outputs(3480);
    layer8_outputs(4754) <= not(layer7_outputs(4136)) or (layer7_outputs(146));
    layer8_outputs(4755) <= '0';
    layer8_outputs(4756) <= not(layer7_outputs(1622));
    layer8_outputs(4757) <= not((layer7_outputs(3892)) and (layer7_outputs(2839)));
    layer8_outputs(4758) <= layer7_outputs(42);
    layer8_outputs(4759) <= layer7_outputs(1586);
    layer8_outputs(4760) <= (layer7_outputs(4915)) and not (layer7_outputs(4680));
    layer8_outputs(4761) <= layer7_outputs(1006);
    layer8_outputs(4762) <= (layer7_outputs(4120)) xor (layer7_outputs(1719));
    layer8_outputs(4763) <= layer7_outputs(1227);
    layer8_outputs(4764) <= not(layer7_outputs(1810));
    layer8_outputs(4765) <= '1';
    layer8_outputs(4766) <= not(layer7_outputs(2383));
    layer8_outputs(4767) <= not((layer7_outputs(1137)) xor (layer7_outputs(1841)));
    layer8_outputs(4768) <= layer7_outputs(3939);
    layer8_outputs(4769) <= not(layer7_outputs(2058)) or (layer7_outputs(3191));
    layer8_outputs(4770) <= (layer7_outputs(5042)) and (layer7_outputs(264));
    layer8_outputs(4771) <= not((layer7_outputs(1757)) xor (layer7_outputs(4957)));
    layer8_outputs(4772) <= not(layer7_outputs(2013));
    layer8_outputs(4773) <= (layer7_outputs(3222)) xor (layer7_outputs(588));
    layer8_outputs(4774) <= layer7_outputs(4035);
    layer8_outputs(4775) <= layer7_outputs(1504);
    layer8_outputs(4776) <= layer7_outputs(798);
    layer8_outputs(4777) <= not(layer7_outputs(2769)) or (layer7_outputs(898));
    layer8_outputs(4778) <= layer7_outputs(3890);
    layer8_outputs(4779) <= not((layer7_outputs(2173)) and (layer7_outputs(1457)));
    layer8_outputs(4780) <= not(layer7_outputs(1417));
    layer8_outputs(4781) <= not(layer7_outputs(631));
    layer8_outputs(4782) <= (layer7_outputs(4009)) and not (layer7_outputs(2545));
    layer8_outputs(4783) <= layer7_outputs(4139);
    layer8_outputs(4784) <= layer7_outputs(1505);
    layer8_outputs(4785) <= not(layer7_outputs(2750));
    layer8_outputs(4786) <= layer7_outputs(4397);
    layer8_outputs(4787) <= not((layer7_outputs(1711)) or (layer7_outputs(2860)));
    layer8_outputs(4788) <= layer7_outputs(3574);
    layer8_outputs(4789) <= (layer7_outputs(396)) xor (layer7_outputs(2215));
    layer8_outputs(4790) <= (layer7_outputs(3012)) and not (layer7_outputs(2369));
    layer8_outputs(4791) <= not(layer7_outputs(3869));
    layer8_outputs(4792) <= not((layer7_outputs(4602)) xor (layer7_outputs(2243)));
    layer8_outputs(4793) <= not(layer7_outputs(1772));
    layer8_outputs(4794) <= not(layer7_outputs(2803));
    layer8_outputs(4795) <= layer7_outputs(2566);
    layer8_outputs(4796) <= not(layer7_outputs(5030));
    layer8_outputs(4797) <= layer7_outputs(1745);
    layer8_outputs(4798) <= not((layer7_outputs(4570)) xor (layer7_outputs(2804)));
    layer8_outputs(4799) <= layer7_outputs(2371);
    layer8_outputs(4800) <= layer7_outputs(4318);
    layer8_outputs(4801) <= not(layer7_outputs(4431));
    layer8_outputs(4802) <= not((layer7_outputs(4801)) xor (layer7_outputs(3260)));
    layer8_outputs(4803) <= (layer7_outputs(2462)) and not (layer7_outputs(2594));
    layer8_outputs(4804) <= not(layer7_outputs(3380));
    layer8_outputs(4805) <= (layer7_outputs(1308)) and not (layer7_outputs(1427));
    layer8_outputs(4806) <= layer7_outputs(4504);
    layer8_outputs(4807) <= (layer7_outputs(2419)) and not (layer7_outputs(2387));
    layer8_outputs(4808) <= (layer7_outputs(2556)) and (layer7_outputs(4351));
    layer8_outputs(4809) <= layer7_outputs(117);
    layer8_outputs(4810) <= not(layer7_outputs(4353)) or (layer7_outputs(3454));
    layer8_outputs(4811) <= (layer7_outputs(1284)) xor (layer7_outputs(1264));
    layer8_outputs(4812) <= layer7_outputs(3922);
    layer8_outputs(4813) <= not((layer7_outputs(676)) xor (layer7_outputs(377)));
    layer8_outputs(4814) <= not(layer7_outputs(3475));
    layer8_outputs(4815) <= layer7_outputs(3141);
    layer8_outputs(4816) <= (layer7_outputs(2719)) and (layer7_outputs(37));
    layer8_outputs(4817) <= layer7_outputs(2393);
    layer8_outputs(4818) <= not((layer7_outputs(795)) xor (layer7_outputs(3323)));
    layer8_outputs(4819) <= layer7_outputs(2045);
    layer8_outputs(4820) <= not(layer7_outputs(1948));
    layer8_outputs(4821) <= (layer7_outputs(2273)) and not (layer7_outputs(2266));
    layer8_outputs(4822) <= not((layer7_outputs(4768)) or (layer7_outputs(3259)));
    layer8_outputs(4823) <= layer7_outputs(2220);
    layer8_outputs(4824) <= not(layer7_outputs(785)) or (layer7_outputs(3060));
    layer8_outputs(4825) <= layer7_outputs(3653);
    layer8_outputs(4826) <= (layer7_outputs(1492)) or (layer7_outputs(4073));
    layer8_outputs(4827) <= (layer7_outputs(2372)) and not (layer7_outputs(3243));
    layer8_outputs(4828) <= not((layer7_outputs(2622)) and (layer7_outputs(4502)));
    layer8_outputs(4829) <= (layer7_outputs(4017)) and not (layer7_outputs(897));
    layer8_outputs(4830) <= not(layer7_outputs(4035));
    layer8_outputs(4831) <= not((layer7_outputs(1030)) or (layer7_outputs(2111)));
    layer8_outputs(4832) <= not(layer7_outputs(1695));
    layer8_outputs(4833) <= (layer7_outputs(3700)) xor (layer7_outputs(4884));
    layer8_outputs(4834) <= layer7_outputs(1066);
    layer8_outputs(4835) <= not(layer7_outputs(3735));
    layer8_outputs(4836) <= layer7_outputs(2333);
    layer8_outputs(4837) <= not(layer7_outputs(1610));
    layer8_outputs(4838) <= not((layer7_outputs(929)) xor (layer7_outputs(4765)));
    layer8_outputs(4839) <= (layer7_outputs(3189)) xor (layer7_outputs(3290));
    layer8_outputs(4840) <= not((layer7_outputs(3234)) xor (layer7_outputs(739)));
    layer8_outputs(4841) <= (layer7_outputs(1070)) xor (layer7_outputs(3015));
    layer8_outputs(4842) <= (layer7_outputs(3040)) xor (layer7_outputs(1656));
    layer8_outputs(4843) <= not(layer7_outputs(493));
    layer8_outputs(4844) <= not(layer7_outputs(2833));
    layer8_outputs(4845) <= layer7_outputs(1592);
    layer8_outputs(4846) <= layer7_outputs(4394);
    layer8_outputs(4847) <= not(layer7_outputs(2926));
    layer8_outputs(4848) <= not(layer7_outputs(4204));
    layer8_outputs(4849) <= not(layer7_outputs(3185));
    layer8_outputs(4850) <= layer7_outputs(4780);
    layer8_outputs(4851) <= not((layer7_outputs(2957)) or (layer7_outputs(4111)));
    layer8_outputs(4852) <= not((layer7_outputs(4604)) and (layer7_outputs(2627)));
    layer8_outputs(4853) <= not(layer7_outputs(4422)) or (layer7_outputs(4228));
    layer8_outputs(4854) <= not((layer7_outputs(2844)) xor (layer7_outputs(717)));
    layer8_outputs(4855) <= not(layer7_outputs(4955));
    layer8_outputs(4856) <= not((layer7_outputs(4249)) and (layer7_outputs(1466)));
    layer8_outputs(4857) <= layer7_outputs(5023);
    layer8_outputs(4858) <= layer7_outputs(2797);
    layer8_outputs(4859) <= (layer7_outputs(1886)) and not (layer7_outputs(598));
    layer8_outputs(4860) <= (layer7_outputs(2822)) xor (layer7_outputs(2720));
    layer8_outputs(4861) <= not(layer7_outputs(2921));
    layer8_outputs(4862) <= (layer7_outputs(5096)) and (layer7_outputs(1454));
    layer8_outputs(4863) <= (layer7_outputs(4769)) xor (layer7_outputs(5057));
    layer8_outputs(4864) <= (layer7_outputs(784)) and not (layer7_outputs(1557));
    layer8_outputs(4865) <= not(layer7_outputs(3684)) or (layer7_outputs(4995));
    layer8_outputs(4866) <= not(layer7_outputs(635)) or (layer7_outputs(3679));
    layer8_outputs(4867) <= layer7_outputs(1984);
    layer8_outputs(4868) <= not(layer7_outputs(5110));
    layer8_outputs(4869) <= not(layer7_outputs(4696));
    layer8_outputs(4870) <= '0';
    layer8_outputs(4871) <= not(layer7_outputs(394)) or (layer7_outputs(4506));
    layer8_outputs(4872) <= (layer7_outputs(2296)) or (layer7_outputs(894));
    layer8_outputs(4873) <= (layer7_outputs(2794)) xor (layer7_outputs(929));
    layer8_outputs(4874) <= not(layer7_outputs(4809)) or (layer7_outputs(3987));
    layer8_outputs(4875) <= layer7_outputs(1560);
    layer8_outputs(4876) <= (layer7_outputs(4887)) and not (layer7_outputs(2809));
    layer8_outputs(4877) <= layer7_outputs(2959);
    layer8_outputs(4878) <= '1';
    layer8_outputs(4879) <= layer7_outputs(3932);
    layer8_outputs(4880) <= (layer7_outputs(1900)) xor (layer7_outputs(4263));
    layer8_outputs(4881) <= (layer7_outputs(131)) and not (layer7_outputs(2541));
    layer8_outputs(4882) <= not((layer7_outputs(338)) xor (layer7_outputs(3714)));
    layer8_outputs(4883) <= not((layer7_outputs(3437)) and (layer7_outputs(623)));
    layer8_outputs(4884) <= (layer7_outputs(4455)) and not (layer7_outputs(1147));
    layer8_outputs(4885) <= not((layer7_outputs(252)) xor (layer7_outputs(1135)));
    layer8_outputs(4886) <= not(layer7_outputs(3983));
    layer8_outputs(4887) <= layer7_outputs(3028);
    layer8_outputs(4888) <= not(layer7_outputs(3778));
    layer8_outputs(4889) <= not((layer7_outputs(2501)) xor (layer7_outputs(3389)));
    layer8_outputs(4890) <= not(layer7_outputs(896));
    layer8_outputs(4891) <= not((layer7_outputs(3097)) xor (layer7_outputs(1428)));
    layer8_outputs(4892) <= layer7_outputs(2656);
    layer8_outputs(4893) <= not(layer7_outputs(2960));
    layer8_outputs(4894) <= layer7_outputs(4046);
    layer8_outputs(4895) <= layer7_outputs(4568);
    layer8_outputs(4896) <= not(layer7_outputs(3068)) or (layer7_outputs(1268));
    layer8_outputs(4897) <= (layer7_outputs(829)) xor (layer7_outputs(4346));
    layer8_outputs(4898) <= '0';
    layer8_outputs(4899) <= layer7_outputs(2095);
    layer8_outputs(4900) <= (layer7_outputs(4324)) or (layer7_outputs(346));
    layer8_outputs(4901) <= (layer7_outputs(3557)) and (layer7_outputs(4933));
    layer8_outputs(4902) <= not(layer7_outputs(3609)) or (layer7_outputs(2631));
    layer8_outputs(4903) <= layer7_outputs(532);
    layer8_outputs(4904) <= layer7_outputs(1474);
    layer8_outputs(4905) <= not(layer7_outputs(2428));
    layer8_outputs(4906) <= not((layer7_outputs(271)) or (layer7_outputs(4472)));
    layer8_outputs(4907) <= layer7_outputs(2894);
    layer8_outputs(4908) <= layer7_outputs(4598);
    layer8_outputs(4909) <= (layer7_outputs(2277)) xor (layer7_outputs(853));
    layer8_outputs(4910) <= not(layer7_outputs(2715));
    layer8_outputs(4911) <= layer7_outputs(1320);
    layer8_outputs(4912) <= not(layer7_outputs(414));
    layer8_outputs(4913) <= layer7_outputs(3902);
    layer8_outputs(4914) <= layer7_outputs(3774);
    layer8_outputs(4915) <= not(layer7_outputs(3270));
    layer8_outputs(4916) <= not(layer7_outputs(4408));
    layer8_outputs(4917) <= (layer7_outputs(4597)) or (layer7_outputs(2748));
    layer8_outputs(4918) <= not((layer7_outputs(2737)) xor (layer7_outputs(334)));
    layer8_outputs(4919) <= layer7_outputs(3076);
    layer8_outputs(4920) <= (layer7_outputs(45)) xor (layer7_outputs(1412));
    layer8_outputs(4921) <= not((layer7_outputs(1533)) and (layer7_outputs(1860)));
    layer8_outputs(4922) <= (layer7_outputs(4417)) or (layer7_outputs(755));
    layer8_outputs(4923) <= (layer7_outputs(2524)) and not (layer7_outputs(1580));
    layer8_outputs(4924) <= (layer7_outputs(4362)) xor (layer7_outputs(1129));
    layer8_outputs(4925) <= not(layer7_outputs(1919));
    layer8_outputs(4926) <= not(layer7_outputs(1716)) or (layer7_outputs(5037));
    layer8_outputs(4927) <= layer7_outputs(3110);
    layer8_outputs(4928) <= not(layer7_outputs(2442));
    layer8_outputs(4929) <= (layer7_outputs(1116)) and not (layer7_outputs(189));
    layer8_outputs(4930) <= layer7_outputs(1712);
    layer8_outputs(4931) <= layer7_outputs(2606);
    layer8_outputs(4932) <= (layer7_outputs(3511)) and not (layer7_outputs(2492));
    layer8_outputs(4933) <= layer7_outputs(3856);
    layer8_outputs(4934) <= not(layer7_outputs(2865));
    layer8_outputs(4935) <= layer7_outputs(4808);
    layer8_outputs(4936) <= not((layer7_outputs(185)) and (layer7_outputs(3909)));
    layer8_outputs(4937) <= layer7_outputs(752);
    layer8_outputs(4938) <= layer7_outputs(4925);
    layer8_outputs(4939) <= (layer7_outputs(3670)) xor (layer7_outputs(1224));
    layer8_outputs(4940) <= layer7_outputs(4998);
    layer8_outputs(4941) <= (layer7_outputs(3294)) and not (layer7_outputs(2290));
    layer8_outputs(4942) <= not((layer7_outputs(4469)) xor (layer7_outputs(860)));
    layer8_outputs(4943) <= (layer7_outputs(4412)) xor (layer7_outputs(2852));
    layer8_outputs(4944) <= not(layer7_outputs(4549));
    layer8_outputs(4945) <= not((layer7_outputs(1390)) or (layer7_outputs(924)));
    layer8_outputs(4946) <= not(layer7_outputs(488));
    layer8_outputs(4947) <= (layer7_outputs(3296)) and not (layer7_outputs(1702));
    layer8_outputs(4948) <= not(layer7_outputs(873));
    layer8_outputs(4949) <= (layer7_outputs(3054)) xor (layer7_outputs(5104));
    layer8_outputs(4950) <= not(layer7_outputs(4348));
    layer8_outputs(4951) <= layer7_outputs(2401);
    layer8_outputs(4952) <= layer7_outputs(956);
    layer8_outputs(4953) <= (layer7_outputs(4608)) xor (layer7_outputs(2673));
    layer8_outputs(4954) <= not((layer7_outputs(1152)) and (layer7_outputs(2229)));
    layer8_outputs(4955) <= not(layer7_outputs(2672));
    layer8_outputs(4956) <= '1';
    layer8_outputs(4957) <= (layer7_outputs(3764)) and not (layer7_outputs(3470));
    layer8_outputs(4958) <= not(layer7_outputs(1334)) or (layer7_outputs(3605));
    layer8_outputs(4959) <= not(layer7_outputs(2624));
    layer8_outputs(4960) <= (layer7_outputs(1797)) and (layer7_outputs(1859));
    layer8_outputs(4961) <= layer7_outputs(1961);
    layer8_outputs(4962) <= layer7_outputs(3137);
    layer8_outputs(4963) <= (layer7_outputs(4454)) and not (layer7_outputs(2304));
    layer8_outputs(4964) <= not((layer7_outputs(1251)) xor (layer7_outputs(4156)));
    layer8_outputs(4965) <= (layer7_outputs(991)) and not (layer7_outputs(4733));
    layer8_outputs(4966) <= not(layer7_outputs(4632));
    layer8_outputs(4967) <= (layer7_outputs(4864)) and not (layer7_outputs(1854));
    layer8_outputs(4968) <= layer7_outputs(2209);
    layer8_outputs(4969) <= not(layer7_outputs(2719)) or (layer7_outputs(5047));
    layer8_outputs(4970) <= layer7_outputs(22);
    layer8_outputs(4971) <= layer7_outputs(1568);
    layer8_outputs(4972) <= not((layer7_outputs(625)) xor (layer7_outputs(2196)));
    layer8_outputs(4973) <= not(layer7_outputs(4995));
    layer8_outputs(4974) <= not(layer7_outputs(4958)) or (layer7_outputs(3402));
    layer8_outputs(4975) <= not(layer7_outputs(4565));
    layer8_outputs(4976) <= layer7_outputs(4228);
    layer8_outputs(4977) <= (layer7_outputs(4173)) xor (layer7_outputs(3832));
    layer8_outputs(4978) <= not(layer7_outputs(1056));
    layer8_outputs(4979) <= layer7_outputs(2327);
    layer8_outputs(4980) <= layer7_outputs(4577);
    layer8_outputs(4981) <= (layer7_outputs(823)) and not (layer7_outputs(1965));
    layer8_outputs(4982) <= not((layer7_outputs(4266)) or (layer7_outputs(3118)));
    layer8_outputs(4983) <= layer7_outputs(439);
    layer8_outputs(4984) <= not(layer7_outputs(910));
    layer8_outputs(4985) <= not(layer7_outputs(1614));
    layer8_outputs(4986) <= (layer7_outputs(130)) xor (layer7_outputs(1282));
    layer8_outputs(4987) <= layer7_outputs(3556);
    layer8_outputs(4988) <= (layer7_outputs(938)) and not (layer7_outputs(1621));
    layer8_outputs(4989) <= '0';
    layer8_outputs(4990) <= layer7_outputs(2990);
    layer8_outputs(4991) <= not((layer7_outputs(1133)) xor (layer7_outputs(2115)));
    layer8_outputs(4992) <= layer7_outputs(4555);
    layer8_outputs(4993) <= not(layer7_outputs(2366)) or (layer7_outputs(3874));
    layer8_outputs(4994) <= (layer7_outputs(1723)) xor (layer7_outputs(1510));
    layer8_outputs(4995) <= layer7_outputs(32);
    layer8_outputs(4996) <= (layer7_outputs(972)) and not (layer7_outputs(1024));
    layer8_outputs(4997) <= not(layer7_outputs(404));
    layer8_outputs(4998) <= (layer7_outputs(864)) xor (layer7_outputs(4494));
    layer8_outputs(4999) <= not(layer7_outputs(3721));
    layer8_outputs(5000) <= not((layer7_outputs(4238)) and (layer7_outputs(1305)));
    layer8_outputs(5001) <= (layer7_outputs(2114)) or (layer7_outputs(421));
    layer8_outputs(5002) <= (layer7_outputs(4293)) and (layer7_outputs(306));
    layer8_outputs(5003) <= (layer7_outputs(515)) and not (layer7_outputs(4452));
    layer8_outputs(5004) <= layer7_outputs(1685);
    layer8_outputs(5005) <= (layer7_outputs(3087)) xor (layer7_outputs(96));
    layer8_outputs(5006) <= (layer7_outputs(1833)) or (layer7_outputs(356));
    layer8_outputs(5007) <= layer7_outputs(1451);
    layer8_outputs(5008) <= not((layer7_outputs(2638)) xor (layer7_outputs(2884)));
    layer8_outputs(5009) <= (layer7_outputs(4931)) and not (layer7_outputs(1937));
    layer8_outputs(5010) <= not((layer7_outputs(2927)) xor (layer7_outputs(390)));
    layer8_outputs(5011) <= layer7_outputs(4590);
    layer8_outputs(5012) <= layer7_outputs(1583);
    layer8_outputs(5013) <= not(layer7_outputs(3566));
    layer8_outputs(5014) <= not((layer7_outputs(4994)) xor (layer7_outputs(2337)));
    layer8_outputs(5015) <= layer7_outputs(5026);
    layer8_outputs(5016) <= (layer7_outputs(4920)) xor (layer7_outputs(3925));
    layer8_outputs(5017) <= layer7_outputs(3113);
    layer8_outputs(5018) <= not((layer7_outputs(2981)) xor (layer7_outputs(1913)));
    layer8_outputs(5019) <= not((layer7_outputs(19)) xor (layer7_outputs(713)));
    layer8_outputs(5020) <= not((layer7_outputs(3050)) xor (layer7_outputs(746)));
    layer8_outputs(5021) <= layer7_outputs(1846);
    layer8_outputs(5022) <= not((layer7_outputs(1401)) xor (layer7_outputs(986)));
    layer8_outputs(5023) <= (layer7_outputs(4727)) and (layer7_outputs(4062));
    layer8_outputs(5024) <= not((layer7_outputs(69)) xor (layer7_outputs(2321)));
    layer8_outputs(5025) <= layer7_outputs(1103);
    layer8_outputs(5026) <= layer7_outputs(2661);
    layer8_outputs(5027) <= (layer7_outputs(1631)) or (layer7_outputs(1921));
    layer8_outputs(5028) <= (layer7_outputs(3385)) xor (layer7_outputs(2535));
    layer8_outputs(5029) <= not((layer7_outputs(24)) or (layer7_outputs(4056)));
    layer8_outputs(5030) <= not(layer7_outputs(119));
    layer8_outputs(5031) <= layer7_outputs(4987);
    layer8_outputs(5032) <= not(layer7_outputs(2743));
    layer8_outputs(5033) <= (layer7_outputs(3764)) or (layer7_outputs(3373));
    layer8_outputs(5034) <= not((layer7_outputs(979)) xor (layer7_outputs(2034)));
    layer8_outputs(5035) <= not(layer7_outputs(1170));
    layer8_outputs(5036) <= not(layer7_outputs(2896));
    layer8_outputs(5037) <= (layer7_outputs(2455)) xor (layer7_outputs(2065));
    layer8_outputs(5038) <= layer7_outputs(771);
    layer8_outputs(5039) <= (layer7_outputs(856)) and (layer7_outputs(910));
    layer8_outputs(5040) <= not(layer7_outputs(284)) or (layer7_outputs(4354));
    layer8_outputs(5041) <= not((layer7_outputs(3499)) xor (layer7_outputs(2362)));
    layer8_outputs(5042) <= layer7_outputs(193);
    layer8_outputs(5043) <= not(layer7_outputs(969));
    layer8_outputs(5044) <= not((layer7_outputs(4218)) and (layer7_outputs(1726)));
    layer8_outputs(5045) <= (layer7_outputs(2285)) xor (layer7_outputs(2509));
    layer8_outputs(5046) <= not(layer7_outputs(856));
    layer8_outputs(5047) <= (layer7_outputs(4276)) and not (layer7_outputs(883));
    layer8_outputs(5048) <= layer7_outputs(1314);
    layer8_outputs(5049) <= not((layer7_outputs(3092)) and (layer7_outputs(3001)));
    layer8_outputs(5050) <= not((layer7_outputs(4545)) xor (layer7_outputs(389)));
    layer8_outputs(5051) <= layer7_outputs(4769);
    layer8_outputs(5052) <= not((layer7_outputs(4338)) xor (layer7_outputs(1883)));
    layer8_outputs(5053) <= not((layer7_outputs(2416)) xor (layer7_outputs(1339)));
    layer8_outputs(5054) <= not(layer7_outputs(1071));
    layer8_outputs(5055) <= layer7_outputs(1983);
    layer8_outputs(5056) <= not((layer7_outputs(3192)) xor (layer7_outputs(2770)));
    layer8_outputs(5057) <= not(layer7_outputs(1735));
    layer8_outputs(5058) <= layer7_outputs(1049);
    layer8_outputs(5059) <= layer7_outputs(1601);
    layer8_outputs(5060) <= not(layer7_outputs(5107));
    layer8_outputs(5061) <= (layer7_outputs(1963)) and not (layer7_outputs(1555));
    layer8_outputs(5062) <= not((layer7_outputs(3340)) and (layer7_outputs(2019)));
    layer8_outputs(5063) <= (layer7_outputs(4057)) and not (layer7_outputs(4055));
    layer8_outputs(5064) <= (layer7_outputs(1937)) or (layer7_outputs(1119));
    layer8_outputs(5065) <= (layer7_outputs(780)) xor (layer7_outputs(3857));
    layer8_outputs(5066) <= not((layer7_outputs(527)) or (layer7_outputs(2619)));
    layer8_outputs(5067) <= layer7_outputs(221);
    layer8_outputs(5068) <= not((layer7_outputs(4723)) or (layer7_outputs(3662)));
    layer8_outputs(5069) <= layer7_outputs(1419);
    layer8_outputs(5070) <= not(layer7_outputs(1820));
    layer8_outputs(5071) <= layer7_outputs(3571);
    layer8_outputs(5072) <= layer7_outputs(2827);
    layer8_outputs(5073) <= not(layer7_outputs(1652));
    layer8_outputs(5074) <= (layer7_outputs(1747)) xor (layer7_outputs(3907));
    layer8_outputs(5075) <= (layer7_outputs(518)) xor (layer7_outputs(2436));
    layer8_outputs(5076) <= (layer7_outputs(3588)) xor (layer7_outputs(4292));
    layer8_outputs(5077) <= layer7_outputs(4429);
    layer8_outputs(5078) <= not((layer7_outputs(2618)) xor (layer7_outputs(2792)));
    layer8_outputs(5079) <= layer7_outputs(1757);
    layer8_outputs(5080) <= layer7_outputs(3927);
    layer8_outputs(5081) <= not(layer7_outputs(2729)) or (layer7_outputs(1121));
    layer8_outputs(5082) <= not((layer7_outputs(4960)) or (layer7_outputs(4771)));
    layer8_outputs(5083) <= not(layer7_outputs(4401));
    layer8_outputs(5084) <= (layer7_outputs(1782)) and (layer7_outputs(4750));
    layer8_outputs(5085) <= (layer7_outputs(1086)) or (layer7_outputs(2761));
    layer8_outputs(5086) <= (layer7_outputs(3522)) and (layer7_outputs(4361));
    layer8_outputs(5087) <= (layer7_outputs(1966)) and not (layer7_outputs(1738));
    layer8_outputs(5088) <= (layer7_outputs(2766)) and not (layer7_outputs(1168));
    layer8_outputs(5089) <= not(layer7_outputs(1364));
    layer8_outputs(5090) <= not(layer7_outputs(3761));
    layer8_outputs(5091) <= (layer7_outputs(3196)) xor (layer7_outputs(1361));
    layer8_outputs(5092) <= not(layer7_outputs(2382)) or (layer7_outputs(1982));
    layer8_outputs(5093) <= not(layer7_outputs(3456));
    layer8_outputs(5094) <= not(layer7_outputs(1344));
    layer8_outputs(5095) <= (layer7_outputs(2480)) and not (layer7_outputs(2573));
    layer8_outputs(5096) <= not(layer7_outputs(751));
    layer8_outputs(5097) <= not(layer7_outputs(4585));
    layer8_outputs(5098) <= not(layer7_outputs(1168));
    layer8_outputs(5099) <= (layer7_outputs(2167)) and not (layer7_outputs(822));
    layer8_outputs(5100) <= layer7_outputs(400);
    layer8_outputs(5101) <= (layer7_outputs(3527)) xor (layer7_outputs(2031));
    layer8_outputs(5102) <= layer7_outputs(2742);
    layer8_outputs(5103) <= (layer7_outputs(4247)) and not (layer7_outputs(4548));
    layer8_outputs(5104) <= layer7_outputs(5092);
    layer8_outputs(5105) <= (layer7_outputs(1106)) and (layer7_outputs(1415));
    layer8_outputs(5106) <= not((layer7_outputs(4379)) xor (layer7_outputs(2985)));
    layer8_outputs(5107) <= (layer7_outputs(4180)) xor (layer7_outputs(4886));
    layer8_outputs(5108) <= (layer7_outputs(3971)) xor (layer7_outputs(2799));
    layer8_outputs(5109) <= not(layer7_outputs(4465)) or (layer7_outputs(630));
    layer8_outputs(5110) <= not((layer7_outputs(1920)) xor (layer7_outputs(1205)));
    layer8_outputs(5111) <= '0';
    layer8_outputs(5112) <= not(layer7_outputs(3897));
    layer8_outputs(5113) <= layer7_outputs(4347);
    layer8_outputs(5114) <= (layer7_outputs(1201)) and (layer7_outputs(4916));
    layer8_outputs(5115) <= (layer7_outputs(1857)) xor (layer7_outputs(2464));
    layer8_outputs(5116) <= '0';
    layer8_outputs(5117) <= (layer7_outputs(4793)) and not (layer7_outputs(3479));
    layer8_outputs(5118) <= not(layer7_outputs(2339));
    layer8_outputs(5119) <= not(layer7_outputs(4875));
    outputs(0) <= (layer8_outputs(1745)) or (layer8_outputs(930));
    outputs(1) <= not(layer8_outputs(4509));
    outputs(2) <= layer8_outputs(184);
    outputs(3) <= not((layer8_outputs(2100)) xor (layer8_outputs(2475)));
    outputs(4) <= not(layer8_outputs(2719));
    outputs(5) <= layer8_outputs(3485);
    outputs(6) <= not(layer8_outputs(1741));
    outputs(7) <= layer8_outputs(3122);
    outputs(8) <= layer8_outputs(2425);
    outputs(9) <= (layer8_outputs(1345)) and (layer8_outputs(2845));
    outputs(10) <= layer8_outputs(2100);
    outputs(11) <= not(layer8_outputs(2656));
    outputs(12) <= not(layer8_outputs(696));
    outputs(13) <= not(layer8_outputs(4948));
    outputs(14) <= layer8_outputs(1706);
    outputs(15) <= (layer8_outputs(1308)) xor (layer8_outputs(1081));
    outputs(16) <= layer8_outputs(3382);
    outputs(17) <= not(layer8_outputs(1059));
    outputs(18) <= not((layer8_outputs(336)) or (layer8_outputs(85)));
    outputs(19) <= layer8_outputs(2583);
    outputs(20) <= not(layer8_outputs(3572));
    outputs(21) <= not(layer8_outputs(4546)) or (layer8_outputs(86));
    outputs(22) <= layer8_outputs(1038);
    outputs(23) <= not((layer8_outputs(3830)) and (layer8_outputs(1553)));
    outputs(24) <= not((layer8_outputs(3538)) xor (layer8_outputs(4157)));
    outputs(25) <= layer8_outputs(1403);
    outputs(26) <= not((layer8_outputs(653)) xor (layer8_outputs(3961)));
    outputs(27) <= layer8_outputs(2124);
    outputs(28) <= (layer8_outputs(872)) and (layer8_outputs(515));
    outputs(29) <= (layer8_outputs(521)) and not (layer8_outputs(3146));
    outputs(30) <= (layer8_outputs(3234)) or (layer8_outputs(2850));
    outputs(31) <= layer8_outputs(3131);
    outputs(32) <= not(layer8_outputs(1091));
    outputs(33) <= not((layer8_outputs(4029)) xor (layer8_outputs(2322)));
    outputs(34) <= not(layer8_outputs(4885));
    outputs(35) <= not((layer8_outputs(4277)) or (layer8_outputs(3509)));
    outputs(36) <= layer8_outputs(2204);
    outputs(37) <= not(layer8_outputs(3775));
    outputs(38) <= layer8_outputs(2700);
    outputs(39) <= not(layer8_outputs(632)) or (layer8_outputs(3799));
    outputs(40) <= layer8_outputs(3408);
    outputs(41) <= not(layer8_outputs(3173)) or (layer8_outputs(2582));
    outputs(42) <= not(layer8_outputs(1486));
    outputs(43) <= not(layer8_outputs(1085)) or (layer8_outputs(3661));
    outputs(44) <= layer8_outputs(1040);
    outputs(45) <= not(layer8_outputs(4226));
    outputs(46) <= (layer8_outputs(1569)) xor (layer8_outputs(2301));
    outputs(47) <= not(layer8_outputs(4106));
    outputs(48) <= (layer8_outputs(660)) xor (layer8_outputs(2037));
    outputs(49) <= layer8_outputs(4471);
    outputs(50) <= layer8_outputs(1379);
    outputs(51) <= not(layer8_outputs(565));
    outputs(52) <= (layer8_outputs(4290)) xor (layer8_outputs(4051));
    outputs(53) <= not(layer8_outputs(3289));
    outputs(54) <= not(layer8_outputs(387));
    outputs(55) <= not((layer8_outputs(2350)) xor (layer8_outputs(623)));
    outputs(56) <= not(layer8_outputs(3125)) or (layer8_outputs(2760));
    outputs(57) <= layer8_outputs(281);
    outputs(58) <= not((layer8_outputs(688)) or (layer8_outputs(487)));
    outputs(59) <= (layer8_outputs(2598)) and not (layer8_outputs(398));
    outputs(60) <= (layer8_outputs(1686)) and not (layer8_outputs(4234));
    outputs(61) <= not((layer8_outputs(3926)) xor (layer8_outputs(2893)));
    outputs(62) <= (layer8_outputs(1350)) xor (layer8_outputs(1185));
    outputs(63) <= not((layer8_outputs(2574)) and (layer8_outputs(4490)));
    outputs(64) <= not(layer8_outputs(1980));
    outputs(65) <= (layer8_outputs(168)) xor (layer8_outputs(1807));
    outputs(66) <= not(layer8_outputs(476)) or (layer8_outputs(4724));
    outputs(67) <= (layer8_outputs(2771)) xor (layer8_outputs(656));
    outputs(68) <= not((layer8_outputs(2159)) xor (layer8_outputs(3720)));
    outputs(69) <= not(layer8_outputs(4873));
    outputs(70) <= not((layer8_outputs(282)) and (layer8_outputs(1022)));
    outputs(71) <= not((layer8_outputs(1264)) xor (layer8_outputs(841)));
    outputs(72) <= layer8_outputs(277);
    outputs(73) <= layer8_outputs(3023);
    outputs(74) <= not(layer8_outputs(306));
    outputs(75) <= (layer8_outputs(1614)) xor (layer8_outputs(1285));
    outputs(76) <= layer8_outputs(3460);
    outputs(77) <= not(layer8_outputs(3045));
    outputs(78) <= layer8_outputs(1228);
    outputs(79) <= layer8_outputs(3018);
    outputs(80) <= not((layer8_outputs(2198)) xor (layer8_outputs(1291)));
    outputs(81) <= layer8_outputs(3170);
    outputs(82) <= not((layer8_outputs(737)) or (layer8_outputs(2794)));
    outputs(83) <= (layer8_outputs(459)) xor (layer8_outputs(1054));
    outputs(84) <= not(layer8_outputs(1861));
    outputs(85) <= layer8_outputs(1793);
    outputs(86) <= not((layer8_outputs(427)) xor (layer8_outputs(3166)));
    outputs(87) <= not(layer8_outputs(154));
    outputs(88) <= layer8_outputs(4807);
    outputs(89) <= not((layer8_outputs(1381)) xor (layer8_outputs(3355)));
    outputs(90) <= not(layer8_outputs(1183));
    outputs(91) <= layer8_outputs(514);
    outputs(92) <= layer8_outputs(3875);
    outputs(93) <= layer8_outputs(1069);
    outputs(94) <= layer8_outputs(4109);
    outputs(95) <= not(layer8_outputs(4565));
    outputs(96) <= layer8_outputs(665);
    outputs(97) <= not((layer8_outputs(1382)) xor (layer8_outputs(2810)));
    outputs(98) <= not((layer8_outputs(853)) xor (layer8_outputs(3371)));
    outputs(99) <= layer8_outputs(1469);
    outputs(100) <= layer8_outputs(2174);
    outputs(101) <= (layer8_outputs(802)) xor (layer8_outputs(2778));
    outputs(102) <= layer8_outputs(4994);
    outputs(103) <= layer8_outputs(4093);
    outputs(104) <= not((layer8_outputs(625)) xor (layer8_outputs(1271)));
    outputs(105) <= (layer8_outputs(1208)) and not (layer8_outputs(377));
    outputs(106) <= not(layer8_outputs(121));
    outputs(107) <= (layer8_outputs(2711)) and not (layer8_outputs(4010));
    outputs(108) <= not((layer8_outputs(1954)) xor (layer8_outputs(4707)));
    outputs(109) <= not(layer8_outputs(3019));
    outputs(110) <= layer8_outputs(2921);
    outputs(111) <= not(layer8_outputs(2176));
    outputs(112) <= layer8_outputs(3109);
    outputs(113) <= layer8_outputs(705);
    outputs(114) <= (layer8_outputs(3429)) or (layer8_outputs(4373));
    outputs(115) <= not(layer8_outputs(4826));
    outputs(116) <= not((layer8_outputs(622)) xor (layer8_outputs(4948)));
    outputs(117) <= layer8_outputs(1693);
    outputs(118) <= layer8_outputs(2197);
    outputs(119) <= not(layer8_outputs(1109));
    outputs(120) <= not(layer8_outputs(2060));
    outputs(121) <= not(layer8_outputs(3652));
    outputs(122) <= (layer8_outputs(663)) xor (layer8_outputs(487));
    outputs(123) <= layer8_outputs(3225);
    outputs(124) <= layer8_outputs(3123);
    outputs(125) <= not(layer8_outputs(1971));
    outputs(126) <= not((layer8_outputs(2858)) xor (layer8_outputs(4596)));
    outputs(127) <= not((layer8_outputs(4464)) or (layer8_outputs(314)));
    outputs(128) <= (layer8_outputs(2857)) xor (layer8_outputs(1447));
    outputs(129) <= (layer8_outputs(3079)) and not (layer8_outputs(4231));
    outputs(130) <= layer8_outputs(277);
    outputs(131) <= layer8_outputs(1126);
    outputs(132) <= not(layer8_outputs(1448));
    outputs(133) <= not(layer8_outputs(3280));
    outputs(134) <= not(layer8_outputs(2062));
    outputs(135) <= layer8_outputs(4503);
    outputs(136) <= (layer8_outputs(5100)) and not (layer8_outputs(4361));
    outputs(137) <= not(layer8_outputs(2572)) or (layer8_outputs(4989));
    outputs(138) <= not((layer8_outputs(1056)) or (layer8_outputs(3243)));
    outputs(139) <= (layer8_outputs(2597)) xor (layer8_outputs(485));
    outputs(140) <= not(layer8_outputs(4155));
    outputs(141) <= not(layer8_outputs(4461));
    outputs(142) <= not((layer8_outputs(2987)) or (layer8_outputs(3879)));
    outputs(143) <= layer8_outputs(3377);
    outputs(144) <= not(layer8_outputs(702));
    outputs(145) <= layer8_outputs(907);
    outputs(146) <= not(layer8_outputs(2355));
    outputs(147) <= layer8_outputs(3204);
    outputs(148) <= layer8_outputs(1814);
    outputs(149) <= not((layer8_outputs(2872)) xor (layer8_outputs(4655)));
    outputs(150) <= layer8_outputs(2362);
    outputs(151) <= not(layer8_outputs(1990));
    outputs(152) <= not(layer8_outputs(4602));
    outputs(153) <= (layer8_outputs(3638)) and (layer8_outputs(437));
    outputs(154) <= layer8_outputs(5051);
    outputs(155) <= (layer8_outputs(402)) and not (layer8_outputs(4305));
    outputs(156) <= (layer8_outputs(1943)) xor (layer8_outputs(4423));
    outputs(157) <= not(layer8_outputs(2814));
    outputs(158) <= layer8_outputs(5013);
    outputs(159) <= not(layer8_outputs(1270));
    outputs(160) <= (layer8_outputs(2839)) xor (layer8_outputs(962));
    outputs(161) <= not(layer8_outputs(4339));
    outputs(162) <= not((layer8_outputs(2610)) xor (layer8_outputs(3770)));
    outputs(163) <= (layer8_outputs(2148)) xor (layer8_outputs(327));
    outputs(164) <= not((layer8_outputs(2006)) xor (layer8_outputs(4316)));
    outputs(165) <= layer8_outputs(3984);
    outputs(166) <= not((layer8_outputs(2786)) xor (layer8_outputs(4117)));
    outputs(167) <= layer8_outputs(1019);
    outputs(168) <= not((layer8_outputs(4667)) or (layer8_outputs(2521)));
    outputs(169) <= layer8_outputs(450);
    outputs(170) <= layer8_outputs(4960);
    outputs(171) <= layer8_outputs(3440);
    outputs(172) <= not((layer8_outputs(4344)) xor (layer8_outputs(135)));
    outputs(173) <= not((layer8_outputs(4374)) and (layer8_outputs(4974)));
    outputs(174) <= not(layer8_outputs(4723));
    outputs(175) <= (layer8_outputs(1537)) xor (layer8_outputs(31));
    outputs(176) <= not((layer8_outputs(396)) xor (layer8_outputs(3597)));
    outputs(177) <= not(layer8_outputs(1127));
    outputs(178) <= layer8_outputs(933);
    outputs(179) <= layer8_outputs(249);
    outputs(180) <= not(layer8_outputs(2468));
    outputs(181) <= not(layer8_outputs(3477));
    outputs(182) <= layer8_outputs(3525);
    outputs(183) <= not((layer8_outputs(2269)) and (layer8_outputs(4668)));
    outputs(184) <= (layer8_outputs(1858)) and (layer8_outputs(338));
    outputs(185) <= not(layer8_outputs(3662));
    outputs(186) <= layer8_outputs(355);
    outputs(187) <= (layer8_outputs(1163)) and not (layer8_outputs(130));
    outputs(188) <= not((layer8_outputs(4107)) xor (layer8_outputs(2590)));
    outputs(189) <= not(layer8_outputs(3973));
    outputs(190) <= (layer8_outputs(288)) and not (layer8_outputs(2367));
    outputs(191) <= layer8_outputs(1424);
    outputs(192) <= not(layer8_outputs(4657));
    outputs(193) <= not((layer8_outputs(1996)) xor (layer8_outputs(4245)));
    outputs(194) <= not(layer8_outputs(1463));
    outputs(195) <= layer8_outputs(228);
    outputs(196) <= not((layer8_outputs(74)) or (layer8_outputs(1547)));
    outputs(197) <= not(layer8_outputs(1838));
    outputs(198) <= (layer8_outputs(984)) xor (layer8_outputs(4212));
    outputs(199) <= layer8_outputs(3491);
    outputs(200) <= not(layer8_outputs(132));
    outputs(201) <= not(layer8_outputs(4694));
    outputs(202) <= not(layer8_outputs(2130));
    outputs(203) <= layer8_outputs(1322);
    outputs(204) <= (layer8_outputs(4248)) or (layer8_outputs(938));
    outputs(205) <= not((layer8_outputs(3465)) xor (layer8_outputs(1623)));
    outputs(206) <= layer8_outputs(141);
    outputs(207) <= not(layer8_outputs(3068));
    outputs(208) <= layer8_outputs(3050);
    outputs(209) <= layer8_outputs(2653);
    outputs(210) <= (layer8_outputs(4023)) and not (layer8_outputs(4140));
    outputs(211) <= layer8_outputs(2958);
    outputs(212) <= not(layer8_outputs(2951));
    outputs(213) <= not(layer8_outputs(2805));
    outputs(214) <= layer8_outputs(3582);
    outputs(215) <= not(layer8_outputs(3844));
    outputs(216) <= layer8_outputs(4517);
    outputs(217) <= layer8_outputs(3726);
    outputs(218) <= layer8_outputs(1418);
    outputs(219) <= not(layer8_outputs(3135));
    outputs(220) <= not((layer8_outputs(4589)) or (layer8_outputs(1913)));
    outputs(221) <= not(layer8_outputs(3645));
    outputs(222) <= not(layer8_outputs(1768));
    outputs(223) <= not((layer8_outputs(2045)) and (layer8_outputs(1873)));
    outputs(224) <= layer8_outputs(873);
    outputs(225) <= layer8_outputs(3076);
    outputs(226) <= not(layer8_outputs(70));
    outputs(227) <= layer8_outputs(5080);
    outputs(228) <= not(layer8_outputs(1352));
    outputs(229) <= (layer8_outputs(2307)) xor (layer8_outputs(3893));
    outputs(230) <= not(layer8_outputs(3236));
    outputs(231) <= not(layer8_outputs(1079));
    outputs(232) <= not((layer8_outputs(2576)) or (layer8_outputs(2231)));
    outputs(233) <= layer8_outputs(1839);
    outputs(234) <= layer8_outputs(1790);
    outputs(235) <= layer8_outputs(3741);
    outputs(236) <= layer8_outputs(4802);
    outputs(237) <= not((layer8_outputs(4728)) xor (layer8_outputs(1739)));
    outputs(238) <= layer8_outputs(976);
    outputs(239) <= layer8_outputs(3574);
    outputs(240) <= (layer8_outputs(4195)) and not (layer8_outputs(1310));
    outputs(241) <= not(layer8_outputs(3102));
    outputs(242) <= not(layer8_outputs(1359));
    outputs(243) <= not((layer8_outputs(4782)) or (layer8_outputs(106)));
    outputs(244) <= layer8_outputs(2494);
    outputs(245) <= layer8_outputs(451);
    outputs(246) <= not(layer8_outputs(798));
    outputs(247) <= not(layer8_outputs(2854));
    outputs(248) <= not(layer8_outputs(742));
    outputs(249) <= layer8_outputs(2976);
    outputs(250) <= not(layer8_outputs(130));
    outputs(251) <= layer8_outputs(3786);
    outputs(252) <= not(layer8_outputs(3672));
    outputs(253) <= not(layer8_outputs(4295));
    outputs(254) <= not((layer8_outputs(1707)) xor (layer8_outputs(1158)));
    outputs(255) <= layer8_outputs(225);
    outputs(256) <= (layer8_outputs(3790)) xor (layer8_outputs(4097));
    outputs(257) <= not(layer8_outputs(1895));
    outputs(258) <= (layer8_outputs(1346)) xor (layer8_outputs(2351));
    outputs(259) <= not(layer8_outputs(4040));
    outputs(260) <= layer8_outputs(1042);
    outputs(261) <= layer8_outputs(837);
    outputs(262) <= layer8_outputs(4855);
    outputs(263) <= not(layer8_outputs(1953));
    outputs(264) <= not(layer8_outputs(1850));
    outputs(265) <= not(layer8_outputs(1899));
    outputs(266) <= not(layer8_outputs(507)) or (layer8_outputs(1323));
    outputs(267) <= not(layer8_outputs(1495));
    outputs(268) <= not((layer8_outputs(2698)) xor (layer8_outputs(175)));
    outputs(269) <= not(layer8_outputs(1997));
    outputs(270) <= layer8_outputs(1036);
    outputs(271) <= layer8_outputs(4649);
    outputs(272) <= layer8_outputs(1160);
    outputs(273) <= not(layer8_outputs(827));
    outputs(274) <= (layer8_outputs(1422)) xor (layer8_outputs(1917));
    outputs(275) <= not(layer8_outputs(3209));
    outputs(276) <= not(layer8_outputs(3996));
    outputs(277) <= layer8_outputs(3823);
    outputs(278) <= layer8_outputs(2156);
    outputs(279) <= layer8_outputs(3882);
    outputs(280) <= not(layer8_outputs(1484));
    outputs(281) <= not((layer8_outputs(1869)) or (layer8_outputs(3424)));
    outputs(282) <= not((layer8_outputs(965)) xor (layer8_outputs(1940)));
    outputs(283) <= layer8_outputs(2440);
    outputs(284) <= layer8_outputs(1915);
    outputs(285) <= layer8_outputs(3984);
    outputs(286) <= not((layer8_outputs(1488)) xor (layer8_outputs(2512)));
    outputs(287) <= not(layer8_outputs(88));
    outputs(288) <= (layer8_outputs(259)) and not (layer8_outputs(856));
    outputs(289) <= not((layer8_outputs(1957)) or (layer8_outputs(4971)));
    outputs(290) <= (layer8_outputs(4858)) xor (layer8_outputs(3199));
    outputs(291) <= not(layer8_outputs(4277));
    outputs(292) <= not(layer8_outputs(261));
    outputs(293) <= layer8_outputs(1069);
    outputs(294) <= layer8_outputs(2595);
    outputs(295) <= not((layer8_outputs(4827)) xor (layer8_outputs(438)));
    outputs(296) <= not(layer8_outputs(4551));
    outputs(297) <= not(layer8_outputs(3406));
    outputs(298) <= not(layer8_outputs(3618));
    outputs(299) <= layer8_outputs(4371);
    outputs(300) <= not((layer8_outputs(2264)) xor (layer8_outputs(2784)));
    outputs(301) <= layer8_outputs(1104);
    outputs(302) <= not(layer8_outputs(3842)) or (layer8_outputs(2848));
    outputs(303) <= not((layer8_outputs(2741)) xor (layer8_outputs(4476)));
    outputs(304) <= layer8_outputs(4130);
    outputs(305) <= not(layer8_outputs(4500));
    outputs(306) <= (layer8_outputs(2025)) or (layer8_outputs(4652));
    outputs(307) <= not((layer8_outputs(3959)) xor (layer8_outputs(3868)));
    outputs(308) <= (layer8_outputs(1592)) xor (layer8_outputs(4926));
    outputs(309) <= not((layer8_outputs(4421)) xor (layer8_outputs(2564)));
    outputs(310) <= layer8_outputs(1164);
    outputs(311) <= (layer8_outputs(2687)) xor (layer8_outputs(76));
    outputs(312) <= not(layer8_outputs(2267));
    outputs(313) <= not(layer8_outputs(3425));
    outputs(314) <= (layer8_outputs(1819)) and (layer8_outputs(3237));
    outputs(315) <= layer8_outputs(878);
    outputs(316) <= not((layer8_outputs(311)) xor (layer8_outputs(509)));
    outputs(317) <= layer8_outputs(353);
    outputs(318) <= layer8_outputs(4293);
    outputs(319) <= not(layer8_outputs(2418)) or (layer8_outputs(815));
    outputs(320) <= (layer8_outputs(669)) or (layer8_outputs(4584));
    outputs(321) <= layer8_outputs(1469);
    outputs(322) <= (layer8_outputs(571)) xor (layer8_outputs(362));
    outputs(323) <= not((layer8_outputs(1083)) xor (layer8_outputs(4592)));
    outputs(324) <= layer8_outputs(4618);
    outputs(325) <= not(layer8_outputs(1056));
    outputs(326) <= (layer8_outputs(5117)) xor (layer8_outputs(4753));
    outputs(327) <= not((layer8_outputs(3810)) xor (layer8_outputs(2431)));
    outputs(328) <= not(layer8_outputs(4645));
    outputs(329) <= not(layer8_outputs(1744));
    outputs(330) <= layer8_outputs(3908);
    outputs(331) <= (layer8_outputs(1464)) and not (layer8_outputs(3343));
    outputs(332) <= layer8_outputs(2329);
    outputs(333) <= layer8_outputs(2177);
    outputs(334) <= (layer8_outputs(300)) xor (layer8_outputs(1250));
    outputs(335) <= not(layer8_outputs(1133));
    outputs(336) <= not((layer8_outputs(1109)) xor (layer8_outputs(4506)));
    outputs(337) <= not((layer8_outputs(4143)) xor (layer8_outputs(2617)));
    outputs(338) <= not(layer8_outputs(1590)) or (layer8_outputs(4233));
    outputs(339) <= not(layer8_outputs(2120));
    outputs(340) <= (layer8_outputs(823)) xor (layer8_outputs(875));
    outputs(341) <= not((layer8_outputs(2032)) or (layer8_outputs(4138)));
    outputs(342) <= layer8_outputs(349);
    outputs(343) <= not(layer8_outputs(2294));
    outputs(344) <= layer8_outputs(642);
    outputs(345) <= not(layer8_outputs(2854));
    outputs(346) <= not((layer8_outputs(169)) xor (layer8_outputs(1888)));
    outputs(347) <= not(layer8_outputs(2062));
    outputs(348) <= layer8_outputs(3479);
    outputs(349) <= (layer8_outputs(3619)) xor (layer8_outputs(2141));
    outputs(350) <= not(layer8_outputs(4190));
    outputs(351) <= not(layer8_outputs(194));
    outputs(352) <= not((layer8_outputs(17)) xor (layer8_outputs(4691)));
    outputs(353) <= not(layer8_outputs(1957));
    outputs(354) <= not(layer8_outputs(3685));
    outputs(355) <= not(layer8_outputs(1016)) or (layer8_outputs(770));
    outputs(356) <= (layer8_outputs(514)) and not (layer8_outputs(2317));
    outputs(357) <= layer8_outputs(741);
    outputs(358) <= not(layer8_outputs(3640));
    outputs(359) <= not((layer8_outputs(3278)) xor (layer8_outputs(3688)));
    outputs(360) <= (layer8_outputs(4121)) and not (layer8_outputs(1941));
    outputs(361) <= not(layer8_outputs(1127));
    outputs(362) <= not((layer8_outputs(161)) xor (layer8_outputs(1223)));
    outputs(363) <= not(layer8_outputs(2514));
    outputs(364) <= layer8_outputs(3957);
    outputs(365) <= not((layer8_outputs(619)) or (layer8_outputs(4438)));
    outputs(366) <= layer8_outputs(957);
    outputs(367) <= not(layer8_outputs(547));
    outputs(368) <= (layer8_outputs(327)) xor (layer8_outputs(4715));
    outputs(369) <= not(layer8_outputs(3683));
    outputs(370) <= not(layer8_outputs(2547));
    outputs(371) <= layer8_outputs(1403);
    outputs(372) <= layer8_outputs(2052);
    outputs(373) <= (layer8_outputs(3449)) and (layer8_outputs(3611));
    outputs(374) <= (layer8_outputs(4709)) xor (layer8_outputs(1183));
    outputs(375) <= layer8_outputs(1070);
    outputs(376) <= not((layer8_outputs(710)) xor (layer8_outputs(2292)));
    outputs(377) <= not(layer8_outputs(2980));
    outputs(378) <= not(layer8_outputs(1237));
    outputs(379) <= layer8_outputs(3869);
    outputs(380) <= not((layer8_outputs(2684)) xor (layer8_outputs(3678)));
    outputs(381) <= not((layer8_outputs(3961)) xor (layer8_outputs(1158)));
    outputs(382) <= layer8_outputs(3317);
    outputs(383) <= (layer8_outputs(4878)) and not (layer8_outputs(3659));
    outputs(384) <= not(layer8_outputs(3017));
    outputs(385) <= (layer8_outputs(764)) xor (layer8_outputs(3172));
    outputs(386) <= (layer8_outputs(426)) xor (layer8_outputs(4841));
    outputs(387) <= (layer8_outputs(1289)) and not (layer8_outputs(3118));
    outputs(388) <= not(layer8_outputs(3113));
    outputs(389) <= not((layer8_outputs(4026)) xor (layer8_outputs(1588)));
    outputs(390) <= not(layer8_outputs(2627)) or (layer8_outputs(4506));
    outputs(391) <= not((layer8_outputs(5097)) or (layer8_outputs(4884)));
    outputs(392) <= not((layer8_outputs(2238)) and (layer8_outputs(3596)));
    outputs(393) <= layer8_outputs(3954);
    outputs(394) <= (layer8_outputs(1139)) and (layer8_outputs(4089));
    outputs(395) <= not(layer8_outputs(1714));
    outputs(396) <= layer8_outputs(4388);
    outputs(397) <= layer8_outputs(1233);
    outputs(398) <= not((layer8_outputs(4829)) xor (layer8_outputs(861)));
    outputs(399) <= not((layer8_outputs(616)) xor (layer8_outputs(2188)));
    outputs(400) <= not((layer8_outputs(2450)) xor (layer8_outputs(2936)));
    outputs(401) <= not(layer8_outputs(3432));
    outputs(402) <= not((layer8_outputs(29)) or (layer8_outputs(1851)));
    outputs(403) <= not((layer8_outputs(4032)) or (layer8_outputs(541)));
    outputs(404) <= (layer8_outputs(2782)) xor (layer8_outputs(1867));
    outputs(405) <= (layer8_outputs(5038)) xor (layer8_outputs(2411));
    outputs(406) <= not(layer8_outputs(2416));
    outputs(407) <= layer8_outputs(921);
    outputs(408) <= not((layer8_outputs(3836)) or (layer8_outputs(3314)));
    outputs(409) <= not((layer8_outputs(1955)) xor (layer8_outputs(2479)));
    outputs(410) <= (layer8_outputs(4580)) xor (layer8_outputs(4651));
    outputs(411) <= not(layer8_outputs(12)) or (layer8_outputs(4722));
    outputs(412) <= not(layer8_outputs(4817));
    outputs(413) <= not(layer8_outputs(28));
    outputs(414) <= not(layer8_outputs(1063));
    outputs(415) <= not(layer8_outputs(4868));
    outputs(416) <= (layer8_outputs(4383)) xor (layer8_outputs(448));
    outputs(417) <= not((layer8_outputs(3858)) or (layer8_outputs(575)));
    outputs(418) <= layer8_outputs(2830);
    outputs(419) <= layer8_outputs(4094);
    outputs(420) <= not(layer8_outputs(3524));
    outputs(421) <= (layer8_outputs(238)) or (layer8_outputs(771));
    outputs(422) <= (layer8_outputs(3213)) xor (layer8_outputs(3494));
    outputs(423) <= layer8_outputs(451);
    outputs(424) <= not(layer8_outputs(2203));
    outputs(425) <= not((layer8_outputs(1966)) xor (layer8_outputs(4875)));
    outputs(426) <= (layer8_outputs(3089)) xor (layer8_outputs(792));
    outputs(427) <= not(layer8_outputs(3248));
    outputs(428) <= not((layer8_outputs(3339)) xor (layer8_outputs(1703)));
    outputs(429) <= not(layer8_outputs(2601)) or (layer8_outputs(2497));
    outputs(430) <= layer8_outputs(3009);
    outputs(431) <= (layer8_outputs(4797)) and not (layer8_outputs(1017));
    outputs(432) <= not(layer8_outputs(4189));
    outputs(433) <= not((layer8_outputs(1151)) xor (layer8_outputs(2158)));
    outputs(434) <= (layer8_outputs(2816)) and (layer8_outputs(2685));
    outputs(435) <= (layer8_outputs(2832)) and not (layer8_outputs(417));
    outputs(436) <= layer8_outputs(4984);
    outputs(437) <= not(layer8_outputs(1797));
    outputs(438) <= not((layer8_outputs(1788)) xor (layer8_outputs(903)));
    outputs(439) <= layer8_outputs(1527);
    outputs(440) <= not(layer8_outputs(3174)) or (layer8_outputs(2921));
    outputs(441) <= (layer8_outputs(2732)) xor (layer8_outputs(3572));
    outputs(442) <= layer8_outputs(4913);
    outputs(443) <= not((layer8_outputs(326)) xor (layer8_outputs(2414)));
    outputs(444) <= not(layer8_outputs(3773));
    outputs(445) <= not((layer8_outputs(331)) or (layer8_outputs(2553)));
    outputs(446) <= (layer8_outputs(3197)) and not (layer8_outputs(1776));
    outputs(447) <= (layer8_outputs(670)) xor (layer8_outputs(2911));
    outputs(448) <= (layer8_outputs(2943)) xor (layer8_outputs(4573));
    outputs(449) <= (layer8_outputs(4708)) xor (layer8_outputs(1148));
    outputs(450) <= (layer8_outputs(3196)) and not (layer8_outputs(781));
    outputs(451) <= (layer8_outputs(2755)) xor (layer8_outputs(4633));
    outputs(452) <= not(layer8_outputs(4345));
    outputs(453) <= layer8_outputs(2391);
    outputs(454) <= (layer8_outputs(1906)) xor (layer8_outputs(4884));
    outputs(455) <= layer8_outputs(3226);
    outputs(456) <= not(layer8_outputs(3565));
    outputs(457) <= not(layer8_outputs(4081));
    outputs(458) <= layer8_outputs(3951);
    outputs(459) <= not(layer8_outputs(1825));
    outputs(460) <= not((layer8_outputs(4011)) xor (layer8_outputs(2708)));
    outputs(461) <= layer8_outputs(2549);
    outputs(462) <= not((layer8_outputs(5040)) or (layer8_outputs(656)));
    outputs(463) <= (layer8_outputs(4921)) xor (layer8_outputs(4845));
    outputs(464) <= not((layer8_outputs(250)) xor (layer8_outputs(1465)));
    outputs(465) <= (layer8_outputs(4803)) xor (layer8_outputs(4172));
    outputs(466) <= not((layer8_outputs(83)) xor (layer8_outputs(4847)));
    outputs(467) <= not((layer8_outputs(716)) and (layer8_outputs(2776)));
    outputs(468) <= layer8_outputs(1052);
    outputs(469) <= (layer8_outputs(3513)) and not (layer8_outputs(2828));
    outputs(470) <= not((layer8_outputs(2863)) xor (layer8_outputs(4141)));
    outputs(471) <= not(layer8_outputs(2714));
    outputs(472) <= layer8_outputs(5003);
    outputs(473) <= layer8_outputs(1221);
    outputs(474) <= not((layer8_outputs(1147)) or (layer8_outputs(3824)));
    outputs(475) <= not(layer8_outputs(2695));
    outputs(476) <= not((layer8_outputs(3960)) xor (layer8_outputs(4937)));
    outputs(477) <= not((layer8_outputs(4576)) xor (layer8_outputs(2947)));
    outputs(478) <= not(layer8_outputs(4889));
    outputs(479) <= (layer8_outputs(3202)) and not (layer8_outputs(2564));
    outputs(480) <= not(layer8_outputs(2077));
    outputs(481) <= not(layer8_outputs(3585));
    outputs(482) <= not(layer8_outputs(81));
    outputs(483) <= layer8_outputs(4353);
    outputs(484) <= layer8_outputs(852);
    outputs(485) <= layer8_outputs(1630);
    outputs(486) <= not(layer8_outputs(2738));
    outputs(487) <= layer8_outputs(2641);
    outputs(488) <= not(layer8_outputs(2366));
    outputs(489) <= layer8_outputs(1075);
    outputs(490) <= not((layer8_outputs(2036)) xor (layer8_outputs(3193)));
    outputs(491) <= layer8_outputs(1870);
    outputs(492) <= (layer8_outputs(4314)) and not (layer8_outputs(4986));
    outputs(493) <= not(layer8_outputs(995));
    outputs(494) <= layer8_outputs(225);
    outputs(495) <= (layer8_outputs(1351)) xor (layer8_outputs(1699));
    outputs(496) <= (layer8_outputs(4221)) xor (layer8_outputs(1761));
    outputs(497) <= layer8_outputs(2819);
    outputs(498) <= (layer8_outputs(2163)) xor (layer8_outputs(3660));
    outputs(499) <= not((layer8_outputs(4738)) xor (layer8_outputs(2674)));
    outputs(500) <= not((layer8_outputs(3680)) xor (layer8_outputs(2752)));
    outputs(501) <= not(layer8_outputs(1438));
    outputs(502) <= not(layer8_outputs(2537));
    outputs(503) <= layer8_outputs(2631);
    outputs(504) <= not(layer8_outputs(886));
    outputs(505) <= not(layer8_outputs(1705));
    outputs(506) <= (layer8_outputs(929)) and not (layer8_outputs(400));
    outputs(507) <= not(layer8_outputs(3703));
    outputs(508) <= layer8_outputs(125);
    outputs(509) <= not(layer8_outputs(325));
    outputs(510) <= not(layer8_outputs(1830)) or (layer8_outputs(3632));
    outputs(511) <= not(layer8_outputs(4866));
    outputs(512) <= layer8_outputs(1947);
    outputs(513) <= not((layer8_outputs(819)) and (layer8_outputs(800)));
    outputs(514) <= (layer8_outputs(4352)) and not (layer8_outputs(2549));
    outputs(515) <= (layer8_outputs(1454)) and not (layer8_outputs(805));
    outputs(516) <= layer8_outputs(2043);
    outputs(517) <= not(layer8_outputs(4265));
    outputs(518) <= layer8_outputs(4346);
    outputs(519) <= not(layer8_outputs(3004)) or (layer8_outputs(3999));
    outputs(520) <= not((layer8_outputs(2647)) xor (layer8_outputs(2046)));
    outputs(521) <= not(layer8_outputs(3013));
    outputs(522) <= layer8_outputs(637);
    outputs(523) <= (layer8_outputs(3779)) and (layer8_outputs(1937));
    outputs(524) <= layer8_outputs(1903);
    outputs(525) <= layer8_outputs(2074);
    outputs(526) <= layer8_outputs(1339);
    outputs(527) <= not(layer8_outputs(1406));
    outputs(528) <= layer8_outputs(1998);
    outputs(529) <= not(layer8_outputs(843));
    outputs(530) <= not((layer8_outputs(2477)) xor (layer8_outputs(3988)));
    outputs(531) <= not(layer8_outputs(1975));
    outputs(532) <= not(layer8_outputs(4735));
    outputs(533) <= (layer8_outputs(1065)) xor (layer8_outputs(1539));
    outputs(534) <= not((layer8_outputs(1529)) or (layer8_outputs(3081)));
    outputs(535) <= not(layer8_outputs(431));
    outputs(536) <= (layer8_outputs(2491)) and not (layer8_outputs(4424));
    outputs(537) <= layer8_outputs(4328);
    outputs(538) <= (layer8_outputs(4073)) xor (layer8_outputs(2037));
    outputs(539) <= not((layer8_outputs(4540)) or (layer8_outputs(3890)));
    outputs(540) <= layer8_outputs(5017);
    outputs(541) <= not((layer8_outputs(2129)) or (layer8_outputs(2216)));
    outputs(542) <= layer8_outputs(232);
    outputs(543) <= (layer8_outputs(3016)) and (layer8_outputs(1439));
    outputs(544) <= layer8_outputs(3141);
    outputs(545) <= not(layer8_outputs(532));
    outputs(546) <= layer8_outputs(3993);
    outputs(547) <= not(layer8_outputs(807));
    outputs(548) <= not((layer8_outputs(3933)) xor (layer8_outputs(5001)));
    outputs(549) <= layer8_outputs(4965);
    outputs(550) <= not((layer8_outputs(1229)) xor (layer8_outputs(1529)));
    outputs(551) <= not((layer8_outputs(3814)) xor (layer8_outputs(3569)));
    outputs(552) <= not(layer8_outputs(1601));
    outputs(553) <= not(layer8_outputs(271));
    outputs(554) <= not(layer8_outputs(3558));
    outputs(555) <= not(layer8_outputs(1600));
    outputs(556) <= not((layer8_outputs(4499)) xor (layer8_outputs(904)));
    outputs(557) <= layer8_outputs(3398);
    outputs(558) <= (layer8_outputs(2291)) xor (layer8_outputs(4118));
    outputs(559) <= (layer8_outputs(4680)) and (layer8_outputs(74));
    outputs(560) <= not((layer8_outputs(1398)) xor (layer8_outputs(539)));
    outputs(561) <= not(layer8_outputs(405));
    outputs(562) <= layer8_outputs(2543);
    outputs(563) <= not(layer8_outputs(3911));
    outputs(564) <= (layer8_outputs(2941)) and not (layer8_outputs(4914));
    outputs(565) <= not(layer8_outputs(3967));
    outputs(566) <= layer8_outputs(200);
    outputs(567) <= not(layer8_outputs(1357));
    outputs(568) <= layer8_outputs(951);
    outputs(569) <= layer8_outputs(1395);
    outputs(570) <= layer8_outputs(1288);
    outputs(571) <= (layer8_outputs(4923)) and (layer8_outputs(2521));
    outputs(572) <= not((layer8_outputs(3843)) xor (layer8_outputs(4429)));
    outputs(573) <= not((layer8_outputs(3873)) xor (layer8_outputs(1784)));
    outputs(574) <= not(layer8_outputs(1517));
    outputs(575) <= not((layer8_outputs(4303)) or (layer8_outputs(2832)));
    outputs(576) <= (layer8_outputs(2720)) and not (layer8_outputs(2072));
    outputs(577) <= layer8_outputs(2370);
    outputs(578) <= not((layer8_outputs(1558)) xor (layer8_outputs(3200)));
    outputs(579) <= not((layer8_outputs(1632)) or (layer8_outputs(3934)));
    outputs(580) <= layer8_outputs(4120);
    outputs(581) <= not(layer8_outputs(2533));
    outputs(582) <= layer8_outputs(3499);
    outputs(583) <= (layer8_outputs(3730)) and not (layer8_outputs(1047));
    outputs(584) <= layer8_outputs(1964);
    outputs(585) <= layer8_outputs(1274);
    outputs(586) <= not(layer8_outputs(3356));
    outputs(587) <= not(layer8_outputs(3615));
    outputs(588) <= layer8_outputs(562);
    outputs(589) <= not(layer8_outputs(4895));
    outputs(590) <= layer8_outputs(1207);
    outputs(591) <= layer8_outputs(742);
    outputs(592) <= layer8_outputs(4788);
    outputs(593) <= layer8_outputs(960);
    outputs(594) <= layer8_outputs(1277);
    outputs(595) <= not((layer8_outputs(3463)) xor (layer8_outputs(112)));
    outputs(596) <= (layer8_outputs(4021)) and not (layer8_outputs(3418));
    outputs(597) <= layer8_outputs(490);
    outputs(598) <= (layer8_outputs(2556)) xor (layer8_outputs(4136));
    outputs(599) <= layer8_outputs(4812);
    outputs(600) <= layer8_outputs(2408);
    outputs(601) <= (layer8_outputs(1680)) xor (layer8_outputs(4382));
    outputs(602) <= not(layer8_outputs(2843)) or (layer8_outputs(2901));
    outputs(603) <= layer8_outputs(94);
    outputs(604) <= not((layer8_outputs(881)) xor (layer8_outputs(2798)));
    outputs(605) <= not(layer8_outputs(1383));
    outputs(606) <= layer8_outputs(3180);
    outputs(607) <= not(layer8_outputs(1050));
    outputs(608) <= layer8_outputs(1133);
    outputs(609) <= layer8_outputs(2231);
    outputs(610) <= not(layer8_outputs(4198));
    outputs(611) <= not(layer8_outputs(3718)) or (layer8_outputs(2759));
    outputs(612) <= (layer8_outputs(4610)) and not (layer8_outputs(2053));
    outputs(613) <= layer8_outputs(613);
    outputs(614) <= not(layer8_outputs(3613));
    outputs(615) <= layer8_outputs(1165);
    outputs(616) <= not((layer8_outputs(2963)) or (layer8_outputs(971)));
    outputs(617) <= layer8_outputs(1787);
    outputs(618) <= layer8_outputs(4941);
    outputs(619) <= layer8_outputs(3600);
    outputs(620) <= layer8_outputs(3602);
    outputs(621) <= (layer8_outputs(1890)) and (layer8_outputs(4232));
    outputs(622) <= not((layer8_outputs(2399)) xor (layer8_outputs(4315)));
    outputs(623) <= (layer8_outputs(3452)) xor (layer8_outputs(2680));
    outputs(624) <= not(layer8_outputs(3490));
    outputs(625) <= (layer8_outputs(3331)) xor (layer8_outputs(4267));
    outputs(626) <= not(layer8_outputs(310));
    outputs(627) <= (layer8_outputs(2019)) and (layer8_outputs(1925));
    outputs(628) <= layer8_outputs(2121);
    outputs(629) <= (layer8_outputs(4373)) xor (layer8_outputs(4489));
    outputs(630) <= (layer8_outputs(145)) xor (layer8_outputs(2726));
    outputs(631) <= layer8_outputs(2199);
    outputs(632) <= layer8_outputs(1442);
    outputs(633) <= layer8_outputs(3298);
    outputs(634) <= layer8_outputs(3147);
    outputs(635) <= not(layer8_outputs(4544));
    outputs(636) <= (layer8_outputs(1627)) xor (layer8_outputs(2648));
    outputs(637) <= not(layer8_outputs(791));
    outputs(638) <= not(layer8_outputs(1632));
    outputs(639) <= layer8_outputs(2067);
    outputs(640) <= layer8_outputs(146);
    outputs(641) <= (layer8_outputs(3945)) and not (layer8_outputs(1532));
    outputs(642) <= not(layer8_outputs(3946));
    outputs(643) <= layer8_outputs(2455);
    outputs(644) <= layer8_outputs(1390);
    outputs(645) <= not(layer8_outputs(604));
    outputs(646) <= (layer8_outputs(3970)) and not (layer8_outputs(2353));
    outputs(647) <= not(layer8_outputs(540));
    outputs(648) <= layer8_outputs(1134);
    outputs(649) <= (layer8_outputs(3069)) and not (layer8_outputs(3927));
    outputs(650) <= not((layer8_outputs(4397)) or (layer8_outputs(3054)));
    outputs(651) <= layer8_outputs(5090);
    outputs(652) <= layer8_outputs(1511);
    outputs(653) <= layer8_outputs(230);
    outputs(654) <= layer8_outputs(5066);
    outputs(655) <= not(layer8_outputs(1201));
    outputs(656) <= layer8_outputs(2661);
    outputs(657) <= layer8_outputs(1826);
    outputs(658) <= layer8_outputs(3639);
    outputs(659) <= not(layer8_outputs(2493));
    outputs(660) <= layer8_outputs(2214);
    outputs(661) <= layer8_outputs(2697);
    outputs(662) <= layer8_outputs(4779);
    outputs(663) <= not((layer8_outputs(4259)) xor (layer8_outputs(4413)));
    outputs(664) <= layer8_outputs(1475);
    outputs(665) <= not(layer8_outputs(515));
    outputs(666) <= not((layer8_outputs(2375)) or (layer8_outputs(4821)));
    outputs(667) <= not(layer8_outputs(35));
    outputs(668) <= not((layer8_outputs(1513)) xor (layer8_outputs(3331)));
    outputs(669) <= layer8_outputs(2212);
    outputs(670) <= not((layer8_outputs(2707)) xor (layer8_outputs(1360)));
    outputs(671) <= (layer8_outputs(381)) and not (layer8_outputs(197));
    outputs(672) <= not(layer8_outputs(4900));
    outputs(673) <= not(layer8_outputs(1139));
    outputs(674) <= (layer8_outputs(1103)) and (layer8_outputs(1769));
    outputs(675) <= not((layer8_outputs(1645)) or (layer8_outputs(5015)));
    outputs(676) <= not(layer8_outputs(2421));
    outputs(677) <= not(layer8_outputs(3495));
    outputs(678) <= not(layer8_outputs(3638)) or (layer8_outputs(1053));
    outputs(679) <= (layer8_outputs(3709)) xor (layer8_outputs(3932));
    outputs(680) <= (layer8_outputs(215)) and (layer8_outputs(3781));
    outputs(681) <= (layer8_outputs(1904)) xor (layer8_outputs(3534));
    outputs(682) <= (layer8_outputs(4936)) xor (layer8_outputs(4166));
    outputs(683) <= layer8_outputs(4204);
    outputs(684) <= not(layer8_outputs(578));
    outputs(685) <= not(layer8_outputs(3790));
    outputs(686) <= layer8_outputs(4868);
    outputs(687) <= not(layer8_outputs(3894));
    outputs(688) <= (layer8_outputs(3916)) and not (layer8_outputs(453));
    outputs(689) <= (layer8_outputs(2573)) and not (layer8_outputs(4179));
    outputs(690) <= (layer8_outputs(1249)) xor (layer8_outputs(3451));
    outputs(691) <= layer8_outputs(3363);
    outputs(692) <= not((layer8_outputs(4362)) xor (layer8_outputs(1617)));
    outputs(693) <= layer8_outputs(1575);
    outputs(694) <= layer8_outputs(831);
    outputs(695) <= not(layer8_outputs(1347));
    outputs(696) <= not((layer8_outputs(4357)) xor (layer8_outputs(5011)));
    outputs(697) <= not((layer8_outputs(61)) xor (layer8_outputs(3548)));
    outputs(698) <= (layer8_outputs(2527)) and not (layer8_outputs(3489));
    outputs(699) <= layer8_outputs(4036);
    outputs(700) <= (layer8_outputs(582)) xor (layer8_outputs(346));
    outputs(701) <= not((layer8_outputs(3761)) xor (layer8_outputs(3707)));
    outputs(702) <= not(layer8_outputs(391));
    outputs(703) <= not(layer8_outputs(2500));
    outputs(704) <= layer8_outputs(3976);
    outputs(705) <= (layer8_outputs(165)) and not (layer8_outputs(1324));
    outputs(706) <= (layer8_outputs(967)) xor (layer8_outputs(3167));
    outputs(707) <= layer8_outputs(2467);
    outputs(708) <= (layer8_outputs(953)) and not (layer8_outputs(614));
    outputs(709) <= not((layer8_outputs(1557)) xor (layer8_outputs(3431)));
    outputs(710) <= layer8_outputs(1239);
    outputs(711) <= layer8_outputs(4014);
    outputs(712) <= layer8_outputs(3714);
    outputs(713) <= layer8_outputs(4445);
    outputs(714) <= layer8_outputs(378);
    outputs(715) <= not(layer8_outputs(2230));
    outputs(716) <= not((layer8_outputs(95)) xor (layer8_outputs(4700)));
    outputs(717) <= (layer8_outputs(1508)) and not (layer8_outputs(1391));
    outputs(718) <= not((layer8_outputs(2834)) xor (layer8_outputs(4765)));
    outputs(719) <= layer8_outputs(503);
    outputs(720) <= layer8_outputs(3859);
    outputs(721) <= not(layer8_outputs(3139));
    outputs(722) <= layer8_outputs(1717);
    outputs(723) <= (layer8_outputs(2670)) and not (layer8_outputs(2451));
    outputs(724) <= (layer8_outputs(2013)) xor (layer8_outputs(3066));
    outputs(725) <= not(layer8_outputs(2785));
    outputs(726) <= (layer8_outputs(3306)) and (layer8_outputs(855));
    outputs(727) <= not(layer8_outputs(1765));
    outputs(728) <= (layer8_outputs(4722)) xor (layer8_outputs(2437));
    outputs(729) <= layer8_outputs(1479);
    outputs(730) <= (layer8_outputs(1533)) and not (layer8_outputs(205));
    outputs(731) <= not((layer8_outputs(2245)) xor (layer8_outputs(3492)));
    outputs(732) <= (layer8_outputs(3205)) and not (layer8_outputs(950));
    outputs(733) <= not(layer8_outputs(1519));
    outputs(734) <= layer8_outputs(4361);
    outputs(735) <= (layer8_outputs(1169)) and (layer8_outputs(3370));
    outputs(736) <= (layer8_outputs(3676)) and (layer8_outputs(4074));
    outputs(737) <= layer8_outputs(3874);
    outputs(738) <= not((layer8_outputs(4490)) xor (layer8_outputs(710)));
    outputs(739) <= (layer8_outputs(3967)) and (layer8_outputs(3947));
    outputs(740) <= layer8_outputs(4472);
    outputs(741) <= not((layer8_outputs(3781)) xor (layer8_outputs(1426)));
    outputs(742) <= not((layer8_outputs(4266)) or (layer8_outputs(1823)));
    outputs(743) <= (layer8_outputs(1141)) and not (layer8_outputs(3161));
    outputs(744) <= not(layer8_outputs(3690)) or (layer8_outputs(5047));
    outputs(745) <= not(layer8_outputs(667));
    outputs(746) <= not(layer8_outputs(4272));
    outputs(747) <= (layer8_outputs(2678)) xor (layer8_outputs(4442));
    outputs(748) <= (layer8_outputs(2793)) xor (layer8_outputs(1886));
    outputs(749) <= not(layer8_outputs(3856));
    outputs(750) <= not(layer8_outputs(1265));
    outputs(751) <= not(layer8_outputs(4235));
    outputs(752) <= not(layer8_outputs(4045));
    outputs(753) <= layer8_outputs(4165);
    outputs(754) <= layer8_outputs(240);
    outputs(755) <= not(layer8_outputs(3407));
    outputs(756) <= not(layer8_outputs(3385)) or (layer8_outputs(3562));
    outputs(757) <= not(layer8_outputs(1138));
    outputs(758) <= layer8_outputs(4919);
    outputs(759) <= not(layer8_outputs(2838));
    outputs(760) <= not((layer8_outputs(1641)) xor (layer8_outputs(1842)));
    outputs(761) <= not((layer8_outputs(771)) or (layer8_outputs(2122)));
    outputs(762) <= (layer8_outputs(4525)) and (layer8_outputs(4142));
    outputs(763) <= layer8_outputs(1922);
    outputs(764) <= layer8_outputs(1121);
    outputs(765) <= not((layer8_outputs(2766)) or (layer8_outputs(4684)));
    outputs(766) <= not(layer8_outputs(3307));
    outputs(767) <= (layer8_outputs(1679)) and not (layer8_outputs(2905));
    outputs(768) <= (layer8_outputs(4350)) xor (layer8_outputs(1701));
    outputs(769) <= not(layer8_outputs(2693));
    outputs(770) <= layer8_outputs(1154);
    outputs(771) <= (layer8_outputs(3271)) xor (layer8_outputs(5003));
    outputs(772) <= not(layer8_outputs(808));
    outputs(773) <= layer8_outputs(4461);
    outputs(774) <= not(layer8_outputs(2027));
    outputs(775) <= not(layer8_outputs(1142));
    outputs(776) <= (layer8_outputs(2085)) and not (layer8_outputs(2874));
    outputs(777) <= (layer8_outputs(2988)) and not (layer8_outputs(628));
    outputs(778) <= not(layer8_outputs(3121));
    outputs(779) <= (layer8_outputs(2252)) xor (layer8_outputs(5058));
    outputs(780) <= not((layer8_outputs(2322)) xor (layer8_outputs(2634)));
    outputs(781) <= (layer8_outputs(4677)) and not (layer8_outputs(3684));
    outputs(782) <= not((layer8_outputs(3381)) xor (layer8_outputs(21)));
    outputs(783) <= (layer8_outputs(80)) and not (layer8_outputs(491));
    outputs(784) <= (layer8_outputs(2015)) xor (layer8_outputs(4012));
    outputs(785) <= (layer8_outputs(1944)) and not (layer8_outputs(3953));
    outputs(786) <= not(layer8_outputs(4701));
    outputs(787) <= not(layer8_outputs(2156));
    outputs(788) <= not(layer8_outputs(4759));
    outputs(789) <= layer8_outputs(4831);
    outputs(790) <= (layer8_outputs(2350)) and not (layer8_outputs(389));
    outputs(791) <= layer8_outputs(4472);
    outputs(792) <= not(layer8_outputs(5013));
    outputs(793) <= (layer8_outputs(4925)) xor (layer8_outputs(2441));
    outputs(794) <= not(layer8_outputs(3173)) or (layer8_outputs(4876));
    outputs(795) <= layer8_outputs(1235);
    outputs(796) <= (layer8_outputs(4609)) xor (layer8_outputs(4268));
    outputs(797) <= not(layer8_outputs(2942));
    outputs(798) <= (layer8_outputs(1197)) xor (layer8_outputs(3784));
    outputs(799) <= (layer8_outputs(2054)) and not (layer8_outputs(3791));
    outputs(800) <= layer8_outputs(309);
    outputs(801) <= (layer8_outputs(900)) and not (layer8_outputs(3806));
    outputs(802) <= (layer8_outputs(4415)) xor (layer8_outputs(383));
    outputs(803) <= (layer8_outputs(2040)) and (layer8_outputs(217));
    outputs(804) <= (layer8_outputs(1633)) and not (layer8_outputs(2498));
    outputs(805) <= (layer8_outputs(1728)) xor (layer8_outputs(133));
    outputs(806) <= not(layer8_outputs(1543));
    outputs(807) <= layer8_outputs(1637);
    outputs(808) <= (layer8_outputs(1840)) xor (layer8_outputs(2342));
    outputs(809) <= not((layer8_outputs(3383)) or (layer8_outputs(18)));
    outputs(810) <= layer8_outputs(3581);
    outputs(811) <= not((layer8_outputs(2683)) or (layer8_outputs(2173)));
    outputs(812) <= not((layer8_outputs(4560)) xor (layer8_outputs(2194)));
    outputs(813) <= not((layer8_outputs(1199)) xor (layer8_outputs(2421)));
    outputs(814) <= not(layer8_outputs(239));
    outputs(815) <= layer8_outputs(688);
    outputs(816) <= layer8_outputs(2459);
    outputs(817) <= not((layer8_outputs(2943)) xor (layer8_outputs(3457)));
    outputs(818) <= not((layer8_outputs(3682)) or (layer8_outputs(42)));
    outputs(819) <= not(layer8_outputs(3708)) or (layer8_outputs(104));
    outputs(820) <= not((layer8_outputs(1931)) or (layer8_outputs(2177)));
    outputs(821) <= (layer8_outputs(3496)) and (layer8_outputs(547));
    outputs(822) <= layer8_outputs(3227);
    outputs(823) <= not(layer8_outputs(592)) or (layer8_outputs(2187));
    outputs(824) <= layer8_outputs(3793);
    outputs(825) <= (layer8_outputs(2318)) xor (layer8_outputs(16));
    outputs(826) <= layer8_outputs(1893);
    outputs(827) <= layer8_outputs(146);
    outputs(828) <= not(layer8_outputs(1273));
    outputs(829) <= not(layer8_outputs(540));
    outputs(830) <= not(layer8_outputs(2694));
    outputs(831) <= not(layer8_outputs(5110));
    outputs(832) <= (layer8_outputs(3224)) xor (layer8_outputs(3681));
    outputs(833) <= (layer8_outputs(1906)) and (layer8_outputs(1785));
    outputs(834) <= not((layer8_outputs(988)) xor (layer8_outputs(1468)));
    outputs(835) <= not(layer8_outputs(3729));
    outputs(836) <= not(layer8_outputs(3355));
    outputs(837) <= (layer8_outputs(3567)) and not (layer8_outputs(1889));
    outputs(838) <= (layer8_outputs(1851)) and (layer8_outputs(329));
    outputs(839) <= not(layer8_outputs(4273));
    outputs(840) <= (layer8_outputs(3458)) xor (layer8_outputs(1546));
    outputs(841) <= layer8_outputs(236);
    outputs(842) <= not((layer8_outputs(399)) or (layer8_outputs(1047)));
    outputs(843) <= (layer8_outputs(1079)) and (layer8_outputs(3441));
    outputs(844) <= (layer8_outputs(4835)) or (layer8_outputs(102));
    outputs(845) <= not((layer8_outputs(1284)) xor (layer8_outputs(4947)));
    outputs(846) <= layer8_outputs(4516);
    outputs(847) <= layer8_outputs(2956);
    outputs(848) <= not((layer8_outputs(2427)) or (layer8_outputs(4402)));
    outputs(849) <= layer8_outputs(2719);
    outputs(850) <= not(layer8_outputs(3310));
    outputs(851) <= (layer8_outputs(536)) xor (layer8_outputs(5053));
    outputs(852) <= (layer8_outputs(2115)) xor (layer8_outputs(2395));
    outputs(853) <= not((layer8_outputs(3502)) xor (layer8_outputs(869)));
    outputs(854) <= not((layer8_outputs(198)) xor (layer8_outputs(4665)));
    outputs(855) <= (layer8_outputs(1345)) and (layer8_outputs(1110));
    outputs(856) <= not((layer8_outputs(788)) xor (layer8_outputs(3801)));
    outputs(857) <= not((layer8_outputs(1654)) or (layer8_outputs(242)));
    outputs(858) <= layer8_outputs(4238);
    outputs(859) <= (layer8_outputs(4768)) xor (layer8_outputs(4464));
    outputs(860) <= not(layer8_outputs(5005));
    outputs(861) <= (layer8_outputs(230)) xor (layer8_outputs(3516));
    outputs(862) <= (layer8_outputs(3466)) and (layer8_outputs(3648));
    outputs(863) <= layer8_outputs(4217);
    outputs(864) <= layer8_outputs(1136);
    outputs(865) <= layer8_outputs(253);
    outputs(866) <= (layer8_outputs(1155)) and not (layer8_outputs(3806));
    outputs(867) <= layer8_outputs(4083);
    outputs(868) <= layer8_outputs(1835);
    outputs(869) <= (layer8_outputs(533)) xor (layer8_outputs(317));
    outputs(870) <= layer8_outputs(3160);
    outputs(871) <= layer8_outputs(1395);
    outputs(872) <= not(layer8_outputs(2616));
    outputs(873) <= not((layer8_outputs(3500)) and (layer8_outputs(111)));
    outputs(874) <= (layer8_outputs(3979)) and not (layer8_outputs(4371));
    outputs(875) <= layer8_outputs(2125);
    outputs(876) <= not(layer8_outputs(1898));
    outputs(877) <= (layer8_outputs(584)) and (layer8_outputs(522));
    outputs(878) <= (layer8_outputs(376)) and (layer8_outputs(1713));
    outputs(879) <= not(layer8_outputs(5089));
    outputs(880) <= not(layer8_outputs(1228));
    outputs(881) <= not(layer8_outputs(4446));
    outputs(882) <= layer8_outputs(1150);
    outputs(883) <= layer8_outputs(3472);
    outputs(884) <= not(layer8_outputs(2694));
    outputs(885) <= (layer8_outputs(744)) and (layer8_outputs(2417));
    outputs(886) <= (layer8_outputs(3036)) and (layer8_outputs(2266));
    outputs(887) <= layer8_outputs(3907);
    outputs(888) <= not(layer8_outputs(1241));
    outputs(889) <= not(layer8_outputs(1293));
    outputs(890) <= not((layer8_outputs(3210)) or (layer8_outputs(62)));
    outputs(891) <= (layer8_outputs(4430)) and not (layer8_outputs(4161));
    outputs(892) <= layer8_outputs(4261);
    outputs(893) <= (layer8_outputs(123)) xor (layer8_outputs(1634));
    outputs(894) <= not((layer8_outputs(139)) xor (layer8_outputs(583)));
    outputs(895) <= (layer8_outputs(3885)) and not (layer8_outputs(1594));
    outputs(896) <= layer8_outputs(1779);
    outputs(897) <= (layer8_outputs(616)) or (layer8_outputs(2155));
    outputs(898) <= not(layer8_outputs(1994));
    outputs(899) <= not((layer8_outputs(322)) or (layer8_outputs(2159)));
    outputs(900) <= layer8_outputs(4082);
    outputs(901) <= not((layer8_outputs(3981)) xor (layer8_outputs(2125)));
    outputs(902) <= not(layer8_outputs(3197));
    outputs(903) <= layer8_outputs(82);
    outputs(904) <= not(layer8_outputs(911));
    outputs(905) <= layer8_outputs(2273);
    outputs(906) <= layer8_outputs(491);
    outputs(907) <= (layer8_outputs(851)) and not (layer8_outputs(1397));
    outputs(908) <= (layer8_outputs(212)) and (layer8_outputs(280));
    outputs(909) <= not(layer8_outputs(2916));
    outputs(910) <= layer8_outputs(2715);
    outputs(911) <= not((layer8_outputs(554)) xor (layer8_outputs(3013)));
    outputs(912) <= (layer8_outputs(1856)) xor (layer8_outputs(3286));
    outputs(913) <= (layer8_outputs(4218)) and not (layer8_outputs(1921));
    outputs(914) <= not((layer8_outputs(1498)) or (layer8_outputs(2463)));
    outputs(915) <= (layer8_outputs(4972)) and not (layer8_outputs(3437));
    outputs(916) <= not((layer8_outputs(4215)) xor (layer8_outputs(3384)));
    outputs(917) <= not((layer8_outputs(156)) and (layer8_outputs(863)));
    outputs(918) <= not((layer8_outputs(1844)) xor (layer8_outputs(2602)));
    outputs(919) <= not(layer8_outputs(3058));
    outputs(920) <= not(layer8_outputs(3583));
    outputs(921) <= not(layer8_outputs(3487));
    outputs(922) <= (layer8_outputs(523)) and (layer8_outputs(3305));
    outputs(923) <= (layer8_outputs(577)) and not (layer8_outputs(650));
    outputs(924) <= layer8_outputs(4917);
    outputs(925) <= layer8_outputs(3248);
    outputs(926) <= not((layer8_outputs(4281)) or (layer8_outputs(3335)));
    outputs(927) <= not(layer8_outputs(1374));
    outputs(928) <= not(layer8_outputs(505)) or (layer8_outputs(2314));
    outputs(929) <= not(layer8_outputs(785));
    outputs(930) <= not((layer8_outputs(683)) xor (layer8_outputs(1171)));
    outputs(931) <= layer8_outputs(315);
    outputs(932) <= layer8_outputs(184);
    outputs(933) <= not((layer8_outputs(3360)) xor (layer8_outputs(2115)));
    outputs(934) <= (layer8_outputs(1459)) and not (layer8_outputs(1331));
    outputs(935) <= not(layer8_outputs(803));
    outputs(936) <= (layer8_outputs(3701)) xor (layer8_outputs(2690));
    outputs(937) <= not(layer8_outputs(4926)) or (layer8_outputs(4822));
    outputs(938) <= (layer8_outputs(4906)) xor (layer8_outputs(51));
    outputs(939) <= layer8_outputs(1867);
    outputs(940) <= not((layer8_outputs(1611)) xor (layer8_outputs(2305)));
    outputs(941) <= layer8_outputs(775);
    outputs(942) <= layer8_outputs(1369);
    outputs(943) <= not((layer8_outputs(3500)) and (layer8_outputs(1600)));
    outputs(944) <= not(layer8_outputs(1973));
    outputs(945) <= not((layer8_outputs(1106)) or (layer8_outputs(4838)));
    outputs(946) <= not(layer8_outputs(53));
    outputs(947) <= layer8_outputs(259);
    outputs(948) <= not(layer8_outputs(3225));
    outputs(949) <= not(layer8_outputs(961));
    outputs(950) <= (layer8_outputs(1112)) xor (layer8_outputs(4923));
    outputs(951) <= not(layer8_outputs(604)) or (layer8_outputs(5077));
    outputs(952) <= layer8_outputs(4848);
    outputs(953) <= layer8_outputs(5084);
    outputs(954) <= (layer8_outputs(4673)) and (layer8_outputs(435));
    outputs(955) <= layer8_outputs(4549);
    outputs(956) <= (layer8_outputs(1774)) xor (layer8_outputs(4257));
    outputs(957) <= not((layer8_outputs(2660)) xor (layer8_outputs(3995)));
    outputs(958) <= not(layer8_outputs(1629));
    outputs(959) <= layer8_outputs(2572);
    outputs(960) <= layer8_outputs(2674);
    outputs(961) <= not(layer8_outputs(2968));
    outputs(962) <= '0';
    outputs(963) <= layer8_outputs(1572);
    outputs(964) <= layer8_outputs(2657);
    outputs(965) <= not(layer8_outputs(3811));
    outputs(966) <= not((layer8_outputs(1490)) xor (layer8_outputs(2054)));
    outputs(967) <= not((layer8_outputs(3809)) xor (layer8_outputs(963)));
    outputs(968) <= not(layer8_outputs(2545));
    outputs(969) <= (layer8_outputs(4790)) xor (layer8_outputs(2035));
    outputs(970) <= not((layer8_outputs(2834)) xor (layer8_outputs(3686)));
    outputs(971) <= not((layer8_outputs(3379)) xor (layer8_outputs(0)));
    outputs(972) <= (layer8_outputs(313)) xor (layer8_outputs(3053));
    outputs(973) <= '0';
    outputs(974) <= (layer8_outputs(4484)) and (layer8_outputs(134));
    outputs(975) <= not((layer8_outputs(3905)) xor (layer8_outputs(4452)));
    outputs(976) <= (layer8_outputs(445)) and not (layer8_outputs(411));
    outputs(977) <= layer8_outputs(4069);
    outputs(978) <= layer8_outputs(3388);
    outputs(979) <= not((layer8_outputs(612)) or (layer8_outputs(3246)));
    outputs(980) <= not((layer8_outputs(2548)) xor (layer8_outputs(4962)));
    outputs(981) <= not(layer8_outputs(650));
    outputs(982) <= not((layer8_outputs(700)) xor (layer8_outputs(2095)));
    outputs(983) <= '0';
    outputs(984) <= not((layer8_outputs(3884)) xor (layer8_outputs(129)));
    outputs(985) <= not(layer8_outputs(1081));
    outputs(986) <= (layer8_outputs(2268)) xor (layer8_outputs(61));
    outputs(987) <= not(layer8_outputs(2886));
    outputs(988) <= (layer8_outputs(1148)) and (layer8_outputs(1959));
    outputs(989) <= layer8_outputs(3284);
    outputs(990) <= not(layer8_outputs(3533));
    outputs(991) <= (layer8_outputs(1832)) xor (layer8_outputs(2516));
    outputs(992) <= not(layer8_outputs(785));
    outputs(993) <= layer8_outputs(4077);
    outputs(994) <= not((layer8_outputs(3189)) xor (layer8_outputs(578)));
    outputs(995) <= not(layer8_outputs(1405));
    outputs(996) <= not(layer8_outputs(1951));
    outputs(997) <= not((layer8_outputs(410)) or (layer8_outputs(5028)));
    outputs(998) <= layer8_outputs(2663);
    outputs(999) <= layer8_outputs(2004);
    outputs(1000) <= not(layer8_outputs(1355));
    outputs(1001) <= not((layer8_outputs(833)) or (layer8_outputs(1032)));
    outputs(1002) <= not(layer8_outputs(2284));
    outputs(1003) <= not(layer8_outputs(4043));
    outputs(1004) <= not(layer8_outputs(3073));
    outputs(1005) <= not(layer8_outputs(1854));
    outputs(1006) <= layer8_outputs(5039);
    outputs(1007) <= not(layer8_outputs(213));
    outputs(1008) <= (layer8_outputs(3337)) xor (layer8_outputs(3717));
    outputs(1009) <= not(layer8_outputs(1030));
    outputs(1010) <= (layer8_outputs(3201)) xor (layer8_outputs(5110));
    outputs(1011) <= layer8_outputs(845);
    outputs(1012) <= layer8_outputs(3679);
    outputs(1013) <= layer8_outputs(2256);
    outputs(1014) <= layer8_outputs(4089);
    outputs(1015) <= (layer8_outputs(3364)) xor (layer8_outputs(2843));
    outputs(1016) <= not(layer8_outputs(3318)) or (layer8_outputs(3738));
    outputs(1017) <= layer8_outputs(1095);
    outputs(1018) <= (layer8_outputs(1531)) and (layer8_outputs(2116));
    outputs(1019) <= not((layer8_outputs(4449)) or (layer8_outputs(4805)));
    outputs(1020) <= not((layer8_outputs(5055)) xor (layer8_outputs(4738)));
    outputs(1021) <= not(layer8_outputs(1686));
    outputs(1022) <= (layer8_outputs(3105)) xor (layer8_outputs(1399));
    outputs(1023) <= not(layer8_outputs(603));
    outputs(1024) <= (layer8_outputs(1177)) xor (layer8_outputs(768));
    outputs(1025) <= not(layer8_outputs(4047));
    outputs(1026) <= not(layer8_outputs(2043));
    outputs(1027) <= (layer8_outputs(2058)) and not (layer8_outputs(1641));
    outputs(1028) <= not(layer8_outputs(492));
    outputs(1029) <= layer8_outputs(1772);
    outputs(1030) <= (layer8_outputs(3968)) or (layer8_outputs(138));
    outputs(1031) <= layer8_outputs(3737);
    outputs(1032) <= (layer8_outputs(3626)) xor (layer8_outputs(1809));
    outputs(1033) <= (layer8_outputs(943)) and not (layer8_outputs(3230));
    outputs(1034) <= layer8_outputs(29);
    outputs(1035) <= not(layer8_outputs(3662));
    outputs(1036) <= (layer8_outputs(2074)) xor (layer8_outputs(2908));
    outputs(1037) <= layer8_outputs(4602);
    outputs(1038) <= layer8_outputs(1155);
    outputs(1039) <= not(layer8_outputs(318)) or (layer8_outputs(4211));
    outputs(1040) <= not(layer8_outputs(2302));
    outputs(1041) <= not((layer8_outputs(2297)) xor (layer8_outputs(1928)));
    outputs(1042) <= (layer8_outputs(712)) or (layer8_outputs(3290));
    outputs(1043) <= (layer8_outputs(769)) or (layer8_outputs(1411));
    outputs(1044) <= (layer8_outputs(4224)) xor (layer8_outputs(691));
    outputs(1045) <= not(layer8_outputs(990));
    outputs(1046) <= not(layer8_outputs(363));
    outputs(1047) <= layer8_outputs(1879);
    outputs(1048) <= not(layer8_outputs(4049));
    outputs(1049) <= layer8_outputs(1254);
    outputs(1050) <= not(layer8_outputs(96));
    outputs(1051) <= (layer8_outputs(3263)) xor (layer8_outputs(3826));
    outputs(1052) <= not(layer8_outputs(121));
    outputs(1053) <= layer8_outputs(3135);
    outputs(1054) <= (layer8_outputs(4426)) xor (layer8_outputs(1954));
    outputs(1055) <= layer8_outputs(2087);
    outputs(1056) <= not((layer8_outputs(3421)) or (layer8_outputs(4733)));
    outputs(1057) <= (layer8_outputs(3745)) xor (layer8_outputs(560));
    outputs(1058) <= not(layer8_outputs(2932));
    outputs(1059) <= (layer8_outputs(5092)) or (layer8_outputs(2201));
    outputs(1060) <= layer8_outputs(2663);
    outputs(1061) <= not((layer8_outputs(4596)) xor (layer8_outputs(947)));
    outputs(1062) <= layer8_outputs(1756);
    outputs(1063) <= not(layer8_outputs(120));
    outputs(1064) <= not((layer8_outputs(4244)) xor (layer8_outputs(4024)));
    outputs(1065) <= layer8_outputs(1876);
    outputs(1066) <= layer8_outputs(3426);
    outputs(1067) <= not(layer8_outputs(971));
    outputs(1068) <= not(layer8_outputs(4055));
    outputs(1069) <= not(layer8_outputs(513));
    outputs(1070) <= layer8_outputs(644);
    outputs(1071) <= not(layer8_outputs(4279)) or (layer8_outputs(4131));
    outputs(1072) <= not(layer8_outputs(163));
    outputs(1073) <= (layer8_outputs(2894)) xor (layer8_outputs(4967));
    outputs(1074) <= not(layer8_outputs(1974));
    outputs(1075) <= layer8_outputs(3962);
    outputs(1076) <= not(layer8_outputs(4535));
    outputs(1077) <= not((layer8_outputs(2113)) xor (layer8_outputs(3244)));
    outputs(1078) <= layer8_outputs(1817);
    outputs(1079) <= not(layer8_outputs(4651));
    outputs(1080) <= not(layer8_outputs(1128));
    outputs(1081) <= not(layer8_outputs(2351));
    outputs(1082) <= layer8_outputs(943);
    outputs(1083) <= layer8_outputs(2724);
    outputs(1084) <= layer8_outputs(3892);
    outputs(1085) <= layer8_outputs(1161);
    outputs(1086) <= (layer8_outputs(4655)) xor (layer8_outputs(2846));
    outputs(1087) <= not(layer8_outputs(1269));
    outputs(1088) <= not(layer8_outputs(246));
    outputs(1089) <= (layer8_outputs(3055)) and not (layer8_outputs(1230));
    outputs(1090) <= not(layer8_outputs(2463));
    outputs(1091) <= layer8_outputs(803);
    outputs(1092) <= not(layer8_outputs(4186));
    outputs(1093) <= not(layer8_outputs(91));
    outputs(1094) <= not(layer8_outputs(273));
    outputs(1095) <= layer8_outputs(58);
    outputs(1096) <= not(layer8_outputs(4406));
    outputs(1097) <= not(layer8_outputs(2387));
    outputs(1098) <= not((layer8_outputs(3417)) xor (layer8_outputs(5072)));
    outputs(1099) <= not((layer8_outputs(1539)) xor (layer8_outputs(4001)));
    outputs(1100) <= not(layer8_outputs(3780));
    outputs(1101) <= layer8_outputs(3356);
    outputs(1102) <= not((layer8_outputs(1629)) xor (layer8_outputs(702)));
    outputs(1103) <= not((layer8_outputs(1738)) xor (layer8_outputs(2594)));
    outputs(1104) <= (layer8_outputs(1666)) xor (layer8_outputs(974));
    outputs(1105) <= layer8_outputs(854);
    outputs(1106) <= layer8_outputs(2841);
    outputs(1107) <= layer8_outputs(4616);
    outputs(1108) <= layer8_outputs(1555);
    outputs(1109) <= not(layer8_outputs(3450));
    outputs(1110) <= not((layer8_outputs(3542)) or (layer8_outputs(395)));
    outputs(1111) <= (layer8_outputs(3261)) xor (layer8_outputs(227));
    outputs(1112) <= not(layer8_outputs(4246));
    outputs(1113) <= not((layer8_outputs(3702)) xor (layer8_outputs(599)));
    outputs(1114) <= not((layer8_outputs(3492)) xor (layer8_outputs(2104)));
    outputs(1115) <= not(layer8_outputs(3521)) or (layer8_outputs(2093));
    outputs(1116) <= layer8_outputs(2069);
    outputs(1117) <= (layer8_outputs(4993)) xor (layer8_outputs(1972));
    outputs(1118) <= not(layer8_outputs(657));
    outputs(1119) <= not((layer8_outputs(3820)) or (layer8_outputs(4469)));
    outputs(1120) <= layer8_outputs(5117);
    outputs(1121) <= not(layer8_outputs(2452));
    outputs(1122) <= layer8_outputs(261);
    outputs(1123) <= not((layer8_outputs(903)) xor (layer8_outputs(1894)));
    outputs(1124) <= not(layer8_outputs(3274));
    outputs(1125) <= not((layer8_outputs(2418)) xor (layer8_outputs(3270)));
    outputs(1126) <= not(layer8_outputs(4091));
    outputs(1127) <= layer8_outputs(3277);
    outputs(1128) <= not((layer8_outputs(4448)) xor (layer8_outputs(4792)));
    outputs(1129) <= not(layer8_outputs(4723));
    outputs(1130) <= layer8_outputs(2152);
    outputs(1131) <= layer8_outputs(4994);
    outputs(1132) <= not((layer8_outputs(3407)) xor (layer8_outputs(2565)));
    outputs(1133) <= not((layer8_outputs(284)) xor (layer8_outputs(2102)));
    outputs(1134) <= not(layer8_outputs(3474));
    outputs(1135) <= layer8_outputs(2081);
    outputs(1136) <= layer8_outputs(2092);
    outputs(1137) <= not(layer8_outputs(632)) or (layer8_outputs(3419));
    outputs(1138) <= layer8_outputs(2390);
    outputs(1139) <= not((layer8_outputs(2867)) xor (layer8_outputs(3184)));
    outputs(1140) <= layer8_outputs(4719);
    outputs(1141) <= (layer8_outputs(5010)) xor (layer8_outputs(4002));
    outputs(1142) <= layer8_outputs(3657);
    outputs(1143) <= not((layer8_outputs(698)) xor (layer8_outputs(5052)));
    outputs(1144) <= layer8_outputs(4337);
    outputs(1145) <= (layer8_outputs(4808)) xor (layer8_outputs(905));
    outputs(1146) <= not((layer8_outputs(759)) and (layer8_outputs(1521)));
    outputs(1147) <= not(layer8_outputs(1688));
    outputs(1148) <= not(layer8_outputs(3549)) or (layer8_outputs(4369));
    outputs(1149) <= layer8_outputs(4467);
    outputs(1150) <= layer8_outputs(1437);
    outputs(1151) <= layer8_outputs(2994);
    outputs(1152) <= not(layer8_outputs(5029));
    outputs(1153) <= (layer8_outputs(3467)) and not (layer8_outputs(952));
    outputs(1154) <= not(layer8_outputs(3268));
    outputs(1155) <= layer8_outputs(3848);
    outputs(1156) <= not(layer8_outputs(1961));
    outputs(1157) <= layer8_outputs(4149);
    outputs(1158) <= not((layer8_outputs(2985)) xor (layer8_outputs(229)));
    outputs(1159) <= not(layer8_outputs(23));
    outputs(1160) <= not(layer8_outputs(1512));
    outputs(1161) <= layer8_outputs(1003);
    outputs(1162) <= layer8_outputs(3157);
    outputs(1163) <= not(layer8_outputs(3470));
    outputs(1164) <= not(layer8_outputs(456));
    outputs(1165) <= not(layer8_outputs(3123));
    outputs(1166) <= layer8_outputs(2576);
    outputs(1167) <= layer8_outputs(49);
    outputs(1168) <= (layer8_outputs(5081)) xor (layer8_outputs(3743));
    outputs(1169) <= not(layer8_outputs(2710));
    outputs(1170) <= not(layer8_outputs(2539)) or (layer8_outputs(609));
    outputs(1171) <= not(layer8_outputs(3615));
    outputs(1172) <= (layer8_outputs(1691)) xor (layer8_outputs(2068));
    outputs(1173) <= not((layer8_outputs(1523)) xor (layer8_outputs(1533)));
    outputs(1174) <= not(layer8_outputs(786));
    outputs(1175) <= not(layer8_outputs(1530));
    outputs(1176) <= not(layer8_outputs(925));
    outputs(1177) <= not((layer8_outputs(956)) xor (layer8_outputs(888)));
    outputs(1178) <= layer8_outputs(3906);
    outputs(1179) <= (layer8_outputs(1846)) xor (layer8_outputs(3482));
    outputs(1180) <= not(layer8_outputs(5109));
    outputs(1181) <= not(layer8_outputs(2864));
    outputs(1182) <= not((layer8_outputs(3798)) xor (layer8_outputs(4294)));
    outputs(1183) <= (layer8_outputs(4635)) xor (layer8_outputs(1520));
    outputs(1184) <= not((layer8_outputs(287)) xor (layer8_outputs(1046)));
    outputs(1185) <= not(layer8_outputs(2757));
    outputs(1186) <= layer8_outputs(1985);
    outputs(1187) <= not((layer8_outputs(1452)) and (layer8_outputs(319)));
    outputs(1188) <= (layer8_outputs(2589)) and not (layer8_outputs(3483));
    outputs(1189) <= (layer8_outputs(4098)) xor (layer8_outputs(4775));
    outputs(1190) <= layer8_outputs(1999);
    outputs(1191) <= not(layer8_outputs(4033));
    outputs(1192) <= not(layer8_outputs(2736));
    outputs(1193) <= not(layer8_outputs(3132)) or (layer8_outputs(915));
    outputs(1194) <= (layer8_outputs(2941)) xor (layer8_outputs(5103));
    outputs(1195) <= not(layer8_outputs(4793));
    outputs(1196) <= not(layer8_outputs(868));
    outputs(1197) <= not(layer8_outputs(1388));
    outputs(1198) <= (layer8_outputs(2338)) or (layer8_outputs(2453));
    outputs(1199) <= not((layer8_outputs(1428)) and (layer8_outputs(1445)));
    outputs(1200) <= not((layer8_outputs(2328)) xor (layer8_outputs(4501)));
    outputs(1201) <= (layer8_outputs(3939)) xor (layer8_outputs(997));
    outputs(1202) <= layer8_outputs(155);
    outputs(1203) <= not(layer8_outputs(3262));
    outputs(1204) <= (layer8_outputs(3990)) xor (layer8_outputs(2274));
    outputs(1205) <= (layer8_outputs(1896)) and not (layer8_outputs(2578));
    outputs(1206) <= not((layer8_outputs(1670)) and (layer8_outputs(3015)));
    outputs(1207) <= not((layer8_outputs(892)) or (layer8_outputs(3279)));
    outputs(1208) <= (layer8_outputs(2317)) xor (layer8_outputs(4689));
    outputs(1209) <= not(layer8_outputs(1972));
    outputs(1210) <= layer8_outputs(3467);
    outputs(1211) <= not((layer8_outputs(2341)) or (layer8_outputs(4047)));
    outputs(1212) <= not((layer8_outputs(4127)) xor (layer8_outputs(3668)));
    outputs(1213) <= not(layer8_outputs(3924)) or (layer8_outputs(3000));
    outputs(1214) <= not(layer8_outputs(2779));
    outputs(1215) <= layer8_outputs(674);
    outputs(1216) <= layer8_outputs(3124);
    outputs(1217) <= (layer8_outputs(949)) xor (layer8_outputs(4323));
    outputs(1218) <= (layer8_outputs(2774)) xor (layer8_outputs(2255));
    outputs(1219) <= not((layer8_outputs(390)) xor (layer8_outputs(8)));
    outputs(1220) <= (layer8_outputs(1580)) xor (layer8_outputs(2419));
    outputs(1221) <= not((layer8_outputs(3041)) or (layer8_outputs(2962)));
    outputs(1222) <= not(layer8_outputs(1602));
    outputs(1223) <= not(layer8_outputs(687));
    outputs(1224) <= layer8_outputs(518);
    outputs(1225) <= not(layer8_outputs(2476));
    outputs(1226) <= (layer8_outputs(2677)) xor (layer8_outputs(4944));
    outputs(1227) <= layer8_outputs(1232);
    outputs(1228) <= not(layer8_outputs(2740));
    outputs(1229) <= not(layer8_outputs(142));
    outputs(1230) <= (layer8_outputs(1688)) xor (layer8_outputs(3359));
    outputs(1231) <= not((layer8_outputs(3583)) xor (layer8_outputs(638)));
    outputs(1232) <= not((layer8_outputs(4297)) or (layer8_outputs(3393)));
    outputs(1233) <= not(layer8_outputs(1708));
    outputs(1234) <= layer8_outputs(3788);
    outputs(1235) <= (layer8_outputs(517)) and not (layer8_outputs(1097));
    outputs(1236) <= (layer8_outputs(3212)) and (layer8_outputs(2193));
    outputs(1237) <= layer8_outputs(2795);
    outputs(1238) <= not((layer8_outputs(2489)) xor (layer8_outputs(2002)));
    outputs(1239) <= layer8_outputs(178);
    outputs(1240) <= (layer8_outputs(4269)) xor (layer8_outputs(920));
    outputs(1241) <= not((layer8_outputs(2706)) xor (layer8_outputs(4531)));
    outputs(1242) <= not(layer8_outputs(582));
    outputs(1243) <= not((layer8_outputs(4036)) xor (layer8_outputs(1579)));
    outputs(1244) <= layer8_outputs(5015);
    outputs(1245) <= not(layer8_outputs(2680)) or (layer8_outputs(4497));
    outputs(1246) <= (layer8_outputs(4427)) xor (layer8_outputs(1083));
    outputs(1247) <= (layer8_outputs(1659)) xor (layer8_outputs(3469));
    outputs(1248) <= layer8_outputs(1443);
    outputs(1249) <= layer8_outputs(5056);
    outputs(1250) <= not((layer8_outputs(1329)) and (layer8_outputs(3397)));
    outputs(1251) <= not((layer8_outputs(845)) xor (layer8_outputs(2938)));
    outputs(1252) <= not((layer8_outputs(4063)) xor (layer8_outputs(4949)));
    outputs(1253) <= not(layer8_outputs(3891));
    outputs(1254) <= layer8_outputs(4813);
    outputs(1255) <= layer8_outputs(4088);
    outputs(1256) <= not(layer8_outputs(3666)) or (layer8_outputs(2541));
    outputs(1257) <= (layer8_outputs(3243)) xor (layer8_outputs(4366));
    outputs(1258) <= layer8_outputs(4554);
    outputs(1259) <= not(layer8_outputs(4103));
    outputs(1260) <= not(layer8_outputs(4995));
    outputs(1261) <= not(layer8_outputs(3999)) or (layer8_outputs(4807));
    outputs(1262) <= layer8_outputs(2089);
    outputs(1263) <= layer8_outputs(191);
    outputs(1264) <= (layer8_outputs(4518)) xor (layer8_outputs(4413));
    outputs(1265) <= not((layer8_outputs(3257)) xor (layer8_outputs(4105)));
    outputs(1266) <= not(layer8_outputs(4706));
    outputs(1267) <= layer8_outputs(2246);
    outputs(1268) <= not((layer8_outputs(532)) and (layer8_outputs(4765)));
    outputs(1269) <= (layer8_outputs(1060)) xor (layer8_outputs(2853));
    outputs(1270) <= not(layer8_outputs(610));
    outputs(1271) <= (layer8_outputs(2756)) xor (layer8_outputs(4831));
    outputs(1272) <= (layer8_outputs(3754)) xor (layer8_outputs(881));
    outputs(1273) <= not(layer8_outputs(2995));
    outputs(1274) <= (layer8_outputs(3445)) xor (layer8_outputs(4985));
    outputs(1275) <= (layer8_outputs(3001)) xor (layer8_outputs(864));
    outputs(1276) <= layer8_outputs(3755);
    outputs(1277) <= not(layer8_outputs(728));
    outputs(1278) <= not(layer8_outputs(2167));
    outputs(1279) <= layer8_outputs(2881);
    outputs(1280) <= not(layer8_outputs(4740));
    outputs(1281) <= not((layer8_outputs(1820)) xor (layer8_outputs(2001)));
    outputs(1282) <= (layer8_outputs(2617)) xor (layer8_outputs(2808));
    outputs(1283) <= (layer8_outputs(4760)) or (layer8_outputs(4382));
    outputs(1284) <= not(layer8_outputs(2362));
    outputs(1285) <= not(layer8_outputs(1597));
    outputs(1286) <= not(layer8_outputs(693));
    outputs(1287) <= not((layer8_outputs(4337)) xor (layer8_outputs(3646)));
    outputs(1288) <= not((layer8_outputs(2604)) xor (layer8_outputs(111)));
    outputs(1289) <= (layer8_outputs(1036)) xor (layer8_outputs(3661));
    outputs(1290) <= not(layer8_outputs(2274));
    outputs(1291) <= not(layer8_outputs(4076));
    outputs(1292) <= not(layer8_outputs(4184));
    outputs(1293) <= not(layer8_outputs(4314));
    outputs(1294) <= not(layer8_outputs(291));
    outputs(1295) <= not(layer8_outputs(1708));
    outputs(1296) <= layer8_outputs(2017);
    outputs(1297) <= not(layer8_outputs(4500));
    outputs(1298) <= not((layer8_outputs(4604)) xor (layer8_outputs(1387)));
    outputs(1299) <= not(layer8_outputs(2574));
    outputs(1300) <= not(layer8_outputs(3382));
    outputs(1301) <= not(layer8_outputs(3203)) or (layer8_outputs(480));
    outputs(1302) <= not(layer8_outputs(794));
    outputs(1303) <= layer8_outputs(493);
    outputs(1304) <= (layer8_outputs(2278)) or (layer8_outputs(1045));
    outputs(1305) <= layer8_outputs(4202);
    outputs(1306) <= layer8_outputs(983);
    outputs(1307) <= (layer8_outputs(735)) xor (layer8_outputs(4087));
    outputs(1308) <= not((layer8_outputs(3452)) xor (layer8_outputs(4057)));
    outputs(1309) <= not(layer8_outputs(2619));
    outputs(1310) <= (layer8_outputs(3102)) and (layer8_outputs(4323));
    outputs(1311) <= (layer8_outputs(98)) xor (layer8_outputs(2974));
    outputs(1312) <= layer8_outputs(1796);
    outputs(1313) <= not((layer8_outputs(2623)) xor (layer8_outputs(1303)));
    outputs(1314) <= (layer8_outputs(1946)) and (layer8_outputs(1034));
    outputs(1315) <= layer8_outputs(568);
    outputs(1316) <= layer8_outputs(3587);
    outputs(1317) <= (layer8_outputs(2225)) xor (layer8_outputs(526));
    outputs(1318) <= (layer8_outputs(1685)) and not (layer8_outputs(4757));
    outputs(1319) <= not(layer8_outputs(1132)) or (layer8_outputs(231));
    outputs(1320) <= layer8_outputs(2138);
    outputs(1321) <= not(layer8_outputs(2722)) or (layer8_outputs(2175));
    outputs(1322) <= layer8_outputs(1202);
    outputs(1323) <= not((layer8_outputs(1610)) xor (layer8_outputs(3267)));
    outputs(1324) <= not(layer8_outputs(2571)) or (layer8_outputs(3329));
    outputs(1325) <= layer8_outputs(679);
    outputs(1326) <= not((layer8_outputs(4725)) xor (layer8_outputs(4870)));
    outputs(1327) <= not(layer8_outputs(4248));
    outputs(1328) <= (layer8_outputs(1470)) or (layer8_outputs(78));
    outputs(1329) <= layer8_outputs(749);
    outputs(1330) <= not(layer8_outputs(182));
    outputs(1331) <= (layer8_outputs(3695)) and not (layer8_outputs(473));
    outputs(1332) <= layer8_outputs(2606);
    outputs(1333) <= layer8_outputs(1330);
    outputs(1334) <= layer8_outputs(3828);
    outputs(1335) <= not((layer8_outputs(1212)) xor (layer8_outputs(4570)));
    outputs(1336) <= not(layer8_outputs(3196));
    outputs(1337) <= not(layer8_outputs(4598)) or (layer8_outputs(3497));
    outputs(1338) <= layer8_outputs(3792);
    outputs(1339) <= not(layer8_outputs(3391));
    outputs(1340) <= (layer8_outputs(432)) and not (layer8_outputs(2140));
    outputs(1341) <= not(layer8_outputs(867));
    outputs(1342) <= layer8_outputs(2891);
    outputs(1343) <= not((layer8_outputs(594)) or (layer8_outputs(4051)));
    outputs(1344) <= (layer8_outputs(3063)) and not (layer8_outputs(133));
    outputs(1345) <= not(layer8_outputs(5029));
    outputs(1346) <= layer8_outputs(2709);
    outputs(1347) <= not((layer8_outputs(4850)) and (layer8_outputs(2487)));
    outputs(1348) <= not(layer8_outputs(1246));
    outputs(1349) <= not(layer8_outputs(356));
    outputs(1350) <= not((layer8_outputs(2029)) xor (layer8_outputs(406)));
    outputs(1351) <= not(layer8_outputs(562));
    outputs(1352) <= layer8_outputs(3418);
    outputs(1353) <= (layer8_outputs(4558)) and not (layer8_outputs(4206));
    outputs(1354) <= (layer8_outputs(345)) xor (layer8_outputs(2119));
    outputs(1355) <= layer8_outputs(2530);
    outputs(1356) <= not(layer8_outputs(3322));
    outputs(1357) <= not(layer8_outputs(2473));
    outputs(1358) <= layer8_outputs(4309);
    outputs(1359) <= not(layer8_outputs(4372));
    outputs(1360) <= not(layer8_outputs(3502));
    outputs(1361) <= layer8_outputs(3175);
    outputs(1362) <= layer8_outputs(355);
    outputs(1363) <= (layer8_outputs(241)) xor (layer8_outputs(3296));
    outputs(1364) <= layer8_outputs(3771);
    outputs(1365) <= (layer8_outputs(2339)) or (layer8_outputs(1149));
    outputs(1366) <= not((layer8_outputs(1107)) xor (layer8_outputs(2000)));
    outputs(1367) <= layer8_outputs(4751);
    outputs(1368) <= not((layer8_outputs(1743)) or (layer8_outputs(100)));
    outputs(1369) <= not((layer8_outputs(4436)) xor (layer8_outputs(2147)));
    outputs(1370) <= layer8_outputs(484);
    outputs(1371) <= not((layer8_outputs(2428)) xor (layer8_outputs(4161)));
    outputs(1372) <= (layer8_outputs(937)) xor (layer8_outputs(159));
    outputs(1373) <= not(layer8_outputs(216));
    outputs(1374) <= layer8_outputs(4492);
    outputs(1375) <= (layer8_outputs(3508)) xor (layer8_outputs(2311));
    outputs(1376) <= not((layer8_outputs(955)) xor (layer8_outputs(4729)));
    outputs(1377) <= layer8_outputs(3871);
    outputs(1378) <= layer8_outputs(2697);
    outputs(1379) <= layer8_outputs(138);
    outputs(1380) <= layer8_outputs(1735);
    outputs(1381) <= (layer8_outputs(2165)) xor (layer8_outputs(3910));
    outputs(1382) <= layer8_outputs(2799);
    outputs(1383) <= layer8_outputs(218);
    outputs(1384) <= layer8_outputs(4429);
    outputs(1385) <= not(layer8_outputs(1420));
    outputs(1386) <= layer8_outputs(3843);
    outputs(1387) <= (layer8_outputs(858)) xor (layer8_outputs(2701));
    outputs(1388) <= not(layer8_outputs(5019)) or (layer8_outputs(1827));
    outputs(1389) <= layer8_outputs(3756);
    outputs(1390) <= (layer8_outputs(3091)) xor (layer8_outputs(3181));
    outputs(1391) <= not(layer8_outputs(4347));
    outputs(1392) <= layer8_outputs(1328);
    outputs(1393) <= layer8_outputs(1288);
    outputs(1394) <= layer8_outputs(2804);
    outputs(1395) <= layer8_outputs(2532);
    outputs(1396) <= (layer8_outputs(4524)) and (layer8_outputs(4640));
    outputs(1397) <= not(layer8_outputs(1821));
    outputs(1398) <= layer8_outputs(2500);
    outputs(1399) <= not((layer8_outputs(4742)) xor (layer8_outputs(2382)));
    outputs(1400) <= layer8_outputs(1650);
    outputs(1401) <= (layer8_outputs(2103)) or (layer8_outputs(2328));
    outputs(1402) <= not(layer8_outputs(3265));
    outputs(1403) <= not(layer8_outputs(4480));
    outputs(1404) <= not(layer8_outputs(489));
    outputs(1405) <= not(layer8_outputs(4262));
    outputs(1406) <= layer8_outputs(3955);
    outputs(1407) <= not(layer8_outputs(2609));
    outputs(1408) <= not(layer8_outputs(426));
    outputs(1409) <= (layer8_outputs(2809)) or (layer8_outputs(756));
    outputs(1410) <= not((layer8_outputs(2850)) xor (layer8_outputs(865)));
    outputs(1411) <= not((layer8_outputs(2084)) xor (layer8_outputs(8)));
    outputs(1412) <= layer8_outputs(2851);
    outputs(1413) <= not(layer8_outputs(1577));
    outputs(1414) <= layer8_outputs(1988);
    outputs(1415) <= not(layer8_outputs(625));
    outputs(1416) <= layer8_outputs(1684);
    outputs(1417) <= not(layer8_outputs(3119)) or (layer8_outputs(2186));
    outputs(1418) <= layer8_outputs(2413);
    outputs(1419) <= not((layer8_outputs(1213)) or (layer8_outputs(413)));
    outputs(1420) <= layer8_outputs(2509);
    outputs(1421) <= layer8_outputs(1051);
    outputs(1422) <= not(layer8_outputs(4264));
    outputs(1423) <= layer8_outputs(4198);
    outputs(1424) <= layer8_outputs(3744);
    outputs(1425) <= not(layer8_outputs(924));
    outputs(1426) <= (layer8_outputs(4764)) xor (layer8_outputs(1090));
    outputs(1427) <= layer8_outputs(127);
    outputs(1428) <= layer8_outputs(4452);
    outputs(1429) <= not(layer8_outputs(179));
    outputs(1430) <= layer8_outputs(506);
    outputs(1431) <= not((layer8_outputs(3960)) xor (layer8_outputs(497)));
    outputs(1432) <= not(layer8_outputs(1734)) or (layer8_outputs(795));
    outputs(1433) <= (layer8_outputs(2063)) xor (layer8_outputs(4996));
    outputs(1434) <= not(layer8_outputs(2200));
    outputs(1435) <= not((layer8_outputs(3332)) xor (layer8_outputs(3476)));
    outputs(1436) <= not(layer8_outputs(3930));
    outputs(1437) <= layer8_outputs(27);
    outputs(1438) <= not((layer8_outputs(4263)) xor (layer8_outputs(2578)));
    outputs(1439) <= not(layer8_outputs(424)) or (layer8_outputs(3914));
    outputs(1440) <= not(layer8_outputs(4754));
    outputs(1441) <= not(layer8_outputs(3699));
    outputs(1442) <= not(layer8_outputs(1975));
    outputs(1443) <= not(layer8_outputs(1084));
    outputs(1444) <= (layer8_outputs(2756)) xor (layer8_outputs(4344));
    outputs(1445) <= not(layer8_outputs(4773));
    outputs(1446) <= not((layer8_outputs(1042)) xor (layer8_outputs(2822)));
    outputs(1447) <= not(layer8_outputs(3257));
    outputs(1448) <= layer8_outputs(3221);
    outputs(1449) <= (layer8_outputs(196)) or (layer8_outputs(978));
    outputs(1450) <= layer8_outputs(2860);
    outputs(1451) <= not((layer8_outputs(4055)) and (layer8_outputs(3574)));
    outputs(1452) <= layer8_outputs(4418);
    outputs(1453) <= layer8_outputs(1927);
    outputs(1454) <= not((layer8_outputs(4615)) xor (layer8_outputs(4728)));
    outputs(1455) <= not(layer8_outputs(3762));
    outputs(1456) <= (layer8_outputs(2813)) and not (layer8_outputs(4711));
    outputs(1457) <= layer8_outputs(4975);
    outputs(1458) <= (layer8_outputs(2127)) xor (layer8_outputs(4127));
    outputs(1459) <= (layer8_outputs(423)) xor (layer8_outputs(3410));
    outputs(1460) <= not(layer8_outputs(3751));
    outputs(1461) <= not((layer8_outputs(2435)) xor (layer8_outputs(1993)));
    outputs(1462) <= (layer8_outputs(3426)) or (layer8_outputs(1222));
    outputs(1463) <= (layer8_outputs(4529)) xor (layer8_outputs(4154));
    outputs(1464) <= layer8_outputs(662);
    outputs(1465) <= (layer8_outputs(1014)) xor (layer8_outputs(2948));
    outputs(1466) <= (layer8_outputs(1392)) xor (layer8_outputs(637));
    outputs(1467) <= not((layer8_outputs(263)) xor (layer8_outputs(2213)));
    outputs(1468) <= (layer8_outputs(1611)) xor (layer8_outputs(2129));
    outputs(1469) <= layer8_outputs(2532);
    outputs(1470) <= (layer8_outputs(543)) xor (layer8_outputs(4474));
    outputs(1471) <= layer8_outputs(1258);
    outputs(1472) <= layer8_outputs(1986);
    outputs(1473) <= not(layer8_outputs(4163));
    outputs(1474) <= (layer8_outputs(2542)) xor (layer8_outputs(3796));
    outputs(1475) <= not(layer8_outputs(1253));
    outputs(1476) <= (layer8_outputs(4586)) xor (layer8_outputs(3177));
    outputs(1477) <= layer8_outputs(3655);
    outputs(1478) <= (layer8_outputs(3803)) and not (layer8_outputs(4833));
    outputs(1479) <= not((layer8_outputs(2683)) xor (layer8_outputs(2970)));
    outputs(1480) <= layer8_outputs(857);
    outputs(1481) <= layer8_outputs(2959);
    outputs(1482) <= layer8_outputs(4841);
    outputs(1483) <= (layer8_outputs(2)) xor (layer8_outputs(1451));
    outputs(1484) <= not(layer8_outputs(410));
    outputs(1485) <= layer8_outputs(1727);
    outputs(1486) <= not(layer8_outputs(4252)) or (layer8_outputs(682));
    outputs(1487) <= layer8_outputs(2530);
    outputs(1488) <= not((layer8_outputs(4987)) xor (layer8_outputs(814)));
    outputs(1489) <= layer8_outputs(4880);
    outputs(1490) <= not(layer8_outputs(4101));
    outputs(1491) <= not(layer8_outputs(4789));
    outputs(1492) <= not(layer8_outputs(951));
    outputs(1493) <= layer8_outputs(1483);
    outputs(1494) <= (layer8_outputs(4173)) xor (layer8_outputs(1324));
    outputs(1495) <= not(layer8_outputs(483));
    outputs(1496) <= (layer8_outputs(3797)) xor (layer8_outputs(1912));
    outputs(1497) <= (layer8_outputs(817)) and (layer8_outputs(4536));
    outputs(1498) <= not((layer8_outputs(4369)) xor (layer8_outputs(197)));
    outputs(1499) <= (layer8_outputs(504)) xor (layer8_outputs(3527));
    outputs(1500) <= layer8_outputs(4610);
    outputs(1501) <= not(layer8_outputs(319));
    outputs(1502) <= not((layer8_outputs(4023)) and (layer8_outputs(4493)));
    outputs(1503) <= (layer8_outputs(2111)) xor (layer8_outputs(2265));
    outputs(1504) <= not(layer8_outputs(76)) or (layer8_outputs(1078));
    outputs(1505) <= (layer8_outputs(2651)) and (layer8_outputs(2443));
    outputs(1506) <= layer8_outputs(4853);
    outputs(1507) <= not(layer8_outputs(3659));
    outputs(1508) <= layer8_outputs(2657);
    outputs(1509) <= (layer8_outputs(4177)) xor (layer8_outputs(2003));
    outputs(1510) <= layer8_outputs(3584);
    outputs(1511) <= not(layer8_outputs(4842));
    outputs(1512) <= not((layer8_outputs(2476)) xor (layer8_outputs(1272)));
    outputs(1513) <= layer8_outputs(1417);
    outputs(1514) <= layer8_outputs(63);
    outputs(1515) <= not(layer8_outputs(760));
    outputs(1516) <= (layer8_outputs(811)) xor (layer8_outputs(4379));
    outputs(1517) <= (layer8_outputs(4796)) xor (layer8_outputs(4108));
    outputs(1518) <= not(layer8_outputs(629));
    outputs(1519) <= not(layer8_outputs(1140));
    outputs(1520) <= layer8_outputs(2607);
    outputs(1521) <= (layer8_outputs(3389)) and not (layer8_outputs(4278));
    outputs(1522) <= layer8_outputs(2092);
    outputs(1523) <= layer8_outputs(4145);
    outputs(1524) <= (layer8_outputs(4109)) xor (layer8_outputs(4857));
    outputs(1525) <= not((layer8_outputs(598)) xor (layer8_outputs(3429)));
    outputs(1526) <= not(layer8_outputs(931));
    outputs(1527) <= not((layer8_outputs(1053)) xor (layer8_outputs(120)));
    outputs(1528) <= not((layer8_outputs(4688)) xor (layer8_outputs(4617)));
    outputs(1529) <= not(layer8_outputs(2817));
    outputs(1530) <= not(layer8_outputs(3368));
    outputs(1531) <= layer8_outputs(202);
    outputs(1532) <= not(layer8_outputs(2932));
    outputs(1533) <= layer8_outputs(4777);
    outputs(1534) <= layer8_outputs(5073);
    outputs(1535) <= not(layer8_outputs(2712));
    outputs(1536) <= not((layer8_outputs(2783)) xor (layer8_outputs(3641)));
    outputs(1537) <= layer8_outputs(4524);
    outputs(1538) <= (layer8_outputs(4639)) and not (layer8_outputs(3414));
    outputs(1539) <= not(layer8_outputs(1618));
    outputs(1540) <= not(layer8_outputs(856));
    outputs(1541) <= (layer8_outputs(4005)) and not (layer8_outputs(1326));
    outputs(1542) <= not((layer8_outputs(4496)) xor (layer8_outputs(3065)));
    outputs(1543) <= not((layer8_outputs(549)) xor (layer8_outputs(308)));
    outputs(1544) <= (layer8_outputs(2165)) xor (layer8_outputs(579));
    outputs(1545) <= not(layer8_outputs(3952));
    outputs(1546) <= not(layer8_outputs(934));
    outputs(1547) <= not(layer8_outputs(4343));
    outputs(1548) <= not(layer8_outputs(3040));
    outputs(1549) <= layer8_outputs(97);
    outputs(1550) <= (layer8_outputs(815)) xor (layer8_outputs(465));
    outputs(1551) <= (layer8_outputs(2238)) and not (layer8_outputs(3540));
    outputs(1552) <= layer8_outputs(5069);
    outputs(1553) <= not((layer8_outputs(4405)) xor (layer8_outputs(753)));
    outputs(1554) <= not(layer8_outputs(1448));
    outputs(1555) <= layer8_outputs(2895);
    outputs(1556) <= not(layer8_outputs(1698));
    outputs(1557) <= not(layer8_outputs(4744));
    outputs(1558) <= not(layer8_outputs(1260));
    outputs(1559) <= layer8_outputs(3120);
    outputs(1560) <= layer8_outputs(4692);
    outputs(1561) <= not((layer8_outputs(1555)) or (layer8_outputs(1322)));
    outputs(1562) <= layer8_outputs(58);
    outputs(1563) <= (layer8_outputs(4836)) xor (layer8_outputs(3415));
    outputs(1564) <= not(layer8_outputs(550));
    outputs(1565) <= not(layer8_outputs(1801));
    outputs(1566) <= not(layer8_outputs(2163)) or (layer8_outputs(3643));
    outputs(1567) <= (layer8_outputs(2425)) xor (layer8_outputs(2420));
    outputs(1568) <= (layer8_outputs(2162)) and not (layer8_outputs(4892));
    outputs(1569) <= layer8_outputs(825);
    outputs(1570) <= not(layer8_outputs(4426));
    outputs(1571) <= (layer8_outputs(940)) xor (layer8_outputs(5009));
    outputs(1572) <= (layer8_outputs(72)) xor (layer8_outputs(1818));
    outputs(1573) <= not((layer8_outputs(27)) xor (layer8_outputs(3129)));
    outputs(1574) <= (layer8_outputs(2080)) and (layer8_outputs(1104));
    outputs(1575) <= not(layer8_outputs(528));
    outputs(1576) <= (layer8_outputs(1613)) and not (layer8_outputs(1146));
    outputs(1577) <= (layer8_outputs(3522)) xor (layer8_outputs(358));
    outputs(1578) <= (layer8_outputs(4542)) xor (layer8_outputs(3209));
    outputs(1579) <= layer8_outputs(4366);
    outputs(1580) <= layer8_outputs(4801);
    outputs(1581) <= (layer8_outputs(4887)) xor (layer8_outputs(315));
    outputs(1582) <= (layer8_outputs(4125)) xor (layer8_outputs(1943));
    outputs(1583) <= not(layer8_outputs(2918)) or (layer8_outputs(1823));
    outputs(1584) <= layer8_outputs(899);
    outputs(1585) <= (layer8_outputs(2409)) and (layer8_outputs(2750));
    outputs(1586) <= not((layer8_outputs(144)) xor (layer8_outputs(1320)));
    outputs(1587) <= (layer8_outputs(537)) xor (layer8_outputs(701));
    outputs(1588) <= layer8_outputs(3986);
    outputs(1589) <= not(layer8_outputs(1810));
    outputs(1590) <= not(layer8_outputs(751));
    outputs(1591) <= not(layer8_outputs(301));
    outputs(1592) <= (layer8_outputs(1504)) xor (layer8_outputs(4939));
    outputs(1593) <= not(layer8_outputs(4865));
    outputs(1594) <= layer8_outputs(4834);
    outputs(1595) <= not((layer8_outputs(367)) xor (layer8_outputs(3506)));
    outputs(1596) <= (layer8_outputs(2149)) and not (layer8_outputs(4380));
    outputs(1597) <= not((layer8_outputs(3634)) xor (layer8_outputs(3478)));
    outputs(1598) <= (layer8_outputs(4022)) xor (layer8_outputs(2809));
    outputs(1599) <= not(layer8_outputs(3592)) or (layer8_outputs(2075));
    outputs(1600) <= not(layer8_outputs(3531));
    outputs(1601) <= layer8_outputs(2305);
    outputs(1602) <= (layer8_outputs(297)) xor (layer8_outputs(4332));
    outputs(1603) <= layer8_outputs(53);
    outputs(1604) <= not((layer8_outputs(4324)) or (layer8_outputs(572)));
    outputs(1605) <= (layer8_outputs(4879)) xor (layer8_outputs(1642));
    outputs(1606) <= not(layer8_outputs(1482));
    outputs(1607) <= (layer8_outputs(2792)) and not (layer8_outputs(3312));
    outputs(1608) <= not(layer8_outputs(2307));
    outputs(1609) <= layer8_outputs(2402);
    outputs(1610) <= (layer8_outputs(2472)) or (layer8_outputs(2924));
    outputs(1611) <= not(layer8_outputs(4933));
    outputs(1612) <= (layer8_outputs(661)) xor (layer8_outputs(826));
    outputs(1613) <= layer8_outputs(5024);
    outputs(1614) <= not(layer8_outputs(2825));
    outputs(1615) <= layer8_outputs(1204);
    outputs(1616) <= (layer8_outputs(1290)) xor (layer8_outputs(725));
    outputs(1617) <= layer8_outputs(2171);
    outputs(1618) <= layer8_outputs(4257);
    outputs(1619) <= (layer8_outputs(3487)) and (layer8_outputs(2397));
    outputs(1620) <= layer8_outputs(3440);
    outputs(1621) <= not((layer8_outputs(3731)) xor (layer8_outputs(4810)));
    outputs(1622) <= not(layer8_outputs(2589));
    outputs(1623) <= not((layer8_outputs(3910)) or (layer8_outputs(2056)));
    outputs(1624) <= layer8_outputs(3101);
    outputs(1625) <= (layer8_outputs(2386)) xor (layer8_outputs(247));
    outputs(1626) <= not(layer8_outputs(2183));
    outputs(1627) <= layer8_outputs(2575);
    outputs(1628) <= layer8_outputs(5090);
    outputs(1629) <= (layer8_outputs(1631)) or (layer8_outputs(5063));
    outputs(1630) <= layer8_outputs(2446);
    outputs(1631) <= not((layer8_outputs(2966)) xor (layer8_outputs(1837)));
    outputs(1632) <= not(layer8_outputs(118));
    outputs(1633) <= (layer8_outputs(1205)) and not (layer8_outputs(385));
    outputs(1634) <= not(layer8_outputs(1991));
    outputs(1635) <= not((layer8_outputs(3516)) xor (layer8_outputs(1956)));
    outputs(1636) <= (layer8_outputs(5073)) and (layer8_outputs(493));
    outputs(1637) <= layer8_outputs(687);
    outputs(1638) <= layer8_outputs(3256);
    outputs(1639) <= not(layer8_outputs(2721));
    outputs(1640) <= layer8_outputs(4278);
    outputs(1641) <= not(layer8_outputs(5078));
    outputs(1642) <= layer8_outputs(4969);
    outputs(1643) <= not((layer8_outputs(3997)) xor (layer8_outputs(4003)));
    outputs(1644) <= (layer8_outputs(4007)) xor (layer8_outputs(774));
    outputs(1645) <= not(layer8_outputs(2513));
    outputs(1646) <= not(layer8_outputs(3272)) or (layer8_outputs(810));
    outputs(1647) <= not(layer8_outputs(2226));
    outputs(1648) <= layer8_outputs(3792);
    outputs(1649) <= not(layer8_outputs(2652));
    outputs(1650) <= not(layer8_outputs(1934));
    outputs(1651) <= not((layer8_outputs(1481)) xor (layer8_outputs(1696)));
    outputs(1652) <= layer8_outputs(712);
    outputs(1653) <= not((layer8_outputs(4643)) xor (layer8_outputs(433)));
    outputs(1654) <= not(layer8_outputs(3710));
    outputs(1655) <= not(layer8_outputs(304)) or (layer8_outputs(1981));
    outputs(1656) <= layer8_outputs(3128);
    outputs(1657) <= not((layer8_outputs(2325)) or (layer8_outputs(665)));
    outputs(1658) <= layer8_outputs(2788);
    outputs(1659) <= not(layer8_outputs(1433));
    outputs(1660) <= (layer8_outputs(1005)) and (layer8_outputs(4574));
    outputs(1661) <= (layer8_outputs(2022)) or (layer8_outputs(2450));
    outputs(1662) <= layer8_outputs(4253);
    outputs(1663) <= (layer8_outputs(4991)) or (layer8_outputs(1718));
    outputs(1664) <= layer8_outputs(1289);
    outputs(1665) <= not((layer8_outputs(1726)) xor (layer8_outputs(1736)));
    outputs(1666) <= layer8_outputs(420);
    outputs(1667) <= layer8_outputs(2639);
    outputs(1668) <= (layer8_outputs(262)) and not (layer8_outputs(449));
    outputs(1669) <= layer8_outputs(3928);
    outputs(1670) <= not(layer8_outputs(1862));
    outputs(1671) <= not((layer8_outputs(4254)) xor (layer8_outputs(1932)));
    outputs(1672) <= layer8_outputs(2773);
    outputs(1673) <= layer8_outputs(3559);
    outputs(1674) <= layer8_outputs(2372);
    outputs(1675) <= layer8_outputs(4028);
    outputs(1676) <= (layer8_outputs(939)) and (layer8_outputs(860));
    outputs(1677) <= not(layer8_outputs(2344));
    outputs(1678) <= not(layer8_outputs(2662));
    outputs(1679) <= not(layer8_outputs(2433));
    outputs(1680) <= not(layer8_outputs(574));
    outputs(1681) <= not(layer8_outputs(310));
    outputs(1682) <= not(layer8_outputs(681));
    outputs(1683) <= (layer8_outputs(185)) xor (layer8_outputs(171));
    outputs(1684) <= not(layer8_outputs(2219));
    outputs(1685) <= layer8_outputs(4450);
    outputs(1686) <= layer8_outputs(2661);
    outputs(1687) <= not((layer8_outputs(1754)) or (layer8_outputs(4922)));
    outputs(1688) <= not((layer8_outputs(3877)) xor (layer8_outputs(3395)));
    outputs(1689) <= not(layer8_outputs(1240));
    outputs(1690) <= layer8_outputs(5036);
    outputs(1691) <= layer8_outputs(4027);
    outputs(1692) <= not(layer8_outputs(3974));
    outputs(1693) <= not(layer8_outputs(4422));
    outputs(1694) <= not((layer8_outputs(2974)) or (layer8_outputs(480)));
    outputs(1695) <= not((layer8_outputs(4318)) xor (layer8_outputs(2150)));
    outputs(1696) <= layer8_outputs(1809);
    outputs(1697) <= not(layer8_outputs(3282));
    outputs(1698) <= not((layer8_outputs(3927)) xor (layer8_outputs(2447)));
    outputs(1699) <= (layer8_outputs(3891)) and not (layer8_outputs(4907));
    outputs(1700) <= layer8_outputs(1613);
    outputs(1701) <= (layer8_outputs(3415)) xor (layer8_outputs(519));
    outputs(1702) <= not(layer8_outputs(2899));
    outputs(1703) <= not((layer8_outputs(1472)) and (layer8_outputs(2970)));
    outputs(1704) <= not(layer8_outputs(599));
    outputs(1705) <= (layer8_outputs(4393)) and not (layer8_outputs(4686));
    outputs(1706) <= (layer8_outputs(4830)) xor (layer8_outputs(2783));
    outputs(1707) <= not(layer8_outputs(2249));
    outputs(1708) <= (layer8_outputs(914)) and not (layer8_outputs(1458));
    outputs(1709) <= (layer8_outputs(4639)) and not (layer8_outputs(4285));
    outputs(1710) <= layer8_outputs(2086);
    outputs(1711) <= layer8_outputs(467);
    outputs(1712) <= layer8_outputs(4241);
    outputs(1713) <= layer8_outputs(2837);
    outputs(1714) <= not(layer8_outputs(443));
    outputs(1715) <= not(layer8_outputs(303));
    outputs(1716) <= layer8_outputs(3103);
    outputs(1717) <= not(layer8_outputs(4558));
    outputs(1718) <= not((layer8_outputs(2280)) xor (layer8_outputs(1560)));
    outputs(1719) <= (layer8_outputs(3777)) and (layer8_outputs(2444));
    outputs(1720) <= not((layer8_outputs(4729)) xor (layer8_outputs(2885)));
    outputs(1721) <= not(layer8_outputs(1135));
    outputs(1722) <= not((layer8_outputs(4902)) or (layer8_outputs(2232)));
    outputs(1723) <= not(layer8_outputs(2502));
    outputs(1724) <= (layer8_outputs(3060)) xor (layer8_outputs(490));
    outputs(1725) <= (layer8_outputs(553)) and (layer8_outputs(3120));
    outputs(1726) <= layer8_outputs(2023);
    outputs(1727) <= (layer8_outputs(4752)) and not (layer8_outputs(3252));
    outputs(1728) <= not(layer8_outputs(3303));
    outputs(1729) <= (layer8_outputs(3157)) and not (layer8_outputs(4340));
    outputs(1730) <= not((layer8_outputs(4478)) xor (layer8_outputs(730)));
    outputs(1731) <= not(layer8_outputs(4319));
    outputs(1732) <= not((layer8_outputs(4534)) or (layer8_outputs(4983)));
    outputs(1733) <= not(layer8_outputs(1174));
    outputs(1734) <= layer8_outputs(3439);
    outputs(1735) <= (layer8_outputs(1001)) and not (layer8_outputs(906));
    outputs(1736) <= not((layer8_outputs(2659)) xor (layer8_outputs(2806)));
    outputs(1737) <= not((layer8_outputs(3594)) and (layer8_outputs(2381)));
    outputs(1738) <= layer8_outputs(2797);
    outputs(1739) <= layer8_outputs(941);
    outputs(1740) <= not(layer8_outputs(3682));
    outputs(1741) <= not((layer8_outputs(3974)) xor (layer8_outputs(2679)));
    outputs(1742) <= (layer8_outputs(1014)) xor (layer8_outputs(622));
    outputs(1743) <= not(layer8_outputs(3882));
    outputs(1744) <= (layer8_outputs(152)) xor (layer8_outputs(3047));
    outputs(1745) <= layer8_outputs(1378);
    outputs(1746) <= not(layer8_outputs(1835));
    outputs(1747) <= not((layer8_outputs(1683)) and (layer8_outputs(408)));
    outputs(1748) <= not(layer8_outputs(5079));
    outputs(1749) <= layer8_outputs(2150);
    outputs(1750) <= not(layer8_outputs(2520));
    outputs(1751) <= not(layer8_outputs(466));
    outputs(1752) <= not((layer8_outputs(3518)) xor (layer8_outputs(3669)));
    outputs(1753) <= layer8_outputs(1078);
    outputs(1754) <= layer8_outputs(4769);
    outputs(1755) <= (layer8_outputs(811)) and (layer8_outputs(2515));
    outputs(1756) <= not(layer8_outputs(2951));
    outputs(1757) <= not((layer8_outputs(3704)) or (layer8_outputs(529)));
    outputs(1758) <= not(layer8_outputs(4680));
    outputs(1759) <= layer8_outputs(472);
    outputs(1760) <= layer8_outputs(4696);
    outputs(1761) <= (layer8_outputs(3220)) and (layer8_outputs(981));
    outputs(1762) <= layer8_outputs(4099);
    outputs(1763) <= not(layer8_outputs(3258));
    outputs(1764) <= layer8_outputs(3417);
    outputs(1765) <= not(layer8_outputs(2557));
    outputs(1766) <= not(layer8_outputs(2064));
    outputs(1767) <= layer8_outputs(1410);
    outputs(1768) <= layer8_outputs(2205);
    outputs(1769) <= not((layer8_outputs(708)) xor (layer8_outputs(3353)));
    outputs(1770) <= not((layer8_outputs(4003)) or (layer8_outputs(2052)));
    outputs(1771) <= (layer8_outputs(203)) xor (layer8_outputs(2641));
    outputs(1772) <= not(layer8_outputs(1494));
    outputs(1773) <= not((layer8_outputs(4086)) xor (layer8_outputs(4766)));
    outputs(1774) <= not(layer8_outputs(4933));
    outputs(1775) <= not(layer8_outputs(4896));
    outputs(1776) <= layer8_outputs(452);
    outputs(1777) <= layer8_outputs(3062);
    outputs(1778) <= layer8_outputs(4063);
    outputs(1779) <= (layer8_outputs(2856)) or (layer8_outputs(4112));
    outputs(1780) <= layer8_outputs(3006);
    outputs(1781) <= layer8_outputs(2923);
    outputs(1782) <= layer8_outputs(3558);
    outputs(1783) <= not(layer8_outputs(2765));
    outputs(1784) <= layer8_outputs(1102);
    outputs(1785) <= layer8_outputs(2157);
    outputs(1786) <= not((layer8_outputs(4279)) or (layer8_outputs(2618)));
    outputs(1787) <= not((layer8_outputs(198)) xor (layer8_outputs(3559)));
    outputs(1788) <= not((layer8_outputs(3110)) or (layer8_outputs(930)));
    outputs(1789) <= (layer8_outputs(2179)) and not (layer8_outputs(3668));
    outputs(1790) <= layer8_outputs(4717);
    outputs(1791) <= not(layer8_outputs(4809));
    outputs(1792) <= layer8_outputs(5112);
    outputs(1793) <= not(layer8_outputs(2909));
    outputs(1794) <= not(layer8_outputs(4090));
    outputs(1795) <= not(layer8_outputs(4975));
    outputs(1796) <= not(layer8_outputs(2512));
    outputs(1797) <= layer8_outputs(1918);
    outputs(1798) <= layer8_outputs(1336);
    outputs(1799) <= not((layer8_outputs(1607)) xor (layer8_outputs(1981)));
    outputs(1800) <= not(layer8_outputs(4984)) or (layer8_outputs(2654));
    outputs(1801) <= not((layer8_outputs(789)) xor (layer8_outputs(3260)));
    outputs(1802) <= not((layer8_outputs(2360)) or (layer8_outputs(1226)));
    outputs(1803) <= not((layer8_outputs(377)) or (layer8_outputs(3758)));
    outputs(1804) <= not(layer8_outputs(4798));
    outputs(1805) <= (layer8_outputs(4111)) xor (layer8_outputs(4901));
    outputs(1806) <= not((layer8_outputs(940)) xor (layer8_outputs(3623)));
    outputs(1807) <= not((layer8_outputs(1368)) xor (layer8_outputs(852)));
    outputs(1808) <= layer8_outputs(1830);
    outputs(1809) <= layer8_outputs(1887);
    outputs(1810) <= (layer8_outputs(2189)) and not (layer8_outputs(5026));
    outputs(1811) <= not(layer8_outputs(4169));
    outputs(1812) <= layer8_outputs(2269);
    outputs(1813) <= layer8_outputs(2172);
    outputs(1814) <= not(layer8_outputs(2736));
    outputs(1815) <= (layer8_outputs(3206)) xor (layer8_outputs(3480));
    outputs(1816) <= not(layer8_outputs(3316));
    outputs(1817) <= layer8_outputs(783);
    outputs(1818) <= layer8_outputs(4033);
    outputs(1819) <= (layer8_outputs(2835)) or (layer8_outputs(2325));
    outputs(1820) <= not(layer8_outputs(5056));
    outputs(1821) <= layer8_outputs(3396);
    outputs(1822) <= not(layer8_outputs(1755));
    outputs(1823) <= not((layer8_outputs(783)) xor (layer8_outputs(1052)));
    outputs(1824) <= (layer8_outputs(2876)) xor (layer8_outputs(3348));
    outputs(1825) <= layer8_outputs(2001);
    outputs(1826) <= not(layer8_outputs(2137));
    outputs(1827) <= (layer8_outputs(1093)) and (layer8_outputs(1770));
    outputs(1828) <= layer8_outputs(3017);
    outputs(1829) <= not((layer8_outputs(4537)) xor (layer8_outputs(288)));
    outputs(1830) <= (layer8_outputs(973)) xor (layer8_outputs(1400));
    outputs(1831) <= (layer8_outputs(4194)) xor (layer8_outputs(1507));
    outputs(1832) <= layer8_outputs(900);
    outputs(1833) <= not(layer8_outputs(1550));
    outputs(1834) <= layer8_outputs(2016);
    outputs(1835) <= not((layer8_outputs(203)) xor (layer8_outputs(527)));
    outputs(1836) <= layer8_outputs(2912);
    outputs(1837) <= layer8_outputs(848);
    outputs(1838) <= (layer8_outputs(24)) and (layer8_outputs(3872));
    outputs(1839) <= not(layer8_outputs(1130));
    outputs(1840) <= not(layer8_outputs(2379));
    outputs(1841) <= (layer8_outputs(2929)) xor (layer8_outputs(155));
    outputs(1842) <= layer8_outputs(5022);
    outputs(1843) <= layer8_outputs(3391);
    outputs(1844) <= (layer8_outputs(2948)) xor (layer8_outputs(4899));
    outputs(1845) <= (layer8_outputs(3052)) xor (layer8_outputs(4938));
    outputs(1846) <= layer8_outputs(2684);
    outputs(1847) <= (layer8_outputs(71)) or (layer8_outputs(624));
    outputs(1848) <= layer8_outputs(3504);
    outputs(1849) <= not(layer8_outputs(4916));
    outputs(1850) <= not((layer8_outputs(652)) xor (layer8_outputs(1499)));
    outputs(1851) <= layer8_outputs(220);
    outputs(1852) <= not(layer8_outputs(3401));
    outputs(1853) <= (layer8_outputs(5072)) xor (layer8_outputs(3126));
    outputs(1854) <= (layer8_outputs(4687)) xor (layer8_outputs(3183));
    outputs(1855) <= not(layer8_outputs(3929));
    outputs(1856) <= (layer8_outputs(2299)) xor (layer8_outputs(5002));
    outputs(1857) <= not(layer8_outputs(1576));
    outputs(1858) <= not(layer8_outputs(4862));
    outputs(1859) <= not(layer8_outputs(859));
    outputs(1860) <= (layer8_outputs(499)) and not (layer8_outputs(2259));
    outputs(1861) <= (layer8_outputs(3995)) or (layer8_outputs(1640));
    outputs(1862) <= layer8_outputs(714);
    outputs(1863) <= (layer8_outputs(636)) xor (layer8_outputs(4599));
    outputs(1864) <= layer8_outputs(4987);
    outputs(1865) <= not(layer8_outputs(2713));
    outputs(1866) <= not((layer8_outputs(2161)) xor (layer8_outputs(1340)));
    outputs(1867) <= (layer8_outputs(2051)) or (layer8_outputs(872));
    outputs(1868) <= not(layer8_outputs(2980));
    outputs(1869) <= (layer8_outputs(825)) and not (layer8_outputs(4088));
    outputs(1870) <= not(layer8_outputs(3565));
    outputs(1871) <= not((layer8_outputs(1100)) xor (layer8_outputs(2571)));
    outputs(1872) <= (layer8_outputs(4352)) and not (layer8_outputs(136));
    outputs(1873) <= not(layer8_outputs(1771));
    outputs(1874) <= not(layer8_outputs(2266));
    outputs(1875) <= layer8_outputs(1111);
    outputs(1876) <= not(layer8_outputs(212));
    outputs(1877) <= not(layer8_outputs(4094)) or (layer8_outputs(1015));
    outputs(1878) <= (layer8_outputs(1918)) and not (layer8_outputs(4552));
    outputs(1879) <= not((layer8_outputs(1792)) xor (layer8_outputs(928)));
    outputs(1880) <= layer8_outputs(4050);
    outputs(1881) <= (layer8_outputs(4857)) xor (layer8_outputs(3169));
    outputs(1882) <= layer8_outputs(2342);
    outputs(1883) <= (layer8_outputs(3306)) and not (layer8_outputs(3032));
    outputs(1884) <= (layer8_outputs(3403)) and (layer8_outputs(3142));
    outputs(1885) <= not((layer8_outputs(421)) xor (layer8_outputs(3734)));
    outputs(1886) <= not((layer8_outputs(2323)) or (layer8_outputs(3992)));
    outputs(1887) <= not((layer8_outputs(1070)) xor (layer8_outputs(1431)));
    outputs(1888) <= (layer8_outputs(366)) and (layer8_outputs(4261));
    outputs(1889) <= not((layer8_outputs(5058)) xor (layer8_outputs(218)));
    outputs(1890) <= layer8_outputs(3112);
    outputs(1891) <= (layer8_outputs(4969)) xor (layer8_outputs(4258));
    outputs(1892) <= (layer8_outputs(4952)) xor (layer8_outputs(3859));
    outputs(1893) <= not((layer8_outputs(2275)) xor (layer8_outputs(2971)));
    outputs(1894) <= not(layer8_outputs(2676));
    outputs(1895) <= not(layer8_outputs(2983));
    outputs(1896) <= (layer8_outputs(323)) xor (layer8_outputs(3218));
    outputs(1897) <= layer8_outputs(3561);
    outputs(1898) <= not((layer8_outputs(1124)) xor (layer8_outputs(2584)));
    outputs(1899) <= not(layer8_outputs(4715));
    outputs(1900) <= not(layer8_outputs(4124));
    outputs(1901) <= not(layer8_outputs(1152));
    outputs(1902) <= layer8_outputs(868);
    outputs(1903) <= (layer8_outputs(2840)) xor (layer8_outputs(1509));
    outputs(1904) <= not(layer8_outputs(4730));
    outputs(1905) <= (layer8_outputs(1311)) and (layer8_outputs(855));
    outputs(1906) <= not(layer8_outputs(2655));
    outputs(1907) <= not((layer8_outputs(1010)) xor (layer8_outputs(4571)));
    outputs(1908) <= (layer8_outputs(3230)) or (layer8_outputs(2757));
    outputs(1909) <= not(layer8_outputs(3831));
    outputs(1910) <= not((layer8_outputs(3770)) xor (layer8_outputs(4873)));
    outputs(1911) <= not(layer8_outputs(4059));
    outputs(1912) <= layer8_outputs(516);
    outputs(1913) <= layer8_outputs(4530);
    outputs(1914) <= (layer8_outputs(590)) xor (layer8_outputs(5068));
    outputs(1915) <= not(layer8_outputs(1869));
    outputs(1916) <= not(layer8_outputs(766));
    outputs(1917) <= not((layer8_outputs(3033)) xor (layer8_outputs(3845)));
    outputs(1918) <= layer8_outputs(4013);
    outputs(1919) <= not(layer8_outputs(3476));
    outputs(1920) <= layer8_outputs(942);
    outputs(1921) <= layer8_outputs(551);
    outputs(1922) <= not((layer8_outputs(1386)) or (layer8_outputs(3616)));
    outputs(1923) <= (layer8_outputs(345)) and (layer8_outputs(2061));
    outputs(1924) <= layer8_outputs(1775);
    outputs(1925) <= not(layer8_outputs(2954));
    outputs(1926) <= not(layer8_outputs(3635));
    outputs(1927) <= layer8_outputs(704);
    outputs(1928) <= layer8_outputs(3892);
    outputs(1929) <= (layer8_outputs(4624)) xor (layer8_outputs(4794));
    outputs(1930) <= not(layer8_outputs(2581));
    outputs(1931) <= (layer8_outputs(3491)) and not (layer8_outputs(938));
    outputs(1932) <= layer8_outputs(3343);
    outputs(1933) <= not((layer8_outputs(1330)) xor (layer8_outputs(4291)));
    outputs(1934) <= layer8_outputs(5097);
    outputs(1935) <= (layer8_outputs(2234)) xor (layer8_outputs(109));
    outputs(1936) <= not(layer8_outputs(4095));
    outputs(1937) <= layer8_outputs(2691);
    outputs(1938) <= not(layer8_outputs(3917));
    outputs(1939) <= layer8_outputs(1677);
    outputs(1940) <= (layer8_outputs(3847)) and not (layer8_outputs(1623));
    outputs(1941) <= layer8_outputs(2345);
    outputs(1942) <= not(layer8_outputs(2301));
    outputs(1943) <= (layer8_outputs(2544)) xor (layer8_outputs(3442));
    outputs(1944) <= not((layer8_outputs(1846)) xor (layer8_outputs(3319)));
    outputs(1945) <= not((layer8_outputs(1576)) and (layer8_outputs(3357)));
    outputs(1946) <= not(layer8_outputs(4409));
    outputs(1947) <= not(layer8_outputs(1129));
    outputs(1948) <= layer8_outputs(1492);
    outputs(1949) <= not((layer8_outputs(3374)) or (layer8_outputs(3675)));
    outputs(1950) <= not((layer8_outputs(2878)) xor (layer8_outputs(1460)));
    outputs(1951) <= layer8_outputs(1399);
    outputs(1952) <= layer8_outputs(3621);
    outputs(1953) <= not(layer8_outputs(4970));
    outputs(1954) <= (layer8_outputs(3950)) and not (layer8_outputs(337));
    outputs(1955) <= (layer8_outputs(3195)) and not (layer8_outputs(3782));
    outputs(1956) <= layer8_outputs(351);
    outputs(1957) <= not(layer8_outputs(4570));
    outputs(1958) <= (layer8_outputs(3866)) xor (layer8_outputs(3281));
    outputs(1959) <= not(layer8_outputs(1365));
    outputs(1960) <= layer8_outputs(71);
    outputs(1961) <= not(layer8_outputs(1224));
    outputs(1962) <= not((layer8_outputs(2707)) xor (layer8_outputs(933)));
    outputs(1963) <= layer8_outputs(4363);
    outputs(1964) <= not(layer8_outputs(131));
    outputs(1965) <= layer8_outputs(1775);
    outputs(1966) <= not((layer8_outputs(1916)) xor (layer8_outputs(1679)));
    outputs(1967) <= (layer8_outputs(2560)) xor (layer8_outputs(1295));
    outputs(1968) <= layer8_outputs(2016);
    outputs(1969) <= layer8_outputs(1393);
    outputs(1970) <= (layer8_outputs(4056)) and not (layer8_outputs(2096));
    outputs(1971) <= layer8_outputs(1787);
    outputs(1972) <= layer8_outputs(4747);
    outputs(1973) <= not(layer8_outputs(4992));
    outputs(1974) <= layer8_outputs(4523);
    outputs(1975) <= not(layer8_outputs(4517));
    outputs(1976) <= not((layer8_outputs(2880)) and (layer8_outputs(1412)));
    outputs(1977) <= layer8_outputs(746);
    outputs(1978) <= not(layer8_outputs(592));
    outputs(1979) <= not((layer8_outputs(37)) xor (layer8_outputs(3852)));
    outputs(1980) <= not(layer8_outputs(584));
    outputs(1981) <= layer8_outputs(3031);
    outputs(1982) <= not(layer8_outputs(3485));
    outputs(1983) <= (layer8_outputs(1822)) xor (layer8_outputs(1573));
    outputs(1984) <= (layer8_outputs(4819)) xor (layer8_outputs(4599));
    outputs(1985) <= not((layer8_outputs(3633)) xor (layer8_outputs(3229)));
    outputs(1986) <= not(layer8_outputs(658));
    outputs(1987) <= layer8_outputs(3987);
    outputs(1988) <= layer8_outputs(849);
    outputs(1989) <= (layer8_outputs(4824)) xor (layer8_outputs(3745));
    outputs(1990) <= (layer8_outputs(4301)) xor (layer8_outputs(1367));
    outputs(1991) <= not(layer8_outputs(1797));
    outputs(1992) <= layer8_outputs(17);
    outputs(1993) <= layer8_outputs(3199);
    outputs(1994) <= not(layer8_outputs(1910));
    outputs(1995) <= (layer8_outputs(3207)) and (layer8_outputs(4028));
    outputs(1996) <= (layer8_outputs(4562)) xor (layer8_outputs(2884));
    outputs(1997) <= (layer8_outputs(1911)) and not (layer8_outputs(5064));
    outputs(1998) <= not((layer8_outputs(4989)) or (layer8_outputs(4135)));
    outputs(1999) <= not((layer8_outputs(3404)) xor (layer8_outputs(454)));
    outputs(2000) <= (layer8_outputs(1377)) xor (layer8_outputs(1402));
    outputs(2001) <= not(layer8_outputs(4449));
    outputs(2002) <= layer8_outputs(1107);
    outputs(2003) <= not(layer8_outputs(4820));
    outputs(2004) <= not(layer8_outputs(85));
    outputs(2005) <= (layer8_outputs(3096)) or (layer8_outputs(2879));
    outputs(2006) <= (layer8_outputs(617)) xor (layer8_outputs(3164));
    outputs(2007) <= layer8_outputs(3664);
    outputs(2008) <= layer8_outputs(3865);
    outputs(2009) <= not((layer8_outputs(829)) or (layer8_outputs(346)));
    outputs(2010) <= not((layer8_outputs(195)) or (layer8_outputs(5045)));
    outputs(2011) <= layer8_outputs(446);
    outputs(2012) <= not(layer8_outputs(1477));
    outputs(2013) <= not(layer8_outputs(4726));
    outputs(2014) <= not((layer8_outputs(4867)) or (layer8_outputs(2765)));
    outputs(2015) <= layer8_outputs(2620);
    outputs(2016) <= layer8_outputs(1256);
    outputs(2017) <= not(layer8_outputs(38));
    outputs(2018) <= (layer8_outputs(1746)) and not (layer8_outputs(483));
    outputs(2019) <= layer8_outputs(1378);
    outputs(2020) <= not((layer8_outputs(4439)) xor (layer8_outputs(2944)));
    outputs(2021) <= layer8_outputs(1705);
    outputs(2022) <= not(layer8_outputs(3730));
    outputs(2023) <= not((layer8_outputs(109)) xor (layer8_outputs(3925)));
    outputs(2024) <= not(layer8_outputs(1516));
    outputs(2025) <= not(layer8_outputs(635));
    outputs(2026) <= (layer8_outputs(3938)) and (layer8_outputs(4551));
    outputs(2027) <= (layer8_outputs(4762)) or (layer8_outputs(2091));
    outputs(2028) <= not((layer8_outputs(4776)) xor (layer8_outputs(4462)));
    outputs(2029) <= not((layer8_outputs(2742)) or (layer8_outputs(1894)));
    outputs(2030) <= not(layer8_outputs(724));
    outputs(2031) <= layer8_outputs(4871);
    outputs(2032) <= not(layer8_outputs(5095));
    outputs(2033) <= (layer8_outputs(4973)) and (layer8_outputs(3132));
    outputs(2034) <= layer8_outputs(2032);
    outputs(2035) <= not(layer8_outputs(3535));
    outputs(2036) <= not((layer8_outputs(1612)) xor (layer8_outputs(4959)));
    outputs(2037) <= (layer8_outputs(4561)) and not (layer8_outputs(3130));
    outputs(2038) <= (layer8_outputs(4092)) xor (layer8_outputs(4648));
    outputs(2039) <= (layer8_outputs(919)) and (layer8_outputs(2160));
    outputs(2040) <= layer8_outputs(3655);
    outputs(2041) <= not(layer8_outputs(1802));
    outputs(2042) <= not((layer8_outputs(1603)) xor (layer8_outputs(5065)));
    outputs(2043) <= (layer8_outputs(876)) xor (layer8_outputs(4789));
    outputs(2044) <= layer8_outputs(647);
    outputs(2045) <= not((layer8_outputs(2012)) xor (layer8_outputs(1938)));
    outputs(2046) <= not((layer8_outputs(3918)) and (layer8_outputs(3767)));
    outputs(2047) <= (layer8_outputs(3566)) xor (layer8_outputs(1310));
    outputs(2048) <= '0';
    outputs(2049) <= not(layer8_outputs(685));
    outputs(2050) <= layer8_outputs(4795);
    outputs(2051) <= not(layer8_outputs(1767)) or (layer8_outputs(818));
    outputs(2052) <= (layer8_outputs(1638)) xor (layer8_outputs(1294));
    outputs(2053) <= (layer8_outputs(4749)) xor (layer8_outputs(2883));
    outputs(2054) <= not(layer8_outputs(3390));
    outputs(2055) <= (layer8_outputs(1626)) xor (layer8_outputs(2705));
    outputs(2056) <= (layer8_outputs(1637)) xor (layer8_outputs(4961));
    outputs(2057) <= not(layer8_outputs(3526));
    outputs(2058) <= not((layer8_outputs(4311)) xor (layer8_outputs(2187)));
    outputs(2059) <= (layer8_outputs(576)) and (layer8_outputs(4740));
    outputs(2060) <= not(layer8_outputs(3049));
    outputs(2061) <= not((layer8_outputs(3185)) and (layer8_outputs(3217)));
    outputs(2062) <= layer8_outputs(1466);
    outputs(2063) <= layer8_outputs(4286);
    outputs(2064) <= not(layer8_outputs(4313));
    outputs(2065) <= layer8_outputs(3042);
    outputs(2066) <= not((layer8_outputs(3387)) xor (layer8_outputs(1384)));
    outputs(2067) <= not(layer8_outputs(2875));
    outputs(2068) <= not(layer8_outputs(4011));
    outputs(2069) <= layer8_outputs(3351);
    outputs(2070) <= layer8_outputs(3831);
    outputs(2071) <= layer8_outputs(766);
    outputs(2072) <= layer8_outputs(2646);
    outputs(2073) <= (layer8_outputs(801)) and not (layer8_outputs(2075));
    outputs(2074) <= (layer8_outputs(4170)) and not (layer8_outputs(4531));
    outputs(2075) <= (layer8_outputs(5083)) xor (layer8_outputs(2168));
    outputs(2076) <= (layer8_outputs(3435)) and not (layer8_outputs(222));
    outputs(2077) <= (layer8_outputs(3463)) xor (layer8_outputs(4897));
    outputs(2078) <= not(layer8_outputs(3541));
    outputs(2079) <= (layer8_outputs(1528)) or (layer8_outputs(3278));
    outputs(2080) <= not(layer8_outputs(4260));
    outputs(2081) <= (layer8_outputs(4881)) or (layer8_outputs(423));
    outputs(2082) <= layer8_outputs(1950);
    outputs(2083) <= layer8_outputs(3814);
    outputs(2084) <= not(layer8_outputs(2835));
    outputs(2085) <= not(layer8_outputs(4315));
    outputs(2086) <= not((layer8_outputs(980)) xor (layer8_outputs(4759)));
    outputs(2087) <= layer8_outputs(2128);
    outputs(2088) <= layer8_outputs(4809);
    outputs(2089) <= not(layer8_outputs(3763));
    outputs(2090) <= not((layer8_outputs(780)) xor (layer8_outputs(4414)));
    outputs(2091) <= not(layer8_outputs(668));
    outputs(2092) <= layer8_outputs(1994);
    outputs(2093) <= not((layer8_outputs(842)) xor (layer8_outputs(2154)));
    outputs(2094) <= not(layer8_outputs(4976));
    outputs(2095) <= (layer8_outputs(3648)) and not (layer8_outputs(4864));
    outputs(2096) <= not(layer8_outputs(3239));
    outputs(2097) <= layer8_outputs(2215);
    outputs(2098) <= (layer8_outputs(2781)) xor (layer8_outputs(3956));
    outputs(2099) <= not(layer8_outputs(476));
    outputs(2100) <= not(layer8_outputs(4802));
    outputs(2101) <= not(layer8_outputs(1143));
    outputs(2102) <= layer8_outputs(2143);
    outputs(2103) <= not((layer8_outputs(4771)) xor (layer8_outputs(3597)));
    outputs(2104) <= not((layer8_outputs(2465)) xor (layer8_outputs(4164)));
    outputs(2105) <= not(layer8_outputs(1951));
    outputs(2106) <= layer8_outputs(3624);
    outputs(2107) <= (layer8_outputs(2831)) and (layer8_outputs(134));
    outputs(2108) <= (layer8_outputs(2702)) xor (layer8_outputs(1118));
    outputs(2109) <= layer8_outputs(4103);
    outputs(2110) <= layer8_outputs(1702);
    outputs(2111) <= (layer8_outputs(234)) xor (layer8_outputs(2192));
    outputs(2112) <= not((layer8_outputs(1208)) xor (layer8_outputs(4675)));
    outputs(2113) <= (layer8_outputs(4568)) and (layer8_outputs(5115));
    outputs(2114) <= (layer8_outputs(3590)) and not (layer8_outputs(2668));
    outputs(2115) <= layer8_outputs(4745);
    outputs(2116) <= not((layer8_outputs(4622)) xor (layer8_outputs(1857)));
    outputs(2117) <= layer8_outputs(4408);
    outputs(2118) <= not(layer8_outputs(3271));
    outputs(2119) <= not(layer8_outputs(4259));
    outputs(2120) <= layer8_outputs(2787);
    outputs(2121) <= layer8_outputs(3555);
    outputs(2122) <= not(layer8_outputs(1574));
    outputs(2123) <= (layer8_outputs(1307)) and (layer8_outputs(3610));
    outputs(2124) <= not(layer8_outputs(769));
    outputs(2125) <= layer8_outputs(2285);
    outputs(2126) <= not(layer8_outputs(499));
    outputs(2127) <= layer8_outputs(2261);
    outputs(2128) <= (layer8_outputs(2666)) xor (layer8_outputs(1209));
    outputs(2129) <= not(layer8_outputs(516));
    outputs(2130) <= not(layer8_outputs(2347)) or (layer8_outputs(1802));
    outputs(2131) <= not(layer8_outputs(1854));
    outputs(2132) <= not(layer8_outputs(3986));
    outputs(2133) <= layer8_outputs(1434);
    outputs(2134) <= (layer8_outputs(4626)) or (layer8_outputs(1624));
    outputs(2135) <= not(layer8_outputs(3737)) or (layer8_outputs(4934));
    outputs(2136) <= not((layer8_outputs(3111)) and (layer8_outputs(4999)));
    outputs(2137) <= not(layer8_outputs(4120));
    outputs(2138) <= not((layer8_outputs(4333)) xor (layer8_outputs(1502)));
    outputs(2139) <= not((layer8_outputs(2766)) and (layer8_outputs(5091)));
    outputs(2140) <= not(layer8_outputs(1977)) or (layer8_outputs(246));
    outputs(2141) <= not(layer8_outputs(3100));
    outputs(2142) <= layer8_outputs(241);
    outputs(2143) <= (layer8_outputs(3733)) xor (layer8_outputs(831));
    outputs(2144) <= (layer8_outputs(1159)) or (layer8_outputs(1188));
    outputs(2145) <= (layer8_outputs(1865)) xor (layer8_outputs(1923));
    outputs(2146) <= layer8_outputs(4733);
    outputs(2147) <= not((layer8_outputs(3372)) xor (layer8_outputs(4262)));
    outputs(2148) <= not(layer8_outputs(2983));
    outputs(2149) <= not(layer8_outputs(641));
    outputs(2150) <= layer8_outputs(73);
    outputs(2151) <= layer8_outputs(3304);
    outputs(2152) <= not((layer8_outputs(3338)) xor (layer8_outputs(907)));
    outputs(2153) <= not(layer8_outputs(3108));
    outputs(2154) <= (layer8_outputs(1009)) and (layer8_outputs(3138));
    outputs(2155) <= not((layer8_outputs(2857)) xor (layer8_outputs(2516)));
    outputs(2156) <= not(layer8_outputs(4411));
    outputs(2157) <= not(layer8_outputs(2290));
    outputs(2158) <= layer8_outputs(2104);
    outputs(2159) <= (layer8_outputs(1263)) xor (layer8_outputs(4918));
    outputs(2160) <= layer8_outputs(3454);
    outputs(2161) <= layer8_outputs(2934);
    outputs(2162) <= layer8_outputs(4761);
    outputs(2163) <= not((layer8_outputs(4019)) xor (layer8_outputs(748)));
    outputs(2164) <= not((layer8_outputs(4482)) xor (layer8_outputs(4546)));
    outputs(2165) <= layer8_outputs(373);
    outputs(2166) <= layer8_outputs(321);
    outputs(2167) <= not(layer8_outputs(778));
    outputs(2168) <= not(layer8_outputs(678));
    outputs(2169) <= (layer8_outputs(4052)) xor (layer8_outputs(4675));
    outputs(2170) <= not(layer8_outputs(5049));
    outputs(2171) <= layer8_outputs(2353);
    outputs(2172) <= not(layer8_outputs(3057));
    outputs(2173) <= not(layer8_outputs(2717));
    outputs(2174) <= not(layer8_outputs(5));
    outputs(2175) <= layer8_outputs(3226);
    outputs(2176) <= not(layer8_outputs(4597));
    outputs(2177) <= not((layer8_outputs(2063)) xor (layer8_outputs(418)));
    outputs(2178) <= not(layer8_outputs(4566));
    outputs(2179) <= not(layer8_outputs(3563));
    outputs(2180) <= (layer8_outputs(1257)) and not (layer8_outputs(6));
    outputs(2181) <= not(layer8_outputs(2984));
    outputs(2182) <= (layer8_outputs(1536)) and (layer8_outputs(4396));
    outputs(2183) <= layer8_outputs(2315);
    outputs(2184) <= layer8_outputs(89);
    outputs(2185) <= not(layer8_outputs(2179));
    outputs(2186) <= not((layer8_outputs(537)) xor (layer8_outputs(3178)));
    outputs(2187) <= not(layer8_outputs(3057));
    outputs(2188) <= not(layer8_outputs(4230));
    outputs(2189) <= not(layer8_outputs(1336));
    outputs(2190) <= layer8_outputs(4195);
    outputs(2191) <= not(layer8_outputs(3054));
    outputs(2192) <= not(layer8_outputs(172));
    outputs(2193) <= (layer8_outputs(1956)) or (layer8_outputs(166));
    outputs(2194) <= layer8_outputs(4419);
    outputs(2195) <= layer8_outputs(4335);
    outputs(2196) <= layer8_outputs(1597);
    outputs(2197) <= (layer8_outputs(83)) xor (layer8_outputs(2393));
    outputs(2198) <= not(layer8_outputs(3270));
    outputs(2199) <= layer8_outputs(4508);
    outputs(2200) <= not((layer8_outputs(574)) xor (layer8_outputs(4750)));
    outputs(2201) <= not(layer8_outputs(1921));
    outputs(2202) <= layer8_outputs(3099);
    outputs(2203) <= (layer8_outputs(2310)) xor (layer8_outputs(1473));
    outputs(2204) <= not(layer8_outputs(1748));
    outputs(2205) <= not((layer8_outputs(1274)) xor (layer8_outputs(2141)));
    outputs(2206) <= layer8_outputs(3457);
    outputs(2207) <= not((layer8_outputs(726)) xor (layer8_outputs(1010)));
    outputs(2208) <= (layer8_outputs(737)) xor (layer8_outputs(2059));
    outputs(2209) <= (layer8_outputs(4591)) and not (layer8_outputs(4990));
    outputs(2210) <= (layer8_outputs(266)) and not (layer8_outputs(4979));
    outputs(2211) <= not(layer8_outputs(5071));
    outputs(2212) <= not((layer8_outputs(147)) xor (layer8_outputs(3149)));
    outputs(2213) <= layer8_outputs(3433);
    outputs(2214) <= not(layer8_outputs(2430));
    outputs(2215) <= not((layer8_outputs(177)) xor (layer8_outputs(1323)));
    outputs(2216) <= (layer8_outputs(531)) xor (layer8_outputs(4326));
    outputs(2217) <= (layer8_outputs(3542)) xor (layer8_outputs(3456));
    outputs(2218) <= not(layer8_outputs(4358));
    outputs(2219) <= not(layer8_outputs(2053));
    outputs(2220) <= not((layer8_outputs(275)) xor (layer8_outputs(1543)));
    outputs(2221) <= not(layer8_outputs(4560));
    outputs(2222) <= (layer8_outputs(1455)) and (layer8_outputs(2482));
    outputs(2223) <= not(layer8_outputs(193));
    outputs(2224) <= layer8_outputs(4955);
    outputs(2225) <= not((layer8_outputs(3023)) or (layer8_outputs(3494)));
    outputs(2226) <= not(layer8_outputs(4930));
    outputs(2227) <= (layer8_outputs(2506)) xor (layer8_outputs(559));
    outputs(2228) <= not(layer8_outputs(67));
    outputs(2229) <= (layer8_outputs(2673)) xor (layer8_outputs(4333));
    outputs(2230) <= not(layer8_outputs(458)) or (layer8_outputs(2399));
    outputs(2231) <= not(layer8_outputs(844));
    outputs(2232) <= not(layer8_outputs(2384));
    outputs(2233) <= layer8_outputs(557);
    outputs(2234) <= not((layer8_outputs(2645)) xor (layer8_outputs(279)));
    outputs(2235) <= layer8_outputs(4837);
    outputs(2236) <= not(layer8_outputs(755));
    outputs(2237) <= layer8_outputs(2097);
    outputs(2238) <= (layer8_outputs(2611)) and not (layer8_outputs(3514));
    outputs(2239) <= not(layer8_outputs(4532));
    outputs(2240) <= layer8_outputs(1230);
    outputs(2241) <= (layer8_outputs(3191)) xor (layer8_outputs(1864));
    outputs(2242) <= (layer8_outputs(4243)) and not (layer8_outputs(220));
    outputs(2243) <= layer8_outputs(5063);
    outputs(2244) <= (layer8_outputs(1394)) xor (layer8_outputs(3388));
    outputs(2245) <= layer8_outputs(4435);
    outputs(2246) <= layer8_outputs(1121);
    outputs(2247) <= not(layer8_outputs(3801));
    outputs(2248) <= layer8_outputs(2394);
    outputs(2249) <= not((layer8_outputs(180)) xor (layer8_outputs(1039)));
    outputs(2250) <= not(layer8_outputs(1992));
    outputs(2251) <= (layer8_outputs(1764)) xor (layer8_outputs(2915));
    outputs(2252) <= layer8_outputs(2967);
    outputs(2253) <= not(layer8_outputs(1905));
    outputs(2254) <= not((layer8_outputs(2392)) xor (layer8_outputs(4370)));
    outputs(2255) <= not(layer8_outputs(3216));
    outputs(2256) <= (layer8_outputs(3477)) and not (layer8_outputs(470));
    outputs(2257) <= not(layer8_outputs(1131));
    outputs(2258) <= (layer8_outputs(4377)) and not (layer8_outputs(4470));
    outputs(2259) <= (layer8_outputs(1440)) xor (layer8_outputs(3099));
    outputs(2260) <= not(layer8_outputs(3031));
    outputs(2261) <= not(layer8_outputs(1860));
    outputs(2262) <= (layer8_outputs(285)) xor (layer8_outputs(192));
    outputs(2263) <= (layer8_outputs(1887)) xor (layer8_outputs(1974));
    outputs(2264) <= (layer8_outputs(3804)) xor (layer8_outputs(4839));
    outputs(2265) <= (layer8_outputs(906)) and not (layer8_outputs(2430));
    outputs(2266) <= not((layer8_outputs(1440)) xor (layer8_outputs(4502)));
    outputs(2267) <= layer8_outputs(3041);
    outputs(2268) <= (layer8_outputs(136)) and not (layer8_outputs(4801));
    outputs(2269) <= not(layer8_outputs(4751)) or (layer8_outputs(4105));
    outputs(2270) <= layer8_outputs(5094);
    outputs(2271) <= (layer8_outputs(2469)) and not (layer8_outputs(2688));
    outputs(2272) <= not(layer8_outputs(3422));
    outputs(2273) <= layer8_outputs(2403);
    outputs(2274) <= not(layer8_outputs(2204));
    outputs(2275) <= layer8_outputs(2158);
    outputs(2276) <= (layer8_outputs(4881)) or (layer8_outputs(501));
    outputs(2277) <= not(layer8_outputs(2514));
    outputs(2278) <= (layer8_outputs(4048)) and not (layer8_outputs(1398));
    outputs(2279) <= not(layer8_outputs(2186));
    outputs(2280) <= layer8_outputs(4391);
    outputs(2281) <= layer8_outputs(602);
    outputs(2282) <= layer8_outputs(412);
    outputs(2283) <= layer8_outputs(329);
    outputs(2284) <= (layer8_outputs(167)) xor (layer8_outputs(22));
    outputs(2285) <= not(layer8_outputs(4769));
    outputs(2286) <= (layer8_outputs(2595)) xor (layer8_outputs(1451));
    outputs(2287) <= layer8_outputs(615);
    outputs(2288) <= layer8_outputs(4015);
    outputs(2289) <= layer8_outputs(4016);
    outputs(2290) <= layer8_outputs(1718);
    outputs(2291) <= not(layer8_outputs(4168));
    outputs(2292) <= not(layer8_outputs(757));
    outputs(2293) <= not((layer8_outputs(3000)) and (layer8_outputs(361)));
    outputs(2294) <= (layer8_outputs(3977)) or (layer8_outputs(4970));
    outputs(2295) <= layer8_outputs(2731);
    outputs(2296) <= layer8_outputs(1627);
    outputs(2297) <= not((layer8_outputs(2478)) or (layer8_outputs(2653)));
    outputs(2298) <= (layer8_outputs(90)) xor (layer8_outputs(3371));
    outputs(2299) <= (layer8_outputs(4133)) and (layer8_outputs(3214));
    outputs(2300) <= layer8_outputs(370);
    outputs(2301) <= not(layer8_outputs(2996));
    outputs(2302) <= layer8_outputs(1848);
    outputs(2303) <= not((layer8_outputs(4684)) xor (layer8_outputs(1072)));
    outputs(2304) <= layer8_outputs(645);
    outputs(2305) <= (layer8_outputs(1563)) xor (layer8_outputs(1648));
    outputs(2306) <= layer8_outputs(4381);
    outputs(2307) <= layer8_outputs(4465);
    outputs(2308) <= (layer8_outputs(4176)) xor (layer8_outputs(1818));
    outputs(2309) <= not(layer8_outputs(1249));
    outputs(2310) <= not((layer8_outputs(1073)) xor (layer8_outputs(4649)));
    outputs(2311) <= layer8_outputs(4516);
    outputs(2312) <= (layer8_outputs(3779)) xor (layer8_outputs(1449));
    outputs(2313) <= layer8_outputs(3978);
    outputs(2314) <= (layer8_outputs(2682)) and not (layer8_outputs(2080));
    outputs(2315) <= not((layer8_outputs(1970)) xor (layer8_outputs(3397)));
    outputs(2316) <= not((layer8_outputs(4353)) xor (layer8_outputs(1987)));
    outputs(2317) <= (layer8_outputs(4140)) xor (layer8_outputs(1868));
    outputs(2318) <= not((layer8_outputs(5087)) xor (layer8_outputs(1449)));
    outputs(2319) <= (layer8_outputs(1720)) xor (layer8_outputs(1979));
    outputs(2320) <= not((layer8_outputs(1161)) or (layer8_outputs(758)));
    outputs(2321) <= layer8_outputs(3536);
    outputs(2322) <= not(layer8_outputs(3276));
    outputs(2323) <= layer8_outputs(1313);
    outputs(2324) <= (layer8_outputs(1277)) and not (layer8_outputs(4298));
    outputs(2325) <= not(layer8_outputs(231));
    outputs(2326) <= not(layer8_outputs(3694));
    outputs(2327) <= not((layer8_outputs(2784)) xor (layer8_outputs(3474)));
    outputs(2328) <= not((layer8_outputs(54)) xor (layer8_outputs(4666)));
    outputs(2329) <= not(layer8_outputs(2426));
    outputs(2330) <= not(layer8_outputs(1190)) or (layer8_outputs(1599));
    outputs(2331) <= (layer8_outputs(2264)) xor (layer8_outputs(1258));
    outputs(2332) <= not(layer8_outputs(531));
    outputs(2333) <= layer8_outputs(3709);
    outputs(2334) <= layer8_outputs(4299);
    outputs(2335) <= not(layer8_outputs(2216));
    outputs(2336) <= not(layer8_outputs(4450));
    outputs(2337) <= layer8_outputs(4342);
    outputs(2338) <= (layer8_outputs(1915)) and not (layer8_outputs(1359));
    outputs(2339) <= not(layer8_outputs(3581));
    outputs(2340) <= layer8_outputs(1284);
    outputs(2341) <= not(layer8_outputs(609));
    outputs(2342) <= not((layer8_outputs(1909)) xor (layer8_outputs(4496)));
    outputs(2343) <= not(layer8_outputs(2256));
    outputs(2344) <= not((layer8_outputs(2343)) xor (layer8_outputs(4804)));
    outputs(2345) <= not((layer8_outputs(1901)) xor (layer8_outputs(4305)));
    outputs(2346) <= not(layer8_outputs(3647));
    outputs(2347) <= not(layer8_outputs(1007));
    outputs(2348) <= layer8_outputs(2210);
    outputs(2349) <= not(layer8_outputs(3308));
    outputs(2350) <= not(layer8_outputs(4156));
    outputs(2351) <= not(layer8_outputs(1808));
    outputs(2352) <= layer8_outputs(1246);
    outputs(2353) <= (layer8_outputs(2755)) or (layer8_outputs(148));
    outputs(2354) <= (layer8_outputs(4727)) or (layer8_outputs(649));
    outputs(2355) <= not((layer8_outputs(3805)) xor (layer8_outputs(4816)));
    outputs(2356) <= not((layer8_outputs(4455)) and (layer8_outputs(4139)));
    outputs(2357) <= (layer8_outputs(3294)) and not (layer8_outputs(565));
    outputs(2358) <= (layer8_outputs(573)) xor (layer8_outputs(420));
    outputs(2359) <= layer8_outputs(4068);
    outputs(2360) <= not(layer8_outputs(2626));
    outputs(2361) <= not((layer8_outputs(2597)) xor (layer8_outputs(3283)));
    outputs(2362) <= layer8_outputs(2400);
    outputs(2363) <= not(layer8_outputs(2575));
    outputs(2364) <= layer8_outputs(4280);
    outputs(2365) <= not(layer8_outputs(2146));
    outputs(2366) <= not((layer8_outputs(728)) or (layer8_outputs(3095)));
    outputs(2367) <= layer8_outputs(3373);
    outputs(2368) <= (layer8_outputs(3065)) xor (layer8_outputs(1008));
    outputs(2369) <= (layer8_outputs(332)) xor (layer8_outputs(4128));
    outputs(2370) <= (layer8_outputs(2705)) xor (layer8_outputs(796));
    outputs(2371) <= not(layer8_outputs(5071));
    outputs(2372) <= not((layer8_outputs(4822)) or (layer8_outputs(4223)));
    outputs(2373) <= layer8_outputs(4163);
    outputs(2374) <= layer8_outputs(4265);
    outputs(2375) <= not((layer8_outputs(5104)) xor (layer8_outputs(3994)));
    outputs(2376) <= not(layer8_outputs(4778));
    outputs(2377) <= not((layer8_outputs(456)) xor (layer8_outputs(4743)));
    outputs(2378) <= not((layer8_outputs(3857)) xor (layer8_outputs(4830)));
    outputs(2379) <= (layer8_outputs(2340)) xor (layer8_outputs(5085));
    outputs(2380) <= not(layer8_outputs(4301));
    outputs(2381) <= not((layer8_outputs(680)) xor (layer8_outputs(3568)));
    outputs(2382) <= (layer8_outputs(691)) or (layer8_outputs(4190));
    outputs(2383) <= not(layer8_outputs(5006));
    outputs(2384) <= layer8_outputs(2299);
    outputs(2385) <= layer8_outputs(2501);
    outputs(2386) <= not(layer8_outputs(1142));
    outputs(2387) <= not(layer8_outputs(2096));
    outputs(2388) <= not(layer8_outputs(654));
    outputs(2389) <= (layer8_outputs(4178)) xor (layer8_outputs(5100));
    outputs(2390) <= not(layer8_outputs(4685));
    outputs(2391) <= (layer8_outputs(43)) xor (layer8_outputs(1337));
    outputs(2392) <= not(layer8_outputs(1570));
    outputs(2393) <= not(layer8_outputs(3752)) or (layer8_outputs(2523));
    outputs(2394) <= not(layer8_outputs(3846)) or (layer8_outputs(1144));
    outputs(2395) <= (layer8_outputs(2105)) and not (layer8_outputs(3763));
    outputs(2396) <= (layer8_outputs(1930)) xor (layer8_outputs(2946));
    outputs(2397) <= (layer8_outputs(3760)) xor (layer8_outputs(2955));
    outputs(2398) <= (layer8_outputs(2579)) and not (layer8_outputs(3863));
    outputs(2399) <= not((layer8_outputs(2800)) xor (layer8_outputs(3725)));
    outputs(2400) <= not((layer8_outputs(3717)) xor (layer8_outputs(444)));
    outputs(2401) <= layer8_outputs(4648);
    outputs(2402) <= (layer8_outputs(3874)) xor (layer8_outputs(1360));
    outputs(2403) <= not(layer8_outputs(3187));
    outputs(2404) <= (layer8_outputs(5050)) and (layer8_outputs(1505));
    outputs(2405) <= (layer8_outputs(2349)) and (layer8_outputs(2267));
    outputs(2406) <= layer8_outputs(4031);
    outputs(2407) <= layer8_outputs(566);
    outputs(2408) <= layer8_outputs(2934);
    outputs(2409) <= not(layer8_outputs(4316));
    outputs(2410) <= not((layer8_outputs(292)) xor (layer8_outputs(1200)));
    outputs(2411) <= layer8_outputs(3700);
    outputs(2412) <= (layer8_outputs(2209)) and not (layer8_outputs(4481));
    outputs(2413) <= (layer8_outputs(2018)) xor (layer8_outputs(4898));
    outputs(2414) <= (layer8_outputs(1864)) xor (layer8_outputs(4191));
    outputs(2415) <= not(layer8_outputs(4364));
    outputs(2416) <= not(layer8_outputs(630));
    outputs(2417) <= not(layer8_outputs(3332));
    outputs(2418) <= layer8_outputs(1319);
    outputs(2419) <= (layer8_outputs(1865)) xor (layer8_outputs(4509));
    outputs(2420) <= not(layer8_outputs(1041));
    outputs(2421) <= not((layer8_outputs(2529)) xor (layer8_outputs(2930)));
    outputs(2422) <= not((layer8_outputs(1767)) xor (layer8_outputs(4849)));
    outputs(2423) <= layer8_outputs(3979);
    outputs(2424) <= not(layer8_outputs(2861));
    outputs(2425) <= layer8_outputs(3989);
    outputs(2426) <= layer8_outputs(5067);
    outputs(2427) <= not((layer8_outputs(290)) xor (layer8_outputs(4718)));
    outputs(2428) <= layer8_outputs(4644);
    outputs(2429) <= not(layer8_outputs(3510));
    outputs(2430) <= layer8_outputs(4445);
    outputs(2431) <= (layer8_outputs(3268)) and not (layer8_outputs(1233));
    outputs(2432) <= not((layer8_outputs(4431)) xor (layer8_outputs(3934)));
    outputs(2433) <= not(layer8_outputs(1168));
    outputs(2434) <= not(layer8_outputs(3312));
    outputs(2435) <= not(layer8_outputs(1116)) or (layer8_outputs(1836));
    outputs(2436) <= (layer8_outputs(1313)) xor (layer8_outputs(4700));
    outputs(2437) <= not(layer8_outputs(1730));
    outputs(2438) <= (layer8_outputs(2884)) xor (layer8_outputs(43));
    outputs(2439) <= layer8_outputs(2021);
    outputs(2440) <= not((layer8_outputs(1571)) xor (layer8_outputs(1251)));
    outputs(2441) <= layer8_outputs(4929);
    outputs(2442) <= not((layer8_outputs(763)) xor (layer8_outputs(1704)));
    outputs(2443) <= (layer8_outputs(833)) xor (layer8_outputs(4454));
    outputs(2444) <= layer8_outputs(2070);
    outputs(2445) <= not(layer8_outputs(461));
    outputs(2446) <= layer8_outputs(4440);
    outputs(2447) <= not(layer8_outputs(2518));
    outputs(2448) <= not(layer8_outputs(1317));
    outputs(2449) <= (layer8_outputs(389)) xor (layer8_outputs(3719));
    outputs(2450) <= (layer8_outputs(1349)) xor (layer8_outputs(1285));
    outputs(2451) <= not((layer8_outputs(3242)) xor (layer8_outputs(1191)));
    outputs(2452) <= layer8_outputs(3496);
    outputs(2453) <= not(layer8_outputs(4778));
    outputs(2454) <= not((layer8_outputs(4475)) xor (layer8_outputs(2686)));
    outputs(2455) <= not(layer8_outputs(2643)) or (layer8_outputs(4683));
    outputs(2456) <= (layer8_outputs(108)) or (layer8_outputs(192));
    outputs(2457) <= not(layer8_outputs(3107));
    outputs(2458) <= not((layer8_outputs(4521)) xor (layer8_outputs(3247)));
    outputs(2459) <= (layer8_outputs(3140)) and (layer8_outputs(2309));
    outputs(2460) <= not(layer8_outputs(947));
    outputs(2461) <= (layer8_outputs(2559)) xor (layer8_outputs(139));
    outputs(2462) <= (layer8_outputs(4186)) and not (layer8_outputs(959));
    outputs(2463) <= not(layer8_outputs(425)) or (layer8_outputs(3035));
    outputs(2464) <= (layer8_outputs(3532)) xor (layer8_outputs(1373));
    outputs(2465) <= (layer8_outputs(1853)) xor (layer8_outputs(1761));
    outputs(2466) <= (layer8_outputs(3803)) and (layer8_outputs(913));
    outputs(2467) <= not(layer8_outputs(24));
    outputs(2468) <= (layer8_outputs(5092)) xor (layer8_outputs(2235));
    outputs(2469) <= (layer8_outputs(1437)) and not (layer8_outputs(2733));
    outputs(2470) <= not((layer8_outputs(926)) and (layer8_outputs(390)));
    outputs(2471) <= not(layer8_outputs(3687));
    outputs(2472) <= layer8_outputs(1542);
    outputs(2473) <= layer8_outputs(3750);
    outputs(2474) <= layer8_outputs(1461);
    outputs(2475) <= layer8_outputs(4319);
    outputs(2476) <= layer8_outputs(2417);
    outputs(2477) <= layer8_outputs(196);
    outputs(2478) <= layer8_outputs(4518);
    outputs(2479) <= not((layer8_outputs(4630)) xor (layer8_outputs(3647)));
    outputs(2480) <= not(layer8_outputs(5048));
    outputs(2481) <= not(layer8_outputs(895));
    outputs(2482) <= not((layer8_outputs(3603)) xor (layer8_outputs(107)));
    outputs(2483) <= (layer8_outputs(5112)) xor (layer8_outputs(5000));
    outputs(2484) <= layer8_outputs(1278);
    outputs(2485) <= layer8_outputs(2066);
    outputs(2486) <= (layer8_outputs(3650)) xor (layer8_outputs(2319));
    outputs(2487) <= (layer8_outputs(1434)) and (layer8_outputs(2787));
    outputs(2488) <= not(layer8_outputs(1453)) or (layer8_outputs(5086));
    outputs(2489) <= (layer8_outputs(1162)) xor (layer8_outputs(2859));
    outputs(2490) <= not((layer8_outputs(1430)) xor (layer8_outputs(4513)));
    outputs(2491) <= not(layer8_outputs(4295)) or (layer8_outputs(380));
    outputs(2492) <= not((layer8_outputs(4006)) or (layer8_outputs(3269)));
    outputs(2493) <= layer8_outputs(1068);
    outputs(2494) <= not(layer8_outputs(335));
    outputs(2495) <= not((layer8_outputs(4670)) xor (layer8_outputs(3736)));
    outputs(2496) <= (layer8_outputs(3712)) and not (layer8_outputs(3014));
    outputs(2497) <= layer8_outputs(1561);
    outputs(2498) <= (layer8_outputs(151)) xor (layer8_outputs(1089));
    outputs(2499) <= layer8_outputs(3380);
    outputs(2500) <= layer8_outputs(892);
    outputs(2501) <= not((layer8_outputs(4322)) or (layer8_outputs(4082)));
    outputs(2502) <= (layer8_outputs(221)) and (layer8_outputs(4932));
    outputs(2503) <= layer8_outputs(3917);
    outputs(2504) <= not((layer8_outputs(1172)) xor (layer8_outputs(1656)));
    outputs(2505) <= layer8_outputs(954);
    outputs(2506) <= not(layer8_outputs(3829));
    outputs(2507) <= (layer8_outputs(208)) xor (layer8_outputs(839));
    outputs(2508) <= layer8_outputs(2070);
    outputs(2509) <= layer8_outputs(4530);
    outputs(2510) <= layer8_outputs(729);
    outputs(2511) <= not(layer8_outputs(3333));
    outputs(2512) <= not(layer8_outputs(2368));
    outputs(2513) <= not(layer8_outputs(3840));
    outputs(2514) <= not(layer8_outputs(4321));
    outputs(2515) <= (layer8_outputs(882)) and (layer8_outputs(3862));
    outputs(2516) <= (layer8_outputs(2910)) and not (layer8_outputs(1409));
    outputs(2517) <= layer8_outputs(1891);
    outputs(2518) <= not(layer8_outputs(713)) or (layer8_outputs(368));
    outputs(2519) <= layer8_outputs(4533);
    outputs(2520) <= not(layer8_outputs(4645));
    outputs(2521) <= layer8_outputs(2059);
    outputs(2522) <= layer8_outputs(2315);
    outputs(2523) <= (layer8_outputs(587)) xor (layer8_outputs(1419));
    outputs(2524) <= layer8_outputs(882);
    outputs(2525) <= (layer8_outputs(2057)) xor (layer8_outputs(3764));
    outputs(2526) <= not(layer8_outputs(2431));
    outputs(2527) <= (layer8_outputs(2114)) xor (layer8_outputs(2775));
    outputs(2528) <= not(layer8_outputs(5054));
    outputs(2529) <= layer8_outputs(3612);
    outputs(2530) <= not(layer8_outputs(4149));
    outputs(2531) <= (layer8_outputs(1094)) xor (layer8_outputs(1799));
    outputs(2532) <= layer8_outputs(5076);
    outputs(2533) <= layer8_outputs(201);
    outputs(2534) <= not(layer8_outputs(4216));
    outputs(2535) <= not(layer8_outputs(830));
    outputs(2536) <= layer8_outputs(69);
    outputs(2537) <= layer8_outputs(4297);
    outputs(2538) <= layer8_outputs(822);
    outputs(2539) <= (layer8_outputs(4909)) xor (layer8_outputs(3644));
    outputs(2540) <= not(layer8_outputs(860));
    outputs(2541) <= layer8_outputs(796);
    outputs(2542) <= (layer8_outputs(1423)) and not (layer8_outputs(620));
    outputs(2543) <= layer8_outputs(4968);
    outputs(2544) <= (layer8_outputs(48)) xor (layer8_outputs(2410));
    outputs(2545) <= (layer8_outputs(1892)) xor (layer8_outputs(2489));
    outputs(2546) <= layer8_outputs(2360);
    outputs(2547) <= layer8_outputs(645);
    outputs(2548) <= not(layer8_outputs(328));
    outputs(2549) <= not(layer8_outputs(1765));
    outputs(2550) <= (layer8_outputs(2665)) xor (layer8_outputs(2439));
    outputs(2551) <= layer8_outputs(2820);
    outputs(2552) <= not((layer8_outputs(4663)) xor (layer8_outputs(4154)));
    outputs(2553) <= not(layer8_outputs(1011)) or (layer8_outputs(2672));
    outputs(2554) <= not((layer8_outputs(884)) xor (layer8_outputs(3087)));
    outputs(2555) <= (layer8_outputs(4379)) and not (layer8_outputs(2559));
    outputs(2556) <= not(layer8_outputs(4418)) or (layer8_outputs(1944));
    outputs(2557) <= not(layer8_outputs(2823));
    outputs(2558) <= layer8_outputs(3383);
    outputs(2559) <= not(layer8_outputs(506));
    outputs(2560) <= not(layer8_outputs(2105)) or (layer8_outputs(4973));
    outputs(2561) <= not(layer8_outputs(1302));
    outputs(2562) <= (layer8_outputs(4856)) xor (layer8_outputs(694));
    outputs(2563) <= (layer8_outputs(3548)) xor (layer8_outputs(4631));
    outputs(2564) <= not(layer8_outputs(2599));
    outputs(2565) <= not((layer8_outputs(1206)) xor (layer8_outputs(1262)));
    outputs(2566) <= (layer8_outputs(4779)) xor (layer8_outputs(1729));
    outputs(2567) <= not(layer8_outputs(3411));
    outputs(2568) <= (layer8_outputs(4061)) xor (layer8_outputs(131));
    outputs(2569) <= not(layer8_outputs(1297));
    outputs(2570) <= (layer8_outputs(1793)) and (layer8_outputs(2897));
    outputs(2571) <= not((layer8_outputs(3134)) xor (layer8_outputs(912)));
    outputs(2572) <= not((layer8_outputs(4207)) xor (layer8_outputs(4812)));
    outputs(2573) <= layer8_outputs(5036);
    outputs(2574) <= not((layer8_outputs(1247)) xor (layer8_outputs(159)));
    outputs(2575) <= not((layer8_outputs(3698)) xor (layer8_outputs(3493)));
    outputs(2576) <= not(layer8_outputs(4568));
    outputs(2577) <= not(layer8_outputs(250)) or (layer8_outputs(2079));
    outputs(2578) <= (layer8_outputs(2505)) xor (layer8_outputs(1074));
    outputs(2579) <= layer8_outputs(1456);
    outputs(2580) <= not(layer8_outputs(498)) or (layer8_outputs(2240));
    outputs(2581) <= (layer8_outputs(4495)) xor (layer8_outputs(4598));
    outputs(2582) <= (layer8_outputs(3579)) or (layer8_outputs(4197));
    outputs(2583) <= not(layer8_outputs(2279));
    outputs(2584) <= layer8_outputs(3464);
    outputs(2585) <= not(layer8_outputs(488));
    outputs(2586) <= not(layer8_outputs(2717));
    outputs(2587) <= not((layer8_outputs(2395)) xor (layer8_outputs(2107)));
    outputs(2588) <= not((layer8_outputs(1560)) xor (layer8_outputs(3241)));
    outputs(2589) <= layer8_outputs(3926);
    outputs(2590) <= layer8_outputs(4349);
    outputs(2591) <= layer8_outputs(117);
    outputs(2592) <= not(layer8_outputs(4890));
    outputs(2593) <= not(layer8_outputs(1685));
    outputs(2594) <= (layer8_outputs(2145)) xor (layer8_outputs(57));
    outputs(2595) <= layer8_outputs(4492);
    outputs(2596) <= not(layer8_outputs(4922));
    outputs(2597) <= (layer8_outputs(4842)) xor (layer8_outputs(3086));
    outputs(2598) <= not((layer8_outputs(4041)) xor (layer8_outputs(4256)));
    outputs(2599) <= not(layer8_outputs(982));
    outputs(2600) <= (layer8_outputs(2546)) xor (layer8_outputs(4698));
    outputs(2601) <= (layer8_outputs(802)) xor (layer8_outputs(3073));
    outputs(2602) <= not(layer8_outputs(2487));
    outputs(2603) <= layer8_outputs(3158);
    outputs(2604) <= (layer8_outputs(3003)) and not (layer8_outputs(973));
    outputs(2605) <= not(layer8_outputs(3673));
    outputs(2606) <= not((layer8_outputs(3179)) and (layer8_outputs(897)));
    outputs(2607) <= layer8_outputs(335);
    outputs(2608) <= layer8_outputs(3206);
    outputs(2609) <= (layer8_outputs(2628)) xor (layer8_outputs(2534));
    outputs(2610) <= not(layer8_outputs(762));
    outputs(2611) <= layer8_outputs(1201);
    outputs(2612) <= not(layer8_outputs(4345));
    outputs(2613) <= not(layer8_outputs(1883));
    outputs(2614) <= layer8_outputs(137);
    outputs(2615) <= layer8_outputs(3024);
    outputs(2616) <= layer8_outputs(3131);
    outputs(2617) <= not(layer8_outputs(4513));
    outputs(2618) <= not((layer8_outputs(3090)) xor (layer8_outputs(2499)));
    outputs(2619) <= not(layer8_outputs(3498));
    outputs(2620) <= layer8_outputs(4960);
    outputs(2621) <= not(layer8_outputs(3310));
    outputs(2622) <= not(layer8_outputs(452));
    outputs(2623) <= not((layer8_outputs(736)) xor (layer8_outputs(4328)));
    outputs(2624) <= not((layer8_outputs(4291)) or (layer8_outputs(3399)));
    outputs(2625) <= not(layer8_outputs(3649));
    outputs(2626) <= not(layer8_outputs(3744));
    outputs(2627) <= not(layer8_outputs(3128));
    outputs(2628) <= not((layer8_outputs(4502)) xor (layer8_outputs(1799)));
    outputs(2629) <= layer8_outputs(1758);
    outputs(2630) <= layer8_outputs(5076);
    outputs(2631) <= (layer8_outputs(1098)) xor (layer8_outputs(2320));
    outputs(2632) <= (layer8_outputs(2347)) xor (layer8_outputs(3176));
    outputs(2633) <= not((layer8_outputs(66)) xor (layer8_outputs(3352)));
    outputs(2634) <= (layer8_outputs(1875)) and not (layer8_outputs(1621));
    outputs(2635) <= not(layer8_outputs(97));
    outputs(2636) <= not(layer8_outputs(2569));
    outputs(2637) <= (layer8_outputs(4885)) xor (layer8_outputs(4453));
    outputs(2638) <= (layer8_outputs(3833)) xor (layer8_outputs(1027));
    outputs(2639) <= not(layer8_outputs(611));
    outputs(2640) <= not(layer8_outputs(658));
    outputs(2641) <= (layer8_outputs(3454)) xor (layer8_outputs(4804));
    outputs(2642) <= (layer8_outputs(3150)) xor (layer8_outputs(4566));
    outputs(2643) <= not((layer8_outputs(334)) xor (layer8_outputs(160)));
    outputs(2644) <= not((layer8_outputs(1875)) xor (layer8_outputs(3471)));
    outputs(2645) <= not(layer8_outputs(1682));
    outputs(2646) <= not((layer8_outputs(1169)) xor (layer8_outputs(2535)));
    outputs(2647) <= not(layer8_outputs(110));
    outputs(2648) <= layer8_outputs(3222);
    outputs(2649) <= (layer8_outputs(4824)) xor (layer8_outputs(2786));
    outputs(2650) <= not((layer8_outputs(1502)) xor (layer8_outputs(4423)));
    outputs(2651) <= not(layer8_outputs(1790));
    outputs(2652) <= not(layer8_outputs(1062)) or (layer8_outputs(298));
    outputs(2653) <= layer8_outputs(4153);
    outputs(2654) <= layer8_outputs(2964);
    outputs(2655) <= not(layer8_outputs(988));
    outputs(2656) <= layer8_outputs(407);
    outputs(2657) <= (layer8_outputs(1441)) xor (layer8_outputs(304));
    outputs(2658) <= layer8_outputs(2811);
    outputs(2659) <= not(layer8_outputs(1849));
    outputs(2660) <= not((layer8_outputs(1791)) or (layer8_outputs(4607)));
    outputs(2661) <= not(layer8_outputs(2403));
    outputs(2662) <= not(layer8_outputs(2775));
    outputs(2663) <= not((layer8_outputs(3860)) xor (layer8_outputs(1049)));
    outputs(2664) <= layer8_outputs(1033);
    outputs(2665) <= layer8_outputs(3136);
    outputs(2666) <= not(layer8_outputs(1050)) or (layer8_outputs(773));
    outputs(2667) <= not(layer8_outputs(4148));
    outputs(2668) <= (layer8_outputs(986)) xor (layer8_outputs(1770));
    outputs(2669) <= (layer8_outputs(4074)) and (layer8_outputs(285));
    outputs(2670) <= layer8_outputs(4695);
    outputs(2671) <= layer8_outputs(589);
    outputs(2672) <= not((layer8_outputs(3067)) xor (layer8_outputs(4387)));
    outputs(2673) <= (layer8_outputs(672)) and not (layer8_outputs(396));
    outputs(2674) <= layer8_outputs(1325);
    outputs(2675) <= not(layer8_outputs(1242));
    outputs(2676) <= not(layer8_outputs(268));
    outputs(2677) <= not((layer8_outputs(2772)) xor (layer8_outputs(351)));
    outputs(2678) <= not((layer8_outputs(3991)) and (layer8_outputs(4962)));
    outputs(2679) <= layer8_outputs(824);
    outputs(2680) <= not(layer8_outputs(3867));
    outputs(2681) <= (layer8_outputs(4044)) xor (layer8_outputs(3895));
    outputs(2682) <= (layer8_outputs(40)) and not (layer8_outputs(2140));
    outputs(2683) <= not(layer8_outputs(1259));
    outputs(2684) <= not(layer8_outputs(1102)) or (layer8_outputs(3006));
    outputs(2685) <= not(layer8_outputs(4078));
    outputs(2686) <= not(layer8_outputs(44)) or (layer8_outputs(1467));
    outputs(2687) <= layer8_outputs(2650);
    outputs(2688) <= not((layer8_outputs(1387)) xor (layer8_outputs(4814)));
    outputs(2689) <= not((layer8_outputs(1261)) xor (layer8_outputs(1715)));
    outputs(2690) <= layer8_outputs(4656);
    outputs(2691) <= layer8_outputs(2188);
    outputs(2692) <= (layer8_outputs(719)) xor (layer8_outputs(3887));
    outputs(2693) <= not((layer8_outputs(3930)) xor (layer8_outputs(1001)));
    outputs(2694) <= layer8_outputs(3114);
    outputs(2695) <= not(layer8_outputs(732));
    outputs(2696) <= (layer8_outputs(2703)) and not (layer8_outputs(3919));
    outputs(2697) <= not(layer8_outputs(4536));
    outputs(2698) <= not((layer8_outputs(2861)) or (layer8_outputs(2827)));
    outputs(2699) <= not((layer8_outputs(4410)) xor (layer8_outputs(2402)));
    outputs(2700) <= not((layer8_outputs(2802)) xor (layer8_outputs(5025)));
    outputs(2701) <= not(layer8_outputs(1192));
    outputs(2702) <= (layer8_outputs(505)) and not (layer8_outputs(4827));
    outputs(2703) <= (layer8_outputs(4741)) and not (layer8_outputs(1210));
    outputs(2704) <= not(layer8_outputs(2753)) or (layer8_outputs(3921));
    outputs(2705) <= not(layer8_outputs(219));
    outputs(2706) <= (layer8_outputs(1953)) and not (layer8_outputs(68));
    outputs(2707) <= layer8_outputs(2272);
    outputs(2708) <= layer8_outputs(4191);
    outputs(2709) <= not(layer8_outputs(4144));
    outputs(2710) <= layer8_outputs(641);
    outputs(2711) <= not(layer8_outputs(2871));
    outputs(2712) <= (layer8_outputs(2354)) xor (layer8_outputs(4942));
    outputs(2713) <= layer8_outputs(2745);
    outputs(2714) <= layer8_outputs(3101);
    outputs(2715) <= not(layer8_outputs(647));
    outputs(2716) <= not(layer8_outputs(4629));
    outputs(2717) <= not((layer8_outputs(1016)) xor (layer8_outputs(1344)));
    outputs(2718) <= not(layer8_outputs(549)) or (layer8_outputs(3350));
    outputs(2719) <= not((layer8_outputs(793)) xor (layer8_outputs(1375)));
    outputs(2720) <= not(layer8_outputs(2965));
    outputs(2721) <= not(layer8_outputs(1005));
    outputs(2722) <= not((layer8_outputs(2780)) xor (layer8_outputs(464)));
    outputs(2723) <= not(layer8_outputs(2008));
    outputs(2724) <= not((layer8_outputs(2993)) xor (layer8_outputs(4395)));
    outputs(2725) <= not((layer8_outputs(3653)) xor (layer8_outputs(1272)));
    outputs(2726) <= not(layer8_outputs(37));
    outputs(2727) <= not((layer8_outputs(3335)) xor (layer8_outputs(3809)));
    outputs(2728) <= not(layer8_outputs(92));
    outputs(2729) <= not(layer8_outputs(2689));
    outputs(2730) <= not(layer8_outputs(4308));
    outputs(2731) <= not(layer8_outputs(1791));
    outputs(2732) <= (layer8_outputs(3115)) xor (layer8_outputs(3588));
    outputs(2733) <= not(layer8_outputs(2626));
    outputs(2734) <= layer8_outputs(5075);
    outputs(2735) <= (layer8_outputs(2621)) xor (layer8_outputs(2015));
    outputs(2736) <= layer8_outputs(2419);
    outputs(2737) <= not((layer8_outputs(4430)) or (layer8_outputs(3557)));
    outputs(2738) <= layer8_outputs(3420);
    outputs(2739) <= layer8_outputs(181);
    outputs(2740) <= not(layer8_outputs(3692));
    outputs(2741) <= not((layer8_outputs(4783)) xor (layer8_outputs(1901)));
    outputs(2742) <= layer8_outputs(2638);
    outputs(2743) <= layer8_outputs(2896);
    outputs(2744) <= not((layer8_outputs(1229)) xor (layer8_outputs(2445)));
    outputs(2745) <= (layer8_outputs(1178)) xor (layer8_outputs(60));
    outputs(2746) <= not(layer8_outputs(1998));
    outputs(2747) <= layer8_outputs(2609);
    outputs(2748) <= not(layer8_outputs(1444));
    outputs(2749) <= not(layer8_outputs(340));
    outputs(2750) <= not(layer8_outputs(2738));
    outputs(2751) <= not(layer8_outputs(1383));
    outputs(2752) <= (layer8_outputs(4980)) xor (layer8_outputs(2993));
    outputs(2753) <= not(layer8_outputs(3735));
    outputs(2754) <= not((layer8_outputs(570)) xor (layer8_outputs(4646)));
    outputs(2755) <= not((layer8_outputs(3912)) xor (layer8_outputs(1676)));
    outputs(2756) <= layer8_outputs(3433);
    outputs(2757) <= not(layer8_outputs(1826));
    outputs(2758) <= not(layer8_outputs(89));
    outputs(2759) <= layer8_outputs(2926);
    outputs(2760) <= not((layer8_outputs(896)) xor (layer8_outputs(3070)));
    outputs(2761) <= (layer8_outputs(205)) xor (layer8_outputs(3956));
    outputs(2762) <= not((layer8_outputs(784)) xor (layer8_outputs(4396)));
    outputs(2763) <= not((layer8_outputs(1806)) xor (layer8_outputs(545)));
    outputs(2764) <= (layer8_outputs(4920)) and not (layer8_outputs(404));
    outputs(2765) <= layer8_outputs(974);
    outputs(2766) <= (layer8_outputs(1194)) xor (layer8_outputs(4017));
    outputs(2767) <= layer8_outputs(992);
    outputs(2768) <= not(layer8_outputs(496));
    outputs(2769) <= (layer8_outputs(3521)) xor (layer8_outputs(1384));
    outputs(2770) <= not(layer8_outputs(2282));
    outputs(2771) <= not((layer8_outputs(3378)) or (layer8_outputs(3620)));
    outputs(2772) <= layer8_outputs(4079);
    outputs(2773) <= layer8_outputs(176);
    outputs(2774) <= layer8_outputs(3889);
    outputs(2775) <= (layer8_outputs(2511)) xor (layer8_outputs(2357));
    outputs(2776) <= not((layer8_outputs(1299)) and (layer8_outputs(2600)));
    outputs(2777) <= not((layer8_outputs(4208)) or (layer8_outputs(1908)));
    outputs(2778) <= (layer8_outputs(1579)) and not (layer8_outputs(1302));
    outputs(2779) <= not(layer8_outputs(4397));
    outputs(2780) <= not(layer8_outputs(4606));
    outputs(2781) <= not(layer8_outputs(1087));
    outputs(2782) <= not(layer8_outputs(1681));
    outputs(2783) <= (layer8_outputs(3265)) and not (layer8_outputs(1251));
    outputs(2784) <= layer8_outputs(898);
    outputs(2785) <= layer8_outputs(5114);
    outputs(2786) <= layer8_outputs(5022);
    outputs(2787) <= not(layer8_outputs(272));
    outputs(2788) <= layer8_outputs(2824);
    outputs(2789) <= (layer8_outputs(4136)) xor (layer8_outputs(1463));
    outputs(2790) <= not((layer8_outputs(2955)) xor (layer8_outputs(588)));
    outputs(2791) <= layer8_outputs(4394);
    outputs(2792) <= not((layer8_outputs(916)) xor (layer8_outputs(4307)));
    outputs(2793) <= layer8_outputs(1418);
    outputs(2794) <= not(layer8_outputs(4324));
    outputs(2795) <= not((layer8_outputs(84)) or (layer8_outputs(1092)));
    outputs(2796) <= not(layer8_outputs(2071));
    outputs(2797) <= not(layer8_outputs(4293));
    outputs(2798) <= (layer8_outputs(3915)) xor (layer8_outputs(4654));
    outputs(2799) <= not((layer8_outputs(2428)) or (layer8_outputs(4522)));
    outputs(2800) <= (layer8_outputs(4787)) xor (layer8_outputs(1414));
    outputs(2801) <= not(layer8_outputs(419));
    outputs(2802) <= layer8_outputs(3555);
    outputs(2803) <= not(layer8_outputs(3182));
    outputs(2804) <= layer8_outputs(1530);
    outputs(2805) <= (layer8_outputs(2196)) xor (layer8_outputs(1506));
    outputs(2806) <= (layer8_outputs(2944)) and not (layer8_outputs(4053));
    outputs(2807) <= not(layer8_outputs(628));
    outputs(2808) <= (layer8_outputs(2182)) xor (layer8_outputs(1281));
    outputs(2809) <= not(layer8_outputs(2162));
    outputs(2810) <= (layer8_outputs(1514)) xor (layer8_outputs(4443));
    outputs(2811) <= not((layer8_outputs(9)) xor (layer8_outputs(2396)));
    outputs(2812) <= not(layer8_outputs(3286));
    outputs(2813) <= layer8_outputs(2851);
    outputs(2814) <= (layer8_outputs(118)) and not (layer8_outputs(1589));
    outputs(2815) <= not(layer8_outputs(3300));
    outputs(2816) <= not(layer8_outputs(5027));
    outputs(2817) <= layer8_outputs(1480);
    outputs(2818) <= layer8_outputs(1485);
    outputs(2819) <= not(layer8_outputs(3256));
    outputs(2820) <= not(layer8_outputs(1123));
    outputs(2821) <= layer8_outputs(417);
    outputs(2822) <= layer8_outputs(2306);
    outputs(2823) <= not(layer8_outputs(3182));
    outputs(2824) <= not((layer8_outputs(3311)) xor (layer8_outputs(468)));
    outputs(2825) <= not((layer8_outputs(630)) xor (layer8_outputs(101)));
    outputs(2826) <= layer8_outputs(302);
    outputs(2827) <= not(layer8_outputs(2723));
    outputs(2828) <= not(layer8_outputs(976));
    outputs(2829) <= (layer8_outputs(4102)) and not (layer8_outputs(2805));
    outputs(2830) <= layer8_outputs(2005);
    outputs(2831) <= layer8_outputs(3082);
    outputs(2832) <= layer8_outputs(3766);
    outputs(2833) <= not((layer8_outputs(836)) xor (layer8_outputs(2033)));
    outputs(2834) <= not(layer8_outputs(3963));
    outputs(2835) <= not(layer8_outputs(2881));
    outputs(2836) <= (layer8_outputs(3983)) xor (layer8_outputs(1760));
    outputs(2837) <= layer8_outputs(3623);
    outputs(2838) <= layer8_outputs(4132);
    outputs(2839) <= (layer8_outputs(972)) or (layer8_outputs(4785));
    outputs(2840) <= layer8_outputs(2214);
    outputs(2841) <= layer8_outputs(2446);
    outputs(2842) <= not(layer8_outputs(2089));
    outputs(2843) <= (layer8_outputs(117)) and not (layer8_outputs(4951));
    outputs(2844) <= not((layer8_outputs(1122)) xor (layer8_outputs(119)));
    outputs(2845) <= not((layer8_outputs(2975)) xor (layer8_outputs(4833)));
    outputs(2846) <= not((layer8_outputs(1528)) or (layer8_outputs(4533)));
    outputs(2847) <= not(layer8_outputs(2094));
    outputs(2848) <= not(layer8_outputs(1542));
    outputs(2849) <= (layer8_outputs(1671)) xor (layer8_outputs(3078));
    outputs(2850) <= (layer8_outputs(3886)) xor (layer8_outputs(5070));
    outputs(2851) <= layer8_outputs(2405);
    outputs(2852) <= not(layer8_outputs(558));
    outputs(2853) <= (layer8_outputs(4782)) xor (layer8_outputs(873));
    outputs(2854) <= not(layer8_outputs(3728));
    outputs(2855) <= not(layer8_outputs(4276));
    outputs(2856) <= (layer8_outputs(2359)) xor (layer8_outputs(4274));
    outputs(2857) <= not((layer8_outputs(3526)) xor (layer8_outputs(4084)));
    outputs(2858) <= (layer8_outputs(320)) and not (layer8_outputs(4210));
    outputs(2859) <= layer8_outputs(4029);
    outputs(2860) <= layer8_outputs(4679);
    outputs(2861) <= not((layer8_outputs(435)) xor (layer8_outputs(4486)));
    outputs(2862) <= (layer8_outputs(2271)) xor (layer8_outputs(4122));
    outputs(2863) <= (layer8_outputs(2927)) xor (layer8_outputs(1636));
    outputs(2864) <= not((layer8_outputs(1086)) or (layer8_outputs(621)));
    outputs(2865) <= layer8_outputs(2180);
    outputs(2866) <= layer8_outputs(3513);
    outputs(2867) <= (layer8_outputs(40)) and not (layer8_outputs(3180));
    outputs(2868) <= layer8_outputs(740);
    outputs(2869) <= (layer8_outputs(4026)) xor (layer8_outputs(2018));
    outputs(2870) <= not(layer8_outputs(2222));
    outputs(2871) <= not(layer8_outputs(3716));
    outputs(2872) <= not(layer8_outputs(3325));
    outputs(2873) <= (layer8_outputs(3939)) xor (layer8_outputs(1315));
    outputs(2874) <= (layer8_outputs(502)) and (layer8_outputs(365));
    outputs(2875) <= layer8_outputs(4893);
    outputs(2876) <= (layer8_outputs(2321)) xor (layer8_outputs(3713));
    outputs(2877) <= layer8_outputs(1481);
    outputs(2878) <= layer8_outputs(2027);
    outputs(2879) <= layer8_outputs(1348);
    outputs(2880) <= (layer8_outputs(966)) xor (layer8_outputs(4162));
    outputs(2881) <= (layer8_outputs(3010)) xor (layer8_outputs(4882));
    outputs(2882) <= not(layer8_outputs(5080));
    outputs(2883) <= (layer8_outputs(2296)) xor (layer8_outputs(1586));
    outputs(2884) <= (layer8_outputs(4815)) xor (layer8_outputs(843));
    outputs(2885) <= not((layer8_outputs(1361)) xor (layer8_outputs(312)));
    outputs(2886) <= not(layer8_outputs(5033));
    outputs(2887) <= not((layer8_outputs(4693)) xor (layer8_outputs(3362)));
    outputs(2888) <= (layer8_outputs(2181)) and (layer8_outputs(1742));
    outputs(2889) <= not(layer8_outputs(2492));
    outputs(2890) <= (layer8_outputs(1143)) xor (layer8_outputs(4590));
    outputs(2891) <= layer8_outputs(378);
    outputs(2892) <= not((layer8_outputs(1518)) xor (layer8_outputs(2283)));
    outputs(2893) <= not(layer8_outputs(4900));
    outputs(2894) <= layer8_outputs(4756);
    outputs(2895) <= layer8_outputs(966);
    outputs(2896) <= layer8_outputs(150);
    outputs(2897) <= layer8_outputs(1511);
    outputs(2898) <= (layer8_outputs(462)) xor (layer8_outputs(2110));
    outputs(2899) <= (layer8_outputs(1853)) xor (layer8_outputs(780));
    outputs(2900) <= not(layer8_outputs(257));
    outputs(2901) <= (layer8_outputs(3143)) and (layer8_outputs(5041));
    outputs(2902) <= layer8_outputs(4896);
    outputs(2903) <= not(layer8_outputs(1436));
    outputs(2904) <= not(layer8_outputs(526));
    outputs(2905) <= not((layer8_outputs(957)) xor (layer8_outputs(4383)));
    outputs(2906) <= layer8_outputs(5019);
    outputs(2907) <= not(layer8_outputs(1520)) or (layer8_outputs(980));
    outputs(2908) <= (layer8_outputs(2099)) xor (layer8_outputs(3677));
    outputs(2909) <= layer8_outputs(1728);
    outputs(2910) <= not((layer8_outputs(2195)) xor (layer8_outputs(538)));
    outputs(2911) <= layer8_outputs(3321);
    outputs(2912) <= layer8_outputs(4187);
    outputs(2913) <= not(layer8_outputs(3692));
    outputs(2914) <= (layer8_outputs(934)) and not (layer8_outputs(2081));
    outputs(2915) <= not(layer8_outputs(3443));
    outputs(2916) <= not((layer8_outputs(2708)) or (layer8_outputs(240)));
    outputs(2917) <= (layer8_outputs(2712)) xor (layer8_outputs(1214));
    outputs(2918) <= not(layer8_outputs(1335));
    outputs(2919) <= not(layer8_outputs(4915));
    outputs(2920) <= not(layer8_outputs(4341));
    outputs(2921) <= (layer8_outputs(4310)) and not (layer8_outputs(4493));
    outputs(2922) <= not((layer8_outputs(3471)) xor (layer8_outputs(4856)));
    outputs(2923) <= (layer8_outputs(2078)) and not (layer8_outputs(3147));
    outputs(2924) <= (layer8_outputs(4637)) and not (layer8_outputs(939));
    outputs(2925) <= not(layer8_outputs(172));
    outputs(2926) <= (layer8_outputs(1096)) xor (layer8_outputs(2363));
    outputs(2927) <= layer8_outputs(1855);
    outputs(2928) <= not(layer8_outputs(4701)) or (layer8_outputs(399));
    outputs(2929) <= not((layer8_outputs(2954)) or (layer8_outputs(4992)));
    outputs(2930) <= not(layer8_outputs(427));
    outputs(2931) <= layer8_outputs(4505);
    outputs(2932) <= (layer8_outputs(4968)) and not (layer8_outputs(486));
    outputs(2933) <= not((layer8_outputs(4207)) xor (layer8_outputs(861)));
    outputs(2934) <= (layer8_outputs(1428)) xor (layer8_outputs(4545));
    outputs(2935) <= layer8_outputs(2178);
    outputs(2936) <= (layer8_outputs(4108)) xor (layer8_outputs(1416));
    outputs(2937) <= (layer8_outputs(3060)) xor (layer8_outputs(3118));
    outputs(2938) <= layer8_outputs(1731);
    outputs(2939) <= layer8_outputs(525);
    outputs(2940) <= not(layer8_outputs(3366));
    outputs(2941) <= not(layer8_outputs(3635));
    outputs(2942) <= not(layer8_outputs(4521));
    outputs(2943) <= not((layer8_outputs(640)) xor (layer8_outputs(3212)));
    outputs(2944) <= (layer8_outputs(189)) and (layer8_outputs(4241));
    outputs(2945) <= (layer8_outputs(267)) xor (layer8_outputs(3446));
    outputs(2946) <= not(layer8_outputs(4762));
    outputs(2947) <= not(layer8_outputs(1176));
    outputs(2948) <= (layer8_outputs(116)) and not (layer8_outputs(4246));
    outputs(2949) <= layer8_outputs(4932);
    outputs(2950) <= not(layer8_outputs(3867));
    outputs(2951) <= not((layer8_outputs(1394)) xor (layer8_outputs(5108)));
    outputs(2952) <= not((layer8_outputs(4818)) xor (layer8_outputs(471)));
    outputs(2953) <= (layer8_outputs(2746)) xor (layer8_outputs(1484));
    outputs(2954) <= layer8_outputs(2650);
    outputs(2955) <= not(layer8_outputs(1392));
    outputs(2956) <= not(layer8_outputs(4955));
    outputs(2957) <= not(layer8_outputs(1967)) or (layer8_outputs(1153));
    outputs(2958) <= (layer8_outputs(1858)) xor (layer8_outputs(586));
    outputs(2959) <= layer8_outputs(1664);
    outputs(2960) <= not(layer8_outputs(260));
    outputs(2961) <= (layer8_outputs(223)) xor (layer8_outputs(2244));
    outputs(2962) <= not(layer8_outputs(2953));
    outputs(2963) <= (layer8_outputs(1722)) and not (layer8_outputs(1997));
    outputs(2964) <= layer8_outputs(4440);
    outputs(2965) <= not((layer8_outputs(4308)) xor (layer8_outputs(3161)));
    outputs(2966) <= not(layer8_outputs(1266));
    outputs(2967) <= not((layer8_outputs(844)) or (layer8_outputs(2291)));
    outputs(2968) <= (layer8_outputs(4162)) xor (layer8_outputs(1913));
    outputs(2969) <= not((layer8_outputs(4245)) and (layer8_outputs(3665)));
    outputs(2970) <= (layer8_outputs(2485)) xor (layer8_outputs(4038));
    outputs(2971) <= (layer8_outputs(2153)) and not (layer8_outputs(1432));
    outputs(2972) <= layer8_outputs(1435);
    outputs(2973) <= not((layer8_outputs(1034)) xor (layer8_outputs(3713)));
    outputs(2974) <= (layer8_outputs(4864)) or (layer8_outputs(2142));
    outputs(2975) <= (layer8_outputs(4115)) xor (layer8_outputs(3059));
    outputs(2976) <= not(layer8_outputs(1989));
    outputs(2977) <= not((layer8_outputs(128)) xor (layer8_outputs(4057)));
    outputs(2978) <= not(layer8_outputs(375));
    outputs(2979) <= not(layer8_outputs(1092));
    outputs(2980) <= not(layer8_outputs(2208));
    outputs(2981) <= not((layer8_outputs(286)) or (layer8_outputs(4534)));
    outputs(2982) <= not((layer8_outputs(3693)) or (layer8_outputs(4835)));
    outputs(2983) <= layer8_outputs(2060);
    outputs(2984) <= layer8_outputs(3014);
    outputs(2985) <= (layer8_outputs(2202)) xor (layer8_outputs(3509));
    outputs(2986) <= not(layer8_outputs(2510)) or (layer8_outputs(4746));
    outputs(2987) <= not(layer8_outputs(875));
    outputs(2988) <= not(layer8_outputs(1572));
    outputs(2989) <= not((layer8_outputs(1156)) xor (layer8_outputs(3392)));
    outputs(2990) <= not(layer8_outputs(4171));
    outputs(2991) <= not(layer8_outputs(669));
    outputs(2992) <= layer8_outputs(1170);
    outputs(2993) <= (layer8_outputs(3958)) xor (layer8_outputs(3528));
    outputs(2994) <= not(layer8_outputs(1190));
    outputs(2995) <= layer8_outputs(2889);
    outputs(2996) <= not((layer8_outputs(78)) or (layer8_outputs(3564)));
    outputs(2997) <= not(layer8_outputs(5032));
    outputs(2998) <= not((layer8_outputs(12)) and (layer8_outputs(663)));
    outputs(2999) <= not(layer8_outputs(1068));
    outputs(3000) <= not((layer8_outputs(1690)) xor (layer8_outputs(1936)));
    outputs(3001) <= not(layer8_outputs(4636));
    outputs(3002) <= (layer8_outputs(401)) xor (layer8_outputs(122));
    outputs(3003) <= layer8_outputs(2251);
    outputs(3004) <= not((layer8_outputs(4360)) xor (layer8_outputs(270)));
    outputs(3005) <= (layer8_outputs(461)) and (layer8_outputs(983));
    outputs(3006) <= not(layer8_outputs(3575));
    outputs(3007) <= not((layer8_outputs(3617)) and (layer8_outputs(2416)));
    outputs(3008) <= not(layer8_outputs(2494));
    outputs(3009) <= layer8_outputs(2212);
    outputs(3010) <= (layer8_outputs(140)) and not (layer8_outputs(2031));
    outputs(3011) <= (layer8_outputs(3546)) xor (layer8_outputs(536));
    outputs(3012) <= (layer8_outputs(1212)) and not (layer8_outputs(226));
    outputs(3013) <= layer8_outputs(4637);
    outputs(3014) <= not(layer8_outputs(4375));
    outputs(3015) <= not(layer8_outputs(888));
    outputs(3016) <= (layer8_outputs(3223)) xor (layer8_outputs(2762));
    outputs(3017) <= not(layer8_outputs(4264));
    outputs(3018) <= (layer8_outputs(3045)) xor (layer8_outputs(2793));
    outputs(3019) <= layer8_outputs(4750);
    outputs(3020) <= not(layer8_outputs(2651)) or (layer8_outputs(3273));
    outputs(3021) <= not(layer8_outputs(3996));
    outputs(3022) <= not(layer8_outputs(4273));
    outputs(3023) <= not(layer8_outputs(4341));
    outputs(3024) <= (layer8_outputs(2249)) and (layer8_outputs(4623));
    outputs(3025) <= layer8_outputs(4871);
    outputs(3026) <= layer8_outputs(597);
    outputs(3027) <= not((layer8_outputs(1367)) xor (layer8_outputs(987)));
    outputs(3028) <= not(layer8_outputs(2254));
    outputs(3029) <= layer8_outputs(1495);
    outputs(3030) <= (layer8_outputs(4704)) or (layer8_outputs(3820));
    outputs(3031) <= not((layer8_outputs(3501)) xor (layer8_outputs(2385)));
    outputs(3032) <= (layer8_outputs(4974)) and (layer8_outputs(1341));
    outputs(3033) <= not((layer8_outputs(2696)) xor (layer8_outputs(2190)));
    outputs(3034) <= layer8_outputs(2880);
    outputs(3035) <= not(layer8_outputs(2130));
    outputs(3036) <= layer8_outputs(4946);
    outputs(3037) <= (layer8_outputs(4797)) xor (layer8_outputs(3952));
    outputs(3038) <= layer8_outputs(1673);
    outputs(3039) <= not(layer8_outputs(1908));
    outputs(3040) <= layer8_outputs(4840);
    outputs(3041) <= (layer8_outputs(2244)) xor (layer8_outputs(4386));
    outputs(3042) <= layer8_outputs(1952);
    outputs(3043) <= not(layer8_outputs(2998));
    outputs(3044) <= not(layer8_outputs(2973));
    outputs(3045) <= layer8_outputs(509);
    outputs(3046) <= not(layer8_outputs(1684));
    outputs(3047) <= not((layer8_outputs(2772)) xor (layer8_outputs(381)));
    outputs(3048) <= (layer8_outputs(2996)) and not (layer8_outputs(3949));
    outputs(3049) <= layer8_outputs(32);
    outputs(3050) <= layer8_outputs(2726);
    outputs(3051) <= not((layer8_outputs(2562)) xor (layer8_outputs(1305)));
    outputs(3052) <= not(layer8_outputs(1518));
    outputs(3053) <= not(layer8_outputs(2108));
    outputs(3054) <= (layer8_outputs(3756)) xor (layer8_outputs(2553));
    outputs(3055) <= layer8_outputs(1174);
    outputs(3056) <= not((layer8_outputs(2669)) xor (layer8_outputs(2596)));
    outputs(3057) <= layer8_outputs(3556);
    outputs(3058) <= not((layer8_outputs(210)) or (layer8_outputs(4157)));
    outputs(3059) <= (layer8_outputs(3403)) xor (layer8_outputs(3656));
    outputs(3060) <= not(layer8_outputs(2217));
    outputs(3061) <= layer8_outputs(4402);
    outputs(3062) <= (layer8_outputs(1101)) xor (layer8_outputs(1964));
    outputs(3063) <= not((layer8_outputs(3336)) xor (layer8_outputs(2997)));
    outputs(3064) <= not(layer8_outputs(832));
    outputs(3065) <= not(layer8_outputs(982));
    outputs(3066) <= not(layer8_outputs(1544));
    outputs(3067) <= not((layer8_outputs(1026)) xor (layer8_outputs(761)));
    outputs(3068) <= not(layer8_outputs(2544));
    outputs(3069) <= layer8_outputs(4808);
    outputs(3070) <= (layer8_outputs(3965)) xor (layer8_outputs(2950));
    outputs(3071) <= not(layer8_outputs(3985));
    outputs(3072) <= (layer8_outputs(2333)) or (layer8_outputs(2890));
    outputs(3073) <= layer8_outputs(3699);
    outputs(3074) <= not(layer8_outputs(3697));
    outputs(3075) <= layer8_outputs(4662);
    outputs(3076) <= layer8_outputs(2503);
    outputs(3077) <= not(layer8_outputs(2101));
    outputs(3078) <= not(layer8_outputs(4863));
    outputs(3079) <= not(layer8_outputs(989));
    outputs(3080) <= not(layer8_outputs(1182));
    outputs(3081) <= layer8_outputs(3651);
    outputs(3082) <= not(layer8_outputs(741));
    outputs(3083) <= not(layer8_outputs(2157));
    outputs(3084) <= (layer8_outputs(4066)) or (layer8_outputs(689));
    outputs(3085) <= layer8_outputs(2917);
    outputs(3086) <= layer8_outputs(1207);
    outputs(3087) <= layer8_outputs(3323);
    outputs(3088) <= not(layer8_outputs(2466)) or (layer8_outputs(3030));
    outputs(3089) <= not(layer8_outputs(2423));
    outputs(3090) <= not(layer8_outputs(3281));
    outputs(3091) <= (layer8_outputs(1614)) and not (layer8_outputs(1301));
    outputs(3092) <= not(layer8_outputs(1920));
    outputs(3093) <= layer8_outputs(1716);
    outputs(3094) <= (layer8_outputs(5024)) and not (layer8_outputs(3613));
    outputs(3095) <= not(layer8_outputs(1273));
    outputs(3096) <= not((layer8_outputs(2497)) xor (layer8_outputs(1552)));
    outputs(3097) <= layer8_outputs(879);
    outputs(3098) <= not(layer8_outputs(3051));
    outputs(3099) <= not(layer8_outputs(2493));
    outputs(3100) <= not(layer8_outputs(1978));
    outputs(3101) <= layer8_outputs(4918);
    outputs(3102) <= not(layer8_outputs(1388));
    outputs(3103) <= not(layer8_outputs(672));
    outputs(3104) <= (layer8_outputs(5043)) xor (layer8_outputs(4021));
    outputs(3105) <= layer8_outputs(4336);
    outputs(3106) <= layer8_outputs(970);
    outputs(3107) <= not(layer8_outputs(3116));
    outputs(3108) <= not(layer8_outputs(3904));
    outputs(3109) <= (layer8_outputs(3716)) and not (layer8_outputs(4950));
    outputs(3110) <= (layer8_outputs(2973)) and not (layer8_outputs(5099));
    outputs(3111) <= layer8_outputs(1960);
    outputs(3112) <= not(layer8_outputs(635));
    outputs(3113) <= layer8_outputs(924);
    outputs(3114) <= (layer8_outputs(4743)) xor (layer8_outputs(1115));
    outputs(3115) <= (layer8_outputs(4428)) xor (layer8_outputs(4330));
    outputs(3116) <= (layer8_outputs(557)) xor (layer8_outputs(2034));
    outputs(3117) <= (layer8_outputs(3673)) and (layer8_outputs(4290));
    outputs(3118) <= not((layer8_outputs(1505)) and (layer8_outputs(13)));
    outputs(3119) <= layer8_outputs(4820);
    outputs(3120) <= not((layer8_outputs(2376)) xor (layer8_outputs(3151)));
    outputs(3121) <= not((layer8_outputs(2247)) xor (layer8_outputs(441)));
    outputs(3122) <= layer8_outputs(1646);
    outputs(3123) <= not(layer8_outputs(3911));
    outputs(3124) <= layer8_outputs(3557);
    outputs(3125) <= not(layer8_outputs(1290));
    outputs(3126) <= not(layer8_outputs(3575));
    outputs(3127) <= not(layer8_outputs(3760));
    outputs(3128) <= (layer8_outputs(1117)) and not (layer8_outputs(2681));
    outputs(3129) <= not(layer8_outputs(3204));
    outputs(3130) <= not(layer8_outputs(3621));
    outputs(3131) <= layer8_outputs(778);
    outputs(3132) <= not(layer8_outputs(4282));
    outputs(3133) <= (layer8_outputs(2033)) and not (layer8_outputs(4690));
    outputs(3134) <= layer8_outputs(3769);
    outputs(3135) <= layer8_outputs(4147);
    outputs(3136) <= layer8_outputs(1093);
    outputs(3137) <= layer8_outputs(2148);
    outputs(3138) <= not((layer8_outputs(5104)) xor (layer8_outputs(107)));
    outputs(3139) <= layer8_outputs(1991);
    outputs(3140) <= layer8_outputs(2171);
    outputs(3141) <= layer8_outputs(1203);
    outputs(3142) <= layer8_outputs(1261);
    outputs(3143) <= not((layer8_outputs(3231)) and (layer8_outputs(3743)));
    outputs(3144) <= not((layer8_outputs(1740)) xor (layer8_outputs(746)));
    outputs(3145) <= not((layer8_outputs(3072)) xor (layer8_outputs(4697)));
    outputs(3146) <= layer8_outputs(2390);
    outputs(3147) <= not(layer8_outputs(242));
    outputs(3148) <= layer8_outputs(1017);
    outputs(3149) <= not(layer8_outputs(3697));
    outputs(3150) <= layer8_outputs(751);
    outputs(3151) <= (layer8_outputs(3592)) and (layer8_outputs(4579));
    outputs(3152) <= not(layer8_outputs(4107));
    outputs(3153) <= not((layer8_outputs(486)) xor (layer8_outputs(711)));
    outputs(3154) <= (layer8_outputs(4741)) and (layer8_outputs(3074));
    outputs(3155) <= not((layer8_outputs(1296)) xor (layer8_outputs(3249)));
    outputs(3156) <= (layer8_outputs(66)) and (layer8_outputs(2853));
    outputs(3157) <= not((layer8_outputs(103)) and (layer8_outputs(1562)));
    outputs(3158) <= not(layer8_outputs(3192));
    outputs(3159) <= not(layer8_outputs(2009));
    outputs(3160) <= layer8_outputs(2454);
    outputs(3161) <= layer8_outputs(544);
    outputs(3162) <= (layer8_outputs(2093)) or (layer8_outputs(4744));
    outputs(3163) <= not(layer8_outputs(2833));
    outputs(3164) <= not(layer8_outputs(1750));
    outputs(3165) <= layer8_outputs(4183);
    outputs(3166) <= (layer8_outputs(4179)) or (layer8_outputs(4168));
    outputs(3167) <= not((layer8_outputs(4823)) or (layer8_outputs(3964)));
    outputs(3168) <= (layer8_outputs(4947)) xor (layer8_outputs(1510));
    outputs(3169) <= layer8_outputs(4658);
    outputs(3170) <= not(layer8_outputs(1332));
    outputs(3171) <= layer8_outputs(1163);
    outputs(3172) <= (layer8_outputs(4717)) xor (layer8_outputs(485));
    outputs(3173) <= not(layer8_outputs(2397));
    outputs(3174) <= not(layer8_outputs(1945));
    outputs(3175) <= not(layer8_outputs(719));
    outputs(3176) <= not(layer8_outputs(32));
    outputs(3177) <= (layer8_outputs(1364)) xor (layer8_outputs(4512));
    outputs(3178) <= not(layer8_outputs(528));
    outputs(3179) <= layer8_outputs(929);
    outputs(3180) <= layer8_outputs(4422);
    outputs(3181) <= not(layer8_outputs(1356));
    outputs(3182) <= not(layer8_outputs(717));
    outputs(3183) <= layer8_outputs(807);
    outputs(3184) <= not(layer8_outputs(4882));
    outputs(3185) <= not(layer8_outputs(2077));
    outputs(3186) <= (layer8_outputs(2041)) xor (layer8_outputs(2482));
    outputs(3187) <= not(layer8_outputs(2698));
    outputs(3188) <= layer8_outputs(189);
    outputs(3189) <= (layer8_outputs(666)) or (layer8_outputs(4406));
    outputs(3190) <= not(layer8_outputs(1682));
    outputs(3191) <= not((layer8_outputs(3292)) xor (layer8_outputs(3175)));
    outputs(3192) <= not((layer8_outputs(4526)) xor (layer8_outputs(360)));
    outputs(3193) <= not(layer8_outputs(1426));
    outputs(3194) <= layer8_outputs(3037);
    outputs(3195) <= not((layer8_outputs(4859)) xor (layer8_outputs(2406)));
    outputs(3196) <= layer8_outputs(1747);
    outputs(3197) <= not((layer8_outputs(3901)) xor (layer8_outputs(1526)));
    outputs(3198) <= not(layer8_outputs(1700));
    outputs(3199) <= (layer8_outputs(2638)) and not (layer8_outputs(3817));
    outputs(3200) <= not(layer8_outputs(3861));
    outputs(3201) <= (layer8_outputs(3633)) xor (layer8_outputs(2483));
    outputs(3202) <= not(layer8_outputs(2375));
    outputs(3203) <= layer8_outputs(1747);
    outputs(3204) <= not(layer8_outputs(365));
    outputs(3205) <= not(layer8_outputs(5083));
    outputs(3206) <= layer8_outputs(2548);
    outputs(3207) <= layer8_outputs(4585);
    outputs(3208) <= layer8_outputs(1547);
    outputs(3209) <= not(layer8_outputs(4943));
    outputs(3210) <= not((layer8_outputs(4998)) and (layer8_outputs(4067)));
    outputs(3211) <= (layer8_outputs(3339)) xor (layer8_outputs(1316));
    outputs(3212) <= not((layer8_outputs(1279)) xor (layer8_outputs(2408)));
    outputs(3213) <= layer8_outputs(4625);
    outputs(3214) <= layer8_outputs(2005);
    outputs(3215) <= not(layer8_outputs(1776));
    outputs(3216) <= not(layer8_outputs(3920));
    outputs(3217) <= not((layer8_outputs(2)) or (layer8_outputs(3681)));
    outputs(3218) <= (layer8_outputs(2377)) and not (layer8_outputs(2761));
    outputs(3219) <= not(layer8_outputs(734));
    outputs(3220) <= not(layer8_outputs(4252)) or (layer8_outputs(382));
    outputs(3221) <= layer8_outputs(2981);
    outputs(3222) <= not(layer8_outputs(2637));
    outputs(3223) <= (layer8_outputs(3497)) and not (layer8_outputs(306));
    outputs(3224) <= layer8_outputs(2437);
    outputs(3225) <= layer8_outputs(4927);
    outputs(3226) <= not(layer8_outputs(2210));
    outputs(3227) <= (layer8_outputs(2519)) xor (layer8_outputs(440));
    outputs(3228) <= not((layer8_outputs(185)) xor (layer8_outputs(4557)));
    outputs(3229) <= not(layer8_outputs(4134));
    outputs(3230) <= not(layer8_outputs(789));
    outputs(3231) <= layer8_outputs(4348);
    outputs(3232) <= not(layer8_outputs(135));
    outputs(3233) <= layer8_outputs(4225);
    outputs(3234) <= layer8_outputs(2740);
    outputs(3235) <= not(layer8_outputs(2539));
    outputs(3236) <= (layer8_outputs(1362)) and not (layer8_outputs(324));
    outputs(3237) <= not((layer8_outputs(2155)) or (layer8_outputs(2175)));
    outputs(3238) <= not(layer8_outputs(1995)) or (layer8_outputs(2673));
    outputs(3239) <= not(layer8_outputs(2443));
    outputs(3240) <= (layer8_outputs(2196)) and (layer8_outputs(1714));
    outputs(3241) <= layer8_outputs(3903);
    outputs(3242) <= not((layer8_outputs(3929)) xor (layer8_outputs(3117)));
    outputs(3243) <= (layer8_outputs(239)) or (layer8_outputs(2890));
    outputs(3244) <= not((layer8_outputs(2628)) xor (layer8_outputs(2891)));
    outputs(3245) <= not((layer8_outputs(985)) xor (layer8_outputs(164)));
    outputs(3246) <= layer8_outputs(1117);
    outputs(3247) <= not(layer8_outputs(2960));
    outputs(3248) <= layer8_outputs(4613);
    outputs(3249) <= layer8_outputs(3);
    outputs(3250) <= not(layer8_outputs(4940));
    outputs(3251) <= not((layer8_outputs(1113)) xor (layer8_outputs(2480)));
    outputs(3252) <= (layer8_outputs(620)) xor (layer8_outputs(1312));
    outputs(3253) <= layer8_outputs(2412);
    outputs(3254) <= (layer8_outputs(3630)) xor (layer8_outputs(149));
    outputs(3255) <= not(layer8_outputs(112));
    outputs(3256) <= not(layer8_outputs(1256));
    outputs(3257) <= layer8_outputs(1179);
    outputs(3258) <= not(layer8_outputs(2700));
    outputs(3259) <= layer8_outputs(2142);
    outputs(3260) <= (layer8_outputs(87)) and not (layer8_outputs(162));
    outputs(3261) <= not((layer8_outputs(2821)) xor (layer8_outputs(3591)));
    outputs(3262) <= layer8_outputs(897);
    outputs(3263) <= not(layer8_outputs(5048));
    outputs(3264) <= layer8_outputs(1816);
    outputs(3265) <= not(layer8_outputs(3921));
    outputs(3266) <= not((layer8_outputs(2999)) or (layer8_outputs(4384)));
    outputs(3267) <= layer8_outputs(2170);
    outputs(3268) <= (layer8_outputs(1665)) and (layer8_outputs(4938));
    outputs(3269) <= not((layer8_outputs(3973)) or (layer8_outputs(488)));
    outputs(3270) <= (layer8_outputs(1754)) and not (layer8_outputs(3544));
    outputs(3271) <= not((layer8_outputs(4131)) xor (layer8_outputs(1144)));
    outputs(3272) <= layer8_outputs(4126);
    outputs(3273) <= layer8_outputs(2501);
    outputs(3274) <= layer8_outputs(4034);
    outputs(3275) <= not(layer8_outputs(2178));
    outputs(3276) <= layer8_outputs(4667);
    outputs(3277) <= not(layer8_outputs(2153));
    outputs(3278) <= layer8_outputs(2781);
    outputs(3279) <= layer8_outputs(3710);
    outputs(3280) <= layer8_outputs(1185);
    outputs(3281) <= not(layer8_outputs(2901));
    outputs(3282) <= not((layer8_outputs(858)) xor (layer8_outputs(1678)));
    outputs(3283) <= not(layer8_outputs(2751));
    outputs(3284) <= layer8_outputs(1003);
    outputs(3285) <= layer8_outputs(4335);
    outputs(3286) <= not(layer8_outputs(1959));
    outputs(3287) <= layer8_outputs(3519);
    outputs(3288) <= not(layer8_outputs(3113));
    outputs(3289) <= layer8_outputs(3290);
    outputs(3290) <= not(layer8_outputs(3202));
    outputs(3291) <= not(layer8_outputs(4605));
    outputs(3292) <= not(layer8_outputs(3694));
    outputs(3293) <= not(layer8_outputs(1622));
    outputs(3294) <= layer8_outputs(4432);
    outputs(3295) <= not((layer8_outputs(4595)) xor (layer8_outputs(5038)));
    outputs(3296) <= (layer8_outputs(2017)) and not (layer8_outputs(3835));
    outputs(3297) <= layer8_outputs(2690);
    outputs(3298) <= not((layer8_outputs(3320)) and (layer8_outputs(2552)));
    outputs(3299) <= not((layer8_outputs(4671)) or (layer8_outputs(470)));
    outputs(3300) <= not((layer8_outputs(3885)) xor (layer8_outputs(2608)));
    outputs(3301) <= layer8_outputs(4342);
    outputs(3302) <= layer8_outputs(5094);
    outputs(3303) <= not(layer8_outputs(1433));
    outputs(3304) <= layer8_outputs(1141);
    outputs(3305) <= (layer8_outputs(548)) and not (layer8_outputs(2547));
    outputs(3306) <= layer8_outputs(3208);
    outputs(3307) <= not(layer8_outputs(1491));
    outputs(3308) <= layer8_outputs(4435);
    outputs(3309) <= not((layer8_outputs(2366)) or (layer8_outputs(1304)));
    outputs(3310) <= layer8_outputs(2898);
    outputs(3311) <= (layer8_outputs(4488)) xor (layer8_outputs(3252));
    outputs(3312) <= not((layer8_outputs(1569)) xor (layer8_outputs(828)));
    outputs(3313) <= not(layer8_outputs(3049));
    outputs(3314) <= not((layer8_outputs(2039)) xor (layer8_outputs(1311)));
    outputs(3315) <= layer8_outputs(5079);
    outputs(3316) <= layer8_outputs(2138);
    outputs(3317) <= layer8_outputs(4079);
    outputs(3318) <= layer8_outputs(1278);
    outputs(3319) <= not(layer8_outputs(80));
    outputs(3320) <= layer8_outputs(359);
    outputs(3321) <= not(layer8_outputs(1625));
    outputs(3322) <= (layer8_outputs(1366)) xor (layer8_outputs(4286));
    outputs(3323) <= (layer8_outputs(3177)) and (layer8_outputs(2468));
    outputs(3324) <= not(layer8_outputs(2226));
    outputs(3325) <= not(layer8_outputs(3011));
    outputs(3326) <= layer8_outputs(2046);
    outputs(3327) <= layer8_outputs(1911);
    outputs(3328) <= not((layer8_outputs(736)) xor (layer8_outputs(211)));
    outputs(3329) <= not((layer8_outputs(4387)) xor (layer8_outputs(3103)));
    outputs(3330) <= layer8_outputs(1960);
    outputs(3331) <= (layer8_outputs(1782)) and not (layer8_outputs(1828));
    outputs(3332) <= layer8_outputs(3703);
    outputs(3333) <= not(layer8_outputs(2739));
    outputs(3334) <= (layer8_outputs(4372)) xor (layer8_outputs(1929));
    outputs(3335) <= layer8_outputs(3714);
    outputs(3336) <= not(layer8_outputs(4607));
    outputs(3337) <= not(layer8_outputs(5086));
    outputs(3338) <= not(layer8_outputs(1045));
    outputs(3339) <= not(layer8_outputs(2749));
    outputs(3340) <= layer8_outputs(2279);
    outputs(3341) <= layer8_outputs(4840);
    outputs(3342) <= layer8_outputs(2344);
    outputs(3343) <= not(layer8_outputs(4062));
    outputs(3344) <= not(layer8_outputs(1989));
    outputs(3345) <= not(layer8_outputs(3536));
    outputs(3346) <= layer8_outputs(4340);
    outputs(3347) <= (layer8_outputs(709)) and not (layer8_outputs(1111));
    outputs(3348) <= not((layer8_outputs(2669)) xor (layer8_outputs(3005)));
    outputs(3349) <= not(layer8_outputs(50));
    outputs(3350) <= layer8_outputs(3870);
    outputs(3351) <= not(layer8_outputs(3517));
    outputs(3352) <= not((layer8_outputs(1847)) xor (layer8_outputs(2202)));
    outputs(3353) <= layer8_outputs(3530);
    outputs(3354) <= layer8_outputs(386);
    outputs(3355) <= (layer8_outputs(4214)) and (layer8_outputs(2262));
    outputs(3356) <= not(layer8_outputs(183)) or (layer8_outputs(5018));
    outputs(3357) <= not(layer8_outputs(1508)) or (layer8_outputs(765));
    outputs(3358) <= (layer8_outputs(2398)) and not (layer8_outputs(4309));
    outputs(3359) <= not((layer8_outputs(849)) and (layer8_outputs(1385)));
    outputs(3360) <= layer8_outputs(3148);
    outputs(3361) <= not(layer8_outputs(4078));
    outputs(3362) <= not(layer8_outputs(2751));
    outputs(3363) <= not(layer8_outputs(706));
    outputs(3364) <= (layer8_outputs(3288)) xor (layer8_outputs(2942));
    outputs(3365) <= not(layer8_outputs(3599));
    outputs(3366) <= (layer8_outputs(4576)) xor (layer8_outputs(3036));
    outputs(3367) <= (layer8_outputs(4031)) xor (layer8_outputs(2282));
    outputs(3368) <= not(layer8_outputs(3108));
    outputs(3369) <= not((layer8_outputs(2977)) xor (layer8_outputs(1086)));
    outputs(3370) <= not(layer8_outputs(1456));
    outputs(3371) <= not(layer8_outputs(3342));
    outputs(3372) <= (layer8_outputs(4102)) and (layer8_outputs(3481));
    outputs(3373) <= layer8_outputs(2524);
    outputs(3374) <= not(layer8_outputs(2990));
    outputs(3375) <= not(layer8_outputs(1454));
    outputs(3376) <= not((layer8_outputs(2448)) and (layer8_outputs(1122)));
    outputs(3377) <= not(layer8_outputs(4211));
    outputs(3378) <= not(layer8_outputs(1059));
    outputs(3379) <= not((layer8_outputs(679)) xor (layer8_outputs(100)));
    outputs(3380) <= not(layer8_outputs(2749));
    outputs(3381) <= (layer8_outputs(400)) and (layer8_outputs(3889));
    outputs(3382) <= layer8_outputs(3029);
    outputs(3383) <= layer8_outputs(2346);
    outputs(3384) <= layer8_outputs(2864);
    outputs(3385) <= layer8_outputs(2276);
    outputs(3386) <= (layer8_outputs(2988)) and not (layer8_outputs(2281));
    outputs(3387) <= layer8_outputs(3059);
    outputs(3388) <= not(layer8_outputs(2491));
    outputs(3389) <= not((layer8_outputs(1810)) xor (layer8_outputs(2525)));
    outputs(3390) <= not(layer8_outputs(2245)) or (layer8_outputs(4070));
    outputs(3391) <= layer8_outputs(238);
    outputs(3392) <= layer8_outputs(2741);
    outputs(3393) <= (layer8_outputs(5001)) and not (layer8_outputs(4417));
    outputs(3394) <= not((layer8_outputs(2593)) xor (layer8_outputs(86)));
    outputs(3395) <= not(layer8_outputs(1883));
    outputs(3396) <= (layer8_outputs(4692)) xor (layer8_outputs(82));
    outputs(3397) <= layer8_outputs(2381);
    outputs(3398) <= (layer8_outputs(1416)) and not (layer8_outputs(3475));
    outputs(3399) <= layer8_outputs(3741);
    outputs(3400) <= (layer8_outputs(1585)) or (layer8_outputs(1556));
    outputs(3401) <= not(layer8_outputs(2365));
    outputs(3402) <= not((layer8_outputs(4237)) xor (layer8_outputs(2055)));
    outputs(3403) <= not((layer8_outputs(2767)) and (layer8_outputs(4229)));
    outputs(3404) <= layer8_outputs(4058);
    outputs(3405) <= layer8_outputs(3445);
    outputs(3406) <= (layer8_outputs(1783)) and not (layer8_outputs(113));
    outputs(3407) <= (layer8_outputs(4999)) and not (layer8_outputs(2383));
    outputs(3408) <= not((layer8_outputs(755)) xor (layer8_outputs(215)));
    outputs(3409) <= not((layer8_outputs(813)) xor (layer8_outputs(3285)));
    outputs(3410) <= not((layer8_outputs(1798)) or (layer8_outputs(2414)));
    outputs(3411) <= not(layer8_outputs(4539));
    outputs(3412) <= (layer8_outputs(2143)) xor (layer8_outputs(2448));
    outputs(3413) <= layer8_outputs(1239);
    outputs(3414) <= not((layer8_outputs(739)) xor (layer8_outputs(513)));
    outputs(3415) <= not(layer8_outputs(3671));
    outputs(3416) <= layer8_outputs(4625);
    outputs(3417) <= layer8_outputs(4477);
    outputs(3418) <= not(layer8_outputs(2241));
    outputs(3419) <= layer8_outputs(2633);
    outputs(3420) <= not(layer8_outputs(768)) or (layer8_outputs(880));
    outputs(3421) <= layer8_outputs(4390);
    outputs(3422) <= (layer8_outputs(2510)) xor (layer8_outputs(4270));
    outputs(3423) <= not((layer8_outputs(3315)) or (layer8_outputs(4489)));
    outputs(3424) <= layer8_outputs(646);
    outputs(3425) <= layer8_outputs(2710);
    outputs(3426) <= not(layer8_outputs(1166));
    outputs(3427) <= not(layer8_outputs(3061));
    outputs(3428) <= not((layer8_outputs(428)) xor (layer8_outputs(4553)));
    outputs(3429) <= not(layer8_outputs(4473));
    outputs(3430) <= layer8_outputs(3229);
    outputs(3431) <= not(layer8_outputs(1713));
    outputs(3432) <= not((layer8_outputs(1647)) xor (layer8_outputs(3130)));
    outputs(3433) <= (layer8_outputs(2355)) xor (layer8_outputs(403));
    outputs(3434) <= not(layer8_outputs(908));
    outputs(3435) <= not(layer8_outputs(115));
    outputs(3436) <= layer8_outputs(2191);
    outputs(3437) <= layer8_outputs(4137);
    outputs(3438) <= (layer8_outputs(368)) xor (layer8_outputs(1935));
    outputs(3439) <= not(layer8_outputs(2405));
    outputs(3440) <= not(layer8_outputs(1861));
    outputs(3441) <= not(layer8_outputs(3933));
    outputs(3442) <= not(layer8_outputs(3081));
    outputs(3443) <= not(layer8_outputs(4582));
    outputs(3444) <= (layer8_outputs(1065)) xor (layer8_outputs(3037));
    outputs(3445) <= not(layer8_outputs(4249));
    outputs(3446) <= not(layer8_outputs(2612));
    outputs(3447) <= (layer8_outputs(1173)) xor (layer8_outputs(4554));
    outputs(3448) <= not(layer8_outputs(1934));
    outputs(3449) <= layer8_outputs(1170);
    outputs(3450) <= layer8_outputs(4294);
    outputs(3451) <= not(layer8_outputs(3807));
    outputs(3452) <= not((layer8_outputs(3815)) xor (layer8_outputs(4588)));
    outputs(3453) <= not(layer8_outputs(214));
    outputs(3454) <= not((layer8_outputs(4092)) xor (layer8_outputs(367)));
    outputs(3455) <= not(layer8_outputs(908));
    outputs(3456) <= (layer8_outputs(738)) and not (layer8_outputs(4569));
    outputs(3457) <= (layer8_outputs(3137)) xor (layer8_outputs(4510));
    outputs(3458) <= layer8_outputs(4564);
    outputs(3459) <= layer8_outputs(3374);
    outputs(3460) <= (layer8_outputs(1301)) xor (layer8_outputs(1914));
    outputs(3461) <= not(layer8_outputs(3114));
    outputs(3462) <= (layer8_outputs(224)) xor (layer8_outputs(4916));
    outputs(3463) <= (layer8_outputs(157)) xor (layer8_outputs(1942));
    outputs(3464) <= layer8_outputs(675);
    outputs(3465) <= not((layer8_outputs(3345)) xor (layer8_outputs(4520)));
    outputs(3466) <= (layer8_outputs(3783)) xor (layer8_outputs(4859));
    outputs(3467) <= not((layer8_outputs(4287)) xor (layer8_outputs(3176)));
    outputs(3468) <= layer8_outputs(4604);
    outputs(3469) <= not(layer8_outputs(2004));
    outputs(3470) <= (layer8_outputs(3766)) xor (layer8_outputs(520));
    outputs(3471) <= layer8_outputs(1850);
    outputs(3472) <= not(layer8_outputs(3778));
    outputs(3473) <= not((layer8_outputs(328)) xor (layer8_outputs(3887)));
    outputs(3474) <= not(layer8_outputs(1842));
    outputs(3475) <= not(layer8_outputs(791));
    outputs(3476) <= not((layer8_outputs(4240)) xor (layer8_outputs(3844)));
    outputs(3477) <= layer8_outputs(2649);
    outputs(3478) <= not(layer8_outputs(2769));
    outputs(3479) <= layer8_outputs(5020);
    outputs(3480) <= not(layer8_outputs(1222));
    outputs(3481) <= (layer8_outputs(2134)) xor (layer8_outputs(3188));
    outputs(3482) <= (layer8_outputs(3448)) xor (layer8_outputs(3797));
    outputs(3483) <= not(layer8_outputs(2263));
    outputs(3484) <= not((layer8_outputs(1695)) xor (layer8_outputs(1334)));
    outputs(3485) <= layer8_outputs(4665);
    outputs(3486) <= (layer8_outputs(4424)) xor (layer8_outputs(4438));
    outputs(3487) <= not((layer8_outputs(1119)) xor (layer8_outputs(4826)));
    outputs(3488) <= layer8_outputs(2206);
    outputs(3489) <= not(layer8_outputs(2271));
    outputs(3490) <= (layer8_outputs(3780)) xor (layer8_outputs(2228));
    outputs(3491) <= not(layer8_outputs(2869));
    outputs(3492) <= not((layer8_outputs(4643)) xor (layer8_outputs(808)));
    outputs(3493) <= not(layer8_outputs(4854));
    outputs(3494) <= not(layer8_outputs(1625));
    outputs(3495) <= not(layer8_outputs(523));
    outputs(3496) <= not(layer8_outputs(668));
    outputs(3497) <= (layer8_outputs(1639)) and not (layer8_outputs(1673));
    outputs(3498) <= layer8_outputs(2205);
    outputs(3499) <= not(layer8_outputs(2627));
    outputs(3500) <= layer8_outputs(3167);
    outputs(3501) <= not(layer8_outputs(2287));
    outputs(3502) <= not(layer8_outputs(3904));
    outputs(3503) <= not(layer8_outputs(3869));
    outputs(3504) <= layer8_outputs(3152);
    outputs(3505) <= layer8_outputs(879);
    outputs(3506) <= (layer8_outputs(4583)) xor (layer8_outputs(3352));
    outputs(3507) <= layer8_outputs(2557);
    outputs(3508) <= layer8_outputs(4222);
    outputs(3509) <= (layer8_outputs(2387)) xor (layer8_outputs(1534));
    outputs(3510) <= not((layer8_outputs(4205)) xor (layer8_outputs(2725)));
    outputs(3511) <= layer8_outputs(744);
    outputs(3512) <= not(layer8_outputs(4125));
    outputs(3513) <= not(layer8_outputs(4048));
    outputs(3514) <= (layer8_outputs(1694)) xor (layer8_outputs(2540));
    outputs(3515) <= not(layer8_outputs(3121));
    outputs(3516) <= layer8_outputs(2824);
    outputs(3517) <= layer8_outputs(2076);
    outputs(3518) <= not(layer8_outputs(49));
    outputs(3519) <= (layer8_outputs(2814)) xor (layer8_outputs(3586));
    outputs(3520) <= (layer8_outputs(1372)) xor (layer8_outputs(3977));
    outputs(3521) <= not(layer8_outputs(3816));
    outputs(3522) <= layer8_outputs(2799);
    outputs(3523) <= not(layer8_outputs(4527));
    outputs(3524) <= not(layer8_outputs(234));
    outputs(3525) <= not(layer8_outputs(1880));
    outputs(3526) <= layer8_outputs(1404);
    outputs(3527) <= layer8_outputs(5070);
    outputs(3528) <= (layer8_outputs(1320)) xor (layer8_outputs(3897));
    outputs(3529) <= not(layer8_outputs(142));
    outputs(3530) <= layer8_outputs(3218);
    outputs(3531) <= not((layer8_outputs(4282)) or (layer8_outputs(2807)));
    outputs(3532) <= not((layer8_outputs(4663)) xor (layer8_outputs(2379)));
    outputs(3533) <= not(layer8_outputs(1405));
    outputs(3534) <= layer8_outputs(1364);
    outputs(3535) <= not(layer8_outputs(527));
    outputs(3536) <= layer8_outputs(2164);
    outputs(3537) <= layer8_outputs(126);
    outputs(3538) <= (layer8_outputs(2321)) xor (layer8_outputs(1551));
    outputs(3539) <= not((layer8_outputs(4982)) xor (layer8_outputs(237)));
    outputs(3540) <= layer8_outputs(678);
    outputs(3541) <= not(layer8_outputs(4914)) or (layer8_outputs(2382));
    outputs(3542) <= not(layer8_outputs(3590));
    outputs(3543) <= layer8_outputs(3126);
    outputs(3544) <= (layer8_outputs(2118)) xor (layer8_outputs(4175));
    outputs(3545) <= (layer8_outputs(342)) xor (layer8_outputs(1011));
    outputs(3546) <= (layer8_outputs(1888)) or (layer8_outputs(2652));
    outputs(3547) <= layer8_outputs(152);
    outputs(3548) <= not(layer8_outputs(199));
    outputs(3549) <= layer8_outputs(3258);
    outputs(3550) <= (layer8_outputs(1180)) xor (layer8_outputs(2359));
    outputs(3551) <= (layer8_outputs(2975)) and not (layer8_outputs(4221));
    outputs(3552) <= not(layer8_outputs(4065));
    outputs(3553) <= layer8_outputs(725);
    outputs(3554) <= not(layer8_outputs(1298));
    outputs(3555) <= (layer8_outputs(2152)) or (layer8_outputs(1327));
    outputs(3556) <= layer8_outputs(2721);
    outputs(3557) <= layer8_outputs(384);
    outputs(3558) <= layer8_outputs(2290);
    outputs(3559) <= layer8_outputs(969);
    outputs(3560) <= layer8_outputs(232);
    outputs(3561) <= (layer8_outputs(3307)) xor (layer8_outputs(2907));
    outputs(3562) <= layer8_outputs(1181);
    outputs(3563) <= not((layer8_outputs(4844)) and (layer8_outputs(4114)));
    outputs(3564) <= not(layer8_outputs(1852));
    outputs(3565) <= layer8_outputs(3074);
    outputs(3566) <= not(layer8_outputs(723));
    outputs(3567) <= not(layer8_outputs(3569));
    outputs(3568) <= not((layer8_outputs(2504)) xor (layer8_outputs(4485)));
    outputs(3569) <= (layer8_outputs(3369)) and not (layer8_outputs(1704));
    outputs(3570) <= not((layer8_outputs(4389)) xor (layer8_outputs(3094)));
    outputs(3571) <= layer8_outputs(4334);
    outputs(3572) <= (layer8_outputs(4832)) xor (layer8_outputs(991));
    outputs(3573) <= layer8_outputs(2882);
    outputs(3574) <= layer8_outputs(1655);
    outputs(3575) <= layer8_outputs(4917);
    outputs(3576) <= not(layer8_outputs(3082));
    outputs(3577) <= not(layer8_outputs(989));
    outputs(3578) <= not(layer8_outputs(4623));
    outputs(3579) <= layer8_outputs(2841);
    outputs(3580) <= (layer8_outputs(1446)) and (layer8_outputs(4336));
    outputs(3581) <= layer8_outputs(4730);
    outputs(3582) <= (layer8_outputs(1590)) xor (layer8_outputs(535));
    outputs(3583) <= (layer8_outputs(4459)) xor (layer8_outputs(2349));
    outputs(3584) <= (layer8_outputs(996)) xor (layer8_outputs(3793));
    outputs(3585) <= not((layer8_outputs(2747)) xor (layer8_outputs(3423)));
    outputs(3586) <= layer8_outputs(5087);
    outputs(3587) <= not(layer8_outputs(1022));
    outputs(3588) <= (layer8_outputs(4098)) xor (layer8_outputs(1180));
    outputs(3589) <= (layer8_outputs(3798)) xor (layer8_outputs(4399));
    outputs(3590) <= not((layer8_outputs(597)) xor (layer8_outputs(2250)));
    outputs(3591) <= not((layer8_outputs(1732)) or (layer8_outputs(4304)));
    outputs(3592) <= layer8_outputs(4734);
    outputs(3593) <= layer8_outputs(4519);
    outputs(3594) <= (layer8_outputs(2273)) xor (layer8_outputs(402));
    outputs(3595) <= (layer8_outputs(4222)) xor (layer8_outputs(4682));
    outputs(3596) <= not((layer8_outputs(3587)) xor (layer8_outputs(753)));
    outputs(3597) <= layer8_outputs(1267);
    outputs(3598) <= not((layer8_outputs(3627)) xor (layer8_outputs(3658)));
    outputs(3599) <= (layer8_outputs(2546)) xor (layer8_outputs(4978));
    outputs(3600) <= (layer8_outputs(5005)) xor (layer8_outputs(1805));
    outputs(3601) <= not(layer8_outputs(3208));
    outputs(3602) <= not(layer8_outputs(3447));
    outputs(3603) <= not(layer8_outputs(3787));
    outputs(3604) <= not(layer8_outputs(1616));
    outputs(3605) <= not(layer8_outputs(3530));
    outputs(3606) <= not(layer8_outputs(1055)) or (layer8_outputs(3732));
    outputs(3607) <= not(layer8_outputs(3700));
    outputs(3608) <= layer8_outputs(2502);
    outputs(3609) <= not(layer8_outputs(4919));
    outputs(3610) <= not((layer8_outputs(3909)) or (layer8_outputs(4567)));
    outputs(3611) <= layer8_outputs(1578);
    outputs(3612) <= not((layer8_outputs(3772)) or (layer8_outputs(3573)));
    outputs(3613) <= layer8_outputs(3748);
    outputs(3614) <= not(layer8_outputs(416));
    outputs(3615) <= not(layer8_outputs(3777));
    outputs(3616) <= not(layer8_outputs(2088));
    outputs(3617) <= not(layer8_outputs(4471));
    outputs(3618) <= (layer8_outputs(3245)) and not (layer8_outputs(4567));
    outputs(3619) <= (layer8_outputs(333)) xor (layer8_outputs(1567));
    outputs(3620) <= (layer8_outputs(2518)) and (layer8_outputs(3145));
    outputs(3621) <= not(layer8_outputs(1917));
    outputs(3622) <= layer8_outputs(2073);
    outputs(3623) <= not(layer8_outputs(612));
    outputs(3624) <= not(layer8_outputs(369));
    outputs(3625) <= (layer8_outputs(4880)) and not (layer8_outputs(915));
    outputs(3626) <= (layer8_outputs(79)) xor (layer8_outputs(3554));
    outputs(3627) <= layer8_outputs(3696);
    outputs(3628) <= (layer8_outputs(4852)) and not (layer8_outputs(4608));
    outputs(3629) <= layer8_outputs(4862);
    outputs(3630) <= (layer8_outputs(3439)) and not (layer8_outputs(4760));
    outputs(3631) <= (layer8_outputs(1831)) xor (layer8_outputs(3420));
    outputs(3632) <= layer8_outputs(2706);
    outputs(3633) <= not((layer8_outputs(2184)) xor (layer8_outputs(4858)));
    outputs(3634) <= not((layer8_outputs(2886)) or (layer8_outputs(4213)));
    outputs(3635) <= layer8_outputs(2451);
    outputs(3636) <= not((layer8_outputs(65)) xor (layer8_outputs(1038)));
    outputs(3637) <= (layer8_outputs(3593)) xor (layer8_outputs(4514));
    outputs(3638) <= not(layer8_outputs(209));
    outputs(3639) <= (layer8_outputs(1756)) and not (layer8_outputs(4239));
    outputs(3640) <= not(layer8_outputs(1952));
    outputs(3641) <= not((layer8_outputs(1429)) xor (layer8_outputs(576)));
    outputs(3642) <= not((layer8_outputs(1412)) xor (layer8_outputs(2010)));
    outputs(3643) <= not(layer8_outputs(2345));
    outputs(3644) <= (layer8_outputs(4617)) xor (layer8_outputs(642));
    outputs(3645) <= not(layer8_outputs(3584));
    outputs(3646) <= (layer8_outputs(99)) and not (layer8_outputs(3611));
    outputs(3647) <= (layer8_outputs(270)) and not (layer8_outputs(3484));
    outputs(3648) <= not(layer8_outputs(1733));
    outputs(3649) <= layer8_outputs(2990);
    outputs(3650) <= not((layer8_outputs(3708)) xor (layer8_outputs(5101)));
    outputs(3651) <= layer8_outputs(3326);
    outputs(3652) <= not((layer8_outputs(1773)) xor (layer8_outputs(3207)));
    outputs(3653) <= not(layer8_outputs(2931)) or (layer8_outputs(3414));
    outputs(3654) <= not(layer8_outputs(3153));
    outputs(3655) <= (layer8_outputs(2734)) or (layer8_outputs(2607));
    outputs(3656) <= layer8_outputs(4019);
    outputs(3657) <= (layer8_outputs(3098)) xor (layer8_outputs(4664));
    outputs(3658) <= layer8_outputs(1619);
    outputs(3659) <= not(layer8_outputs(4964));
    outputs(3660) <= not((layer8_outputs(4498)) xor (layer8_outputs(3740)));
    outputs(3661) <= layer8_outputs(3645);
    outputs(3662) <= not((layer8_outputs(3835)) xor (layer8_outputs(867)));
    outputs(3663) <= not(layer8_outputs(1179));
    outputs(3664) <= not(layer8_outputs(439));
    outputs(3665) <= not((layer8_outputs(4592)) xor (layer8_outputs(2969)));
    outputs(3666) <= layer8_outputs(4296);
    outputs(3667) <= (layer8_outputs(2580)) and not (layer8_outputs(4263));
    outputs(3668) <= (layer8_outputs(1242)) or (layer8_outputs(580));
    outputs(3669) <= layer8_outputs(4942);
    outputs(3670) <= (layer8_outputs(4420)) xor (layer8_outputs(148));
    outputs(3671) <= layer8_outputs(890);
    outputs(3672) <= (layer8_outputs(4939)) xor (layer8_outputs(1709));
    outputs(3673) <= (layer8_outputs(2192)) xor (layer8_outputs(1904));
    outputs(3674) <= (layer8_outputs(4681)) xor (layer8_outputs(4796));
    outputs(3675) <= (layer8_outputs(4653)) xor (layer8_outputs(200));
    outputs(3676) <= not((layer8_outputs(552)) xor (layer8_outputs(3450)));
    outputs(3677) <= not(layer8_outputs(3272));
    outputs(3678) <= not(layer8_outputs(4913));
    outputs(3679) <= not((layer8_outputs(3215)) or (layer8_outputs(2361)));
    outputs(3680) <= not(layer8_outputs(4113));
    outputs(3681) <= not((layer8_outputs(4725)) or (layer8_outputs(1286)));
    outputs(3682) <= not(layer8_outputs(2233));
    outputs(3683) <= layer8_outputs(2855);
    outputs(3684) <= not((layer8_outputs(60)) xor (layer8_outputs(621)));
    outputs(3685) <= (layer8_outputs(1013)) xor (layer8_outputs(463));
    outputs(3686) <= not(layer8_outputs(1650));
    outputs(3687) <= (layer8_outputs(4501)) xor (layer8_outputs(48));
    outputs(3688) <= layer8_outputs(1859);
    outputs(3689) <= not((layer8_outputs(4220)) or (layer8_outputs(3299)));
    outputs(3690) <= layer8_outputs(2065);
    outputs(3691) <= not((layer8_outputs(465)) xor (layer8_outputs(846)));
    outputs(3692) <= layer8_outputs(3110);
    outputs(3693) <= layer8_outputs(2902);
    outputs(3694) <= layer8_outputs(3948);
    outputs(3695) <= not((layer8_outputs(3525)) xor (layer8_outputs(1415)));
    outputs(3696) <= not(layer8_outputs(1634));
    outputs(3697) <= layer8_outputs(3545);
    outputs(3698) <= not(layer8_outputs(2896));
    outputs(3699) <= not(layer8_outputs(2133));
    outputs(3700) <= not(layer8_outputs(170));
    outputs(3701) <= (layer8_outputs(876)) xor (layer8_outputs(163));
    outputs(3702) <= not(layer8_outputs(3993));
    outputs(3703) <= not(layer8_outputs(3481));
    outputs(3704) <= (layer8_outputs(1415)) xor (layer8_outputs(3396));
    outputs(3705) <= layer8_outputs(946);
    outputs(3706) <= (layer8_outputs(1380)) and not (layer8_outputs(3856));
    outputs(3707) <= not((layer8_outputs(167)) or (layer8_outputs(359)));
    outputs(3708) <= not(layer8_outputs(1138));
    outputs(3709) <= not(layer8_outputs(3302));
    outputs(3710) <= not(layer8_outputs(972));
    outputs(3711) <= layer8_outputs(3375);
    outputs(3712) <= (layer8_outputs(2550)) and not (layer8_outputs(874));
    outputs(3713) <= not((layer8_outputs(4326)) xor (layer8_outputs(4075)));
    outputs(3714) <= layer8_outputs(932);
    outputs(3715) <= (layer8_outputs(2658)) xor (layer8_outputs(4116));
    outputs(3716) <= (layer8_outputs(4542)) or (layer8_outputs(651));
    outputs(3717) <= layer8_outputs(4693);
    outputs(3718) <= (layer8_outputs(3149)) and (layer8_outputs(457));
    outputs(3719) <= layer8_outputs(3925);
    outputs(3720) <= (layer8_outputs(1125)) xor (layer8_outputs(147));
    outputs(3721) <= layer8_outputs(3539);
    outputs(3722) <= (layer8_outputs(1344)) and not (layer8_outputs(2248));
    outputs(3723) <= not(layer8_outputs(414)) or (layer8_outputs(3752));
    outputs(3724) <= not((layer8_outputs(3771)) xor (layer8_outputs(4836)));
    outputs(3725) <= (layer8_outputs(4275)) xor (layer8_outputs(1167));
    outputs(3726) <= not(layer8_outputs(4686));
    outputs(3727) <= not(layer8_outputs(3424));
    outputs(3728) <= layer8_outputs(4010);
    outputs(3729) <= layer8_outputs(88);
    outputs(3730) <= (layer8_outputs(585)) xor (layer8_outputs(3421));
    outputs(3731) <= not(layer8_outputs(2415));
    outputs(3732) <= layer8_outputs(4188);
    outputs(3733) <= not(layer8_outputs(4460));
    outputs(3734) <= not(layer8_outputs(2372));
    outputs(3735) <= not((layer8_outputs(2969)) xor (layer8_outputs(474)));
    outputs(3736) <= (layer8_outputs(4110)) xor (layer8_outputs(2676));
    outputs(3737) <= not(layer8_outputs(4990));
    outputs(3738) <= (layer8_outputs(4669)) and (layer8_outputs(2293));
    outputs(3739) <= (layer8_outputs(3612)) xor (layer8_outputs(4226));
    outputs(3740) <= not((layer8_outputs(4861)) xor (layer8_outputs(5047)));
    outputs(3741) <= layer8_outputs(2558);
    outputs(3742) <= not((layer8_outputs(160)) xor (layer8_outputs(158)));
    outputs(3743) <= not(layer8_outputs(1733));
    outputs(3744) <= not(layer8_outputs(1203));
    outputs(3745) <= layer8_outputs(4444);
    outputs(3746) <= not(layer8_outputs(797));
    outputs(3747) <= not(layer8_outputs(2635));
    outputs(3748) <= (layer8_outputs(4121)) xor (layer8_outputs(1422));
    outputs(3749) <= not(layer8_outputs(4694));
    outputs(3750) <= layer8_outputs(104);
    outputs(3751) <= not(layer8_outputs(4662));
    outputs(3752) <= (layer8_outputs(243)) xor (layer8_outputs(1946));
    outputs(3753) <= layer8_outputs(4539);
    outputs(3754) <= (layer8_outputs(848)) and not (layer8_outputs(295));
    outputs(3755) <= not((layer8_outputs(2887)) xor (layer8_outputs(3522)));
    outputs(3756) <= layer8_outputs(3543);
    outputs(3757) <= not((layer8_outputs(3966)) xor (layer8_outputs(126)));
    outputs(3758) <= not(layer8_outputs(2917));
    outputs(3759) <= not(layer8_outputs(3510));
    outputs(3760) <= layer8_outputs(3448);
    outputs(3761) <= layer8_outputs(3495);
    outputs(3762) <= not(layer8_outputs(3870));
    outputs(3763) <= not((layer8_outputs(119)) xor (layer8_outputs(35)));
    outputs(3764) <= (layer8_outputs(387)) xor (layer8_outputs(1006));
    outputs(3765) <= (layer8_outputs(3237)) xor (layer8_outputs(1923));
    outputs(3766) <= layer8_outputs(2924);
    outputs(3767) <= not(layer8_outputs(1493));
    outputs(3768) <= not(layer8_outputs(5025));
    outputs(3769) <= (layer8_outputs(2314)) xor (layer8_outputs(4998));
    outputs(3770) <= layer8_outputs(5023);
    outputs(3771) <= (layer8_outputs(1029)) and not (layer8_outputs(2109));
    outputs(3772) <= not((layer8_outputs(3168)) xor (layer8_outputs(1351)));
    outputs(3773) <= (layer8_outputs(2636)) xor (layer8_outputs(654));
    outputs(3774) <= not(layer8_outputs(3124));
    outputs(3775) <= (layer8_outputs(2573)) xor (layer8_outputs(2922));
    outputs(3776) <= layer8_outputs(4844);
    outputs(3777) <= not((layer8_outputs(2136)) xor (layer8_outputs(1540)));
    outputs(3778) <= (layer8_outputs(2303)) xor (layer8_outputs(3275));
    outputs(3779) <= (layer8_outputs(3139)) xor (layer8_outputs(2587));
    outputs(3780) <= not((layer8_outputs(1407)) xor (layer8_outputs(4114)));
    outputs(3781) <= not(layer8_outputs(2849));
    outputs(3782) <= not((layer8_outputs(4644)) xor (layer8_outputs(3056)));
    outputs(3783) <= not((layer8_outputs(733)) xor (layer8_outputs(2111)));
    outputs(3784) <= not(layer8_outputs(156));
    outputs(3785) <= not(layer8_outputs(1748));
    outputs(3786) <= layer8_outputs(2469);
    outputs(3787) <= not((layer8_outputs(4640)) xor (layer8_outputs(3523)));
    outputs(3788) <= (layer8_outputs(1464)) xor (layer8_outputs(2631));
    outputs(3789) <= not((layer8_outputs(2965)) xor (layer8_outputs(2827)));
    outputs(3790) <= not((layer8_outputs(2528)) xor (layer8_outputs(3302)));
    outputs(3791) <= layer8_outputs(1248);
    outputs(3792) <= not((layer8_outputs(343)) xor (layer8_outputs(542)));
    outputs(3793) <= not(layer8_outputs(46));
    outputs(3794) <= layer8_outputs(1982);
    outputs(3795) <= not(layer8_outputs(5030));
    outputs(3796) <= not(layer8_outputs(13)) or (layer8_outputs(1958));
    outputs(3797) <= not((layer8_outputs(1210)) xor (layer8_outputs(2139)));
    outputs(3798) <= not((layer8_outputs(1979)) xor (layer8_outputs(3361)));
    outputs(3799) <= not(layer8_outputs(4073));
    outputs(3800) <= not(layer8_outputs(2388));
    outputs(3801) <= layer8_outputs(4419);
    outputs(3802) <= not(layer8_outputs(2836));
    outputs(3803) <= layer8_outputs(1884);
    outputs(3804) <= not((layer8_outputs(3155)) xor (layer8_outputs(1912)));
    outputs(3805) <= not((layer8_outputs(2377)) and (layer8_outputs(2490)));
    outputs(3806) <= not(layer8_outputs(3316));
    outputs(3807) <= not(layer8_outputs(3136));
    outputs(3808) <= not(layer8_outputs(5114));
    outputs(3809) <= not((layer8_outputs(3514)) xor (layer8_outputs(1902)));
    outputs(3810) <= not((layer8_outputs(1898)) or (layer8_outputs(3628)));
    outputs(3811) <= layer8_outputs(3937);
    outputs(3812) <= (layer8_outputs(2888)) xor (layer8_outputs(832));
    outputs(3813) <= (layer8_outputs(3589)) xor (layer8_outputs(2308));
    outputs(3814) <= (layer8_outputs(3948)) and not (layer8_outputs(294));
    outputs(3815) <= layer8_outputs(3245);
    outputs(3816) <= not(layer8_outputs(2603));
    outputs(3817) <= layer8_outputs(3358);
    outputs(3818) <= not(layer8_outputs(1089));
    outputs(3819) <= layer8_outputs(4621);
    outputs(3820) <= (layer8_outputs(472)) xor (layer8_outputs(2933));
    outputs(3821) <= (layer8_outputs(1985)) xor (layer8_outputs(4774));
    outputs(3822) <= (layer8_outputs(3112)) xor (layer8_outputs(2693));
    outputs(3823) <= not(layer8_outputs(2407));
    outputs(3824) <= (layer8_outputs(4247)) and not (layer8_outputs(4494));
    outputs(3825) <= (layer8_outputs(2967)) xor (layer8_outputs(3625));
    outputs(3826) <= (layer8_outputs(840)) xor (layer8_outputs(3607));
    outputs(3827) <= (layer8_outputs(2842)) and not (layer8_outputs(2808));
    outputs(3828) <= not(layer8_outputs(3896));
    outputs(3829) <= not((layer8_outputs(3411)) or (layer8_outputs(158)));
    outputs(3830) <= (layer8_outputs(1452)) and (layer8_outputs(799));
    outputs(3831) <= (layer8_outputs(684)) and not (layer8_outputs(1965));
    outputs(3832) <= (layer8_outputs(1516)) xor (layer8_outputs(2144));
    outputs(3833) <= layer8_outputs(1266);
    outputs(3834) <= not(layer8_outputs(883));
    outputs(3835) <= not(layer8_outputs(2181));
    outputs(3836) <= not(layer8_outputs(709));
    outputs(3837) <= layer8_outputs(3532);
    outputs(3838) <= not(layer8_outputs(81));
    outputs(3839) <= (layer8_outputs(1491)) and (layer8_outputs(2599));
    outputs(3840) <= layer8_outputs(2728);
    outputs(3841) <= layer8_outputs(1758);
    outputs(3842) <= (layer8_outputs(2371)) and not (layer8_outputs(648));
    outputs(3843) <= not(layer8_outputs(2556)) or (layer8_outputs(918));
    outputs(3844) <= not(layer8_outputs(339));
    outputs(3845) <= not(layer8_outputs(447));
    outputs(3846) <= not((layer8_outputs(2127)) xor (layer8_outputs(1701)));
    outputs(3847) <= not((layer8_outputs(174)) xor (layer8_outputs(2855)));
    outputs(3848) <= (layer8_outputs(4659)) xor (layer8_outputs(1743));
    outputs(3849) <= not((layer8_outputs(2329)) xor (layer8_outputs(1522)));
    outputs(3850) <= layer8_outputs(4043);
    outputs(3851) <= (layer8_outputs(2203)) xor (layer8_outputs(4757));
    outputs(3852) <= not(layer8_outputs(864));
    outputs(3853) <= not(layer8_outputs(401));
    outputs(3854) <= layer8_outputs(4005);
    outputs(3855) <= not(layer8_outputs(2011));
    outputs(3856) <= not((layer8_outputs(4240)) xor (layer8_outputs(3650)));
    outputs(3857) <= layer8_outputs(59);
    outputs(3858) <= not((layer8_outputs(3775)) xor (layer8_outputs(2928)));
    outputs(3859) <= not(layer8_outputs(2686));
    outputs(3860) <= (layer8_outputs(380)) and not (layer8_outputs(2529));
    outputs(3861) <= layer8_outputs(2145);
    outputs(3862) <= not(layer8_outputs(2021));
    outputs(3863) <= (layer8_outputs(438)) xor (layer8_outputs(2585));
    outputs(3864) <= not(layer8_outputs(1992));
    outputs(3865) <= not(layer8_outputs(3092));
    outputs(3866) <= (layer8_outputs(2940)) xor (layer8_outputs(698));
    outputs(3867) <= (layer8_outputs(2577)) and not (layer8_outputs(73));
    outputs(3868) <= layer8_outputs(2220);
    outputs(3869) <= (layer8_outputs(1167)) xor (layer8_outputs(1581));
    outputs(3870) <= (layer8_outputs(1188)) and not (layer8_outputs(393));
    outputs(3871) <= not((layer8_outputs(1596)) xor (layer8_outputs(4888)));
    outputs(3872) <= (layer8_outputs(4712)) xor (layer8_outputs(3923));
    outputs(3873) <= not((layer8_outputs(2030)) xor (layer8_outputs(2933)));
    outputs(3874) <= layer8_outputs(4934);
    outputs(3875) <= not(layer8_outputs(4358));
    outputs(3876) <= not(layer8_outputs(143)) or (layer8_outputs(4867));
    outputs(3877) <= not((layer8_outputs(1243)) or (layer8_outputs(124)));
    outputs(3878) <= (layer8_outputs(838)) and not (layer8_outputs(4));
    outputs(3879) <= (layer8_outputs(816)) xor (layer8_outputs(1833));
    outputs(3880) <= not(layer8_outputs(1363));
    outputs(3881) <= layer8_outputs(3788);
    outputs(3882) <= (layer8_outputs(1644)) xor (layer8_outputs(4192));
    outputs(3883) <= not((layer8_outputs(2796)) xor (layer8_outputs(960)));
    outputs(3884) <= (layer8_outputs(3629)) and not (layer8_outputs(2185));
    outputs(3885) <= not(layer8_outputs(1814));
    outputs(3886) <= not((layer8_outputs(2338)) or (layer8_outputs(77)));
    outputs(3887) <= not((layer8_outputs(1644)) xor (layer8_outputs(4906)));
    outputs(3888) <= not(layer8_outputs(1339));
    outputs(3889) <= layer8_outputs(2555);
    outputs(3890) <= not((layer8_outputs(1829)) or (layer8_outputs(1263)));
    outputs(3891) <= layer8_outputs(1535);
    outputs(3892) <= layer8_outputs(3963);
    outputs(3893) <= not((layer8_outputs(3515)) xor (layer8_outputs(2591)));
    outputs(3894) <= not(layer8_outputs(2011));
    outputs(3895) <= (layer8_outputs(2902)) and not (layer8_outputs(2000));
    outputs(3896) <= not((layer8_outputs(4223)) and (layer8_outputs(1425)));
    outputs(3897) <= (layer8_outputs(496)) and (layer8_outputs(4181));
    outputs(3898) <= not((layer8_outputs(3055)) xor (layer8_outputs(3818)));
    outputs(3899) <= not(layer8_outputs(4462));
    outputs(3900) <= not(layer8_outputs(269));
    outputs(3901) <= not((layer8_outputs(4958)) xor (layer8_outputs(3472)));
    outputs(3902) <= layer8_outputs(1494);
    outputs(3903) <= layer8_outputs(3913);
    outputs(3904) <= not((layer8_outputs(991)) xor (layer8_outputs(2939)));
    outputs(3905) <= not(layer8_outputs(2452));
    outputs(3906) <= not(layer8_outputs(1876));
    outputs(3907) <= (layer8_outputs(2184)) xor (layer8_outputs(1476));
    outputs(3908) <= not((layer8_outputs(4550)) or (layer8_outputs(1023)));
    outputs(3909) <= not(layer8_outputs(1503)) or (layer8_outputs(4988));
    outputs(3910) <= not(layer8_outputs(2952));
    outputs(3911) <= not(layer8_outputs(2762));
    outputs(3912) <= layer8_outputs(343);
    outputs(3913) <= (layer8_outputs(5106)) xor (layer8_outputs(748));
    outputs(3914) <= not(layer8_outputs(3394));
    outputs(3915) <= not(layer8_outputs(3186));
    outputs(3916) <= not(layer8_outputs(3837)) or (layer8_outputs(106));
    outputs(3917) <= (layer8_outputs(397)) xor (layer8_outputs(370));
    outputs(3918) <= layer8_outputs(4950);
    outputs(3919) <= layer8_outputs(1545);
    outputs(3920) <= layer8_outputs(4930);
    outputs(3921) <= not(layer8_outputs(2495)) or (layer8_outputs(585));
    outputs(3922) <= (layer8_outputs(631)) xor (layer8_outputs(3982));
    outputs(3923) <= layer8_outputs(4338);
    outputs(3924) <= (layer8_outputs(4077)) xor (layer8_outputs(3311));
    outputs(3925) <= not(layer8_outputs(2913));
    outputs(3926) <= not((layer8_outputs(1582)) xor (layer8_outputs(5059)));
    outputs(3927) <= not((layer8_outputs(2198)) xor (layer8_outputs(2509)));
    outputs(3928) <= layer8_outputs(644);
    outputs(3929) <= not(layer8_outputs(124));
    outputs(3930) <= (layer8_outputs(2794)) and not (layer8_outputs(1425));
    outputs(3931) <= not(layer8_outputs(3239));
    outputs(3932) <= layer8_outputs(227);
    outputs(3933) <= layer8_outputs(3900);
    outputs(3934) <= not((layer8_outputs(3778)) or (layer8_outputs(3902)));
    outputs(3935) <= not(layer8_outputs(273));
    outputs(3936) <= not((layer8_outputs(3570)) xor (layer8_outputs(171)));
    outputs(3937) <= (layer8_outputs(502)) xor (layer8_outputs(1871));
    outputs(3938) <= layer8_outputs(307);
    outputs(3939) <= not((layer8_outputs(1486)) xor (layer8_outputs(459)));
    outputs(3940) <= (layer8_outputs(782)) xor (layer8_outputs(3330));
    outputs(3941) <= (layer8_outputs(965)) xor (layer8_outputs(3080));
    outputs(3942) <= not((layer8_outputs(3585)) xor (layer8_outputs(3186)));
    outputs(3943) <= layer8_outputs(3900);
    outputs(3944) <= layer8_outputs(918);
    outputs(3945) <= not(layer8_outputs(4579));
    outputs(3946) <= not((layer8_outputs(2947)) xor (layer8_outputs(2107)));
    outputs(3947) <= layer8_outputs(3913);
    outputs(3948) <= layer8_outputs(467);
    outputs(3949) <= layer8_outputs(1601);
    outputs(3950) <= not(layer8_outputs(3008));
    outputs(3951) <= not(layer8_outputs(2281));
    outputs(3952) <= layer8_outputs(1677);
    outputs(3953) <= not(layer8_outputs(4310));
    outputs(3954) <= not(layer8_outputs(4514));
    outputs(3955) <= layer8_outputs(569);
    outputs(3956) <= not((layer8_outputs(2258)) xor (layer8_outputs(1067)));
    outputs(3957) <= not(layer8_outputs(127));
    outputs(3958) <= layer8_outputs(3221);
    outputs(3959) <= (layer8_outputs(2239)) and (layer8_outputs(4754));
    outputs(3960) <= (layer8_outputs(705)) xor (layer8_outputs(919));
    outputs(3961) <= not((layer8_outputs(4561)) xor (layer8_outputs(3871)));
    outputs(3962) <= not(layer8_outputs(2968));
    outputs(3963) <= (layer8_outputs(690)) xor (layer8_outputs(281));
    outputs(3964) <= not((layer8_outputs(3698)) xor (layer8_outputs(2526)));
    outputs(3965) <= (layer8_outputs(1948)) xor (layer8_outputs(3195));
    outputs(3966) <= not((layer8_outputs(3966)) xor (layer8_outputs(703)));
    outputs(3967) <= not((layer8_outputs(4025)) xor (layer8_outputs(1244)));
    outputs(3968) <= not(layer8_outputs(2124));
    outputs(3969) <= (layer8_outputs(1796)) and not (layer8_outputs(5008));
    outputs(3970) <= layer8_outputs(4671);
    outputs(3971) <= layer8_outputs(3604);
    outputs(3972) <= not(layer8_outputs(3091));
    outputs(3973) <= layer8_outputs(1882);
    outputs(3974) <= not(layer8_outputs(2930));
    outputs(3975) <= not((layer8_outputs(4151)) xor (layer8_outputs(4188)));
    outputs(3976) <= layer8_outputs(801);
    outputs(3977) <= (layer8_outputs(2819)) xor (layer8_outputs(3354));
    outputs(3978) <= not((layer8_outputs(3303)) xor (layer8_outputs(3038)));
    outputs(3979) <= (layer8_outputs(4411)) xor (layer8_outputs(2324));
    outputs(3980) <= layer8_outputs(998);
    outputs(3981) <= layer8_outputs(3764);
    outputs(3982) <= not((layer8_outputs(5044)) xor (layer8_outputs(1628)));
    outputs(3983) <= not((layer8_outputs(3380)) xor (layer8_outputs(2471)));
    outputs(3984) <= layer8_outputs(4674);
    outputs(3985) <= (layer8_outputs(692)) xor (layer8_outputs(1631));
    outputs(3986) <= (layer8_outputs(1114)) xor (layer8_outputs(5054));
    outputs(3987) <= (layer8_outputs(762)) and not (layer8_outputs(3639));
    outputs(3988) <= (layer8_outputs(2873)) xor (layer8_outputs(3812));
    outputs(3989) <= layer8_outputs(4083);
    outputs(3990) <= (layer8_outputs(1700)) and not (layer8_outputs(4046));
    outputs(3991) <= not(layer8_outputs(4370));
    outputs(3992) <= not(layer8_outputs(415));
    outputs(3993) <= not(layer8_outputs(2624));
    outputs(3994) <= not((layer8_outputs(5078)) xor (layer8_outputs(2022)));
    outputs(3995) <= layer8_outputs(3222);
    outputs(3996) <= layer8_outputs(1778);
    outputs(3997) <= not(layer8_outputs(1564));
    outputs(3998) <= (layer8_outputs(3384)) xor (layer8_outputs(1192));
    outputs(3999) <= not(layer8_outputs(936));
    outputs(4000) <= layer8_outputs(443);
    outputs(4001) <= layer8_outputs(2709);
    outputs(4002) <= not(layer8_outputs(952));
    outputs(4003) <= not(layer8_outputs(1553));
    outputs(4004) <= not((layer8_outputs(4401)) xor (layer8_outputs(3893)));
    outputs(4005) <= layer8_outputs(2180);
    outputs(4006) <= not((layer8_outputs(763)) xor (layer8_outputs(3205)));
    outputs(4007) <= not((layer8_outputs(2682)) xor (layer8_outputs(4851)));
    outputs(4008) <= not((layer8_outputs(4641)) xor (layer8_outputs(2727)));
    outputs(4009) <= not(layer8_outputs(3757));
    outputs(4010) <= layer8_outputs(3430);
    outputs(4011) <= layer8_outputs(2790);
    outputs(4012) <= (layer8_outputs(3679)) and not (layer8_outputs(4474));
    outputs(4013) <= not(layer8_outputs(2447));
    outputs(4014) <= layer8_outputs(1669);
    outputs(4015) <= (layer8_outputs(4784)) and not (layer8_outputs(2952));
    outputs(4016) <= layer8_outputs(3408);
    outputs(4017) <= (layer8_outputs(1523)) or (layer8_outputs(1253));
    outputs(4018) <= not((layer8_outputs(2733)) and (layer8_outputs(223)));
    outputs(4019) <= not(layer8_outputs(3815));
    outputs(4020) <= not(layer8_outputs(2811));
    outputs(4021) <= layer8_outputs(3315);
    outputs(4022) <= (layer8_outputs(3084)) xor (layer8_outputs(3822));
    outputs(4023) <= not(layer8_outputs(4165));
    outputs(4024) <= not(layer8_outputs(3608));
    outputs(4025) <= layer8_outputs(2086);
    outputs(4026) <= not(layer8_outputs(2303));
    outputs(4027) <= layer8_outputs(18);
    outputs(4028) <= layer8_outputs(2444);
    outputs(4029) <= layer8_outputs(3145);
    outputs(4030) <= (layer8_outputs(3291)) and (layer8_outputs(3935));
    outputs(4031) <= (layer8_outputs(2839)) xor (layer8_outputs(4894));
    outputs(4032) <= not((layer8_outputs(1055)) xor (layer8_outputs(2024)));
    outputs(4033) <= not(layer8_outputs(4152));
    outputs(4034) <= not(layer8_outputs(153));
    outputs(4035) <= not((layer8_outputs(4035)) xor (layer8_outputs(3599)));
    outputs(4036) <= not(layer8_outputs(3819));
    outputs(4037) <= (layer8_outputs(2692)) xor (layer8_outputs(1153));
    outputs(4038) <= not((layer8_outputs(1490)) xor (layer8_outputs(1478)));
    outputs(4039) <= not(layer8_outputs(4392));
    outputs(4040) <= not((layer8_outputs(3754)) xor (layer8_outputs(3641)));
    outputs(4041) <= layer8_outputs(1177);
    outputs(4042) <= (layer8_outputs(1712)) xor (layer8_outputs(3951));
    outputs(4043) <= layer8_outputs(4929);
    outputs(4044) <= (layer8_outputs(2747)) xor (layer8_outputs(4276));
    outputs(4045) <= not(layer8_outputs(4638));
    outputs(4046) <= not((layer8_outputs(3025)) xor (layer8_outputs(3461)));
    outputs(4047) <= layer8_outputs(1817);
    outputs(4048) <= not(layer8_outputs(2761));
    outputs(4049) <= not(layer8_outputs(352)) or (layer8_outputs(2612));
    outputs(4050) <= (layer8_outputs(4296)) and not (layer8_outputs(750));
    outputs(4051) <= (layer8_outputs(34)) and not (layer8_outputs(1574));
    outputs(4052) <= layer8_outputs(4904);
    outputs(4053) <= not((layer8_outputs(2972)) or (layer8_outputs(5066)));
    outputs(4054) <= layer8_outputs(63);
    outputs(4055) <= not(layer8_outputs(2945)) or (layer8_outputs(910));
    outputs(4056) <= not((layer8_outputs(405)) xor (layer8_outputs(2084)));
    outputs(4057) <= layer8_outputs(1444);
    outputs(4058) <= not(layer8_outputs(1693));
    outputs(4059) <= not(layer8_outputs(4020));
    outputs(4060) <= layer8_outputs(1402);
    outputs(4061) <= layer8_outputs(2659);
    outputs(4062) <= not(layer8_outputs(1371));
    outputs(4063) <= not(layer8_outputs(2823));
    outputs(4064) <= (layer8_outputs(4481)) xor (layer8_outputs(1897));
    outputs(4065) <= layer8_outputs(4988);
    outputs(4066) <= not(layer8_outputs(4216));
    outputs(4067) <= layer8_outputs(1591);
    outputs(4068) <= not(layer8_outputs(3341));
    outputs(4069) <= layer8_outputs(93);
    outputs(4070) <= not((layer8_outputs(1149)) xor (layer8_outputs(4966)));
    outputs(4071) <= not(layer8_outputs(4164));
    outputs(4072) <= (layer8_outputs(47)) xor (layer8_outputs(1517));
    outputs(4073) <= not((layer8_outputs(1431)) or (layer8_outputs(4803)));
    outputs(4074) <= not(layer8_outputs(1026));
    outputs(4075) <= layer8_outputs(3455);
    outputs(4076) <= not(layer8_outputs(1027));
    outputs(4077) <= (layer8_outputs(2041)) xor (layer8_outputs(4281));
    outputs(4078) <= layer8_outputs(2246);
    outputs(4079) <= layer8_outputs(2691);
    outputs(4080) <= (layer8_outputs(3021)) xor (layer8_outputs(1907));
    outputs(4081) <= not((layer8_outputs(1326)) xor (layer8_outputs(248)));
    outputs(4082) <= not((layer8_outputs(5046)) xor (layer8_outputs(469)));
    outputs(4083) <= layer8_outputs(325);
    outputs(4084) <= (layer8_outputs(123)) and (layer8_outputs(3138));
    outputs(4085) <= not(layer8_outputs(4792));
    outputs(4086) <= not(layer8_outputs(309));
    outputs(4087) <= not((layer8_outputs(3393)) xor (layer8_outputs(4997)));
    outputs(4088) <= layer8_outputs(1043);
    outputs(4089) <= (layer8_outputs(4206)) xor (layer8_outputs(3048));
    outputs(4090) <= not(layer8_outputs(822));
    outputs(4091) <= layer8_outputs(1652);
    outputs(4092) <= layer8_outputs(1931);
    outputs(4093) <= not((layer8_outputs(690)) xor (layer8_outputs(1041)));
    outputs(4094) <= layer8_outputs(219);
    outputs(4095) <= (layer8_outputs(752)) and not (layer8_outputs(4594));
    outputs(4096) <= (layer8_outputs(15)) and (layer8_outputs(1781));
    outputs(4097) <= (layer8_outputs(1926)) xor (layer8_outputs(1643));
    outputs(4098) <= layer8_outputs(3622);
    outputs(4099) <= not((layer8_outputs(2048)) xor (layer8_outputs(1000)));
    outputs(4100) <= not(layer8_outputs(4068));
    outputs(4101) <= not(layer8_outputs(909));
    outputs(4102) <= not((layer8_outputs(4843)) xor (layer8_outputs(4810)));
    outputs(4103) <= not((layer8_outputs(4540)) xor (layer8_outputs(2348)));
    outputs(4104) <= (layer8_outputs(1877)) xor (layer8_outputs(2817));
    outputs(4105) <= (layer8_outputs(4306)) and (layer8_outputs(4786));
    outputs(4106) <= (layer8_outputs(2496)) xor (layer8_outputs(1445));
    outputs(4107) <= layer8_outputs(2737);
    outputs(4108) <= not(layer8_outputs(4924));
    outputs(4109) <= (layer8_outputs(3404)) xor (layer8_outputs(153));
    outputs(4110) <= layer8_outputs(1472);
    outputs(4111) <= layer8_outputs(2259);
    outputs(4112) <= not((layer8_outputs(4096)) or (layer8_outputs(4270)));
    outputs(4113) <= layer8_outputs(816);
    outputs(4114) <= not(layer8_outputs(4527));
    outputs(4115) <= layer8_outputs(3624);
    outputs(4116) <= not(layer8_outputs(1541));
    outputs(4117) <= not(layer8_outputs(2371));
    outputs(4118) <= not(layer8_outputs(969));
    outputs(4119) <= not(layer8_outputs(1051));
    outputs(4120) <= (layer8_outputs(1085)) xor (layer8_outputs(4569));
    outputs(4121) <= layer8_outputs(891);
    outputs(4122) <= not((layer8_outputs(2987)) xor (layer8_outputs(293)));
    outputs(4123) <= (layer8_outputs(1566)) or (layer8_outputs(179));
    outputs(4124) <= (layer8_outputs(2610)) or (layer8_outputs(2614));
    outputs(4125) <= (layer8_outputs(727)) xor (layer8_outputs(4004));
    outputs(4126) <= layer8_outputs(431);
    outputs(4127) <= layer8_outputs(1361);
    outputs(4128) <= not(layer8_outputs(4902));
    outputs(4129) <= (layer8_outputs(3981)) xor (layer8_outputs(2679));
    outputs(4130) <= (layer8_outputs(3922)) and (layer8_outputs(4085));
    outputs(4131) <= (layer8_outputs(1594)) xor (layer8_outputs(4130));
    outputs(4132) <= layer8_outputs(5075);
    outputs(4133) <= not((layer8_outputs(734)) or (layer8_outputs(925)));
    outputs(4134) <= not((layer8_outputs(2283)) xor (layer8_outputs(3658)));
    outputs(4135) <= not(layer8_outputs(4606));
    outputs(4136) <= not((layer8_outputs(5119)) xor (layer8_outputs(2976)));
    outputs(4137) <= layer8_outputs(339);
    outputs(4138) <= layer8_outputs(4331);
    outputs(4139) <= not((layer8_outputs(962)) xor (layer8_outputs(1459)));
    outputs(4140) <= layer8_outputs(703);
    outputs(4141) <= not(layer8_outputs(5004)) or (layer8_outputs(2323));
    outputs(4142) <= (layer8_outputs(4213)) xor (layer8_outputs(4199));
    outputs(4143) <= not((layer8_outputs(4695)) and (layer8_outputs(2643)));
    outputs(4144) <= not(layer8_outputs(4720));
    outputs(4145) <= (layer8_outputs(2958)) or (layer8_outputs(3721));
    outputs(4146) <= (layer8_outputs(2667)) and not (layer8_outputs(2036));
    outputs(4147) <= (layer8_outputs(4155)) xor (layer8_outputs(31));
    outputs(4148) <= (layer8_outputs(2918)) and not (layer8_outputs(4303));
    outputs(4149) <= not((layer8_outputs(731)) xor (layer8_outputs(605)));
    outputs(4150) <= not(layer8_outputs(3507));
    outputs(4151) <= (layer8_outputs(1939)) xor (layer8_outputs(1276));
    outputs(4152) <= not(layer8_outputs(772));
    outputs(4153) <= not(layer8_outputs(745));
    outputs(4154) <= layer8_outputs(2296);
    outputs(4155) <= not((layer8_outputs(3052)) xor (layer8_outputs(4453)));
    outputs(4156) <= layer8_outputs(4943);
    outputs(4157) <= not(layer8_outputs(931));
    outputs(4158) <= (layer8_outputs(1751)) xor (layer8_outputs(5061));
    outputs(4159) <= (layer8_outputs(1658)) xor (layer8_outputs(1773));
    outputs(4160) <= not(layer8_outputs(4716)) or (layer8_outputs(52));
    outputs(4161) <= not(layer8_outputs(2285));
    outputs(4162) <= layer8_outputs(3847);
    outputs(4163) <= not(layer8_outputs(2909));
    outputs(4164) <= not(layer8_outputs(4981));
    outputs(4165) <= layer8_outputs(912);
    outputs(4166) <= (layer8_outputs(1370)) xor (layer8_outputs(1015));
    outputs(4167) <= not((layer8_outputs(572)) xor (layer8_outputs(4605)));
    outputs(4168) <= layer8_outputs(2622);
    outputs(4169) <= not(layer8_outputs(4022));
    outputs(4170) <= not((layer8_outputs(2065)) xor (layer8_outputs(469)));
    outputs(4171) <= (layer8_outputs(1969)) xor (layer8_outputs(287));
    outputs(4172) <= not(layer8_outputs(3191));
    outputs(4173) <= layer8_outputs(3347);
    outputs(4174) <= not(layer8_outputs(4905));
    outputs(4175) <= (layer8_outputs(1764)) or (layer8_outputs(4354));
    outputs(4176) <= not((layer8_outputs(4038)) xor (layer8_outputs(1811)));
    outputs(4177) <= (layer8_outputs(3630)) xor (layer8_outputs(1667));
    outputs(4178) <= (layer8_outputs(905)) xor (layer8_outputs(3531));
    outputs(4179) <= layer8_outputs(4238);
    outputs(4180) <= layer8_outputs(188);
    outputs(4181) <= not(layer8_outputs(2293)) or (layer8_outputs(1137));
    outputs(4182) <= layer8_outputs(1423);
    outputs(4183) <= layer8_outputs(1098);
    outputs(4184) <= (layer8_outputs(1824)) xor (layer8_outputs(165));
    outputs(4185) <= layer8_outputs(1385);
    outputs(4186) <= not(layer8_outputs(2842));
    outputs(4187) <= (layer8_outputs(2801)) xor (layer8_outputs(3133));
    outputs(4188) <= not(layer8_outputs(792));
    outputs(4189) <= layer8_outputs(5030);
    outputs(4190) <= layer8_outputs(2994);
    outputs(4191) <= layer8_outputs(1615);
    outputs(4192) <= not(layer8_outputs(2536)) or (layer8_outputs(3394));
    outputs(4193) <= not(layer8_outputs(4666)) or (layer8_outputs(92));
    outputs(4194) <= not((layer8_outputs(4360)) xor (layer8_outputs(3868)));
    outputs(4195) <= not(layer8_outputs(4095));
    outputs(4196) <= (layer8_outputs(1245)) xor (layer8_outputs(3685));
    outputs(4197) <= not((layer8_outputs(3044)) xor (layer8_outputs(4458)));
    outputs(4198) <= layer8_outputs(4966);
    outputs(4199) <= layer8_outputs(1586);
    outputs(4200) <= not(layer8_outputs(3342));
    outputs(4201) <= layer8_outputs(2103);
    outputs(4202) <= layer8_outputs(3616);
    outputs(4203) <= not(layer8_outputs(776));
    outputs(4204) <= layer8_outputs(1749);
    outputs(4205) <= layer8_outputs(2131);
    outputs(4206) <= not((layer8_outputs(1453)) xor (layer8_outputs(4178)));
    outputs(4207) <= (layer8_outputs(3288)) xor (layer8_outputs(2752));
    outputs(4208) <= layer8_outputs(3942);
    outputs(4209) <= layer8_outputs(2109);
    outputs(4210) <= not(layer8_outputs(1595));
    outputs(4211) <= (layer8_outputs(1891)) xor (layer8_outputs(3317));
    outputs(4212) <= layer8_outputs(1241);
    outputs(4213) <= (layer8_outputs(425)) xor (layer8_outputs(1353));
    outputs(4214) <= (layer8_outputs(2840)) xor (layer8_outputs(447));
    outputs(4215) <= not(layer8_outputs(1550));
    outputs(4216) <= not(layer8_outputs(4550));
    outputs(4217) <= (layer8_outputs(1666)) and not (layer8_outputs(4811));
    outputs(4218) <= layer8_outputs(1135);
    outputs(4219) <= not((layer8_outputs(2998)) xor (layer8_outputs(4069)));
    outputs(4220) <= not(layer8_outputs(4201));
    outputs(4221) <= not(layer8_outputs(2312));
    outputs(4222) <= not((layer8_outputs(2759)) and (layer8_outputs(4414)));
    outputs(4223) <= not(layer8_outputs(2615));
    outputs(4224) <= layer8_outputs(62);
    outputs(4225) <= not(layer8_outputs(681));
    outputs(4226) <= (layer8_outputs(4160)) xor (layer8_outputs(627));
    outputs(4227) <= not(layer8_outputs(4473));
    outputs(4228) <= not(layer8_outputs(422));
    outputs(4229) <= layer8_outputs(3970);
    outputs(4230) <= not(layer8_outputs(408));
    outputs(4231) <= layer8_outputs(1863);
    outputs(4232) <= layer8_outputs(386);
    outputs(4233) <= (layer8_outputs(4668)) xor (layer8_outputs(3001));
    outputs(4234) <= layer8_outputs(3883);
    outputs(4235) <= layer8_outputs(4099);
    outputs(4236) <= (layer8_outputs(4875)) xor (layer8_outputs(350));
    outputs(4237) <= not(layer8_outputs(3489));
    outputs(4238) <= (layer8_outputs(3720)) and not (layer8_outputs(692));
    outputs(4239) <= not(layer8_outputs(773));
    outputs(4240) <= layer8_outputs(2603);
    outputs(4241) <= layer8_outputs(4394);
    outputs(4242) <= (layer8_outputs(1862)) and (layer8_outputs(3266));
    outputs(4243) <= not(layer8_outputs(583));
    outputs(4244) <= not(layer8_outputs(4456));
    outputs(4245) <= (layer8_outputs(161)) xor (layer8_outputs(3134));
    outputs(4246) <= layer8_outputs(188);
    outputs(4247) <= not(layer8_outputs(3169)) or (layer8_outputs(2068));
    outputs(4248) <= (layer8_outputs(4488)) or (layer8_outputs(1752));
    outputs(4249) <= not(layer8_outputs(125));
    outputs(4250) <= not(layer8_outputs(4203));
    outputs(4251) <= not(layer8_outputs(221));
    outputs(4252) <= not(layer8_outputs(4437));
    outputs(4253) <= layer8_outputs(353);
    outputs(4254) <= not((layer8_outputs(2623)) xor (layer8_outputs(2737)));
    outputs(4255) <= layer8_outputs(3607);
    outputs(4256) <= layer8_outputs(1730);
    outputs(4257) <= not((layer8_outputs(3289)) or (layer8_outputs(3077)));
    outputs(4258) <= not(layer8_outputs(4205));
    outputs(4259) <= not((layer8_outputs(1476)) xor (layer8_outputs(3945)));
    outputs(4260) <= not((layer8_outputs(2300)) xor (layer8_outputs(2536)));
    outputs(4261) <= (layer8_outputs(3619)) xor (layer8_outputs(471));
    outputs(4262) <= not((layer8_outputs(666)) xor (layer8_outputs(4915)));
    outputs(4263) <= layer8_outputs(1329);
    outputs(4264) <= (layer8_outputs(6)) and not (layer8_outputs(2768));
    outputs(4265) <= (layer8_outputs(4058)) xor (layer8_outputs(4971));
    outputs(4266) <= layer8_outputs(4274);
    outputs(4267) <= not((layer8_outputs(955)) xor (layer8_outputs(1847)));
    outputs(4268) <= (layer8_outputs(953)) xor (layer8_outputs(3550));
    outputs(4269) <= layer8_outputs(2262);
    outputs(4270) <= layer8_outputs(2126);
    outputs(4271) <= not((layer8_outputs(2563)) xor (layer8_outputs(2038)));
    outputs(4272) <= not(layer8_outputs(4945));
    outputs(4273) <= (layer8_outputs(4381)) xor (layer8_outputs(372));
    outputs(4274) <= layer8_outputs(3706);
    outputs(4275) <= not(layer8_outputs(3358)) or (layer8_outputs(323));
    outputs(4276) <= not((layer8_outputs(1035)) xor (layer8_outputs(798)));
    outputs(4277) <= (layer8_outputs(460)) xor (layer8_outputs(3541));
    outputs(4278) <= not((layer8_outputs(1969)) xor (layer8_outputs(3376)));
    outputs(4279) <= not(layer8_outputs(413));
    outputs(4280) <= layer8_outputs(1655);
    outputs(4281) <= not(layer8_outputs(110));
    outputs(4282) <= (layer8_outputs(1420)) xor (layer8_outputs(3906));
    outputs(4283) <= (layer8_outputs(3028)) xor (layer8_outputs(1549));
    outputs(4284) <= (layer8_outputs(1132)) xor (layer8_outputs(1376));
    outputs(4285) <= layer8_outputs(4597);
    outputs(4286) <= not(layer8_outputs(1421));
    outputs(4287) <= not(layer8_outputs(4));
    outputs(4288) <= layer8_outputs(2758);
    outputs(4289) <= not((layer8_outputs(1919)) xor (layer8_outputs(4111)));
    outputs(4290) <= (layer8_outputs(4724)) xor (layer8_outputs(2211));
    outputs(4291) <= layer8_outputs(1583);
    outputs(4292) <= not((layer8_outputs(4457)) and (layer8_outputs(4895)));
    outputs(4293) <= not((layer8_outputs(1813)) or (layer8_outputs(3198)));
    outputs(4294) <= (layer8_outputs(4581)) xor (layer8_outputs(2462));
    outputs(4295) <= layer8_outputs(305);
    outputs(4296) <= not(layer8_outputs(4720));
    outputs(4297) <= not((layer8_outputs(4834)) xor (layer8_outputs(2069)));
    outputs(4298) <= layer8_outputs(945);
    outputs(4299) <= not(layer8_outputs(2233)) or (layer8_outputs(653));
    outputs(4300) <= (layer8_outputs(926)) xor (layer8_outputs(1318));
    outputs(4301) <= layer8_outputs(4059);
    outputs(4302) <= (layer8_outputs(1243)) xor (layer8_outputs(1327));
    outputs(4303) <= layer8_outputs(2758);
    outputs(4304) <= (layer8_outputs(697)) xor (layer8_outputs(4954));
    outputs(4305) <= layer8_outputs(384);
    outputs(4306) <= not(layer8_outputs(392)) or (layer8_outputs(707));
    outputs(4307) <= not(layer8_outputs(1995));
    outputs(4308) <= not(layer8_outputs(3406));
    outputs(4309) <= layer8_outputs(1786);
    outputs(4310) <= not(layer8_outputs(2538)) or (layer8_outputs(2764));
    outputs(4311) <= (layer8_outputs(3003)) xor (layer8_outputs(2258));
    outputs(4312) <= layer8_outputs(4235);
    outputs(4313) <= not((layer8_outputs(2132)) xor (layer8_outputs(2442)));
    outputs(4314) <= not((layer8_outputs(1691)) xor (layer8_outputs(4543)));
    outputs(4315) <= layer8_outputs(3377);
    outputs(4316) <= layer8_outputs(4523);
    outputs(4317) <= not((layer8_outputs(173)) xor (layer8_outputs(464)));
    outputs(4318) <= not((layer8_outputs(1757)) and (layer8_outputs(3552)));
    outputs(4319) <= not(layer8_outputs(1298)) or (layer8_outputs(670));
    outputs(4320) <= layer8_outputs(1195);
    outputs(4321) <= (layer8_outputs(4582)) xor (layer8_outputs(4959));
    outputs(4322) <= layer8_outputs(2424);
    outputs(4323) <= layer8_outputs(2394);
    outputs(4324) <= layer8_outputs(36);
    outputs(4325) <= not(layer8_outputs(1306));
    outputs(4326) <= not(layer8_outputs(2433));
    outputs(4327) <= (layer8_outputs(600)) xor (layer8_outputs(865));
    outputs(4328) <= not(layer8_outputs(2122));
    outputs(4329) <= not(layer8_outputs(890));
    outputs(4330) <= (layer8_outputs(2505)) xor (layer8_outputs(4878));
    outputs(4331) <= (layer8_outputs(5039)) and not (layer8_outputs(968));
    outputs(4332) <= not((layer8_outputs(4658)) xor (layer8_outputs(403)));
    outputs(4333) <= not(layer8_outputs(4669));
    outputs(4334) <= layer8_outputs(2561);
    outputs(4335) <= layer8_outputs(1032);
    outputs(4336) <= not(layer8_outputs(2995));
    outputs(4337) <= layer8_outputs(305);
    outputs(4338) <= (layer8_outputs(3747)) and not (layer8_outputs(4401));
    outputs(4339) <= not((layer8_outputs(1204)) xor (layer8_outputs(262)));
    outputs(4340) <= (layer8_outputs(2634)) xor (layer8_outputs(902));
    outputs(4341) <= (layer8_outputs(2587)) xor (layer8_outputs(1642));
    outputs(4342) <= not(layer8_outputs(4515));
    outputs(4343) <= not(layer8_outputs(4721)) or (layer8_outputs(3832));
    outputs(4344) <= (layer8_outputs(821)) xor (layer8_outputs(4626));
    outputs(4345) <= (layer8_outputs(3228)) and not (layer8_outputs(4045));
    outputs(4346) <= not(layer8_outputs(2986));
    outputs(4347) <= (layer8_outputs(3350)) xor (layer8_outputs(4951));
    outputs(4348) <= (layer8_outputs(90)) xor (layer8_outputs(149));
    outputs(4349) <= not(layer8_outputs(2739)) or (layer8_outputs(2711));
    outputs(4350) <= not(layer8_outputs(1240));
    outputs(4351) <= not(layer8_outputs(3881)) or (layer8_outputs(3515));
    outputs(4352) <= not(layer8_outputs(4391)) or (layer8_outputs(2592));
    outputs(4353) <= not(layer8_outputs(1286)) or (layer8_outputs(1200));
    outputs(4354) <= layer8_outputs(2848);
    outputs(4355) <= layer8_outputs(4144);
    outputs(4356) <= not(layer8_outputs(2870));
    outputs(4357) <= (layer8_outputs(4060)) and not (layer8_outputs(4210));
    outputs(4358) <= not(layer8_outputs(837));
    outputs(4359) <= layer8_outputs(2583);
    outputs(4360) <= layer8_outputs(1626);
    outputs(4361) <= not(layer8_outputs(2116));
    outputs(4362) <= not(layer8_outputs(5021));
    outputs(4363) <= (layer8_outputs(2569)) xor (layer8_outputs(4209));
    outputs(4364) <= not((layer8_outputs(3602)) xor (layer8_outputs(818)));
    outputs(4365) <= not(layer8_outputs(4090));
    outputs(4366) <= layer8_outputs(2183);
    outputs(4367) <= not((layer8_outputs(4389)) xor (layer8_outputs(1742)));
    outputs(4368) <= layer8_outputs(354);
    outputs(4369) <= layer8_outputs(4978);
    outputs(4370) <= layer8_outputs(4006);
    outputs(4371) <= not(layer8_outputs(482));
    outputs(4372) <= (layer8_outputs(1567)) xor (layer8_outputs(4482));
    outputs(4373) <= not((layer8_outputs(4467)) xor (layer8_outputs(2802)));
    outputs(4374) <= not(layer8_outputs(695));
    outputs(4375) <= layer8_outputs(4441);
    outputs(4376) <= not(layer8_outputs(4498));
    outputs(4377) <= layer8_outputs(3387);
    outputs(4378) <= (layer8_outputs(4800)) and not (layer8_outputs(5042));
    outputs(4379) <= not(layer8_outputs(4242));
    outputs(4380) <= (layer8_outputs(150)) xor (layer8_outputs(108));
    outputs(4381) <= layer8_outputs(3116);
    outputs(4382) <= layer8_outputs(50);
    outputs(4383) <= (layer8_outputs(3773)) xor (layer8_outputs(4710));
    outputs(4384) <= not((layer8_outputs(2034)) xor (layer8_outputs(344)));
    outputs(4385) <= not((layer8_outputs(1620)) xor (layer8_outputs(3589)));
    outputs(4386) <= not((layer8_outputs(1368)) xor (layer8_outputs(4123)));
    outputs(4387) <= layer8_outputs(2748);
    outputs(4388) <= not(layer8_outputs(3085));
    outputs(4389) <= layer8_outputs(689);
    outputs(4390) <= layer8_outputs(4619);
    outputs(4391) <= (layer8_outputs(4806)) and not (layer8_outputs(1305));
    outputs(4392) <= not(layer8_outputs(3535)) or (layer8_outputs(4469));
    outputs(4393) <= not(layer8_outputs(1838)) or (layer8_outputs(2888));
    outputs(4394) <= (layer8_outputs(3451)) xor (layer8_outputs(2147));
    outputs(4395) <= (layer8_outputs(1736)) or (layer8_outputs(5109));
    outputs(4396) <= not(layer8_outputs(2472));
    outputs(4397) <= layer8_outputs(5102);
    outputs(4398) <= layer8_outputs(4565);
    outputs(4399) <= (layer8_outputs(233)) xor (layer8_outputs(3577));
    outputs(4400) <= not((layer8_outputs(3855)) or (layer8_outputs(3862)));
    outputs(4401) <= layer8_outputs(3449);
    outputs(4402) <= (layer8_outputs(3813)) and not (layer8_outputs(2649));
    outputs(4403) <= not(layer8_outputs(1783));
    outputs(4404) <= layer8_outputs(4911);
    outputs(4405) <= not(layer8_outputs(3470));
    outputs(4406) <= not(layer8_outputs(553)) or (layer8_outputs(1160));
    outputs(4407) <= (layer8_outputs(1568)) xor (layer8_outputs(827));
    outputs(4408) <= not(layer8_outputs(4811));
    outputs(4409) <= (layer8_outputs(4080)) xor (layer8_outputs(1651));
    outputs(4410) <= not(layer8_outputs(3811));
    outputs(4411) <= not(layer8_outputs(3683));
    outputs(4412) <= layer8_outputs(3413);
    outputs(4413) <= layer8_outputs(3438);
    outputs(4414) <= layer8_outputs(3747);
    outputs(4415) <= (layer8_outputs(3519)) xor (layer8_outputs(4860));
    outputs(4416) <= not((layer8_outputs(4151)) xor (layer8_outputs(2792)));
    outputs(4417) <= layer8_outputs(3947);
    outputs(4418) <= layer8_outputs(2234);
    outputs(4419) <= not(layer8_outputs(3950));
    outputs(4420) <= not(layer8_outputs(4347));
    outputs(4421) <= not(layer8_outputs(41));
    outputs(4422) <= (layer8_outputs(667)) and (layer8_outputs(1123));
    outputs(4423) <= not((layer8_outputs(894)) xor (layer8_outputs(2767)));
    outputs(4424) <= not((layer8_outputs(2519)) xor (layer8_outputs(1557)));
    outputs(4425) <= not(layer8_outputs(3827));
    outputs(4426) <= (layer8_outputs(835)) xor (layer8_outputs(3562));
    outputs(4427) <= not(layer8_outputs(2946));
    outputs(4428) <= not((layer8_outputs(3301)) xor (layer8_outputs(4702)));
    outputs(4429) <= (layer8_outputs(2031)) xor (layer8_outputs(2558));
    outputs(4430) <= not((layer8_outputs(968)) xor (layer8_outputs(1021)));
    outputs(4431) <= (layer8_outputs(3914)) xor (layer8_outputs(3938));
    outputs(4432) <= not(layer8_outputs(1356));
    outputs(4433) <= not(layer8_outputs(522));
    outputs(4434) <= not(layer8_outputs(1281)) or (layer8_outputs(5088));
    outputs(4435) <= not(layer8_outputs(3192));
    outputs(4436) <= not((layer8_outputs(4299)) xor (layer8_outputs(1028)));
    outputs(4437) <= not((layer8_outputs(3152)) xor (layer8_outputs(2999)));
    outputs(4438) <= (layer8_outputs(3545)) xor (layer8_outputs(1151));
    outputs(4439) <= (layer8_outputs(634)) xor (layer8_outputs(4442));
    outputs(4440) <= (layer8_outputs(4182)) xor (layer8_outputs(765));
    outputs(4441) <= (layer8_outputs(4224)) and not (layer8_outputs(178));
    outputs(4442) <= layer8_outputs(3432);
    outputs(4443) <= layer8_outputs(854);
    outputs(4444) <= not((layer8_outputs(303)) xor (layer8_outputs(497)));
    outputs(4445) <= not(layer8_outputs(28));
    outputs(4446) <= layer8_outputs(4889);
    outputs(4447) <= not(layer8_outputs(3935));
    outputs(4448) <= not((layer8_outputs(1922)) or (layer8_outputs(4817)));
    outputs(4449) <= (layer8_outputs(4563)) xor (layer8_outputs(322));
    outputs(4450) <= layer8_outputs(2045);
    outputs(4451) <= not(layer8_outputs(2455));
    outputs(4452) <= layer8_outputs(3706);
    outputs(4453) <= layer8_outputs(853);
    outputs(4454) <= layer8_outputs(970);
    outputs(4455) <= not((layer8_outputs(3776)) xor (layer8_outputs(455)));
    outputs(4456) <= not(layer8_outputs(4153));
    outputs(4457) <= not(layer8_outputs(4156));
    outputs(4458) <= (layer8_outputs(3902)) and not (layer8_outputs(2615));
    outputs(4459) <= layer8_outputs(4200);
    outputs(4460) <= not((layer8_outputs(3506)) xor (layer8_outputs(2438)));
    outputs(4461) <= not((layer8_outputs(1774)) xor (layer8_outputs(2099)));
    outputs(4462) <= not(layer8_outputs(4249));
    outputs(4463) <= layer8_outputs(2211);
    outputs(4464) <= (layer8_outputs(374)) xor (layer8_outputs(1525));
    outputs(4465) <= layer8_outputs(191);
    outputs(4466) <= not(layer8_outputs(1166));
    outputs(4467) <= not((layer8_outputs(3534)) xor (layer8_outputs(3297)));
    outputs(4468) <= layer8_outputs(2849);
    outputs(4469) <= not((layer8_outputs(4025)) xor (layer8_outputs(3313)));
    outputs(4470) <= layer8_outputs(2537);
    outputs(4471) <= (layer8_outputs(1216)) xor (layer8_outputs(4979));
    outputs(4472) <= not(layer8_outputs(5093)) or (layer8_outputs(21));
    outputs(4473) <= not((layer8_outputs(3962)) xor (layer8_outputs(2404)));
    outputs(4474) <= not(layer8_outputs(4236));
    outputs(4475) <= not(layer8_outputs(4061)) or (layer8_outputs(3360));
    outputs(4476) <= (layer8_outputs(2591)) and not (layer8_outputs(2816));
    outputs(4477) <= not(layer8_outputs(3240));
    outputs(4478) <= not((layer8_outputs(3742)) or (layer8_outputs(3338)));
    outputs(4479) <= not(layer8_outputs(1697)) or (layer8_outputs(1438));
    outputs(4480) <= not(layer8_outputs(2331));
    outputs(4481) <= layer8_outputs(4653);
    outputs(4482) <= not((layer8_outputs(1154)) and (layer8_outputs(3739)));
    outputs(4483) <= (layer8_outputs(3841)) or (layer8_outputs(3804));
    outputs(4484) <= not(layer8_outputs(1292));
    outputs(4485) <= not((layer8_outputs(1307)) xor (layer8_outputs(4673)));
    outputs(4486) <= not((layer8_outputs(5014)) xor (layer8_outputs(5057)));
    outputs(4487) <= not(layer8_outputs(1198));
    outputs(4488) <= not(layer8_outputs(1131));
    outputs(4489) <= layer8_outputs(2685);
    outputs(4490) <= not(layer8_outputs(4863));
    outputs(4491) <= not((layer8_outputs(2713)) xor (layer8_outputs(4080)));
    outputs(4492) <= layer8_outputs(2197);
    outputs(4493) <= not((layer8_outputs(407)) and (layer8_outputs(4193)));
    outputs(4494) <= not(layer8_outputs(3284));
    outputs(4495) <= not(layer8_outputs(3150));
    outputs(4496) <= not(layer8_outputs(2803));
    outputs(4497) <= not((layer8_outputs(4848)) or (layer8_outputs(4608)));
    outputs(4498) <= not((layer8_outputs(1532)) xor (layer8_outputs(2605)));
    outputs(4499) <= (layer8_outputs(278)) xor (layer8_outputs(1662));
    outputs(4500) <= layer8_outputs(4466);
    outputs(4501) <= (layer8_outputs(4847)) xor (layer8_outputs(3596));
    outputs(4502) <= layer8_outputs(2413);
    outputs(4503) <= layer8_outputs(1551);
    outputs(4504) <= not((layer8_outputs(4772)) xor (layer8_outputs(4961)));
    outputs(4505) <= not(layer8_outputs(271));
    outputs(4506) <= (layer8_outputs(606)) or (layer8_outputs(4624));
    outputs(4507) <= (layer8_outputs(1489)) and (layer8_outputs(1999));
    outputs(4508) <= not(layer8_outputs(1500));
    outputs(4509) <= not(layer8_outputs(2860)) or (layer8_outputs(3791));
    outputs(4510) <= (layer8_outputs(4096)) xor (layer8_outputs(2257));
    outputs(4511) <= layer8_outputs(3857);
    outputs(4512) <= not((layer8_outputs(1443)) and (layer8_outputs(5016)));
    outputs(4513) <= not((layer8_outputs(1622)) or (layer8_outputs(1646)));
    outputs(4514) <= layer8_outputs(1475);
    outputs(4515) <= not(layer8_outputs(2838));
    outputs(4516) <= not(layer8_outputs(3824));
    outputs(4517) <= (layer8_outputs(550)) xor (layer8_outputs(3795));
    outputs(4518) <= not(layer8_outputs(555)) or (layer8_outputs(636));
    outputs(4519) <= (layer8_outputs(2223)) xor (layer8_outputs(3736));
    outputs(4520) <= not(layer8_outputs(45));
    outputs(4521) <= layer8_outputs(2524);
    outputs(4522) <= not((layer8_outputs(3556)) xor (layer8_outputs(4030)));
    outputs(4523) <= not((layer8_outputs(2940)) xor (layer8_outputs(886)));
    outputs(4524) <= not((layer8_outputs(4734)) and (layer8_outputs(373)));
    outputs(4525) <= layer8_outputs(664);
    outputs(4526) <= (layer8_outputs(3772)) xor (layer8_outputs(4908));
    outputs(4527) <= layer8_outputs(1473);
    outputs(4528) <= not(layer8_outputs(336));
    outputs(4529) <= not((layer8_outputs(1732)) xor (layer8_outputs(70)));
    outputs(4530) <= not(layer8_outputs(5077)) or (layer8_outputs(3158));
    outputs(4531) <= layer8_outputs(1967);
    outputs(4532) <= not(layer8_outputs(3010));
    outputs(4533) <= (layer8_outputs(2061)) and not (layer8_outputs(2364));
    outputs(4534) <= not((layer8_outputs(2268)) or (layer8_outputs(258)));
    outputs(4535) <= not(layer8_outputs(4388));
    outputs(4536) <= (layer8_outputs(4650)) or (layer8_outputs(1942));
    outputs(4537) <= not((layer8_outputs(3088)) xor (layer8_outputs(3319)));
    outputs(4538) <= (layer8_outputs(4171)) or (layer8_outputs(4735));
    outputs(4539) <= layer8_outputs(885);
    outputs(4540) <= not(layer8_outputs(4845));
    outputs(4541) <= not(layer8_outputs(978));
    outputs(4542) <= (layer8_outputs(5062)) xor (layer8_outputs(2227));
    outputs(4543) <= not((layer8_outputs(4945)) or (layer8_outputs(94)));
    outputs(4544) <= not((layer8_outputs(1058)) xor (layer8_outputs(4674)));
    outputs(4545) <= not(layer8_outputs(3043));
    outputs(4546) <= (layer8_outputs(5002)) xor (layer8_outputs(3125));
    outputs(4547) <= (layer8_outputs(3369)) xor (layer8_outputs(1215));
    outputs(4548) <= (layer8_outputs(2778)) xor (layer8_outputs(349));
    outputs(4549) <= (layer8_outputs(3978)) or (layer8_outputs(4466));
    outputs(4550) <= layer8_outputs(1608);
    outputs(4551) <= layer8_outputs(3345);
    outputs(4552) <= (layer8_outputs(1584)) xor (layer8_outputs(442));
    outputs(4553) <= layer8_outputs(1717);
    outputs(4554) <= layer8_outputs(3499);
    outputs(4555) <= not((layer8_outputs(1878)) xor (layer8_outputs(2009)));
    outputs(4556) <= (layer8_outputs(1618)) xor (layer8_outputs(2936));
    outputs(4557) <= layer8_outputs(2498);
    outputs(4558) <= layer8_outputs(1798);
    outputs(4559) <= layer8_outputs(4392);
    outputs(4560) <= (layer8_outputs(4564)) xor (layer8_outputs(3077));
    outputs(4561) <= layer8_outputs(2687);
    outputs(4562) <= layer8_outputs(3594);
    outputs(4563) <= not((layer8_outputs(2309)) xor (layer8_outputs(4563)));
    outputs(4564) <= not(layer8_outputs(3812));
    outputs(4565) <= layer8_outputs(1);
    outputs(4566) <= not(layer8_outputs(2910));
    outputs(4567) <= layer8_outputs(2038);
    outputs(4568) <= not((layer8_outputs(264)) xor (layer8_outputs(4616)));
    outputs(4569) <= not(layer8_outputs(3998));
    outputs(4570) <= (layer8_outputs(895)) xor (layer8_outputs(151));
    outputs(4571) <= not(layer8_outputs(4957));
    outputs(4572) <= not((layer8_outputs(2714)) xor (layer8_outputs(618)));
    outputs(4573) <= not((layer8_outputs(354)) xor (layer8_outputs(3232)));
    outputs(4574) <= not(layer8_outputs(3865));
    outputs(4575) <= not(layer8_outputs(4289));
    outputs(4576) <= layer8_outputs(2326);
    outputs(4577) <= not(layer8_outputs(4854));
    outputs(4578) <= not(layer8_outputs(3172));
    outputs(4579) <= not(layer8_outputs(2962));
    outputs(4580) <= layer8_outputs(1029);
    outputs(4581) <= not((layer8_outputs(2957)) and (layer8_outputs(5091)));
    outputs(4582) <= not(layer8_outputs(4220));
    outputs(4583) <= layer8_outputs(1147);
    outputs(4584) <= not((layer8_outputs(1250)) xor (layer8_outputs(145)));
    outputs(4585) <= not((layer8_outputs(2672)) xor (layer8_outputs(1376)));
    outputs(4586) <= not(layer8_outputs(2135));
    outputs(4587) <= not(layer8_outputs(1202));
    outputs(4588) <= layer8_outputs(559);
    outputs(4589) <= not(layer8_outputs(1303));
    outputs(4590) <= layer8_outputs(1342);
    outputs(4591) <= not((layer8_outputs(1902)) xor (layer8_outputs(1280)));
    outputs(4592) <= not((layer8_outputs(3058)) xor (layer8_outputs(2144)));
    outputs(4593) <= not(layer8_outputs(257));
    outputs(4594) <= (layer8_outputs(3618)) xor (layer8_outputs(4143));
    outputs(4595) <= not(layer8_outputs(2173));
    outputs(4596) <= (layer8_outputs(3259)) xor (layer8_outputs(1280));
    outputs(4597) <= not((layer8_outputs(4572)) xor (layer8_outputs(4716)));
    outputs(4598) <= not(layer8_outputs(4196)) or (layer8_outputs(1140));
    outputs(4599) <= layer8_outputs(169);
    outputs(4600) <= (layer8_outputs(1570)) and not (layer8_outputs(3170));
    outputs(4601) <= layer8_outputs(1189);
    outputs(4602) <= not(layer8_outputs(2992));
    outputs(4603) <= layer8_outputs(87);
    outputs(4604) <= not(layer8_outputs(1409));
    outputs(4605) <= not(layer8_outputs(3554));
    outputs(4606) <= (layer8_outputs(2227)) xor (layer8_outputs(276));
    outputs(4607) <= layer8_outputs(141);
    outputs(4608) <= not((layer8_outputs(113)) xor (layer8_outputs(1929)));
    outputs(4609) <= layer8_outputs(812);
    outputs(4610) <= layer8_outputs(1043);
    outputs(4611) <= (layer8_outputs(2097)) xor (layer8_outputs(4893));
    outputs(4612) <= layer8_outputs(5105);
    outputs(4613) <= not((layer8_outputs(2337)) xor (layer8_outputs(1831)));
    outputs(4614) <= (layer8_outputs(2565)) xor (layer8_outputs(1268));
    outputs(4615) <= (layer8_outputs(3937)) and not (layer8_outputs(245));
    outputs(4616) <= not(layer8_outputs(3863));
    outputs(4617) <= not(layer8_outputs(2486));
    outputs(4618) <= layer8_outputs(1450);
    outputs(4619) <= not(layer8_outputs(5118));
    outputs(4620) <= not(layer8_outputs(4594));
    outputs(4621) <= (layer8_outputs(1777)) xor (layer8_outputs(1088));
    outputs(4622) <= not((layer8_outputs(1616)) or (layer8_outputs(1734)));
    outputs(4623) <= (layer8_outputs(4571)) xor (layer8_outputs(4795));
    outputs(4624) <= layer8_outputs(2503);
    outputs(4625) <= layer8_outputs(436);
    outputs(4626) <= not(layer8_outputs(1536));
    outputs(4627) <= (layer8_outputs(157)) xor (layer8_outputs(504));
    outputs(4628) <= not(layer8_outputs(3561));
    outputs(4629) <= not(layer8_outputs(2265));
    outputs(4630) <= not((layer8_outputs(3512)) xor (layer8_outputs(4676)));
    outputs(4631) <= (layer8_outputs(3586)) and not (layer8_outputs(4417));
    outputs(4632) <= not((layer8_outputs(3163)) xor (layer8_outputs(619)));
    outputs(4633) <= not((layer8_outputs(473)) xor (layer8_outputs(4289)));
    outputs(4634) <= (layer8_outputs(1680)) and not (layer8_outputs(4380));
    outputs(4635) <= not(layer8_outputs(5008));
    outputs(4636) <= (layer8_outputs(1834)) xor (layer8_outputs(1719));
    outputs(4637) <= not(layer8_outputs(4515));
    outputs(4638) <= layer8_outputs(2662);
    outputs(4639) <= not(layer8_outputs(4367));
    outputs(4640) <= (layer8_outputs(4877)) xor (layer8_outputs(932));
    outputs(4641) <= not(layer8_outputs(1745));
    outputs(4642) <= not(layer8_outputs(3447));
    outputs(4643) <= (layer8_outputs(1895)) and (layer8_outputs(3089));
    outputs(4644) <= (layer8_outputs(4996)) xor (layer8_outputs(4890));
    outputs(4645) <= layer8_outputs(721);
    outputs(4646) <= (layer8_outputs(1725)) xor (layer8_outputs(4312));
    outputs(4647) <= layer8_outputs(1152);
    outputs(4648) <= (layer8_outputs(1254)) and not (layer8_outputs(4139));
    outputs(4649) <= not(layer8_outputs(1546));
    outputs(4650) <= layer8_outputs(3861);
    outputs(4651) <= not((layer8_outputs(2087)) xor (layer8_outputs(3765)));
    outputs(4652) <= not(layer8_outputs(3761));
    outputs(4653) <= layer8_outputs(4580);
    outputs(4654) <= layer8_outputs(5074);
    outputs(4655) <= layer8_outputs(1581);
    outputs(4656) <= not(layer8_outputs(518));
    outputs(4657) <= not(layer8_outputs(458));
    outputs(4658) <= not((layer8_outputs(154)) and (layer8_outputs(3627)));
    outputs(4659) <= (layer8_outputs(3274)) and not (layer8_outputs(1396));
    outputs(4660) <= not(layer8_outputs(1407));
    outputs(4661) <= layer8_outputs(356);
    outputs(4662) <= not((layer8_outputs(2412)) or (layer8_outputs(5115)));
    outputs(4663) <= not(layer8_outputs(909));
    outputs(4664) <= not((layer8_outputs(4682)) or (layer8_outputs(1711)));
    outputs(4665) <= not((layer8_outputs(1227)) and (layer8_outputs(4412)));
    outputs(4666) <= (layer8_outputs(4852)) and not (layer8_outputs(4628));
    outputs(4667) <= (layer8_outputs(564)) and (layer8_outputs(3549));
    outputs(4668) <= not(layer8_outputs(3438));
    outputs(4669) <= not(layer8_outputs(4763));
    outputs(4670) <= layer8_outputs(3434);
    outputs(4671) <= layer8_outputs(4404);
    outputs(4672) <= (layer8_outputs(2324)) xor (layer8_outputs(3111));
    outputs(4673) <= not(layer8_outputs(3787));
    outputs(4674) <= not(layer8_outputs(880));
    outputs(4675) <= layer8_outputs(4184);
    outputs(4676) <= (layer8_outputs(4656)) xor (layer8_outputs(3223));
    outputs(4677) <= (layer8_outputs(1565)) xor (layer8_outputs(2121));
    outputs(4678) <= layer8_outputs(1535);
    outputs(4679) <= layer8_outputs(193);
    outputs(4680) <= not(layer8_outputs(2120));
    outputs(4681) <= not((layer8_outputs(3263)) xor (layer8_outputs(987)));
    outputs(4682) <= not(layer8_outputs(3840));
    outputs(4683) <= not(layer8_outputs(4320));
    outputs(4684) <= layer8_outputs(3877);
    outputs(4685) <= (layer8_outputs(3287)) xor (layer8_outputs(2042));
    outputs(4686) <= layer8_outputs(4250);
    outputs(4687) <= layer8_outputs(4793);
    outputs(4688) <= not(layer8_outputs(3909));
    outputs(4689) <= not(layer8_outputs(4981));
    outputs(4690) <= layer8_outputs(2396);
    outputs(4691) <= not((layer8_outputs(2288)) xor (layer8_outputs(4497)));
    outputs(4692) <= layer8_outputs(561);
    outputs(4693) <= not((layer8_outputs(1582)) xor (layer8_outputs(524)));
    outputs(4694) <= not(layer8_outputs(2972));
    outputs(4695) <= layer8_outputs(33);
    outputs(4696) <= not((layer8_outputs(3579)) xor (layer8_outputs(2248)));
    outputs(4697) <= (layer8_outputs(3151)) xor (layer8_outputs(2306));
    outputs(4698) <= layer8_outputs(2154);
    outputs(4699) <= not(layer8_outputs(1617));
    outputs(4700) <= not((layer8_outputs(4823)) xor (layer8_outputs(289)));
    outputs(4701) <= not(layer8_outputs(2620));
    outputs(4702) <= layer8_outputs(446);
    outputs(4703) <= (layer8_outputs(3988)) and (layer8_outputs(3053));
    outputs(4704) <= not(layer8_outputs(3689));
    outputs(4705) <= layer8_outputs(3034);
    outputs(4706) <= layer8_outputs(4495);
    outputs(4707) <= (layer8_outputs(558)) xor (layer8_outputs(3830));
    outputs(4708) <= not(layer8_outputs(1630));
    outputs(4709) <= layer8_outputs(4661);
    outputs(4710) <= layer8_outputs(2252);
    outputs(4711) <= not((layer8_outputs(3078)) xor (layer8_outputs(2647)));
    outputs(4712) <= layer8_outputs(2656);
    outputs(4713) <= not(layer8_outputs(3007));
    outputs(4714) <= not(layer8_outputs(4921));
    outputs(4715) <= layer8_outputs(885);
    outputs(4716) <= layer8_outputs(1209);
    outputs(4717) <= not(layer8_outputs(3729));
    outputs(4718) <= not((layer8_outputs(3416)) xor (layer8_outputs(1477)));
    outputs(4719) <= not((layer8_outputs(4799)) xor (layer8_outputs(1072)));
    outputs(4720) <= not(layer8_outputs(2358));
    outputs(4721) <= not(layer8_outputs(2754));
    outputs(4722) <= layer8_outputs(4756);
    outputs(4723) <= not(layer8_outputs(269));
    outputs(4724) <= (layer8_outputs(4846)) xor (layer8_outputs(2300));
    outputs(4725) <= not((layer8_outputs(1914)) and (layer8_outputs(1421)));
    outputs(4726) <= (layer8_outputs(5065)) and not (layer8_outputs(1984));
    outputs(4727) <= not((layer8_outputs(1881)) and (layer8_outputs(3455)));
    outputs(4728) <= not(layer8_outputs(1410));
    outputs(4729) <= not((layer8_outputs(790)) or (layer8_outputs(2889)));
    outputs(4730) <= layer8_outputs(1432);
    outputs(4731) <= (layer8_outputs(2729)) xor (layer8_outputs(23));
    outputs(4732) <= layer8_outputs(3459);
    outputs(4733) <= not(layer8_outputs(4034));
    outputs(4734) <= not(layer8_outputs(4714));
    outputs(4735) <= not(layer8_outputs(1257));
    outputs(4736) <= not(layer8_outputs(3895));
    outputs(4737) <= not((layer8_outputs(3767)) xor (layer8_outputs(4355)));
    outputs(4738) <= (layer8_outputs(1661)) xor (layer8_outputs(4007));
    outputs(4739) <= layer8_outputs(2229);
    outputs(4740) <= not(layer8_outputs(2170));
    outputs(4741) <= not(layer8_outputs(3297));
    outputs(4742) <= not(layer8_outputs(1379));
    outputs(4743) <= not((layer8_outputs(958)) and (layer8_outputs(1538)));
    outputs(4744) <= not((layer8_outputs(3231)) xor (layer8_outputs(2112)));
    outputs(4745) <= not(layer8_outputs(245));
    outputs(4746) <= layer8_outputs(2341);
    outputs(4747) <= not((layer8_outputs(3678)) xor (layer8_outputs(4678)));
    outputs(4748) <= (layer8_outputs(2815)) xor (layer8_outputs(1621));
    outputs(4749) <= layer8_outputs(2586);
    outputs(4750) <= layer8_outputs(2542);
    outputs(4751) <= layer8_outputs(2026);
    outputs(4752) <= layer8_outputs(826);
    outputs(4753) <= not(layer8_outputs(2830));
    outputs(4754) <= (layer8_outputs(3637)) or (layer8_outputs(937));
    outputs(4755) <= layer8_outputs(721);
    outputs(4756) <= not((layer8_outputs(1296)) xor (layer8_outputs(4329)));
    outputs(4757) <= layer8_outputs(3203);
    outputs(4758) <= (layer8_outputs(1512)) and not (layer8_outputs(5035));
    outputs(4759) <= (layer8_outputs(1815)) and not (layer8_outputs(1896));
    outputs(4760) <= layer8_outputs(1769);
    outputs(4761) <= not(layer8_outputs(1012));
    outputs(4762) <= not(layer8_outputs(3362));
    outputs(4763) <= not((layer8_outputs(723)) xor (layer8_outputs(3972)));
    outputs(4764) <= not((layer8_outputs(4203)) xor (layer8_outputs(4634)));
    outputs(4765) <= not((layer8_outputs(2616)) and (layer8_outputs(2725)));
    outputs(4766) <= (layer8_outputs(1558)) xor (layer8_outputs(2012));
    outputs(4767) <= layer8_outputs(4183);
    outputs(4768) <= not(layer8_outputs(4600));
    outputs(4769) <= (layer8_outputs(412)) xor (layer8_outputs(5057));
    outputs(4770) <= not(layer8_outputs(568));
    outputs(4771) <= (layer8_outputs(2776)) xor (layer8_outputs(3024));
    outputs(4772) <= not(layer8_outputs(4924));
    outputs(4773) <= (layer8_outputs(1308)) and not (layer8_outputs(1061));
    outputs(4774) <= not((layer8_outputs(4768)) xor (layer8_outputs(1350)));
    outputs(4775) <= layer8_outputs(2753);
    outputs(4776) <= not(layer8_outputs(2495));
    outputs(4777) <= (layer8_outputs(1961)) and not (layer8_outputs(633));
    outputs(4778) <= layer8_outputs(4463);
    outputs(4779) <= not(layer8_outputs(1949));
    outputs(4780) <= not((layer8_outputs(4547)) xor (layer8_outputs(1941)));
    outputs(4781) <= layer8_outputs(1224);
    outputs(4782) <= layer8_outputs(4791);
    outputs(4783) <= not(layer8_outputs(1105));
    outputs(4784) <= not(layer8_outputs(936));
    outputs(4785) <= not(layer8_outputs(2635));
    outputs(4786) <= (layer8_outputs(4000)) xor (layer8_outputs(3160));
    outputs(4787) <= layer8_outputs(2637);
    outputs(4788) <= not(layer8_outputs(3782));
    outputs(4789) <= (layer8_outputs(4883)) and not (layer8_outputs(2701));
    outputs(4790) <= layer8_outputs(440);
    outputs(4791) <= (layer8_outputs(4708)) and not (layer8_outputs(2769));
    outputs(4792) <= not((layer8_outputs(1653)) xor (layer8_outputs(1196)));
    outputs(4793) <= layer8_outputs(1304);
    outputs(4794) <= not(layer8_outputs(1480));
    outputs(4795) <= (layer8_outputs(5000)) xor (layer8_outputs(3098));
    outputs(4796) <= layer8_outputs(4106);
    outputs(4797) <= layer8_outputs(1162);
    outputs(4798) <= layer8_outputs(1702);
    outputs(4799) <= not(layer8_outputs(1381));
    outputs(4800) <= not(layer8_outputs(4364));
    outputs(4801) <= not(layer8_outputs(3344));
    outputs(4802) <= not((layer8_outputs(3912)) or (layer8_outputs(1519)));
    outputs(4803) <= (layer8_outputs(4039)) xor (layer8_outputs(1268));
    outputs(4804) <= not((layer8_outputs(4317)) xor (layer8_outputs(42)));
    outputs(4805) <= not(layer8_outputs(3758));
    outputs(4806) <= not(layer8_outputs(1672));
    outputs(4807) <= not(layer8_outputs(4901));
    outputs(4808) <= layer8_outputs(1899);
    outputs(4809) <= not((layer8_outputs(2937)) xor (layer8_outputs(2837)));
    outputs(4810) <= layer8_outputs(3410);
    outputs(4811) <= not((layer8_outputs(1856)) xor (layer8_outputs(4400)));
    outputs(4812) <= not((layer8_outputs(3879)) xor (layer8_outputs(720)));
    outputs(4813) <= (layer8_outputs(4696)) and (layer8_outputs(2689));
    outputs(4814) <= not(layer8_outputs(1723));
    outputs(4815) <= not(layer8_outputs(921));
    outputs(4816) <= layer8_outputs(5060);
    outputs(4817) <= (layer8_outputs(4910)) and not (layer8_outputs(2461));
    outputs(4818) <= layer8_outputs(3194);
    outputs(4819) <= (layer8_outputs(2567)) xor (layer8_outputs(3674));
    outputs(4820) <= (layer8_outputs(3097)) xor (layer8_outputs(4227));
    outputs(4821) <= not((layer8_outputs(2554)) xor (layer8_outputs(4425)));
    outputs(4822) <= layer8_outputs(4603);
    outputs(4823) <= not((layer8_outputs(4967)) xor (layer8_outputs(4219)));
    outputs(4824) <= not(layer8_outputs(3431));
    outputs(4825) <= (layer8_outputs(964)) xor (layer8_outputs(348));
    outputs(4826) <= not(layer8_outputs(2066));
    outputs(4827) <= (layer8_outputs(2750)) xor (layer8_outputs(1503));
    outputs(4828) <= not(layer8_outputs(4306));
    outputs(4829) <= not(layer8_outputs(4393));
    outputs(4830) <= (layer8_outputs(4232)) xor (layer8_outputs(144));
    outputs(4831) <= layer8_outputs(3829);
    outputs(4832) <= (layer8_outputs(2207)) xor (layer8_outputs(2877));
    outputs(4833) <= not((layer8_outputs(3646)) xor (layer8_outputs(4619)));
    outputs(4834) <= (layer8_outputs(894)) and not (layer8_outputs(5069));
    outputs(4835) <= layer8_outputs(115);
    outputs(4836) <= not(layer8_outputs(1903));
    outputs(4837) <= not(layer8_outputs(207));
    outputs(4838) <= layer8_outputs(4883);
    outputs(4839) <= not((layer8_outputs(5028)) xor (layer8_outputs(3822)));
    outputs(4840) <= not(layer8_outputs(1105));
    outputs(4841) <= (layer8_outputs(3975)) and (layer8_outputs(3090));
    outputs(4842) <= not((layer8_outputs(2621)) xor (layer8_outputs(3104)));
    outputs(4843) <= layer8_outputs(2006);
    outputs(4844) <= layer8_outputs(1482);
    outputs(4845) <= layer8_outputs(3666);
    outputs(4846) <= not(layer8_outputs(3588));
    outputs(4847) <= not(layer8_outputs(301));
    outputs(4848) <= not((layer8_outputs(914)) and (layer8_outputs(99)));
    outputs(4849) <= not(layer8_outputs(3304));
    outputs(4850) <= layer8_outputs(781);
    outputs(4851) <= (layer8_outputs(2189)) xor (layer8_outputs(3663));
    outputs(4852) <= not(layer8_outputs(4952));
    outputs(4853) <= layer8_outputs(2545);
    outputs(4854) <= layer8_outputs(4343);
    outputs(4855) <= not(layer8_outputs(3520));
    outputs(4856) <= not(layer8_outputs(4892));
    outputs(4857) <= layer8_outputs(3511);
    outputs(4858) <= (layer8_outputs(2632)) xor (layer8_outputs(927));
    outputs(4859) <= layer8_outputs(758);
    outputs(4860) <= not(layer8_outputs(2613));
    outputs(4861) <= not((layer8_outputs(556)) xor (layer8_outputs(4480)));
    outputs(4862) <= (layer8_outputs(4062)) and (layer8_outputs(1852));
    outputs(4863) <= not(layer8_outputs(11));
    outputs(4864) <= (layer8_outputs(3012)) and not (layer8_outputs(4320));
    outputs(4865) <= not((layer8_outputs(2436)) xor (layer8_outputs(1393)));
    outputs(4866) <= layer8_outputs(173);
    outputs(4867) <= not(layer8_outputs(1417));
    outputs(4868) <= not((layer8_outputs(3821)) xor (layer8_outputs(4660)));
    outputs(4869) <= layer8_outputs(2137);
    outputs(4870) <= layer8_outputs(1658);
    outputs(4871) <= layer8_outputs(4234);
    outputs(4872) <= not((layer8_outputs(640)) xor (layer8_outputs(3598)));
    outputs(4873) <= not((layer8_outputs(4113)) xor (layer8_outputs(2991)));
    outputs(4874) <= (layer8_outputs(3923)) and not (layer8_outputs(3154));
    outputs(4875) <= (layer8_outputs(1371)) xor (layer8_outputs(1980));
    outputs(4876) <= not(layer8_outputs(3029));
    outputs(4877) <= layer8_outputs(54);
    outputs(4878) <= layer8_outputs(4039);
    outputs(4879) <= layer8_outputs(1130);
    outputs(4880) <= not(layer8_outputs(4266));
    outputs(4881) <= (layer8_outputs(1752)) and (layer8_outputs(216));
    outputs(4882) <= (layer8_outputs(3217)) xor (layer8_outputs(1615));
    outputs(4883) <= (layer8_outputs(3878)) xor (layer8_outputs(2598));
    outputs(4884) <= layer8_outputs(2240);
    outputs(4885) <= not(layer8_outputs(2003));
    outputs(4886) <= not((layer8_outputs(4618)) xor (layer8_outputs(2051)));
    outputs(4887) <= (layer8_outputs(1501)) xor (layer8_outputs(2432));
    outputs(4888) <= not(layer8_outputs(5012));
    outputs(4889) <= layer8_outputs(1457);
    outputs(4890) <= not((layer8_outputs(4691)) or (layer8_outputs(4713)));
    outputs(4891) <= not((layer8_outputs(4632)) or (layer8_outputs(2925)));
    outputs(4892) <= not((layer8_outputs(4269)) xor (layer8_outputs(2356)));
    outputs(4893) <= (layer8_outputs(4037)) and (layer8_outputs(1450));
    outputs(4894) <= layer8_outputs(2879);
    outputs(4895) <= layer8_outputs(437);
    outputs(4896) <= not(layer8_outputs(2894));
    outputs(4897) <= not((layer8_outputs(1886)) xor (layer8_outputs(3941)));
    outputs(4898) <= not(layer8_outputs(685));
    outputs(4899) <= (layer8_outputs(2251)) and not (layer8_outputs(2208));
    outputs(4900) <= not(layer8_outputs(3267));
    outputs(4901) <= not(layer8_outputs(1785));
    outputs(4902) <= not(layer8_outputs(1030));
    outputs(4903) <= (layer8_outputs(2596)) or (layer8_outputs(3601));
    outputs(4904) <= (layer8_outputs(695)) xor (layer8_outputs(1816));
    outputs(4905) <= not(layer8_outputs(4818));
    outputs(4906) <= not(layer8_outputs(1583));
    outputs(4907) <= layer8_outputs(4627);
    outputs(4908) <= not((layer8_outputs(3298)) or (layer8_outputs(3675)));
    outputs(4909) <= (layer8_outputs(3759)) xor (layer8_outputs(3386));
    outputs(4910) <= layer8_outputs(1589);
    outputs(4911) <= not(layer8_outputs(3794));
    outputs(4912) <= layer8_outputs(2655);
    outputs(4913) <= not(layer8_outputs(2648));
    outputs(4914) <= not(layer8_outputs(1571));
    outputs(4915) <= not(layer8_outputs(1232));
    outputs(4916) <= (layer8_outputs(4346)) xor (layer8_outputs(3842));
    outputs(4917) <= layer8_outputs(3093);
    outputs(4918) <= not((layer8_outputs(3802)) xor (layer8_outputs(935)));
    outputs(4919) <= (layer8_outputs(4903)) and not (layer8_outputs(228));
    outputs(4920) <= layer8_outputs(1562);
    outputs(4921) <= layer8_outputs(2868);
    outputs(4922) <= (layer8_outputs(3250)) and not (layer8_outputs(2044));
    outputs(4923) <= not(layer8_outputs(2346));
    outputs(4924) <= not(layer8_outputs(5118));
    outputs(4925) <= not((layer8_outputs(1446)) xor (layer8_outputs(1467)));
    outputs(4926) <= (layer8_outputs(19)) xor (layer8_outputs(2024));
    outputs(4927) <= (layer8_outputs(3459)) xor (layer8_outputs(3660));
    outputs(4928) <= (layer8_outputs(2859)) xor (layer8_outputs(4657));
    outputs(4929) <= layer8_outputs(2821);
    outputs(4930) <= layer8_outputs(2025);
    outputs(4931) <= not(layer8_outputs(4304));
    outputs(4932) <= layer8_outputs(4535);
    outputs(4933) <= layer8_outputs(1461);
    outputs(4934) <= layer8_outputs(2622);
    outputs(4935) <= not(layer8_outputs(2745));
    outputs(4936) <= layer8_outputs(2768);
    outputs(4937) <= layer8_outputs(20);
    outputs(4938) <= layer8_outputs(4629);
    outputs(4939) <= layer8_outputs(331);
    outputs(4940) <= (layer8_outputs(1314)) and not (layer8_outputs(4359));
    outputs(4941) <= layer8_outputs(2963);
    outputs(4942) <= (layer8_outputs(2922)) and (layer8_outputs(2695));
    outputs(4943) <= not((layer8_outputs(4574)) xor (layer8_outputs(498)));
    outputs(4944) <= not(layer8_outputs(3943)) or (layer8_outputs(4180));
    outputs(4945) <= not(layer8_outputs(4015));
    outputs(4946) <= not(layer8_outputs(3344));
    outputs(4947) <= layer8_outputs(4679);
    outputs(4948) <= layer8_outputs(3949);
    outputs(4949) <= not((layer8_outputs(4302)) xor (layer8_outputs(3687)));
    outputs(4950) <= (layer8_outputs(3168)) xor (layer8_outputs(5089));
    outputs(4951) <= not(layer8_outputs(4781));
    outputs(4952) <= layer8_outputs(3253);
    outputs(4953) <= (layer8_outputs(3194)) and not (layer8_outputs(2391));
    outputs(4954) <= layer8_outputs(2213);
    outputs(4955) <= (layer8_outputs(4185)) xor (layer8_outputs(686));
    outputs(4956) <= (layer8_outputs(1064)) xor (layer8_outputs(59));
    outputs(4957) <= layer8_outputs(395);
    outputs(4958) <= (layer8_outputs(1198)) and (layer8_outputs(4707));
    outputs(4959) <= not(layer8_outputs(3651));
    outputs(4960) <= not(layer8_outputs(46));
    outputs(4961) <= layer8_outputs(3159);
    outputs(4962) <= (layer8_outputs(4000)) and not (layer8_outputs(2777));
    outputs(4963) <= layer8_outputs(5017);
    outputs(4964) <= (layer8_outputs(4247)) xor (layer8_outputs(3466));
    outputs(4965) <= not(layer8_outputs(643));
    outputs(4966) <= not((layer8_outputs(1211)) xor (layer8_outputs(2010)));
    outputs(4967) <= layer8_outputs(1031);
    outputs(4968) <= (layer8_outputs(3039)) xor (layer8_outputs(2883));
    outputs(4969) <= layer8_outputs(2833);
    outputs(4970) <= layer8_outputs(4800);
    outputs(4971) <= not(layer8_outputs(4348));
    outputs(4972) <= layer8_outputs(313);
    outputs(4973) <= not(layer8_outputs(1509));
    outputs(4974) <= not(layer8_outputs(942));
    outputs(4975) <= not((layer8_outputs(2681)) xor (layer8_outputs(466)));
    outputs(4976) <= layer8_outputs(598);
    outputs(4977) <= layer8_outputs(1009);
    outputs(4978) <= (layer8_outputs(3971)) xor (layer8_outputs(1541));
    outputs(4979) <= layer8_outputs(820);
    outputs(4980) <= (layer8_outputs(2937)) xor (layer8_outputs(4791));
    outputs(4981) <= layer8_outputs(2298);
    outputs(4982) <= not(layer8_outputs(217));
    outputs(4983) <= layer8_outputs(3250);
    outputs(4984) <= layer8_outputs(4064);
    outputs(4985) <= (layer8_outputs(2311)) xor (layer8_outputs(2803));
    outputs(4986) <= not(layer8_outputs(347));
    outputs(4987) <= not(layer8_outputs(1248));
    outputs(4988) <= layer8_outputs(4465);
    outputs(4989) <= not((layer8_outputs(4615)) or (layer8_outputs(830)));
    outputs(4990) <= not(layer8_outputs(3227));
    outputs(4991) <= (layer8_outputs(4832)) and (layer8_outputs(1103));
    outputs(4992) <= not(layer8_outputs(363));
    outputs(4993) <= layer8_outputs(2831);
    outputs(4994) <= not((layer8_outputs(5096)) xor (layer8_outputs(2378)));
    outputs(4995) <= not(layer8_outputs(3314)) or (layer8_outputs(2978));
    outputs(4996) <= (layer8_outputs(33)) and (layer8_outputs(2729));
    outputs(4997) <= not((layer8_outputs(4356)) or (layer8_outputs(699)));
    outputs(4998) <= layer8_outputs(5095);
    outputs(4999) <= not(layer8_outputs(1711));
    outputs(5000) <= not(layer8_outputs(2230));
    outputs(5001) <= layer8_outputs(4284);
    outputs(5002) <= (layer8_outputs(4869)) xor (layer8_outputs(477));
    outputs(5003) <= (layer8_outputs(4620)) and (layer8_outputs(1575));
    outputs(5004) <= not((layer8_outputs(2082)) xor (layer8_outputs(4037)));
    outputs(5005) <= not((layer8_outputs(4628)) xor (layer8_outputs(675)));
    outputs(5006) <= (layer8_outputs(813)) and not (layer8_outputs(1215));
    outputs(5007) <= layer8_outputs(3524);
    outputs(5008) <= (layer8_outputs(5074)) and not (layer8_outputs(2426));
    outputs(5009) <= not(layer8_outputs(2957)) or (layer8_outputs(923));
    outputs(5010) <= (layer8_outputs(1892)) xor (layer8_outputs(3211));
    outputs(5011) <= not((layer8_outputs(429)) xor (layer8_outputs(4537)));
    outputs(5012) <= (layer8_outputs(1746)) xor (layer8_outputs(4110));
    outputs(5013) <= not((layer8_outputs(602)) xor (layer8_outputs(2336)));
    outputs(5014) <= layer8_outputs(4545);
    outputs(5015) <= (layer8_outputs(233)) xor (layer8_outputs(2040));
    outputs(5016) <= layer8_outputs(3738);
    outputs(5017) <= layer8_outputs(4491);
    outputs(5018) <= not((layer8_outputs(1662)) xor (layer8_outputs(4404)));
    outputs(5019) <= (layer8_outputs(2400)) and not (layer8_outputs(4747));
    outputs(5020) <= (layer8_outputs(794)) and not (layer8_outputs(1094));
    outputs(5021) <= (layer8_outputs(1591)) and not (layer8_outputs(4447));
    outputs(5022) <= (layer8_outputs(2735)) and (layer8_outputs(510));
    outputs(5023) <= (layer8_outputs(4887)) xor (layer8_outputs(2185));
    outputs(5024) <= not((layer8_outputs(776)) or (layer8_outputs(2276)));
    outputs(5025) <= not((layer8_outputs(4230)) xor (layer8_outputs(2239)));
    outputs(5026) <= not(layer8_outputs(4126));
    outputs(5027) <= (layer8_outputs(1885)) xor (layer8_outputs(2956));
    outputs(5028) <= not(layer8_outputs(4780));
    outputs(5029) <= not(layer8_outputs(1665));
    outputs(5030) <= (layer8_outputs(102)) xor (layer8_outputs(4886));
    outputs(5031) <= (layer8_outputs(2560)) and not (layer8_outputs(3796));
    outputs(5032) <= layer8_outputs(4065);
    outputs(5033) <= not(layer8_outputs(4494));
    outputs(5034) <= not(layer8_outputs(258));
    outputs(5035) <= not(layer8_outputs(411));
    outputs(5036) <= not(layer8_outputs(4634)) or (layer8_outputs(593));
    outputs(5037) <= not(layer8_outputs(347));
    outputs(5038) <= (layer8_outputs(3294)) and (layer8_outputs(2785));
    outputs(5039) <= layer8_outputs(1525);
    outputs(5040) <= not(layer8_outputs(1340));
    outputs(5041) <= not(layer8_outputs(2724));
    outputs(5042) <= not(layer8_outputs(2357));
    outputs(5043) <= layer8_outputs(575);
    outputs(5044) <= (layer8_outputs(1283)) xor (layer8_outputs(1457));
    outputs(5045) <= layer8_outputs(1670);
    outputs(5046) <= layer8_outputs(4949);
    outputs(5047) <= not(layer8_outputs(871));
    outputs(5048) <= layer8_outputs(2383);
    outputs(5049) <= (layer8_outputs(3696)) xor (layer8_outputs(2442));
    outputs(5050) <= not((layer8_outputs(2788)) xor (layer8_outputs(994)));
    outputs(5051) <= (layer8_outputs(264)) xor (layer8_outputs(4548));
    outputs(5052) <= (layer8_outputs(4894)) and not (layer8_outputs(2449));
    outputs(5053) <= layer8_outputs(3742);
    outputs(5054) <= layer8_outputs(2209);
    outputs(5055) <= (layer8_outputs(1932)) and not (layer8_outputs(4766));
    outputs(5056) <= layer8_outputs(2415);
    outputs(5057) <= not((layer8_outputs(4018)) xor (layer8_outputs(3735)));
    outputs(5058) <= not(layer8_outputs(415));
    outputs(5059) <= not((layer8_outputs(3580)) xor (layer8_outputs(1521)));
    outputs(5060) <= not((layer8_outputs(3159)) xor (layer8_outputs(4318)));
    outputs(5061) <= layer8_outputs(4672);
    outputs(5062) <= layer8_outputs(2406);
    outputs(5063) <= layer8_outputs(735);
    outputs(5064) <= not((layer8_outputs(3347)) xor (layer8_outputs(996)));
    outputs(5065) <= not((layer8_outputs(3022)) xor (layer8_outputs(1145)));
    outputs(5066) <= (layer8_outputs(3266)) xor (layer8_outputs(3333));
    outputs(5067) <= layer8_outputs(5041);
    outputs(5068) <= not((layer8_outputs(460)) or (layer8_outputs(9)));
    outputs(5069) <= not(layer8_outputs(3946));
    outputs(5070) <= not(layer8_outputs(3722));
    outputs(5071) <= not((layer8_outputs(187)) or (layer8_outputs(2818)));
    outputs(5072) <= layer8_outputs(3740);
    outputs(5073) <= layer8_outputs(4661);
    outputs(5074) <= not((layer8_outputs(2459)) xor (layer8_outputs(4511)));
    outputs(5075) <= not((layer8_outputs(1116)) xor (layer8_outputs(2020)));
    outputs(5076) <= not((layer8_outputs(2117)) xor (layer8_outputs(5034)));
    outputs(5077) <= not(layer8_outputs(729));
    outputs(5078) <= (layer8_outputs(1859)) or (layer8_outputs(1719));
    outputs(5079) <= layer8_outputs(3551);
    outputs(5080) <= layer8_outputs(4529);
    outputs(5081) <= layer8_outputs(341);
    outputs(5082) <= layer8_outputs(3920);
    outputs(5083) <= layer8_outputs(38);
    outputs(5084) <= not(layer8_outputs(1807));
    outputs(5085) <= (layer8_outputs(4017)) xor (layer8_outputs(3359));
    outputs(5086) <= layer8_outputs(1800);
    outputs(5087) <= not((layer8_outputs(5102)) or (layer8_outputs(2950)));
    outputs(5088) <= not((layer8_outputs(959)) xor (layer8_outputs(1455)));
    outputs(5089) <= not(layer8_outputs(3385)) or (layer8_outputs(2916));
    outputs(5090) <= layer8_outputs(521);
    outputs(5091) <= not(layer8_outputs(3295));
    outputs(5092) <= (layer8_outputs(4035)) xor (layer8_outputs(1506));
    outputs(5093) <= layer8_outputs(4642);
    outputs(5094) <= not(layer8_outputs(1604));
    outputs(5095) <= (layer8_outputs(1165)) and not (layer8_outputs(1295));
    outputs(5096) <= (layer8_outputs(2723)) and not (layer8_outputs(923));
    outputs(5097) <= (layer8_outputs(2193)) xor (layer8_outputs(4433));
    outputs(5098) <= layer8_outputs(361);
    outputs(5099) <= (layer8_outputs(3695)) or (layer8_outputs(3715));
    outputs(5100) <= layer8_outputs(3443);
    outputs(5101) <= not(layer8_outputs(4685));
    outputs(5102) <= layer8_outputs(489);
    outputs(5103) <= (layer8_outputs(1978)) and not (layer8_outputs(283));
    outputs(5104) <= layer8_outputs(3858);
    outputs(5105) <= (layer8_outputs(316)) xor (layer8_outputs(1194));
    outputs(5106) <= layer8_outputs(3601);
    outputs(5107) <= not(layer8_outputs(4879));
    outputs(5108) <= not((layer8_outputs(3083)) xor (layer8_outputs(4839)));
    outputs(5109) <= not(layer8_outputs(484));
    outputs(5110) <= layer8_outputs(4681);
    outputs(5111) <= not((layer8_outputs(1002)) xor (layer8_outputs(3027)));
    outputs(5112) <= layer8_outputs(3279);
    outputs(5113) <= not(layer8_outputs(3853));
    outputs(5114) <= not(layer8_outputs(1825));
    outputs(5115) <= (layer8_outputs(4378)) xor (layer8_outputs(4129));
    outputs(5116) <= layer8_outputs(3776);
    outputs(5117) <= (layer8_outputs(2606)) xor (layer8_outputs(1784));
    outputs(5118) <= layer8_outputs(3890);
    outputs(5119) <= not(layer8_outputs(294));

end Behavioral;
