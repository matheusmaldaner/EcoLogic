library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(7679 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(7679 downto 0);
    signal layer1_outputs : std_logic_vector(7679 downto 0);
    signal layer2_outputs : std_logic_vector(7679 downto 0);
    signal layer3_outputs : std_logic_vector(7679 downto 0);
    signal layer4_outputs : std_logic_vector(7679 downto 0);

begin

    layer0_outputs(0) <= inputs(43);
    layer0_outputs(1) <= inputs(99);
    layer0_outputs(2) <= inputs(159);
    layer0_outputs(3) <= not(inputs(16));
    layer0_outputs(4) <= '1';
    layer0_outputs(5) <= not(inputs(236));
    layer0_outputs(6) <= not(inputs(126));
    layer0_outputs(7) <= (inputs(152)) or (inputs(180));
    layer0_outputs(8) <= '1';
    layer0_outputs(9) <= (inputs(19)) or (inputs(155));
    layer0_outputs(10) <= inputs(101);
    layer0_outputs(11) <= (inputs(191)) or (inputs(150));
    layer0_outputs(12) <= (inputs(23)) and not (inputs(164));
    layer0_outputs(13) <= (inputs(128)) and not (inputs(181));
    layer0_outputs(14) <= (inputs(238)) or (inputs(254));
    layer0_outputs(15) <= not(inputs(98));
    layer0_outputs(16) <= not(inputs(230));
    layer0_outputs(17) <= not((inputs(60)) xor (inputs(28)));
    layer0_outputs(18) <= not((inputs(76)) xor (inputs(144)));
    layer0_outputs(19) <= inputs(72);
    layer0_outputs(20) <= (inputs(51)) or (inputs(75));
    layer0_outputs(21) <= not((inputs(167)) or (inputs(169)));
    layer0_outputs(22) <= not(inputs(1));
    layer0_outputs(23) <= (inputs(50)) and not (inputs(18));
    layer0_outputs(24) <= inputs(50);
    layer0_outputs(25) <= not((inputs(105)) or (inputs(253)));
    layer0_outputs(26) <= (inputs(248)) and (inputs(255));
    layer0_outputs(27) <= (inputs(226)) or (inputs(239));
    layer0_outputs(28) <= not(inputs(87));
    layer0_outputs(29) <= (inputs(220)) xor (inputs(187));
    layer0_outputs(30) <= '1';
    layer0_outputs(31) <= (inputs(219)) and (inputs(242));
    layer0_outputs(32) <= not(inputs(83)) or (inputs(231));
    layer0_outputs(33) <= inputs(162);
    layer0_outputs(34) <= (inputs(37)) or (inputs(25));
    layer0_outputs(35) <= not(inputs(124)) or (inputs(144));
    layer0_outputs(36) <= '0';
    layer0_outputs(37) <= '0';
    layer0_outputs(38) <= not((inputs(188)) or (inputs(85)));
    layer0_outputs(39) <= not(inputs(30)) or (inputs(61));
    layer0_outputs(40) <= (inputs(246)) and (inputs(168));
    layer0_outputs(41) <= '1';
    layer0_outputs(42) <= not((inputs(85)) or (inputs(33)));
    layer0_outputs(43) <= not(inputs(76));
    layer0_outputs(44) <= not(inputs(53)) or (inputs(168));
    layer0_outputs(45) <= not(inputs(148));
    layer0_outputs(46) <= inputs(143);
    layer0_outputs(47) <= not((inputs(147)) and (inputs(141)));
    layer0_outputs(48) <= not(inputs(89));
    layer0_outputs(49) <= (inputs(198)) and (inputs(240));
    layer0_outputs(50) <= not((inputs(202)) or (inputs(27)));
    layer0_outputs(51) <= inputs(114);
    layer0_outputs(52) <= inputs(204);
    layer0_outputs(53) <= (inputs(82)) or (inputs(143));
    layer0_outputs(54) <= (inputs(154)) or (inputs(128));
    layer0_outputs(55) <= (inputs(104)) and not (inputs(18));
    layer0_outputs(56) <= not((inputs(115)) and (inputs(36)));
    layer0_outputs(57) <= not(inputs(132));
    layer0_outputs(58) <= not((inputs(14)) or (inputs(255)));
    layer0_outputs(59) <= not((inputs(75)) xor (inputs(28)));
    layer0_outputs(60) <= inputs(146);
    layer0_outputs(61) <= not((inputs(237)) or (inputs(147)));
    layer0_outputs(62) <= not((inputs(172)) xor (inputs(220)));
    layer0_outputs(63) <= not(inputs(140));
    layer0_outputs(64) <= not((inputs(213)) and (inputs(169)));
    layer0_outputs(65) <= not(inputs(25));
    layer0_outputs(66) <= not(inputs(255));
    layer0_outputs(67) <= inputs(42);
    layer0_outputs(68) <= not((inputs(241)) xor (inputs(224)));
    layer0_outputs(69) <= not(inputs(35)) or (inputs(58));
    layer0_outputs(70) <= not((inputs(99)) or (inputs(152)));
    layer0_outputs(71) <= (inputs(196)) or (inputs(6));
    layer0_outputs(72) <= '1';
    layer0_outputs(73) <= inputs(189);
    layer0_outputs(74) <= '0';
    layer0_outputs(75) <= not((inputs(88)) or (inputs(110)));
    layer0_outputs(76) <= (inputs(28)) xor (inputs(3));
    layer0_outputs(77) <= '0';
    layer0_outputs(78) <= not(inputs(33));
    layer0_outputs(79) <= not(inputs(197)) or (inputs(33));
    layer0_outputs(80) <= (inputs(154)) and not (inputs(174));
    layer0_outputs(81) <= (inputs(74)) or (inputs(135));
    layer0_outputs(82) <= not(inputs(42)) or (inputs(171));
    layer0_outputs(83) <= not((inputs(103)) or (inputs(64)));
    layer0_outputs(84) <= not(inputs(127));
    layer0_outputs(85) <= '1';
    layer0_outputs(86) <= not((inputs(248)) and (inputs(80)));
    layer0_outputs(87) <= not((inputs(176)) or (inputs(216)));
    layer0_outputs(88) <= (inputs(9)) xor (inputs(57));
    layer0_outputs(89) <= not(inputs(161));
    layer0_outputs(90) <= not((inputs(31)) xor (inputs(127)));
    layer0_outputs(91) <= '0';
    layer0_outputs(92) <= (inputs(210)) and (inputs(160));
    layer0_outputs(93) <= (inputs(149)) or (inputs(96));
    layer0_outputs(94) <= (inputs(178)) or (inputs(19));
    layer0_outputs(95) <= not(inputs(221)) or (inputs(107));
    layer0_outputs(96) <= not(inputs(67)) or (inputs(156));
    layer0_outputs(97) <= not((inputs(21)) or (inputs(22)));
    layer0_outputs(98) <= inputs(62);
    layer0_outputs(99) <= (inputs(178)) and not (inputs(178));
    layer0_outputs(100) <= (inputs(160)) and not (inputs(232));
    layer0_outputs(101) <= inputs(77);
    layer0_outputs(102) <= (inputs(157)) or (inputs(234));
    layer0_outputs(103) <= '1';
    layer0_outputs(104) <= not(inputs(217)) or (inputs(255));
    layer0_outputs(105) <= not((inputs(163)) xor (inputs(32)));
    layer0_outputs(106) <= not((inputs(194)) and (inputs(177)));
    layer0_outputs(107) <= inputs(36);
    layer0_outputs(108) <= '1';
    layer0_outputs(109) <= inputs(188);
    layer0_outputs(110) <= inputs(135);
    layer0_outputs(111) <= (inputs(68)) and not (inputs(87));
    layer0_outputs(112) <= not((inputs(52)) and (inputs(237)));
    layer0_outputs(113) <= '0';
    layer0_outputs(114) <= (inputs(83)) and not (inputs(162));
    layer0_outputs(115) <= not(inputs(28));
    layer0_outputs(116) <= (inputs(218)) and not (inputs(65));
    layer0_outputs(117) <= (inputs(206)) or (inputs(65));
    layer0_outputs(118) <= '0';
    layer0_outputs(119) <= '1';
    layer0_outputs(120) <= not(inputs(194));
    layer0_outputs(121) <= (inputs(50)) or (inputs(65));
    layer0_outputs(122) <= not((inputs(59)) and (inputs(114)));
    layer0_outputs(123) <= not(inputs(92)) or (inputs(50));
    layer0_outputs(124) <= inputs(177);
    layer0_outputs(125) <= inputs(24);
    layer0_outputs(126) <= (inputs(245)) and not (inputs(183));
    layer0_outputs(127) <= not((inputs(104)) xor (inputs(173)));
    layer0_outputs(128) <= inputs(197);
    layer0_outputs(129) <= '1';
    layer0_outputs(130) <= not(inputs(94));
    layer0_outputs(131) <= '1';
    layer0_outputs(132) <= (inputs(237)) and not (inputs(177));
    layer0_outputs(133) <= not(inputs(101));
    layer0_outputs(134) <= not((inputs(209)) and (inputs(0)));
    layer0_outputs(135) <= '0';
    layer0_outputs(136) <= not((inputs(86)) xor (inputs(115)));
    layer0_outputs(137) <= inputs(74);
    layer0_outputs(138) <= not(inputs(143));
    layer0_outputs(139) <= inputs(177);
    layer0_outputs(140) <= not((inputs(28)) or (inputs(69)));
    layer0_outputs(141) <= (inputs(225)) and (inputs(99));
    layer0_outputs(142) <= not((inputs(132)) or (inputs(230)));
    layer0_outputs(143) <= inputs(46);
    layer0_outputs(144) <= not(inputs(58)) or (inputs(120));
    layer0_outputs(145) <= not((inputs(93)) or (inputs(9)));
    layer0_outputs(146) <= '1';
    layer0_outputs(147) <= not((inputs(226)) or (inputs(210)));
    layer0_outputs(148) <= (inputs(89)) or (inputs(31));
    layer0_outputs(149) <= inputs(235);
    layer0_outputs(150) <= (inputs(245)) and (inputs(254));
    layer0_outputs(151) <= not(inputs(55));
    layer0_outputs(152) <= inputs(123);
    layer0_outputs(153) <= not((inputs(49)) or (inputs(14)));
    layer0_outputs(154) <= '0';
    layer0_outputs(155) <= not((inputs(233)) or (inputs(87)));
    layer0_outputs(156) <= inputs(126);
    layer0_outputs(157) <= (inputs(105)) and not (inputs(169));
    layer0_outputs(158) <= not((inputs(130)) or (inputs(193)));
    layer0_outputs(159) <= (inputs(51)) and (inputs(125));
    layer0_outputs(160) <= not(inputs(116));
    layer0_outputs(161) <= (inputs(250)) and not (inputs(65));
    layer0_outputs(162) <= not(inputs(83)) or (inputs(236));
    layer0_outputs(163) <= not(inputs(102));
    layer0_outputs(164) <= not(inputs(39));
    layer0_outputs(165) <= inputs(119);
    layer0_outputs(166) <= inputs(110);
    layer0_outputs(167) <= not((inputs(115)) or (inputs(144)));
    layer0_outputs(168) <= '1';
    layer0_outputs(169) <= not(inputs(214));
    layer0_outputs(170) <= not(inputs(71));
    layer0_outputs(171) <= not(inputs(98)) or (inputs(61));
    layer0_outputs(172) <= (inputs(212)) and (inputs(253));
    layer0_outputs(173) <= not(inputs(168));
    layer0_outputs(174) <= not(inputs(34));
    layer0_outputs(175) <= inputs(77);
    layer0_outputs(176) <= not(inputs(10));
    layer0_outputs(177) <= inputs(225);
    layer0_outputs(178) <= inputs(231);
    layer0_outputs(179) <= not(inputs(213)) or (inputs(102));
    layer0_outputs(180) <= not(inputs(77));
    layer0_outputs(181) <= not((inputs(206)) or (inputs(134)));
    layer0_outputs(182) <= inputs(56);
    layer0_outputs(183) <= (inputs(208)) and (inputs(35));
    layer0_outputs(184) <= '1';
    layer0_outputs(185) <= not(inputs(238));
    layer0_outputs(186) <= not((inputs(241)) or (inputs(210)));
    layer0_outputs(187) <= (inputs(47)) xor (inputs(73));
    layer0_outputs(188) <= (inputs(154)) or (inputs(161));
    layer0_outputs(189) <= not((inputs(20)) xor (inputs(255)));
    layer0_outputs(190) <= (inputs(96)) or (inputs(147));
    layer0_outputs(191) <= not(inputs(206)) or (inputs(154));
    layer0_outputs(192) <= not(inputs(165));
    layer0_outputs(193) <= not((inputs(210)) and (inputs(35)));
    layer0_outputs(194) <= '1';
    layer0_outputs(195) <= not((inputs(208)) or (inputs(73)));
    layer0_outputs(196) <= (inputs(179)) and not (inputs(48));
    layer0_outputs(197) <= not((inputs(227)) or (inputs(170)));
    layer0_outputs(198) <= not(inputs(229)) or (inputs(20));
    layer0_outputs(199) <= '0';
    layer0_outputs(200) <= '1';
    layer0_outputs(201) <= not(inputs(65)) or (inputs(80));
    layer0_outputs(202) <= inputs(90);
    layer0_outputs(203) <= not(inputs(203));
    layer0_outputs(204) <= inputs(44);
    layer0_outputs(205) <= not((inputs(249)) or (inputs(7)));
    layer0_outputs(206) <= not(inputs(21));
    layer0_outputs(207) <= not((inputs(164)) or (inputs(206)));
    layer0_outputs(208) <= inputs(238);
    layer0_outputs(209) <= inputs(95);
    layer0_outputs(210) <= (inputs(135)) and not (inputs(27));
    layer0_outputs(211) <= not(inputs(129)) or (inputs(201));
    layer0_outputs(212) <= not((inputs(186)) and (inputs(243)));
    layer0_outputs(213) <= not(inputs(194));
    layer0_outputs(214) <= '0';
    layer0_outputs(215) <= (inputs(147)) and not (inputs(79));
    layer0_outputs(216) <= (inputs(158)) or (inputs(231));
    layer0_outputs(217) <= not(inputs(160));
    layer0_outputs(218) <= (inputs(3)) or (inputs(150));
    layer0_outputs(219) <= not(inputs(185));
    layer0_outputs(220) <= not(inputs(2));
    layer0_outputs(221) <= (inputs(166)) and (inputs(83));
    layer0_outputs(222) <= not((inputs(209)) or (inputs(98)));
    layer0_outputs(223) <= '0';
    layer0_outputs(224) <= (inputs(204)) and not (inputs(197));
    layer0_outputs(225) <= not((inputs(66)) or (inputs(148)));
    layer0_outputs(226) <= (inputs(13)) and (inputs(9));
    layer0_outputs(227) <= not(inputs(109)) or (inputs(133));
    layer0_outputs(228) <= '1';
    layer0_outputs(229) <= not(inputs(91));
    layer0_outputs(230) <= inputs(104);
    layer0_outputs(231) <= (inputs(94)) and (inputs(159));
    layer0_outputs(232) <= inputs(135);
    layer0_outputs(233) <= not(inputs(9));
    layer0_outputs(234) <= not(inputs(239));
    layer0_outputs(235) <= (inputs(149)) xor (inputs(248));
    layer0_outputs(236) <= inputs(51);
    layer0_outputs(237) <= '0';
    layer0_outputs(238) <= (inputs(252)) and (inputs(223));
    layer0_outputs(239) <= inputs(201);
    layer0_outputs(240) <= not((inputs(41)) and (inputs(108)));
    layer0_outputs(241) <= not((inputs(133)) or (inputs(100)));
    layer0_outputs(242) <= not((inputs(224)) xor (inputs(101)));
    layer0_outputs(243) <= inputs(162);
    layer0_outputs(244) <= inputs(59);
    layer0_outputs(245) <= '0';
    layer0_outputs(246) <= '1';
    layer0_outputs(247) <= (inputs(2)) and not (inputs(82));
    layer0_outputs(248) <= '0';
    layer0_outputs(249) <= (inputs(158)) or (inputs(72));
    layer0_outputs(250) <= not(inputs(22)) or (inputs(219));
    layer0_outputs(251) <= (inputs(108)) or (inputs(98));
    layer0_outputs(252) <= '1';
    layer0_outputs(253) <= (inputs(249)) or (inputs(103));
    layer0_outputs(254) <= (inputs(31)) and not (inputs(174));
    layer0_outputs(255) <= not(inputs(36)) or (inputs(158));
    layer0_outputs(256) <= inputs(237);
    layer0_outputs(257) <= inputs(190);
    layer0_outputs(258) <= inputs(178);
    layer0_outputs(259) <= (inputs(145)) and not (inputs(31));
    layer0_outputs(260) <= (inputs(167)) or (inputs(102));
    layer0_outputs(261) <= '1';
    layer0_outputs(262) <= not(inputs(139)) or (inputs(41));
    layer0_outputs(263) <= not(inputs(172));
    layer0_outputs(264) <= (inputs(8)) and not (inputs(216));
    layer0_outputs(265) <= not((inputs(9)) xor (inputs(205)));
    layer0_outputs(266) <= (inputs(61)) and (inputs(15));
    layer0_outputs(267) <= not(inputs(122)) or (inputs(190));
    layer0_outputs(268) <= not(inputs(33));
    layer0_outputs(269) <= inputs(108);
    layer0_outputs(270) <= not((inputs(204)) and (inputs(5)));
    layer0_outputs(271) <= (inputs(121)) and not (inputs(7));
    layer0_outputs(272) <= inputs(195);
    layer0_outputs(273) <= not(inputs(155)) or (inputs(90));
    layer0_outputs(274) <= (inputs(193)) or (inputs(119));
    layer0_outputs(275) <= inputs(127);
    layer0_outputs(276) <= (inputs(138)) or (inputs(247));
    layer0_outputs(277) <= not(inputs(129));
    layer0_outputs(278) <= (inputs(135)) and not (inputs(253));
    layer0_outputs(279) <= not((inputs(219)) xor (inputs(145)));
    layer0_outputs(280) <= (inputs(16)) and (inputs(72));
    layer0_outputs(281) <= not(inputs(49)) or (inputs(199));
    layer0_outputs(282) <= (inputs(10)) and not (inputs(26));
    layer0_outputs(283) <= not((inputs(217)) and (inputs(18)));
    layer0_outputs(284) <= inputs(143);
    layer0_outputs(285) <= not((inputs(140)) or (inputs(216)));
    layer0_outputs(286) <= (inputs(143)) or (inputs(198));
    layer0_outputs(287) <= (inputs(217)) or (inputs(125));
    layer0_outputs(288) <= (inputs(71)) and (inputs(116));
    layer0_outputs(289) <= not((inputs(218)) and (inputs(138)));
    layer0_outputs(290) <= (inputs(119)) and not (inputs(98));
    layer0_outputs(291) <= (inputs(52)) or (inputs(113));
    layer0_outputs(292) <= inputs(132);
    layer0_outputs(293) <= (inputs(60)) and not (inputs(69));
    layer0_outputs(294) <= not(inputs(130));
    layer0_outputs(295) <= not(inputs(100));
    layer0_outputs(296) <= not((inputs(140)) or (inputs(144)));
    layer0_outputs(297) <= '0';
    layer0_outputs(298) <= not((inputs(11)) or (inputs(22)));
    layer0_outputs(299) <= inputs(75);
    layer0_outputs(300) <= not((inputs(89)) and (inputs(102)));
    layer0_outputs(301) <= not(inputs(84));
    layer0_outputs(302) <= '0';
    layer0_outputs(303) <= '1';
    layer0_outputs(304) <= (inputs(245)) or (inputs(243));
    layer0_outputs(305) <= inputs(189);
    layer0_outputs(306) <= not(inputs(6)) or (inputs(53));
    layer0_outputs(307) <= (inputs(236)) or (inputs(221));
    layer0_outputs(308) <= (inputs(174)) or (inputs(118));
    layer0_outputs(309) <= inputs(254);
    layer0_outputs(310) <= inputs(49);
    layer0_outputs(311) <= inputs(101);
    layer0_outputs(312) <= inputs(125);
    layer0_outputs(313) <= not(inputs(74));
    layer0_outputs(314) <= (inputs(246)) or (inputs(144));
    layer0_outputs(315) <= not(inputs(229));
    layer0_outputs(316) <= not((inputs(156)) xor (inputs(190)));
    layer0_outputs(317) <= inputs(245);
    layer0_outputs(318) <= (inputs(254)) xor (inputs(19));
    layer0_outputs(319) <= not((inputs(122)) or (inputs(81)));
    layer0_outputs(320) <= not((inputs(207)) and (inputs(187)));
    layer0_outputs(321) <= not(inputs(55));
    layer0_outputs(322) <= '0';
    layer0_outputs(323) <= not(inputs(2)) or (inputs(219));
    layer0_outputs(324) <= '1';
    layer0_outputs(325) <= inputs(59);
    layer0_outputs(326) <= not(inputs(7)) or (inputs(13));
    layer0_outputs(327) <= '1';
    layer0_outputs(328) <= (inputs(65)) and not (inputs(235));
    layer0_outputs(329) <= '0';
    layer0_outputs(330) <= (inputs(38)) xor (inputs(217));
    layer0_outputs(331) <= not((inputs(9)) and (inputs(44)));
    layer0_outputs(332) <= '1';
    layer0_outputs(333) <= inputs(187);
    layer0_outputs(334) <= inputs(119);
    layer0_outputs(335) <= (inputs(243)) and not (inputs(90));
    layer0_outputs(336) <= inputs(18);
    layer0_outputs(337) <= not(inputs(152));
    layer0_outputs(338) <= inputs(250);
    layer0_outputs(339) <= not((inputs(81)) xor (inputs(84)));
    layer0_outputs(340) <= (inputs(162)) or (inputs(182));
    layer0_outputs(341) <= '0';
    layer0_outputs(342) <= not(inputs(10)) or (inputs(116));
    layer0_outputs(343) <= not(inputs(121));
    layer0_outputs(344) <= not(inputs(120)) or (inputs(138));
    layer0_outputs(345) <= not(inputs(246));
    layer0_outputs(346) <= inputs(98);
    layer0_outputs(347) <= not(inputs(109)) or (inputs(175));
    layer0_outputs(348) <= not((inputs(57)) or (inputs(26)));
    layer0_outputs(349) <= not(inputs(58)) or (inputs(162));
    layer0_outputs(350) <= (inputs(144)) or (inputs(240));
    layer0_outputs(351) <= not(inputs(34));
    layer0_outputs(352) <= not((inputs(77)) or (inputs(233)));
    layer0_outputs(353) <= not(inputs(247)) or (inputs(49));
    layer0_outputs(354) <= inputs(148);
    layer0_outputs(355) <= (inputs(27)) and not (inputs(58));
    layer0_outputs(356) <= not(inputs(186));
    layer0_outputs(357) <= not((inputs(6)) or (inputs(227)));
    layer0_outputs(358) <= inputs(190);
    layer0_outputs(359) <= not((inputs(23)) or (inputs(233)));
    layer0_outputs(360) <= (inputs(132)) and not (inputs(89));
    layer0_outputs(361) <= not(inputs(250)) or (inputs(51));
    layer0_outputs(362) <= not(inputs(84));
    layer0_outputs(363) <= not(inputs(72)) or (inputs(142));
    layer0_outputs(364) <= '1';
    layer0_outputs(365) <= (inputs(97)) and not (inputs(139));
    layer0_outputs(366) <= not(inputs(73));
    layer0_outputs(367) <= not((inputs(233)) or (inputs(246)));
    layer0_outputs(368) <= inputs(81);
    layer0_outputs(369) <= (inputs(175)) or (inputs(192));
    layer0_outputs(370) <= '1';
    layer0_outputs(371) <= not((inputs(78)) xor (inputs(3)));
    layer0_outputs(372) <= not(inputs(117));
    layer0_outputs(373) <= not(inputs(162));
    layer0_outputs(374) <= not((inputs(79)) or (inputs(101)));
    layer0_outputs(375) <= (inputs(107)) and not (inputs(147));
    layer0_outputs(376) <= not(inputs(40));
    layer0_outputs(377) <= not(inputs(165));
    layer0_outputs(378) <= '0';
    layer0_outputs(379) <= not(inputs(35));
    layer0_outputs(380) <= not((inputs(190)) and (inputs(201)));
    layer0_outputs(381) <= inputs(211);
    layer0_outputs(382) <= (inputs(215)) and not (inputs(34));
    layer0_outputs(383) <= inputs(87);
    layer0_outputs(384) <= not(inputs(196));
    layer0_outputs(385) <= (inputs(6)) and (inputs(6));
    layer0_outputs(386) <= '0';
    layer0_outputs(387) <= '1';
    layer0_outputs(388) <= (inputs(201)) xor (inputs(182));
    layer0_outputs(389) <= not((inputs(73)) and (inputs(251)));
    layer0_outputs(390) <= not((inputs(201)) or (inputs(53)));
    layer0_outputs(391) <= inputs(114);
    layer0_outputs(392) <= not(inputs(144));
    layer0_outputs(393) <= (inputs(179)) or (inputs(236));
    layer0_outputs(394) <= (inputs(113)) and not (inputs(133));
    layer0_outputs(395) <= not(inputs(76));
    layer0_outputs(396) <= (inputs(55)) and not (inputs(20));
    layer0_outputs(397) <= (inputs(242)) or (inputs(49));
    layer0_outputs(398) <= not(inputs(66));
    layer0_outputs(399) <= inputs(194);
    layer0_outputs(400) <= not(inputs(54)) or (inputs(182));
    layer0_outputs(401) <= (inputs(222)) or (inputs(151));
    layer0_outputs(402) <= inputs(192);
    layer0_outputs(403) <= (inputs(32)) or (inputs(213));
    layer0_outputs(404) <= not(inputs(164));
    layer0_outputs(405) <= (inputs(212)) or (inputs(4));
    layer0_outputs(406) <= inputs(127);
    layer0_outputs(407) <= (inputs(183)) and not (inputs(73));
    layer0_outputs(408) <= not(inputs(211));
    layer0_outputs(409) <= (inputs(250)) and not (inputs(107));
    layer0_outputs(410) <= not(inputs(197));
    layer0_outputs(411) <= (inputs(199)) xor (inputs(162));
    layer0_outputs(412) <= not((inputs(253)) xor (inputs(48)));
    layer0_outputs(413) <= not(inputs(238));
    layer0_outputs(414) <= inputs(238);
    layer0_outputs(415) <= not(inputs(63)) or (inputs(64));
    layer0_outputs(416) <= '0';
    layer0_outputs(417) <= not(inputs(134));
    layer0_outputs(418) <= not(inputs(26)) or (inputs(141));
    layer0_outputs(419) <= (inputs(27)) and not (inputs(251));
    layer0_outputs(420) <= not(inputs(162));
    layer0_outputs(421) <= '0';
    layer0_outputs(422) <= inputs(122);
    layer0_outputs(423) <= (inputs(245)) and not (inputs(142));
    layer0_outputs(424) <= (inputs(27)) or (inputs(52));
    layer0_outputs(425) <= (inputs(198)) or (inputs(239));
    layer0_outputs(426) <= not(inputs(17));
    layer0_outputs(427) <= inputs(100);
    layer0_outputs(428) <= (inputs(47)) and not (inputs(129));
    layer0_outputs(429) <= not(inputs(22));
    layer0_outputs(430) <= (inputs(213)) or (inputs(63));
    layer0_outputs(431) <= (inputs(196)) or (inputs(254));
    layer0_outputs(432) <= not((inputs(255)) or (inputs(201)));
    layer0_outputs(433) <= (inputs(14)) xor (inputs(107));
    layer0_outputs(434) <= '0';
    layer0_outputs(435) <= (inputs(6)) or (inputs(196));
    layer0_outputs(436) <= not(inputs(246));
    layer0_outputs(437) <= not((inputs(145)) or (inputs(2)));
    layer0_outputs(438) <= inputs(82);
    layer0_outputs(439) <= not(inputs(30)) or (inputs(197));
    layer0_outputs(440) <= (inputs(180)) and not (inputs(140));
    layer0_outputs(441) <= inputs(59);
    layer0_outputs(442) <= not(inputs(231));
    layer0_outputs(443) <= '1';
    layer0_outputs(444) <= not(inputs(41)) or (inputs(255));
    layer0_outputs(445) <= not(inputs(149)) or (inputs(74));
    layer0_outputs(446) <= '1';
    layer0_outputs(447) <= inputs(8);
    layer0_outputs(448) <= not(inputs(31));
    layer0_outputs(449) <= not(inputs(196)) or (inputs(93));
    layer0_outputs(450) <= (inputs(160)) and not (inputs(212));
    layer0_outputs(451) <= not(inputs(39)) or (inputs(87));
    layer0_outputs(452) <= inputs(163);
    layer0_outputs(453) <= inputs(179);
    layer0_outputs(454) <= not(inputs(36)) or (inputs(250));
    layer0_outputs(455) <= not((inputs(117)) or (inputs(132)));
    layer0_outputs(456) <= (inputs(7)) and not (inputs(18));
    layer0_outputs(457) <= not(inputs(212));
    layer0_outputs(458) <= inputs(186);
    layer0_outputs(459) <= (inputs(225)) xor (inputs(231));
    layer0_outputs(460) <= (inputs(127)) or (inputs(166));
    layer0_outputs(461) <= (inputs(237)) or (inputs(53));
    layer0_outputs(462) <= not((inputs(165)) and (inputs(213)));
    layer0_outputs(463) <= (inputs(51)) or (inputs(61));
    layer0_outputs(464) <= inputs(73);
    layer0_outputs(465) <= not((inputs(204)) or (inputs(40)));
    layer0_outputs(466) <= (inputs(30)) and (inputs(126));
    layer0_outputs(467) <= (inputs(19)) xor (inputs(156));
    layer0_outputs(468) <= inputs(228);
    layer0_outputs(469) <= not(inputs(40)) or (inputs(251));
    layer0_outputs(470) <= inputs(89);
    layer0_outputs(471) <= not(inputs(102)) or (inputs(241));
    layer0_outputs(472) <= (inputs(232)) and not (inputs(0));
    layer0_outputs(473) <= not(inputs(197));
    layer0_outputs(474) <= (inputs(193)) or (inputs(214));
    layer0_outputs(475) <= inputs(79);
    layer0_outputs(476) <= inputs(193);
    layer0_outputs(477) <= not(inputs(60)) or (inputs(73));
    layer0_outputs(478) <= inputs(120);
    layer0_outputs(479) <= not(inputs(135));
    layer0_outputs(480) <= (inputs(23)) and not (inputs(184));
    layer0_outputs(481) <= not(inputs(26));
    layer0_outputs(482) <= (inputs(9)) xor (inputs(189));
    layer0_outputs(483) <= inputs(229);
    layer0_outputs(484) <= (inputs(141)) and not (inputs(155));
    layer0_outputs(485) <= '1';
    layer0_outputs(486) <= not((inputs(145)) and (inputs(192)));
    layer0_outputs(487) <= not(inputs(54));
    layer0_outputs(488) <= not(inputs(128));
    layer0_outputs(489) <= not(inputs(158)) or (inputs(131));
    layer0_outputs(490) <= not(inputs(129));
    layer0_outputs(491) <= not((inputs(107)) or (inputs(157)));
    layer0_outputs(492) <= (inputs(32)) or (inputs(106));
    layer0_outputs(493) <= (inputs(40)) and not (inputs(252));
    layer0_outputs(494) <= (inputs(237)) and (inputs(93));
    layer0_outputs(495) <= inputs(161);
    layer0_outputs(496) <= (inputs(29)) or (inputs(46));
    layer0_outputs(497) <= not((inputs(109)) or (inputs(191)));
    layer0_outputs(498) <= not((inputs(229)) or (inputs(16)));
    layer0_outputs(499) <= (inputs(158)) and not (inputs(151));
    layer0_outputs(500) <= not((inputs(111)) or (inputs(56)));
    layer0_outputs(501) <= not(inputs(60)) or (inputs(251));
    layer0_outputs(502) <= (inputs(95)) or (inputs(61));
    layer0_outputs(503) <= '1';
    layer0_outputs(504) <= '1';
    layer0_outputs(505) <= not((inputs(59)) xor (inputs(135)));
    layer0_outputs(506) <= not(inputs(42));
    layer0_outputs(507) <= (inputs(223)) and not (inputs(7));
    layer0_outputs(508) <= '1';
    layer0_outputs(509) <= not(inputs(197));
    layer0_outputs(510) <= (inputs(65)) or (inputs(95));
    layer0_outputs(511) <= inputs(135);
    layer0_outputs(512) <= inputs(179);
    layer0_outputs(513) <= (inputs(189)) and not (inputs(239));
    layer0_outputs(514) <= inputs(94);
    layer0_outputs(515) <= (inputs(3)) and not (inputs(107));
    layer0_outputs(516) <= (inputs(242)) and not (inputs(128));
    layer0_outputs(517) <= (inputs(16)) xor (inputs(90));
    layer0_outputs(518) <= not((inputs(148)) or (inputs(94)));
    layer0_outputs(519) <= not(inputs(233)) or (inputs(158));
    layer0_outputs(520) <= (inputs(206)) or (inputs(151));
    layer0_outputs(521) <= '0';
    layer0_outputs(522) <= inputs(37);
    layer0_outputs(523) <= '0';
    layer0_outputs(524) <= not(inputs(83));
    layer0_outputs(525) <= not((inputs(235)) xor (inputs(161)));
    layer0_outputs(526) <= (inputs(66)) and not (inputs(207));
    layer0_outputs(527) <= (inputs(164)) or (inputs(218));
    layer0_outputs(528) <= not(inputs(167));
    layer0_outputs(529) <= '1';
    layer0_outputs(530) <= not((inputs(168)) or (inputs(182)));
    layer0_outputs(531) <= not((inputs(224)) or (inputs(6)));
    layer0_outputs(532) <= not((inputs(193)) or (inputs(56)));
    layer0_outputs(533) <= not((inputs(155)) and (inputs(20)));
    layer0_outputs(534) <= (inputs(78)) and (inputs(65));
    layer0_outputs(535) <= not(inputs(180)) or (inputs(170));
    layer0_outputs(536) <= not(inputs(199)) or (inputs(31));
    layer0_outputs(537) <= (inputs(45)) and not (inputs(161));
    layer0_outputs(538) <= inputs(181);
    layer0_outputs(539) <= inputs(145);
    layer0_outputs(540) <= (inputs(115)) and (inputs(115));
    layer0_outputs(541) <= inputs(72);
    layer0_outputs(542) <= '0';
    layer0_outputs(543) <= not(inputs(61));
    layer0_outputs(544) <= (inputs(131)) or (inputs(195));
    layer0_outputs(545) <= not((inputs(2)) and (inputs(188)));
    layer0_outputs(546) <= not((inputs(14)) or (inputs(75)));
    layer0_outputs(547) <= '0';
    layer0_outputs(548) <= (inputs(106)) xor (inputs(96));
    layer0_outputs(549) <= (inputs(39)) or (inputs(7));
    layer0_outputs(550) <= not(inputs(234)) or (inputs(154));
    layer0_outputs(551) <= (inputs(74)) and not (inputs(143));
    layer0_outputs(552) <= '0';
    layer0_outputs(553) <= not((inputs(114)) or (inputs(157)));
    layer0_outputs(554) <= not((inputs(43)) and (inputs(250)));
    layer0_outputs(555) <= not((inputs(168)) or (inputs(199)));
    layer0_outputs(556) <= inputs(104);
    layer0_outputs(557) <= (inputs(47)) xor (inputs(13));
    layer0_outputs(558) <= inputs(190);
    layer0_outputs(559) <= (inputs(74)) and not (inputs(166));
    layer0_outputs(560) <= not(inputs(101)) or (inputs(174));
    layer0_outputs(561) <= not((inputs(6)) or (inputs(7)));
    layer0_outputs(562) <= not(inputs(2));
    layer0_outputs(563) <= not((inputs(199)) or (inputs(251)));
    layer0_outputs(564) <= not(inputs(95));
    layer0_outputs(565) <= not(inputs(136));
    layer0_outputs(566) <= not((inputs(196)) or (inputs(116)));
    layer0_outputs(567) <= not(inputs(104));
    layer0_outputs(568) <= not(inputs(79)) or (inputs(25));
    layer0_outputs(569) <= (inputs(251)) or (inputs(22));
    layer0_outputs(570) <= inputs(104);
    layer0_outputs(571) <= not((inputs(55)) or (inputs(244)));
    layer0_outputs(572) <= '1';
    layer0_outputs(573) <= '1';
    layer0_outputs(574) <= (inputs(134)) or (inputs(85));
    layer0_outputs(575) <= (inputs(239)) and not (inputs(251));
    layer0_outputs(576) <= not(inputs(204));
    layer0_outputs(577) <= (inputs(165)) or (inputs(166));
    layer0_outputs(578) <= inputs(78);
    layer0_outputs(579) <= not(inputs(22)) or (inputs(183));
    layer0_outputs(580) <= not((inputs(227)) and (inputs(243)));
    layer0_outputs(581) <= not((inputs(12)) or (inputs(80)));
    layer0_outputs(582) <= inputs(157);
    layer0_outputs(583) <= not((inputs(149)) or (inputs(44)));
    layer0_outputs(584) <= (inputs(23)) and not (inputs(163));
    layer0_outputs(585) <= (inputs(82)) or (inputs(43));
    layer0_outputs(586) <= not(inputs(203)) or (inputs(14));
    layer0_outputs(587) <= inputs(178);
    layer0_outputs(588) <= inputs(150);
    layer0_outputs(589) <= not((inputs(225)) or (inputs(163)));
    layer0_outputs(590) <= not(inputs(65)) or (inputs(232));
    layer0_outputs(591) <= '1';
    layer0_outputs(592) <= not(inputs(198)) or (inputs(226));
    layer0_outputs(593) <= not((inputs(76)) or (inputs(94)));
    layer0_outputs(594) <= (inputs(2)) and (inputs(149));
    layer0_outputs(595) <= (inputs(133)) and not (inputs(95));
    layer0_outputs(596) <= '0';
    layer0_outputs(597) <= inputs(153);
    layer0_outputs(598) <= inputs(79);
    layer0_outputs(599) <= not(inputs(198)) or (inputs(34));
    layer0_outputs(600) <= not(inputs(111)) or (inputs(87));
    layer0_outputs(601) <= not((inputs(55)) xor (inputs(102)));
    layer0_outputs(602) <= (inputs(10)) and not (inputs(30));
    layer0_outputs(603) <= not(inputs(6));
    layer0_outputs(604) <= not(inputs(188)) or (inputs(89));
    layer0_outputs(605) <= (inputs(104)) and not (inputs(108));
    layer0_outputs(606) <= not((inputs(198)) or (inputs(227)));
    layer0_outputs(607) <= not(inputs(62));
    layer0_outputs(608) <= not(inputs(182));
    layer0_outputs(609) <= not((inputs(0)) or (inputs(138)));
    layer0_outputs(610) <= not((inputs(79)) xor (inputs(28)));
    layer0_outputs(611) <= '1';
    layer0_outputs(612) <= not(inputs(242)) or (inputs(114));
    layer0_outputs(613) <= not(inputs(139));
    layer0_outputs(614) <= (inputs(102)) or (inputs(68));
    layer0_outputs(615) <= (inputs(43)) and not (inputs(123));
    layer0_outputs(616) <= (inputs(178)) and not (inputs(191));
    layer0_outputs(617) <= inputs(217);
    layer0_outputs(618) <= (inputs(232)) and not (inputs(242));
    layer0_outputs(619) <= '1';
    layer0_outputs(620) <= '1';
    layer0_outputs(621) <= (inputs(187)) or (inputs(171));
    layer0_outputs(622) <= '1';
    layer0_outputs(623) <= not(inputs(51));
    layer0_outputs(624) <= inputs(133);
    layer0_outputs(625) <= not(inputs(183)) or (inputs(135));
    layer0_outputs(626) <= inputs(20);
    layer0_outputs(627) <= (inputs(142)) and (inputs(99));
    layer0_outputs(628) <= not(inputs(196)) or (inputs(22));
    layer0_outputs(629) <= (inputs(28)) or (inputs(44));
    layer0_outputs(630) <= not(inputs(232));
    layer0_outputs(631) <= (inputs(38)) or (inputs(5));
    layer0_outputs(632) <= (inputs(25)) and not (inputs(248));
    layer0_outputs(633) <= (inputs(88)) or (inputs(9));
    layer0_outputs(634) <= '0';
    layer0_outputs(635) <= not(inputs(168)) or (inputs(238));
    layer0_outputs(636) <= not(inputs(45));
    layer0_outputs(637) <= not(inputs(27));
    layer0_outputs(638) <= inputs(168);
    layer0_outputs(639) <= inputs(119);
    layer0_outputs(640) <= not((inputs(23)) xor (inputs(209)));
    layer0_outputs(641) <= '1';
    layer0_outputs(642) <= not((inputs(149)) or (inputs(161)));
    layer0_outputs(643) <= '1';
    layer0_outputs(644) <= not(inputs(228)) or (inputs(48));
    layer0_outputs(645) <= not((inputs(3)) and (inputs(200)));
    layer0_outputs(646) <= inputs(97);
    layer0_outputs(647) <= not(inputs(154)) or (inputs(127));
    layer0_outputs(648) <= inputs(69);
    layer0_outputs(649) <= not(inputs(163));
    layer0_outputs(650) <= not((inputs(252)) or (inputs(137)));
    layer0_outputs(651) <= inputs(72);
    layer0_outputs(652) <= (inputs(86)) or (inputs(61));
    layer0_outputs(653) <= not(inputs(128));
    layer0_outputs(654) <= (inputs(79)) and not (inputs(220));
    layer0_outputs(655) <= not(inputs(218));
    layer0_outputs(656) <= inputs(105);
    layer0_outputs(657) <= '0';
    layer0_outputs(658) <= not(inputs(58));
    layer0_outputs(659) <= (inputs(176)) and not (inputs(245));
    layer0_outputs(660) <= not((inputs(34)) and (inputs(225)));
    layer0_outputs(661) <= inputs(163);
    layer0_outputs(662) <= inputs(176);
    layer0_outputs(663) <= inputs(125);
    layer0_outputs(664) <= (inputs(187)) and (inputs(245));
    layer0_outputs(665) <= not(inputs(45));
    layer0_outputs(666) <= '0';
    layer0_outputs(667) <= (inputs(110)) or (inputs(247));
    layer0_outputs(668) <= inputs(114);
    layer0_outputs(669) <= (inputs(177)) and not (inputs(75));
    layer0_outputs(670) <= not((inputs(57)) or (inputs(163)));
    layer0_outputs(671) <= (inputs(175)) and not (inputs(240));
    layer0_outputs(672) <= (inputs(28)) and not (inputs(41));
    layer0_outputs(673) <= (inputs(138)) and (inputs(114));
    layer0_outputs(674) <= (inputs(160)) or (inputs(215));
    layer0_outputs(675) <= inputs(231);
    layer0_outputs(676) <= inputs(119);
    layer0_outputs(677) <= (inputs(108)) and not (inputs(243));
    layer0_outputs(678) <= (inputs(62)) or (inputs(60));
    layer0_outputs(679) <= not((inputs(176)) or (inputs(236)));
    layer0_outputs(680) <= (inputs(76)) and not (inputs(149));
    layer0_outputs(681) <= (inputs(117)) and not (inputs(134));
    layer0_outputs(682) <= (inputs(186)) and not (inputs(202));
    layer0_outputs(683) <= '0';
    layer0_outputs(684) <= inputs(112);
    layer0_outputs(685) <= not((inputs(67)) or (inputs(90)));
    layer0_outputs(686) <= (inputs(89)) and (inputs(124));
    layer0_outputs(687) <= '1';
    layer0_outputs(688) <= not((inputs(182)) xor (inputs(95)));
    layer0_outputs(689) <= inputs(24);
    layer0_outputs(690) <= (inputs(84)) or (inputs(67));
    layer0_outputs(691) <= not(inputs(133)) or (inputs(114));
    layer0_outputs(692) <= inputs(162);
    layer0_outputs(693) <= inputs(93);
    layer0_outputs(694) <= (inputs(78)) and not (inputs(4));
    layer0_outputs(695) <= not((inputs(252)) or (inputs(15)));
    layer0_outputs(696) <= not((inputs(205)) or (inputs(180)));
    layer0_outputs(697) <= not((inputs(118)) xor (inputs(129)));
    layer0_outputs(698) <= not(inputs(162)) or (inputs(9));
    layer0_outputs(699) <= inputs(61);
    layer0_outputs(700) <= (inputs(90)) or (inputs(19));
    layer0_outputs(701) <= (inputs(69)) or (inputs(164));
    layer0_outputs(702) <= inputs(37);
    layer0_outputs(703) <= inputs(77);
    layer0_outputs(704) <= not(inputs(253));
    layer0_outputs(705) <= not(inputs(92));
    layer0_outputs(706) <= inputs(13);
    layer0_outputs(707) <= inputs(247);
    layer0_outputs(708) <= (inputs(188)) and not (inputs(110));
    layer0_outputs(709) <= not((inputs(103)) and (inputs(207)));
    layer0_outputs(710) <= '1';
    layer0_outputs(711) <= '1';
    layer0_outputs(712) <= '0';
    layer0_outputs(713) <= inputs(110);
    layer0_outputs(714) <= not(inputs(145)) or (inputs(226));
    layer0_outputs(715) <= inputs(75);
    layer0_outputs(716) <= not(inputs(52));
    layer0_outputs(717) <= '0';
    layer0_outputs(718) <= '1';
    layer0_outputs(719) <= not(inputs(145)) or (inputs(47));
    layer0_outputs(720) <= (inputs(149)) or (inputs(17));
    layer0_outputs(721) <= not(inputs(31)) or (inputs(184));
    layer0_outputs(722) <= not(inputs(164)) or (inputs(179));
    layer0_outputs(723) <= (inputs(88)) and not (inputs(5));
    layer0_outputs(724) <= inputs(192);
    layer0_outputs(725) <= not((inputs(121)) or (inputs(30)));
    layer0_outputs(726) <= inputs(120);
    layer0_outputs(727) <= not((inputs(24)) xor (inputs(28)));
    layer0_outputs(728) <= not(inputs(30)) or (inputs(16));
    layer0_outputs(729) <= not(inputs(195));
    layer0_outputs(730) <= (inputs(84)) and not (inputs(197));
    layer0_outputs(731) <= (inputs(53)) and not (inputs(211));
    layer0_outputs(732) <= (inputs(238)) and not (inputs(82));
    layer0_outputs(733) <= not(inputs(193)) or (inputs(187));
    layer0_outputs(734) <= not((inputs(59)) and (inputs(160)));
    layer0_outputs(735) <= not(inputs(91));
    layer0_outputs(736) <= '1';
    layer0_outputs(737) <= not((inputs(233)) xor (inputs(56)));
    layer0_outputs(738) <= not(inputs(32));
    layer0_outputs(739) <= not(inputs(184)) or (inputs(47));
    layer0_outputs(740) <= inputs(248);
    layer0_outputs(741) <= not((inputs(199)) and (inputs(42)));
    layer0_outputs(742) <= not(inputs(30)) or (inputs(101));
    layer0_outputs(743) <= not((inputs(20)) or (inputs(42)));
    layer0_outputs(744) <= not(inputs(174)) or (inputs(150));
    layer0_outputs(745) <= not(inputs(42));
    layer0_outputs(746) <= not(inputs(193));
    layer0_outputs(747) <= '0';
    layer0_outputs(748) <= not((inputs(236)) xor (inputs(28)));
    layer0_outputs(749) <= '0';
    layer0_outputs(750) <= '0';
    layer0_outputs(751) <= not((inputs(67)) or (inputs(57)));
    layer0_outputs(752) <= not((inputs(12)) or (inputs(43)));
    layer0_outputs(753) <= '0';
    layer0_outputs(754) <= not(inputs(206)) or (inputs(185));
    layer0_outputs(755) <= '1';
    layer0_outputs(756) <= not(inputs(28)) or (inputs(43));
    layer0_outputs(757) <= not((inputs(78)) or (inputs(79)));
    layer0_outputs(758) <= inputs(170);
    layer0_outputs(759) <= (inputs(73)) and not (inputs(18));
    layer0_outputs(760) <= not(inputs(176));
    layer0_outputs(761) <= not((inputs(126)) or (inputs(22)));
    layer0_outputs(762) <= '1';
    layer0_outputs(763) <= '1';
    layer0_outputs(764) <= not(inputs(157));
    layer0_outputs(765) <= not(inputs(178));
    layer0_outputs(766) <= not((inputs(73)) or (inputs(128)));
    layer0_outputs(767) <= not((inputs(113)) or (inputs(95)));
    layer0_outputs(768) <= (inputs(83)) or (inputs(37));
    layer0_outputs(769) <= not(inputs(123));
    layer0_outputs(770) <= not(inputs(147)) or (inputs(69));
    layer0_outputs(771) <= not(inputs(178));
    layer0_outputs(772) <= '0';
    layer0_outputs(773) <= not((inputs(149)) or (inputs(154)));
    layer0_outputs(774) <= not((inputs(234)) or (inputs(103)));
    layer0_outputs(775) <= not(inputs(184));
    layer0_outputs(776) <= not(inputs(105)) or (inputs(196));
    layer0_outputs(777) <= (inputs(21)) and not (inputs(176));
    layer0_outputs(778) <= not(inputs(230));
    layer0_outputs(779) <= not((inputs(204)) or (inputs(40)));
    layer0_outputs(780) <= inputs(236);
    layer0_outputs(781) <= (inputs(173)) and not (inputs(121));
    layer0_outputs(782) <= not((inputs(8)) or (inputs(29)));
    layer0_outputs(783) <= (inputs(88)) or (inputs(102));
    layer0_outputs(784) <= not(inputs(33)) or (inputs(82));
    layer0_outputs(785) <= (inputs(199)) and not (inputs(162));
    layer0_outputs(786) <= (inputs(212)) and not (inputs(62));
    layer0_outputs(787) <= not(inputs(199)) or (inputs(133));
    layer0_outputs(788) <= (inputs(9)) or (inputs(192));
    layer0_outputs(789) <= (inputs(78)) or (inputs(203));
    layer0_outputs(790) <= not((inputs(32)) and (inputs(141)));
    layer0_outputs(791) <= not(inputs(236)) or (inputs(140));
    layer0_outputs(792) <= (inputs(234)) and not (inputs(243));
    layer0_outputs(793) <= not((inputs(146)) xor (inputs(65)));
    layer0_outputs(794) <= inputs(167);
    layer0_outputs(795) <= '0';
    layer0_outputs(796) <= (inputs(48)) and not (inputs(47));
    layer0_outputs(797) <= inputs(17);
    layer0_outputs(798) <= inputs(121);
    layer0_outputs(799) <= not(inputs(61)) or (inputs(239));
    layer0_outputs(800) <= inputs(91);
    layer0_outputs(801) <= not(inputs(8)) or (inputs(103));
    layer0_outputs(802) <= not(inputs(131)) or (inputs(61));
    layer0_outputs(803) <= not(inputs(209)) or (inputs(250));
    layer0_outputs(804) <= (inputs(100)) and not (inputs(18));
    layer0_outputs(805) <= inputs(232);
    layer0_outputs(806) <= inputs(122);
    layer0_outputs(807) <= inputs(26);
    layer0_outputs(808) <= not((inputs(63)) xor (inputs(191)));
    layer0_outputs(809) <= (inputs(20)) or (inputs(207));
    layer0_outputs(810) <= (inputs(249)) or (inputs(89));
    layer0_outputs(811) <= not((inputs(81)) or (inputs(171)));
    layer0_outputs(812) <= (inputs(223)) and (inputs(13));
    layer0_outputs(813) <= inputs(159);
    layer0_outputs(814) <= inputs(3);
    layer0_outputs(815) <= not(inputs(114));
    layer0_outputs(816) <= (inputs(193)) and not (inputs(116));
    layer0_outputs(817) <= '0';
    layer0_outputs(818) <= not((inputs(245)) or (inputs(77)));
    layer0_outputs(819) <= '1';
    layer0_outputs(820) <= not(inputs(103));
    layer0_outputs(821) <= not(inputs(59));
    layer0_outputs(822) <= not((inputs(35)) xor (inputs(107)));
    layer0_outputs(823) <= (inputs(190)) or (inputs(215));
    layer0_outputs(824) <= not((inputs(94)) or (inputs(203)));
    layer0_outputs(825) <= not(inputs(91)) or (inputs(209));
    layer0_outputs(826) <= (inputs(248)) and not (inputs(213));
    layer0_outputs(827) <= not((inputs(164)) or (inputs(127)));
    layer0_outputs(828) <= (inputs(93)) and (inputs(100));
    layer0_outputs(829) <= not((inputs(170)) or (inputs(165)));
    layer0_outputs(830) <= not(inputs(203));
    layer0_outputs(831) <= (inputs(119)) or (inputs(191));
    layer0_outputs(832) <= (inputs(137)) or (inputs(253));
    layer0_outputs(833) <= (inputs(245)) or (inputs(143));
    layer0_outputs(834) <= (inputs(151)) or (inputs(177));
    layer0_outputs(835) <= (inputs(79)) and not (inputs(162));
    layer0_outputs(836) <= inputs(197);
    layer0_outputs(837) <= (inputs(21)) and not (inputs(107));
    layer0_outputs(838) <= (inputs(157)) or (inputs(86));
    layer0_outputs(839) <= (inputs(117)) and not (inputs(207));
    layer0_outputs(840) <= (inputs(97)) or (inputs(164));
    layer0_outputs(841) <= not(inputs(61));
    layer0_outputs(842) <= not(inputs(98)) or (inputs(211));
    layer0_outputs(843) <= '0';
    layer0_outputs(844) <= (inputs(172)) or (inputs(229));
    layer0_outputs(845) <= not(inputs(145)) or (inputs(14));
    layer0_outputs(846) <= '0';
    layer0_outputs(847) <= inputs(102);
    layer0_outputs(848) <= (inputs(153)) or (inputs(238));
    layer0_outputs(849) <= not(inputs(132));
    layer0_outputs(850) <= not((inputs(131)) or (inputs(67)));
    layer0_outputs(851) <= (inputs(206)) and not (inputs(17));
    layer0_outputs(852) <= not(inputs(118));
    layer0_outputs(853) <= '0';
    layer0_outputs(854) <= inputs(199);
    layer0_outputs(855) <= not((inputs(233)) and (inputs(113)));
    layer0_outputs(856) <= inputs(135);
    layer0_outputs(857) <= inputs(96);
    layer0_outputs(858) <= not((inputs(65)) or (inputs(29)));
    layer0_outputs(859) <= not(inputs(74));
    layer0_outputs(860) <= '0';
    layer0_outputs(861) <= inputs(59);
    layer0_outputs(862) <= '0';
    layer0_outputs(863) <= not((inputs(121)) or (inputs(219)));
    layer0_outputs(864) <= not(inputs(72));
    layer0_outputs(865) <= not(inputs(71));
    layer0_outputs(866) <= (inputs(85)) and not (inputs(207));
    layer0_outputs(867) <= not(inputs(53));
    layer0_outputs(868) <= not((inputs(53)) xor (inputs(34)));
    layer0_outputs(869) <= not((inputs(191)) xor (inputs(47)));
    layer0_outputs(870) <= not(inputs(94));
    layer0_outputs(871) <= not((inputs(108)) and (inputs(103)));
    layer0_outputs(872) <= inputs(163);
    layer0_outputs(873) <= '0';
    layer0_outputs(874) <= not((inputs(179)) or (inputs(34)));
    layer0_outputs(875) <= not(inputs(197)) or (inputs(107));
    layer0_outputs(876) <= not((inputs(173)) or (inputs(176)));
    layer0_outputs(877) <= not(inputs(86));
    layer0_outputs(878) <= (inputs(6)) or (inputs(37));
    layer0_outputs(879) <= not((inputs(228)) or (inputs(211)));
    layer0_outputs(880) <= inputs(132);
    layer0_outputs(881) <= (inputs(195)) and not (inputs(154));
    layer0_outputs(882) <= (inputs(18)) or (inputs(83));
    layer0_outputs(883) <= '0';
    layer0_outputs(884) <= (inputs(96)) or (inputs(167));
    layer0_outputs(885) <= not(inputs(238));
    layer0_outputs(886) <= '0';
    layer0_outputs(887) <= (inputs(3)) xor (inputs(121));
    layer0_outputs(888) <= (inputs(212)) and not (inputs(153));
    layer0_outputs(889) <= not(inputs(168)) or (inputs(130));
    layer0_outputs(890) <= not((inputs(238)) or (inputs(21)));
    layer0_outputs(891) <= (inputs(108)) and not (inputs(151));
    layer0_outputs(892) <= not(inputs(17));
    layer0_outputs(893) <= not(inputs(145));
    layer0_outputs(894) <= (inputs(76)) and not (inputs(14));
    layer0_outputs(895) <= not(inputs(138)) or (inputs(204));
    layer0_outputs(896) <= not((inputs(0)) or (inputs(24)));
    layer0_outputs(897) <= not((inputs(113)) or (inputs(98)));
    layer0_outputs(898) <= (inputs(150)) and not (inputs(242));
    layer0_outputs(899) <= (inputs(104)) and not (inputs(181));
    layer0_outputs(900) <= inputs(178);
    layer0_outputs(901) <= (inputs(239)) or (inputs(2));
    layer0_outputs(902) <= not((inputs(226)) xor (inputs(62)));
    layer0_outputs(903) <= (inputs(59)) or (inputs(163));
    layer0_outputs(904) <= not((inputs(170)) or (inputs(115)));
    layer0_outputs(905) <= (inputs(122)) or (inputs(82));
    layer0_outputs(906) <= not(inputs(207));
    layer0_outputs(907) <= '0';
    layer0_outputs(908) <= '0';
    layer0_outputs(909) <= (inputs(84)) and not (inputs(19));
    layer0_outputs(910) <= not((inputs(161)) xor (inputs(34)));
    layer0_outputs(911) <= not(inputs(39));
    layer0_outputs(912) <= not(inputs(117)) or (inputs(208));
    layer0_outputs(913) <= not(inputs(184));
    layer0_outputs(914) <= (inputs(24)) xor (inputs(252));
    layer0_outputs(915) <= '0';
    layer0_outputs(916) <= (inputs(47)) and not (inputs(19));
    layer0_outputs(917) <= not((inputs(198)) or (inputs(161)));
    layer0_outputs(918) <= '1';
    layer0_outputs(919) <= not((inputs(140)) and (inputs(173)));
    layer0_outputs(920) <= not(inputs(172));
    layer0_outputs(921) <= inputs(76);
    layer0_outputs(922) <= '0';
    layer0_outputs(923) <= (inputs(196)) xor (inputs(177));
    layer0_outputs(924) <= inputs(39);
    layer0_outputs(925) <= not((inputs(38)) or (inputs(142)));
    layer0_outputs(926) <= not((inputs(69)) xor (inputs(97)));
    layer0_outputs(927) <= not(inputs(83)) or (inputs(113));
    layer0_outputs(928) <= (inputs(50)) and not (inputs(46));
    layer0_outputs(929) <= '0';
    layer0_outputs(930) <= not(inputs(127));
    layer0_outputs(931) <= (inputs(124)) or (inputs(137));
    layer0_outputs(932) <= '1';
    layer0_outputs(933) <= not(inputs(112)) or (inputs(176));
    layer0_outputs(934) <= (inputs(148)) or (inputs(63));
    layer0_outputs(935) <= not(inputs(43)) or (inputs(244));
    layer0_outputs(936) <= (inputs(176)) or (inputs(211));
    layer0_outputs(937) <= not(inputs(68)) or (inputs(153));
    layer0_outputs(938) <= not(inputs(139));
    layer0_outputs(939) <= inputs(244);
    layer0_outputs(940) <= (inputs(236)) or (inputs(85));
    layer0_outputs(941) <= (inputs(42)) or (inputs(88));
    layer0_outputs(942) <= not(inputs(171));
    layer0_outputs(943) <= not(inputs(69));
    layer0_outputs(944) <= not(inputs(22));
    layer0_outputs(945) <= not((inputs(101)) or (inputs(227)));
    layer0_outputs(946) <= '0';
    layer0_outputs(947) <= inputs(33);
    layer0_outputs(948) <= (inputs(161)) and not (inputs(173));
    layer0_outputs(949) <= not(inputs(207)) or (inputs(112));
    layer0_outputs(950) <= not(inputs(155));
    layer0_outputs(951) <= not(inputs(159));
    layer0_outputs(952) <= not(inputs(118)) or (inputs(9));
    layer0_outputs(953) <= (inputs(43)) and not (inputs(178));
    layer0_outputs(954) <= not(inputs(102)) or (inputs(7));
    layer0_outputs(955) <= inputs(0);
    layer0_outputs(956) <= (inputs(118)) and not (inputs(2));
    layer0_outputs(957) <= inputs(233);
    layer0_outputs(958) <= (inputs(169)) or (inputs(156));
    layer0_outputs(959) <= not((inputs(125)) or (inputs(35)));
    layer0_outputs(960) <= '1';
    layer0_outputs(961) <= not(inputs(219)) or (inputs(99));
    layer0_outputs(962) <= not(inputs(88));
    layer0_outputs(963) <= not((inputs(204)) and (inputs(0)));
    layer0_outputs(964) <= inputs(193);
    layer0_outputs(965) <= (inputs(168)) and not (inputs(40));
    layer0_outputs(966) <= not(inputs(4)) or (inputs(40));
    layer0_outputs(967) <= not((inputs(28)) xor (inputs(33)));
    layer0_outputs(968) <= '1';
    layer0_outputs(969) <= not(inputs(139)) or (inputs(234));
    layer0_outputs(970) <= (inputs(202)) and (inputs(247));
    layer0_outputs(971) <= inputs(169);
    layer0_outputs(972) <= not(inputs(2));
    layer0_outputs(973) <= not(inputs(226)) or (inputs(211));
    layer0_outputs(974) <= not(inputs(220));
    layer0_outputs(975) <= not(inputs(68)) or (inputs(46));
    layer0_outputs(976) <= not((inputs(156)) and (inputs(181)));
    layer0_outputs(977) <= not((inputs(209)) or (inputs(40)));
    layer0_outputs(978) <= (inputs(213)) or (inputs(59));
    layer0_outputs(979) <= not(inputs(245)) or (inputs(251));
    layer0_outputs(980) <= '1';
    layer0_outputs(981) <= inputs(109);
    layer0_outputs(982) <= (inputs(49)) and not (inputs(238));
    layer0_outputs(983) <= '1';
    layer0_outputs(984) <= (inputs(159)) and not (inputs(69));
    layer0_outputs(985) <= inputs(231);
    layer0_outputs(986) <= not(inputs(128));
    layer0_outputs(987) <= inputs(123);
    layer0_outputs(988) <= not((inputs(166)) xor (inputs(147)));
    layer0_outputs(989) <= not((inputs(99)) or (inputs(204)));
    layer0_outputs(990) <= inputs(101);
    layer0_outputs(991) <= '1';
    layer0_outputs(992) <= inputs(177);
    layer0_outputs(993) <= not(inputs(77));
    layer0_outputs(994) <= (inputs(116)) xor (inputs(86));
    layer0_outputs(995) <= (inputs(66)) or (inputs(84));
    layer0_outputs(996) <= inputs(195);
    layer0_outputs(997) <= not(inputs(93));
    layer0_outputs(998) <= not(inputs(37)) or (inputs(178));
    layer0_outputs(999) <= not(inputs(161)) or (inputs(64));
    layer0_outputs(1000) <= inputs(136);
    layer0_outputs(1001) <= (inputs(157)) or (inputs(187));
    layer0_outputs(1002) <= inputs(252);
    layer0_outputs(1003) <= not((inputs(171)) or (inputs(85)));
    layer0_outputs(1004) <= not(inputs(60)) or (inputs(240));
    layer0_outputs(1005) <= (inputs(170)) and not (inputs(113));
    layer0_outputs(1006) <= not(inputs(244)) or (inputs(1));
    layer0_outputs(1007) <= (inputs(125)) and not (inputs(179));
    layer0_outputs(1008) <= inputs(81);
    layer0_outputs(1009) <= not((inputs(104)) and (inputs(224)));
    layer0_outputs(1010) <= inputs(54);
    layer0_outputs(1011) <= (inputs(117)) and not (inputs(34));
    layer0_outputs(1012) <= (inputs(105)) and (inputs(221));
    layer0_outputs(1013) <= not(inputs(179));
    layer0_outputs(1014) <= not(inputs(221));
    layer0_outputs(1015) <= '0';
    layer0_outputs(1016) <= not((inputs(16)) or (inputs(172)));
    layer0_outputs(1017) <= inputs(38);
    layer0_outputs(1018) <= inputs(67);
    layer0_outputs(1019) <= inputs(223);
    layer0_outputs(1020) <= (inputs(91)) and not (inputs(117));
    layer0_outputs(1021) <= not((inputs(229)) or (inputs(72)));
    layer0_outputs(1022) <= not(inputs(52)) or (inputs(214));
    layer0_outputs(1023) <= not(inputs(93));
    layer0_outputs(1024) <= not((inputs(54)) and (inputs(17)));
    layer0_outputs(1025) <= (inputs(109)) and not (inputs(230));
    layer0_outputs(1026) <= (inputs(207)) xor (inputs(31));
    layer0_outputs(1027) <= not(inputs(188));
    layer0_outputs(1028) <= (inputs(13)) and (inputs(16));
    layer0_outputs(1029) <= (inputs(144)) xor (inputs(99));
    layer0_outputs(1030) <= not(inputs(83)) or (inputs(29));
    layer0_outputs(1031) <= inputs(126);
    layer0_outputs(1032) <= inputs(251);
    layer0_outputs(1033) <= not(inputs(116));
    layer0_outputs(1034) <= not((inputs(66)) or (inputs(19)));
    layer0_outputs(1035) <= not((inputs(47)) or (inputs(22)));
    layer0_outputs(1036) <= '1';
    layer0_outputs(1037) <= inputs(21);
    layer0_outputs(1038) <= not(inputs(22)) or (inputs(90));
    layer0_outputs(1039) <= not((inputs(62)) or (inputs(245)));
    layer0_outputs(1040) <= (inputs(120)) and not (inputs(186));
    layer0_outputs(1041) <= (inputs(105)) and not (inputs(99));
    layer0_outputs(1042) <= inputs(247);
    layer0_outputs(1043) <= not((inputs(140)) or (inputs(218)));
    layer0_outputs(1044) <= not(inputs(91));
    layer0_outputs(1045) <= not(inputs(23)) or (inputs(143));
    layer0_outputs(1046) <= (inputs(100)) and not (inputs(136));
    layer0_outputs(1047) <= not((inputs(234)) or (inputs(216)));
    layer0_outputs(1048) <= not(inputs(44));
    layer0_outputs(1049) <= '1';
    layer0_outputs(1050) <= not((inputs(2)) or (inputs(207)));
    layer0_outputs(1051) <= not(inputs(127)) or (inputs(20));
    layer0_outputs(1052) <= (inputs(227)) or (inputs(97));
    layer0_outputs(1053) <= inputs(230);
    layer0_outputs(1054) <= inputs(54);
    layer0_outputs(1055) <= not((inputs(176)) and (inputs(124)));
    layer0_outputs(1056) <= inputs(172);
    layer0_outputs(1057) <= (inputs(176)) xor (inputs(232));
    layer0_outputs(1058) <= (inputs(10)) and not (inputs(72));
    layer0_outputs(1059) <= not((inputs(9)) or (inputs(230)));
    layer0_outputs(1060) <= not(inputs(180));
    layer0_outputs(1061) <= not((inputs(16)) xor (inputs(208)));
    layer0_outputs(1062) <= (inputs(58)) xor (inputs(130));
    layer0_outputs(1063) <= inputs(104);
    layer0_outputs(1064) <= (inputs(214)) and (inputs(48));
    layer0_outputs(1065) <= (inputs(30)) and (inputs(3));
    layer0_outputs(1066) <= inputs(113);
    layer0_outputs(1067) <= not(inputs(146));
    layer0_outputs(1068) <= not((inputs(28)) or (inputs(201)));
    layer0_outputs(1069) <= not(inputs(39));
    layer0_outputs(1070) <= not(inputs(211));
    layer0_outputs(1071) <= (inputs(226)) xor (inputs(73));
    layer0_outputs(1072) <= (inputs(33)) and (inputs(14));
    layer0_outputs(1073) <= not((inputs(181)) xor (inputs(144)));
    layer0_outputs(1074) <= not(inputs(78));
    layer0_outputs(1075) <= not(inputs(34)) or (inputs(221));
    layer0_outputs(1076) <= '1';
    layer0_outputs(1077) <= inputs(206);
    layer0_outputs(1078) <= not(inputs(226)) or (inputs(31));
    layer0_outputs(1079) <= not((inputs(153)) xor (inputs(146)));
    layer0_outputs(1080) <= (inputs(122)) and not (inputs(221));
    layer0_outputs(1081) <= not((inputs(32)) or (inputs(65)));
    layer0_outputs(1082) <= not((inputs(208)) xor (inputs(51)));
    layer0_outputs(1083) <= (inputs(185)) and not (inputs(141));
    layer0_outputs(1084) <= not(inputs(21));
    layer0_outputs(1085) <= not((inputs(80)) and (inputs(77)));
    layer0_outputs(1086) <= not((inputs(85)) and (inputs(35)));
    layer0_outputs(1087) <= not(inputs(52));
    layer0_outputs(1088) <= not(inputs(76));
    layer0_outputs(1089) <= (inputs(198)) and not (inputs(106));
    layer0_outputs(1090) <= not(inputs(231));
    layer0_outputs(1091) <= (inputs(56)) or (inputs(147));
    layer0_outputs(1092) <= not(inputs(14));
    layer0_outputs(1093) <= not(inputs(187));
    layer0_outputs(1094) <= inputs(162);
    layer0_outputs(1095) <= inputs(5);
    layer0_outputs(1096) <= inputs(206);
    layer0_outputs(1097) <= not((inputs(205)) and (inputs(249)));
    layer0_outputs(1098) <= not((inputs(191)) or (inputs(233)));
    layer0_outputs(1099) <= inputs(104);
    layer0_outputs(1100) <= not(inputs(190)) or (inputs(159));
    layer0_outputs(1101) <= inputs(166);
    layer0_outputs(1102) <= (inputs(37)) and not (inputs(181));
    layer0_outputs(1103) <= (inputs(85)) or (inputs(38));
    layer0_outputs(1104) <= inputs(193);
    layer0_outputs(1105) <= '0';
    layer0_outputs(1106) <= not(inputs(105));
    layer0_outputs(1107) <= (inputs(160)) or (inputs(114));
    layer0_outputs(1108) <= not(inputs(208));
    layer0_outputs(1109) <= not(inputs(7)) or (inputs(16));
    layer0_outputs(1110) <= not(inputs(147)) or (inputs(5));
    layer0_outputs(1111) <= not((inputs(85)) xor (inputs(19)));
    layer0_outputs(1112) <= (inputs(190)) and (inputs(201));
    layer0_outputs(1113) <= not(inputs(218));
    layer0_outputs(1114) <= inputs(249);
    layer0_outputs(1115) <= (inputs(13)) or (inputs(29));
    layer0_outputs(1116) <= not(inputs(0));
    layer0_outputs(1117) <= not((inputs(199)) or (inputs(253)));
    layer0_outputs(1118) <= not((inputs(138)) or (inputs(235)));
    layer0_outputs(1119) <= not(inputs(218)) or (inputs(227));
    layer0_outputs(1120) <= (inputs(127)) or (inputs(88));
    layer0_outputs(1121) <= not(inputs(251)) or (inputs(209));
    layer0_outputs(1122) <= (inputs(255)) and (inputs(173));
    layer0_outputs(1123) <= (inputs(122)) and not (inputs(204));
    layer0_outputs(1124) <= (inputs(13)) xor (inputs(120));
    layer0_outputs(1125) <= (inputs(217)) or (inputs(134));
    layer0_outputs(1126) <= inputs(39);
    layer0_outputs(1127) <= not(inputs(86)) or (inputs(156));
    layer0_outputs(1128) <= (inputs(130)) or (inputs(183));
    layer0_outputs(1129) <= not(inputs(75)) or (inputs(158));
    layer0_outputs(1130) <= '0';
    layer0_outputs(1131) <= (inputs(86)) and not (inputs(49));
    layer0_outputs(1132) <= not(inputs(134)) or (inputs(66));
    layer0_outputs(1133) <= (inputs(130)) and not (inputs(33));
    layer0_outputs(1134) <= not((inputs(61)) and (inputs(18)));
    layer0_outputs(1135) <= (inputs(29)) and (inputs(11));
    layer0_outputs(1136) <= (inputs(92)) and not (inputs(48));
    layer0_outputs(1137) <= (inputs(123)) and not (inputs(73));
    layer0_outputs(1138) <= not(inputs(182));
    layer0_outputs(1139) <= (inputs(150)) and not (inputs(184));
    layer0_outputs(1140) <= '0';
    layer0_outputs(1141) <= not(inputs(91));
    layer0_outputs(1142) <= inputs(130);
    layer0_outputs(1143) <= not(inputs(45)) or (inputs(202));
    layer0_outputs(1144) <= not(inputs(220));
    layer0_outputs(1145) <= not((inputs(210)) and (inputs(200)));
    layer0_outputs(1146) <= '0';
    layer0_outputs(1147) <= '0';
    layer0_outputs(1148) <= not((inputs(204)) and (inputs(141)));
    layer0_outputs(1149) <= not(inputs(234));
    layer0_outputs(1150) <= inputs(85);
    layer0_outputs(1151) <= (inputs(16)) and not (inputs(223));
    layer0_outputs(1152) <= not((inputs(183)) xor (inputs(221)));
    layer0_outputs(1153) <= not((inputs(186)) or (inputs(159)));
    layer0_outputs(1154) <= not((inputs(209)) xor (inputs(206)));
    layer0_outputs(1155) <= (inputs(93)) and not (inputs(48));
    layer0_outputs(1156) <= not((inputs(1)) or (inputs(23)));
    layer0_outputs(1157) <= inputs(177);
    layer0_outputs(1158) <= not((inputs(230)) or (inputs(208)));
    layer0_outputs(1159) <= not((inputs(105)) and (inputs(232)));
    layer0_outputs(1160) <= not(inputs(105));
    layer0_outputs(1161) <= not(inputs(231));
    layer0_outputs(1162) <= not(inputs(241)) or (inputs(54));
    layer0_outputs(1163) <= not(inputs(175));
    layer0_outputs(1164) <= not(inputs(90));
    layer0_outputs(1165) <= not(inputs(162));
    layer0_outputs(1166) <= not((inputs(109)) and (inputs(65)));
    layer0_outputs(1167) <= not(inputs(223));
    layer0_outputs(1168) <= (inputs(92)) or (inputs(51));
    layer0_outputs(1169) <= (inputs(110)) and not (inputs(252));
    layer0_outputs(1170) <= not((inputs(74)) and (inputs(19)));
    layer0_outputs(1171) <= (inputs(180)) and not (inputs(81));
    layer0_outputs(1172) <= (inputs(198)) xor (inputs(181));
    layer0_outputs(1173) <= not(inputs(150));
    layer0_outputs(1174) <= not(inputs(53)) or (inputs(236));
    layer0_outputs(1175) <= not((inputs(1)) or (inputs(111)));
    layer0_outputs(1176) <= not(inputs(77));
    layer0_outputs(1177) <= (inputs(253)) or (inputs(10));
    layer0_outputs(1178) <= inputs(182);
    layer0_outputs(1179) <= not(inputs(93)) or (inputs(125));
    layer0_outputs(1180) <= not(inputs(250)) or (inputs(38));
    layer0_outputs(1181) <= (inputs(84)) xor (inputs(36));
    layer0_outputs(1182) <= not(inputs(165));
    layer0_outputs(1183) <= (inputs(109)) or (inputs(153));
    layer0_outputs(1184) <= not(inputs(132));
    layer0_outputs(1185) <= not((inputs(62)) or (inputs(4)));
    layer0_outputs(1186) <= not(inputs(135));
    layer0_outputs(1187) <= '1';
    layer0_outputs(1188) <= not(inputs(130));
    layer0_outputs(1189) <= (inputs(230)) and (inputs(130));
    layer0_outputs(1190) <= '0';
    layer0_outputs(1191) <= (inputs(44)) and not (inputs(142));
    layer0_outputs(1192) <= not(inputs(135)) or (inputs(96));
    layer0_outputs(1193) <= inputs(121);
    layer0_outputs(1194) <= not(inputs(246));
    layer0_outputs(1195) <= not(inputs(209));
    layer0_outputs(1196) <= inputs(195);
    layer0_outputs(1197) <= inputs(156);
    layer0_outputs(1198) <= not((inputs(117)) and (inputs(40)));
    layer0_outputs(1199) <= '1';
    layer0_outputs(1200) <= inputs(26);
    layer0_outputs(1201) <= not(inputs(76)) or (inputs(240));
    layer0_outputs(1202) <= (inputs(102)) and not (inputs(33));
    layer0_outputs(1203) <= not((inputs(213)) or (inputs(193)));
    layer0_outputs(1204) <= not((inputs(166)) xor (inputs(148)));
    layer0_outputs(1205) <= not(inputs(60)) or (inputs(126));
    layer0_outputs(1206) <= (inputs(45)) xor (inputs(11));
    layer0_outputs(1207) <= not(inputs(48));
    layer0_outputs(1208) <= '0';
    layer0_outputs(1209) <= not((inputs(235)) xor (inputs(210)));
    layer0_outputs(1210) <= (inputs(162)) and not (inputs(94));
    layer0_outputs(1211) <= not(inputs(111));
    layer0_outputs(1212) <= not(inputs(121));
    layer0_outputs(1213) <= (inputs(77)) or (inputs(234));
    layer0_outputs(1214) <= not(inputs(71));
    layer0_outputs(1215) <= inputs(103);
    layer0_outputs(1216) <= inputs(26);
    layer0_outputs(1217) <= (inputs(96)) or (inputs(171));
    layer0_outputs(1218) <= '0';
    layer0_outputs(1219) <= not(inputs(25));
    layer0_outputs(1220) <= (inputs(204)) or (inputs(223));
    layer0_outputs(1221) <= not((inputs(192)) or (inputs(191)));
    layer0_outputs(1222) <= not(inputs(133)) or (inputs(180));
    layer0_outputs(1223) <= not(inputs(150)) or (inputs(2));
    layer0_outputs(1224) <= not(inputs(179));
    layer0_outputs(1225) <= not(inputs(157)) or (inputs(157));
    layer0_outputs(1226) <= not((inputs(193)) or (inputs(218)));
    layer0_outputs(1227) <= not(inputs(213));
    layer0_outputs(1228) <= '0';
    layer0_outputs(1229) <= not((inputs(46)) xor (inputs(20)));
    layer0_outputs(1230) <= not(inputs(213));
    layer0_outputs(1231) <= (inputs(73)) or (inputs(237));
    layer0_outputs(1232) <= not((inputs(203)) and (inputs(118)));
    layer0_outputs(1233) <= inputs(9);
    layer0_outputs(1234) <= '0';
    layer0_outputs(1235) <= inputs(76);
    layer0_outputs(1236) <= (inputs(53)) or (inputs(16));
    layer0_outputs(1237) <= not(inputs(105)) or (inputs(0));
    layer0_outputs(1238) <= not(inputs(22)) or (inputs(112));
    layer0_outputs(1239) <= not((inputs(144)) and (inputs(205)));
    layer0_outputs(1240) <= (inputs(70)) and not (inputs(190));
    layer0_outputs(1241) <= (inputs(14)) xor (inputs(196));
    layer0_outputs(1242) <= inputs(72);
    layer0_outputs(1243) <= not(inputs(232));
    layer0_outputs(1244) <= (inputs(143)) and not (inputs(9));
    layer0_outputs(1245) <= not((inputs(76)) or (inputs(77)));
    layer0_outputs(1246) <= '1';
    layer0_outputs(1247) <= not(inputs(165)) or (inputs(206));
    layer0_outputs(1248) <= '1';
    layer0_outputs(1249) <= not((inputs(51)) or (inputs(65)));
    layer0_outputs(1250) <= not((inputs(184)) or (inputs(255)));
    layer0_outputs(1251) <= inputs(2);
    layer0_outputs(1252) <= (inputs(187)) and not (inputs(18));
    layer0_outputs(1253) <= not(inputs(90)) or (inputs(128));
    layer0_outputs(1254) <= not(inputs(25));
    layer0_outputs(1255) <= '0';
    layer0_outputs(1256) <= not((inputs(191)) or (inputs(229)));
    layer0_outputs(1257) <= not(inputs(36)) or (inputs(196));
    layer0_outputs(1258) <= not(inputs(213));
    layer0_outputs(1259) <= not(inputs(100));
    layer0_outputs(1260) <= not(inputs(6)) or (inputs(101));
    layer0_outputs(1261) <= not(inputs(230));
    layer0_outputs(1262) <= (inputs(241)) and (inputs(206));
    layer0_outputs(1263) <= not(inputs(168)) or (inputs(92));
    layer0_outputs(1264) <= (inputs(115)) and (inputs(178));
    layer0_outputs(1265) <= not(inputs(1));
    layer0_outputs(1266) <= not((inputs(115)) or (inputs(255)));
    layer0_outputs(1267) <= inputs(37);
    layer0_outputs(1268) <= not(inputs(220)) or (inputs(87));
    layer0_outputs(1269) <= not(inputs(119));
    layer0_outputs(1270) <= (inputs(69)) or (inputs(129));
    layer0_outputs(1271) <= (inputs(155)) or (inputs(96));
    layer0_outputs(1272) <= (inputs(93)) or (inputs(163));
    layer0_outputs(1273) <= (inputs(193)) xor (inputs(84));
    layer0_outputs(1274) <= not(inputs(139)) or (inputs(66));
    layer0_outputs(1275) <= not(inputs(7)) or (inputs(130));
    layer0_outputs(1276) <= (inputs(83)) or (inputs(21));
    layer0_outputs(1277) <= not((inputs(38)) xor (inputs(146)));
    layer0_outputs(1278) <= not((inputs(185)) xor (inputs(44)));
    layer0_outputs(1279) <= '1';
    layer0_outputs(1280) <= not((inputs(31)) or (inputs(138)));
    layer0_outputs(1281) <= not(inputs(159));
    layer0_outputs(1282) <= not(inputs(130));
    layer0_outputs(1283) <= not(inputs(155)) or (inputs(204));
    layer0_outputs(1284) <= not(inputs(194)) or (inputs(10));
    layer0_outputs(1285) <= (inputs(195)) and not (inputs(44));
    layer0_outputs(1286) <= not(inputs(200)) or (inputs(110));
    layer0_outputs(1287) <= (inputs(127)) and not (inputs(251));
    layer0_outputs(1288) <= not((inputs(133)) or (inputs(237)));
    layer0_outputs(1289) <= inputs(224);
    layer0_outputs(1290) <= not((inputs(250)) or (inputs(244)));
    layer0_outputs(1291) <= not(inputs(90));
    layer0_outputs(1292) <= (inputs(3)) and not (inputs(77));
    layer0_outputs(1293) <= (inputs(195)) and (inputs(192));
    layer0_outputs(1294) <= not(inputs(158));
    layer0_outputs(1295) <= '1';
    layer0_outputs(1296) <= (inputs(151)) and not (inputs(46));
    layer0_outputs(1297) <= (inputs(226)) xor (inputs(205));
    layer0_outputs(1298) <= not(inputs(34));
    layer0_outputs(1299) <= (inputs(86)) and not (inputs(20));
    layer0_outputs(1300) <= not((inputs(255)) and (inputs(240)));
    layer0_outputs(1301) <= inputs(230);
    layer0_outputs(1302) <= (inputs(2)) or (inputs(121));
    layer0_outputs(1303) <= not(inputs(124)) or (inputs(167));
    layer0_outputs(1304) <= not(inputs(91));
    layer0_outputs(1305) <= not(inputs(157)) or (inputs(82));
    layer0_outputs(1306) <= (inputs(129)) and not (inputs(0));
    layer0_outputs(1307) <= (inputs(253)) or (inputs(44));
    layer0_outputs(1308) <= not(inputs(89)) or (inputs(27));
    layer0_outputs(1309) <= (inputs(227)) and not (inputs(126));
    layer0_outputs(1310) <= (inputs(176)) xor (inputs(96));
    layer0_outputs(1311) <= (inputs(166)) or (inputs(85));
    layer0_outputs(1312) <= '1';
    layer0_outputs(1313) <= '0';
    layer0_outputs(1314) <= not((inputs(215)) and (inputs(37)));
    layer0_outputs(1315) <= not((inputs(141)) and (inputs(191)));
    layer0_outputs(1316) <= (inputs(134)) and not (inputs(157));
    layer0_outputs(1317) <= '0';
    layer0_outputs(1318) <= inputs(26);
    layer0_outputs(1319) <= not((inputs(253)) or (inputs(222)));
    layer0_outputs(1320) <= not(inputs(1));
    layer0_outputs(1321) <= (inputs(253)) and not (inputs(95));
    layer0_outputs(1322) <= not(inputs(198));
    layer0_outputs(1323) <= not(inputs(224));
    layer0_outputs(1324) <= (inputs(126)) and not (inputs(92));
    layer0_outputs(1325) <= not(inputs(199)) or (inputs(88));
    layer0_outputs(1326) <= (inputs(25)) and not (inputs(250));
    layer0_outputs(1327) <= '1';
    layer0_outputs(1328) <= inputs(126);
    layer0_outputs(1329) <= '1';
    layer0_outputs(1330) <= (inputs(15)) or (inputs(177));
    layer0_outputs(1331) <= not((inputs(155)) or (inputs(190)));
    layer0_outputs(1332) <= inputs(234);
    layer0_outputs(1333) <= (inputs(84)) or (inputs(79));
    layer0_outputs(1334) <= not((inputs(75)) and (inputs(25)));
    layer0_outputs(1335) <= inputs(197);
    layer0_outputs(1336) <= inputs(2);
    layer0_outputs(1337) <= not(inputs(57)) or (inputs(219));
    layer0_outputs(1338) <= not(inputs(213)) or (inputs(45));
    layer0_outputs(1339) <= not((inputs(220)) xor (inputs(47)));
    layer0_outputs(1340) <= not(inputs(52)) or (inputs(103));
    layer0_outputs(1341) <= (inputs(131)) xor (inputs(144));
    layer0_outputs(1342) <= not((inputs(77)) or (inputs(5)));
    layer0_outputs(1343) <= not((inputs(109)) or (inputs(133)));
    layer0_outputs(1344) <= not(inputs(103));
    layer0_outputs(1345) <= not(inputs(145));
    layer0_outputs(1346) <= not(inputs(200)) or (inputs(86));
    layer0_outputs(1347) <= not((inputs(191)) or (inputs(215)));
    layer0_outputs(1348) <= '0';
    layer0_outputs(1349) <= (inputs(87)) xor (inputs(116));
    layer0_outputs(1350) <= (inputs(147)) and not (inputs(26));
    layer0_outputs(1351) <= '0';
    layer0_outputs(1352) <= not(inputs(109));
    layer0_outputs(1353) <= not((inputs(121)) or (inputs(35)));
    layer0_outputs(1354) <= (inputs(59)) and not (inputs(231));
    layer0_outputs(1355) <= (inputs(172)) or (inputs(187));
    layer0_outputs(1356) <= not((inputs(74)) and (inputs(128)));
    layer0_outputs(1357) <= (inputs(235)) or (inputs(230));
    layer0_outputs(1358) <= inputs(56);
    layer0_outputs(1359) <= (inputs(78)) and not (inputs(254));
    layer0_outputs(1360) <= inputs(159);
    layer0_outputs(1361) <= '1';
    layer0_outputs(1362) <= inputs(49);
    layer0_outputs(1363) <= not(inputs(222));
    layer0_outputs(1364) <= '0';
    layer0_outputs(1365) <= not(inputs(73));
    layer0_outputs(1366) <= not(inputs(233));
    layer0_outputs(1367) <= not((inputs(208)) and (inputs(66)));
    layer0_outputs(1368) <= (inputs(214)) and (inputs(202));
    layer0_outputs(1369) <= not(inputs(218)) or (inputs(154));
    layer0_outputs(1370) <= not((inputs(226)) or (inputs(25)));
    layer0_outputs(1371) <= not(inputs(114));
    layer0_outputs(1372) <= inputs(212);
    layer0_outputs(1373) <= inputs(49);
    layer0_outputs(1374) <= (inputs(229)) or (inputs(175));
    layer0_outputs(1375) <= not(inputs(173)) or (inputs(156));
    layer0_outputs(1376) <= (inputs(54)) xor (inputs(7));
    layer0_outputs(1377) <= inputs(113);
    layer0_outputs(1378) <= not(inputs(123));
    layer0_outputs(1379) <= not(inputs(48));
    layer0_outputs(1380) <= '0';
    layer0_outputs(1381) <= (inputs(62)) or (inputs(151));
    layer0_outputs(1382) <= (inputs(106)) and not (inputs(57));
    layer0_outputs(1383) <= (inputs(45)) and (inputs(47));
    layer0_outputs(1384) <= not((inputs(151)) and (inputs(184)));
    layer0_outputs(1385) <= not(inputs(210));
    layer0_outputs(1386) <= (inputs(182)) and not (inputs(228));
    layer0_outputs(1387) <= not((inputs(250)) xor (inputs(19)));
    layer0_outputs(1388) <= '0';
    layer0_outputs(1389) <= inputs(253);
    layer0_outputs(1390) <= not((inputs(221)) xor (inputs(157)));
    layer0_outputs(1391) <= (inputs(251)) and not (inputs(49));
    layer0_outputs(1392) <= not(inputs(165)) or (inputs(63));
    layer0_outputs(1393) <= not(inputs(32)) or (inputs(50));
    layer0_outputs(1394) <= inputs(13);
    layer0_outputs(1395) <= inputs(40);
    layer0_outputs(1396) <= (inputs(85)) and not (inputs(18));
    layer0_outputs(1397) <= (inputs(53)) and not (inputs(132));
    layer0_outputs(1398) <= not(inputs(97)) or (inputs(147));
    layer0_outputs(1399) <= '0';
    layer0_outputs(1400) <= (inputs(78)) or (inputs(91));
    layer0_outputs(1401) <= (inputs(121)) or (inputs(83));
    layer0_outputs(1402) <= not(inputs(162));
    layer0_outputs(1403) <= inputs(25);
    layer0_outputs(1404) <= not(inputs(59)) or (inputs(113));
    layer0_outputs(1405) <= not((inputs(13)) or (inputs(116)));
    layer0_outputs(1406) <= not(inputs(109)) or (inputs(140));
    layer0_outputs(1407) <= (inputs(205)) xor (inputs(13));
    layer0_outputs(1408) <= not((inputs(241)) xor (inputs(188)));
    layer0_outputs(1409) <= '0';
    layer0_outputs(1410) <= inputs(66);
    layer0_outputs(1411) <= not((inputs(184)) or (inputs(129)));
    layer0_outputs(1412) <= not(inputs(127)) or (inputs(240));
    layer0_outputs(1413) <= not(inputs(239)) or (inputs(81));
    layer0_outputs(1414) <= not(inputs(37));
    layer0_outputs(1415) <= (inputs(253)) and not (inputs(30));
    layer0_outputs(1416) <= (inputs(66)) and not (inputs(12));
    layer0_outputs(1417) <= not((inputs(67)) or (inputs(161)));
    layer0_outputs(1418) <= (inputs(8)) and not (inputs(226));
    layer0_outputs(1419) <= (inputs(225)) and not (inputs(125));
    layer0_outputs(1420) <= not(inputs(63));
    layer0_outputs(1421) <= not((inputs(189)) or (inputs(98)));
    layer0_outputs(1422) <= not((inputs(128)) or (inputs(97)));
    layer0_outputs(1423) <= not(inputs(118));
    layer0_outputs(1424) <= (inputs(26)) and not (inputs(188));
    layer0_outputs(1425) <= not(inputs(86));
    layer0_outputs(1426) <= '0';
    layer0_outputs(1427) <= not(inputs(29)) or (inputs(162));
    layer0_outputs(1428) <= (inputs(183)) and not (inputs(52));
    layer0_outputs(1429) <= not((inputs(242)) xor (inputs(219)));
    layer0_outputs(1430) <= not((inputs(129)) or (inputs(149)));
    layer0_outputs(1431) <= not(inputs(114));
    layer0_outputs(1432) <= inputs(70);
    layer0_outputs(1433) <= (inputs(36)) or (inputs(241));
    layer0_outputs(1434) <= not((inputs(83)) or (inputs(123)));
    layer0_outputs(1435) <= inputs(100);
    layer0_outputs(1436) <= not((inputs(214)) and (inputs(101)));
    layer0_outputs(1437) <= not((inputs(242)) xor (inputs(79)));
    layer0_outputs(1438) <= (inputs(223)) xor (inputs(94));
    layer0_outputs(1439) <= not(inputs(132)) or (inputs(236));
    layer0_outputs(1440) <= not((inputs(91)) or (inputs(185)));
    layer0_outputs(1441) <= not(inputs(248));
    layer0_outputs(1442) <= (inputs(103)) and (inputs(81));
    layer0_outputs(1443) <= not(inputs(127));
    layer0_outputs(1444) <= (inputs(190)) or (inputs(119));
    layer0_outputs(1445) <= inputs(128);
    layer0_outputs(1446) <= (inputs(201)) and (inputs(65));
    layer0_outputs(1447) <= not(inputs(220));
    layer0_outputs(1448) <= not((inputs(181)) xor (inputs(105)));
    layer0_outputs(1449) <= not(inputs(33));
    layer0_outputs(1450) <= inputs(14);
    layer0_outputs(1451) <= (inputs(94)) and not (inputs(251));
    layer0_outputs(1452) <= not((inputs(50)) or (inputs(56)));
    layer0_outputs(1453) <= not(inputs(62)) or (inputs(119));
    layer0_outputs(1454) <= '1';
    layer0_outputs(1455) <= inputs(51);
    layer0_outputs(1456) <= (inputs(108)) and (inputs(19));
    layer0_outputs(1457) <= (inputs(20)) or (inputs(174));
    layer0_outputs(1458) <= inputs(168);
    layer0_outputs(1459) <= (inputs(66)) or (inputs(32));
    layer0_outputs(1460) <= not((inputs(50)) and (inputs(216)));
    layer0_outputs(1461) <= '0';
    layer0_outputs(1462) <= not(inputs(2));
    layer0_outputs(1463) <= not(inputs(91));
    layer0_outputs(1464) <= (inputs(203)) and not (inputs(239));
    layer0_outputs(1465) <= (inputs(248)) and not (inputs(29));
    layer0_outputs(1466) <= not(inputs(69)) or (inputs(17));
    layer0_outputs(1467) <= '1';
    layer0_outputs(1468) <= not((inputs(214)) or (inputs(37)));
    layer0_outputs(1469) <= not((inputs(233)) xor (inputs(187)));
    layer0_outputs(1470) <= inputs(24);
    layer0_outputs(1471) <= not((inputs(40)) or (inputs(156)));
    layer0_outputs(1472) <= '0';
    layer0_outputs(1473) <= inputs(226);
    layer0_outputs(1474) <= '0';
    layer0_outputs(1475) <= inputs(246);
    layer0_outputs(1476) <= not(inputs(231));
    layer0_outputs(1477) <= (inputs(158)) and (inputs(233));
    layer0_outputs(1478) <= not((inputs(110)) or (inputs(70)));
    layer0_outputs(1479) <= not(inputs(70));
    layer0_outputs(1480) <= not(inputs(143));
    layer0_outputs(1481) <= (inputs(56)) and (inputs(11));
    layer0_outputs(1482) <= inputs(198);
    layer0_outputs(1483) <= not((inputs(237)) or (inputs(228)));
    layer0_outputs(1484) <= (inputs(61)) and (inputs(113));
    layer0_outputs(1485) <= (inputs(141)) and not (inputs(162));
    layer0_outputs(1486) <= not(inputs(161));
    layer0_outputs(1487) <= not(inputs(169)) or (inputs(223));
    layer0_outputs(1488) <= not(inputs(24));
    layer0_outputs(1489) <= (inputs(103)) and (inputs(68));
    layer0_outputs(1490) <= inputs(26);
    layer0_outputs(1491) <= not(inputs(62));
    layer0_outputs(1492) <= not((inputs(251)) xor (inputs(86)));
    layer0_outputs(1493) <= inputs(60);
    layer0_outputs(1494) <= not((inputs(115)) or (inputs(239)));
    layer0_outputs(1495) <= not(inputs(123));
    layer0_outputs(1496) <= (inputs(93)) xor (inputs(19));
    layer0_outputs(1497) <= inputs(230);
    layer0_outputs(1498) <= not(inputs(166));
    layer0_outputs(1499) <= not(inputs(136)) or (inputs(216));
    layer0_outputs(1500) <= not(inputs(121)) or (inputs(200));
    layer0_outputs(1501) <= (inputs(180)) and not (inputs(192));
    layer0_outputs(1502) <= inputs(22);
    layer0_outputs(1503) <= inputs(32);
    layer0_outputs(1504) <= not(inputs(235));
    layer0_outputs(1505) <= not((inputs(45)) and (inputs(206)));
    layer0_outputs(1506) <= (inputs(29)) and not (inputs(125));
    layer0_outputs(1507) <= inputs(214);
    layer0_outputs(1508) <= (inputs(225)) or (inputs(99));
    layer0_outputs(1509) <= (inputs(71)) and not (inputs(168));
    layer0_outputs(1510) <= not(inputs(210)) or (inputs(113));
    layer0_outputs(1511) <= inputs(99);
    layer0_outputs(1512) <= not((inputs(67)) or (inputs(119)));
    layer0_outputs(1513) <= (inputs(105)) and not (inputs(244));
    layer0_outputs(1514) <= '0';
    layer0_outputs(1515) <= not((inputs(46)) or (inputs(24)));
    layer0_outputs(1516) <= not(inputs(91)) or (inputs(19));
    layer0_outputs(1517) <= inputs(231);
    layer0_outputs(1518) <= not((inputs(90)) or (inputs(77)));
    layer0_outputs(1519) <= (inputs(46)) or (inputs(165));
    layer0_outputs(1520) <= (inputs(63)) and not (inputs(167));
    layer0_outputs(1521) <= (inputs(153)) or (inputs(242));
    layer0_outputs(1522) <= not((inputs(211)) and (inputs(27)));
    layer0_outputs(1523) <= not(inputs(235));
    layer0_outputs(1524) <= not((inputs(218)) xor (inputs(64)));
    layer0_outputs(1525) <= inputs(181);
    layer0_outputs(1526) <= (inputs(76)) or (inputs(126));
    layer0_outputs(1527) <= (inputs(103)) and not (inputs(219));
    layer0_outputs(1528) <= inputs(130);
    layer0_outputs(1529) <= (inputs(33)) and (inputs(69));
    layer0_outputs(1530) <= inputs(79);
    layer0_outputs(1531) <= not(inputs(110));
    layer0_outputs(1532) <= inputs(118);
    layer0_outputs(1533) <= (inputs(127)) or (inputs(63));
    layer0_outputs(1534) <= (inputs(106)) and not (inputs(133));
    layer0_outputs(1535) <= (inputs(135)) and not (inputs(127));
    layer0_outputs(1536) <= (inputs(45)) and (inputs(34));
    layer0_outputs(1537) <= (inputs(200)) xor (inputs(0));
    layer0_outputs(1538) <= inputs(98);
    layer0_outputs(1539) <= '0';
    layer0_outputs(1540) <= not((inputs(209)) and (inputs(141)));
    layer0_outputs(1541) <= (inputs(215)) and not (inputs(240));
    layer0_outputs(1542) <= not((inputs(57)) or (inputs(44)));
    layer0_outputs(1543) <= inputs(179);
    layer0_outputs(1544) <= not(inputs(151));
    layer0_outputs(1545) <= '0';
    layer0_outputs(1546) <= not((inputs(93)) xor (inputs(114)));
    layer0_outputs(1547) <= not(inputs(130)) or (inputs(185));
    layer0_outputs(1548) <= inputs(135);
    layer0_outputs(1549) <= '0';
    layer0_outputs(1550) <= not(inputs(164)) or (inputs(221));
    layer0_outputs(1551) <= not((inputs(223)) or (inputs(239)));
    layer0_outputs(1552) <= inputs(104);
    layer0_outputs(1553) <= '0';
    layer0_outputs(1554) <= (inputs(85)) or (inputs(113));
    layer0_outputs(1555) <= inputs(8);
    layer0_outputs(1556) <= (inputs(149)) and not (inputs(240));
    layer0_outputs(1557) <= (inputs(18)) or (inputs(49));
    layer0_outputs(1558) <= (inputs(254)) and not (inputs(237));
    layer0_outputs(1559) <= '1';
    layer0_outputs(1560) <= not(inputs(131));
    layer0_outputs(1561) <= inputs(131);
    layer0_outputs(1562) <= inputs(83);
    layer0_outputs(1563) <= (inputs(203)) and not (inputs(147));
    layer0_outputs(1564) <= not(inputs(192)) or (inputs(233));
    layer0_outputs(1565) <= (inputs(165)) or (inputs(70));
    layer0_outputs(1566) <= inputs(131);
    layer0_outputs(1567) <= not(inputs(137)) or (inputs(195));
    layer0_outputs(1568) <= not((inputs(9)) xor (inputs(41)));
    layer0_outputs(1569) <= not((inputs(78)) xor (inputs(217)));
    layer0_outputs(1570) <= not(inputs(236)) or (inputs(94));
    layer0_outputs(1571) <= not(inputs(248));
    layer0_outputs(1572) <= (inputs(245)) xor (inputs(214));
    layer0_outputs(1573) <= not((inputs(61)) xor (inputs(154)));
    layer0_outputs(1574) <= (inputs(61)) or (inputs(152));
    layer0_outputs(1575) <= (inputs(194)) or (inputs(104));
    layer0_outputs(1576) <= inputs(118);
    layer0_outputs(1577) <= '1';
    layer0_outputs(1578) <= '0';
    layer0_outputs(1579) <= (inputs(97)) or (inputs(32));
    layer0_outputs(1580) <= not(inputs(47));
    layer0_outputs(1581) <= (inputs(139)) or (inputs(117));
    layer0_outputs(1582) <= not((inputs(116)) or (inputs(118)));
    layer0_outputs(1583) <= '0';
    layer0_outputs(1584) <= not(inputs(39)) or (inputs(174));
    layer0_outputs(1585) <= (inputs(41)) or (inputs(64));
    layer0_outputs(1586) <= '0';
    layer0_outputs(1587) <= not(inputs(208)) or (inputs(48));
    layer0_outputs(1588) <= (inputs(62)) and not (inputs(31));
    layer0_outputs(1589) <= not(inputs(210)) or (inputs(146));
    layer0_outputs(1590) <= (inputs(218)) and (inputs(15));
    layer0_outputs(1591) <= not(inputs(147));
    layer0_outputs(1592) <= not(inputs(164));
    layer0_outputs(1593) <= inputs(62);
    layer0_outputs(1594) <= (inputs(209)) xor (inputs(233));
    layer0_outputs(1595) <= (inputs(174)) and (inputs(36));
    layer0_outputs(1596) <= not(inputs(239));
    layer0_outputs(1597) <= not(inputs(157));
    layer0_outputs(1598) <= inputs(251);
    layer0_outputs(1599) <= not(inputs(157)) or (inputs(134));
    layer0_outputs(1600) <= not(inputs(156)) or (inputs(224));
    layer0_outputs(1601) <= not(inputs(105));
    layer0_outputs(1602) <= (inputs(79)) or (inputs(89));
    layer0_outputs(1603) <= '0';
    layer0_outputs(1604) <= not(inputs(248)) or (inputs(133));
    layer0_outputs(1605) <= '1';
    layer0_outputs(1606) <= not(inputs(112));
    layer0_outputs(1607) <= not(inputs(229));
    layer0_outputs(1608) <= (inputs(86)) or (inputs(172));
    layer0_outputs(1609) <= not(inputs(3)) or (inputs(249));
    layer0_outputs(1610) <= not(inputs(120)) or (inputs(62));
    layer0_outputs(1611) <= inputs(60);
    layer0_outputs(1612) <= not(inputs(104));
    layer0_outputs(1613) <= (inputs(115)) or (inputs(131));
    layer0_outputs(1614) <= (inputs(200)) and not (inputs(126));
    layer0_outputs(1615) <= inputs(199);
    layer0_outputs(1616) <= (inputs(229)) and (inputs(105));
    layer0_outputs(1617) <= not(inputs(109)) or (inputs(64));
    layer0_outputs(1618) <= not((inputs(34)) or (inputs(218)));
    layer0_outputs(1619) <= not(inputs(72)) or (inputs(94));
    layer0_outputs(1620) <= not((inputs(87)) or (inputs(173)));
    layer0_outputs(1621) <= not((inputs(63)) xor (inputs(108)));
    layer0_outputs(1622) <= inputs(234);
    layer0_outputs(1623) <= (inputs(150)) and not (inputs(11));
    layer0_outputs(1624) <= not((inputs(150)) or (inputs(132)));
    layer0_outputs(1625) <= not(inputs(202)) or (inputs(12));
    layer0_outputs(1626) <= not((inputs(248)) or (inputs(146)));
    layer0_outputs(1627) <= not(inputs(117));
    layer0_outputs(1628) <= '0';
    layer0_outputs(1629) <= inputs(159);
    layer0_outputs(1630) <= not(inputs(25)) or (inputs(73));
    layer0_outputs(1631) <= (inputs(43)) or (inputs(191));
    layer0_outputs(1632) <= not(inputs(153));
    layer0_outputs(1633) <= not(inputs(211));
    layer0_outputs(1634) <= inputs(2);
    layer0_outputs(1635) <= not(inputs(101)) or (inputs(187));
    layer0_outputs(1636) <= (inputs(245)) or (inputs(98));
    layer0_outputs(1637) <= inputs(68);
    layer0_outputs(1638) <= not((inputs(123)) or (inputs(37)));
    layer0_outputs(1639) <= not(inputs(248));
    layer0_outputs(1640) <= inputs(143);
    layer0_outputs(1641) <= inputs(104);
    layer0_outputs(1642) <= (inputs(162)) or (inputs(159));
    layer0_outputs(1643) <= not((inputs(75)) or (inputs(92)));
    layer0_outputs(1644) <= inputs(172);
    layer0_outputs(1645) <= '0';
    layer0_outputs(1646) <= inputs(88);
    layer0_outputs(1647) <= (inputs(227)) and (inputs(252));
    layer0_outputs(1648) <= not(inputs(17)) or (inputs(199));
    layer0_outputs(1649) <= (inputs(215)) or (inputs(55));
    layer0_outputs(1650) <= (inputs(67)) or (inputs(97));
    layer0_outputs(1651) <= not(inputs(246));
    layer0_outputs(1652) <= inputs(120);
    layer0_outputs(1653) <= not(inputs(69));
    layer0_outputs(1654) <= inputs(76);
    layer0_outputs(1655) <= (inputs(189)) or (inputs(85));
    layer0_outputs(1656) <= not(inputs(33)) or (inputs(89));
    layer0_outputs(1657) <= (inputs(221)) or (inputs(132));
    layer0_outputs(1658) <= not(inputs(47)) or (inputs(70));
    layer0_outputs(1659) <= (inputs(91)) and not (inputs(144));
    layer0_outputs(1660) <= not((inputs(232)) and (inputs(73)));
    layer0_outputs(1661) <= not((inputs(89)) and (inputs(86)));
    layer0_outputs(1662) <= not(inputs(144));
    layer0_outputs(1663) <= not(inputs(247));
    layer0_outputs(1664) <= (inputs(109)) and not (inputs(37));
    layer0_outputs(1665) <= not(inputs(161)) or (inputs(188));
    layer0_outputs(1666) <= not(inputs(60));
    layer0_outputs(1667) <= not((inputs(28)) or (inputs(178)));
    layer0_outputs(1668) <= (inputs(95)) and (inputs(76));
    layer0_outputs(1669) <= inputs(123);
    layer0_outputs(1670) <= not(inputs(71));
    layer0_outputs(1671) <= not(inputs(46)) or (inputs(65));
    layer0_outputs(1672) <= inputs(125);
    layer0_outputs(1673) <= not((inputs(85)) xor (inputs(22)));
    layer0_outputs(1674) <= not(inputs(179));
    layer0_outputs(1675) <= inputs(100);
    layer0_outputs(1676) <= inputs(194);
    layer0_outputs(1677) <= not(inputs(214)) or (inputs(247));
    layer0_outputs(1678) <= (inputs(79)) or (inputs(62));
    layer0_outputs(1679) <= not(inputs(64));
    layer0_outputs(1680) <= not(inputs(24)) or (inputs(179));
    layer0_outputs(1681) <= not(inputs(140)) or (inputs(244));
    layer0_outputs(1682) <= (inputs(26)) or (inputs(243));
    layer0_outputs(1683) <= (inputs(46)) xor (inputs(171));
    layer0_outputs(1684) <= not((inputs(33)) and (inputs(94)));
    layer0_outputs(1685) <= not(inputs(244)) or (inputs(167));
    layer0_outputs(1686) <= not((inputs(225)) or (inputs(235)));
    layer0_outputs(1687) <= not((inputs(133)) xor (inputs(188)));
    layer0_outputs(1688) <= (inputs(150)) and not (inputs(249));
    layer0_outputs(1689) <= not(inputs(238));
    layer0_outputs(1690) <= inputs(228);
    layer0_outputs(1691) <= (inputs(219)) and not (inputs(59));
    layer0_outputs(1692) <= not((inputs(221)) or (inputs(254)));
    layer0_outputs(1693) <= (inputs(67)) or (inputs(86));
    layer0_outputs(1694) <= '0';
    layer0_outputs(1695) <= inputs(60);
    layer0_outputs(1696) <= (inputs(165)) and (inputs(175));
    layer0_outputs(1697) <= (inputs(209)) or (inputs(125));
    layer0_outputs(1698) <= not(inputs(82));
    layer0_outputs(1699) <= (inputs(162)) and (inputs(86));
    layer0_outputs(1700) <= '1';
    layer0_outputs(1701) <= not(inputs(164));
    layer0_outputs(1702) <= '0';
    layer0_outputs(1703) <= (inputs(238)) and not (inputs(34));
    layer0_outputs(1704) <= (inputs(118)) and (inputs(158));
    layer0_outputs(1705) <= not(inputs(238)) or (inputs(27));
    layer0_outputs(1706) <= (inputs(232)) or (inputs(35));
    layer0_outputs(1707) <= not(inputs(88));
    layer0_outputs(1708) <= '0';
    layer0_outputs(1709) <= not((inputs(54)) and (inputs(42)));
    layer0_outputs(1710) <= not(inputs(146)) or (inputs(29));
    layer0_outputs(1711) <= not(inputs(106));
    layer0_outputs(1712) <= inputs(18);
    layer0_outputs(1713) <= inputs(121);
    layer0_outputs(1714) <= '1';
    layer0_outputs(1715) <= inputs(162);
    layer0_outputs(1716) <= not(inputs(49));
    layer0_outputs(1717) <= (inputs(107)) or (inputs(58));
    layer0_outputs(1718) <= not(inputs(72));
    layer0_outputs(1719) <= inputs(174);
    layer0_outputs(1720) <= '1';
    layer0_outputs(1721) <= inputs(15);
    layer0_outputs(1722) <= not(inputs(131)) or (inputs(212));
    layer0_outputs(1723) <= not(inputs(12)) or (inputs(104));
    layer0_outputs(1724) <= not((inputs(98)) or (inputs(65)));
    layer0_outputs(1725) <= not((inputs(205)) or (inputs(174)));
    layer0_outputs(1726) <= (inputs(33)) and (inputs(251));
    layer0_outputs(1727) <= (inputs(159)) and not (inputs(19));
    layer0_outputs(1728) <= not(inputs(40));
    layer0_outputs(1729) <= (inputs(114)) and (inputs(137));
    layer0_outputs(1730) <= inputs(222);
    layer0_outputs(1731) <= (inputs(166)) and not (inputs(112));
    layer0_outputs(1732) <= (inputs(218)) and not (inputs(15));
    layer0_outputs(1733) <= not((inputs(99)) or (inputs(29)));
    layer0_outputs(1734) <= not((inputs(109)) and (inputs(155)));
    layer0_outputs(1735) <= not((inputs(220)) and (inputs(171)));
    layer0_outputs(1736) <= inputs(180);
    layer0_outputs(1737) <= '1';
    layer0_outputs(1738) <= not(inputs(83));
    layer0_outputs(1739) <= (inputs(222)) or (inputs(253));
    layer0_outputs(1740) <= (inputs(238)) and not (inputs(190));
    layer0_outputs(1741) <= (inputs(45)) and (inputs(251));
    layer0_outputs(1742) <= not(inputs(10));
    layer0_outputs(1743) <= inputs(21);
    layer0_outputs(1744) <= not(inputs(173));
    layer0_outputs(1745) <= not(inputs(182)) or (inputs(32));
    layer0_outputs(1746) <= (inputs(245)) or (inputs(143));
    layer0_outputs(1747) <= (inputs(36)) or (inputs(125));
    layer0_outputs(1748) <= (inputs(173)) and not (inputs(13));
    layer0_outputs(1749) <= not((inputs(133)) and (inputs(171)));
    layer0_outputs(1750) <= not(inputs(248));
    layer0_outputs(1751) <= not(inputs(174));
    layer0_outputs(1752) <= not(inputs(91));
    layer0_outputs(1753) <= (inputs(37)) and not (inputs(98));
    layer0_outputs(1754) <= not(inputs(166));
    layer0_outputs(1755) <= (inputs(25)) xor (inputs(192));
    layer0_outputs(1756) <= not((inputs(217)) and (inputs(16)));
    layer0_outputs(1757) <= '1';
    layer0_outputs(1758) <= not((inputs(68)) or (inputs(20)));
    layer0_outputs(1759) <= not(inputs(186)) or (inputs(169));
    layer0_outputs(1760) <= (inputs(42)) or (inputs(24));
    layer0_outputs(1761) <= (inputs(99)) or (inputs(98));
    layer0_outputs(1762) <= (inputs(92)) and not (inputs(200));
    layer0_outputs(1763) <= '0';
    layer0_outputs(1764) <= (inputs(218)) and not (inputs(109));
    layer0_outputs(1765) <= (inputs(140)) xor (inputs(240));
    layer0_outputs(1766) <= not((inputs(218)) and (inputs(168)));
    layer0_outputs(1767) <= not(inputs(8));
    layer0_outputs(1768) <= inputs(109);
    layer0_outputs(1769) <= not((inputs(240)) xor (inputs(177)));
    layer0_outputs(1770) <= not(inputs(251)) or (inputs(23));
    layer0_outputs(1771) <= not((inputs(184)) and (inputs(155)));
    layer0_outputs(1772) <= not((inputs(23)) or (inputs(126)));
    layer0_outputs(1773) <= (inputs(222)) and not (inputs(209));
    layer0_outputs(1774) <= not(inputs(119));
    layer0_outputs(1775) <= (inputs(66)) and not (inputs(215));
    layer0_outputs(1776) <= inputs(230);
    layer0_outputs(1777) <= not(inputs(84));
    layer0_outputs(1778) <= (inputs(148)) and not (inputs(236));
    layer0_outputs(1779) <= not(inputs(162));
    layer0_outputs(1780) <= '1';
    layer0_outputs(1781) <= '0';
    layer0_outputs(1782) <= not(inputs(145));
    layer0_outputs(1783) <= (inputs(108)) and (inputs(170));
    layer0_outputs(1784) <= (inputs(194)) or (inputs(80));
    layer0_outputs(1785) <= (inputs(34)) or (inputs(192));
    layer0_outputs(1786) <= not(inputs(162));
    layer0_outputs(1787) <= not((inputs(108)) or (inputs(117)));
    layer0_outputs(1788) <= not((inputs(106)) or (inputs(6)));
    layer0_outputs(1789) <= not(inputs(155));
    layer0_outputs(1790) <= not((inputs(173)) or (inputs(21)));
    layer0_outputs(1791) <= (inputs(21)) and not (inputs(82));
    layer0_outputs(1792) <= (inputs(94)) and not (inputs(217));
    layer0_outputs(1793) <= inputs(10);
    layer0_outputs(1794) <= not(inputs(93)) or (inputs(15));
    layer0_outputs(1795) <= not(inputs(233));
    layer0_outputs(1796) <= '0';
    layer0_outputs(1797) <= inputs(81);
    layer0_outputs(1798) <= inputs(152);
    layer0_outputs(1799) <= (inputs(88)) xor (inputs(62));
    layer0_outputs(1800) <= inputs(120);
    layer0_outputs(1801) <= (inputs(231)) and not (inputs(15));
    layer0_outputs(1802) <= not((inputs(139)) xor (inputs(139)));
    layer0_outputs(1803) <= (inputs(49)) and not (inputs(82));
    layer0_outputs(1804) <= not(inputs(226)) or (inputs(175));
    layer0_outputs(1805) <= not(inputs(98)) or (inputs(130));
    layer0_outputs(1806) <= (inputs(41)) or (inputs(226));
    layer0_outputs(1807) <= (inputs(132)) and not (inputs(139));
    layer0_outputs(1808) <= (inputs(145)) xor (inputs(8));
    layer0_outputs(1809) <= not((inputs(79)) or (inputs(8)));
    layer0_outputs(1810) <= (inputs(103)) or (inputs(249));
    layer0_outputs(1811) <= not((inputs(144)) and (inputs(36)));
    layer0_outputs(1812) <= not(inputs(101));
    layer0_outputs(1813) <= not((inputs(72)) and (inputs(69)));
    layer0_outputs(1814) <= inputs(161);
    layer0_outputs(1815) <= (inputs(41)) or (inputs(62));
    layer0_outputs(1816) <= not(inputs(165));
    layer0_outputs(1817) <= not(inputs(219)) or (inputs(244));
    layer0_outputs(1818) <= not((inputs(120)) or (inputs(114)));
    layer0_outputs(1819) <= not((inputs(59)) or (inputs(74)));
    layer0_outputs(1820) <= inputs(116);
    layer0_outputs(1821) <= '1';
    layer0_outputs(1822) <= (inputs(38)) or (inputs(152));
    layer0_outputs(1823) <= '1';
    layer0_outputs(1824) <= not(inputs(120));
    layer0_outputs(1825) <= not(inputs(157)) or (inputs(18));
    layer0_outputs(1826) <= '0';
    layer0_outputs(1827) <= inputs(25);
    layer0_outputs(1828) <= not(inputs(119));
    layer0_outputs(1829) <= not((inputs(97)) or (inputs(100)));
    layer0_outputs(1830) <= not(inputs(207));
    layer0_outputs(1831) <= inputs(245);
    layer0_outputs(1832) <= (inputs(205)) and not (inputs(7));
    layer0_outputs(1833) <= (inputs(125)) and (inputs(59));
    layer0_outputs(1834) <= not(inputs(186));
    layer0_outputs(1835) <= not(inputs(118)) or (inputs(241));
    layer0_outputs(1836) <= not(inputs(2));
    layer0_outputs(1837) <= (inputs(173)) or (inputs(7));
    layer0_outputs(1838) <= (inputs(228)) and not (inputs(7));
    layer0_outputs(1839) <= inputs(44);
    layer0_outputs(1840) <= not(inputs(68)) or (inputs(103));
    layer0_outputs(1841) <= inputs(226);
    layer0_outputs(1842) <= (inputs(103)) xor (inputs(80));
    layer0_outputs(1843) <= not(inputs(191)) or (inputs(209));
    layer0_outputs(1844) <= inputs(229);
    layer0_outputs(1845) <= not(inputs(213)) or (inputs(87));
    layer0_outputs(1846) <= inputs(71);
    layer0_outputs(1847) <= not(inputs(197));
    layer0_outputs(1848) <= inputs(41);
    layer0_outputs(1849) <= not(inputs(30));
    layer0_outputs(1850) <= not(inputs(80)) or (inputs(151));
    layer0_outputs(1851) <= (inputs(50)) or (inputs(25));
    layer0_outputs(1852) <= inputs(249);
    layer0_outputs(1853) <= inputs(130);
    layer0_outputs(1854) <= (inputs(18)) and not (inputs(32));
    layer0_outputs(1855) <= not((inputs(136)) xor (inputs(2)));
    layer0_outputs(1856) <= (inputs(233)) or (inputs(53));
    layer0_outputs(1857) <= not(inputs(123)) or (inputs(188));
    layer0_outputs(1858) <= (inputs(37)) and not (inputs(2));
    layer0_outputs(1859) <= not((inputs(222)) or (inputs(230)));
    layer0_outputs(1860) <= not(inputs(193));
    layer0_outputs(1861) <= (inputs(105)) and not (inputs(111));
    layer0_outputs(1862) <= (inputs(182)) or (inputs(220));
    layer0_outputs(1863) <= inputs(231);
    layer0_outputs(1864) <= inputs(231);
    layer0_outputs(1865) <= not(inputs(138));
    layer0_outputs(1866) <= (inputs(170)) and not (inputs(21));
    layer0_outputs(1867) <= not(inputs(213)) or (inputs(63));
    layer0_outputs(1868) <= not((inputs(70)) xor (inputs(26)));
    layer0_outputs(1869) <= not(inputs(5));
    layer0_outputs(1870) <= inputs(141);
    layer0_outputs(1871) <= inputs(190);
    layer0_outputs(1872) <= not(inputs(95));
    layer0_outputs(1873) <= not(inputs(236)) or (inputs(243));
    layer0_outputs(1874) <= (inputs(135)) and not (inputs(197));
    layer0_outputs(1875) <= (inputs(156)) or (inputs(75));
    layer0_outputs(1876) <= '1';
    layer0_outputs(1877) <= (inputs(217)) and not (inputs(3));
    layer0_outputs(1878) <= not((inputs(215)) and (inputs(250)));
    layer0_outputs(1879) <= (inputs(52)) or (inputs(48));
    layer0_outputs(1880) <= not((inputs(177)) xor (inputs(235)));
    layer0_outputs(1881) <= inputs(188);
    layer0_outputs(1882) <= not(inputs(137));
    layer0_outputs(1883) <= (inputs(225)) or (inputs(141));
    layer0_outputs(1884) <= '0';
    layer0_outputs(1885) <= not(inputs(170));
    layer0_outputs(1886) <= (inputs(64)) or (inputs(95));
    layer0_outputs(1887) <= (inputs(14)) and (inputs(64));
    layer0_outputs(1888) <= not((inputs(18)) or (inputs(246)));
    layer0_outputs(1889) <= not(inputs(213));
    layer0_outputs(1890) <= not(inputs(76));
    layer0_outputs(1891) <= inputs(83);
    layer0_outputs(1892) <= not((inputs(131)) or (inputs(93)));
    layer0_outputs(1893) <= not(inputs(164));
    layer0_outputs(1894) <= not(inputs(163)) or (inputs(139));
    layer0_outputs(1895) <= not((inputs(66)) or (inputs(123)));
    layer0_outputs(1896) <= (inputs(104)) or (inputs(90));
    layer0_outputs(1897) <= not(inputs(98));
    layer0_outputs(1898) <= (inputs(195)) or (inputs(240));
    layer0_outputs(1899) <= (inputs(220)) or (inputs(146));
    layer0_outputs(1900) <= inputs(217);
    layer0_outputs(1901) <= (inputs(234)) or (inputs(246));
    layer0_outputs(1902) <= (inputs(225)) and (inputs(63));
    layer0_outputs(1903) <= (inputs(107)) and not (inputs(15));
    layer0_outputs(1904) <= not(inputs(36));
    layer0_outputs(1905) <= (inputs(36)) and not (inputs(131));
    layer0_outputs(1906) <= (inputs(120)) or (inputs(106));
    layer0_outputs(1907) <= (inputs(12)) xor (inputs(25));
    layer0_outputs(1908) <= (inputs(136)) xor (inputs(34));
    layer0_outputs(1909) <= (inputs(84)) xor (inputs(148));
    layer0_outputs(1910) <= not(inputs(130));
    layer0_outputs(1911) <= not(inputs(92));
    layer0_outputs(1912) <= (inputs(30)) xor (inputs(172));
    layer0_outputs(1913) <= (inputs(148)) and not (inputs(186));
    layer0_outputs(1914) <= inputs(201);
    layer0_outputs(1915) <= (inputs(143)) and not (inputs(158));
    layer0_outputs(1916) <= inputs(42);
    layer0_outputs(1917) <= (inputs(180)) and not (inputs(229));
    layer0_outputs(1918) <= (inputs(226)) or (inputs(87));
    layer0_outputs(1919) <= inputs(253);
    layer0_outputs(1920) <= not(inputs(84));
    layer0_outputs(1921) <= (inputs(167)) or (inputs(189));
    layer0_outputs(1922) <= inputs(146);
    layer0_outputs(1923) <= not(inputs(124));
    layer0_outputs(1924) <= not(inputs(191));
    layer0_outputs(1925) <= (inputs(193)) and not (inputs(148));
    layer0_outputs(1926) <= (inputs(11)) and not (inputs(83));
    layer0_outputs(1927) <= not(inputs(214));
    layer0_outputs(1928) <= '1';
    layer0_outputs(1929) <= not(inputs(99)) or (inputs(115));
    layer0_outputs(1930) <= not(inputs(196));
    layer0_outputs(1931) <= (inputs(145)) or (inputs(66));
    layer0_outputs(1932) <= inputs(87);
    layer0_outputs(1933) <= not(inputs(83));
    layer0_outputs(1934) <= (inputs(209)) and (inputs(104));
    layer0_outputs(1935) <= not((inputs(182)) or (inputs(84)));
    layer0_outputs(1936) <= '1';
    layer0_outputs(1937) <= inputs(24);
    layer0_outputs(1938) <= (inputs(194)) and not (inputs(201));
    layer0_outputs(1939) <= not(inputs(111));
    layer0_outputs(1940) <= inputs(58);
    layer0_outputs(1941) <= (inputs(175)) and not (inputs(208));
    layer0_outputs(1942) <= not((inputs(48)) xor (inputs(176)));
    layer0_outputs(1943) <= '1';
    layer0_outputs(1944) <= '1';
    layer0_outputs(1945) <= not(inputs(94));
    layer0_outputs(1946) <= '0';
    layer0_outputs(1947) <= not(inputs(78));
    layer0_outputs(1948) <= (inputs(53)) or (inputs(37));
    layer0_outputs(1949) <= (inputs(1)) or (inputs(71));
    layer0_outputs(1950) <= (inputs(220)) or (inputs(115));
    layer0_outputs(1951) <= inputs(15);
    layer0_outputs(1952) <= (inputs(244)) or (inputs(33));
    layer0_outputs(1953) <= inputs(219);
    layer0_outputs(1954) <= not(inputs(154)) or (inputs(115));
    layer0_outputs(1955) <= inputs(28);
    layer0_outputs(1956) <= inputs(66);
    layer0_outputs(1957) <= (inputs(203)) or (inputs(189));
    layer0_outputs(1958) <= '1';
    layer0_outputs(1959) <= inputs(83);
    layer0_outputs(1960) <= inputs(108);
    layer0_outputs(1961) <= not(inputs(206)) or (inputs(80));
    layer0_outputs(1962) <= inputs(8);
    layer0_outputs(1963) <= not(inputs(131));
    layer0_outputs(1964) <= (inputs(231)) and not (inputs(65));
    layer0_outputs(1965) <= not(inputs(131)) or (inputs(223));
    layer0_outputs(1966) <= not(inputs(169)) or (inputs(47));
    layer0_outputs(1967) <= not(inputs(71)) or (inputs(32));
    layer0_outputs(1968) <= '1';
    layer0_outputs(1969) <= (inputs(71)) and not (inputs(148));
    layer0_outputs(1970) <= not(inputs(24)) or (inputs(131));
    layer0_outputs(1971) <= not((inputs(178)) or (inputs(199)));
    layer0_outputs(1972) <= not(inputs(14));
    layer0_outputs(1973) <= not((inputs(197)) and (inputs(8)));
    layer0_outputs(1974) <= inputs(72);
    layer0_outputs(1975) <= inputs(25);
    layer0_outputs(1976) <= not(inputs(85)) or (inputs(210));
    layer0_outputs(1977) <= inputs(211);
    layer0_outputs(1978) <= '0';
    layer0_outputs(1979) <= inputs(101);
    layer0_outputs(1980) <= '1';
    layer0_outputs(1981) <= not((inputs(203)) or (inputs(194)));
    layer0_outputs(1982) <= not(inputs(133));
    layer0_outputs(1983) <= not(inputs(219));
    layer0_outputs(1984) <= not(inputs(55)) or (inputs(3));
    layer0_outputs(1985) <= inputs(27);
    layer0_outputs(1986) <= not(inputs(96));
    layer0_outputs(1987) <= (inputs(109)) xor (inputs(158));
    layer0_outputs(1988) <= not((inputs(219)) or (inputs(185)));
    layer0_outputs(1989) <= not(inputs(37));
    layer0_outputs(1990) <= not(inputs(24));
    layer0_outputs(1991) <= not((inputs(49)) or (inputs(241)));
    layer0_outputs(1992) <= inputs(115);
    layer0_outputs(1993) <= (inputs(30)) or (inputs(241));
    layer0_outputs(1994) <= not((inputs(211)) or (inputs(173)));
    layer0_outputs(1995) <= not(inputs(188));
    layer0_outputs(1996) <= (inputs(17)) or (inputs(74));
    layer0_outputs(1997) <= not((inputs(71)) and (inputs(146)));
    layer0_outputs(1998) <= (inputs(26)) and not (inputs(157));
    layer0_outputs(1999) <= (inputs(6)) or (inputs(23));
    layer0_outputs(2000) <= (inputs(194)) and (inputs(175));
    layer0_outputs(2001) <= not(inputs(197)) or (inputs(166));
    layer0_outputs(2002) <= not(inputs(67));
    layer0_outputs(2003) <= not((inputs(76)) xor (inputs(198)));
    layer0_outputs(2004) <= not((inputs(44)) or (inputs(43)));
    layer0_outputs(2005) <= not(inputs(157)) or (inputs(83));
    layer0_outputs(2006) <= not((inputs(149)) and (inputs(85)));
    layer0_outputs(2007) <= not((inputs(84)) or (inputs(78)));
    layer0_outputs(2008) <= not(inputs(124));
    layer0_outputs(2009) <= not((inputs(137)) and (inputs(48)));
    layer0_outputs(2010) <= (inputs(205)) or (inputs(179));
    layer0_outputs(2011) <= (inputs(247)) and not (inputs(125));
    layer0_outputs(2012) <= (inputs(218)) and not (inputs(108));
    layer0_outputs(2013) <= not((inputs(38)) or (inputs(176)));
    layer0_outputs(2014) <= not((inputs(138)) or (inputs(104)));
    layer0_outputs(2015) <= (inputs(152)) and not (inputs(74));
    layer0_outputs(2016) <= not(inputs(178));
    layer0_outputs(2017) <= not(inputs(144)) or (inputs(236));
    layer0_outputs(2018) <= (inputs(125)) and not (inputs(31));
    layer0_outputs(2019) <= not(inputs(184));
    layer0_outputs(2020) <= not(inputs(120)) or (inputs(206));
    layer0_outputs(2021) <= not(inputs(131));
    layer0_outputs(2022) <= not(inputs(159)) or (inputs(74));
    layer0_outputs(2023) <= (inputs(98)) and (inputs(18));
    layer0_outputs(2024) <= inputs(70);
    layer0_outputs(2025) <= (inputs(32)) or (inputs(25));
    layer0_outputs(2026) <= inputs(184);
    layer0_outputs(2027) <= not(inputs(230));
    layer0_outputs(2028) <= not(inputs(43));
    layer0_outputs(2029) <= '1';
    layer0_outputs(2030) <= not((inputs(101)) xor (inputs(108)));
    layer0_outputs(2031) <= not(inputs(65)) or (inputs(21));
    layer0_outputs(2032) <= not((inputs(238)) and (inputs(22)));
    layer0_outputs(2033) <= (inputs(136)) or (inputs(222));
    layer0_outputs(2034) <= not((inputs(77)) or (inputs(69)));
    layer0_outputs(2035) <= (inputs(136)) or (inputs(55));
    layer0_outputs(2036) <= not((inputs(164)) xor (inputs(128)));
    layer0_outputs(2037) <= not(inputs(253)) or (inputs(222));
    layer0_outputs(2038) <= not(inputs(75));
    layer0_outputs(2039) <= not((inputs(14)) or (inputs(245)));
    layer0_outputs(2040) <= inputs(168);
    layer0_outputs(2041) <= not(inputs(25)) or (inputs(210));
    layer0_outputs(2042) <= not(inputs(18)) or (inputs(76));
    layer0_outputs(2043) <= '0';
    layer0_outputs(2044) <= not(inputs(107));
    layer0_outputs(2045) <= inputs(83);
    layer0_outputs(2046) <= inputs(80);
    layer0_outputs(2047) <= not(inputs(27));
    layer0_outputs(2048) <= not((inputs(72)) and (inputs(65)));
    layer0_outputs(2049) <= not(inputs(241));
    layer0_outputs(2050) <= not((inputs(142)) or (inputs(156)));
    layer0_outputs(2051) <= not(inputs(79)) or (inputs(87));
    layer0_outputs(2052) <= not((inputs(21)) or (inputs(0)));
    layer0_outputs(2053) <= not((inputs(181)) or (inputs(151)));
    layer0_outputs(2054) <= not((inputs(237)) or (inputs(166)));
    layer0_outputs(2055) <= not((inputs(236)) xor (inputs(218)));
    layer0_outputs(2056) <= (inputs(12)) and not (inputs(3));
    layer0_outputs(2057) <= not((inputs(32)) and (inputs(14)));
    layer0_outputs(2058) <= (inputs(178)) or (inputs(52));
    layer0_outputs(2059) <= (inputs(33)) and (inputs(216));
    layer0_outputs(2060) <= (inputs(136)) xor (inputs(255));
    layer0_outputs(2061) <= (inputs(205)) or (inputs(206));
    layer0_outputs(2062) <= not(inputs(42));
    layer0_outputs(2063) <= (inputs(162)) and not (inputs(215));
    layer0_outputs(2064) <= not((inputs(79)) and (inputs(80)));
    layer0_outputs(2065) <= not(inputs(22));
    layer0_outputs(2066) <= not((inputs(46)) xor (inputs(27)));
    layer0_outputs(2067) <= not(inputs(62)) or (inputs(255));
    layer0_outputs(2068) <= (inputs(240)) and not (inputs(15));
    layer0_outputs(2069) <= not((inputs(4)) or (inputs(240)));
    layer0_outputs(2070) <= not(inputs(252));
    layer0_outputs(2071) <= inputs(102);
    layer0_outputs(2072) <= not(inputs(143));
    layer0_outputs(2073) <= '0';
    layer0_outputs(2074) <= (inputs(117)) or (inputs(98));
    layer0_outputs(2075) <= inputs(139);
    layer0_outputs(2076) <= '0';
    layer0_outputs(2077) <= not(inputs(187));
    layer0_outputs(2078) <= not(inputs(129));
    layer0_outputs(2079) <= inputs(139);
    layer0_outputs(2080) <= (inputs(185)) xor (inputs(232));
    layer0_outputs(2081) <= '0';
    layer0_outputs(2082) <= not(inputs(37)) or (inputs(131));
    layer0_outputs(2083) <= not(inputs(110));
    layer0_outputs(2084) <= not(inputs(193));
    layer0_outputs(2085) <= '1';
    layer0_outputs(2086) <= not((inputs(65)) and (inputs(150)));
    layer0_outputs(2087) <= inputs(100);
    layer0_outputs(2088) <= not((inputs(222)) or (inputs(206)));
    layer0_outputs(2089) <= not(inputs(53)) or (inputs(155));
    layer0_outputs(2090) <= inputs(172);
    layer0_outputs(2091) <= inputs(147);
    layer0_outputs(2092) <= (inputs(237)) or (inputs(52));
    layer0_outputs(2093) <= not(inputs(236)) or (inputs(67));
    layer0_outputs(2094) <= not(inputs(148));
    layer0_outputs(2095) <= inputs(57);
    layer0_outputs(2096) <= inputs(126);
    layer0_outputs(2097) <= '0';
    layer0_outputs(2098) <= not(inputs(158)) or (inputs(53));
    layer0_outputs(2099) <= (inputs(152)) and not (inputs(188));
    layer0_outputs(2100) <= not((inputs(16)) or (inputs(42)));
    layer0_outputs(2101) <= (inputs(254)) and not (inputs(15));
    layer0_outputs(2102) <= (inputs(83)) or (inputs(101));
    layer0_outputs(2103) <= not(inputs(123)) or (inputs(86));
    layer0_outputs(2104) <= inputs(142);
    layer0_outputs(2105) <= (inputs(230)) and not (inputs(97));
    layer0_outputs(2106) <= not((inputs(133)) or (inputs(161)));
    layer0_outputs(2107) <= not(inputs(166));
    layer0_outputs(2108) <= not(inputs(79)) or (inputs(214));
    layer0_outputs(2109) <= '0';
    layer0_outputs(2110) <= not((inputs(55)) or (inputs(69)));
    layer0_outputs(2111) <= '0';
    layer0_outputs(2112) <= (inputs(64)) or (inputs(82));
    layer0_outputs(2113) <= (inputs(31)) or (inputs(134));
    layer0_outputs(2114) <= (inputs(197)) and not (inputs(57));
    layer0_outputs(2115) <= not((inputs(6)) xor (inputs(10)));
    layer0_outputs(2116) <= inputs(178);
    layer0_outputs(2117) <= '1';
    layer0_outputs(2118) <= (inputs(81)) and not (inputs(118));
    layer0_outputs(2119) <= not((inputs(250)) and (inputs(0)));
    layer0_outputs(2120) <= '0';
    layer0_outputs(2121) <= not((inputs(12)) xor (inputs(45)));
    layer0_outputs(2122) <= '1';
    layer0_outputs(2123) <= not(inputs(156)) or (inputs(80));
    layer0_outputs(2124) <= not(inputs(72));
    layer0_outputs(2125) <= not(inputs(57));
    layer0_outputs(2126) <= '0';
    layer0_outputs(2127) <= (inputs(138)) or (inputs(80));
    layer0_outputs(2128) <= not(inputs(104));
    layer0_outputs(2129) <= not(inputs(199)) or (inputs(63));
    layer0_outputs(2130) <= (inputs(21)) xor (inputs(205));
    layer0_outputs(2131) <= not(inputs(180)) or (inputs(13));
    layer0_outputs(2132) <= not(inputs(8)) or (inputs(25));
    layer0_outputs(2133) <= not(inputs(197));
    layer0_outputs(2134) <= (inputs(95)) xor (inputs(99));
    layer0_outputs(2135) <= (inputs(172)) and not (inputs(94));
    layer0_outputs(2136) <= not(inputs(118));
    layer0_outputs(2137) <= (inputs(181)) xor (inputs(183));
    layer0_outputs(2138) <= not((inputs(118)) or (inputs(133)));
    layer0_outputs(2139) <= not((inputs(112)) or (inputs(223)));
    layer0_outputs(2140) <= not(inputs(35)) or (inputs(199));
    layer0_outputs(2141) <= (inputs(128)) xor (inputs(146));
    layer0_outputs(2142) <= (inputs(100)) and not (inputs(245));
    layer0_outputs(2143) <= not(inputs(91)) or (inputs(55));
    layer0_outputs(2144) <= inputs(89);
    layer0_outputs(2145) <= not((inputs(136)) or (inputs(134)));
    layer0_outputs(2146) <= not(inputs(47)) or (inputs(7));
    layer0_outputs(2147) <= not(inputs(118)) or (inputs(18));
    layer0_outputs(2148) <= (inputs(187)) and not (inputs(149));
    layer0_outputs(2149) <= inputs(158);
    layer0_outputs(2150) <= '1';
    layer0_outputs(2151) <= (inputs(182)) and not (inputs(185));
    layer0_outputs(2152) <= (inputs(48)) or (inputs(126));
    layer0_outputs(2153) <= (inputs(128)) and (inputs(156));
    layer0_outputs(2154) <= not(inputs(181)) or (inputs(169));
    layer0_outputs(2155) <= inputs(44);
    layer0_outputs(2156) <= (inputs(161)) xor (inputs(244));
    layer0_outputs(2157) <= '0';
    layer0_outputs(2158) <= (inputs(12)) and not (inputs(200));
    layer0_outputs(2159) <= inputs(77);
    layer0_outputs(2160) <= inputs(150);
    layer0_outputs(2161) <= inputs(145);
    layer0_outputs(2162) <= not((inputs(143)) or (inputs(218)));
    layer0_outputs(2163) <= not(inputs(30));
    layer0_outputs(2164) <= (inputs(78)) xor (inputs(0));
    layer0_outputs(2165) <= not(inputs(206));
    layer0_outputs(2166) <= not((inputs(88)) and (inputs(96)));
    layer0_outputs(2167) <= (inputs(146)) and not (inputs(43));
    layer0_outputs(2168) <= not(inputs(65));
    layer0_outputs(2169) <= (inputs(119)) and not (inputs(233));
    layer0_outputs(2170) <= (inputs(33)) and not (inputs(62));
    layer0_outputs(2171) <= not(inputs(245));
    layer0_outputs(2172) <= (inputs(22)) and not (inputs(183));
    layer0_outputs(2173) <= not((inputs(245)) and (inputs(149)));
    layer0_outputs(2174) <= not(inputs(114)) or (inputs(49));
    layer0_outputs(2175) <= not(inputs(8)) or (inputs(32));
    layer0_outputs(2176) <= inputs(75);
    layer0_outputs(2177) <= not(inputs(193));
    layer0_outputs(2178) <= '0';
    layer0_outputs(2179) <= not((inputs(229)) or (inputs(251)));
    layer0_outputs(2180) <= not(inputs(4));
    layer0_outputs(2181) <= inputs(105);
    layer0_outputs(2182) <= inputs(167);
    layer0_outputs(2183) <= not((inputs(67)) xor (inputs(70)));
    layer0_outputs(2184) <= not(inputs(129));
    layer0_outputs(2185) <= not(inputs(199));
    layer0_outputs(2186) <= '1';
    layer0_outputs(2187) <= (inputs(33)) and (inputs(214));
    layer0_outputs(2188) <= inputs(99);
    layer0_outputs(2189) <= not(inputs(104));
    layer0_outputs(2190) <= not((inputs(211)) or (inputs(67)));
    layer0_outputs(2191) <= (inputs(96)) and not (inputs(222));
    layer0_outputs(2192) <= not(inputs(239));
    layer0_outputs(2193) <= inputs(249);
    layer0_outputs(2194) <= not((inputs(101)) xor (inputs(99)));
    layer0_outputs(2195) <= inputs(14);
    layer0_outputs(2196) <= not(inputs(180));
    layer0_outputs(2197) <= not(inputs(19));
    layer0_outputs(2198) <= not(inputs(224));
    layer0_outputs(2199) <= not(inputs(243));
    layer0_outputs(2200) <= not(inputs(31));
    layer0_outputs(2201) <= not(inputs(191)) or (inputs(143));
    layer0_outputs(2202) <= not(inputs(174));
    layer0_outputs(2203) <= not(inputs(126));
    layer0_outputs(2204) <= (inputs(202)) or (inputs(254));
    layer0_outputs(2205) <= not(inputs(161));
    layer0_outputs(2206) <= (inputs(153)) and not (inputs(42));
    layer0_outputs(2207) <= inputs(147);
    layer0_outputs(2208) <= not((inputs(20)) and (inputs(185)));
    layer0_outputs(2209) <= '0';
    layer0_outputs(2210) <= '1';
    layer0_outputs(2211) <= not(inputs(84));
    layer0_outputs(2212) <= not((inputs(158)) and (inputs(214)));
    layer0_outputs(2213) <= not(inputs(241)) or (inputs(42));
    layer0_outputs(2214) <= not(inputs(150));
    layer0_outputs(2215) <= (inputs(119)) or (inputs(122));
    layer0_outputs(2216) <= '0';
    layer0_outputs(2217) <= (inputs(27)) and not (inputs(146));
    layer0_outputs(2218) <= not((inputs(38)) or (inputs(165)));
    layer0_outputs(2219) <= not((inputs(17)) or (inputs(192)));
    layer0_outputs(2220) <= not((inputs(156)) or (inputs(118)));
    layer0_outputs(2221) <= not(inputs(68));
    layer0_outputs(2222) <= not(inputs(7)) or (inputs(106));
    layer0_outputs(2223) <= not(inputs(234));
    layer0_outputs(2224) <= not((inputs(51)) and (inputs(179)));
    layer0_outputs(2225) <= not(inputs(230)) or (inputs(79));
    layer0_outputs(2226) <= inputs(58);
    layer0_outputs(2227) <= inputs(148);
    layer0_outputs(2228) <= not(inputs(27));
    layer0_outputs(2229) <= (inputs(24)) and not (inputs(103));
    layer0_outputs(2230) <= (inputs(208)) or (inputs(205));
    layer0_outputs(2231) <= (inputs(233)) or (inputs(224));
    layer0_outputs(2232) <= inputs(84);
    layer0_outputs(2233) <= (inputs(126)) and not (inputs(19));
    layer0_outputs(2234) <= not((inputs(43)) or (inputs(17)));
    layer0_outputs(2235) <= (inputs(191)) and not (inputs(11));
    layer0_outputs(2236) <= not(inputs(210));
    layer0_outputs(2237) <= not(inputs(161));
    layer0_outputs(2238) <= (inputs(147)) and not (inputs(122));
    layer0_outputs(2239) <= not((inputs(227)) xor (inputs(78)));
    layer0_outputs(2240) <= (inputs(4)) or (inputs(19));
    layer0_outputs(2241) <= (inputs(219)) and not (inputs(151));
    layer0_outputs(2242) <= inputs(4);
    layer0_outputs(2243) <= (inputs(21)) and not (inputs(54));
    layer0_outputs(2244) <= not(inputs(177));
    layer0_outputs(2245) <= not(inputs(232));
    layer0_outputs(2246) <= (inputs(47)) and not (inputs(71));
    layer0_outputs(2247) <= not(inputs(139)) or (inputs(27));
    layer0_outputs(2248) <= (inputs(237)) xor (inputs(149));
    layer0_outputs(2249) <= (inputs(95)) and not (inputs(251));
    layer0_outputs(2250) <= '0';
    layer0_outputs(2251) <= not(inputs(34));
    layer0_outputs(2252) <= not(inputs(153));
    layer0_outputs(2253) <= inputs(145);
    layer0_outputs(2254) <= inputs(89);
    layer0_outputs(2255) <= not(inputs(182)) or (inputs(177));
    layer0_outputs(2256) <= '0';
    layer0_outputs(2257) <= not(inputs(90));
    layer0_outputs(2258) <= inputs(231);
    layer0_outputs(2259) <= (inputs(160)) and not (inputs(152));
    layer0_outputs(2260) <= inputs(90);
    layer0_outputs(2261) <= (inputs(18)) and not (inputs(92));
    layer0_outputs(2262) <= (inputs(139)) and not (inputs(95));
    layer0_outputs(2263) <= inputs(97);
    layer0_outputs(2264) <= not(inputs(104)) or (inputs(208));
    layer0_outputs(2265) <= not((inputs(101)) or (inputs(249)));
    layer0_outputs(2266) <= (inputs(60)) and (inputs(147));
    layer0_outputs(2267) <= not(inputs(123));
    layer0_outputs(2268) <= not((inputs(174)) xor (inputs(223)));
    layer0_outputs(2269) <= (inputs(46)) or (inputs(17));
    layer0_outputs(2270) <= not(inputs(111));
    layer0_outputs(2271) <= (inputs(83)) and not (inputs(143));
    layer0_outputs(2272) <= (inputs(193)) and not (inputs(101));
    layer0_outputs(2273) <= '1';
    layer0_outputs(2274) <= not(inputs(29));
    layer0_outputs(2275) <= not(inputs(19));
    layer0_outputs(2276) <= inputs(220);
    layer0_outputs(2277) <= not((inputs(242)) or (inputs(43)));
    layer0_outputs(2278) <= not((inputs(75)) xor (inputs(92)));
    layer0_outputs(2279) <= (inputs(216)) xor (inputs(207));
    layer0_outputs(2280) <= '0';
    layer0_outputs(2281) <= (inputs(209)) or (inputs(4));
    layer0_outputs(2282) <= (inputs(171)) or (inputs(31));
    layer0_outputs(2283) <= not((inputs(149)) or (inputs(107)));
    layer0_outputs(2284) <= '1';
    layer0_outputs(2285) <= not(inputs(119)) or (inputs(218));
    layer0_outputs(2286) <= '1';
    layer0_outputs(2287) <= not(inputs(164));
    layer0_outputs(2288) <= not(inputs(4));
    layer0_outputs(2289) <= not((inputs(87)) and (inputs(215)));
    layer0_outputs(2290) <= not((inputs(158)) and (inputs(19)));
    layer0_outputs(2291) <= not((inputs(17)) and (inputs(225)));
    layer0_outputs(2292) <= not(inputs(131));
    layer0_outputs(2293) <= not(inputs(212)) or (inputs(105));
    layer0_outputs(2294) <= not(inputs(176)) or (inputs(5));
    layer0_outputs(2295) <= not((inputs(253)) or (inputs(245)));
    layer0_outputs(2296) <= not(inputs(177));
    layer0_outputs(2297) <= (inputs(139)) and not (inputs(206));
    layer0_outputs(2298) <= not(inputs(211)) or (inputs(88));
    layer0_outputs(2299) <= not(inputs(21));
    layer0_outputs(2300) <= not(inputs(193));
    layer0_outputs(2301) <= not((inputs(210)) and (inputs(250)));
    layer0_outputs(2302) <= inputs(223);
    layer0_outputs(2303) <= not((inputs(220)) or (inputs(207)));
    layer0_outputs(2304) <= not((inputs(47)) or (inputs(129)));
    layer0_outputs(2305) <= not(inputs(84)) or (inputs(195));
    layer0_outputs(2306) <= inputs(2);
    layer0_outputs(2307) <= (inputs(28)) xor (inputs(82));
    layer0_outputs(2308) <= (inputs(26)) or (inputs(153));
    layer0_outputs(2309) <= not((inputs(150)) xor (inputs(148)));
    layer0_outputs(2310) <= inputs(246);
    layer0_outputs(2311) <= not(inputs(86)) or (inputs(62));
    layer0_outputs(2312) <= not(inputs(223));
    layer0_outputs(2313) <= not(inputs(193));
    layer0_outputs(2314) <= (inputs(157)) or (inputs(179));
    layer0_outputs(2315) <= inputs(108);
    layer0_outputs(2316) <= (inputs(223)) xor (inputs(121));
    layer0_outputs(2317) <= not(inputs(52));
    layer0_outputs(2318) <= inputs(82);
    layer0_outputs(2319) <= not(inputs(183));
    layer0_outputs(2320) <= (inputs(8)) or (inputs(91));
    layer0_outputs(2321) <= (inputs(249)) or (inputs(216));
    layer0_outputs(2322) <= not((inputs(68)) or (inputs(71)));
    layer0_outputs(2323) <= (inputs(242)) xor (inputs(43));
    layer0_outputs(2324) <= not((inputs(222)) or (inputs(79)));
    layer0_outputs(2325) <= not((inputs(247)) or (inputs(106)));
    layer0_outputs(2326) <= not((inputs(197)) xor (inputs(107)));
    layer0_outputs(2327) <= not((inputs(243)) or (inputs(57)));
    layer0_outputs(2328) <= inputs(110);
    layer0_outputs(2329) <= not(inputs(133));
    layer0_outputs(2330) <= '0';
    layer0_outputs(2331) <= (inputs(209)) and (inputs(202));
    layer0_outputs(2332) <= '1';
    layer0_outputs(2333) <= (inputs(174)) or (inputs(186));
    layer0_outputs(2334) <= inputs(79);
    layer0_outputs(2335) <= not(inputs(56)) or (inputs(101));
    layer0_outputs(2336) <= not((inputs(120)) or (inputs(16)));
    layer0_outputs(2337) <= not(inputs(140));
    layer0_outputs(2338) <= (inputs(186)) or (inputs(173));
    layer0_outputs(2339) <= not((inputs(29)) and (inputs(71)));
    layer0_outputs(2340) <= '0';
    layer0_outputs(2341) <= (inputs(204)) and not (inputs(255));
    layer0_outputs(2342) <= (inputs(244)) and not (inputs(96));
    layer0_outputs(2343) <= (inputs(81)) or (inputs(117));
    layer0_outputs(2344) <= not(inputs(198));
    layer0_outputs(2345) <= (inputs(241)) or (inputs(80));
    layer0_outputs(2346) <= (inputs(155)) and (inputs(139));
    layer0_outputs(2347) <= not(inputs(211)) or (inputs(243));
    layer0_outputs(2348) <= not((inputs(30)) and (inputs(111)));
    layer0_outputs(2349) <= not(inputs(146));
    layer0_outputs(2350) <= not(inputs(27)) or (inputs(214));
    layer0_outputs(2351) <= not(inputs(148));
    layer0_outputs(2352) <= inputs(23);
    layer0_outputs(2353) <= (inputs(138)) or (inputs(189));
    layer0_outputs(2354) <= (inputs(246)) and not (inputs(205));
    layer0_outputs(2355) <= not(inputs(89)) or (inputs(15));
    layer0_outputs(2356) <= not(inputs(129)) or (inputs(35));
    layer0_outputs(2357) <= inputs(27);
    layer0_outputs(2358) <= not((inputs(95)) and (inputs(56)));
    layer0_outputs(2359) <= not(inputs(118)) or (inputs(167));
    layer0_outputs(2360) <= not(inputs(233));
    layer0_outputs(2361) <= inputs(95);
    layer0_outputs(2362) <= (inputs(183)) and not (inputs(6));
    layer0_outputs(2363) <= inputs(133);
    layer0_outputs(2364) <= inputs(122);
    layer0_outputs(2365) <= inputs(231);
    layer0_outputs(2366) <= not(inputs(216));
    layer0_outputs(2367) <= not(inputs(231));
    layer0_outputs(2368) <= not(inputs(100)) or (inputs(111));
    layer0_outputs(2369) <= (inputs(233)) or (inputs(159));
    layer0_outputs(2370) <= (inputs(216)) and (inputs(48));
    layer0_outputs(2371) <= not(inputs(172)) or (inputs(249));
    layer0_outputs(2372) <= not(inputs(160));
    layer0_outputs(2373) <= inputs(101);
    layer0_outputs(2374) <= not(inputs(68)) or (inputs(127));
    layer0_outputs(2375) <= (inputs(143)) and not (inputs(6));
    layer0_outputs(2376) <= '1';
    layer0_outputs(2377) <= (inputs(9)) or (inputs(81));
    layer0_outputs(2378) <= (inputs(231)) and not (inputs(120));
    layer0_outputs(2379) <= not(inputs(231));
    layer0_outputs(2380) <= inputs(118);
    layer0_outputs(2381) <= (inputs(118)) and (inputs(159));
    layer0_outputs(2382) <= inputs(179);
    layer0_outputs(2383) <= not((inputs(247)) or (inputs(190)));
    layer0_outputs(2384) <= not(inputs(123)) or (inputs(14));
    layer0_outputs(2385) <= not(inputs(101)) or (inputs(71));
    layer0_outputs(2386) <= inputs(73);
    layer0_outputs(2387) <= not(inputs(213));
    layer0_outputs(2388) <= inputs(153);
    layer0_outputs(2389) <= (inputs(236)) xor (inputs(180));
    layer0_outputs(2390) <= (inputs(239)) or (inputs(106));
    layer0_outputs(2391) <= (inputs(100)) and not (inputs(72));
    layer0_outputs(2392) <= (inputs(181)) and (inputs(216));
    layer0_outputs(2393) <= not(inputs(183));
    layer0_outputs(2394) <= inputs(239);
    layer0_outputs(2395) <= not(inputs(134)) or (inputs(16));
    layer0_outputs(2396) <= (inputs(150)) and not (inputs(62));
    layer0_outputs(2397) <= not((inputs(111)) and (inputs(21)));
    layer0_outputs(2398) <= not(inputs(131));
    layer0_outputs(2399) <= not(inputs(189)) or (inputs(128));
    layer0_outputs(2400) <= (inputs(174)) xor (inputs(238));
    layer0_outputs(2401) <= not((inputs(138)) or (inputs(192)));
    layer0_outputs(2402) <= (inputs(22)) or (inputs(223));
    layer0_outputs(2403) <= not(inputs(73));
    layer0_outputs(2404) <= not((inputs(204)) and (inputs(112)));
    layer0_outputs(2405) <= not(inputs(44)) or (inputs(207));
    layer0_outputs(2406) <= (inputs(184)) or (inputs(167));
    layer0_outputs(2407) <= (inputs(134)) and not (inputs(223));
    layer0_outputs(2408) <= not(inputs(134)) or (inputs(39));
    layer0_outputs(2409) <= not((inputs(170)) xor (inputs(123)));
    layer0_outputs(2410) <= '1';
    layer0_outputs(2411) <= inputs(255);
    layer0_outputs(2412) <= not(inputs(74));
    layer0_outputs(2413) <= (inputs(37)) or (inputs(38));
    layer0_outputs(2414) <= not(inputs(183)) or (inputs(122));
    layer0_outputs(2415) <= (inputs(9)) and not (inputs(20));
    layer0_outputs(2416) <= not((inputs(78)) or (inputs(79)));
    layer0_outputs(2417) <= not(inputs(234));
    layer0_outputs(2418) <= '0';
    layer0_outputs(2419) <= inputs(103);
    layer0_outputs(2420) <= not((inputs(136)) or (inputs(242)));
    layer0_outputs(2421) <= '0';
    layer0_outputs(2422) <= inputs(97);
    layer0_outputs(2423) <= not(inputs(4)) or (inputs(213));
    layer0_outputs(2424) <= not(inputs(116));
    layer0_outputs(2425) <= (inputs(145)) or (inputs(130));
    layer0_outputs(2426) <= not(inputs(177));
    layer0_outputs(2427) <= '0';
    layer0_outputs(2428) <= not(inputs(139));
    layer0_outputs(2429) <= (inputs(224)) or (inputs(144));
    layer0_outputs(2430) <= inputs(104);
    layer0_outputs(2431) <= inputs(17);
    layer0_outputs(2432) <= (inputs(187)) xor (inputs(142));
    layer0_outputs(2433) <= (inputs(113)) and not (inputs(120));
    layer0_outputs(2434) <= not(inputs(194));
    layer0_outputs(2435) <= not(inputs(28)) or (inputs(17));
    layer0_outputs(2436) <= (inputs(112)) xor (inputs(141));
    layer0_outputs(2437) <= not((inputs(197)) and (inputs(53)));
    layer0_outputs(2438) <= inputs(136);
    layer0_outputs(2439) <= (inputs(101)) or (inputs(66));
    layer0_outputs(2440) <= not(inputs(103)) or (inputs(17));
    layer0_outputs(2441) <= '1';
    layer0_outputs(2442) <= '0';
    layer0_outputs(2443) <= not(inputs(232)) or (inputs(7));
    layer0_outputs(2444) <= not(inputs(109));
    layer0_outputs(2445) <= (inputs(6)) or (inputs(60));
    layer0_outputs(2446) <= inputs(228);
    layer0_outputs(2447) <= not((inputs(252)) or (inputs(3)));
    layer0_outputs(2448) <= not(inputs(22)) or (inputs(158));
    layer0_outputs(2449) <= (inputs(12)) or (inputs(197));
    layer0_outputs(2450) <= inputs(141);
    layer0_outputs(2451) <= not(inputs(164));
    layer0_outputs(2452) <= not(inputs(136));
    layer0_outputs(2453) <= not((inputs(115)) or (inputs(192)));
    layer0_outputs(2454) <= not((inputs(222)) xor (inputs(159)));
    layer0_outputs(2455) <= (inputs(114)) and not (inputs(235));
    layer0_outputs(2456) <= not((inputs(114)) or (inputs(181)));
    layer0_outputs(2457) <= not((inputs(180)) or (inputs(56)));
    layer0_outputs(2458) <= not(inputs(183)) or (inputs(121));
    layer0_outputs(2459) <= (inputs(91)) xor (inputs(3));
    layer0_outputs(2460) <= inputs(218);
    layer0_outputs(2461) <= not(inputs(231));
    layer0_outputs(2462) <= (inputs(204)) or (inputs(194));
    layer0_outputs(2463) <= (inputs(89)) and not (inputs(63));
    layer0_outputs(2464) <= (inputs(224)) and (inputs(30));
    layer0_outputs(2465) <= not(inputs(98));
    layer0_outputs(2466) <= not((inputs(145)) or (inputs(202)));
    layer0_outputs(2467) <= inputs(237);
    layer0_outputs(2468) <= (inputs(124)) or (inputs(30));
    layer0_outputs(2469) <= inputs(174);
    layer0_outputs(2470) <= inputs(188);
    layer0_outputs(2471) <= inputs(113);
    layer0_outputs(2472) <= inputs(135);
    layer0_outputs(2473) <= not((inputs(241)) or (inputs(148)));
    layer0_outputs(2474) <= (inputs(16)) or (inputs(1));
    layer0_outputs(2475) <= not(inputs(39));
    layer0_outputs(2476) <= '1';
    layer0_outputs(2477) <= not(inputs(190));
    layer0_outputs(2478) <= (inputs(147)) and (inputs(199));
    layer0_outputs(2479) <= inputs(166);
    layer0_outputs(2480) <= inputs(249);
    layer0_outputs(2481) <= inputs(154);
    layer0_outputs(2482) <= '1';
    layer0_outputs(2483) <= inputs(160);
    layer0_outputs(2484) <= (inputs(49)) or (inputs(33));
    layer0_outputs(2485) <= '0';
    layer0_outputs(2486) <= not((inputs(47)) or (inputs(245)));
    layer0_outputs(2487) <= '0';
    layer0_outputs(2488) <= (inputs(227)) and not (inputs(62));
    layer0_outputs(2489) <= not(inputs(236));
    layer0_outputs(2490) <= inputs(93);
    layer0_outputs(2491) <= not(inputs(222));
    layer0_outputs(2492) <= not(inputs(238));
    layer0_outputs(2493) <= '0';
    layer0_outputs(2494) <= not((inputs(145)) xor (inputs(138)));
    layer0_outputs(2495) <= inputs(8);
    layer0_outputs(2496) <= (inputs(197)) or (inputs(99));
    layer0_outputs(2497) <= not(inputs(31)) or (inputs(46));
    layer0_outputs(2498) <= not(inputs(212));
    layer0_outputs(2499) <= '0';
    layer0_outputs(2500) <= not((inputs(23)) or (inputs(62)));
    layer0_outputs(2501) <= not(inputs(148));
    layer0_outputs(2502) <= (inputs(0)) and not (inputs(15));
    layer0_outputs(2503) <= (inputs(62)) or (inputs(42));
    layer0_outputs(2504) <= (inputs(92)) or (inputs(75));
    layer0_outputs(2505) <= '0';
    layer0_outputs(2506) <= (inputs(20)) or (inputs(202));
    layer0_outputs(2507) <= inputs(242);
    layer0_outputs(2508) <= '0';
    layer0_outputs(2509) <= inputs(125);
    layer0_outputs(2510) <= not(inputs(203));
    layer0_outputs(2511) <= not(inputs(98));
    layer0_outputs(2512) <= (inputs(212)) xor (inputs(224));
    layer0_outputs(2513) <= not(inputs(217)) or (inputs(166));
    layer0_outputs(2514) <= (inputs(196)) and not (inputs(57));
    layer0_outputs(2515) <= inputs(210);
    layer0_outputs(2516) <= (inputs(37)) and not (inputs(236));
    layer0_outputs(2517) <= (inputs(138)) or (inputs(108));
    layer0_outputs(2518) <= (inputs(248)) or (inputs(160));
    layer0_outputs(2519) <= '1';
    layer0_outputs(2520) <= not(inputs(91));
    layer0_outputs(2521) <= (inputs(192)) and not (inputs(214));
    layer0_outputs(2522) <= not(inputs(27)) or (inputs(58));
    layer0_outputs(2523) <= (inputs(4)) xor (inputs(94));
    layer0_outputs(2524) <= '0';
    layer0_outputs(2525) <= (inputs(181)) or (inputs(19));
    layer0_outputs(2526) <= not(inputs(148)) or (inputs(150));
    layer0_outputs(2527) <= not((inputs(157)) or (inputs(126)));
    layer0_outputs(2528) <= not(inputs(249));
    layer0_outputs(2529) <= (inputs(93)) or (inputs(43));
    layer0_outputs(2530) <= '1';
    layer0_outputs(2531) <= not((inputs(55)) or (inputs(23)));
    layer0_outputs(2532) <= not(inputs(175)) or (inputs(15));
    layer0_outputs(2533) <= (inputs(62)) or (inputs(79));
    layer0_outputs(2534) <= inputs(163);
    layer0_outputs(2535) <= not((inputs(66)) xor (inputs(108)));
    layer0_outputs(2536) <= (inputs(246)) and not (inputs(22));
    layer0_outputs(2537) <= inputs(141);
    layer0_outputs(2538) <= not((inputs(169)) or (inputs(88)));
    layer0_outputs(2539) <= not(inputs(211));
    layer0_outputs(2540) <= '0';
    layer0_outputs(2541) <= '0';
    layer0_outputs(2542) <= not(inputs(152));
    layer0_outputs(2543) <= (inputs(222)) xor (inputs(139));
    layer0_outputs(2544) <= '1';
    layer0_outputs(2545) <= inputs(103);
    layer0_outputs(2546) <= not((inputs(177)) or (inputs(88)));
    layer0_outputs(2547) <= not((inputs(45)) or (inputs(120)));
    layer0_outputs(2548) <= not((inputs(67)) or (inputs(175)));
    layer0_outputs(2549) <= inputs(105);
    layer0_outputs(2550) <= (inputs(217)) and not (inputs(75));
    layer0_outputs(2551) <= not(inputs(253));
    layer0_outputs(2552) <= (inputs(136)) and (inputs(219));
    layer0_outputs(2553) <= not(inputs(205));
    layer0_outputs(2554) <= (inputs(41)) and (inputs(37));
    layer0_outputs(2555) <= inputs(57);
    layer0_outputs(2556) <= (inputs(140)) or (inputs(0));
    layer0_outputs(2557) <= not(inputs(75)) or (inputs(254));
    layer0_outputs(2558) <= not((inputs(237)) or (inputs(134)));
    layer0_outputs(2559) <= (inputs(254)) xor (inputs(32));
    layer0_outputs(2560) <= not((inputs(70)) or (inputs(110)));
    layer0_outputs(2561) <= (inputs(24)) and (inputs(238));
    layer0_outputs(2562) <= (inputs(114)) or (inputs(225));
    layer0_outputs(2563) <= inputs(239);
    layer0_outputs(2564) <= (inputs(215)) or (inputs(192));
    layer0_outputs(2565) <= inputs(222);
    layer0_outputs(2566) <= not(inputs(140)) or (inputs(82));
    layer0_outputs(2567) <= inputs(60);
    layer0_outputs(2568) <= (inputs(210)) and not (inputs(23));
    layer0_outputs(2569) <= (inputs(241)) xor (inputs(7));
    layer0_outputs(2570) <= inputs(121);
    layer0_outputs(2571) <= (inputs(170)) and (inputs(178));
    layer0_outputs(2572) <= inputs(162);
    layer0_outputs(2573) <= '1';
    layer0_outputs(2574) <= (inputs(163)) and not (inputs(126));
    layer0_outputs(2575) <= not(inputs(70)) or (inputs(50));
    layer0_outputs(2576) <= (inputs(188)) or (inputs(165));
    layer0_outputs(2577) <= (inputs(210)) xor (inputs(17));
    layer0_outputs(2578) <= (inputs(117)) and not (inputs(180));
    layer0_outputs(2579) <= not((inputs(248)) and (inputs(241)));
    layer0_outputs(2580) <= not(inputs(20));
    layer0_outputs(2581) <= not(inputs(80));
    layer0_outputs(2582) <= not((inputs(47)) or (inputs(160)));
    layer0_outputs(2583) <= inputs(134);
    layer0_outputs(2584) <= inputs(119);
    layer0_outputs(2585) <= not((inputs(156)) xor (inputs(238)));
    layer0_outputs(2586) <= inputs(128);
    layer0_outputs(2587) <= (inputs(160)) and (inputs(65));
    layer0_outputs(2588) <= inputs(81);
    layer0_outputs(2589) <= '0';
    layer0_outputs(2590) <= not(inputs(90));
    layer0_outputs(2591) <= (inputs(21)) and not (inputs(167));
    layer0_outputs(2592) <= not(inputs(137)) or (inputs(8));
    layer0_outputs(2593) <= not(inputs(220));
    layer0_outputs(2594) <= '0';
    layer0_outputs(2595) <= (inputs(240)) and (inputs(51));
    layer0_outputs(2596) <= inputs(90);
    layer0_outputs(2597) <= inputs(217);
    layer0_outputs(2598) <= not((inputs(243)) and (inputs(142)));
    layer0_outputs(2599) <= not(inputs(169)) or (inputs(93));
    layer0_outputs(2600) <= inputs(228);
    layer0_outputs(2601) <= (inputs(81)) and (inputs(24));
    layer0_outputs(2602) <= not((inputs(222)) xor (inputs(69)));
    layer0_outputs(2603) <= not(inputs(214)) or (inputs(227));
    layer0_outputs(2604) <= not((inputs(22)) xor (inputs(26)));
    layer0_outputs(2605) <= (inputs(64)) or (inputs(225));
    layer0_outputs(2606) <= not(inputs(166));
    layer0_outputs(2607) <= not((inputs(207)) xor (inputs(146)));
    layer0_outputs(2608) <= not((inputs(249)) or (inputs(55)));
    layer0_outputs(2609) <= not(inputs(77));
    layer0_outputs(2610) <= not(inputs(100)) or (inputs(48));
    layer0_outputs(2611) <= (inputs(82)) and not (inputs(29));
    layer0_outputs(2612) <= not(inputs(63));
    layer0_outputs(2613) <= '0';
    layer0_outputs(2614) <= (inputs(116)) and not (inputs(254));
    layer0_outputs(2615) <= inputs(137);
    layer0_outputs(2616) <= not((inputs(65)) or (inputs(89)));
    layer0_outputs(2617) <= not(inputs(87));
    layer0_outputs(2618) <= not(inputs(197)) or (inputs(108));
    layer0_outputs(2619) <= not(inputs(244)) or (inputs(15));
    layer0_outputs(2620) <= not((inputs(89)) or (inputs(27)));
    layer0_outputs(2621) <= not((inputs(10)) or (inputs(47)));
    layer0_outputs(2622) <= not(inputs(220));
    layer0_outputs(2623) <= not(inputs(98));
    layer0_outputs(2624) <= (inputs(11)) and not (inputs(234));
    layer0_outputs(2625) <= inputs(157);
    layer0_outputs(2626) <= inputs(43);
    layer0_outputs(2627) <= not(inputs(221));
    layer0_outputs(2628) <= not((inputs(203)) and (inputs(237)));
    layer0_outputs(2629) <= inputs(69);
    layer0_outputs(2630) <= '0';
    layer0_outputs(2631) <= (inputs(142)) and not (inputs(69));
    layer0_outputs(2632) <= not(inputs(130));
    layer0_outputs(2633) <= '1';
    layer0_outputs(2634) <= (inputs(248)) xor (inputs(224));
    layer0_outputs(2635) <= not(inputs(224)) or (inputs(197));
    layer0_outputs(2636) <= not(inputs(182));
    layer0_outputs(2637) <= (inputs(187)) and not (inputs(192));
    layer0_outputs(2638) <= not((inputs(191)) and (inputs(219)));
    layer0_outputs(2639) <= inputs(107);
    layer0_outputs(2640) <= (inputs(176)) and not (inputs(32));
    layer0_outputs(2641) <= (inputs(21)) and not (inputs(82));
    layer0_outputs(2642) <= (inputs(144)) and not (inputs(161));
    layer0_outputs(2643) <= '1';
    layer0_outputs(2644) <= not(inputs(67));
    layer0_outputs(2645) <= (inputs(194)) xor (inputs(150));
    layer0_outputs(2646) <= (inputs(154)) and not (inputs(219));
    layer0_outputs(2647) <= '1';
    layer0_outputs(2648) <= not((inputs(86)) or (inputs(7)));
    layer0_outputs(2649) <= '0';
    layer0_outputs(2650) <= not(inputs(40)) or (inputs(151));
    layer0_outputs(2651) <= (inputs(95)) and (inputs(8));
    layer0_outputs(2652) <= (inputs(122)) and not (inputs(101));
    layer0_outputs(2653) <= (inputs(72)) or (inputs(183));
    layer0_outputs(2654) <= not(inputs(221));
    layer0_outputs(2655) <= (inputs(142)) and (inputs(49));
    layer0_outputs(2656) <= inputs(23);
    layer0_outputs(2657) <= not((inputs(85)) or (inputs(142)));
    layer0_outputs(2658) <= not(inputs(114)) or (inputs(0));
    layer0_outputs(2659) <= not(inputs(80));
    layer0_outputs(2660) <= not((inputs(155)) or (inputs(250)));
    layer0_outputs(2661) <= not(inputs(118));
    layer0_outputs(2662) <= (inputs(43)) or (inputs(61));
    layer0_outputs(2663) <= inputs(123);
    layer0_outputs(2664) <= not((inputs(115)) or (inputs(155)));
    layer0_outputs(2665) <= (inputs(217)) and (inputs(245));
    layer0_outputs(2666) <= (inputs(51)) and not (inputs(126));
    layer0_outputs(2667) <= (inputs(197)) and (inputs(185));
    layer0_outputs(2668) <= not((inputs(119)) or (inputs(87)));
    layer0_outputs(2669) <= inputs(162);
    layer0_outputs(2670) <= (inputs(13)) or (inputs(44));
    layer0_outputs(2671) <= inputs(92);
    layer0_outputs(2672) <= (inputs(40)) and not (inputs(5));
    layer0_outputs(2673) <= not(inputs(156)) or (inputs(223));
    layer0_outputs(2674) <= inputs(146);
    layer0_outputs(2675) <= not(inputs(58));
    layer0_outputs(2676) <= not(inputs(50));
    layer0_outputs(2677) <= not(inputs(70));
    layer0_outputs(2678) <= not(inputs(236));
    layer0_outputs(2679) <= '1';
    layer0_outputs(2680) <= inputs(73);
    layer0_outputs(2681) <= inputs(162);
    layer0_outputs(2682) <= not(inputs(104));
    layer0_outputs(2683) <= not(inputs(195));
    layer0_outputs(2684) <= not(inputs(181));
    layer0_outputs(2685) <= not((inputs(31)) or (inputs(100)));
    layer0_outputs(2686) <= '0';
    layer0_outputs(2687) <= not((inputs(37)) or (inputs(116)));
    layer0_outputs(2688) <= (inputs(243)) xor (inputs(110));
    layer0_outputs(2689) <= not((inputs(44)) or (inputs(249)));
    layer0_outputs(2690) <= '0';
    layer0_outputs(2691) <= (inputs(154)) or (inputs(178));
    layer0_outputs(2692) <= not((inputs(95)) or (inputs(67)));
    layer0_outputs(2693) <= not(inputs(154));
    layer0_outputs(2694) <= (inputs(54)) and not (inputs(16));
    layer0_outputs(2695) <= (inputs(240)) and not (inputs(160));
    layer0_outputs(2696) <= not((inputs(84)) xor (inputs(62)));
    layer0_outputs(2697) <= inputs(49);
    layer0_outputs(2698) <= (inputs(154)) or (inputs(103));
    layer0_outputs(2699) <= not((inputs(178)) or (inputs(204)));
    layer0_outputs(2700) <= (inputs(30)) or (inputs(156));
    layer0_outputs(2701) <= not(inputs(160));
    layer0_outputs(2702) <= '0';
    layer0_outputs(2703) <= not(inputs(108));
    layer0_outputs(2704) <= inputs(136);
    layer0_outputs(2705) <= not(inputs(93));
    layer0_outputs(2706) <= inputs(2);
    layer0_outputs(2707) <= not(inputs(143));
    layer0_outputs(2708) <= not(inputs(51)) or (inputs(112));
    layer0_outputs(2709) <= not(inputs(88));
    layer0_outputs(2710) <= (inputs(166)) and not (inputs(73));
    layer0_outputs(2711) <= inputs(240);
    layer0_outputs(2712) <= inputs(166);
    layer0_outputs(2713) <= not(inputs(57));
    layer0_outputs(2714) <= not((inputs(173)) and (inputs(149)));
    layer0_outputs(2715) <= '0';
    layer0_outputs(2716) <= not((inputs(232)) or (inputs(225)));
    layer0_outputs(2717) <= not(inputs(4));
    layer0_outputs(2718) <= not(inputs(98)) or (inputs(215));
    layer0_outputs(2719) <= not(inputs(81));
    layer0_outputs(2720) <= not(inputs(41));
    layer0_outputs(2721) <= not((inputs(67)) or (inputs(42)));
    layer0_outputs(2722) <= (inputs(19)) or (inputs(207));
    layer0_outputs(2723) <= inputs(206);
    layer0_outputs(2724) <= '0';
    layer0_outputs(2725) <= not(inputs(254)) or (inputs(43));
    layer0_outputs(2726) <= not(inputs(93));
    layer0_outputs(2727) <= '0';
    layer0_outputs(2728) <= not(inputs(124));
    layer0_outputs(2729) <= (inputs(140)) xor (inputs(89));
    layer0_outputs(2730) <= not((inputs(97)) or (inputs(12)));
    layer0_outputs(2731) <= (inputs(1)) and not (inputs(29));
    layer0_outputs(2732) <= (inputs(25)) or (inputs(77));
    layer0_outputs(2733) <= '0';
    layer0_outputs(2734) <= (inputs(193)) or (inputs(194));
    layer0_outputs(2735) <= inputs(141);
    layer0_outputs(2736) <= not(inputs(121)) or (inputs(192));
    layer0_outputs(2737) <= not(inputs(56)) or (inputs(224));
    layer0_outputs(2738) <= (inputs(228)) or (inputs(214));
    layer0_outputs(2739) <= not(inputs(87));
    layer0_outputs(2740) <= not(inputs(140)) or (inputs(225));
    layer0_outputs(2741) <= not(inputs(190));
    layer0_outputs(2742) <= not(inputs(26)) or (inputs(121));
    layer0_outputs(2743) <= (inputs(65)) and not (inputs(128));
    layer0_outputs(2744) <= inputs(24);
    layer0_outputs(2745) <= inputs(1);
    layer0_outputs(2746) <= (inputs(63)) or (inputs(21));
    layer0_outputs(2747) <= not((inputs(73)) and (inputs(123)));
    layer0_outputs(2748) <= (inputs(135)) and not (inputs(248));
    layer0_outputs(2749) <= not(inputs(24));
    layer0_outputs(2750) <= (inputs(208)) or (inputs(69));
    layer0_outputs(2751) <= (inputs(173)) or (inputs(121));
    layer0_outputs(2752) <= (inputs(49)) xor (inputs(95));
    layer0_outputs(2753) <= (inputs(189)) and (inputs(211));
    layer0_outputs(2754) <= inputs(149);
    layer0_outputs(2755) <= inputs(110);
    layer0_outputs(2756) <= (inputs(106)) and not (inputs(186));
    layer0_outputs(2757) <= not(inputs(207));
    layer0_outputs(2758) <= not(inputs(177)) or (inputs(246));
    layer0_outputs(2759) <= (inputs(204)) or (inputs(203));
    layer0_outputs(2760) <= not((inputs(12)) and (inputs(27)));
    layer0_outputs(2761) <= inputs(78);
    layer0_outputs(2762) <= (inputs(150)) and not (inputs(20));
    layer0_outputs(2763) <= (inputs(94)) or (inputs(53));
    layer0_outputs(2764) <= inputs(201);
    layer0_outputs(2765) <= '1';
    layer0_outputs(2766) <= (inputs(173)) or (inputs(94));
    layer0_outputs(2767) <= inputs(47);
    layer0_outputs(2768) <= (inputs(14)) or (inputs(149));
    layer0_outputs(2769) <= (inputs(114)) and (inputs(241));
    layer0_outputs(2770) <= not(inputs(40)) or (inputs(67));
    layer0_outputs(2771) <= not(inputs(26));
    layer0_outputs(2772) <= not((inputs(200)) or (inputs(105)));
    layer0_outputs(2773) <= not(inputs(239));
    layer0_outputs(2774) <= (inputs(116)) and (inputs(151));
    layer0_outputs(2775) <= not((inputs(54)) and (inputs(189)));
    layer0_outputs(2776) <= not((inputs(76)) or (inputs(55)));
    layer0_outputs(2777) <= not(inputs(177));
    layer0_outputs(2778) <= not((inputs(168)) or (inputs(141)));
    layer0_outputs(2779) <= not((inputs(125)) or (inputs(145)));
    layer0_outputs(2780) <= inputs(167);
    layer0_outputs(2781) <= (inputs(190)) and (inputs(143));
    layer0_outputs(2782) <= (inputs(243)) and (inputs(86));
    layer0_outputs(2783) <= not(inputs(116)) or (inputs(126));
    layer0_outputs(2784) <= not((inputs(169)) and (inputs(10)));
    layer0_outputs(2785) <= not((inputs(200)) xor (inputs(197)));
    layer0_outputs(2786) <= inputs(248);
    layer0_outputs(2787) <= inputs(225);
    layer0_outputs(2788) <= not((inputs(149)) xor (inputs(102)));
    layer0_outputs(2789) <= (inputs(197)) or (inputs(255));
    layer0_outputs(2790) <= inputs(28);
    layer0_outputs(2791) <= not(inputs(210));
    layer0_outputs(2792) <= (inputs(184)) or (inputs(43));
    layer0_outputs(2793) <= inputs(72);
    layer0_outputs(2794) <= not((inputs(13)) and (inputs(49)));
    layer0_outputs(2795) <= inputs(213);
    layer0_outputs(2796) <= (inputs(10)) and not (inputs(191));
    layer0_outputs(2797) <= not(inputs(254));
    layer0_outputs(2798) <= inputs(24);
    layer0_outputs(2799) <= not(inputs(140)) or (inputs(168));
    layer0_outputs(2800) <= (inputs(15)) or (inputs(227));
    layer0_outputs(2801) <= (inputs(242)) and not (inputs(253));
    layer0_outputs(2802) <= inputs(194);
    layer0_outputs(2803) <= not((inputs(120)) xor (inputs(255)));
    layer0_outputs(2804) <= (inputs(162)) xor (inputs(180));
    layer0_outputs(2805) <= not((inputs(34)) and (inputs(77)));
    layer0_outputs(2806) <= (inputs(18)) and not (inputs(191));
    layer0_outputs(2807) <= not(inputs(154)) or (inputs(198));
    layer0_outputs(2808) <= not(inputs(238));
    layer0_outputs(2809) <= not(inputs(169));
    layer0_outputs(2810) <= (inputs(26)) and not (inputs(169));
    layer0_outputs(2811) <= (inputs(237)) and not (inputs(200));
    layer0_outputs(2812) <= not(inputs(7)) or (inputs(212));
    layer0_outputs(2813) <= (inputs(239)) or (inputs(25));
    layer0_outputs(2814) <= not(inputs(235));
    layer0_outputs(2815) <= not(inputs(246)) or (inputs(154));
    layer0_outputs(2816) <= '1';
    layer0_outputs(2817) <= (inputs(250)) or (inputs(23));
    layer0_outputs(2818) <= inputs(32);
    layer0_outputs(2819) <= not(inputs(50)) or (inputs(141));
    layer0_outputs(2820) <= inputs(102);
    layer0_outputs(2821) <= not((inputs(112)) and (inputs(124)));
    layer0_outputs(2822) <= '0';
    layer0_outputs(2823) <= not((inputs(135)) or (inputs(58)));
    layer0_outputs(2824) <= (inputs(133)) or (inputs(237));
    layer0_outputs(2825) <= not((inputs(15)) or (inputs(41)));
    layer0_outputs(2826) <= (inputs(214)) and not (inputs(29));
    layer0_outputs(2827) <= not(inputs(230));
    layer0_outputs(2828) <= not(inputs(115));
    layer0_outputs(2829) <= (inputs(132)) and not (inputs(55));
    layer0_outputs(2830) <= not(inputs(179)) or (inputs(17));
    layer0_outputs(2831) <= (inputs(124)) or (inputs(172));
    layer0_outputs(2832) <= not(inputs(35));
    layer0_outputs(2833) <= not(inputs(69));
    layer0_outputs(2834) <= '0';
    layer0_outputs(2835) <= not(inputs(92)) or (inputs(203));
    layer0_outputs(2836) <= not(inputs(102)) or (inputs(2));
    layer0_outputs(2837) <= (inputs(198)) and (inputs(49));
    layer0_outputs(2838) <= not((inputs(175)) or (inputs(106)));
    layer0_outputs(2839) <= (inputs(183)) or (inputs(179));
    layer0_outputs(2840) <= not(inputs(172));
    layer0_outputs(2841) <= (inputs(191)) and not (inputs(212));
    layer0_outputs(2842) <= not((inputs(214)) and (inputs(155)));
    layer0_outputs(2843) <= (inputs(122)) xor (inputs(175));
    layer0_outputs(2844) <= not(inputs(55));
    layer0_outputs(2845) <= (inputs(228)) or (inputs(4));
    layer0_outputs(2846) <= (inputs(82)) and (inputs(90));
    layer0_outputs(2847) <= '0';
    layer0_outputs(2848) <= not(inputs(114));
    layer0_outputs(2849) <= (inputs(3)) and not (inputs(96));
    layer0_outputs(2850) <= (inputs(204)) xor (inputs(176));
    layer0_outputs(2851) <= '1';
    layer0_outputs(2852) <= not(inputs(227)) or (inputs(19));
    layer0_outputs(2853) <= (inputs(216)) xor (inputs(240));
    layer0_outputs(2854) <= inputs(119);
    layer0_outputs(2855) <= not(inputs(161)) or (inputs(168));
    layer0_outputs(2856) <= not((inputs(244)) xor (inputs(60)));
    layer0_outputs(2857) <= '1';
    layer0_outputs(2858) <= not(inputs(215));
    layer0_outputs(2859) <= (inputs(38)) and not (inputs(192));
    layer0_outputs(2860) <= inputs(176);
    layer0_outputs(2861) <= not(inputs(24)) or (inputs(177));
    layer0_outputs(2862) <= not(inputs(230));
    layer0_outputs(2863) <= (inputs(113)) and not (inputs(88));
    layer0_outputs(2864) <= (inputs(145)) or (inputs(228));
    layer0_outputs(2865) <= (inputs(19)) and not (inputs(243));
    layer0_outputs(2866) <= not(inputs(212));
    layer0_outputs(2867) <= (inputs(101)) or (inputs(95));
    layer0_outputs(2868) <= not(inputs(104));
    layer0_outputs(2869) <= not(inputs(117));
    layer0_outputs(2870) <= not(inputs(67));
    layer0_outputs(2871) <= not(inputs(113));
    layer0_outputs(2872) <= (inputs(252)) or (inputs(194));
    layer0_outputs(2873) <= not(inputs(188));
    layer0_outputs(2874) <= (inputs(184)) and (inputs(91));
    layer0_outputs(2875) <= inputs(140);
    layer0_outputs(2876) <= '0';
    layer0_outputs(2877) <= not(inputs(241)) or (inputs(43));
    layer0_outputs(2878) <= not(inputs(219)) or (inputs(129));
    layer0_outputs(2879) <= '1';
    layer0_outputs(2880) <= not(inputs(26));
    layer0_outputs(2881) <= not(inputs(65)) or (inputs(68));
    layer0_outputs(2882) <= not(inputs(221));
    layer0_outputs(2883) <= not((inputs(239)) and (inputs(191)));
    layer0_outputs(2884) <= (inputs(193)) or (inputs(250));
    layer0_outputs(2885) <= not((inputs(180)) or (inputs(50)));
    layer0_outputs(2886) <= not((inputs(195)) or (inputs(230)));
    layer0_outputs(2887) <= not(inputs(139));
    layer0_outputs(2888) <= (inputs(74)) and not (inputs(236));
    layer0_outputs(2889) <= not((inputs(215)) or (inputs(111)));
    layer0_outputs(2890) <= inputs(82);
    layer0_outputs(2891) <= not(inputs(43));
    layer0_outputs(2892) <= (inputs(31)) xor (inputs(50));
    layer0_outputs(2893) <= (inputs(86)) and not (inputs(46));
    layer0_outputs(2894) <= not(inputs(68));
    layer0_outputs(2895) <= '1';
    layer0_outputs(2896) <= not(inputs(157));
    layer0_outputs(2897) <= not(inputs(129));
    layer0_outputs(2898) <= not(inputs(187)) or (inputs(140));
    layer0_outputs(2899) <= not(inputs(44));
    layer0_outputs(2900) <= not(inputs(105));
    layer0_outputs(2901) <= not(inputs(210));
    layer0_outputs(2902) <= '1';
    layer0_outputs(2903) <= (inputs(148)) and not (inputs(57));
    layer0_outputs(2904) <= (inputs(183)) or (inputs(50));
    layer0_outputs(2905) <= not(inputs(5));
    layer0_outputs(2906) <= inputs(130);
    layer0_outputs(2907) <= not(inputs(39));
    layer0_outputs(2908) <= inputs(96);
    layer0_outputs(2909) <= (inputs(27)) or (inputs(101));
    layer0_outputs(2910) <= inputs(138);
    layer0_outputs(2911) <= not((inputs(186)) or (inputs(155)));
    layer0_outputs(2912) <= inputs(210);
    layer0_outputs(2913) <= not((inputs(26)) or (inputs(118)));
    layer0_outputs(2914) <= not(inputs(10)) or (inputs(191));
    layer0_outputs(2915) <= (inputs(171)) or (inputs(177));
    layer0_outputs(2916) <= inputs(15);
    layer0_outputs(2917) <= not((inputs(176)) or (inputs(111)));
    layer0_outputs(2918) <= inputs(148);
    layer0_outputs(2919) <= (inputs(8)) or (inputs(178));
    layer0_outputs(2920) <= not(inputs(196)) or (inputs(64));
    layer0_outputs(2921) <= not((inputs(143)) or (inputs(86)));
    layer0_outputs(2922) <= (inputs(235)) and not (inputs(130));
    layer0_outputs(2923) <= not((inputs(154)) and (inputs(71)));
    layer0_outputs(2924) <= not(inputs(12));
    layer0_outputs(2925) <= not(inputs(194));
    layer0_outputs(2926) <= not((inputs(89)) or (inputs(99)));
    layer0_outputs(2927) <= not((inputs(182)) and (inputs(188)));
    layer0_outputs(2928) <= not((inputs(53)) or (inputs(108)));
    layer0_outputs(2929) <= not(inputs(62));
    layer0_outputs(2930) <= '1';
    layer0_outputs(2931) <= not((inputs(11)) or (inputs(175)));
    layer0_outputs(2932) <= not((inputs(52)) or (inputs(69)));
    layer0_outputs(2933) <= not(inputs(232));
    layer0_outputs(2934) <= '0';
    layer0_outputs(2935) <= (inputs(144)) or (inputs(149));
    layer0_outputs(2936) <= not(inputs(95));
    layer0_outputs(2937) <= not((inputs(18)) or (inputs(238)));
    layer0_outputs(2938) <= not((inputs(186)) or (inputs(138)));
    layer0_outputs(2939) <= (inputs(52)) or (inputs(254));
    layer0_outputs(2940) <= not((inputs(51)) or (inputs(110)));
    layer0_outputs(2941) <= inputs(154);
    layer0_outputs(2942) <= not((inputs(252)) or (inputs(181)));
    layer0_outputs(2943) <= (inputs(252)) or (inputs(233));
    layer0_outputs(2944) <= (inputs(238)) or (inputs(164));
    layer0_outputs(2945) <= (inputs(159)) or (inputs(64));
    layer0_outputs(2946) <= not((inputs(226)) and (inputs(55)));
    layer0_outputs(2947) <= '1';
    layer0_outputs(2948) <= inputs(136);
    layer0_outputs(2949) <= not(inputs(163));
    layer0_outputs(2950) <= not(inputs(228)) or (inputs(117));
    layer0_outputs(2951) <= not((inputs(84)) or (inputs(113)));
    layer0_outputs(2952) <= not((inputs(194)) or (inputs(203)));
    layer0_outputs(2953) <= inputs(142);
    layer0_outputs(2954) <= inputs(153);
    layer0_outputs(2955) <= (inputs(44)) or (inputs(53));
    layer0_outputs(2956) <= not((inputs(157)) and (inputs(188)));
    layer0_outputs(2957) <= inputs(221);
    layer0_outputs(2958) <= not(inputs(113));
    layer0_outputs(2959) <= (inputs(35)) and not (inputs(221));
    layer0_outputs(2960) <= (inputs(190)) and (inputs(34));
    layer0_outputs(2961) <= '1';
    layer0_outputs(2962) <= inputs(101);
    layer0_outputs(2963) <= not((inputs(3)) or (inputs(40)));
    layer0_outputs(2964) <= (inputs(63)) and (inputs(30));
    layer0_outputs(2965) <= not(inputs(213)) or (inputs(96));
    layer0_outputs(2966) <= not(inputs(100));
    layer0_outputs(2967) <= (inputs(80)) or (inputs(43));
    layer0_outputs(2968) <= '1';
    layer0_outputs(2969) <= inputs(234);
    layer0_outputs(2970) <= not(inputs(203)) or (inputs(97));
    layer0_outputs(2971) <= (inputs(178)) xor (inputs(227));
    layer0_outputs(2972) <= not((inputs(248)) or (inputs(129)));
    layer0_outputs(2973) <= '0';
    layer0_outputs(2974) <= inputs(148);
    layer0_outputs(2975) <= not((inputs(228)) or (inputs(215)));
    layer0_outputs(2976) <= not((inputs(191)) and (inputs(50)));
    layer0_outputs(2977) <= inputs(116);
    layer0_outputs(2978) <= not(inputs(215));
    layer0_outputs(2979) <= not((inputs(10)) or (inputs(67)));
    layer0_outputs(2980) <= '1';
    layer0_outputs(2981) <= not((inputs(207)) or (inputs(156)));
    layer0_outputs(2982) <= not(inputs(181)) or (inputs(79));
    layer0_outputs(2983) <= not(inputs(72));
    layer0_outputs(2984) <= '1';
    layer0_outputs(2985) <= not((inputs(74)) or (inputs(115)));
    layer0_outputs(2986) <= not(inputs(143));
    layer0_outputs(2987) <= (inputs(66)) xor (inputs(116));
    layer0_outputs(2988) <= not((inputs(231)) and (inputs(76)));
    layer0_outputs(2989) <= '0';
    layer0_outputs(2990) <= (inputs(33)) or (inputs(245));
    layer0_outputs(2991) <= (inputs(215)) or (inputs(162));
    layer0_outputs(2992) <= not((inputs(99)) xor (inputs(23)));
    layer0_outputs(2993) <= inputs(125);
    layer0_outputs(2994) <= not(inputs(216)) or (inputs(85));
    layer0_outputs(2995) <= (inputs(91)) and not (inputs(159));
    layer0_outputs(2996) <= inputs(187);
    layer0_outputs(2997) <= (inputs(216)) and not (inputs(94));
    layer0_outputs(2998) <= (inputs(119)) and not (inputs(20));
    layer0_outputs(2999) <= '1';
    layer0_outputs(3000) <= not(inputs(83)) or (inputs(133));
    layer0_outputs(3001) <= not((inputs(177)) or (inputs(55)));
    layer0_outputs(3002) <= '0';
    layer0_outputs(3003) <= (inputs(49)) or (inputs(226));
    layer0_outputs(3004) <= (inputs(35)) and not (inputs(232));
    layer0_outputs(3005) <= inputs(124);
    layer0_outputs(3006) <= '1';
    layer0_outputs(3007) <= inputs(111);
    layer0_outputs(3008) <= not(inputs(42)) or (inputs(93));
    layer0_outputs(3009) <= not((inputs(235)) and (inputs(191)));
    layer0_outputs(3010) <= inputs(146);
    layer0_outputs(3011) <= (inputs(197)) or (inputs(70));
    layer0_outputs(3012) <= not((inputs(250)) or (inputs(46)));
    layer0_outputs(3013) <= not((inputs(107)) and (inputs(230)));
    layer0_outputs(3014) <= not((inputs(39)) or (inputs(0)));
    layer0_outputs(3015) <= not((inputs(101)) or (inputs(114)));
    layer0_outputs(3016) <= inputs(122);
    layer0_outputs(3017) <= not(inputs(8));
    layer0_outputs(3018) <= (inputs(0)) or (inputs(34));
    layer0_outputs(3019) <= (inputs(19)) and not (inputs(112));
    layer0_outputs(3020) <= (inputs(100)) and not (inputs(163));
    layer0_outputs(3021) <= not(inputs(107));
    layer0_outputs(3022) <= (inputs(158)) or (inputs(19));
    layer0_outputs(3023) <= '0';
    layer0_outputs(3024) <= (inputs(159)) and not (inputs(93));
    layer0_outputs(3025) <= (inputs(151)) or (inputs(152));
    layer0_outputs(3026) <= inputs(212);
    layer0_outputs(3027) <= not(inputs(234));
    layer0_outputs(3028) <= (inputs(206)) and not (inputs(101));
    layer0_outputs(3029) <= inputs(196);
    layer0_outputs(3030) <= not(inputs(110));
    layer0_outputs(3031) <= (inputs(184)) and (inputs(63));
    layer0_outputs(3032) <= not(inputs(74));
    layer0_outputs(3033) <= not(inputs(246));
    layer0_outputs(3034) <= not((inputs(126)) and (inputs(117)));
    layer0_outputs(3035) <= not(inputs(69));
    layer0_outputs(3036) <= (inputs(57)) or (inputs(67));
    layer0_outputs(3037) <= (inputs(48)) or (inputs(35));
    layer0_outputs(3038) <= not((inputs(85)) xor (inputs(96)));
    layer0_outputs(3039) <= not(inputs(139)) or (inputs(208));
    layer0_outputs(3040) <= not((inputs(195)) or (inputs(162)));
    layer0_outputs(3041) <= not(inputs(102)) or (inputs(199));
    layer0_outputs(3042) <= not(inputs(176));
    layer0_outputs(3043) <= '1';
    layer0_outputs(3044) <= not(inputs(125)) or (inputs(20));
    layer0_outputs(3045) <= (inputs(47)) or (inputs(78));
    layer0_outputs(3046) <= (inputs(233)) and not (inputs(4));
    layer0_outputs(3047) <= not(inputs(179)) or (inputs(242));
    layer0_outputs(3048) <= not((inputs(107)) xor (inputs(142)));
    layer0_outputs(3049) <= inputs(100);
    layer0_outputs(3050) <= (inputs(17)) or (inputs(218));
    layer0_outputs(3051) <= '1';
    layer0_outputs(3052) <= (inputs(122)) and (inputs(60));
    layer0_outputs(3053) <= not(inputs(179));
    layer0_outputs(3054) <= not(inputs(244)) or (inputs(172));
    layer0_outputs(3055) <= (inputs(71)) or (inputs(201));
    layer0_outputs(3056) <= inputs(183);
    layer0_outputs(3057) <= not(inputs(244));
    layer0_outputs(3058) <= not((inputs(190)) and (inputs(188)));
    layer0_outputs(3059) <= not(inputs(148));
    layer0_outputs(3060) <= '1';
    layer0_outputs(3061) <= (inputs(79)) or (inputs(172));
    layer0_outputs(3062) <= (inputs(173)) and not (inputs(30));
    layer0_outputs(3063) <= not(inputs(191)) or (inputs(162));
    layer0_outputs(3064) <= not(inputs(24));
    layer0_outputs(3065) <= not(inputs(209));
    layer0_outputs(3066) <= (inputs(66)) and (inputs(189));
    layer0_outputs(3067) <= (inputs(89)) and not (inputs(112));
    layer0_outputs(3068) <= not((inputs(230)) or (inputs(27)));
    layer0_outputs(3069) <= (inputs(100)) and not (inputs(3));
    layer0_outputs(3070) <= not(inputs(206));
    layer0_outputs(3071) <= inputs(167);
    layer0_outputs(3072) <= (inputs(250)) and (inputs(45));
    layer0_outputs(3073) <= inputs(51);
    layer0_outputs(3074) <= not(inputs(54));
    layer0_outputs(3075) <= not(inputs(241));
    layer0_outputs(3076) <= inputs(126);
    layer0_outputs(3077) <= (inputs(146)) or (inputs(163));
    layer0_outputs(3078) <= not(inputs(57)) or (inputs(13));
    layer0_outputs(3079) <= not((inputs(219)) or (inputs(196)));
    layer0_outputs(3080) <= not((inputs(20)) or (inputs(244)));
    layer0_outputs(3081) <= not(inputs(104)) or (inputs(201));
    layer0_outputs(3082) <= (inputs(24)) and not (inputs(175));
    layer0_outputs(3083) <= (inputs(156)) and not (inputs(198));
    layer0_outputs(3084) <= (inputs(249)) and (inputs(222));
    layer0_outputs(3085) <= not((inputs(56)) or (inputs(1)));
    layer0_outputs(3086) <= '1';
    layer0_outputs(3087) <= not(inputs(237));
    layer0_outputs(3088) <= not(inputs(33));
    layer0_outputs(3089) <= (inputs(169)) or (inputs(60));
    layer0_outputs(3090) <= (inputs(6)) or (inputs(93));
    layer0_outputs(3091) <= not(inputs(181));
    layer0_outputs(3092) <= not(inputs(149)) or (inputs(95));
    layer0_outputs(3093) <= not(inputs(215)) or (inputs(10));
    layer0_outputs(3094) <= (inputs(88)) and not (inputs(250));
    layer0_outputs(3095) <= not(inputs(1));
    layer0_outputs(3096) <= inputs(165);
    layer0_outputs(3097) <= inputs(139);
    layer0_outputs(3098) <= (inputs(28)) xor (inputs(255));
    layer0_outputs(3099) <= (inputs(35)) or (inputs(183));
    layer0_outputs(3100) <= inputs(166);
    layer0_outputs(3101) <= not(inputs(93));
    layer0_outputs(3102) <= not(inputs(174));
    layer0_outputs(3103) <= '0';
    layer0_outputs(3104) <= (inputs(87)) and not (inputs(201));
    layer0_outputs(3105) <= (inputs(163)) and not (inputs(127));
    layer0_outputs(3106) <= not((inputs(109)) or (inputs(74)));
    layer0_outputs(3107) <= not((inputs(3)) or (inputs(137)));
    layer0_outputs(3108) <= not((inputs(44)) or (inputs(186)));
    layer0_outputs(3109) <= not(inputs(94)) or (inputs(185));
    layer0_outputs(3110) <= not(inputs(218));
    layer0_outputs(3111) <= not((inputs(185)) xor (inputs(137)));
    layer0_outputs(3112) <= inputs(208);
    layer0_outputs(3113) <= not(inputs(105));
    layer0_outputs(3114) <= inputs(125);
    layer0_outputs(3115) <= inputs(128);
    layer0_outputs(3116) <= not(inputs(132)) or (inputs(175));
    layer0_outputs(3117) <= not(inputs(211)) or (inputs(94));
    layer0_outputs(3118) <= (inputs(72)) or (inputs(243));
    layer0_outputs(3119) <= not(inputs(177));
    layer0_outputs(3120) <= not(inputs(45));
    layer0_outputs(3121) <= not(inputs(132)) or (inputs(49));
    layer0_outputs(3122) <= (inputs(36)) and not (inputs(155));
    layer0_outputs(3123) <= (inputs(221)) and not (inputs(57));
    layer0_outputs(3124) <= not((inputs(141)) or (inputs(232)));
    layer0_outputs(3125) <= (inputs(219)) and (inputs(252));
    layer0_outputs(3126) <= (inputs(231)) and not (inputs(98));
    layer0_outputs(3127) <= not((inputs(176)) and (inputs(189)));
    layer0_outputs(3128) <= inputs(87);
    layer0_outputs(3129) <= inputs(168);
    layer0_outputs(3130) <= inputs(197);
    layer0_outputs(3131) <= not((inputs(22)) or (inputs(245)));
    layer0_outputs(3132) <= (inputs(72)) and not (inputs(163));
    layer0_outputs(3133) <= (inputs(61)) or (inputs(1));
    layer0_outputs(3134) <= not((inputs(21)) or (inputs(55)));
    layer0_outputs(3135) <= inputs(52);
    layer0_outputs(3136) <= (inputs(22)) or (inputs(64));
    layer0_outputs(3137) <= not(inputs(108)) or (inputs(160));
    layer0_outputs(3138) <= not((inputs(23)) or (inputs(96)));
    layer0_outputs(3139) <= (inputs(25)) and not (inputs(222));
    layer0_outputs(3140) <= not(inputs(34)) or (inputs(236));
    layer0_outputs(3141) <= not(inputs(178));
    layer0_outputs(3142) <= inputs(53);
    layer0_outputs(3143) <= not(inputs(78));
    layer0_outputs(3144) <= not(inputs(213));
    layer0_outputs(3145) <= (inputs(66)) and not (inputs(91));
    layer0_outputs(3146) <= not((inputs(212)) or (inputs(151)));
    layer0_outputs(3147) <= (inputs(131)) or (inputs(132));
    layer0_outputs(3148) <= '0';
    layer0_outputs(3149) <= not(inputs(119)) or (inputs(12));
    layer0_outputs(3150) <= not(inputs(128));
    layer0_outputs(3151) <= inputs(216);
    layer0_outputs(3152) <= not((inputs(163)) or (inputs(149)));
    layer0_outputs(3153) <= (inputs(121)) and not (inputs(163));
    layer0_outputs(3154) <= (inputs(183)) and not (inputs(16));
    layer0_outputs(3155) <= not(inputs(96));
    layer0_outputs(3156) <= inputs(152);
    layer0_outputs(3157) <= not((inputs(211)) or (inputs(101)));
    layer0_outputs(3158) <= not((inputs(79)) or (inputs(200)));
    layer0_outputs(3159) <= (inputs(11)) and not (inputs(65));
    layer0_outputs(3160) <= not(inputs(247)) or (inputs(223));
    layer0_outputs(3161) <= (inputs(204)) or (inputs(227));
    layer0_outputs(3162) <= (inputs(249)) and not (inputs(15));
    layer0_outputs(3163) <= not((inputs(37)) or (inputs(236)));
    layer0_outputs(3164) <= inputs(210);
    layer0_outputs(3165) <= '0';
    layer0_outputs(3166) <= '1';
    layer0_outputs(3167) <= not((inputs(38)) or (inputs(87)));
    layer0_outputs(3168) <= inputs(196);
    layer0_outputs(3169) <= not(inputs(204));
    layer0_outputs(3170) <= (inputs(218)) or (inputs(108));
    layer0_outputs(3171) <= not((inputs(145)) or (inputs(204)));
    layer0_outputs(3172) <= not(inputs(196)) or (inputs(90));
    layer0_outputs(3173) <= not(inputs(186)) or (inputs(111));
    layer0_outputs(3174) <= '0';
    layer0_outputs(3175) <= not((inputs(229)) or (inputs(240)));
    layer0_outputs(3176) <= (inputs(145)) xor (inputs(171));
    layer0_outputs(3177) <= (inputs(192)) xor (inputs(39));
    layer0_outputs(3178) <= inputs(106);
    layer0_outputs(3179) <= not(inputs(255));
    layer0_outputs(3180) <= not((inputs(89)) or (inputs(60)));
    layer0_outputs(3181) <= inputs(116);
    layer0_outputs(3182) <= '0';
    layer0_outputs(3183) <= not((inputs(120)) or (inputs(117)));
    layer0_outputs(3184) <= inputs(88);
    layer0_outputs(3185) <= not(inputs(51));
    layer0_outputs(3186) <= inputs(195);
    layer0_outputs(3187) <= (inputs(122)) and not (inputs(167));
    layer0_outputs(3188) <= inputs(9);
    layer0_outputs(3189) <= '0';
    layer0_outputs(3190) <= (inputs(183)) or (inputs(49));
    layer0_outputs(3191) <= not(inputs(78));
    layer0_outputs(3192) <= '1';
    layer0_outputs(3193) <= inputs(58);
    layer0_outputs(3194) <= '0';
    layer0_outputs(3195) <= (inputs(213)) or (inputs(175));
    layer0_outputs(3196) <= not(inputs(203));
    layer0_outputs(3197) <= not(inputs(181));
    layer0_outputs(3198) <= not(inputs(178)) or (inputs(16));
    layer0_outputs(3199) <= (inputs(127)) or (inputs(124));
    layer0_outputs(3200) <= not(inputs(232)) or (inputs(103));
    layer0_outputs(3201) <= not((inputs(43)) and (inputs(231)));
    layer0_outputs(3202) <= (inputs(37)) xor (inputs(219));
    layer0_outputs(3203) <= not(inputs(79));
    layer0_outputs(3204) <= not((inputs(54)) and (inputs(248)));
    layer0_outputs(3205) <= not(inputs(98));
    layer0_outputs(3206) <= not((inputs(219)) or (inputs(121)));
    layer0_outputs(3207) <= (inputs(220)) and not (inputs(125));
    layer0_outputs(3208) <= not(inputs(13)) or (inputs(121));
    layer0_outputs(3209) <= inputs(135);
    layer0_outputs(3210) <= not(inputs(146));
    layer0_outputs(3211) <= inputs(98);
    layer0_outputs(3212) <= (inputs(235)) or (inputs(28));
    layer0_outputs(3213) <= not(inputs(149));
    layer0_outputs(3214) <= not((inputs(37)) or (inputs(145)));
    layer0_outputs(3215) <= not(inputs(101));
    layer0_outputs(3216) <= not(inputs(235)) or (inputs(37));
    layer0_outputs(3217) <= (inputs(182)) and not (inputs(141));
    layer0_outputs(3218) <= inputs(89);
    layer0_outputs(3219) <= inputs(72);
    layer0_outputs(3220) <= inputs(9);
    layer0_outputs(3221) <= (inputs(126)) and not (inputs(157));
    layer0_outputs(3222) <= not((inputs(111)) or (inputs(204)));
    layer0_outputs(3223) <= not(inputs(174));
    layer0_outputs(3224) <= '1';
    layer0_outputs(3225) <= (inputs(118)) xor (inputs(205));
    layer0_outputs(3226) <= inputs(130);
    layer0_outputs(3227) <= not(inputs(133)) or (inputs(144));
    layer0_outputs(3228) <= not(inputs(247)) or (inputs(110));
    layer0_outputs(3229) <= inputs(124);
    layer0_outputs(3230) <= (inputs(154)) and (inputs(153));
    layer0_outputs(3231) <= not(inputs(185));
    layer0_outputs(3232) <= inputs(35);
    layer0_outputs(3233) <= inputs(205);
    layer0_outputs(3234) <= (inputs(111)) and not (inputs(72));
    layer0_outputs(3235) <= (inputs(12)) xor (inputs(219));
    layer0_outputs(3236) <= (inputs(143)) or (inputs(127));
    layer0_outputs(3237) <= not((inputs(55)) and (inputs(214)));
    layer0_outputs(3238) <= not((inputs(233)) and (inputs(43)));
    layer0_outputs(3239) <= inputs(48);
    layer0_outputs(3240) <= not((inputs(255)) or (inputs(33)));
    layer0_outputs(3241) <= (inputs(212)) and (inputs(253));
    layer0_outputs(3242) <= not((inputs(176)) or (inputs(171)));
    layer0_outputs(3243) <= '1';
    layer0_outputs(3244) <= not(inputs(105));
    layer0_outputs(3245) <= inputs(142);
    layer0_outputs(3246) <= inputs(195);
    layer0_outputs(3247) <= (inputs(54)) and not (inputs(70));
    layer0_outputs(3248) <= not(inputs(3));
    layer0_outputs(3249) <= '1';
    layer0_outputs(3250) <= '0';
    layer0_outputs(3251) <= inputs(241);
    layer0_outputs(3252) <= (inputs(204)) or (inputs(20));
    layer0_outputs(3253) <= not(inputs(138)) or (inputs(15));
    layer0_outputs(3254) <= (inputs(182)) or (inputs(113));
    layer0_outputs(3255) <= '1';
    layer0_outputs(3256) <= not((inputs(211)) or (inputs(43)));
    layer0_outputs(3257) <= (inputs(238)) or (inputs(59));
    layer0_outputs(3258) <= not((inputs(39)) xor (inputs(71)));
    layer0_outputs(3259) <= inputs(178);
    layer0_outputs(3260) <= not((inputs(55)) or (inputs(86)));
    layer0_outputs(3261) <= '1';
    layer0_outputs(3262) <= not((inputs(112)) or (inputs(26)));
    layer0_outputs(3263) <= not((inputs(249)) and (inputs(168)));
    layer0_outputs(3264) <= (inputs(32)) and not (inputs(230));
    layer0_outputs(3265) <= not(inputs(117));
    layer0_outputs(3266) <= (inputs(56)) and not (inputs(38));
    layer0_outputs(3267) <= (inputs(98)) xor (inputs(51));
    layer0_outputs(3268) <= not((inputs(252)) xor (inputs(125)));
    layer0_outputs(3269) <= (inputs(147)) xor (inputs(3));
    layer0_outputs(3270) <= not(inputs(116));
    layer0_outputs(3271) <= (inputs(137)) and not (inputs(191));
    layer0_outputs(3272) <= (inputs(118)) and not (inputs(253));
    layer0_outputs(3273) <= not((inputs(240)) xor (inputs(93)));
    layer0_outputs(3274) <= not(inputs(127));
    layer0_outputs(3275) <= not((inputs(166)) or (inputs(47)));
    layer0_outputs(3276) <= '1';
    layer0_outputs(3277) <= inputs(64);
    layer0_outputs(3278) <= not((inputs(12)) or (inputs(96)));
    layer0_outputs(3279) <= (inputs(252)) or (inputs(255));
    layer0_outputs(3280) <= (inputs(169)) and not (inputs(53));
    layer0_outputs(3281) <= not(inputs(86));
    layer0_outputs(3282) <= '1';
    layer0_outputs(3283) <= '0';
    layer0_outputs(3284) <= not(inputs(193)) or (inputs(112));
    layer0_outputs(3285) <= '1';
    layer0_outputs(3286) <= not((inputs(237)) xor (inputs(164)));
    layer0_outputs(3287) <= not(inputs(27)) or (inputs(104));
    layer0_outputs(3288) <= not(inputs(131));
    layer0_outputs(3289) <= not(inputs(192));
    layer0_outputs(3290) <= '1';
    layer0_outputs(3291) <= inputs(130);
    layer0_outputs(3292) <= not((inputs(160)) or (inputs(130)));
    layer0_outputs(3293) <= (inputs(218)) or (inputs(123));
    layer0_outputs(3294) <= inputs(218);
    layer0_outputs(3295) <= inputs(53);
    layer0_outputs(3296) <= not((inputs(188)) or (inputs(67)));
    layer0_outputs(3297) <= inputs(69);
    layer0_outputs(3298) <= (inputs(152)) xor (inputs(135));
    layer0_outputs(3299) <= not((inputs(55)) and (inputs(2)));
    layer0_outputs(3300) <= not(inputs(105));
    layer0_outputs(3301) <= not(inputs(150));
    layer0_outputs(3302) <= (inputs(9)) or (inputs(94));
    layer0_outputs(3303) <= inputs(250);
    layer0_outputs(3304) <= (inputs(250)) or (inputs(204));
    layer0_outputs(3305) <= '0';
    layer0_outputs(3306) <= (inputs(228)) and not (inputs(14));
    layer0_outputs(3307) <= not(inputs(133)) or (inputs(0));
    layer0_outputs(3308) <= not(inputs(178));
    layer0_outputs(3309) <= (inputs(159)) and not (inputs(17));
    layer0_outputs(3310) <= not((inputs(55)) xor (inputs(119)));
    layer0_outputs(3311) <= not(inputs(131)) or (inputs(17));
    layer0_outputs(3312) <= not((inputs(68)) and (inputs(42)));
    layer0_outputs(3313) <= (inputs(229)) and (inputs(117));
    layer0_outputs(3314) <= not(inputs(187));
    layer0_outputs(3315) <= not(inputs(238));
    layer0_outputs(3316) <= '0';
    layer0_outputs(3317) <= '1';
    layer0_outputs(3318) <= not(inputs(172));
    layer0_outputs(3319) <= inputs(124);
    layer0_outputs(3320) <= inputs(250);
    layer0_outputs(3321) <= '0';
    layer0_outputs(3322) <= (inputs(138)) and not (inputs(185));
    layer0_outputs(3323) <= inputs(190);
    layer0_outputs(3324) <= inputs(243);
    layer0_outputs(3325) <= inputs(201);
    layer0_outputs(3326) <= not((inputs(110)) or (inputs(144)));
    layer0_outputs(3327) <= not((inputs(183)) or (inputs(136)));
    layer0_outputs(3328) <= (inputs(248)) or (inputs(54));
    layer0_outputs(3329) <= not(inputs(41)) or (inputs(72));
    layer0_outputs(3330) <= not(inputs(123)) or (inputs(180));
    layer0_outputs(3331) <= not(inputs(209));
    layer0_outputs(3332) <= (inputs(93)) and (inputs(87));
    layer0_outputs(3333) <= not((inputs(235)) and (inputs(86)));
    layer0_outputs(3334) <= not((inputs(114)) and (inputs(249)));
    layer0_outputs(3335) <= not(inputs(82));
    layer0_outputs(3336) <= not((inputs(179)) or (inputs(145)));
    layer0_outputs(3337) <= inputs(133);
    layer0_outputs(3338) <= not(inputs(158));
    layer0_outputs(3339) <= not(inputs(38));
    layer0_outputs(3340) <= inputs(108);
    layer0_outputs(3341) <= not(inputs(17));
    layer0_outputs(3342) <= (inputs(97)) and (inputs(255));
    layer0_outputs(3343) <= not((inputs(195)) or (inputs(229)));
    layer0_outputs(3344) <= (inputs(7)) xor (inputs(97));
    layer0_outputs(3345) <= (inputs(74)) and (inputs(185));
    layer0_outputs(3346) <= not(inputs(81));
    layer0_outputs(3347) <= (inputs(239)) and not (inputs(226));
    layer0_outputs(3348) <= not(inputs(162));
    layer0_outputs(3349) <= not(inputs(45));
    layer0_outputs(3350) <= '0';
    layer0_outputs(3351) <= (inputs(116)) and (inputs(179));
    layer0_outputs(3352) <= (inputs(24)) and (inputs(121));
    layer0_outputs(3353) <= not(inputs(125));
    layer0_outputs(3354) <= (inputs(167)) xor (inputs(72));
    layer0_outputs(3355) <= (inputs(94)) and not (inputs(91));
    layer0_outputs(3356) <= inputs(48);
    layer0_outputs(3357) <= (inputs(202)) xor (inputs(220));
    layer0_outputs(3358) <= not(inputs(145));
    layer0_outputs(3359) <= inputs(77);
    layer0_outputs(3360) <= inputs(68);
    layer0_outputs(3361) <= not((inputs(118)) xor (inputs(222)));
    layer0_outputs(3362) <= (inputs(108)) xor (inputs(98));
    layer0_outputs(3363) <= not(inputs(175)) or (inputs(192));
    layer0_outputs(3364) <= not(inputs(87));
    layer0_outputs(3365) <= '1';
    layer0_outputs(3366) <= not(inputs(29));
    layer0_outputs(3367) <= (inputs(172)) and (inputs(250));
    layer0_outputs(3368) <= inputs(144);
    layer0_outputs(3369) <= (inputs(1)) xor (inputs(188));
    layer0_outputs(3370) <= not((inputs(69)) or (inputs(180)));
    layer0_outputs(3371) <= (inputs(26)) xor (inputs(203));
    layer0_outputs(3372) <= (inputs(36)) and not (inputs(157));
    layer0_outputs(3373) <= (inputs(189)) or (inputs(224));
    layer0_outputs(3374) <= not((inputs(7)) and (inputs(7)));
    layer0_outputs(3375) <= (inputs(237)) and (inputs(191));
    layer0_outputs(3376) <= not(inputs(115));
    layer0_outputs(3377) <= not(inputs(96));
    layer0_outputs(3378) <= inputs(236);
    layer0_outputs(3379) <= not(inputs(112)) or (inputs(241));
    layer0_outputs(3380) <= not((inputs(30)) or (inputs(30)));
    layer0_outputs(3381) <= not(inputs(8));
    layer0_outputs(3382) <= (inputs(66)) xor (inputs(186));
    layer0_outputs(3383) <= inputs(228);
    layer0_outputs(3384) <= (inputs(150)) and not (inputs(156));
    layer0_outputs(3385) <= (inputs(122)) or (inputs(73));
    layer0_outputs(3386) <= not(inputs(24));
    layer0_outputs(3387) <= not(inputs(39));
    layer0_outputs(3388) <= not((inputs(139)) and (inputs(245)));
    layer0_outputs(3389) <= not(inputs(126));
    layer0_outputs(3390) <= (inputs(81)) or (inputs(100));
    layer0_outputs(3391) <= not(inputs(50));
    layer0_outputs(3392) <= not(inputs(22));
    layer0_outputs(3393) <= not(inputs(191));
    layer0_outputs(3394) <= (inputs(110)) and (inputs(235));
    layer0_outputs(3395) <= inputs(120);
    layer0_outputs(3396) <= (inputs(10)) xor (inputs(75));
    layer0_outputs(3397) <= not((inputs(113)) or (inputs(132)));
    layer0_outputs(3398) <= inputs(116);
    layer0_outputs(3399) <= not(inputs(101)) or (inputs(172));
    layer0_outputs(3400) <= (inputs(198)) and (inputs(155));
    layer0_outputs(3401) <= (inputs(217)) or (inputs(255));
    layer0_outputs(3402) <= not((inputs(53)) xor (inputs(34)));
    layer0_outputs(3403) <= (inputs(95)) xor (inputs(33));
    layer0_outputs(3404) <= not(inputs(78)) or (inputs(92));
    layer0_outputs(3405) <= (inputs(172)) or (inputs(123));
    layer0_outputs(3406) <= not(inputs(46)) or (inputs(5));
    layer0_outputs(3407) <= not((inputs(249)) and (inputs(224)));
    layer0_outputs(3408) <= not(inputs(204));
    layer0_outputs(3409) <= inputs(228);
    layer0_outputs(3410) <= inputs(129);
    layer0_outputs(3411) <= not(inputs(200));
    layer0_outputs(3412) <= (inputs(82)) or (inputs(42));
    layer0_outputs(3413) <= not((inputs(132)) or (inputs(221)));
    layer0_outputs(3414) <= (inputs(162)) or (inputs(255));
    layer0_outputs(3415) <= (inputs(251)) xor (inputs(220));
    layer0_outputs(3416) <= not(inputs(116));
    layer0_outputs(3417) <= (inputs(140)) xor (inputs(67));
    layer0_outputs(3418) <= inputs(219);
    layer0_outputs(3419) <= inputs(1);
    layer0_outputs(3420) <= (inputs(156)) or (inputs(219));
    layer0_outputs(3421) <= (inputs(18)) xor (inputs(154));
    layer0_outputs(3422) <= not(inputs(233)) or (inputs(89));
    layer0_outputs(3423) <= '0';
    layer0_outputs(3424) <= not((inputs(22)) or (inputs(224)));
    layer0_outputs(3425) <= (inputs(219)) and not (inputs(143));
    layer0_outputs(3426) <= inputs(72);
    layer0_outputs(3427) <= inputs(254);
    layer0_outputs(3428) <= not(inputs(113));
    layer0_outputs(3429) <= (inputs(91)) or (inputs(185));
    layer0_outputs(3430) <= not((inputs(130)) or (inputs(4)));
    layer0_outputs(3431) <= not(inputs(202));
    layer0_outputs(3432) <= (inputs(26)) or (inputs(80));
    layer0_outputs(3433) <= (inputs(186)) or (inputs(162));
    layer0_outputs(3434) <= '1';
    layer0_outputs(3435) <= '0';
    layer0_outputs(3436) <= '0';
    layer0_outputs(3437) <= inputs(74);
    layer0_outputs(3438) <= inputs(217);
    layer0_outputs(3439) <= (inputs(11)) or (inputs(81));
    layer0_outputs(3440) <= not((inputs(101)) xor (inputs(96)));
    layer0_outputs(3441) <= (inputs(27)) and not (inputs(121));
    layer0_outputs(3442) <= not(inputs(3)) or (inputs(159));
    layer0_outputs(3443) <= not((inputs(252)) and (inputs(190)));
    layer0_outputs(3444) <= (inputs(212)) and not (inputs(102));
    layer0_outputs(3445) <= (inputs(46)) and (inputs(250));
    layer0_outputs(3446) <= '1';
    layer0_outputs(3447) <= (inputs(125)) or (inputs(126));
    layer0_outputs(3448) <= not(inputs(99));
    layer0_outputs(3449) <= (inputs(131)) and not (inputs(19));
    layer0_outputs(3450) <= not((inputs(107)) or (inputs(51)));
    layer0_outputs(3451) <= not(inputs(185));
    layer0_outputs(3452) <= inputs(245);
    layer0_outputs(3453) <= not(inputs(59)) or (inputs(134));
    layer0_outputs(3454) <= (inputs(115)) and not (inputs(0));
    layer0_outputs(3455) <= '0';
    layer0_outputs(3456) <= (inputs(8)) and not (inputs(112));
    layer0_outputs(3457) <= (inputs(111)) and (inputs(143));
    layer0_outputs(3458) <= not(inputs(109));
    layer0_outputs(3459) <= not(inputs(251));
    layer0_outputs(3460) <= not((inputs(87)) xor (inputs(115)));
    layer0_outputs(3461) <= not((inputs(127)) and (inputs(96)));
    layer0_outputs(3462) <= not((inputs(51)) xor (inputs(103)));
    layer0_outputs(3463) <= (inputs(174)) and not (inputs(42));
    layer0_outputs(3464) <= (inputs(122)) or (inputs(137));
    layer0_outputs(3465) <= not(inputs(163)) or (inputs(238));
    layer0_outputs(3466) <= '1';
    layer0_outputs(3467) <= '0';
    layer0_outputs(3468) <= not(inputs(66));
    layer0_outputs(3469) <= (inputs(195)) and not (inputs(102));
    layer0_outputs(3470) <= (inputs(165)) and not (inputs(51));
    layer0_outputs(3471) <= not((inputs(11)) or (inputs(159)));
    layer0_outputs(3472) <= (inputs(211)) or (inputs(138));
    layer0_outputs(3473) <= inputs(77);
    layer0_outputs(3474) <= not(inputs(137));
    layer0_outputs(3475) <= inputs(44);
    layer0_outputs(3476) <= not((inputs(233)) and (inputs(148)));
    layer0_outputs(3477) <= (inputs(79)) xor (inputs(74));
    layer0_outputs(3478) <= not((inputs(111)) or (inputs(174)));
    layer0_outputs(3479) <= (inputs(42)) or (inputs(162));
    layer0_outputs(3480) <= not((inputs(147)) xor (inputs(136)));
    layer0_outputs(3481) <= (inputs(22)) or (inputs(68));
    layer0_outputs(3482) <= inputs(172);
    layer0_outputs(3483) <= not((inputs(116)) and (inputs(246)));
    layer0_outputs(3484) <= not((inputs(179)) or (inputs(146)));
    layer0_outputs(3485) <= not(inputs(120));
    layer0_outputs(3486) <= inputs(84);
    layer0_outputs(3487) <= not((inputs(38)) or (inputs(67)));
    layer0_outputs(3488) <= (inputs(67)) and (inputs(71));
    layer0_outputs(3489) <= (inputs(250)) and (inputs(248));
    layer0_outputs(3490) <= inputs(164);
    layer0_outputs(3491) <= inputs(143);
    layer0_outputs(3492) <= (inputs(38)) and not (inputs(179));
    layer0_outputs(3493) <= inputs(255);
    layer0_outputs(3494) <= inputs(90);
    layer0_outputs(3495) <= not(inputs(233));
    layer0_outputs(3496) <= inputs(155);
    layer0_outputs(3497) <= not(inputs(248));
    layer0_outputs(3498) <= (inputs(131)) and not (inputs(17));
    layer0_outputs(3499) <= not((inputs(251)) or (inputs(236)));
    layer0_outputs(3500) <= not(inputs(93));
    layer0_outputs(3501) <= not(inputs(48));
    layer0_outputs(3502) <= '1';
    layer0_outputs(3503) <= '1';
    layer0_outputs(3504) <= '0';
    layer0_outputs(3505) <= inputs(161);
    layer0_outputs(3506) <= not(inputs(218)) or (inputs(71));
    layer0_outputs(3507) <= inputs(232);
    layer0_outputs(3508) <= (inputs(246)) and (inputs(233));
    layer0_outputs(3509) <= inputs(212);
    layer0_outputs(3510) <= not(inputs(39)) or (inputs(94));
    layer0_outputs(3511) <= not((inputs(193)) or (inputs(208)));
    layer0_outputs(3512) <= '0';
    layer0_outputs(3513) <= not(inputs(245));
    layer0_outputs(3514) <= not(inputs(103));
    layer0_outputs(3515) <= not(inputs(36)) or (inputs(133));
    layer0_outputs(3516) <= inputs(186);
    layer0_outputs(3517) <= not(inputs(36)) or (inputs(142));
    layer0_outputs(3518) <= '0';
    layer0_outputs(3519) <= '0';
    layer0_outputs(3520) <= (inputs(121)) and (inputs(135));
    layer0_outputs(3521) <= (inputs(32)) xor (inputs(139));
    layer0_outputs(3522) <= inputs(102);
    layer0_outputs(3523) <= not(inputs(239)) or (inputs(82));
    layer0_outputs(3524) <= not(inputs(167)) or (inputs(130));
    layer0_outputs(3525) <= inputs(88);
    layer0_outputs(3526) <= not(inputs(151)) or (inputs(189));
    layer0_outputs(3527) <= (inputs(92)) xor (inputs(48));
    layer0_outputs(3528) <= not(inputs(178));
    layer0_outputs(3529) <= '0';
    layer0_outputs(3530) <= not(inputs(45));
    layer0_outputs(3531) <= '0';
    layer0_outputs(3532) <= (inputs(230)) and not (inputs(105));
    layer0_outputs(3533) <= not(inputs(200));
    layer0_outputs(3534) <= inputs(129);
    layer0_outputs(3535) <= (inputs(41)) or (inputs(146));
    layer0_outputs(3536) <= not((inputs(162)) or (inputs(34)));
    layer0_outputs(3537) <= '0';
    layer0_outputs(3538) <= not(inputs(100));
    layer0_outputs(3539) <= (inputs(213)) and (inputs(57));
    layer0_outputs(3540) <= inputs(105);
    layer0_outputs(3541) <= not(inputs(83));
    layer0_outputs(3542) <= (inputs(197)) or (inputs(179));
    layer0_outputs(3543) <= not(inputs(37)) or (inputs(196));
    layer0_outputs(3544) <= (inputs(154)) and not (inputs(80));
    layer0_outputs(3545) <= inputs(12);
    layer0_outputs(3546) <= not((inputs(180)) and (inputs(173)));
    layer0_outputs(3547) <= not(inputs(60));
    layer0_outputs(3548) <= (inputs(123)) and not (inputs(240));
    layer0_outputs(3549) <= inputs(1);
    layer0_outputs(3550) <= not((inputs(196)) or (inputs(220)));
    layer0_outputs(3551) <= not((inputs(24)) or (inputs(202)));
    layer0_outputs(3552) <= not(inputs(111));
    layer0_outputs(3553) <= not(inputs(160));
    layer0_outputs(3554) <= (inputs(183)) xor (inputs(181));
    layer0_outputs(3555) <= '0';
    layer0_outputs(3556) <= (inputs(198)) and not (inputs(11));
    layer0_outputs(3557) <= inputs(26);
    layer0_outputs(3558) <= (inputs(68)) xor (inputs(80));
    layer0_outputs(3559) <= inputs(171);
    layer0_outputs(3560) <= not(inputs(236)) or (inputs(240));
    layer0_outputs(3561) <= (inputs(87)) and not (inputs(240));
    layer0_outputs(3562) <= not(inputs(115));
    layer0_outputs(3563) <= (inputs(252)) or (inputs(169));
    layer0_outputs(3564) <= not(inputs(61));
    layer0_outputs(3565) <= not((inputs(142)) or (inputs(247)));
    layer0_outputs(3566) <= not(inputs(214)) or (inputs(120));
    layer0_outputs(3567) <= inputs(13);
    layer0_outputs(3568) <= (inputs(230)) and not (inputs(167));
    layer0_outputs(3569) <= (inputs(4)) and not (inputs(66));
    layer0_outputs(3570) <= (inputs(235)) and not (inputs(161));
    layer0_outputs(3571) <= '0';
    layer0_outputs(3572) <= inputs(109);
    layer0_outputs(3573) <= '0';
    layer0_outputs(3574) <= '0';
    layer0_outputs(3575) <= '1';
    layer0_outputs(3576) <= not((inputs(239)) or (inputs(102)));
    layer0_outputs(3577) <= '0';
    layer0_outputs(3578) <= (inputs(166)) or (inputs(18));
    layer0_outputs(3579) <= (inputs(92)) or (inputs(68));
    layer0_outputs(3580) <= (inputs(4)) or (inputs(208));
    layer0_outputs(3581) <= inputs(102);
    layer0_outputs(3582) <= not(inputs(70)) or (inputs(77));
    layer0_outputs(3583) <= '1';
    layer0_outputs(3584) <= not(inputs(129));
    layer0_outputs(3585) <= (inputs(37)) and not (inputs(161));
    layer0_outputs(3586) <= inputs(161);
    layer0_outputs(3587) <= not(inputs(39)) or (inputs(135));
    layer0_outputs(3588) <= (inputs(119)) and not (inputs(176));
    layer0_outputs(3589) <= not(inputs(85));
    layer0_outputs(3590) <= (inputs(117)) and (inputs(59));
    layer0_outputs(3591) <= '0';
    layer0_outputs(3592) <= not(inputs(33));
    layer0_outputs(3593) <= not(inputs(152));
    layer0_outputs(3594) <= not((inputs(113)) or (inputs(125)));
    layer0_outputs(3595) <= not((inputs(83)) xor (inputs(22)));
    layer0_outputs(3596) <= (inputs(5)) or (inputs(91));
    layer0_outputs(3597) <= '0';
    layer0_outputs(3598) <= '1';
    layer0_outputs(3599) <= inputs(103);
    layer0_outputs(3600) <= (inputs(231)) or (inputs(213));
    layer0_outputs(3601) <= not(inputs(14));
    layer0_outputs(3602) <= (inputs(196)) or (inputs(145));
    layer0_outputs(3603) <= not(inputs(104));
    layer0_outputs(3604) <= (inputs(252)) or (inputs(53));
    layer0_outputs(3605) <= not((inputs(35)) or (inputs(63)));
    layer0_outputs(3606) <= (inputs(40)) and not (inputs(185));
    layer0_outputs(3607) <= (inputs(127)) and not (inputs(243));
    layer0_outputs(3608) <= not(inputs(150));
    layer0_outputs(3609) <= not(inputs(64));
    layer0_outputs(3610) <= '0';
    layer0_outputs(3611) <= not((inputs(203)) and (inputs(240)));
    layer0_outputs(3612) <= (inputs(160)) xor (inputs(126));
    layer0_outputs(3613) <= inputs(225);
    layer0_outputs(3614) <= not(inputs(52));
    layer0_outputs(3615) <= inputs(199);
    layer0_outputs(3616) <= not(inputs(155)) or (inputs(7));
    layer0_outputs(3617) <= not(inputs(122));
    layer0_outputs(3618) <= not(inputs(89)) or (inputs(197));
    layer0_outputs(3619) <= not(inputs(16));
    layer0_outputs(3620) <= (inputs(4)) and not (inputs(114));
    layer0_outputs(3621) <= not(inputs(188));
    layer0_outputs(3622) <= (inputs(219)) and not (inputs(66));
    layer0_outputs(3623) <= not(inputs(35));
    layer0_outputs(3624) <= (inputs(177)) and not (inputs(121));
    layer0_outputs(3625) <= not((inputs(91)) or (inputs(141)));
    layer0_outputs(3626) <= (inputs(129)) xor (inputs(20));
    layer0_outputs(3627) <= inputs(163);
    layer0_outputs(3628) <= (inputs(66)) xor (inputs(172));
    layer0_outputs(3629) <= (inputs(20)) or (inputs(47));
    layer0_outputs(3630) <= inputs(62);
    layer0_outputs(3631) <= not((inputs(177)) xor (inputs(217)));
    layer0_outputs(3632) <= (inputs(63)) and (inputs(57));
    layer0_outputs(3633) <= (inputs(237)) and (inputs(223));
    layer0_outputs(3634) <= not(inputs(246)) or (inputs(96));
    layer0_outputs(3635) <= not(inputs(232));
    layer0_outputs(3636) <= '1';
    layer0_outputs(3637) <= (inputs(80)) xor (inputs(235));
    layer0_outputs(3638) <= not(inputs(232));
    layer0_outputs(3639) <= inputs(165);
    layer0_outputs(3640) <= not((inputs(122)) or (inputs(15)));
    layer0_outputs(3641) <= (inputs(130)) or (inputs(113));
    layer0_outputs(3642) <= not(inputs(109));
    layer0_outputs(3643) <= inputs(98);
    layer0_outputs(3644) <= not((inputs(174)) xor (inputs(53)));
    layer0_outputs(3645) <= (inputs(98)) or (inputs(77));
    layer0_outputs(3646) <= not(inputs(46));
    layer0_outputs(3647) <= not(inputs(111)) or (inputs(24));
    layer0_outputs(3648) <= inputs(125);
    layer0_outputs(3649) <= not(inputs(60));
    layer0_outputs(3650) <= not(inputs(21)) or (inputs(185));
    layer0_outputs(3651) <= (inputs(167)) and (inputs(19));
    layer0_outputs(3652) <= not(inputs(146));
    layer0_outputs(3653) <= not(inputs(149));
    layer0_outputs(3654) <= (inputs(123)) or (inputs(85));
    layer0_outputs(3655) <= (inputs(178)) and not (inputs(45));
    layer0_outputs(3656) <= not(inputs(120)) or (inputs(129));
    layer0_outputs(3657) <= (inputs(204)) xor (inputs(146));
    layer0_outputs(3658) <= not((inputs(214)) and (inputs(55)));
    layer0_outputs(3659) <= not(inputs(135));
    layer0_outputs(3660) <= not(inputs(103)) or (inputs(79));
    layer0_outputs(3661) <= '0';
    layer0_outputs(3662) <= not(inputs(214)) or (inputs(14));
    layer0_outputs(3663) <= not(inputs(161)) or (inputs(109));
    layer0_outputs(3664) <= not(inputs(60));
    layer0_outputs(3665) <= inputs(23);
    layer0_outputs(3666) <= not((inputs(229)) or (inputs(177)));
    layer0_outputs(3667) <= (inputs(18)) xor (inputs(116));
    layer0_outputs(3668) <= not(inputs(84));
    layer0_outputs(3669) <= not((inputs(5)) and (inputs(238)));
    layer0_outputs(3670) <= inputs(126);
    layer0_outputs(3671) <= not(inputs(155)) or (inputs(179));
    layer0_outputs(3672) <= not(inputs(14)) or (inputs(62));
    layer0_outputs(3673) <= not(inputs(111));
    layer0_outputs(3674) <= not((inputs(140)) and (inputs(139)));
    layer0_outputs(3675) <= not(inputs(223)) or (inputs(65));
    layer0_outputs(3676) <= not(inputs(182));
    layer0_outputs(3677) <= '0';
    layer0_outputs(3678) <= (inputs(91)) or (inputs(35));
    layer0_outputs(3679) <= inputs(203);
    layer0_outputs(3680) <= not((inputs(109)) or (inputs(2)));
    layer0_outputs(3681) <= not(inputs(15)) or (inputs(16));
    layer0_outputs(3682) <= not(inputs(229)) or (inputs(58));
    layer0_outputs(3683) <= not(inputs(132));
    layer0_outputs(3684) <= '0';
    layer0_outputs(3685) <= not((inputs(120)) or (inputs(93)));
    layer0_outputs(3686) <= not(inputs(116));
    layer0_outputs(3687) <= (inputs(76)) or (inputs(177));
    layer0_outputs(3688) <= '0';
    layer0_outputs(3689) <= (inputs(186)) or (inputs(172));
    layer0_outputs(3690) <= inputs(156);
    layer0_outputs(3691) <= inputs(211);
    layer0_outputs(3692) <= (inputs(224)) and (inputs(254));
    layer0_outputs(3693) <= not(inputs(104)) or (inputs(162));
    layer0_outputs(3694) <= (inputs(63)) and not (inputs(185));
    layer0_outputs(3695) <= '1';
    layer0_outputs(3696) <= not(inputs(125));
    layer0_outputs(3697) <= (inputs(43)) and not (inputs(222));
    layer0_outputs(3698) <= (inputs(72)) and (inputs(209));
    layer0_outputs(3699) <= '0';
    layer0_outputs(3700) <= not(inputs(179)) or (inputs(50));
    layer0_outputs(3701) <= '1';
    layer0_outputs(3702) <= not((inputs(85)) and (inputs(121)));
    layer0_outputs(3703) <= not(inputs(227));
    layer0_outputs(3704) <= inputs(178);
    layer0_outputs(3705) <= not(inputs(160));
    layer0_outputs(3706) <= '0';
    layer0_outputs(3707) <= not(inputs(57)) or (inputs(88));
    layer0_outputs(3708) <= '1';
    layer0_outputs(3709) <= not(inputs(70)) or (inputs(124));
    layer0_outputs(3710) <= '1';
    layer0_outputs(3711) <= (inputs(245)) or (inputs(112));
    layer0_outputs(3712) <= (inputs(162)) and (inputs(162));
    layer0_outputs(3713) <= inputs(19);
    layer0_outputs(3714) <= not((inputs(88)) or (inputs(152)));
    layer0_outputs(3715) <= (inputs(106)) and not (inputs(84));
    layer0_outputs(3716) <= (inputs(221)) and not (inputs(96));
    layer0_outputs(3717) <= not((inputs(222)) xor (inputs(120)));
    layer0_outputs(3718) <= inputs(58);
    layer0_outputs(3719) <= '0';
    layer0_outputs(3720) <= not(inputs(208)) or (inputs(175));
    layer0_outputs(3721) <= not(inputs(178)) or (inputs(253));
    layer0_outputs(3722) <= not(inputs(190));
    layer0_outputs(3723) <= not(inputs(167));
    layer0_outputs(3724) <= not((inputs(104)) or (inputs(193)));
    layer0_outputs(3725) <= inputs(187);
    layer0_outputs(3726) <= not(inputs(170)) or (inputs(199));
    layer0_outputs(3727) <= '1';
    layer0_outputs(3728) <= not(inputs(173));
    layer0_outputs(3729) <= (inputs(45)) and not (inputs(254));
    layer0_outputs(3730) <= not((inputs(100)) and (inputs(212)));
    layer0_outputs(3731) <= (inputs(3)) xor (inputs(171));
    layer0_outputs(3732) <= '1';
    layer0_outputs(3733) <= not((inputs(245)) or (inputs(104)));
    layer0_outputs(3734) <= inputs(44);
    layer0_outputs(3735) <= not(inputs(103)) or (inputs(247));
    layer0_outputs(3736) <= not((inputs(171)) or (inputs(79)));
    layer0_outputs(3737) <= '1';
    layer0_outputs(3738) <= (inputs(89)) and not (inputs(49));
    layer0_outputs(3739) <= (inputs(21)) and not (inputs(179));
    layer0_outputs(3740) <= not(inputs(184));
    layer0_outputs(3741) <= (inputs(14)) and not (inputs(235));
    layer0_outputs(3742) <= not(inputs(165));
    layer0_outputs(3743) <= not(inputs(85)) or (inputs(56));
    layer0_outputs(3744) <= not((inputs(72)) and (inputs(14)));
    layer0_outputs(3745) <= not((inputs(121)) or (inputs(229)));
    layer0_outputs(3746) <= not(inputs(128));
    layer0_outputs(3747) <= inputs(62);
    layer0_outputs(3748) <= (inputs(242)) and (inputs(133));
    layer0_outputs(3749) <= not(inputs(31)) or (inputs(177));
    layer0_outputs(3750) <= '1';
    layer0_outputs(3751) <= not((inputs(181)) xor (inputs(47)));
    layer0_outputs(3752) <= not(inputs(175)) or (inputs(62));
    layer0_outputs(3753) <= (inputs(242)) or (inputs(200));
    layer0_outputs(3754) <= (inputs(59)) and (inputs(61));
    layer0_outputs(3755) <= not((inputs(86)) xor (inputs(102)));
    layer0_outputs(3756) <= (inputs(152)) and (inputs(213));
    layer0_outputs(3757) <= (inputs(197)) and not (inputs(68));
    layer0_outputs(3758) <= not((inputs(47)) xor (inputs(34)));
    layer0_outputs(3759) <= not((inputs(185)) xor (inputs(31)));
    layer0_outputs(3760) <= inputs(49);
    layer0_outputs(3761) <= not((inputs(124)) xor (inputs(31)));
    layer0_outputs(3762) <= (inputs(24)) and (inputs(89));
    layer0_outputs(3763) <= not((inputs(147)) and (inputs(117)));
    layer0_outputs(3764) <= not(inputs(194));
    layer0_outputs(3765) <= not((inputs(152)) or (inputs(74)));
    layer0_outputs(3766) <= (inputs(242)) or (inputs(239));
    layer0_outputs(3767) <= not((inputs(108)) or (inputs(138)));
    layer0_outputs(3768) <= (inputs(73)) and not (inputs(53));
    layer0_outputs(3769) <= not(inputs(122));
    layer0_outputs(3770) <= inputs(8);
    layer0_outputs(3771) <= inputs(93);
    layer0_outputs(3772) <= inputs(159);
    layer0_outputs(3773) <= not((inputs(32)) or (inputs(253)));
    layer0_outputs(3774) <= inputs(97);
    layer0_outputs(3775) <= not((inputs(49)) or (inputs(156)));
    layer0_outputs(3776) <= not((inputs(171)) xor (inputs(236)));
    layer0_outputs(3777) <= (inputs(123)) or (inputs(220));
    layer0_outputs(3778) <= '1';
    layer0_outputs(3779) <= (inputs(213)) and (inputs(124));
    layer0_outputs(3780) <= inputs(203);
    layer0_outputs(3781) <= (inputs(23)) xor (inputs(129));
    layer0_outputs(3782) <= not((inputs(222)) xor (inputs(211)));
    layer0_outputs(3783) <= inputs(2);
    layer0_outputs(3784) <= not(inputs(206)) or (inputs(11));
    layer0_outputs(3785) <= not(inputs(236));
    layer0_outputs(3786) <= (inputs(205)) or (inputs(245));
    layer0_outputs(3787) <= not(inputs(58)) or (inputs(211));
    layer0_outputs(3788) <= inputs(7);
    layer0_outputs(3789) <= '1';
    layer0_outputs(3790) <= not(inputs(121)) or (inputs(222));
    layer0_outputs(3791) <= not(inputs(197)) or (inputs(170));
    layer0_outputs(3792) <= not(inputs(86));
    layer0_outputs(3793) <= (inputs(240)) xor (inputs(223));
    layer0_outputs(3794) <= inputs(107);
    layer0_outputs(3795) <= (inputs(202)) or (inputs(130));
    layer0_outputs(3796) <= (inputs(13)) or (inputs(79));
    layer0_outputs(3797) <= not((inputs(154)) or (inputs(75)));
    layer0_outputs(3798) <= (inputs(195)) or (inputs(164));
    layer0_outputs(3799) <= (inputs(241)) or (inputs(41));
    layer0_outputs(3800) <= '0';
    layer0_outputs(3801) <= (inputs(78)) and not (inputs(47));
    layer0_outputs(3802) <= inputs(108);
    layer0_outputs(3803) <= not(inputs(240)) or (inputs(185));
    layer0_outputs(3804) <= (inputs(149)) and (inputs(171));
    layer0_outputs(3805) <= not(inputs(157)) or (inputs(59));
    layer0_outputs(3806) <= not((inputs(189)) or (inputs(204)));
    layer0_outputs(3807) <= '1';
    layer0_outputs(3808) <= not(inputs(86)) or (inputs(115));
    layer0_outputs(3809) <= not(inputs(120)) or (inputs(146));
    layer0_outputs(3810) <= (inputs(69)) and not (inputs(159));
    layer0_outputs(3811) <= (inputs(46)) and not (inputs(218));
    layer0_outputs(3812) <= (inputs(137)) and not (inputs(188));
    layer0_outputs(3813) <= inputs(237);
    layer0_outputs(3814) <= (inputs(117)) and not (inputs(33));
    layer0_outputs(3815) <= '0';
    layer0_outputs(3816) <= not((inputs(201)) or (inputs(237)));
    layer0_outputs(3817) <= (inputs(29)) and not (inputs(175));
    layer0_outputs(3818) <= (inputs(62)) and (inputs(254));
    layer0_outputs(3819) <= inputs(132);
    layer0_outputs(3820) <= inputs(249);
    layer0_outputs(3821) <= (inputs(189)) or (inputs(40));
    layer0_outputs(3822) <= not((inputs(170)) xor (inputs(104)));
    layer0_outputs(3823) <= '0';
    layer0_outputs(3824) <= (inputs(118)) xor (inputs(115));
    layer0_outputs(3825) <= not((inputs(50)) or (inputs(106)));
    layer0_outputs(3826) <= (inputs(68)) and not (inputs(178));
    layer0_outputs(3827) <= not((inputs(127)) xor (inputs(24)));
    layer0_outputs(3828) <= not(inputs(230)) or (inputs(240));
    layer0_outputs(3829) <= '1';
    layer0_outputs(3830) <= not(inputs(164));
    layer0_outputs(3831) <= not(inputs(238));
    layer0_outputs(3832) <= (inputs(90)) or (inputs(144));
    layer0_outputs(3833) <= (inputs(128)) or (inputs(235));
    layer0_outputs(3834) <= not((inputs(48)) or (inputs(166)));
    layer0_outputs(3835) <= (inputs(45)) or (inputs(40));
    layer0_outputs(3836) <= not(inputs(136));
    layer0_outputs(3837) <= '0';
    layer0_outputs(3838) <= '0';
    layer0_outputs(3839) <= not(inputs(152)) or (inputs(87));
    layer0_outputs(3840) <= '1';
    layer0_outputs(3841) <= '0';
    layer0_outputs(3842) <= inputs(89);
    layer0_outputs(3843) <= not((inputs(187)) or (inputs(61)));
    layer0_outputs(3844) <= (inputs(226)) or (inputs(175));
    layer0_outputs(3845) <= (inputs(180)) and not (inputs(97));
    layer0_outputs(3846) <= not(inputs(118));
    layer0_outputs(3847) <= (inputs(26)) xor (inputs(48));
    layer0_outputs(3848) <= not((inputs(10)) or (inputs(190)));
    layer0_outputs(3849) <= inputs(142);
    layer0_outputs(3850) <= not(inputs(46));
    layer0_outputs(3851) <= (inputs(83)) or (inputs(173));
    layer0_outputs(3852) <= not((inputs(157)) or (inputs(82)));
    layer0_outputs(3853) <= inputs(192);
    layer0_outputs(3854) <= '0';
    layer0_outputs(3855) <= not((inputs(14)) and (inputs(244)));
    layer0_outputs(3856) <= not(inputs(168));
    layer0_outputs(3857) <= not((inputs(254)) or (inputs(138)));
    layer0_outputs(3858) <= inputs(117);
    layer0_outputs(3859) <= not(inputs(94)) or (inputs(14));
    layer0_outputs(3860) <= inputs(104);
    layer0_outputs(3861) <= not((inputs(252)) and (inputs(216)));
    layer0_outputs(3862) <= not(inputs(99));
    layer0_outputs(3863) <= inputs(15);
    layer0_outputs(3864) <= not(inputs(42)) or (inputs(36));
    layer0_outputs(3865) <= (inputs(177)) or (inputs(248));
    layer0_outputs(3866) <= not(inputs(213));
    layer0_outputs(3867) <= (inputs(50)) and not (inputs(214));
    layer0_outputs(3868) <= not((inputs(53)) and (inputs(120)));
    layer0_outputs(3869) <= not(inputs(110));
    layer0_outputs(3870) <= not(inputs(67)) or (inputs(110));
    layer0_outputs(3871) <= not((inputs(28)) xor (inputs(61)));
    layer0_outputs(3872) <= not(inputs(239));
    layer0_outputs(3873) <= not((inputs(10)) or (inputs(45)));
    layer0_outputs(3874) <= (inputs(129)) or (inputs(238));
    layer0_outputs(3875) <= not((inputs(129)) or (inputs(97)));
    layer0_outputs(3876) <= not(inputs(84)) or (inputs(78));
    layer0_outputs(3877) <= (inputs(176)) or (inputs(37));
    layer0_outputs(3878) <= not(inputs(142)) or (inputs(24));
    layer0_outputs(3879) <= (inputs(67)) and not (inputs(170));
    layer0_outputs(3880) <= (inputs(203)) and not (inputs(85));
    layer0_outputs(3881) <= not(inputs(62));
    layer0_outputs(3882) <= '1';
    layer0_outputs(3883) <= (inputs(164)) and not (inputs(28));
    layer0_outputs(3884) <= (inputs(54)) or (inputs(91));
    layer0_outputs(3885) <= not(inputs(42));
    layer0_outputs(3886) <= not(inputs(78));
    layer0_outputs(3887) <= not((inputs(173)) xor (inputs(128)));
    layer0_outputs(3888) <= not((inputs(95)) and (inputs(71)));
    layer0_outputs(3889) <= (inputs(227)) and not (inputs(220));
    layer0_outputs(3890) <= (inputs(36)) and (inputs(219));
    layer0_outputs(3891) <= not(inputs(22));
    layer0_outputs(3892) <= inputs(73);
    layer0_outputs(3893) <= not((inputs(217)) or (inputs(141)));
    layer0_outputs(3894) <= not(inputs(101));
    layer0_outputs(3895) <= not(inputs(96)) or (inputs(167));
    layer0_outputs(3896) <= not((inputs(72)) or (inputs(208)));
    layer0_outputs(3897) <= inputs(84);
    layer0_outputs(3898) <= (inputs(36)) or (inputs(119));
    layer0_outputs(3899) <= not(inputs(244));
    layer0_outputs(3900) <= not(inputs(97)) or (inputs(137));
    layer0_outputs(3901) <= inputs(142);
    layer0_outputs(3902) <= (inputs(108)) and (inputs(209));
    layer0_outputs(3903) <= '1';
    layer0_outputs(3904) <= not(inputs(94)) or (inputs(110));
    layer0_outputs(3905) <= not((inputs(164)) xor (inputs(128)));
    layer0_outputs(3906) <= (inputs(191)) or (inputs(106));
    layer0_outputs(3907) <= not(inputs(182));
    layer0_outputs(3908) <= not((inputs(75)) xor (inputs(4)));
    layer0_outputs(3909) <= '1';
    layer0_outputs(3910) <= inputs(81);
    layer0_outputs(3911) <= (inputs(156)) or (inputs(128));
    layer0_outputs(3912) <= not((inputs(169)) or (inputs(151)));
    layer0_outputs(3913) <= (inputs(153)) and (inputs(212));
    layer0_outputs(3914) <= '0';
    layer0_outputs(3915) <= (inputs(247)) and (inputs(100));
    layer0_outputs(3916) <= (inputs(172)) and not (inputs(224));
    layer0_outputs(3917) <= not(inputs(231));
    layer0_outputs(3918) <= not((inputs(1)) or (inputs(222)));
    layer0_outputs(3919) <= '1';
    layer0_outputs(3920) <= not(inputs(189));
    layer0_outputs(3921) <= not(inputs(176));
    layer0_outputs(3922) <= not((inputs(145)) xor (inputs(247)));
    layer0_outputs(3923) <= not(inputs(90));
    layer0_outputs(3924) <= (inputs(171)) or (inputs(219));
    layer0_outputs(3925) <= (inputs(232)) and not (inputs(125));
    layer0_outputs(3926) <= (inputs(155)) xor (inputs(17));
    layer0_outputs(3927) <= not(inputs(204)) or (inputs(150));
    layer0_outputs(3928) <= inputs(30);
    layer0_outputs(3929) <= inputs(14);
    layer0_outputs(3930) <= (inputs(159)) and not (inputs(182));
    layer0_outputs(3931) <= inputs(33);
    layer0_outputs(3932) <= (inputs(99)) and not (inputs(218));
    layer0_outputs(3933) <= not((inputs(70)) or (inputs(79)));
    layer0_outputs(3934) <= (inputs(51)) and (inputs(224));
    layer0_outputs(3935) <= not((inputs(160)) xor (inputs(6)));
    layer0_outputs(3936) <= not(inputs(168));
    layer0_outputs(3937) <= (inputs(48)) and not (inputs(221));
    layer0_outputs(3938) <= (inputs(237)) and (inputs(217));
    layer0_outputs(3939) <= not(inputs(144)) or (inputs(154));
    layer0_outputs(3940) <= (inputs(178)) and not (inputs(231));
    layer0_outputs(3941) <= (inputs(230)) and not (inputs(130));
    layer0_outputs(3942) <= not(inputs(195)) or (inputs(47));
    layer0_outputs(3943) <= not(inputs(222)) or (inputs(231));
    layer0_outputs(3944) <= not((inputs(175)) or (inputs(228)));
    layer0_outputs(3945) <= (inputs(216)) and not (inputs(132));
    layer0_outputs(3946) <= not((inputs(251)) or (inputs(135)));
    layer0_outputs(3947) <= not((inputs(44)) or (inputs(5)));
    layer0_outputs(3948) <= (inputs(172)) or (inputs(188));
    layer0_outputs(3949) <= inputs(238);
    layer0_outputs(3950) <= '0';
    layer0_outputs(3951) <= '0';
    layer0_outputs(3952) <= (inputs(145)) or (inputs(227));
    layer0_outputs(3953) <= not(inputs(152));
    layer0_outputs(3954) <= not((inputs(221)) or (inputs(146)));
    layer0_outputs(3955) <= not(inputs(204)) or (inputs(45));
    layer0_outputs(3956) <= not((inputs(181)) or (inputs(129)));
    layer0_outputs(3957) <= not((inputs(250)) or (inputs(223)));
    layer0_outputs(3958) <= not(inputs(126));
    layer0_outputs(3959) <= inputs(112);
    layer0_outputs(3960) <= not(inputs(114)) or (inputs(39));
    layer0_outputs(3961) <= inputs(77);
    layer0_outputs(3962) <= not(inputs(229)) or (inputs(1));
    layer0_outputs(3963) <= not(inputs(44)) or (inputs(138));
    layer0_outputs(3964) <= '1';
    layer0_outputs(3965) <= not(inputs(160));
    layer0_outputs(3966) <= '0';
    layer0_outputs(3967) <= not((inputs(191)) or (inputs(155)));
    layer0_outputs(3968) <= not(inputs(243)) or (inputs(14));
    layer0_outputs(3969) <= not((inputs(106)) or (inputs(90)));
    layer0_outputs(3970) <= (inputs(46)) or (inputs(186));
    layer0_outputs(3971) <= (inputs(92)) or (inputs(128));
    layer0_outputs(3972) <= (inputs(48)) or (inputs(33));
    layer0_outputs(3973) <= (inputs(73)) and (inputs(174));
    layer0_outputs(3974) <= not(inputs(89)) or (inputs(106));
    layer0_outputs(3975) <= not(inputs(13));
    layer0_outputs(3976) <= inputs(90);
    layer0_outputs(3977) <= not((inputs(122)) and (inputs(155)));
    layer0_outputs(3978) <= inputs(48);
    layer0_outputs(3979) <= '1';
    layer0_outputs(3980) <= (inputs(71)) and (inputs(184));
    layer0_outputs(3981) <= inputs(166);
    layer0_outputs(3982) <= '1';
    layer0_outputs(3983) <= (inputs(10)) and (inputs(91));
    layer0_outputs(3984) <= inputs(60);
    layer0_outputs(3985) <= (inputs(230)) and not (inputs(165));
    layer0_outputs(3986) <= inputs(88);
    layer0_outputs(3987) <= inputs(102);
    layer0_outputs(3988) <= (inputs(145)) or (inputs(176));
    layer0_outputs(3989) <= not((inputs(208)) and (inputs(28)));
    layer0_outputs(3990) <= inputs(231);
    layer0_outputs(3991) <= inputs(92);
    layer0_outputs(3992) <= not(inputs(74)) or (inputs(202));
    layer0_outputs(3993) <= not(inputs(138));
    layer0_outputs(3994) <= not(inputs(132)) or (inputs(180));
    layer0_outputs(3995) <= not((inputs(159)) or (inputs(103)));
    layer0_outputs(3996) <= (inputs(145)) or (inputs(246));
    layer0_outputs(3997) <= '0';
    layer0_outputs(3998) <= not(inputs(171)) or (inputs(92));
    layer0_outputs(3999) <= (inputs(76)) xor (inputs(78));
    layer0_outputs(4000) <= inputs(253);
    layer0_outputs(4001) <= not(inputs(41));
    layer0_outputs(4002) <= (inputs(104)) and not (inputs(254));
    layer0_outputs(4003) <= '1';
    layer0_outputs(4004) <= (inputs(100)) and not (inputs(73));
    layer0_outputs(4005) <= (inputs(210)) or (inputs(252));
    layer0_outputs(4006) <= (inputs(255)) xor (inputs(191));
    layer0_outputs(4007) <= not(inputs(199)) or (inputs(27));
    layer0_outputs(4008) <= not((inputs(237)) or (inputs(118)));
    layer0_outputs(4009) <= inputs(148);
    layer0_outputs(4010) <= not(inputs(237)) or (inputs(50));
    layer0_outputs(4011) <= not(inputs(61));
    layer0_outputs(4012) <= inputs(205);
    layer0_outputs(4013) <= (inputs(93)) xor (inputs(0));
    layer0_outputs(4014) <= (inputs(41)) or (inputs(83));
    layer0_outputs(4015) <= not(inputs(202));
    layer0_outputs(4016) <= (inputs(15)) xor (inputs(126));
    layer0_outputs(4017) <= (inputs(122)) and (inputs(60));
    layer0_outputs(4018) <= not((inputs(62)) or (inputs(141)));
    layer0_outputs(4019) <= inputs(49);
    layer0_outputs(4020) <= not(inputs(152)) or (inputs(24));
    layer0_outputs(4021) <= not(inputs(26));
    layer0_outputs(4022) <= '0';
    layer0_outputs(4023) <= not((inputs(243)) or (inputs(223)));
    layer0_outputs(4024) <= not(inputs(221)) or (inputs(221));
    layer0_outputs(4025) <= '0';
    layer0_outputs(4026) <= not(inputs(92)) or (inputs(117));
    layer0_outputs(4027) <= not((inputs(160)) or (inputs(175)));
    layer0_outputs(4028) <= not(inputs(129));
    layer0_outputs(4029) <= (inputs(119)) and not (inputs(127));
    layer0_outputs(4030) <= (inputs(85)) and (inputs(151));
    layer0_outputs(4031) <= '1';
    layer0_outputs(4032) <= (inputs(54)) and not (inputs(135));
    layer0_outputs(4033) <= (inputs(136)) and not (inputs(112));
    layer0_outputs(4034) <= inputs(157);
    layer0_outputs(4035) <= not((inputs(174)) or (inputs(50)));
    layer0_outputs(4036) <= not((inputs(63)) or (inputs(229)));
    layer0_outputs(4037) <= not(inputs(82));
    layer0_outputs(4038) <= not(inputs(220));
    layer0_outputs(4039) <= not((inputs(85)) or (inputs(192)));
    layer0_outputs(4040) <= inputs(176);
    layer0_outputs(4041) <= inputs(82);
    layer0_outputs(4042) <= not((inputs(176)) or (inputs(233)));
    layer0_outputs(4043) <= (inputs(140)) or (inputs(20));
    layer0_outputs(4044) <= (inputs(170)) or (inputs(92));
    layer0_outputs(4045) <= not(inputs(163));
    layer0_outputs(4046) <= (inputs(223)) or (inputs(184));
    layer0_outputs(4047) <= '1';
    layer0_outputs(4048) <= not((inputs(210)) and (inputs(154)));
    layer0_outputs(4049) <= not((inputs(30)) or (inputs(186)));
    layer0_outputs(4050) <= not(inputs(210));
    layer0_outputs(4051) <= (inputs(203)) and not (inputs(79));
    layer0_outputs(4052) <= not(inputs(199)) or (inputs(92));
    layer0_outputs(4053) <= (inputs(44)) and not (inputs(108));
    layer0_outputs(4054) <= inputs(1);
    layer0_outputs(4055) <= (inputs(117)) or (inputs(14));
    layer0_outputs(4056) <= (inputs(95)) or (inputs(145));
    layer0_outputs(4057) <= inputs(81);
    layer0_outputs(4058) <= not(inputs(203));
    layer0_outputs(4059) <= not((inputs(45)) or (inputs(102)));
    layer0_outputs(4060) <= (inputs(81)) and not (inputs(123));
    layer0_outputs(4061) <= not(inputs(126));
    layer0_outputs(4062) <= inputs(176);
    layer0_outputs(4063) <= (inputs(77)) or (inputs(216));
    layer0_outputs(4064) <= (inputs(203)) or (inputs(161));
    layer0_outputs(4065) <= not(inputs(28)) or (inputs(28));
    layer0_outputs(4066) <= '1';
    layer0_outputs(4067) <= (inputs(219)) or (inputs(158));
    layer0_outputs(4068) <= inputs(68);
    layer0_outputs(4069) <= not(inputs(202));
    layer0_outputs(4070) <= not(inputs(23)) or (inputs(135));
    layer0_outputs(4071) <= inputs(35);
    layer0_outputs(4072) <= (inputs(70)) xor (inputs(255));
    layer0_outputs(4073) <= not((inputs(63)) and (inputs(5)));
    layer0_outputs(4074) <= (inputs(239)) or (inputs(146));
    layer0_outputs(4075) <= not((inputs(18)) xor (inputs(18)));
    layer0_outputs(4076) <= (inputs(230)) and not (inputs(103));
    layer0_outputs(4077) <= not((inputs(190)) or (inputs(178)));
    layer0_outputs(4078) <= not(inputs(117)) or (inputs(78));
    layer0_outputs(4079) <= not((inputs(78)) xor (inputs(124)));
    layer0_outputs(4080) <= inputs(24);
    layer0_outputs(4081) <= (inputs(16)) and not (inputs(168));
    layer0_outputs(4082) <= not(inputs(132));
    layer0_outputs(4083) <= not(inputs(188));
    layer0_outputs(4084) <= (inputs(179)) and not (inputs(78));
    layer0_outputs(4085) <= '1';
    layer0_outputs(4086) <= inputs(146);
    layer0_outputs(4087) <= not(inputs(46)) or (inputs(236));
    layer0_outputs(4088) <= inputs(227);
    layer0_outputs(4089) <= inputs(95);
    layer0_outputs(4090) <= '0';
    layer0_outputs(4091) <= not(inputs(149)) or (inputs(18));
    layer0_outputs(4092) <= not(inputs(244)) or (inputs(131));
    layer0_outputs(4093) <= '0';
    layer0_outputs(4094) <= (inputs(168)) and not (inputs(222));
    layer0_outputs(4095) <= (inputs(73)) and not (inputs(68));
    layer0_outputs(4096) <= inputs(90);
    layer0_outputs(4097) <= inputs(186);
    layer0_outputs(4098) <= not((inputs(95)) or (inputs(100)));
    layer0_outputs(4099) <= inputs(164);
    layer0_outputs(4100) <= '1';
    layer0_outputs(4101) <= '0';
    layer0_outputs(4102) <= '1';
    layer0_outputs(4103) <= not(inputs(97));
    layer0_outputs(4104) <= not(inputs(164));
    layer0_outputs(4105) <= inputs(46);
    layer0_outputs(4106) <= not((inputs(217)) and (inputs(205)));
    layer0_outputs(4107) <= (inputs(177)) xor (inputs(144));
    layer0_outputs(4108) <= '1';
    layer0_outputs(4109) <= (inputs(239)) and not (inputs(175));
    layer0_outputs(4110) <= inputs(169);
    layer0_outputs(4111) <= not(inputs(187));
    layer0_outputs(4112) <= not(inputs(128));
    layer0_outputs(4113) <= (inputs(119)) or (inputs(233));
    layer0_outputs(4114) <= not(inputs(189)) or (inputs(192));
    layer0_outputs(4115) <= inputs(89);
    layer0_outputs(4116) <= (inputs(205)) xor (inputs(4));
    layer0_outputs(4117) <= inputs(215);
    layer0_outputs(4118) <= not(inputs(70));
    layer0_outputs(4119) <= not(inputs(234));
    layer0_outputs(4120) <= not(inputs(58)) or (inputs(110));
    layer0_outputs(4121) <= (inputs(219)) and not (inputs(174));
    layer0_outputs(4122) <= not(inputs(129));
    layer0_outputs(4123) <= inputs(84);
    layer0_outputs(4124) <= '0';
    layer0_outputs(4125) <= not((inputs(252)) or (inputs(117)));
    layer0_outputs(4126) <= not(inputs(63));
    layer0_outputs(4127) <= inputs(163);
    layer0_outputs(4128) <= not((inputs(173)) or (inputs(32)));
    layer0_outputs(4129) <= not(inputs(173));
    layer0_outputs(4130) <= not(inputs(93));
    layer0_outputs(4131) <= not(inputs(11));
    layer0_outputs(4132) <= not(inputs(46));
    layer0_outputs(4133) <= not(inputs(99));
    layer0_outputs(4134) <= '0';
    layer0_outputs(4135) <= not(inputs(46)) or (inputs(28));
    layer0_outputs(4136) <= (inputs(7)) or (inputs(45));
    layer0_outputs(4137) <= inputs(20);
    layer0_outputs(4138) <= not((inputs(143)) or (inputs(17)));
    layer0_outputs(4139) <= not((inputs(168)) and (inputs(119)));
    layer0_outputs(4140) <= inputs(97);
    layer0_outputs(4141) <= not((inputs(67)) or (inputs(1)));
    layer0_outputs(4142) <= not(inputs(27)) or (inputs(82));
    layer0_outputs(4143) <= (inputs(55)) or (inputs(50));
    layer0_outputs(4144) <= not(inputs(106));
    layer0_outputs(4145) <= not((inputs(170)) or (inputs(218)));
    layer0_outputs(4146) <= not((inputs(159)) or (inputs(53)));
    layer0_outputs(4147) <= (inputs(118)) and not (inputs(16));
    layer0_outputs(4148) <= not(inputs(115)) or (inputs(154));
    layer0_outputs(4149) <= inputs(65);
    layer0_outputs(4150) <= (inputs(101)) xor (inputs(154));
    layer0_outputs(4151) <= (inputs(205)) or (inputs(149));
    layer0_outputs(4152) <= not((inputs(165)) or (inputs(182)));
    layer0_outputs(4153) <= (inputs(19)) and not (inputs(107));
    layer0_outputs(4154) <= inputs(22);
    layer0_outputs(4155) <= '1';
    layer0_outputs(4156) <= inputs(227);
    layer0_outputs(4157) <= (inputs(22)) and not (inputs(129));
    layer0_outputs(4158) <= '0';
    layer0_outputs(4159) <= not(inputs(41));
    layer0_outputs(4160) <= (inputs(39)) xor (inputs(22));
    layer0_outputs(4161) <= '0';
    layer0_outputs(4162) <= '1';
    layer0_outputs(4163) <= not(inputs(240)) or (inputs(128));
    layer0_outputs(4164) <= not((inputs(110)) xor (inputs(35)));
    layer0_outputs(4165) <= (inputs(254)) or (inputs(183));
    layer0_outputs(4166) <= not((inputs(170)) or (inputs(238)));
    layer0_outputs(4167) <= (inputs(123)) and not (inputs(210));
    layer0_outputs(4168) <= inputs(82);
    layer0_outputs(4169) <= '0';
    layer0_outputs(4170) <= (inputs(229)) and not (inputs(66));
    layer0_outputs(4171) <= not((inputs(169)) or (inputs(36)));
    layer0_outputs(4172) <= (inputs(14)) xor (inputs(20));
    layer0_outputs(4173) <= not(inputs(172));
    layer0_outputs(4174) <= (inputs(143)) and (inputs(3));
    layer0_outputs(4175) <= not(inputs(165));
    layer0_outputs(4176) <= not((inputs(120)) or (inputs(64)));
    layer0_outputs(4177) <= (inputs(87)) and (inputs(137));
    layer0_outputs(4178) <= not((inputs(158)) or (inputs(65)));
    layer0_outputs(4179) <= inputs(143);
    layer0_outputs(4180) <= (inputs(67)) and not (inputs(54));
    layer0_outputs(4181) <= inputs(24);
    layer0_outputs(4182) <= (inputs(210)) or (inputs(51));
    layer0_outputs(4183) <= (inputs(221)) xor (inputs(155));
    layer0_outputs(4184) <= inputs(249);
    layer0_outputs(4185) <= (inputs(94)) or (inputs(105));
    layer0_outputs(4186) <= (inputs(137)) and not (inputs(245));
    layer0_outputs(4187) <= (inputs(24)) and not (inputs(144));
    layer0_outputs(4188) <= (inputs(217)) and not (inputs(30));
    layer0_outputs(4189) <= inputs(0);
    layer0_outputs(4190) <= (inputs(78)) or (inputs(138));
    layer0_outputs(4191) <= not(inputs(63)) or (inputs(230));
    layer0_outputs(4192) <= inputs(195);
    layer0_outputs(4193) <= not((inputs(31)) or (inputs(15)));
    layer0_outputs(4194) <= (inputs(21)) and not (inputs(54));
    layer0_outputs(4195) <= (inputs(164)) or (inputs(120));
    layer0_outputs(4196) <= not(inputs(158)) or (inputs(253));
    layer0_outputs(4197) <= (inputs(161)) and (inputs(238));
    layer0_outputs(4198) <= inputs(69);
    layer0_outputs(4199) <= not((inputs(201)) or (inputs(166)));
    layer0_outputs(4200) <= inputs(27);
    layer0_outputs(4201) <= inputs(222);
    layer0_outputs(4202) <= not(inputs(97));
    layer0_outputs(4203) <= (inputs(247)) and not (inputs(157));
    layer0_outputs(4204) <= not(inputs(220));
    layer0_outputs(4205) <= not(inputs(61));
    layer0_outputs(4206) <= not((inputs(193)) xor (inputs(8)));
    layer0_outputs(4207) <= not(inputs(80));
    layer0_outputs(4208) <= (inputs(243)) and not (inputs(121));
    layer0_outputs(4209) <= (inputs(21)) and not (inputs(183));
    layer0_outputs(4210) <= not((inputs(171)) xor (inputs(21)));
    layer0_outputs(4211) <= not((inputs(161)) or (inputs(204)));
    layer0_outputs(4212) <= (inputs(66)) and (inputs(88));
    layer0_outputs(4213) <= not(inputs(182));
    layer0_outputs(4214) <= '1';
    layer0_outputs(4215) <= not(inputs(106));
    layer0_outputs(4216) <= not(inputs(105));
    layer0_outputs(4217) <= not((inputs(147)) and (inputs(225)));
    layer0_outputs(4218) <= '1';
    layer0_outputs(4219) <= not(inputs(162));
    layer0_outputs(4220) <= '1';
    layer0_outputs(4221) <= (inputs(55)) and not (inputs(34));
    layer0_outputs(4222) <= not((inputs(90)) and (inputs(211)));
    layer0_outputs(4223) <= not((inputs(202)) xor (inputs(112)));
    layer0_outputs(4224) <= not(inputs(43));
    layer0_outputs(4225) <= not(inputs(192)) or (inputs(93));
    layer0_outputs(4226) <= not((inputs(163)) or (inputs(95)));
    layer0_outputs(4227) <= inputs(38);
    layer0_outputs(4228) <= inputs(61);
    layer0_outputs(4229) <= '1';
    layer0_outputs(4230) <= not((inputs(18)) or (inputs(20)));
    layer0_outputs(4231) <= (inputs(251)) xor (inputs(53));
    layer0_outputs(4232) <= '1';
    layer0_outputs(4233) <= '1';
    layer0_outputs(4234) <= (inputs(75)) or (inputs(161));
    layer0_outputs(4235) <= not(inputs(14)) or (inputs(175));
    layer0_outputs(4236) <= (inputs(85)) or (inputs(219));
    layer0_outputs(4237) <= inputs(232);
    layer0_outputs(4238) <= (inputs(23)) and not (inputs(184));
    layer0_outputs(4239) <= inputs(62);
    layer0_outputs(4240) <= (inputs(25)) and not (inputs(159));
    layer0_outputs(4241) <= (inputs(143)) and not (inputs(165));
    layer0_outputs(4242) <= (inputs(206)) or (inputs(195));
    layer0_outputs(4243) <= inputs(141);
    layer0_outputs(4244) <= not((inputs(135)) and (inputs(1)));
    layer0_outputs(4245) <= '1';
    layer0_outputs(4246) <= not((inputs(87)) and (inputs(131)));
    layer0_outputs(4247) <= not(inputs(144));
    layer0_outputs(4248) <= (inputs(211)) or (inputs(2));
    layer0_outputs(4249) <= not((inputs(170)) or (inputs(149)));
    layer0_outputs(4250) <= inputs(89);
    layer0_outputs(4251) <= not(inputs(184));
    layer0_outputs(4252) <= '0';
    layer0_outputs(4253) <= not(inputs(142));
    layer0_outputs(4254) <= (inputs(180)) and not (inputs(87));
    layer0_outputs(4255) <= (inputs(27)) xor (inputs(14));
    layer0_outputs(4256) <= (inputs(188)) and not (inputs(60));
    layer0_outputs(4257) <= (inputs(178)) and not (inputs(10));
    layer0_outputs(4258) <= (inputs(51)) and (inputs(170));
    layer0_outputs(4259) <= not(inputs(194));
    layer0_outputs(4260) <= inputs(228);
    layer0_outputs(4261) <= (inputs(57)) or (inputs(238));
    layer0_outputs(4262) <= (inputs(212)) and not (inputs(54));
    layer0_outputs(4263) <= not(inputs(163));
    layer0_outputs(4264) <= not(inputs(139)) or (inputs(63));
    layer0_outputs(4265) <= not(inputs(136)) or (inputs(252));
    layer0_outputs(4266) <= (inputs(230)) and not (inputs(106));
    layer0_outputs(4267) <= not(inputs(19));
    layer0_outputs(4268) <= (inputs(75)) and not (inputs(142));
    layer0_outputs(4269) <= not(inputs(110));
    layer0_outputs(4270) <= not(inputs(179));
    layer0_outputs(4271) <= not(inputs(97));
    layer0_outputs(4272) <= inputs(186);
    layer0_outputs(4273) <= inputs(98);
    layer0_outputs(4274) <= (inputs(90)) and not (inputs(96));
    layer0_outputs(4275) <= not(inputs(3));
    layer0_outputs(4276) <= (inputs(84)) and not (inputs(136));
    layer0_outputs(4277) <= (inputs(83)) and (inputs(239));
    layer0_outputs(4278) <= not(inputs(133)) or (inputs(108));
    layer0_outputs(4279) <= not(inputs(119));
    layer0_outputs(4280) <= not(inputs(94));
    layer0_outputs(4281) <= (inputs(154)) or (inputs(155));
    layer0_outputs(4282) <= not(inputs(1));
    layer0_outputs(4283) <= not((inputs(28)) or (inputs(0)));
    layer0_outputs(4284) <= not((inputs(206)) or (inputs(219)));
    layer0_outputs(4285) <= not(inputs(192)) or (inputs(141));
    layer0_outputs(4286) <= '0';
    layer0_outputs(4287) <= not(inputs(246)) or (inputs(206));
    layer0_outputs(4288) <= not(inputs(196));
    layer0_outputs(4289) <= not(inputs(156));
    layer0_outputs(4290) <= (inputs(142)) or (inputs(163));
    layer0_outputs(4291) <= '1';
    layer0_outputs(4292) <= inputs(121);
    layer0_outputs(4293) <= not(inputs(47)) or (inputs(102));
    layer0_outputs(4294) <= inputs(22);
    layer0_outputs(4295) <= not((inputs(51)) or (inputs(25)));
    layer0_outputs(4296) <= not(inputs(202)) or (inputs(36));
    layer0_outputs(4297) <= inputs(225);
    layer0_outputs(4298) <= (inputs(255)) and not (inputs(232));
    layer0_outputs(4299) <= not(inputs(143));
    layer0_outputs(4300) <= not(inputs(211));
    layer0_outputs(4301) <= (inputs(206)) or (inputs(228));
    layer0_outputs(4302) <= '0';
    layer0_outputs(4303) <= inputs(83);
    layer0_outputs(4304) <= (inputs(233)) and (inputs(31));
    layer0_outputs(4305) <= not(inputs(132));
    layer0_outputs(4306) <= not(inputs(37));
    layer0_outputs(4307) <= inputs(254);
    layer0_outputs(4308) <= inputs(128);
    layer0_outputs(4309) <= inputs(89);
    layer0_outputs(4310) <= not((inputs(4)) xor (inputs(101)));
    layer0_outputs(4311) <= '1';
    layer0_outputs(4312) <= not((inputs(13)) or (inputs(226)));
    layer0_outputs(4313) <= (inputs(98)) or (inputs(124));
    layer0_outputs(4314) <= (inputs(43)) or (inputs(76));
    layer0_outputs(4315) <= not(inputs(104)) or (inputs(250));
    layer0_outputs(4316) <= not(inputs(198));
    layer0_outputs(4317) <= not(inputs(51));
    layer0_outputs(4318) <= not(inputs(72));
    layer0_outputs(4319) <= not((inputs(130)) or (inputs(14)));
    layer0_outputs(4320) <= '1';
    layer0_outputs(4321) <= not(inputs(73)) or (inputs(254));
    layer0_outputs(4322) <= not(inputs(168)) or (inputs(207));
    layer0_outputs(4323) <= '1';
    layer0_outputs(4324) <= inputs(182);
    layer0_outputs(4325) <= not((inputs(7)) xor (inputs(227)));
    layer0_outputs(4326) <= not((inputs(34)) or (inputs(36)));
    layer0_outputs(4327) <= not(inputs(97));
    layer0_outputs(4328) <= not(inputs(49)) or (inputs(15));
    layer0_outputs(4329) <= inputs(250);
    layer0_outputs(4330) <= not(inputs(5));
    layer0_outputs(4331) <= (inputs(245)) and not (inputs(207));
    layer0_outputs(4332) <= not((inputs(41)) and (inputs(206)));
    layer0_outputs(4333) <= not(inputs(251)) or (inputs(193));
    layer0_outputs(4334) <= inputs(166);
    layer0_outputs(4335) <= inputs(168);
    layer0_outputs(4336) <= (inputs(3)) xor (inputs(90));
    layer0_outputs(4337) <= inputs(195);
    layer0_outputs(4338) <= (inputs(99)) or (inputs(115));
    layer0_outputs(4339) <= not(inputs(118));
    layer0_outputs(4340) <= (inputs(122)) xor (inputs(124));
    layer0_outputs(4341) <= not((inputs(33)) or (inputs(58)));
    layer0_outputs(4342) <= not(inputs(193));
    layer0_outputs(4343) <= (inputs(172)) and not (inputs(14));
    layer0_outputs(4344) <= '0';
    layer0_outputs(4345) <= inputs(223);
    layer0_outputs(4346) <= not((inputs(2)) xor (inputs(43)));
    layer0_outputs(4347) <= (inputs(20)) or (inputs(219));
    layer0_outputs(4348) <= (inputs(171)) and not (inputs(34));
    layer0_outputs(4349) <= not(inputs(13)) or (inputs(12));
    layer0_outputs(4350) <= not((inputs(131)) or (inputs(125)));
    layer0_outputs(4351) <= not(inputs(38));
    layer0_outputs(4352) <= not(inputs(108));
    layer0_outputs(4353) <= not(inputs(61));
    layer0_outputs(4354) <= not(inputs(120)) or (inputs(97));
    layer0_outputs(4355) <= not((inputs(227)) xor (inputs(175)));
    layer0_outputs(4356) <= not(inputs(113));
    layer0_outputs(4357) <= not(inputs(102));
    layer0_outputs(4358) <= inputs(3);
    layer0_outputs(4359) <= (inputs(32)) xor (inputs(78));
    layer0_outputs(4360) <= inputs(192);
    layer0_outputs(4361) <= (inputs(36)) or (inputs(237));
    layer0_outputs(4362) <= not(inputs(144)) or (inputs(198));
    layer0_outputs(4363) <= not((inputs(227)) or (inputs(185)));
    layer0_outputs(4364) <= inputs(80);
    layer0_outputs(4365) <= not((inputs(148)) xor (inputs(97)));
    layer0_outputs(4366) <= not(inputs(118)) or (inputs(111));
    layer0_outputs(4367) <= not(inputs(62));
    layer0_outputs(4368) <= (inputs(198)) or (inputs(207));
    layer0_outputs(4369) <= not(inputs(113));
    layer0_outputs(4370) <= not((inputs(100)) or (inputs(115)));
    layer0_outputs(4371) <= '1';
    layer0_outputs(4372) <= (inputs(166)) or (inputs(135));
    layer0_outputs(4373) <= (inputs(163)) and (inputs(196));
    layer0_outputs(4374) <= inputs(213);
    layer0_outputs(4375) <= not(inputs(147));
    layer0_outputs(4376) <= (inputs(36)) and not (inputs(222));
    layer0_outputs(4377) <= not(inputs(85));
    layer0_outputs(4378) <= (inputs(214)) or (inputs(112));
    layer0_outputs(4379) <= (inputs(39)) and (inputs(109));
    layer0_outputs(4380) <= (inputs(230)) or (inputs(203));
    layer0_outputs(4381) <= inputs(79);
    layer0_outputs(4382) <= not(inputs(59));
    layer0_outputs(4383) <= not((inputs(204)) and (inputs(147)));
    layer0_outputs(4384) <= (inputs(196)) xor (inputs(143));
    layer0_outputs(4385) <= not(inputs(143)) or (inputs(134));
    layer0_outputs(4386) <= not((inputs(91)) and (inputs(135)));
    layer0_outputs(4387) <= not((inputs(7)) xor (inputs(106)));
    layer0_outputs(4388) <= (inputs(124)) and (inputs(96));
    layer0_outputs(4389) <= not((inputs(135)) or (inputs(220)));
    layer0_outputs(4390) <= (inputs(226)) and not (inputs(81));
    layer0_outputs(4391) <= not(inputs(168)) or (inputs(0));
    layer0_outputs(4392) <= not((inputs(167)) or (inputs(165)));
    layer0_outputs(4393) <= (inputs(53)) or (inputs(83));
    layer0_outputs(4394) <= not((inputs(200)) or (inputs(240)));
    layer0_outputs(4395) <= '0';
    layer0_outputs(4396) <= not(inputs(157));
    layer0_outputs(4397) <= '1';
    layer0_outputs(4398) <= not((inputs(246)) or (inputs(114)));
    layer0_outputs(4399) <= not(inputs(88));
    layer0_outputs(4400) <= not(inputs(40)) or (inputs(177));
    layer0_outputs(4401) <= (inputs(234)) or (inputs(250));
    layer0_outputs(4402) <= (inputs(123)) or (inputs(65));
    layer0_outputs(4403) <= (inputs(140)) and not (inputs(136));
    layer0_outputs(4404) <= (inputs(79)) and not (inputs(224));
    layer0_outputs(4405) <= inputs(197);
    layer0_outputs(4406) <= not(inputs(102)) or (inputs(169));
    layer0_outputs(4407) <= (inputs(107)) and not (inputs(29));
    layer0_outputs(4408) <= inputs(155);
    layer0_outputs(4409) <= not((inputs(61)) or (inputs(197)));
    layer0_outputs(4410) <= (inputs(187)) and not (inputs(32));
    layer0_outputs(4411) <= not((inputs(133)) or (inputs(202)));
    layer0_outputs(4412) <= (inputs(224)) and (inputs(109));
    layer0_outputs(4413) <= not(inputs(189));
    layer0_outputs(4414) <= '1';
    layer0_outputs(4415) <= inputs(18);
    layer0_outputs(4416) <= not(inputs(193)) or (inputs(138));
    layer0_outputs(4417) <= not((inputs(216)) and (inputs(205)));
    layer0_outputs(4418) <= (inputs(97)) or (inputs(23));
    layer0_outputs(4419) <= not((inputs(91)) or (inputs(38)));
    layer0_outputs(4420) <= inputs(114);
    layer0_outputs(4421) <= (inputs(99)) and (inputs(170));
    layer0_outputs(4422) <= inputs(128);
    layer0_outputs(4423) <= not((inputs(41)) xor (inputs(73)));
    layer0_outputs(4424) <= not(inputs(84)) or (inputs(223));
    layer0_outputs(4425) <= not(inputs(146)) or (inputs(21));
    layer0_outputs(4426) <= not(inputs(120));
    layer0_outputs(4427) <= '0';
    layer0_outputs(4428) <= not(inputs(132)) or (inputs(39));
    layer0_outputs(4429) <= not(inputs(212));
    layer0_outputs(4430) <= not((inputs(233)) or (inputs(64)));
    layer0_outputs(4431) <= inputs(205);
    layer0_outputs(4432) <= (inputs(212)) and (inputs(108));
    layer0_outputs(4433) <= not(inputs(44));
    layer0_outputs(4434) <= not((inputs(209)) or (inputs(114)));
    layer0_outputs(4435) <= not((inputs(152)) or (inputs(150)));
    layer0_outputs(4436) <= inputs(117);
    layer0_outputs(4437) <= inputs(209);
    layer0_outputs(4438) <= not(inputs(56));
    layer0_outputs(4439) <= '0';
    layer0_outputs(4440) <= (inputs(99)) and not (inputs(57));
    layer0_outputs(4441) <= not(inputs(146)) or (inputs(80));
    layer0_outputs(4442) <= '1';
    layer0_outputs(4443) <= (inputs(227)) and not (inputs(98));
    layer0_outputs(4444) <= not(inputs(185)) or (inputs(133));
    layer0_outputs(4445) <= (inputs(71)) and (inputs(20));
    layer0_outputs(4446) <= inputs(159);
    layer0_outputs(4447) <= '0';
    layer0_outputs(4448) <= not(inputs(247)) or (inputs(49));
    layer0_outputs(4449) <= (inputs(78)) and not (inputs(212));
    layer0_outputs(4450) <= not(inputs(151));
    layer0_outputs(4451) <= not((inputs(100)) or (inputs(4)));
    layer0_outputs(4452) <= not(inputs(174));
    layer0_outputs(4453) <= (inputs(202)) and (inputs(151));
    layer0_outputs(4454) <= not(inputs(126));
    layer0_outputs(4455) <= inputs(167);
    layer0_outputs(4456) <= inputs(99);
    layer0_outputs(4457) <= inputs(94);
    layer0_outputs(4458) <= not(inputs(175)) or (inputs(129));
    layer0_outputs(4459) <= (inputs(182)) or (inputs(150));
    layer0_outputs(4460) <= inputs(126);
    layer0_outputs(4461) <= not(inputs(6)) or (inputs(173));
    layer0_outputs(4462) <= (inputs(155)) and not (inputs(201));
    layer0_outputs(4463) <= not((inputs(196)) or (inputs(220)));
    layer0_outputs(4464) <= not(inputs(109)) or (inputs(6));
    layer0_outputs(4465) <= not(inputs(116));
    layer0_outputs(4466) <= not((inputs(134)) or (inputs(18)));
    layer0_outputs(4467) <= not((inputs(135)) and (inputs(8)));
    layer0_outputs(4468) <= inputs(233);
    layer0_outputs(4469) <= not(inputs(216));
    layer0_outputs(4470) <= inputs(63);
    layer0_outputs(4471) <= (inputs(190)) and (inputs(86));
    layer0_outputs(4472) <= not((inputs(38)) xor (inputs(145)));
    layer0_outputs(4473) <= (inputs(19)) and (inputs(11));
    layer0_outputs(4474) <= (inputs(243)) or (inputs(234));
    layer0_outputs(4475) <= (inputs(232)) or (inputs(160));
    layer0_outputs(4476) <= inputs(107);
    layer0_outputs(4477) <= '1';
    layer0_outputs(4478) <= (inputs(241)) or (inputs(191));
    layer0_outputs(4479) <= not(inputs(10));
    layer0_outputs(4480) <= not(inputs(14));
    layer0_outputs(4481) <= (inputs(90)) xor (inputs(40));
    layer0_outputs(4482) <= inputs(26);
    layer0_outputs(4483) <= not(inputs(84));
    layer0_outputs(4484) <= not(inputs(212));
    layer0_outputs(4485) <= (inputs(239)) xor (inputs(28));
    layer0_outputs(4486) <= not(inputs(130));
    layer0_outputs(4487) <= (inputs(38)) and (inputs(39));
    layer0_outputs(4488) <= '1';
    layer0_outputs(4489) <= (inputs(135)) and not (inputs(38));
    layer0_outputs(4490) <= not(inputs(127));
    layer0_outputs(4491) <= not(inputs(105));
    layer0_outputs(4492) <= inputs(186);
    layer0_outputs(4493) <= (inputs(57)) and (inputs(82));
    layer0_outputs(4494) <= not(inputs(169));
    layer0_outputs(4495) <= inputs(30);
    layer0_outputs(4496) <= (inputs(150)) or (inputs(39));
    layer0_outputs(4497) <= not(inputs(246));
    layer0_outputs(4498) <= '1';
    layer0_outputs(4499) <= '0';
    layer0_outputs(4500) <= not((inputs(160)) or (inputs(231)));
    layer0_outputs(4501) <= not(inputs(213));
    layer0_outputs(4502) <= not(inputs(230));
    layer0_outputs(4503) <= not(inputs(197));
    layer0_outputs(4504) <= not((inputs(228)) xor (inputs(208)));
    layer0_outputs(4505) <= inputs(122);
    layer0_outputs(4506) <= not((inputs(103)) or (inputs(195)));
    layer0_outputs(4507) <= (inputs(60)) and not (inputs(182));
    layer0_outputs(4508) <= inputs(121);
    layer0_outputs(4509) <= inputs(217);
    layer0_outputs(4510) <= not(inputs(50));
    layer0_outputs(4511) <= not(inputs(226)) or (inputs(27));
    layer0_outputs(4512) <= not((inputs(24)) or (inputs(34)));
    layer0_outputs(4513) <= (inputs(235)) and not (inputs(51));
    layer0_outputs(4514) <= '0';
    layer0_outputs(4515) <= inputs(114);
    layer0_outputs(4516) <= not((inputs(235)) and (inputs(223)));
    layer0_outputs(4517) <= not(inputs(254)) or (inputs(253));
    layer0_outputs(4518) <= not(inputs(83)) or (inputs(93));
    layer0_outputs(4519) <= not((inputs(206)) xor (inputs(208)));
    layer0_outputs(4520) <= not(inputs(157));
    layer0_outputs(4521) <= not(inputs(122)) or (inputs(15));
    layer0_outputs(4522) <= not((inputs(245)) and (inputs(91)));
    layer0_outputs(4523) <= (inputs(25)) and not (inputs(185));
    layer0_outputs(4524) <= not(inputs(242)) or (inputs(229));
    layer0_outputs(4525) <= (inputs(83)) xor (inputs(200));
    layer0_outputs(4526) <= (inputs(162)) xor (inputs(219));
    layer0_outputs(4527) <= (inputs(209)) and not (inputs(29));
    layer0_outputs(4528) <= not((inputs(174)) xor (inputs(234)));
    layer0_outputs(4529) <= not(inputs(209));
    layer0_outputs(4530) <= '1';
    layer0_outputs(4531) <= not((inputs(255)) xor (inputs(104)));
    layer0_outputs(4532) <= (inputs(8)) and (inputs(133));
    layer0_outputs(4533) <= not((inputs(185)) xor (inputs(239)));
    layer0_outputs(4534) <= not(inputs(164));
    layer0_outputs(4535) <= not(inputs(182));
    layer0_outputs(4536) <= not(inputs(234));
    layer0_outputs(4537) <= (inputs(239)) or (inputs(16));
    layer0_outputs(4538) <= (inputs(69)) xor (inputs(7));
    layer0_outputs(4539) <= not(inputs(7)) or (inputs(147));
    layer0_outputs(4540) <= inputs(180);
    layer0_outputs(4541) <= (inputs(70)) or (inputs(40));
    layer0_outputs(4542) <= not((inputs(240)) and (inputs(137)));
    layer0_outputs(4543) <= inputs(70);
    layer0_outputs(4544) <= (inputs(134)) and not (inputs(120));
    layer0_outputs(4545) <= not((inputs(36)) and (inputs(53)));
    layer0_outputs(4546) <= not((inputs(148)) and (inputs(16)));
    layer0_outputs(4547) <= inputs(149);
    layer0_outputs(4548) <= (inputs(44)) or (inputs(154));
    layer0_outputs(4549) <= not((inputs(162)) and (inputs(138)));
    layer0_outputs(4550) <= (inputs(247)) or (inputs(40));
    layer0_outputs(4551) <= (inputs(180)) and not (inputs(27));
    layer0_outputs(4552) <= not(inputs(0)) or (inputs(186));
    layer0_outputs(4553) <= not(inputs(15));
    layer0_outputs(4554) <= (inputs(81)) xor (inputs(139));
    layer0_outputs(4555) <= inputs(130);
    layer0_outputs(4556) <= not((inputs(5)) or (inputs(134)));
    layer0_outputs(4557) <= not(inputs(73));
    layer0_outputs(4558) <= not(inputs(227));
    layer0_outputs(4559) <= inputs(153);
    layer0_outputs(4560) <= inputs(237);
    layer0_outputs(4561) <= inputs(124);
    layer0_outputs(4562) <= not(inputs(153));
    layer0_outputs(4563) <= not(inputs(182));
    layer0_outputs(4564) <= not(inputs(202));
    layer0_outputs(4565) <= inputs(151);
    layer0_outputs(4566) <= '0';
    layer0_outputs(4567) <= not(inputs(54)) or (inputs(27));
    layer0_outputs(4568) <= not((inputs(48)) or (inputs(8)));
    layer0_outputs(4569) <= not(inputs(97));
    layer0_outputs(4570) <= not((inputs(197)) or (inputs(78)));
    layer0_outputs(4571) <= not(inputs(244));
    layer0_outputs(4572) <= '0';
    layer0_outputs(4573) <= not(inputs(153));
    layer0_outputs(4574) <= not(inputs(19));
    layer0_outputs(4575) <= inputs(204);
    layer0_outputs(4576) <= (inputs(94)) or (inputs(198));
    layer0_outputs(4577) <= '1';
    layer0_outputs(4578) <= (inputs(23)) and (inputs(74));
    layer0_outputs(4579) <= not(inputs(185)) or (inputs(100));
    layer0_outputs(4580) <= not(inputs(30)) or (inputs(26));
    layer0_outputs(4581) <= (inputs(18)) or (inputs(31));
    layer0_outputs(4582) <= (inputs(11)) or (inputs(44));
    layer0_outputs(4583) <= not(inputs(97));
    layer0_outputs(4584) <= not((inputs(112)) or (inputs(54)));
    layer0_outputs(4585) <= not(inputs(42));
    layer0_outputs(4586) <= not(inputs(24));
    layer0_outputs(4587) <= (inputs(167)) and not (inputs(154));
    layer0_outputs(4588) <= (inputs(106)) and not (inputs(248));
    layer0_outputs(4589) <= not(inputs(92)) or (inputs(219));
    layer0_outputs(4590) <= not((inputs(98)) or (inputs(31)));
    layer0_outputs(4591) <= inputs(117);
    layer0_outputs(4592) <= not(inputs(84));
    layer0_outputs(4593) <= inputs(208);
    layer0_outputs(4594) <= not((inputs(80)) xor (inputs(235)));
    layer0_outputs(4595) <= not(inputs(101));
    layer0_outputs(4596) <= (inputs(120)) and not (inputs(129));
    layer0_outputs(4597) <= inputs(121);
    layer0_outputs(4598) <= not((inputs(18)) or (inputs(41)));
    layer0_outputs(4599) <= not(inputs(209));
    layer0_outputs(4600) <= (inputs(11)) and (inputs(243));
    layer0_outputs(4601) <= not(inputs(156)) or (inputs(96));
    layer0_outputs(4602) <= not(inputs(120));
    layer0_outputs(4603) <= not(inputs(195)) or (inputs(28));
    layer0_outputs(4604) <= inputs(18);
    layer0_outputs(4605) <= not(inputs(101));
    layer0_outputs(4606) <= '0';
    layer0_outputs(4607) <= inputs(216);
    layer0_outputs(4608) <= inputs(240);
    layer0_outputs(4609) <= (inputs(150)) and not (inputs(154));
    layer0_outputs(4610) <= (inputs(159)) and not (inputs(228));
    layer0_outputs(4611) <= (inputs(26)) and not (inputs(131));
    layer0_outputs(4612) <= not((inputs(82)) or (inputs(168)));
    layer0_outputs(4613) <= '1';
    layer0_outputs(4614) <= (inputs(232)) and not (inputs(109));
    layer0_outputs(4615) <= '0';
    layer0_outputs(4616) <= not((inputs(182)) or (inputs(148)));
    layer0_outputs(4617) <= (inputs(218)) and not (inputs(29));
    layer0_outputs(4618) <= not((inputs(194)) or (inputs(165)));
    layer0_outputs(4619) <= inputs(127);
    layer0_outputs(4620) <= not(inputs(184)) or (inputs(245));
    layer0_outputs(4621) <= (inputs(191)) or (inputs(254));
    layer0_outputs(4622) <= '1';
    layer0_outputs(4623) <= not(inputs(79)) or (inputs(96));
    layer0_outputs(4624) <= not((inputs(34)) xor (inputs(52)));
    layer0_outputs(4625) <= (inputs(75)) or (inputs(142));
    layer0_outputs(4626) <= (inputs(207)) or (inputs(192));
    layer0_outputs(4627) <= not(inputs(101));
    layer0_outputs(4628) <= inputs(113);
    layer0_outputs(4629) <= not(inputs(100));
    layer0_outputs(4630) <= (inputs(215)) and (inputs(18));
    layer0_outputs(4631) <= not(inputs(193)) or (inputs(158));
    layer0_outputs(4632) <= '1';
    layer0_outputs(4633) <= (inputs(174)) and not (inputs(13));
    layer0_outputs(4634) <= (inputs(152)) or (inputs(71));
    layer0_outputs(4635) <= not((inputs(246)) and (inputs(148)));
    layer0_outputs(4636) <= not((inputs(100)) or (inputs(84)));
    layer0_outputs(4637) <= not(inputs(136)) or (inputs(91));
    layer0_outputs(4638) <= not(inputs(35));
    layer0_outputs(4639) <= not((inputs(62)) and (inputs(201)));
    layer0_outputs(4640) <= inputs(182);
    layer0_outputs(4641) <= inputs(98);
    layer0_outputs(4642) <= not((inputs(55)) xor (inputs(50)));
    layer0_outputs(4643) <= (inputs(21)) or (inputs(43));
    layer0_outputs(4644) <= not((inputs(90)) or (inputs(59)));
    layer0_outputs(4645) <= not(inputs(119)) or (inputs(236));
    layer0_outputs(4646) <= not(inputs(145)) or (inputs(6));
    layer0_outputs(4647) <= inputs(198);
    layer0_outputs(4648) <= (inputs(52)) and not (inputs(201));
    layer0_outputs(4649) <= not(inputs(56)) or (inputs(35));
    layer0_outputs(4650) <= not(inputs(216));
    layer0_outputs(4651) <= not(inputs(172)) or (inputs(137));
    layer0_outputs(4652) <= not(inputs(253));
    layer0_outputs(4653) <= not((inputs(208)) and (inputs(113)));
    layer0_outputs(4654) <= not((inputs(94)) or (inputs(149)));
    layer0_outputs(4655) <= not(inputs(31));
    layer0_outputs(4656) <= '0';
    layer0_outputs(4657) <= (inputs(252)) or (inputs(10));
    layer0_outputs(4658) <= (inputs(137)) and not (inputs(54));
    layer0_outputs(4659) <= (inputs(167)) xor (inputs(92));
    layer0_outputs(4660) <= not(inputs(139));
    layer0_outputs(4661) <= not(inputs(88)) or (inputs(196));
    layer0_outputs(4662) <= inputs(113);
    layer0_outputs(4663) <= not(inputs(184));
    layer0_outputs(4664) <= inputs(42);
    layer0_outputs(4665) <= (inputs(183)) and (inputs(220));
    layer0_outputs(4666) <= not((inputs(79)) and (inputs(192)));
    layer0_outputs(4667) <= not(inputs(64)) or (inputs(55));
    layer0_outputs(4668) <= (inputs(110)) and not (inputs(221));
    layer0_outputs(4669) <= '0';
    layer0_outputs(4670) <= '1';
    layer0_outputs(4671) <= inputs(163);
    layer0_outputs(4672) <= not((inputs(94)) or (inputs(149)));
    layer0_outputs(4673) <= (inputs(83)) and (inputs(96));
    layer0_outputs(4674) <= inputs(137);
    layer0_outputs(4675) <= '1';
    layer0_outputs(4676) <= inputs(225);
    layer0_outputs(4677) <= (inputs(151)) or (inputs(133));
    layer0_outputs(4678) <= not((inputs(14)) or (inputs(144)));
    layer0_outputs(4679) <= '0';
    layer0_outputs(4680) <= not(inputs(108));
    layer0_outputs(4681) <= not(inputs(72));
    layer0_outputs(4682) <= inputs(83);
    layer0_outputs(4683) <= not(inputs(219));
    layer0_outputs(4684) <= not((inputs(8)) and (inputs(74)));
    layer0_outputs(4685) <= '0';
    layer0_outputs(4686) <= not(inputs(118)) or (inputs(60));
    layer0_outputs(4687) <= not((inputs(246)) or (inputs(113)));
    layer0_outputs(4688) <= not(inputs(81));
    layer0_outputs(4689) <= not(inputs(246)) or (inputs(187));
    layer0_outputs(4690) <= not((inputs(220)) or (inputs(191)));
    layer0_outputs(4691) <= (inputs(72)) or (inputs(97));
    layer0_outputs(4692) <= not(inputs(206));
    layer0_outputs(4693) <= '0';
    layer0_outputs(4694) <= not((inputs(245)) and (inputs(203)));
    layer0_outputs(4695) <= '1';
    layer0_outputs(4696) <= '1';
    layer0_outputs(4697) <= not(inputs(236));
    layer0_outputs(4698) <= not((inputs(154)) or (inputs(169)));
    layer0_outputs(4699) <= inputs(70);
    layer0_outputs(4700) <= '1';
    layer0_outputs(4701) <= not(inputs(135));
    layer0_outputs(4702) <= '0';
    layer0_outputs(4703) <= inputs(204);
    layer0_outputs(4704) <= not(inputs(52));
    layer0_outputs(4705) <= '0';
    layer0_outputs(4706) <= not(inputs(166));
    layer0_outputs(4707) <= (inputs(115)) and not (inputs(4));
    layer0_outputs(4708) <= not(inputs(12));
    layer0_outputs(4709) <= inputs(15);
    layer0_outputs(4710) <= (inputs(32)) and not (inputs(95));
    layer0_outputs(4711) <= (inputs(127)) and not (inputs(89));
    layer0_outputs(4712) <= not((inputs(65)) xor (inputs(229)));
    layer0_outputs(4713) <= not((inputs(132)) and (inputs(38)));
    layer0_outputs(4714) <= not((inputs(203)) and (inputs(103)));
    layer0_outputs(4715) <= inputs(227);
    layer0_outputs(4716) <= not(inputs(176));
    layer0_outputs(4717) <= not((inputs(16)) or (inputs(117)));
    layer0_outputs(4718) <= not(inputs(150)) or (inputs(246));
    layer0_outputs(4719) <= not((inputs(161)) xor (inputs(116)));
    layer0_outputs(4720) <= inputs(240);
    layer0_outputs(4721) <= (inputs(151)) and not (inputs(38));
    layer0_outputs(4722) <= inputs(230);
    layer0_outputs(4723) <= not(inputs(61)) or (inputs(147));
    layer0_outputs(4724) <= (inputs(247)) and not (inputs(209));
    layer0_outputs(4725) <= (inputs(145)) or (inputs(113));
    layer0_outputs(4726) <= (inputs(151)) or (inputs(226));
    layer0_outputs(4727) <= not(inputs(202));
    layer0_outputs(4728) <= not(inputs(144));
    layer0_outputs(4729) <= not(inputs(203)) or (inputs(76));
    layer0_outputs(4730) <= not(inputs(89)) or (inputs(204));
    layer0_outputs(4731) <= (inputs(58)) or (inputs(153));
    layer0_outputs(4732) <= not(inputs(224)) or (inputs(59));
    layer0_outputs(4733) <= '1';
    layer0_outputs(4734) <= not((inputs(106)) or (inputs(63)));
    layer0_outputs(4735) <= not((inputs(98)) or (inputs(11)));
    layer0_outputs(4736) <= not(inputs(101));
    layer0_outputs(4737) <= not((inputs(128)) xor (inputs(131)));
    layer0_outputs(4738) <= (inputs(164)) or (inputs(111));
    layer0_outputs(4739) <= (inputs(94)) xor (inputs(171));
    layer0_outputs(4740) <= (inputs(93)) and not (inputs(134));
    layer0_outputs(4741) <= not(inputs(8));
    layer0_outputs(4742) <= '0';
    layer0_outputs(4743) <= not(inputs(58)) or (inputs(115));
    layer0_outputs(4744) <= (inputs(163)) or (inputs(37));
    layer0_outputs(4745) <= not(inputs(223)) or (inputs(25));
    layer0_outputs(4746) <= not(inputs(106));
    layer0_outputs(4747) <= not(inputs(230));
    layer0_outputs(4748) <= not(inputs(71)) or (inputs(36));
    layer0_outputs(4749) <= inputs(183);
    layer0_outputs(4750) <= not(inputs(64)) or (inputs(39));
    layer0_outputs(4751) <= not(inputs(151));
    layer0_outputs(4752) <= not((inputs(80)) xor (inputs(48)));
    layer0_outputs(4753) <= not((inputs(103)) xor (inputs(128)));
    layer0_outputs(4754) <= not((inputs(21)) and (inputs(215)));
    layer0_outputs(4755) <= (inputs(6)) xor (inputs(192));
    layer0_outputs(4756) <= not(inputs(107)) or (inputs(51));
    layer0_outputs(4757) <= not(inputs(163));
    layer0_outputs(4758) <= not((inputs(140)) or (inputs(63)));
    layer0_outputs(4759) <= not(inputs(100)) or (inputs(3));
    layer0_outputs(4760) <= (inputs(182)) or (inputs(253));
    layer0_outputs(4761) <= not(inputs(179)) or (inputs(80));
    layer0_outputs(4762) <= not(inputs(85));
    layer0_outputs(4763) <= inputs(136);
    layer0_outputs(4764) <= not(inputs(213)) or (inputs(38));
    layer0_outputs(4765) <= (inputs(225)) xor (inputs(158));
    layer0_outputs(4766) <= '1';
    layer0_outputs(4767) <= not(inputs(56)) or (inputs(105));
    layer0_outputs(4768) <= '0';
    layer0_outputs(4769) <= not(inputs(16));
    layer0_outputs(4770) <= '0';
    layer0_outputs(4771) <= (inputs(147)) and not (inputs(224));
    layer0_outputs(4772) <= not((inputs(73)) xor (inputs(105)));
    layer0_outputs(4773) <= not(inputs(54));
    layer0_outputs(4774) <= (inputs(26)) or (inputs(61));
    layer0_outputs(4775) <= '1';
    layer0_outputs(4776) <= not(inputs(23)) or (inputs(85));
    layer0_outputs(4777) <= not((inputs(194)) and (inputs(188)));
    layer0_outputs(4778) <= (inputs(205)) and not (inputs(10));
    layer0_outputs(4779) <= not(inputs(97));
    layer0_outputs(4780) <= (inputs(107)) or (inputs(241));
    layer0_outputs(4781) <= (inputs(117)) and (inputs(128));
    layer0_outputs(4782) <= not((inputs(223)) or (inputs(97)));
    layer0_outputs(4783) <= not(inputs(176));
    layer0_outputs(4784) <= not(inputs(223)) or (inputs(251));
    layer0_outputs(4785) <= inputs(86);
    layer0_outputs(4786) <= not(inputs(170)) or (inputs(154));
    layer0_outputs(4787) <= not(inputs(182)) or (inputs(78));
    layer0_outputs(4788) <= not(inputs(94));
    layer0_outputs(4789) <= (inputs(159)) xor (inputs(69));
    layer0_outputs(4790) <= '1';
    layer0_outputs(4791) <= not(inputs(242));
    layer0_outputs(4792) <= inputs(103);
    layer0_outputs(4793) <= not(inputs(130)) or (inputs(12));
    layer0_outputs(4794) <= not(inputs(75)) or (inputs(197));
    layer0_outputs(4795) <= not((inputs(25)) and (inputs(165)));
    layer0_outputs(4796) <= not(inputs(229));
    layer0_outputs(4797) <= not((inputs(80)) or (inputs(116)));
    layer0_outputs(4798) <= not(inputs(127));
    layer0_outputs(4799) <= not((inputs(209)) and (inputs(54)));
    layer0_outputs(4800) <= inputs(6);
    layer0_outputs(4801) <= not(inputs(117)) or (inputs(8));
    layer0_outputs(4802) <= not((inputs(4)) xor (inputs(39)));
    layer0_outputs(4803) <= not((inputs(177)) or (inputs(7)));
    layer0_outputs(4804) <= not(inputs(170));
    layer0_outputs(4805) <= not((inputs(173)) or (inputs(56)));
    layer0_outputs(4806) <= not(inputs(83));
    layer0_outputs(4807) <= (inputs(244)) and (inputs(25));
    layer0_outputs(4808) <= '1';
    layer0_outputs(4809) <= (inputs(239)) and (inputs(217));
    layer0_outputs(4810) <= inputs(168);
    layer0_outputs(4811) <= inputs(112);
    layer0_outputs(4812) <= inputs(21);
    layer0_outputs(4813) <= not(inputs(63)) or (inputs(124));
    layer0_outputs(4814) <= not(inputs(7)) or (inputs(163));
    layer0_outputs(4815) <= (inputs(155)) or (inputs(111));
    layer0_outputs(4816) <= '1';
    layer0_outputs(4817) <= (inputs(11)) and (inputs(238));
    layer0_outputs(4818) <= not((inputs(152)) or (inputs(75)));
    layer0_outputs(4819) <= not(inputs(127));
    layer0_outputs(4820) <= not(inputs(91)) or (inputs(152));
    layer0_outputs(4821) <= inputs(14);
    layer0_outputs(4822) <= '0';
    layer0_outputs(4823) <= not(inputs(99));
    layer0_outputs(4824) <= not(inputs(189)) or (inputs(214));
    layer0_outputs(4825) <= (inputs(167)) or (inputs(83));
    layer0_outputs(4826) <= inputs(79);
    layer0_outputs(4827) <= not(inputs(223)) or (inputs(47));
    layer0_outputs(4828) <= '0';
    layer0_outputs(4829) <= not(inputs(111));
    layer0_outputs(4830) <= not(inputs(212)) or (inputs(168));
    layer0_outputs(4831) <= (inputs(149)) and not (inputs(3));
    layer0_outputs(4832) <= not(inputs(85)) or (inputs(79));
    layer0_outputs(4833) <= (inputs(99)) and (inputs(200));
    layer0_outputs(4834) <= (inputs(95)) or (inputs(232));
    layer0_outputs(4835) <= not((inputs(46)) xor (inputs(59)));
    layer0_outputs(4836) <= not(inputs(188));
    layer0_outputs(4837) <= not(inputs(123));
    layer0_outputs(4838) <= not((inputs(252)) or (inputs(38)));
    layer0_outputs(4839) <= not(inputs(246)) or (inputs(154));
    layer0_outputs(4840) <= inputs(23);
    layer0_outputs(4841) <= inputs(62);
    layer0_outputs(4842) <= (inputs(131)) or (inputs(77));
    layer0_outputs(4843) <= (inputs(64)) or (inputs(150));
    layer0_outputs(4844) <= not((inputs(10)) or (inputs(109)));
    layer0_outputs(4845) <= not((inputs(96)) or (inputs(189)));
    layer0_outputs(4846) <= (inputs(24)) and (inputs(167));
    layer0_outputs(4847) <= not(inputs(211)) or (inputs(253));
    layer0_outputs(4848) <= not(inputs(149));
    layer0_outputs(4849) <= inputs(40);
    layer0_outputs(4850) <= inputs(161);
    layer0_outputs(4851) <= '0';
    layer0_outputs(4852) <= '0';
    layer0_outputs(4853) <= (inputs(129)) and not (inputs(250));
    layer0_outputs(4854) <= not(inputs(165));
    layer0_outputs(4855) <= inputs(8);
    layer0_outputs(4856) <= inputs(195);
    layer0_outputs(4857) <= '0';
    layer0_outputs(4858) <= not(inputs(179)) or (inputs(192));
    layer0_outputs(4859) <= not(inputs(23));
    layer0_outputs(4860) <= (inputs(124)) or (inputs(242));
    layer0_outputs(4861) <= inputs(114);
    layer0_outputs(4862) <= (inputs(232)) and not (inputs(4));
    layer0_outputs(4863) <= not(inputs(194)) or (inputs(240));
    layer0_outputs(4864) <= not((inputs(153)) or (inputs(130)));
    layer0_outputs(4865) <= not((inputs(173)) or (inputs(133)));
    layer0_outputs(4866) <= (inputs(236)) xor (inputs(206));
    layer0_outputs(4867) <= not((inputs(22)) and (inputs(52)));
    layer0_outputs(4868) <= not(inputs(211));
    layer0_outputs(4869) <= not((inputs(122)) xor (inputs(238)));
    layer0_outputs(4870) <= '0';
    layer0_outputs(4871) <= inputs(146);
    layer0_outputs(4872) <= not(inputs(21));
    layer0_outputs(4873) <= (inputs(137)) and not (inputs(150));
    layer0_outputs(4874) <= not(inputs(22));
    layer0_outputs(4875) <= not((inputs(28)) or (inputs(2)));
    layer0_outputs(4876) <= (inputs(189)) and not (inputs(247));
    layer0_outputs(4877) <= (inputs(132)) and (inputs(178));
    layer0_outputs(4878) <= inputs(19);
    layer0_outputs(4879) <= not((inputs(147)) xor (inputs(240)));
    layer0_outputs(4880) <= not(inputs(15));
    layer0_outputs(4881) <= (inputs(67)) and not (inputs(30));
    layer0_outputs(4882) <= not(inputs(130));
    layer0_outputs(4883) <= (inputs(38)) or (inputs(39));
    layer0_outputs(4884) <= inputs(183);
    layer0_outputs(4885) <= '0';
    layer0_outputs(4886) <= not(inputs(214)) or (inputs(64));
    layer0_outputs(4887) <= not((inputs(210)) or (inputs(31)));
    layer0_outputs(4888) <= not(inputs(141)) or (inputs(181));
    layer0_outputs(4889) <= inputs(99);
    layer0_outputs(4890) <= inputs(179);
    layer0_outputs(4891) <= inputs(147);
    layer0_outputs(4892) <= (inputs(247)) and not (inputs(66));
    layer0_outputs(4893) <= not((inputs(194)) and (inputs(76)));
    layer0_outputs(4894) <= (inputs(108)) or (inputs(69));
    layer0_outputs(4895) <= inputs(148);
    layer0_outputs(4896) <= inputs(115);
    layer0_outputs(4897) <= '1';
    layer0_outputs(4898) <= inputs(105);
    layer0_outputs(4899) <= not(inputs(210)) or (inputs(95));
    layer0_outputs(4900) <= not(inputs(62));
    layer0_outputs(4901) <= inputs(22);
    layer0_outputs(4902) <= not(inputs(132)) or (inputs(3));
    layer0_outputs(4903) <= inputs(126);
    layer0_outputs(4904) <= (inputs(231)) and not (inputs(70));
    layer0_outputs(4905) <= (inputs(131)) and not (inputs(190));
    layer0_outputs(4906) <= (inputs(188)) and not (inputs(244));
    layer0_outputs(4907) <= (inputs(232)) or (inputs(160));
    layer0_outputs(4908) <= not((inputs(94)) or (inputs(107)));
    layer0_outputs(4909) <= (inputs(158)) and not (inputs(155));
    layer0_outputs(4910) <= inputs(87);
    layer0_outputs(4911) <= inputs(110);
    layer0_outputs(4912) <= '0';
    layer0_outputs(4913) <= (inputs(180)) or (inputs(179));
    layer0_outputs(4914) <= not((inputs(85)) or (inputs(112)));
    layer0_outputs(4915) <= not(inputs(105)) or (inputs(199));
    layer0_outputs(4916) <= inputs(72);
    layer0_outputs(4917) <= (inputs(175)) and not (inputs(246));
    layer0_outputs(4918) <= not((inputs(180)) xor (inputs(129)));
    layer0_outputs(4919) <= not((inputs(103)) xor (inputs(145)));
    layer0_outputs(4920) <= (inputs(80)) and (inputs(241));
    layer0_outputs(4921) <= inputs(138);
    layer0_outputs(4922) <= inputs(144);
    layer0_outputs(4923) <= inputs(135);
    layer0_outputs(4924) <= (inputs(45)) and (inputs(120));
    layer0_outputs(4925) <= inputs(234);
    layer0_outputs(4926) <= '1';
    layer0_outputs(4927) <= (inputs(61)) xor (inputs(59));
    layer0_outputs(4928) <= (inputs(177)) and not (inputs(174));
    layer0_outputs(4929) <= inputs(23);
    layer0_outputs(4930) <= not(inputs(36)) or (inputs(255));
    layer0_outputs(4931) <= (inputs(141)) or (inputs(169));
    layer0_outputs(4932) <= inputs(211);
    layer0_outputs(4933) <= (inputs(157)) or (inputs(171));
    layer0_outputs(4934) <= not((inputs(65)) or (inputs(254)));
    layer0_outputs(4935) <= (inputs(119)) and not (inputs(209));
    layer0_outputs(4936) <= (inputs(182)) and not (inputs(92));
    layer0_outputs(4937) <= not(inputs(110));
    layer0_outputs(4938) <= inputs(141);
    layer0_outputs(4939) <= (inputs(23)) and not (inputs(78));
    layer0_outputs(4940) <= (inputs(64)) or (inputs(177));
    layer0_outputs(4941) <= not((inputs(101)) or (inputs(145)));
    layer0_outputs(4942) <= not(inputs(229));
    layer0_outputs(4943) <= not(inputs(86));
    layer0_outputs(4944) <= '1';
    layer0_outputs(4945) <= not(inputs(60)) or (inputs(137));
    layer0_outputs(4946) <= not(inputs(86)) or (inputs(255));
    layer0_outputs(4947) <= '0';
    layer0_outputs(4948) <= (inputs(186)) xor (inputs(185));
    layer0_outputs(4949) <= not(inputs(110)) or (inputs(168));
    layer0_outputs(4950) <= not(inputs(53));
    layer0_outputs(4951) <= not(inputs(92));
    layer0_outputs(4952) <= '1';
    layer0_outputs(4953) <= (inputs(81)) and (inputs(208));
    layer0_outputs(4954) <= (inputs(98)) or (inputs(31));
    layer0_outputs(4955) <= not(inputs(77));
    layer0_outputs(4956) <= (inputs(249)) xor (inputs(71));
    layer0_outputs(4957) <= not(inputs(209)) or (inputs(22));
    layer0_outputs(4958) <= not(inputs(172));
    layer0_outputs(4959) <= not(inputs(29));
    layer0_outputs(4960) <= inputs(8);
    layer0_outputs(4961) <= not(inputs(50)) or (inputs(225));
    layer0_outputs(4962) <= inputs(229);
    layer0_outputs(4963) <= '0';
    layer0_outputs(4964) <= not(inputs(138));
    layer0_outputs(4965) <= not((inputs(127)) or (inputs(189)));
    layer0_outputs(4966) <= not((inputs(147)) or (inputs(92)));
    layer0_outputs(4967) <= (inputs(188)) and not (inputs(32));
    layer0_outputs(4968) <= not((inputs(37)) or (inputs(142)));
    layer0_outputs(4969) <= inputs(145);
    layer0_outputs(4970) <= inputs(111);
    layer0_outputs(4971) <= inputs(215);
    layer0_outputs(4972) <= not(inputs(200));
    layer0_outputs(4973) <= (inputs(110)) and not (inputs(78));
    layer0_outputs(4974) <= not(inputs(77));
    layer0_outputs(4975) <= inputs(160);
    layer0_outputs(4976) <= inputs(144);
    layer0_outputs(4977) <= (inputs(202)) and (inputs(163));
    layer0_outputs(4978) <= (inputs(222)) and not (inputs(77));
    layer0_outputs(4979) <= inputs(13);
    layer0_outputs(4980) <= inputs(19);
    layer0_outputs(4981) <= '1';
    layer0_outputs(4982) <= inputs(181);
    layer0_outputs(4983) <= (inputs(241)) and (inputs(234));
    layer0_outputs(4984) <= inputs(125);
    layer0_outputs(4985) <= not((inputs(252)) and (inputs(202)));
    layer0_outputs(4986) <= (inputs(57)) and not (inputs(186));
    layer0_outputs(4987) <= not((inputs(227)) or (inputs(42)));
    layer0_outputs(4988) <= not(inputs(195)) or (inputs(108));
    layer0_outputs(4989) <= not(inputs(116));
    layer0_outputs(4990) <= '1';
    layer0_outputs(4991) <= '1';
    layer0_outputs(4992) <= not(inputs(120));
    layer0_outputs(4993) <= (inputs(70)) and not (inputs(1));
    layer0_outputs(4994) <= not(inputs(119));
    layer0_outputs(4995) <= not((inputs(195)) or (inputs(239)));
    layer0_outputs(4996) <= not((inputs(250)) and (inputs(189)));
    layer0_outputs(4997) <= not(inputs(214)) or (inputs(253));
    layer0_outputs(4998) <= not((inputs(204)) xor (inputs(42)));
    layer0_outputs(4999) <= '0';
    layer0_outputs(5000) <= (inputs(107)) and not (inputs(1));
    layer0_outputs(5001) <= not(inputs(207));
    layer0_outputs(5002) <= inputs(242);
    layer0_outputs(5003) <= inputs(196);
    layer0_outputs(5004) <= '1';
    layer0_outputs(5005) <= (inputs(130)) and not (inputs(17));
    layer0_outputs(5006) <= not((inputs(239)) or (inputs(165)));
    layer0_outputs(5007) <= not((inputs(94)) and (inputs(117)));
    layer0_outputs(5008) <= not(inputs(225));
    layer0_outputs(5009) <= not((inputs(170)) or (inputs(167)));
    layer0_outputs(5010) <= not((inputs(55)) and (inputs(203)));
    layer0_outputs(5011) <= not(inputs(195)) or (inputs(252));
    layer0_outputs(5012) <= (inputs(55)) and not (inputs(169));
    layer0_outputs(5013) <= not((inputs(115)) or (inputs(230)));
    layer0_outputs(5014) <= not((inputs(175)) and (inputs(201)));
    layer0_outputs(5015) <= inputs(118);
    layer0_outputs(5016) <= inputs(165);
    layer0_outputs(5017) <= (inputs(170)) and not (inputs(71));
    layer0_outputs(5018) <= (inputs(146)) or (inputs(108));
    layer0_outputs(5019) <= inputs(59);
    layer0_outputs(5020) <= (inputs(68)) xor (inputs(71));
    layer0_outputs(5021) <= not(inputs(238));
    layer0_outputs(5022) <= (inputs(92)) xor (inputs(51));
    layer0_outputs(5023) <= inputs(248);
    layer0_outputs(5024) <= not(inputs(177)) or (inputs(153));
    layer0_outputs(5025) <= inputs(191);
    layer0_outputs(5026) <= (inputs(34)) and not (inputs(161));
    layer0_outputs(5027) <= not(inputs(204));
    layer0_outputs(5028) <= inputs(208);
    layer0_outputs(5029) <= not((inputs(182)) xor (inputs(31)));
    layer0_outputs(5030) <= not(inputs(231));
    layer0_outputs(5031) <= '1';
    layer0_outputs(5032) <= inputs(167);
    layer0_outputs(5033) <= (inputs(139)) xor (inputs(79));
    layer0_outputs(5034) <= '0';
    layer0_outputs(5035) <= not(inputs(17)) or (inputs(238));
    layer0_outputs(5036) <= (inputs(135)) and not (inputs(5));
    layer0_outputs(5037) <= inputs(191);
    layer0_outputs(5038) <= inputs(183);
    layer0_outputs(5039) <= (inputs(204)) and not (inputs(11));
    layer0_outputs(5040) <= not(inputs(201));
    layer0_outputs(5041) <= '1';
    layer0_outputs(5042) <= (inputs(149)) and (inputs(221));
    layer0_outputs(5043) <= (inputs(18)) and not (inputs(59));
    layer0_outputs(5044) <= (inputs(138)) or (inputs(70));
    layer0_outputs(5045) <= inputs(115);
    layer0_outputs(5046) <= not(inputs(254)) or (inputs(162));
    layer0_outputs(5047) <= not(inputs(88)) or (inputs(226));
    layer0_outputs(5048) <= not(inputs(189)) or (inputs(117));
    layer0_outputs(5049) <= not(inputs(153)) or (inputs(47));
    layer0_outputs(5050) <= not((inputs(219)) or (inputs(180)));
    layer0_outputs(5051) <= not(inputs(135));
    layer0_outputs(5052) <= (inputs(36)) and (inputs(169));
    layer0_outputs(5053) <= (inputs(168)) xor (inputs(198));
    layer0_outputs(5054) <= (inputs(153)) and not (inputs(222));
    layer0_outputs(5055) <= not(inputs(197)) or (inputs(102));
    layer0_outputs(5056) <= not(inputs(49)) or (inputs(45));
    layer0_outputs(5057) <= inputs(27);
    layer0_outputs(5058) <= inputs(39);
    layer0_outputs(5059) <= not((inputs(221)) or (inputs(207)));
    layer0_outputs(5060) <= (inputs(194)) xor (inputs(210));
    layer0_outputs(5061) <= (inputs(67)) and not (inputs(40));
    layer0_outputs(5062) <= not(inputs(188)) or (inputs(215));
    layer0_outputs(5063) <= '0';
    layer0_outputs(5064) <= (inputs(170)) and not (inputs(235));
    layer0_outputs(5065) <= not(inputs(103)) or (inputs(130));
    layer0_outputs(5066) <= '0';
    layer0_outputs(5067) <= not((inputs(94)) xor (inputs(52)));
    layer0_outputs(5068) <= (inputs(28)) and not (inputs(237));
    layer0_outputs(5069) <= (inputs(82)) and not (inputs(71));
    layer0_outputs(5070) <= not(inputs(146));
    layer0_outputs(5071) <= not(inputs(50));
    layer0_outputs(5072) <= (inputs(164)) or (inputs(30));
    layer0_outputs(5073) <= (inputs(196)) xor (inputs(243));
    layer0_outputs(5074) <= '1';
    layer0_outputs(5075) <= not((inputs(41)) and (inputs(92)));
    layer0_outputs(5076) <= (inputs(202)) and not (inputs(153));
    layer0_outputs(5077) <= not(inputs(95));
    layer0_outputs(5078) <= (inputs(5)) or (inputs(35));
    layer0_outputs(5079) <= (inputs(21)) and not (inputs(130));
    layer0_outputs(5080) <= (inputs(182)) and (inputs(101));
    layer0_outputs(5081) <= (inputs(11)) xor (inputs(254));
    layer0_outputs(5082) <= not(inputs(252));
    layer0_outputs(5083) <= not((inputs(255)) or (inputs(106)));
    layer0_outputs(5084) <= '0';
    layer0_outputs(5085) <= (inputs(247)) and not (inputs(184));
    layer0_outputs(5086) <= (inputs(233)) and not (inputs(45));
    layer0_outputs(5087) <= not((inputs(23)) or (inputs(142)));
    layer0_outputs(5088) <= (inputs(18)) or (inputs(33));
    layer0_outputs(5089) <= '1';
    layer0_outputs(5090) <= '0';
    layer0_outputs(5091) <= (inputs(248)) and (inputs(196));
    layer0_outputs(5092) <= not((inputs(1)) and (inputs(52)));
    layer0_outputs(5093) <= '0';
    layer0_outputs(5094) <= not((inputs(251)) or (inputs(102)));
    layer0_outputs(5095) <= inputs(148);
    layer0_outputs(5096) <= not((inputs(44)) xor (inputs(5)));
    layer0_outputs(5097) <= not((inputs(134)) or (inputs(171)));
    layer0_outputs(5098) <= (inputs(110)) and (inputs(169));
    layer0_outputs(5099) <= '1';
    layer0_outputs(5100) <= inputs(169);
    layer0_outputs(5101) <= (inputs(81)) or (inputs(248));
    layer0_outputs(5102) <= not(inputs(26));
    layer0_outputs(5103) <= not((inputs(208)) and (inputs(143)));
    layer0_outputs(5104) <= (inputs(220)) or (inputs(176));
    layer0_outputs(5105) <= not(inputs(39));
    layer0_outputs(5106) <= not(inputs(197));
    layer0_outputs(5107) <= inputs(122);
    layer0_outputs(5108) <= not(inputs(81));
    layer0_outputs(5109) <= not(inputs(157));
    layer0_outputs(5110) <= inputs(27);
    layer0_outputs(5111) <= not(inputs(228));
    layer0_outputs(5112) <= not(inputs(167)) or (inputs(0));
    layer0_outputs(5113) <= (inputs(15)) or (inputs(128));
    layer0_outputs(5114) <= inputs(108);
    layer0_outputs(5115) <= not(inputs(8)) or (inputs(176));
    layer0_outputs(5116) <= (inputs(21)) and (inputs(90));
    layer0_outputs(5117) <= not(inputs(50));
    layer0_outputs(5118) <= not((inputs(207)) or (inputs(117)));
    layer0_outputs(5119) <= (inputs(234)) or (inputs(213));
    layer0_outputs(5120) <= (inputs(81)) or (inputs(112));
    layer0_outputs(5121) <= inputs(210);
    layer0_outputs(5122) <= inputs(47);
    layer0_outputs(5123) <= not((inputs(147)) or (inputs(1)));
    layer0_outputs(5124) <= inputs(231);
    layer0_outputs(5125) <= inputs(153);
    layer0_outputs(5126) <= (inputs(36)) or (inputs(203));
    layer0_outputs(5127) <= (inputs(137)) or (inputs(24));
    layer0_outputs(5128) <= (inputs(248)) and not (inputs(218));
    layer0_outputs(5129) <= (inputs(173)) and not (inputs(88));
    layer0_outputs(5130) <= (inputs(77)) and not (inputs(234));
    layer0_outputs(5131) <= not(inputs(59));
    layer0_outputs(5132) <= '0';
    layer0_outputs(5133) <= not(inputs(255));
    layer0_outputs(5134) <= not(inputs(164)) or (inputs(88));
    layer0_outputs(5135) <= not((inputs(90)) or (inputs(107)));
    layer0_outputs(5136) <= '1';
    layer0_outputs(5137) <= inputs(119);
    layer0_outputs(5138) <= not(inputs(76));
    layer0_outputs(5139) <= inputs(40);
    layer0_outputs(5140) <= (inputs(194)) or (inputs(144));
    layer0_outputs(5141) <= inputs(114);
    layer0_outputs(5142) <= not(inputs(203)) or (inputs(223));
    layer0_outputs(5143) <= not(inputs(31)) or (inputs(79));
    layer0_outputs(5144) <= (inputs(241)) and (inputs(226));
    layer0_outputs(5145) <= not(inputs(195)) or (inputs(81));
    layer0_outputs(5146) <= not(inputs(118)) or (inputs(15));
    layer0_outputs(5147) <= not((inputs(24)) or (inputs(190)));
    layer0_outputs(5148) <= (inputs(35)) and not (inputs(255));
    layer0_outputs(5149) <= (inputs(193)) or (inputs(189));
    layer0_outputs(5150) <= not(inputs(70));
    layer0_outputs(5151) <= (inputs(157)) or (inputs(228));
    layer0_outputs(5152) <= not(inputs(162));
    layer0_outputs(5153) <= inputs(244);
    layer0_outputs(5154) <= (inputs(204)) and (inputs(115));
    layer0_outputs(5155) <= not(inputs(86));
    layer0_outputs(5156) <= not(inputs(179)) or (inputs(20));
    layer0_outputs(5157) <= not((inputs(221)) or (inputs(194)));
    layer0_outputs(5158) <= '0';
    layer0_outputs(5159) <= not((inputs(42)) and (inputs(74)));
    layer0_outputs(5160) <= (inputs(28)) or (inputs(239));
    layer0_outputs(5161) <= (inputs(63)) xor (inputs(87));
    layer0_outputs(5162) <= '0';
    layer0_outputs(5163) <= inputs(102);
    layer0_outputs(5164) <= not(inputs(232));
    layer0_outputs(5165) <= inputs(108);
    layer0_outputs(5166) <= not(inputs(183));
    layer0_outputs(5167) <= not(inputs(55));
    layer0_outputs(5168) <= (inputs(212)) xor (inputs(209));
    layer0_outputs(5169) <= (inputs(71)) and not (inputs(1));
    layer0_outputs(5170) <= inputs(26);
    layer0_outputs(5171) <= (inputs(43)) or (inputs(32));
    layer0_outputs(5172) <= inputs(63);
    layer0_outputs(5173) <= not(inputs(188));
    layer0_outputs(5174) <= (inputs(82)) and not (inputs(32));
    layer0_outputs(5175) <= not(inputs(120));
    layer0_outputs(5176) <= inputs(58);
    layer0_outputs(5177) <= (inputs(79)) and not (inputs(46));
    layer0_outputs(5178) <= (inputs(196)) xor (inputs(228));
    layer0_outputs(5179) <= not(inputs(35)) or (inputs(147));
    layer0_outputs(5180) <= not(inputs(203));
    layer0_outputs(5181) <= '0';
    layer0_outputs(5182) <= (inputs(123)) and not (inputs(22));
    layer0_outputs(5183) <= (inputs(176)) or (inputs(228));
    layer0_outputs(5184) <= not((inputs(38)) or (inputs(202)));
    layer0_outputs(5185) <= not((inputs(174)) or (inputs(144)));
    layer0_outputs(5186) <= (inputs(177)) and not (inputs(226));
    layer0_outputs(5187) <= not(inputs(148));
    layer0_outputs(5188) <= not(inputs(197)) or (inputs(13));
    layer0_outputs(5189) <= not(inputs(142)) or (inputs(208));
    layer0_outputs(5190) <= not(inputs(211)) or (inputs(133));
    layer0_outputs(5191) <= not((inputs(99)) or (inputs(55)));
    layer0_outputs(5192) <= not(inputs(99)) or (inputs(175));
    layer0_outputs(5193) <= not(inputs(149)) or (inputs(231));
    layer0_outputs(5194) <= (inputs(100)) and not (inputs(41));
    layer0_outputs(5195) <= not(inputs(150));
    layer0_outputs(5196) <= not(inputs(45));
    layer0_outputs(5197) <= '0';
    layer0_outputs(5198) <= inputs(144);
    layer0_outputs(5199) <= not((inputs(42)) or (inputs(70)));
    layer0_outputs(5200) <= not((inputs(190)) or (inputs(4)));
    layer0_outputs(5201) <= '0';
    layer0_outputs(5202) <= not(inputs(49));
    layer0_outputs(5203) <= not(inputs(136)) or (inputs(185));
    layer0_outputs(5204) <= not((inputs(227)) or (inputs(0)));
    layer0_outputs(5205) <= inputs(131);
    layer0_outputs(5206) <= (inputs(106)) or (inputs(94));
    layer0_outputs(5207) <= not(inputs(84)) or (inputs(63));
    layer0_outputs(5208) <= '1';
    layer0_outputs(5209) <= '0';
    layer0_outputs(5210) <= inputs(121);
    layer0_outputs(5211) <= not((inputs(206)) xor (inputs(21)));
    layer0_outputs(5212) <= (inputs(2)) xor (inputs(46));
    layer0_outputs(5213) <= inputs(175);
    layer0_outputs(5214) <= not((inputs(81)) or (inputs(247)));
    layer0_outputs(5215) <= (inputs(61)) or (inputs(120));
    layer0_outputs(5216) <= (inputs(38)) and not (inputs(30));
    layer0_outputs(5217) <= not((inputs(227)) xor (inputs(152)));
    layer0_outputs(5218) <= (inputs(129)) and not (inputs(161));
    layer0_outputs(5219) <= not(inputs(205)) or (inputs(92));
    layer0_outputs(5220) <= (inputs(31)) and (inputs(67));
    layer0_outputs(5221) <= inputs(175);
    layer0_outputs(5222) <= (inputs(139)) and not (inputs(0));
    layer0_outputs(5223) <= not(inputs(179));
    layer0_outputs(5224) <= (inputs(19)) and (inputs(14));
    layer0_outputs(5225) <= not((inputs(68)) xor (inputs(225)));
    layer0_outputs(5226) <= not((inputs(113)) and (inputs(179)));
    layer0_outputs(5227) <= not(inputs(231));
    layer0_outputs(5228) <= '0';
    layer0_outputs(5229) <= (inputs(110)) xor (inputs(14));
    layer0_outputs(5230) <= inputs(230);
    layer0_outputs(5231) <= inputs(180);
    layer0_outputs(5232) <= (inputs(254)) and not (inputs(83));
    layer0_outputs(5233) <= (inputs(252)) or (inputs(127));
    layer0_outputs(5234) <= not((inputs(198)) and (inputs(126)));
    layer0_outputs(5235) <= (inputs(65)) xor (inputs(54));
    layer0_outputs(5236) <= inputs(208);
    layer0_outputs(5237) <= not(inputs(190));
    layer0_outputs(5238) <= not((inputs(142)) and (inputs(76)));
    layer0_outputs(5239) <= (inputs(88)) and not (inputs(224));
    layer0_outputs(5240) <= not(inputs(151));
    layer0_outputs(5241) <= (inputs(17)) or (inputs(113));
    layer0_outputs(5242) <= inputs(1);
    layer0_outputs(5243) <= not((inputs(136)) xor (inputs(240)));
    layer0_outputs(5244) <= not((inputs(248)) or (inputs(114)));
    layer0_outputs(5245) <= '0';
    layer0_outputs(5246) <= not(inputs(212));
    layer0_outputs(5247) <= not(inputs(9)) or (inputs(163));
    layer0_outputs(5248) <= not(inputs(217)) or (inputs(65));
    layer0_outputs(5249) <= (inputs(251)) and not (inputs(10));
    layer0_outputs(5250) <= (inputs(225)) or (inputs(196));
    layer0_outputs(5251) <= (inputs(87)) or (inputs(103));
    layer0_outputs(5252) <= (inputs(242)) and not (inputs(64));
    layer0_outputs(5253) <= (inputs(58)) and not (inputs(2));
    layer0_outputs(5254) <= not(inputs(106));
    layer0_outputs(5255) <= inputs(189);
    layer0_outputs(5256) <= not((inputs(131)) or (inputs(78)));
    layer0_outputs(5257) <= (inputs(172)) and not (inputs(65));
    layer0_outputs(5258) <= '1';
    layer0_outputs(5259) <= not(inputs(55));
    layer0_outputs(5260) <= (inputs(233)) and (inputs(215));
    layer0_outputs(5261) <= '1';
    layer0_outputs(5262) <= not(inputs(221)) or (inputs(57));
    layer0_outputs(5263) <= not(inputs(36));
    layer0_outputs(5264) <= not((inputs(9)) or (inputs(167)));
    layer0_outputs(5265) <= (inputs(145)) or (inputs(157));
    layer0_outputs(5266) <= not((inputs(56)) or (inputs(181)));
    layer0_outputs(5267) <= (inputs(150)) xor (inputs(68));
    layer0_outputs(5268) <= not(inputs(210)) or (inputs(14));
    layer0_outputs(5269) <= inputs(60);
    layer0_outputs(5270) <= (inputs(246)) and (inputs(170));
    layer0_outputs(5271) <= '1';
    layer0_outputs(5272) <= not(inputs(227)) or (inputs(34));
    layer0_outputs(5273) <= not((inputs(153)) xor (inputs(174)));
    layer0_outputs(5274) <= inputs(134);
    layer0_outputs(5275) <= not((inputs(49)) xor (inputs(202)));
    layer0_outputs(5276) <= not(inputs(24)) or (inputs(130));
    layer0_outputs(5277) <= (inputs(47)) and (inputs(39));
    layer0_outputs(5278) <= not(inputs(104)) or (inputs(205));
    layer0_outputs(5279) <= not((inputs(15)) xor (inputs(92)));
    layer0_outputs(5280) <= inputs(19);
    layer0_outputs(5281) <= not(inputs(32)) or (inputs(249));
    layer0_outputs(5282) <= '1';
    layer0_outputs(5283) <= (inputs(184)) and (inputs(184));
    layer0_outputs(5284) <= '0';
    layer0_outputs(5285) <= '1';
    layer0_outputs(5286) <= '1';
    layer0_outputs(5287) <= (inputs(42)) and not (inputs(211));
    layer0_outputs(5288) <= (inputs(228)) and not (inputs(4));
    layer0_outputs(5289) <= (inputs(25)) and not (inputs(238));
    layer0_outputs(5290) <= not(inputs(96));
    layer0_outputs(5291) <= (inputs(142)) or (inputs(84));
    layer0_outputs(5292) <= not(inputs(46)) or (inputs(240));
    layer0_outputs(5293) <= (inputs(226)) and not (inputs(39));
    layer0_outputs(5294) <= not(inputs(37));
    layer0_outputs(5295) <= not((inputs(100)) or (inputs(144)));
    layer0_outputs(5296) <= (inputs(183)) and (inputs(223));
    layer0_outputs(5297) <= not(inputs(112));
    layer0_outputs(5298) <= not(inputs(41));
    layer0_outputs(5299) <= '0';
    layer0_outputs(5300) <= not(inputs(122)) or (inputs(166));
    layer0_outputs(5301) <= '1';
    layer0_outputs(5302) <= not(inputs(133)) or (inputs(196));
    layer0_outputs(5303) <= not((inputs(202)) xor (inputs(205)));
    layer0_outputs(5304) <= (inputs(166)) and not (inputs(218));
    layer0_outputs(5305) <= inputs(210);
    layer0_outputs(5306) <= not(inputs(202)) or (inputs(36));
    layer0_outputs(5307) <= not(inputs(41)) or (inputs(106));
    layer0_outputs(5308) <= not(inputs(59)) or (inputs(252));
    layer0_outputs(5309) <= (inputs(139)) and not (inputs(178));
    layer0_outputs(5310) <= inputs(99);
    layer0_outputs(5311) <= not((inputs(156)) or (inputs(99)));
    layer0_outputs(5312) <= (inputs(186)) or (inputs(143));
    layer0_outputs(5313) <= not((inputs(109)) or (inputs(154)));
    layer0_outputs(5314) <= not(inputs(153));
    layer0_outputs(5315) <= '1';
    layer0_outputs(5316) <= '1';
    layer0_outputs(5317) <= (inputs(75)) and (inputs(26));
    layer0_outputs(5318) <= not(inputs(184));
    layer0_outputs(5319) <= not(inputs(52)) or (inputs(114));
    layer0_outputs(5320) <= (inputs(65)) or (inputs(211));
    layer0_outputs(5321) <= inputs(14);
    layer0_outputs(5322) <= not((inputs(160)) or (inputs(190)));
    layer0_outputs(5323) <= '1';
    layer0_outputs(5324) <= not(inputs(7));
    layer0_outputs(5325) <= (inputs(141)) or (inputs(33));
    layer0_outputs(5326) <= not(inputs(6));
    layer0_outputs(5327) <= not(inputs(100)) or (inputs(17));
    layer0_outputs(5328) <= (inputs(3)) and (inputs(50));
    layer0_outputs(5329) <= (inputs(229)) xor (inputs(6));
    layer0_outputs(5330) <= inputs(142);
    layer0_outputs(5331) <= '1';
    layer0_outputs(5332) <= not(inputs(26)) or (inputs(199));
    layer0_outputs(5333) <= not(inputs(41));
    layer0_outputs(5334) <= not(inputs(184));
    layer0_outputs(5335) <= (inputs(185)) and (inputs(206));
    layer0_outputs(5336) <= not(inputs(249));
    layer0_outputs(5337) <= (inputs(109)) or (inputs(123));
    layer0_outputs(5338) <= (inputs(205)) or (inputs(18));
    layer0_outputs(5339) <= not((inputs(37)) xor (inputs(15)));
    layer0_outputs(5340) <= not((inputs(193)) xor (inputs(248)));
    layer0_outputs(5341) <= inputs(235);
    layer0_outputs(5342) <= not((inputs(169)) xor (inputs(186)));
    layer0_outputs(5343) <= not(inputs(251)) or (inputs(51));
    layer0_outputs(5344) <= inputs(198);
    layer0_outputs(5345) <= inputs(69);
    layer0_outputs(5346) <= inputs(214);
    layer0_outputs(5347) <= not((inputs(228)) xor (inputs(250)));
    layer0_outputs(5348) <= (inputs(202)) and (inputs(183));
    layer0_outputs(5349) <= not(inputs(110));
    layer0_outputs(5350) <= (inputs(44)) and not (inputs(236));
    layer0_outputs(5351) <= not(inputs(171));
    layer0_outputs(5352) <= not(inputs(107));
    layer0_outputs(5353) <= not(inputs(170)) or (inputs(106));
    layer0_outputs(5354) <= (inputs(180)) and not (inputs(242));
    layer0_outputs(5355) <= not(inputs(1)) or (inputs(78));
    layer0_outputs(5356) <= (inputs(181)) and not (inputs(108));
    layer0_outputs(5357) <= inputs(255);
    layer0_outputs(5358) <= not(inputs(106));
    layer0_outputs(5359) <= (inputs(75)) and not (inputs(194));
    layer0_outputs(5360) <= (inputs(98)) or (inputs(16));
    layer0_outputs(5361) <= not((inputs(227)) or (inputs(36)));
    layer0_outputs(5362) <= (inputs(83)) and (inputs(35));
    layer0_outputs(5363) <= (inputs(45)) or (inputs(25));
    layer0_outputs(5364) <= inputs(245);
    layer0_outputs(5365) <= inputs(191);
    layer0_outputs(5366) <= '0';
    layer0_outputs(5367) <= not((inputs(248)) and (inputs(79)));
    layer0_outputs(5368) <= not((inputs(0)) and (inputs(235)));
    layer0_outputs(5369) <= (inputs(199)) or (inputs(224));
    layer0_outputs(5370) <= (inputs(189)) or (inputs(205));
    layer0_outputs(5371) <= (inputs(33)) and not (inputs(254));
    layer0_outputs(5372) <= inputs(78);
    layer0_outputs(5373) <= not(inputs(101));
    layer0_outputs(5374) <= not(inputs(103));
    layer0_outputs(5375) <= inputs(188);
    layer0_outputs(5376) <= '1';
    layer0_outputs(5377) <= '1';
    layer0_outputs(5378) <= '0';
    layer0_outputs(5379) <= inputs(255);
    layer0_outputs(5380) <= inputs(87);
    layer0_outputs(5381) <= (inputs(2)) or (inputs(2));
    layer0_outputs(5382) <= not(inputs(21));
    layer0_outputs(5383) <= not(inputs(115));
    layer0_outputs(5384) <= (inputs(217)) or (inputs(32));
    layer0_outputs(5385) <= (inputs(50)) and (inputs(67));
    layer0_outputs(5386) <= not(inputs(69)) or (inputs(42));
    layer0_outputs(5387) <= (inputs(243)) and not (inputs(74));
    layer0_outputs(5388) <= (inputs(85)) and not (inputs(36));
    layer0_outputs(5389) <= not(inputs(198)) or (inputs(167));
    layer0_outputs(5390) <= '1';
    layer0_outputs(5391) <= (inputs(113)) or (inputs(210));
    layer0_outputs(5392) <= inputs(192);
    layer0_outputs(5393) <= not(inputs(225));
    layer0_outputs(5394) <= '1';
    layer0_outputs(5395) <= not((inputs(173)) and (inputs(215)));
    layer0_outputs(5396) <= '0';
    layer0_outputs(5397) <= inputs(226);
    layer0_outputs(5398) <= not((inputs(148)) or (inputs(253)));
    layer0_outputs(5399) <= not(inputs(155));
    layer0_outputs(5400) <= (inputs(88)) and not (inputs(83));
    layer0_outputs(5401) <= inputs(162);
    layer0_outputs(5402) <= inputs(137);
    layer0_outputs(5403) <= not(inputs(44));
    layer0_outputs(5404) <= not(inputs(159));
    layer0_outputs(5405) <= not(inputs(208)) or (inputs(208));
    layer0_outputs(5406) <= not(inputs(88)) or (inputs(217));
    layer0_outputs(5407) <= (inputs(30)) and not (inputs(234));
    layer0_outputs(5408) <= not((inputs(110)) or (inputs(219)));
    layer0_outputs(5409) <= not(inputs(89));
    layer0_outputs(5410) <= '0';
    layer0_outputs(5411) <= not(inputs(35));
    layer0_outputs(5412) <= not(inputs(248));
    layer0_outputs(5413) <= not((inputs(233)) or (inputs(96)));
    layer0_outputs(5414) <= '0';
    layer0_outputs(5415) <= not(inputs(130));
    layer0_outputs(5416) <= '1';
    layer0_outputs(5417) <= inputs(166);
    layer0_outputs(5418) <= '0';
    layer0_outputs(5419) <= not(inputs(205)) or (inputs(184));
    layer0_outputs(5420) <= (inputs(35)) or (inputs(109));
    layer0_outputs(5421) <= not(inputs(180));
    layer0_outputs(5422) <= '1';
    layer0_outputs(5423) <= (inputs(214)) and (inputs(41));
    layer0_outputs(5424) <= not(inputs(213));
    layer0_outputs(5425) <= not((inputs(10)) or (inputs(23)));
    layer0_outputs(5426) <= inputs(204);
    layer0_outputs(5427) <= inputs(237);
    layer0_outputs(5428) <= not((inputs(140)) or (inputs(102)));
    layer0_outputs(5429) <= (inputs(235)) xor (inputs(226));
    layer0_outputs(5430) <= not((inputs(133)) xor (inputs(120)));
    layer0_outputs(5431) <= (inputs(243)) or (inputs(210));
    layer0_outputs(5432) <= '1';
    layer0_outputs(5433) <= not(inputs(137)) or (inputs(93));
    layer0_outputs(5434) <= (inputs(171)) xor (inputs(195));
    layer0_outputs(5435) <= not(inputs(68));
    layer0_outputs(5436) <= not((inputs(30)) and (inputs(89)));
    layer0_outputs(5437) <= '0';
    layer0_outputs(5438) <= inputs(124);
    layer0_outputs(5439) <= not(inputs(219));
    layer0_outputs(5440) <= (inputs(61)) and not (inputs(153));
    layer0_outputs(5441) <= not(inputs(34)) or (inputs(249));
    layer0_outputs(5442) <= not(inputs(126)) or (inputs(58));
    layer0_outputs(5443) <= not(inputs(57));
    layer0_outputs(5444) <= '0';
    layer0_outputs(5445) <= not((inputs(88)) xor (inputs(151)));
    layer0_outputs(5446) <= not(inputs(147));
    layer0_outputs(5447) <= '1';
    layer0_outputs(5448) <= not(inputs(119));
    layer0_outputs(5449) <= '1';
    layer0_outputs(5450) <= not((inputs(55)) xor (inputs(56)));
    layer0_outputs(5451) <= not((inputs(152)) or (inputs(132)));
    layer0_outputs(5452) <= not((inputs(124)) or (inputs(173)));
    layer0_outputs(5453) <= (inputs(99)) xor (inputs(87));
    layer0_outputs(5454) <= not(inputs(107)) or (inputs(160));
    layer0_outputs(5455) <= inputs(90);
    layer0_outputs(5456) <= not(inputs(41));
    layer0_outputs(5457) <= not((inputs(184)) or (inputs(135)));
    layer0_outputs(5458) <= not(inputs(85)) or (inputs(222));
    layer0_outputs(5459) <= (inputs(127)) or (inputs(110));
    layer0_outputs(5460) <= (inputs(7)) or (inputs(175));
    layer0_outputs(5461) <= (inputs(61)) or (inputs(15));
    layer0_outputs(5462) <= not((inputs(23)) xor (inputs(211)));
    layer0_outputs(5463) <= '0';
    layer0_outputs(5464) <= not((inputs(175)) or (inputs(211)));
    layer0_outputs(5465) <= inputs(36);
    layer0_outputs(5466) <= '1';
    layer0_outputs(5467) <= (inputs(183)) or (inputs(175));
    layer0_outputs(5468) <= not(inputs(211));
    layer0_outputs(5469) <= inputs(74);
    layer0_outputs(5470) <= not(inputs(146));
    layer0_outputs(5471) <= not(inputs(40)) or (inputs(102));
    layer0_outputs(5472) <= not(inputs(217));
    layer0_outputs(5473) <= not((inputs(242)) or (inputs(190)));
    layer0_outputs(5474) <= not(inputs(214));
    layer0_outputs(5475) <= inputs(130);
    layer0_outputs(5476) <= inputs(196);
    layer0_outputs(5477) <= not((inputs(106)) or (inputs(5)));
    layer0_outputs(5478) <= (inputs(251)) xor (inputs(207));
    layer0_outputs(5479) <= not((inputs(111)) or (inputs(40)));
    layer0_outputs(5480) <= (inputs(184)) xor (inputs(137));
    layer0_outputs(5481) <= (inputs(231)) and not (inputs(112));
    layer0_outputs(5482) <= '1';
    layer0_outputs(5483) <= '1';
    layer0_outputs(5484) <= (inputs(162)) and not (inputs(109));
    layer0_outputs(5485) <= not(inputs(201)) or (inputs(130));
    layer0_outputs(5486) <= '1';
    layer0_outputs(5487) <= not((inputs(50)) or (inputs(18)));
    layer0_outputs(5488) <= inputs(231);
    layer0_outputs(5489) <= not(inputs(106));
    layer0_outputs(5490) <= (inputs(199)) and (inputs(202));
    layer0_outputs(5491) <= not(inputs(27));
    layer0_outputs(5492) <= inputs(74);
    layer0_outputs(5493) <= not((inputs(97)) or (inputs(112)));
    layer0_outputs(5494) <= not(inputs(138)) or (inputs(197));
    layer0_outputs(5495) <= not(inputs(150));
    layer0_outputs(5496) <= not(inputs(176));
    layer0_outputs(5497) <= inputs(110);
    layer0_outputs(5498) <= not(inputs(136)) or (inputs(179));
    layer0_outputs(5499) <= inputs(78);
    layer0_outputs(5500) <= not((inputs(97)) xor (inputs(255)));
    layer0_outputs(5501) <= not(inputs(198));
    layer0_outputs(5502) <= inputs(23);
    layer0_outputs(5503) <= (inputs(234)) or (inputs(137));
    layer0_outputs(5504) <= not(inputs(151)) or (inputs(211));
    layer0_outputs(5505) <= '0';
    layer0_outputs(5506) <= inputs(39);
    layer0_outputs(5507) <= not(inputs(238)) or (inputs(29));
    layer0_outputs(5508) <= not(inputs(77));
    layer0_outputs(5509) <= not((inputs(151)) or (inputs(52)));
    layer0_outputs(5510) <= (inputs(20)) and not (inputs(211));
    layer0_outputs(5511) <= not(inputs(105));
    layer0_outputs(5512) <= inputs(164);
    layer0_outputs(5513) <= '0';
    layer0_outputs(5514) <= (inputs(48)) xor (inputs(136));
    layer0_outputs(5515) <= (inputs(4)) and not (inputs(164));
    layer0_outputs(5516) <= (inputs(146)) and not (inputs(79));
    layer0_outputs(5517) <= '0';
    layer0_outputs(5518) <= (inputs(20)) and not (inputs(212));
    layer0_outputs(5519) <= not((inputs(229)) or (inputs(36)));
    layer0_outputs(5520) <= not((inputs(110)) or (inputs(86)));
    layer0_outputs(5521) <= inputs(108);
    layer0_outputs(5522) <= not((inputs(158)) or (inputs(142)));
    layer0_outputs(5523) <= not((inputs(79)) or (inputs(158)));
    layer0_outputs(5524) <= not(inputs(133)) or (inputs(196));
    layer0_outputs(5525) <= not(inputs(11)) or (inputs(90));
    layer0_outputs(5526) <= not((inputs(40)) or (inputs(135)));
    layer0_outputs(5527) <= (inputs(85)) and not (inputs(252));
    layer0_outputs(5528) <= '1';
    layer0_outputs(5529) <= not((inputs(5)) and (inputs(154)));
    layer0_outputs(5530) <= '0';
    layer0_outputs(5531) <= (inputs(107)) and not (inputs(128));
    layer0_outputs(5532) <= not(inputs(166)) or (inputs(4));
    layer0_outputs(5533) <= not((inputs(41)) xor (inputs(57)));
    layer0_outputs(5534) <= not(inputs(94));
    layer0_outputs(5535) <= inputs(63);
    layer0_outputs(5536) <= (inputs(15)) or (inputs(22));
    layer0_outputs(5537) <= (inputs(19)) and not (inputs(7));
    layer0_outputs(5538) <= (inputs(74)) and not (inputs(133));
    layer0_outputs(5539) <= (inputs(91)) and not (inputs(84));
    layer0_outputs(5540) <= not(inputs(193));
    layer0_outputs(5541) <= (inputs(168)) and not (inputs(86));
    layer0_outputs(5542) <= inputs(82);
    layer0_outputs(5543) <= not(inputs(79)) or (inputs(158));
    layer0_outputs(5544) <= (inputs(131)) xor (inputs(221));
    layer0_outputs(5545) <= '1';
    layer0_outputs(5546) <= not(inputs(143));
    layer0_outputs(5547) <= inputs(103);
    layer0_outputs(5548) <= (inputs(168)) and (inputs(59));
    layer0_outputs(5549) <= (inputs(115)) or (inputs(6));
    layer0_outputs(5550) <= (inputs(102)) and not (inputs(148));
    layer0_outputs(5551) <= not(inputs(215));
    layer0_outputs(5552) <= not((inputs(103)) and (inputs(112)));
    layer0_outputs(5553) <= (inputs(124)) and not (inputs(239));
    layer0_outputs(5554) <= not(inputs(254));
    layer0_outputs(5555) <= (inputs(185)) or (inputs(178));
    layer0_outputs(5556) <= not(inputs(133));
    layer0_outputs(5557) <= inputs(146);
    layer0_outputs(5558) <= (inputs(192)) or (inputs(178));
    layer0_outputs(5559) <= (inputs(131)) and not (inputs(67));
    layer0_outputs(5560) <= not(inputs(255));
    layer0_outputs(5561) <= not((inputs(82)) and (inputs(130)));
    layer0_outputs(5562) <= not((inputs(251)) xor (inputs(179)));
    layer0_outputs(5563) <= (inputs(117)) or (inputs(221));
    layer0_outputs(5564) <= (inputs(88)) xor (inputs(153));
    layer0_outputs(5565) <= '0';
    layer0_outputs(5566) <= inputs(85);
    layer0_outputs(5567) <= not(inputs(131)) or (inputs(42));
    layer0_outputs(5568) <= (inputs(241)) or (inputs(122));
    layer0_outputs(5569) <= (inputs(124)) or (inputs(206));
    layer0_outputs(5570) <= not((inputs(150)) xor (inputs(104)));
    layer0_outputs(5571) <= not(inputs(51)) or (inputs(48));
    layer0_outputs(5572) <= inputs(189);
    layer0_outputs(5573) <= not(inputs(14)) or (inputs(46));
    layer0_outputs(5574) <= not((inputs(165)) and (inputs(187)));
    layer0_outputs(5575) <= not((inputs(18)) or (inputs(192)));
    layer0_outputs(5576) <= not(inputs(17)) or (inputs(209));
    layer0_outputs(5577) <= inputs(52);
    layer0_outputs(5578) <= not((inputs(95)) xor (inputs(174)));
    layer0_outputs(5579) <= (inputs(30)) or (inputs(70));
    layer0_outputs(5580) <= (inputs(139)) and not (inputs(125));
    layer0_outputs(5581) <= (inputs(25)) and not (inputs(16));
    layer0_outputs(5582) <= inputs(41);
    layer0_outputs(5583) <= not(inputs(195)) or (inputs(31));
    layer0_outputs(5584) <= not(inputs(145)) or (inputs(214));
    layer0_outputs(5585) <= inputs(183);
    layer0_outputs(5586) <= (inputs(129)) xor (inputs(171));
    layer0_outputs(5587) <= not((inputs(245)) xor (inputs(52)));
    layer0_outputs(5588) <= (inputs(247)) and not (inputs(225));
    layer0_outputs(5589) <= (inputs(158)) and not (inputs(156));
    layer0_outputs(5590) <= not((inputs(56)) and (inputs(211)));
    layer0_outputs(5591) <= (inputs(50)) and not (inputs(160));
    layer0_outputs(5592) <= not(inputs(25)) or (inputs(153));
    layer0_outputs(5593) <= not(inputs(3));
    layer0_outputs(5594) <= not(inputs(162));
    layer0_outputs(5595) <= (inputs(42)) and not (inputs(209));
    layer0_outputs(5596) <= not((inputs(209)) and (inputs(197)));
    layer0_outputs(5597) <= (inputs(77)) xor (inputs(35));
    layer0_outputs(5598) <= not(inputs(123)) or (inputs(153));
    layer0_outputs(5599) <= (inputs(86)) or (inputs(158));
    layer0_outputs(5600) <= not((inputs(65)) or (inputs(147)));
    layer0_outputs(5601) <= not((inputs(164)) and (inputs(28)));
    layer0_outputs(5602) <= inputs(222);
    layer0_outputs(5603) <= inputs(127);
    layer0_outputs(5604) <= inputs(214);
    layer0_outputs(5605) <= not(inputs(95));
    layer0_outputs(5606) <= not((inputs(10)) and (inputs(251)));
    layer0_outputs(5607) <= inputs(142);
    layer0_outputs(5608) <= not(inputs(32));
    layer0_outputs(5609) <= not(inputs(162)) or (inputs(34));
    layer0_outputs(5610) <= not(inputs(122));
    layer0_outputs(5611) <= (inputs(196)) and not (inputs(31));
    layer0_outputs(5612) <= (inputs(187)) and (inputs(187));
    layer0_outputs(5613) <= not((inputs(86)) or (inputs(149)));
    layer0_outputs(5614) <= inputs(202);
    layer0_outputs(5615) <= (inputs(239)) or (inputs(235));
    layer0_outputs(5616) <= inputs(11);
    layer0_outputs(5617) <= not((inputs(198)) and (inputs(200)));
    layer0_outputs(5618) <= not((inputs(243)) and (inputs(44)));
    layer0_outputs(5619) <= '0';
    layer0_outputs(5620) <= (inputs(69)) and (inputs(6));
    layer0_outputs(5621) <= not((inputs(21)) xor (inputs(90)));
    layer0_outputs(5622) <= (inputs(54)) or (inputs(50));
    layer0_outputs(5623) <= '0';
    layer0_outputs(5624) <= not(inputs(120));
    layer0_outputs(5625) <= not((inputs(130)) and (inputs(119)));
    layer0_outputs(5626) <= not(inputs(209)) or (inputs(208));
    layer0_outputs(5627) <= '0';
    layer0_outputs(5628) <= (inputs(214)) or (inputs(160));
    layer0_outputs(5629) <= not(inputs(70)) or (inputs(160));
    layer0_outputs(5630) <= (inputs(200)) or (inputs(111));
    layer0_outputs(5631) <= (inputs(184)) and not (inputs(29));
    layer0_outputs(5632) <= not((inputs(13)) or (inputs(241)));
    layer0_outputs(5633) <= not(inputs(245));
    layer0_outputs(5634) <= not((inputs(136)) and (inputs(153)));
    layer0_outputs(5635) <= (inputs(160)) and not (inputs(146));
    layer0_outputs(5636) <= not(inputs(133));
    layer0_outputs(5637) <= (inputs(245)) and not (inputs(236));
    layer0_outputs(5638) <= not(inputs(107)) or (inputs(248));
    layer0_outputs(5639) <= '1';
    layer0_outputs(5640) <= not((inputs(207)) and (inputs(225)));
    layer0_outputs(5641) <= (inputs(93)) and not (inputs(185));
    layer0_outputs(5642) <= (inputs(206)) or (inputs(160));
    layer0_outputs(5643) <= '0';
    layer0_outputs(5644) <= inputs(125);
    layer0_outputs(5645) <= inputs(117);
    layer0_outputs(5646) <= (inputs(234)) or (inputs(200));
    layer0_outputs(5647) <= not(inputs(96)) or (inputs(114));
    layer0_outputs(5648) <= (inputs(83)) and not (inputs(191));
    layer0_outputs(5649) <= '1';
    layer0_outputs(5650) <= not(inputs(92)) or (inputs(153));
    layer0_outputs(5651) <= inputs(48);
    layer0_outputs(5652) <= not(inputs(191));
    layer0_outputs(5653) <= not((inputs(222)) or (inputs(35)));
    layer0_outputs(5654) <= (inputs(71)) and not (inputs(158));
    layer0_outputs(5655) <= not(inputs(206)) or (inputs(193));
    layer0_outputs(5656) <= '0';
    layer0_outputs(5657) <= not((inputs(98)) and (inputs(96)));
    layer0_outputs(5658) <= (inputs(178)) and not (inputs(208));
    layer0_outputs(5659) <= not(inputs(205));
    layer0_outputs(5660) <= not(inputs(98)) or (inputs(70));
    layer0_outputs(5661) <= not(inputs(128));
    layer0_outputs(5662) <= (inputs(160)) and not (inputs(254));
    layer0_outputs(5663) <= (inputs(25)) or (inputs(29));
    layer0_outputs(5664) <= not(inputs(68));
    layer0_outputs(5665) <= (inputs(42)) or (inputs(94));
    layer0_outputs(5666) <= '0';
    layer0_outputs(5667) <= not((inputs(126)) or (inputs(182)));
    layer0_outputs(5668) <= (inputs(195)) and not (inputs(0));
    layer0_outputs(5669) <= not(inputs(37));
    layer0_outputs(5670) <= (inputs(35)) and not (inputs(239));
    layer0_outputs(5671) <= inputs(15);
    layer0_outputs(5672) <= not((inputs(171)) or (inputs(172)));
    layer0_outputs(5673) <= (inputs(171)) and (inputs(152));
    layer0_outputs(5674) <= not((inputs(21)) and (inputs(26)));
    layer0_outputs(5675) <= '1';
    layer0_outputs(5676) <= not(inputs(142));
    layer0_outputs(5677) <= not(inputs(180));
    layer0_outputs(5678) <= '1';
    layer0_outputs(5679) <= (inputs(170)) or (inputs(127));
    layer0_outputs(5680) <= not(inputs(106));
    layer0_outputs(5681) <= inputs(140);
    layer0_outputs(5682) <= not(inputs(64));
    layer0_outputs(5683) <= inputs(253);
    layer0_outputs(5684) <= (inputs(139)) or (inputs(234));
    layer0_outputs(5685) <= not(inputs(195));
    layer0_outputs(5686) <= not(inputs(179)) or (inputs(229));
    layer0_outputs(5687) <= '0';
    layer0_outputs(5688) <= not(inputs(204)) or (inputs(170));
    layer0_outputs(5689) <= '1';
    layer0_outputs(5690) <= (inputs(212)) or (inputs(222));
    layer0_outputs(5691) <= inputs(136);
    layer0_outputs(5692) <= not((inputs(252)) or (inputs(136)));
    layer0_outputs(5693) <= inputs(143);
    layer0_outputs(5694) <= not((inputs(174)) or (inputs(151)));
    layer0_outputs(5695) <= '0';
    layer0_outputs(5696) <= not((inputs(196)) or (inputs(189)));
    layer0_outputs(5697) <= not(inputs(29));
    layer0_outputs(5698) <= not(inputs(65));
    layer0_outputs(5699) <= '0';
    layer0_outputs(5700) <= (inputs(122)) xor (inputs(253));
    layer0_outputs(5701) <= '0';
    layer0_outputs(5702) <= (inputs(148)) and (inputs(212));
    layer0_outputs(5703) <= not((inputs(23)) or (inputs(39)));
    layer0_outputs(5704) <= not(inputs(231));
    layer0_outputs(5705) <= not(inputs(35)) or (inputs(208));
    layer0_outputs(5706) <= inputs(121);
    layer0_outputs(5707) <= (inputs(105)) and not (inputs(84));
    layer0_outputs(5708) <= (inputs(43)) and not (inputs(183));
    layer0_outputs(5709) <= (inputs(180)) and not (inputs(107));
    layer0_outputs(5710) <= inputs(158);
    layer0_outputs(5711) <= not(inputs(25)) or (inputs(181));
    layer0_outputs(5712) <= not((inputs(66)) and (inputs(24)));
    layer0_outputs(5713) <= not(inputs(124));
    layer0_outputs(5714) <= inputs(203);
    layer0_outputs(5715) <= not((inputs(217)) and (inputs(56)));
    layer0_outputs(5716) <= (inputs(36)) and not (inputs(68));
    layer0_outputs(5717) <= not((inputs(215)) and (inputs(107)));
    layer0_outputs(5718) <= (inputs(198)) or (inputs(246));
    layer0_outputs(5719) <= not(inputs(199)) or (inputs(118));
    layer0_outputs(5720) <= not((inputs(229)) xor (inputs(208)));
    layer0_outputs(5721) <= not(inputs(49));
    layer0_outputs(5722) <= not(inputs(194));
    layer0_outputs(5723) <= not((inputs(51)) xor (inputs(20)));
    layer0_outputs(5724) <= (inputs(199)) and not (inputs(187));
    layer0_outputs(5725) <= not(inputs(119)) or (inputs(13));
    layer0_outputs(5726) <= not(inputs(127)) or (inputs(112));
    layer0_outputs(5727) <= not(inputs(75)) or (inputs(28));
    layer0_outputs(5728) <= (inputs(26)) and not (inputs(239));
    layer0_outputs(5729) <= (inputs(205)) and (inputs(244));
    layer0_outputs(5730) <= (inputs(106)) xor (inputs(111));
    layer0_outputs(5731) <= (inputs(80)) and not (inputs(57));
    layer0_outputs(5732) <= (inputs(167)) and not (inputs(194));
    layer0_outputs(5733) <= not(inputs(131)) or (inputs(202));
    layer0_outputs(5734) <= not(inputs(24));
    layer0_outputs(5735) <= not(inputs(254));
    layer0_outputs(5736) <= inputs(165);
    layer0_outputs(5737) <= inputs(80);
    layer0_outputs(5738) <= (inputs(63)) xor (inputs(176));
    layer0_outputs(5739) <= not(inputs(211)) or (inputs(53));
    layer0_outputs(5740) <= inputs(115);
    layer0_outputs(5741) <= not((inputs(55)) and (inputs(47)));
    layer0_outputs(5742) <= '1';
    layer0_outputs(5743) <= (inputs(86)) and not (inputs(107));
    layer0_outputs(5744) <= not(inputs(96));
    layer0_outputs(5745) <= '0';
    layer0_outputs(5746) <= (inputs(50)) and (inputs(109));
    layer0_outputs(5747) <= inputs(97);
    layer0_outputs(5748) <= inputs(181);
    layer0_outputs(5749) <= not((inputs(226)) xor (inputs(163)));
    layer0_outputs(5750) <= not((inputs(35)) and (inputs(202)));
    layer0_outputs(5751) <= '1';
    layer0_outputs(5752) <= not((inputs(152)) or (inputs(164)));
    layer0_outputs(5753) <= (inputs(105)) or (inputs(181));
    layer0_outputs(5754) <= (inputs(106)) or (inputs(90));
    layer0_outputs(5755) <= (inputs(61)) or (inputs(245));
    layer0_outputs(5756) <= not((inputs(214)) or (inputs(238)));
    layer0_outputs(5757) <= (inputs(68)) and (inputs(3));
    layer0_outputs(5758) <= (inputs(129)) or (inputs(188));
    layer0_outputs(5759) <= not(inputs(144));
    layer0_outputs(5760) <= (inputs(81)) and not (inputs(251));
    layer0_outputs(5761) <= '1';
    layer0_outputs(5762) <= (inputs(126)) and not (inputs(140));
    layer0_outputs(5763) <= not(inputs(118)) or (inputs(255));
    layer0_outputs(5764) <= '0';
    layer0_outputs(5765) <= not(inputs(69)) or (inputs(63));
    layer0_outputs(5766) <= '1';
    layer0_outputs(5767) <= (inputs(94)) or (inputs(204));
    layer0_outputs(5768) <= not((inputs(199)) or (inputs(254)));
    layer0_outputs(5769) <= inputs(29);
    layer0_outputs(5770) <= not((inputs(134)) xor (inputs(57)));
    layer0_outputs(5771) <= not(inputs(243));
    layer0_outputs(5772) <= inputs(115);
    layer0_outputs(5773) <= (inputs(112)) and not (inputs(255));
    layer0_outputs(5774) <= not(inputs(52));
    layer0_outputs(5775) <= (inputs(194)) or (inputs(67));
    layer0_outputs(5776) <= inputs(73);
    layer0_outputs(5777) <= (inputs(95)) and (inputs(74));
    layer0_outputs(5778) <= '1';
    layer0_outputs(5779) <= (inputs(195)) or (inputs(194));
    layer0_outputs(5780) <= (inputs(41)) and not (inputs(251));
    layer0_outputs(5781) <= '0';
    layer0_outputs(5782) <= (inputs(19)) or (inputs(107));
    layer0_outputs(5783) <= (inputs(73)) and (inputs(19));
    layer0_outputs(5784) <= not((inputs(255)) or (inputs(199)));
    layer0_outputs(5785) <= not((inputs(38)) and (inputs(126)));
    layer0_outputs(5786) <= (inputs(4)) and not (inputs(121));
    layer0_outputs(5787) <= not(inputs(250)) or (inputs(152));
    layer0_outputs(5788) <= inputs(105);
    layer0_outputs(5789) <= not(inputs(53)) or (inputs(17));
    layer0_outputs(5790) <= inputs(171);
    layer0_outputs(5791) <= (inputs(226)) and not (inputs(150));
    layer0_outputs(5792) <= (inputs(21)) and not (inputs(77));
    layer0_outputs(5793) <= '0';
    layer0_outputs(5794) <= not(inputs(145)) or (inputs(105));
    layer0_outputs(5795) <= not(inputs(77));
    layer0_outputs(5796) <= (inputs(128)) xor (inputs(4));
    layer0_outputs(5797) <= not(inputs(160));
    layer0_outputs(5798) <= not(inputs(77));
    layer0_outputs(5799) <= '1';
    layer0_outputs(5800) <= (inputs(132)) or (inputs(165));
    layer0_outputs(5801) <= inputs(202);
    layer0_outputs(5802) <= not(inputs(18));
    layer0_outputs(5803) <= not((inputs(80)) xor (inputs(34)));
    layer0_outputs(5804) <= not((inputs(174)) or (inputs(79)));
    layer0_outputs(5805) <= '1';
    layer0_outputs(5806) <= '0';
    layer0_outputs(5807) <= (inputs(176)) xor (inputs(10));
    layer0_outputs(5808) <= not(inputs(102)) or (inputs(108));
    layer0_outputs(5809) <= not(inputs(107));
    layer0_outputs(5810) <= not((inputs(194)) or (inputs(95)));
    layer0_outputs(5811) <= not(inputs(230));
    layer0_outputs(5812) <= inputs(147);
    layer0_outputs(5813) <= not(inputs(214));
    layer0_outputs(5814) <= (inputs(48)) xor (inputs(92));
    layer0_outputs(5815) <= (inputs(65)) or (inputs(21));
    layer0_outputs(5816) <= inputs(23);
    layer0_outputs(5817) <= (inputs(174)) or (inputs(243));
    layer0_outputs(5818) <= not((inputs(161)) xor (inputs(213)));
    layer0_outputs(5819) <= (inputs(160)) or (inputs(144));
    layer0_outputs(5820) <= (inputs(164)) and not (inputs(92));
    layer0_outputs(5821) <= (inputs(142)) or (inputs(233));
    layer0_outputs(5822) <= not(inputs(122)) or (inputs(147));
    layer0_outputs(5823) <= (inputs(210)) or (inputs(214));
    layer0_outputs(5824) <= (inputs(241)) and not (inputs(63));
    layer0_outputs(5825) <= '0';
    layer0_outputs(5826) <= '0';
    layer0_outputs(5827) <= '1';
    layer0_outputs(5828) <= not(inputs(78)) or (inputs(169));
    layer0_outputs(5829) <= not(inputs(13)) or (inputs(61));
    layer0_outputs(5830) <= not((inputs(45)) or (inputs(7)));
    layer0_outputs(5831) <= (inputs(86)) and not (inputs(222));
    layer0_outputs(5832) <= '1';
    layer0_outputs(5833) <= not(inputs(58));
    layer0_outputs(5834) <= not((inputs(196)) xor (inputs(127)));
    layer0_outputs(5835) <= not((inputs(224)) and (inputs(97)));
    layer0_outputs(5836) <= (inputs(95)) and not (inputs(228));
    layer0_outputs(5837) <= (inputs(81)) and not (inputs(12));
    layer0_outputs(5838) <= not(inputs(132)) or (inputs(196));
    layer0_outputs(5839) <= (inputs(136)) and (inputs(167));
    layer0_outputs(5840) <= inputs(78);
    layer0_outputs(5841) <= not(inputs(211)) or (inputs(29));
    layer0_outputs(5842) <= not((inputs(112)) or (inputs(246)));
    layer0_outputs(5843) <= inputs(194);
    layer0_outputs(5844) <= (inputs(180)) or (inputs(221));
    layer0_outputs(5845) <= not((inputs(134)) or (inputs(81)));
    layer0_outputs(5846) <= (inputs(232)) xor (inputs(216));
    layer0_outputs(5847) <= '1';
    layer0_outputs(5848) <= inputs(25);
    layer0_outputs(5849) <= (inputs(237)) and not (inputs(168));
    layer0_outputs(5850) <= inputs(8);
    layer0_outputs(5851) <= (inputs(159)) and not (inputs(101));
    layer0_outputs(5852) <= not((inputs(140)) and (inputs(215)));
    layer0_outputs(5853) <= not(inputs(11));
    layer0_outputs(5854) <= not((inputs(241)) xor (inputs(8)));
    layer0_outputs(5855) <= not(inputs(97));
    layer0_outputs(5856) <= not((inputs(62)) or (inputs(241)));
    layer0_outputs(5857) <= not((inputs(222)) or (inputs(32)));
    layer0_outputs(5858) <= inputs(206);
    layer0_outputs(5859) <= not(inputs(137));
    layer0_outputs(5860) <= not((inputs(41)) and (inputs(15)));
    layer0_outputs(5861) <= (inputs(18)) or (inputs(62));
    layer0_outputs(5862) <= (inputs(193)) or (inputs(192));
    layer0_outputs(5863) <= not(inputs(30));
    layer0_outputs(5864) <= not((inputs(66)) xor (inputs(163)));
    layer0_outputs(5865) <= not((inputs(93)) xor (inputs(19)));
    layer0_outputs(5866) <= not(inputs(122));
    layer0_outputs(5867) <= not(inputs(241));
    layer0_outputs(5868) <= (inputs(235)) or (inputs(26));
    layer0_outputs(5869) <= not((inputs(88)) and (inputs(103)));
    layer0_outputs(5870) <= not(inputs(147)) or (inputs(215));
    layer0_outputs(5871) <= (inputs(234)) and not (inputs(138));
    layer0_outputs(5872) <= inputs(117);
    layer0_outputs(5873) <= (inputs(66)) xor (inputs(20));
    layer0_outputs(5874) <= (inputs(68)) and not (inputs(126));
    layer0_outputs(5875) <= not(inputs(254));
    layer0_outputs(5876) <= inputs(88);
    layer0_outputs(5877) <= not(inputs(100));
    layer0_outputs(5878) <= not(inputs(102));
    layer0_outputs(5879) <= not((inputs(108)) xor (inputs(234)));
    layer0_outputs(5880) <= not(inputs(70)) or (inputs(201));
    layer0_outputs(5881) <= not(inputs(102)) or (inputs(148));
    layer0_outputs(5882) <= (inputs(186)) and (inputs(212));
    layer0_outputs(5883) <= not((inputs(191)) xor (inputs(181)));
    layer0_outputs(5884) <= (inputs(111)) or (inputs(75));
    layer0_outputs(5885) <= (inputs(166)) and not (inputs(119));
    layer0_outputs(5886) <= not(inputs(199));
    layer0_outputs(5887) <= not(inputs(102));
    layer0_outputs(5888) <= not(inputs(182));
    layer0_outputs(5889) <= (inputs(43)) or (inputs(50));
    layer0_outputs(5890) <= not(inputs(115)) or (inputs(15));
    layer0_outputs(5891) <= inputs(218);
    layer0_outputs(5892) <= '0';
    layer0_outputs(5893) <= not(inputs(156)) or (inputs(61));
    layer0_outputs(5894) <= '0';
    layer0_outputs(5895) <= inputs(90);
    layer0_outputs(5896) <= (inputs(64)) and not (inputs(62));
    layer0_outputs(5897) <= (inputs(228)) xor (inputs(251));
    layer0_outputs(5898) <= not(inputs(106));
    layer0_outputs(5899) <= not(inputs(141));
    layer0_outputs(5900) <= (inputs(114)) and not (inputs(10));
    layer0_outputs(5901) <= not(inputs(105)) or (inputs(239));
    layer0_outputs(5902) <= inputs(209);
    layer0_outputs(5903) <= not(inputs(164)) or (inputs(176));
    layer0_outputs(5904) <= '1';
    layer0_outputs(5905) <= inputs(200);
    layer0_outputs(5906) <= not(inputs(245)) or (inputs(65));
    layer0_outputs(5907) <= inputs(63);
    layer0_outputs(5908) <= (inputs(171)) or (inputs(112));
    layer0_outputs(5909) <= not(inputs(128));
    layer0_outputs(5910) <= inputs(81);
    layer0_outputs(5911) <= (inputs(170)) or (inputs(111));
    layer0_outputs(5912) <= not(inputs(233)) or (inputs(217));
    layer0_outputs(5913) <= not((inputs(58)) xor (inputs(29)));
    layer0_outputs(5914) <= not(inputs(166)) or (inputs(62));
    layer0_outputs(5915) <= '0';
    layer0_outputs(5916) <= (inputs(246)) or (inputs(100));
    layer0_outputs(5917) <= not(inputs(140));
    layer0_outputs(5918) <= not((inputs(171)) and (inputs(218)));
    layer0_outputs(5919) <= not((inputs(29)) or (inputs(97)));
    layer0_outputs(5920) <= inputs(226);
    layer0_outputs(5921) <= '0';
    layer0_outputs(5922) <= '0';
    layer0_outputs(5923) <= (inputs(184)) and not (inputs(172));
    layer0_outputs(5924) <= not(inputs(141));
    layer0_outputs(5925) <= inputs(130);
    layer0_outputs(5926) <= inputs(182);
    layer0_outputs(5927) <= inputs(76);
    layer0_outputs(5928) <= '1';
    layer0_outputs(5929) <= (inputs(90)) and not (inputs(193));
    layer0_outputs(5930) <= not(inputs(98));
    layer0_outputs(5931) <= (inputs(235)) or (inputs(151));
    layer0_outputs(5932) <= inputs(95);
    layer0_outputs(5933) <= not(inputs(220));
    layer0_outputs(5934) <= inputs(23);
    layer0_outputs(5935) <= not(inputs(230));
    layer0_outputs(5936) <= not(inputs(57)) or (inputs(23));
    layer0_outputs(5937) <= inputs(59);
    layer0_outputs(5938) <= '0';
    layer0_outputs(5939) <= (inputs(113)) or (inputs(141));
    layer0_outputs(5940) <= (inputs(130)) xor (inputs(220));
    layer0_outputs(5941) <= (inputs(253)) and not (inputs(122));
    layer0_outputs(5942) <= not(inputs(205));
    layer0_outputs(5943) <= not(inputs(127));
    layer0_outputs(5944) <= '1';
    layer0_outputs(5945) <= (inputs(89)) and (inputs(224));
    layer0_outputs(5946) <= inputs(31);
    layer0_outputs(5947) <= (inputs(75)) and not (inputs(176));
    layer0_outputs(5948) <= inputs(41);
    layer0_outputs(5949) <= (inputs(165)) and not (inputs(75));
    layer0_outputs(5950) <= not((inputs(146)) xor (inputs(104)));
    layer0_outputs(5951) <= (inputs(254)) and not (inputs(47));
    layer0_outputs(5952) <= (inputs(89)) and not (inputs(48));
    layer0_outputs(5953) <= '0';
    layer0_outputs(5954) <= '1';
    layer0_outputs(5955) <= not(inputs(249)) or (inputs(208));
    layer0_outputs(5956) <= '1';
    layer0_outputs(5957) <= not((inputs(47)) xor (inputs(250)));
    layer0_outputs(5958) <= not(inputs(195));
    layer0_outputs(5959) <= (inputs(223)) and (inputs(14));
    layer0_outputs(5960) <= (inputs(80)) xor (inputs(68));
    layer0_outputs(5961) <= not((inputs(46)) and (inputs(175)));
    layer0_outputs(5962) <= '0';
    layer0_outputs(5963) <= (inputs(141)) or (inputs(224));
    layer0_outputs(5964) <= not((inputs(147)) or (inputs(189)));
    layer0_outputs(5965) <= (inputs(231)) or (inputs(192));
    layer0_outputs(5966) <= not(inputs(234));
    layer0_outputs(5967) <= (inputs(146)) and not (inputs(46));
    layer0_outputs(5968) <= '1';
    layer0_outputs(5969) <= (inputs(222)) or (inputs(229));
    layer0_outputs(5970) <= (inputs(245)) and not (inputs(189));
    layer0_outputs(5971) <= not(inputs(135)) or (inputs(24));
    layer0_outputs(5972) <= not((inputs(149)) xor (inputs(144)));
    layer0_outputs(5973) <= inputs(243);
    layer0_outputs(5974) <= not((inputs(194)) or (inputs(6)));
    layer0_outputs(5975) <= (inputs(132)) and not (inputs(237));
    layer0_outputs(5976) <= not(inputs(181));
    layer0_outputs(5977) <= (inputs(132)) and not (inputs(14));
    layer0_outputs(5978) <= not((inputs(237)) and (inputs(165)));
    layer0_outputs(5979) <= (inputs(229)) and not (inputs(131));
    layer0_outputs(5980) <= not(inputs(234)) or (inputs(116));
    layer0_outputs(5981) <= not((inputs(51)) or (inputs(168)));
    layer0_outputs(5982) <= not((inputs(8)) or (inputs(230)));
    layer0_outputs(5983) <= not((inputs(31)) or (inputs(153)));
    layer0_outputs(5984) <= (inputs(109)) or (inputs(95));
    layer0_outputs(5985) <= inputs(151);
    layer0_outputs(5986) <= '0';
    layer0_outputs(5987) <= (inputs(182)) and (inputs(157));
    layer0_outputs(5988) <= (inputs(53)) and not (inputs(134));
    layer0_outputs(5989) <= not(inputs(173)) or (inputs(111));
    layer0_outputs(5990) <= (inputs(219)) xor (inputs(179));
    layer0_outputs(5991) <= (inputs(236)) and not (inputs(66));
    layer0_outputs(5992) <= not(inputs(138)) or (inputs(36));
    layer0_outputs(5993) <= inputs(140);
    layer0_outputs(5994) <= not(inputs(141));
    layer0_outputs(5995) <= not(inputs(254));
    layer0_outputs(5996) <= not(inputs(105));
    layer0_outputs(5997) <= inputs(147);
    layer0_outputs(5998) <= not(inputs(230)) or (inputs(0));
    layer0_outputs(5999) <= not(inputs(95));
    layer0_outputs(6000) <= not((inputs(231)) or (inputs(159)));
    layer0_outputs(6001) <= not(inputs(149));
    layer0_outputs(6002) <= inputs(92);
    layer0_outputs(6003) <= not((inputs(51)) and (inputs(224)));
    layer0_outputs(6004) <= (inputs(232)) and not (inputs(247));
    layer0_outputs(6005) <= not((inputs(44)) or (inputs(201)));
    layer0_outputs(6006) <= (inputs(93)) or (inputs(32));
    layer0_outputs(6007) <= (inputs(5)) or (inputs(28));
    layer0_outputs(6008) <= not(inputs(220));
    layer0_outputs(6009) <= not(inputs(225));
    layer0_outputs(6010) <= inputs(13);
    layer0_outputs(6011) <= '1';
    layer0_outputs(6012) <= (inputs(100)) and not (inputs(64));
    layer0_outputs(6013) <= not((inputs(201)) or (inputs(3)));
    layer0_outputs(6014) <= not(inputs(231));
    layer0_outputs(6015) <= inputs(227);
    layer0_outputs(6016) <= (inputs(27)) and not (inputs(163));
    layer0_outputs(6017) <= (inputs(189)) and not (inputs(65));
    layer0_outputs(6018) <= '1';
    layer0_outputs(6019) <= not(inputs(43));
    layer0_outputs(6020) <= not((inputs(179)) or (inputs(116)));
    layer0_outputs(6021) <= '1';
    layer0_outputs(6022) <= not((inputs(94)) and (inputs(81)));
    layer0_outputs(6023) <= not(inputs(229));
    layer0_outputs(6024) <= inputs(131);
    layer0_outputs(6025) <= (inputs(76)) or (inputs(114));
    layer0_outputs(6026) <= not(inputs(253));
    layer0_outputs(6027) <= not(inputs(103));
    layer0_outputs(6028) <= (inputs(148)) and not (inputs(55));
    layer0_outputs(6029) <= not(inputs(100));
    layer0_outputs(6030) <= not(inputs(49)) or (inputs(127));
    layer0_outputs(6031) <= (inputs(23)) or (inputs(96));
    layer0_outputs(6032) <= (inputs(98)) and not (inputs(115));
    layer0_outputs(6033) <= (inputs(76)) and not (inputs(169));
    layer0_outputs(6034) <= inputs(164);
    layer0_outputs(6035) <= inputs(29);
    layer0_outputs(6036) <= not(inputs(117));
    layer0_outputs(6037) <= '1';
    layer0_outputs(6038) <= (inputs(181)) xor (inputs(109));
    layer0_outputs(6039) <= not((inputs(241)) or (inputs(241)));
    layer0_outputs(6040) <= (inputs(168)) and (inputs(190));
    layer0_outputs(6041) <= not((inputs(193)) xor (inputs(195)));
    layer0_outputs(6042) <= '1';
    layer0_outputs(6043) <= (inputs(168)) and not (inputs(94));
    layer0_outputs(6044) <= not(inputs(213)) or (inputs(239));
    layer0_outputs(6045) <= (inputs(144)) and not (inputs(245));
    layer0_outputs(6046) <= not(inputs(24));
    layer0_outputs(6047) <= not(inputs(0));
    layer0_outputs(6048) <= (inputs(202)) or (inputs(67));
    layer0_outputs(6049) <= inputs(225);
    layer0_outputs(6050) <= not(inputs(248));
    layer0_outputs(6051) <= not((inputs(111)) and (inputs(105)));
    layer0_outputs(6052) <= inputs(56);
    layer0_outputs(6053) <= not((inputs(116)) or (inputs(53)));
    layer0_outputs(6054) <= not((inputs(162)) or (inputs(169)));
    layer0_outputs(6055) <= (inputs(157)) xor (inputs(119));
    layer0_outputs(6056) <= not(inputs(99));
    layer0_outputs(6057) <= '1';
    layer0_outputs(6058) <= (inputs(140)) and (inputs(93));
    layer0_outputs(6059) <= not(inputs(199)) or (inputs(152));
    layer0_outputs(6060) <= not(inputs(6));
    layer0_outputs(6061) <= (inputs(104)) xor (inputs(236));
    layer0_outputs(6062) <= (inputs(65)) and not (inputs(107));
    layer0_outputs(6063) <= not(inputs(87));
    layer0_outputs(6064) <= not((inputs(199)) or (inputs(245)));
    layer0_outputs(6065) <= not(inputs(151)) or (inputs(128));
    layer0_outputs(6066) <= not((inputs(148)) xor (inputs(86)));
    layer0_outputs(6067) <= not((inputs(91)) or (inputs(99)));
    layer0_outputs(6068) <= not(inputs(106));
    layer0_outputs(6069) <= (inputs(110)) and not (inputs(56));
    layer0_outputs(6070) <= (inputs(66)) and (inputs(243));
    layer0_outputs(6071) <= inputs(247);
    layer0_outputs(6072) <= (inputs(80)) or (inputs(24));
    layer0_outputs(6073) <= '0';
    layer0_outputs(6074) <= (inputs(86)) and (inputs(22));
    layer0_outputs(6075) <= (inputs(134)) or (inputs(185));
    layer0_outputs(6076) <= (inputs(77)) and not (inputs(88));
    layer0_outputs(6077) <= (inputs(23)) and not (inputs(171));
    layer0_outputs(6078) <= (inputs(210)) or (inputs(186));
    layer0_outputs(6079) <= not(inputs(22));
    layer0_outputs(6080) <= '0';
    layer0_outputs(6081) <= (inputs(173)) and not (inputs(153));
    layer0_outputs(6082) <= (inputs(243)) and not (inputs(35));
    layer0_outputs(6083) <= inputs(49);
    layer0_outputs(6084) <= inputs(120);
    layer0_outputs(6085) <= not(inputs(178)) or (inputs(184));
    layer0_outputs(6086) <= not((inputs(144)) or (inputs(130)));
    layer0_outputs(6087) <= not((inputs(161)) xor (inputs(53)));
    layer0_outputs(6088) <= (inputs(194)) or (inputs(177));
    layer0_outputs(6089) <= not(inputs(155));
    layer0_outputs(6090) <= not((inputs(82)) or (inputs(99)));
    layer0_outputs(6091) <= (inputs(212)) and not (inputs(239));
    layer0_outputs(6092) <= not(inputs(16)) or (inputs(41));
    layer0_outputs(6093) <= not(inputs(38)) or (inputs(205));
    layer0_outputs(6094) <= not((inputs(189)) and (inputs(72)));
    layer0_outputs(6095) <= '0';
    layer0_outputs(6096) <= (inputs(191)) and not (inputs(208));
    layer0_outputs(6097) <= not(inputs(52)) or (inputs(57));
    layer0_outputs(6098) <= not((inputs(177)) or (inputs(16)));
    layer0_outputs(6099) <= (inputs(237)) or (inputs(234));
    layer0_outputs(6100) <= inputs(249);
    layer0_outputs(6101) <= '0';
    layer0_outputs(6102) <= (inputs(114)) and not (inputs(73));
    layer0_outputs(6103) <= not(inputs(195)) or (inputs(63));
    layer0_outputs(6104) <= inputs(223);
    layer0_outputs(6105) <= not((inputs(58)) and (inputs(116)));
    layer0_outputs(6106) <= (inputs(101)) or (inputs(98));
    layer0_outputs(6107) <= not(inputs(142)) or (inputs(165));
    layer0_outputs(6108) <= (inputs(109)) and not (inputs(46));
    layer0_outputs(6109) <= (inputs(217)) and not (inputs(124));
    layer0_outputs(6110) <= inputs(105);
    layer0_outputs(6111) <= (inputs(154)) and not (inputs(9));
    layer0_outputs(6112) <= not(inputs(64));
    layer0_outputs(6113) <= inputs(1);
    layer0_outputs(6114) <= not(inputs(116));
    layer0_outputs(6115) <= (inputs(127)) and not (inputs(215));
    layer0_outputs(6116) <= not(inputs(99));
    layer0_outputs(6117) <= '0';
    layer0_outputs(6118) <= not(inputs(155));
    layer0_outputs(6119) <= inputs(105);
    layer0_outputs(6120) <= (inputs(107)) xor (inputs(94));
    layer0_outputs(6121) <= inputs(33);
    layer0_outputs(6122) <= not((inputs(207)) xor (inputs(241)));
    layer0_outputs(6123) <= not((inputs(68)) xor (inputs(184)));
    layer0_outputs(6124) <= inputs(152);
    layer0_outputs(6125) <= inputs(40);
    layer0_outputs(6126) <= (inputs(135)) and not (inputs(13));
    layer0_outputs(6127) <= (inputs(32)) or (inputs(222));
    layer0_outputs(6128) <= not((inputs(20)) xor (inputs(187)));
    layer0_outputs(6129) <= not(inputs(72)) or (inputs(69));
    layer0_outputs(6130) <= (inputs(1)) xor (inputs(157));
    layer0_outputs(6131) <= not((inputs(87)) or (inputs(13)));
    layer0_outputs(6132) <= (inputs(248)) and not (inputs(80));
    layer0_outputs(6133) <= not(inputs(112)) or (inputs(174));
    layer0_outputs(6134) <= '1';
    layer0_outputs(6135) <= not(inputs(77));
    layer0_outputs(6136) <= inputs(25);
    layer0_outputs(6137) <= not((inputs(170)) or (inputs(54)));
    layer0_outputs(6138) <= (inputs(102)) and (inputs(141));
    layer0_outputs(6139) <= not(inputs(245));
    layer0_outputs(6140) <= not((inputs(222)) xor (inputs(134)));
    layer0_outputs(6141) <= not(inputs(73)) or (inputs(36));
    layer0_outputs(6142) <= not(inputs(153));
    layer0_outputs(6143) <= (inputs(158)) or (inputs(190));
    layer0_outputs(6144) <= not(inputs(180));
    layer0_outputs(6145) <= (inputs(2)) xor (inputs(85));
    layer0_outputs(6146) <= not(inputs(123));
    layer0_outputs(6147) <= not(inputs(246));
    layer0_outputs(6148) <= not(inputs(67));
    layer0_outputs(6149) <= not((inputs(243)) and (inputs(240)));
    layer0_outputs(6150) <= inputs(212);
    layer0_outputs(6151) <= (inputs(17)) and not (inputs(217));
    layer0_outputs(6152) <= not(inputs(195)) or (inputs(124));
    layer0_outputs(6153) <= '0';
    layer0_outputs(6154) <= not((inputs(134)) and (inputs(193)));
    layer0_outputs(6155) <= not(inputs(104)) or (inputs(139));
    layer0_outputs(6156) <= not(inputs(238));
    layer0_outputs(6157) <= not(inputs(112)) or (inputs(29));
    layer0_outputs(6158) <= not(inputs(215)) or (inputs(238));
    layer0_outputs(6159) <= not(inputs(3));
    layer0_outputs(6160) <= '1';
    layer0_outputs(6161) <= inputs(43);
    layer0_outputs(6162) <= (inputs(147)) or (inputs(158));
    layer0_outputs(6163) <= inputs(205);
    layer0_outputs(6164) <= inputs(152);
    layer0_outputs(6165) <= not(inputs(33)) or (inputs(148));
    layer0_outputs(6166) <= not(inputs(224));
    layer0_outputs(6167) <= '1';
    layer0_outputs(6168) <= (inputs(30)) or (inputs(216));
    layer0_outputs(6169) <= (inputs(27)) and (inputs(38));
    layer0_outputs(6170) <= not(inputs(216)) or (inputs(92));
    layer0_outputs(6171) <= not((inputs(229)) and (inputs(201)));
    layer0_outputs(6172) <= not((inputs(201)) xor (inputs(233)));
    layer0_outputs(6173) <= not(inputs(184)) or (inputs(139));
    layer0_outputs(6174) <= not(inputs(208));
    layer0_outputs(6175) <= not((inputs(129)) and (inputs(179)));
    layer0_outputs(6176) <= not(inputs(29));
    layer0_outputs(6177) <= not(inputs(250)) or (inputs(203));
    layer0_outputs(6178) <= not(inputs(163));
    layer0_outputs(6179) <= not(inputs(189));
    layer0_outputs(6180) <= inputs(235);
    layer0_outputs(6181) <= (inputs(166)) or (inputs(83));
    layer0_outputs(6182) <= inputs(209);
    layer0_outputs(6183) <= '1';
    layer0_outputs(6184) <= (inputs(201)) and (inputs(194));
    layer0_outputs(6185) <= (inputs(13)) or (inputs(15));
    layer0_outputs(6186) <= not(inputs(214));
    layer0_outputs(6187) <= (inputs(173)) and not (inputs(70));
    layer0_outputs(6188) <= inputs(227);
    layer0_outputs(6189) <= inputs(114);
    layer0_outputs(6190) <= inputs(146);
    layer0_outputs(6191) <= not(inputs(38)) or (inputs(190));
    layer0_outputs(6192) <= not((inputs(122)) or (inputs(237)));
    layer0_outputs(6193) <= (inputs(208)) and not (inputs(142));
    layer0_outputs(6194) <= '1';
    layer0_outputs(6195) <= not(inputs(223)) or (inputs(141));
    layer0_outputs(6196) <= not(inputs(251)) or (inputs(26));
    layer0_outputs(6197) <= '1';
    layer0_outputs(6198) <= not(inputs(162)) or (inputs(109));
    layer0_outputs(6199) <= not((inputs(253)) or (inputs(134)));
    layer0_outputs(6200) <= not(inputs(10)) or (inputs(180));
    layer0_outputs(6201) <= not((inputs(205)) or (inputs(44)));
    layer0_outputs(6202) <= not(inputs(147));
    layer0_outputs(6203) <= inputs(165);
    layer0_outputs(6204) <= not(inputs(187)) or (inputs(109));
    layer0_outputs(6205) <= not(inputs(66));
    layer0_outputs(6206) <= inputs(89);
    layer0_outputs(6207) <= (inputs(71)) and (inputs(199));
    layer0_outputs(6208) <= not(inputs(25));
    layer0_outputs(6209) <= not((inputs(60)) or (inputs(205)));
    layer0_outputs(6210) <= not(inputs(88));
    layer0_outputs(6211) <= not((inputs(221)) and (inputs(41)));
    layer0_outputs(6212) <= inputs(26);
    layer0_outputs(6213) <= not((inputs(146)) and (inputs(17)));
    layer0_outputs(6214) <= not(inputs(103));
    layer0_outputs(6215) <= (inputs(128)) and not (inputs(214));
    layer0_outputs(6216) <= not(inputs(165)) or (inputs(107));
    layer0_outputs(6217) <= not(inputs(83)) or (inputs(206));
    layer0_outputs(6218) <= not((inputs(32)) and (inputs(109)));
    layer0_outputs(6219) <= not(inputs(212));
    layer0_outputs(6220) <= '0';
    layer0_outputs(6221) <= not(inputs(230));
    layer0_outputs(6222) <= (inputs(237)) and not (inputs(169));
    layer0_outputs(6223) <= (inputs(143)) and not (inputs(59));
    layer0_outputs(6224) <= (inputs(9)) or (inputs(174));
    layer0_outputs(6225) <= inputs(23);
    layer0_outputs(6226) <= not(inputs(68));
    layer0_outputs(6227) <= not(inputs(37));
    layer0_outputs(6228) <= not(inputs(85)) or (inputs(18));
    layer0_outputs(6229) <= inputs(168);
    layer0_outputs(6230) <= not((inputs(203)) or (inputs(220)));
    layer0_outputs(6231) <= not(inputs(133));
    layer0_outputs(6232) <= not((inputs(105)) or (inputs(181)));
    layer0_outputs(6233) <= not(inputs(109));
    layer0_outputs(6234) <= not(inputs(215)) or (inputs(77));
    layer0_outputs(6235) <= not((inputs(148)) or (inputs(142)));
    layer0_outputs(6236) <= inputs(172);
    layer0_outputs(6237) <= inputs(231);
    layer0_outputs(6238) <= not(inputs(230)) or (inputs(13));
    layer0_outputs(6239) <= not(inputs(117)) or (inputs(89));
    layer0_outputs(6240) <= inputs(163);
    layer0_outputs(6241) <= (inputs(36)) and (inputs(142));
    layer0_outputs(6242) <= not(inputs(120));
    layer0_outputs(6243) <= '1';
    layer0_outputs(6244) <= not((inputs(247)) or (inputs(248)));
    layer0_outputs(6245) <= not(inputs(28)) or (inputs(67));
    layer0_outputs(6246) <= inputs(75);
    layer0_outputs(6247) <= (inputs(35)) and not (inputs(128));
    layer0_outputs(6248) <= not(inputs(228)) or (inputs(74));
    layer0_outputs(6249) <= '0';
    layer0_outputs(6250) <= inputs(61);
    layer0_outputs(6251) <= not(inputs(52));
    layer0_outputs(6252) <= not(inputs(146));
    layer0_outputs(6253) <= not(inputs(70)) or (inputs(232));
    layer0_outputs(6254) <= not(inputs(242)) or (inputs(29));
    layer0_outputs(6255) <= (inputs(137)) or (inputs(191));
    layer0_outputs(6256) <= inputs(110);
    layer0_outputs(6257) <= inputs(173);
    layer0_outputs(6258) <= inputs(114);
    layer0_outputs(6259) <= '0';
    layer0_outputs(6260) <= not(inputs(177));
    layer0_outputs(6261) <= not(inputs(118)) or (inputs(112));
    layer0_outputs(6262) <= inputs(129);
    layer0_outputs(6263) <= not(inputs(38));
    layer0_outputs(6264) <= not(inputs(244));
    layer0_outputs(6265) <= '1';
    layer0_outputs(6266) <= (inputs(81)) and not (inputs(253));
    layer0_outputs(6267) <= '0';
    layer0_outputs(6268) <= (inputs(161)) and not (inputs(141));
    layer0_outputs(6269) <= not(inputs(83));
    layer0_outputs(6270) <= '1';
    layer0_outputs(6271) <= (inputs(187)) or (inputs(95));
    layer0_outputs(6272) <= not((inputs(172)) xor (inputs(158)));
    layer0_outputs(6273) <= inputs(75);
    layer0_outputs(6274) <= not(inputs(131));
    layer0_outputs(6275) <= '0';
    layer0_outputs(6276) <= inputs(74);
    layer0_outputs(6277) <= inputs(129);
    layer0_outputs(6278) <= (inputs(191)) xor (inputs(17));
    layer0_outputs(6279) <= not((inputs(193)) or (inputs(113)));
    layer0_outputs(6280) <= (inputs(204)) or (inputs(203));
    layer0_outputs(6281) <= inputs(231);
    layer0_outputs(6282) <= not((inputs(26)) or (inputs(209)));
    layer0_outputs(6283) <= (inputs(9)) and not (inputs(184));
    layer0_outputs(6284) <= '1';
    layer0_outputs(6285) <= not(inputs(30));
    layer0_outputs(6286) <= (inputs(4)) and not (inputs(28));
    layer0_outputs(6287) <= inputs(250);
    layer0_outputs(6288) <= not((inputs(41)) or (inputs(209)));
    layer0_outputs(6289) <= inputs(4);
    layer0_outputs(6290) <= not(inputs(38));
    layer0_outputs(6291) <= not(inputs(4));
    layer0_outputs(6292) <= (inputs(67)) or (inputs(126));
    layer0_outputs(6293) <= '1';
    layer0_outputs(6294) <= inputs(58);
    layer0_outputs(6295) <= (inputs(229)) and not (inputs(60));
    layer0_outputs(6296) <= not(inputs(202));
    layer0_outputs(6297) <= not((inputs(11)) and (inputs(3)));
    layer0_outputs(6298) <= '0';
    layer0_outputs(6299) <= inputs(224);
    layer0_outputs(6300) <= not((inputs(78)) and (inputs(162)));
    layer0_outputs(6301) <= not((inputs(178)) xor (inputs(203)));
    layer0_outputs(6302) <= not(inputs(213));
    layer0_outputs(6303) <= inputs(12);
    layer0_outputs(6304) <= (inputs(144)) and not (inputs(63));
    layer0_outputs(6305) <= inputs(67);
    layer0_outputs(6306) <= not((inputs(169)) or (inputs(61)));
    layer0_outputs(6307) <= (inputs(176)) and not (inputs(116));
    layer0_outputs(6308) <= inputs(178);
    layer0_outputs(6309) <= not(inputs(197)) or (inputs(19));
    layer0_outputs(6310) <= '1';
    layer0_outputs(6311) <= not((inputs(87)) xor (inputs(134)));
    layer0_outputs(6312) <= not(inputs(109));
    layer0_outputs(6313) <= (inputs(157)) xor (inputs(19));
    layer0_outputs(6314) <= not(inputs(158));
    layer0_outputs(6315) <= inputs(27);
    layer0_outputs(6316) <= (inputs(193)) and not (inputs(30));
    layer0_outputs(6317) <= '0';
    layer0_outputs(6318) <= not(inputs(93)) or (inputs(112));
    layer0_outputs(6319) <= (inputs(86)) or (inputs(163));
    layer0_outputs(6320) <= not(inputs(83)) or (inputs(16));
    layer0_outputs(6321) <= inputs(62);
    layer0_outputs(6322) <= not(inputs(66));
    layer0_outputs(6323) <= (inputs(141)) and not (inputs(44));
    layer0_outputs(6324) <= (inputs(51)) and not (inputs(244));
    layer0_outputs(6325) <= inputs(83);
    layer0_outputs(6326) <= inputs(102);
    layer0_outputs(6327) <= (inputs(43)) and not (inputs(121));
    layer0_outputs(6328) <= not((inputs(87)) or (inputs(11)));
    layer0_outputs(6329) <= inputs(139);
    layer0_outputs(6330) <= inputs(155);
    layer0_outputs(6331) <= not(inputs(123));
    layer0_outputs(6332) <= (inputs(139)) xor (inputs(78));
    layer0_outputs(6333) <= (inputs(62)) xor (inputs(69));
    layer0_outputs(6334) <= (inputs(174)) and not (inputs(77));
    layer0_outputs(6335) <= '0';
    layer0_outputs(6336) <= inputs(229);
    layer0_outputs(6337) <= not(inputs(18));
    layer0_outputs(6338) <= (inputs(173)) or (inputs(180));
    layer0_outputs(6339) <= not(inputs(12));
    layer0_outputs(6340) <= inputs(85);
    layer0_outputs(6341) <= not((inputs(12)) and (inputs(63)));
    layer0_outputs(6342) <= not((inputs(242)) or (inputs(166)));
    layer0_outputs(6343) <= not(inputs(110));
    layer0_outputs(6344) <= '0';
    layer0_outputs(6345) <= not((inputs(202)) or (inputs(143)));
    layer0_outputs(6346) <= (inputs(25)) and not (inputs(85));
    layer0_outputs(6347) <= not(inputs(28));
    layer0_outputs(6348) <= '1';
    layer0_outputs(6349) <= not(inputs(93));
    layer0_outputs(6350) <= not(inputs(128)) or (inputs(8));
    layer0_outputs(6351) <= (inputs(210)) and (inputs(36));
    layer0_outputs(6352) <= (inputs(233)) or (inputs(176));
    layer0_outputs(6353) <= (inputs(5)) and (inputs(248));
    layer0_outputs(6354) <= not((inputs(235)) or (inputs(232)));
    layer0_outputs(6355) <= inputs(77);
    layer0_outputs(6356) <= not(inputs(91));
    layer0_outputs(6357) <= not((inputs(184)) and (inputs(255)));
    layer0_outputs(6358) <= not(inputs(120));
    layer0_outputs(6359) <= not(inputs(16));
    layer0_outputs(6360) <= not((inputs(228)) and (inputs(17)));
    layer0_outputs(6361) <= (inputs(233)) and not (inputs(210));
    layer0_outputs(6362) <= not(inputs(157)) or (inputs(49));
    layer0_outputs(6363) <= inputs(208);
    layer0_outputs(6364) <= (inputs(200)) or (inputs(214));
    layer0_outputs(6365) <= '1';
    layer0_outputs(6366) <= '1';
    layer0_outputs(6367) <= not((inputs(32)) xor (inputs(236)));
    layer0_outputs(6368) <= (inputs(36)) and not (inputs(39));
    layer0_outputs(6369) <= not(inputs(26)) or (inputs(1));
    layer0_outputs(6370) <= inputs(70);
    layer0_outputs(6371) <= inputs(123);
    layer0_outputs(6372) <= not((inputs(129)) or (inputs(169)));
    layer0_outputs(6373) <= not(inputs(94));
    layer0_outputs(6374) <= not(inputs(118));
    layer0_outputs(6375) <= (inputs(20)) and not (inputs(28));
    layer0_outputs(6376) <= not(inputs(149));
    layer0_outputs(6377) <= not(inputs(221)) or (inputs(113));
    layer0_outputs(6378) <= (inputs(41)) or (inputs(231));
    layer0_outputs(6379) <= not(inputs(171)) or (inputs(20));
    layer0_outputs(6380) <= (inputs(26)) and not (inputs(135));
    layer0_outputs(6381) <= not(inputs(140));
    layer0_outputs(6382) <= inputs(116);
    layer0_outputs(6383) <= (inputs(124)) and not (inputs(66));
    layer0_outputs(6384) <= '0';
    layer0_outputs(6385) <= inputs(160);
    layer0_outputs(6386) <= (inputs(43)) and (inputs(185));
    layer0_outputs(6387) <= '0';
    layer0_outputs(6388) <= (inputs(217)) and not (inputs(253));
    layer0_outputs(6389) <= not(inputs(240));
    layer0_outputs(6390) <= not((inputs(225)) xor (inputs(195)));
    layer0_outputs(6391) <= inputs(198);
    layer0_outputs(6392) <= inputs(48);
    layer0_outputs(6393) <= not(inputs(173));
    layer0_outputs(6394) <= (inputs(200)) and not (inputs(53));
    layer0_outputs(6395) <= (inputs(27)) or (inputs(60));
    layer0_outputs(6396) <= not(inputs(209));
    layer0_outputs(6397) <= inputs(115);
    layer0_outputs(6398) <= '1';
    layer0_outputs(6399) <= (inputs(5)) and (inputs(225));
    layer0_outputs(6400) <= not(inputs(163)) or (inputs(144));
    layer0_outputs(6401) <= inputs(9);
    layer0_outputs(6402) <= not(inputs(46));
    layer0_outputs(6403) <= not((inputs(224)) and (inputs(96)));
    layer0_outputs(6404) <= not((inputs(133)) or (inputs(206)));
    layer0_outputs(6405) <= (inputs(240)) and not (inputs(190));
    layer0_outputs(6406) <= inputs(73);
    layer0_outputs(6407) <= inputs(93);
    layer0_outputs(6408) <= not((inputs(116)) and (inputs(44)));
    layer0_outputs(6409) <= not(inputs(201));
    layer0_outputs(6410) <= (inputs(122)) and not (inputs(240));
    layer0_outputs(6411) <= inputs(133);
    layer0_outputs(6412) <= not(inputs(154));
    layer0_outputs(6413) <= not(inputs(207));
    layer0_outputs(6414) <= inputs(83);
    layer0_outputs(6415) <= not(inputs(223)) or (inputs(228));
    layer0_outputs(6416) <= not(inputs(164));
    layer0_outputs(6417) <= (inputs(4)) and not (inputs(158));
    layer0_outputs(6418) <= not(inputs(50));
    layer0_outputs(6419) <= inputs(68);
    layer0_outputs(6420) <= (inputs(242)) and not (inputs(242));
    layer0_outputs(6421) <= inputs(161);
    layer0_outputs(6422) <= (inputs(192)) and (inputs(2));
    layer0_outputs(6423) <= not(inputs(244));
    layer0_outputs(6424) <= inputs(175);
    layer0_outputs(6425) <= (inputs(105)) and not (inputs(220));
    layer0_outputs(6426) <= inputs(22);
    layer0_outputs(6427) <= (inputs(228)) or (inputs(56));
    layer0_outputs(6428) <= inputs(112);
    layer0_outputs(6429) <= not(inputs(114));
    layer0_outputs(6430) <= (inputs(216)) and (inputs(200));
    layer0_outputs(6431) <= not((inputs(53)) or (inputs(53)));
    layer0_outputs(6432) <= inputs(224);
    layer0_outputs(6433) <= '1';
    layer0_outputs(6434) <= '0';
    layer0_outputs(6435) <= (inputs(58)) and not (inputs(246));
    layer0_outputs(6436) <= not((inputs(236)) or (inputs(147)));
    layer0_outputs(6437) <= '0';
    layer0_outputs(6438) <= (inputs(220)) and (inputs(51));
    layer0_outputs(6439) <= (inputs(40)) or (inputs(255));
    layer0_outputs(6440) <= inputs(101);
    layer0_outputs(6441) <= not(inputs(215));
    layer0_outputs(6442) <= (inputs(225)) and (inputs(104));
    layer0_outputs(6443) <= not(inputs(99));
    layer0_outputs(6444) <= not((inputs(253)) and (inputs(70)));
    layer0_outputs(6445) <= (inputs(134)) or (inputs(248));
    layer0_outputs(6446) <= inputs(231);
    layer0_outputs(6447) <= not((inputs(156)) or (inputs(157)));
    layer0_outputs(6448) <= not((inputs(222)) xor (inputs(53)));
    layer0_outputs(6449) <= not(inputs(124));
    layer0_outputs(6450) <= not((inputs(12)) or (inputs(7)));
    layer0_outputs(6451) <= not(inputs(81));
    layer0_outputs(6452) <= not(inputs(133)) or (inputs(140));
    layer0_outputs(6453) <= inputs(234);
    layer0_outputs(6454) <= not((inputs(54)) or (inputs(189)));
    layer0_outputs(6455) <= (inputs(248)) or (inputs(177));
    layer0_outputs(6456) <= (inputs(208)) or (inputs(194));
    layer0_outputs(6457) <= not(inputs(165));
    layer0_outputs(6458) <= inputs(228);
    layer0_outputs(6459) <= (inputs(223)) or (inputs(56));
    layer0_outputs(6460) <= not(inputs(249));
    layer0_outputs(6461) <= not(inputs(156)) or (inputs(132));
    layer0_outputs(6462) <= (inputs(0)) and (inputs(173));
    layer0_outputs(6463) <= not((inputs(203)) and (inputs(115)));
    layer0_outputs(6464) <= not(inputs(243)) or (inputs(227));
    layer0_outputs(6465) <= not((inputs(145)) xor (inputs(163)));
    layer0_outputs(6466) <= '1';
    layer0_outputs(6467) <= inputs(106);
    layer0_outputs(6468) <= not(inputs(61)) or (inputs(190));
    layer0_outputs(6469) <= inputs(136);
    layer0_outputs(6470) <= '0';
    layer0_outputs(6471) <= (inputs(205)) and not (inputs(11));
    layer0_outputs(6472) <= not((inputs(82)) xor (inputs(75)));
    layer0_outputs(6473) <= not(inputs(56));
    layer0_outputs(6474) <= not(inputs(156)) or (inputs(123));
    layer0_outputs(6475) <= not(inputs(208));
    layer0_outputs(6476) <= not(inputs(199));
    layer0_outputs(6477) <= '0';
    layer0_outputs(6478) <= not(inputs(23));
    layer0_outputs(6479) <= (inputs(160)) and not (inputs(64));
    layer0_outputs(6480) <= '1';
    layer0_outputs(6481) <= not((inputs(251)) or (inputs(252)));
    layer0_outputs(6482) <= (inputs(3)) and not (inputs(52));
    layer0_outputs(6483) <= inputs(33);
    layer0_outputs(6484) <= not(inputs(126));
    layer0_outputs(6485) <= not(inputs(153));
    layer0_outputs(6486) <= not((inputs(9)) xor (inputs(20)));
    layer0_outputs(6487) <= (inputs(66)) and not (inputs(187));
    layer0_outputs(6488) <= inputs(220);
    layer0_outputs(6489) <= not(inputs(57));
    layer0_outputs(6490) <= (inputs(247)) and not (inputs(106));
    layer0_outputs(6491) <= inputs(186);
    layer0_outputs(6492) <= inputs(97);
    layer0_outputs(6493) <= not(inputs(81));
    layer0_outputs(6494) <= not(inputs(144));
    layer0_outputs(6495) <= (inputs(171)) and not (inputs(163));
    layer0_outputs(6496) <= (inputs(167)) and not (inputs(164));
    layer0_outputs(6497) <= not(inputs(59));
    layer0_outputs(6498) <= not((inputs(108)) xor (inputs(187)));
    layer0_outputs(6499) <= '0';
    layer0_outputs(6500) <= not(inputs(44));
    layer0_outputs(6501) <= not(inputs(41)) or (inputs(0));
    layer0_outputs(6502) <= (inputs(206)) and not (inputs(232));
    layer0_outputs(6503) <= (inputs(160)) or (inputs(175));
    layer0_outputs(6504) <= not(inputs(82)) or (inputs(242));
    layer0_outputs(6505) <= not((inputs(65)) and (inputs(129)));
    layer0_outputs(6506) <= inputs(165);
    layer0_outputs(6507) <= not(inputs(246)) or (inputs(34));
    layer0_outputs(6508) <= inputs(210);
    layer0_outputs(6509) <= inputs(163);
    layer0_outputs(6510) <= (inputs(16)) or (inputs(98));
    layer0_outputs(6511) <= not(inputs(173));
    layer0_outputs(6512) <= inputs(23);
    layer0_outputs(6513) <= (inputs(180)) and not (inputs(166));
    layer0_outputs(6514) <= inputs(245);
    layer0_outputs(6515) <= not(inputs(40));
    layer0_outputs(6516) <= inputs(177);
    layer0_outputs(6517) <= not((inputs(29)) or (inputs(90)));
    layer0_outputs(6518) <= inputs(23);
    layer0_outputs(6519) <= inputs(76);
    layer0_outputs(6520) <= not((inputs(3)) xor (inputs(119)));
    layer0_outputs(6521) <= inputs(238);
    layer0_outputs(6522) <= inputs(165);
    layer0_outputs(6523) <= not(inputs(159));
    layer0_outputs(6524) <= not(inputs(167)) or (inputs(48));
    layer0_outputs(6525) <= not(inputs(91));
    layer0_outputs(6526) <= (inputs(76)) or (inputs(90));
    layer0_outputs(6527) <= not((inputs(47)) or (inputs(123)));
    layer0_outputs(6528) <= not(inputs(76)) or (inputs(32));
    layer0_outputs(6529) <= not(inputs(154));
    layer0_outputs(6530) <= not(inputs(197));
    layer0_outputs(6531) <= not(inputs(61));
    layer0_outputs(6532) <= inputs(54);
    layer0_outputs(6533) <= not(inputs(228)) or (inputs(183));
    layer0_outputs(6534) <= not(inputs(73));
    layer0_outputs(6535) <= (inputs(137)) and (inputs(44));
    layer0_outputs(6536) <= (inputs(20)) or (inputs(237));
    layer0_outputs(6537) <= (inputs(248)) or (inputs(100));
    layer0_outputs(6538) <= '1';
    layer0_outputs(6539) <= not(inputs(145));
    layer0_outputs(6540) <= not(inputs(161));
    layer0_outputs(6541) <= inputs(131);
    layer0_outputs(6542) <= not(inputs(182));
    layer0_outputs(6543) <= not((inputs(202)) or (inputs(212)));
    layer0_outputs(6544) <= inputs(125);
    layer0_outputs(6545) <= (inputs(137)) xor (inputs(76));
    layer0_outputs(6546) <= inputs(199);
    layer0_outputs(6547) <= inputs(187);
    layer0_outputs(6548) <= (inputs(124)) and not (inputs(122));
    layer0_outputs(6549) <= inputs(81);
    layer0_outputs(6550) <= not(inputs(1)) or (inputs(68));
    layer0_outputs(6551) <= (inputs(188)) or (inputs(101));
    layer0_outputs(6552) <= '1';
    layer0_outputs(6553) <= '1';
    layer0_outputs(6554) <= inputs(40);
    layer0_outputs(6555) <= not((inputs(246)) or (inputs(62)));
    layer0_outputs(6556) <= (inputs(77)) and not (inputs(130));
    layer0_outputs(6557) <= (inputs(253)) or (inputs(32));
    layer0_outputs(6558) <= inputs(48);
    layer0_outputs(6559) <= not(inputs(14)) or (inputs(61));
    layer0_outputs(6560) <= (inputs(246)) and not (inputs(54));
    layer0_outputs(6561) <= (inputs(48)) or (inputs(195));
    layer0_outputs(6562) <= '0';
    layer0_outputs(6563) <= not((inputs(49)) or (inputs(103)));
    layer0_outputs(6564) <= not(inputs(182)) or (inputs(167));
    layer0_outputs(6565) <= inputs(82);
    layer0_outputs(6566) <= not((inputs(94)) or (inputs(21)));
    layer0_outputs(6567) <= (inputs(93)) or (inputs(39));
    layer0_outputs(6568) <= (inputs(138)) or (inputs(190));
    layer0_outputs(6569) <= (inputs(88)) or (inputs(87));
    layer0_outputs(6570) <= not(inputs(248));
    layer0_outputs(6571) <= not(inputs(149));
    layer0_outputs(6572) <= inputs(252);
    layer0_outputs(6573) <= (inputs(220)) xor (inputs(235));
    layer0_outputs(6574) <= (inputs(53)) and not (inputs(103));
    layer0_outputs(6575) <= not(inputs(56)) or (inputs(31));
    layer0_outputs(6576) <= (inputs(5)) or (inputs(118));
    layer0_outputs(6577) <= (inputs(150)) and not (inputs(218));
    layer0_outputs(6578) <= '1';
    layer0_outputs(6579) <= '0';
    layer0_outputs(6580) <= '0';
    layer0_outputs(6581) <= not(inputs(145));
    layer0_outputs(6582) <= (inputs(44)) and (inputs(40));
    layer0_outputs(6583) <= not((inputs(144)) or (inputs(47)));
    layer0_outputs(6584) <= (inputs(141)) or (inputs(172));
    layer0_outputs(6585) <= not(inputs(110));
    layer0_outputs(6586) <= inputs(196);
    layer0_outputs(6587) <= not((inputs(30)) or (inputs(173)));
    layer0_outputs(6588) <= not((inputs(226)) or (inputs(242)));
    layer0_outputs(6589) <= not(inputs(62));
    layer0_outputs(6590) <= (inputs(207)) or (inputs(139));
    layer0_outputs(6591) <= inputs(168);
    layer0_outputs(6592) <= (inputs(149)) xor (inputs(226));
    layer0_outputs(6593) <= inputs(44);
    layer0_outputs(6594) <= (inputs(29)) or (inputs(82));
    layer0_outputs(6595) <= (inputs(121)) and not (inputs(16));
    layer0_outputs(6596) <= (inputs(186)) or (inputs(125));
    layer0_outputs(6597) <= not(inputs(55));
    layer0_outputs(6598) <= inputs(148);
    layer0_outputs(6599) <= (inputs(28)) and (inputs(162));
    layer0_outputs(6600) <= inputs(195);
    layer0_outputs(6601) <= (inputs(60)) and not (inputs(226));
    layer0_outputs(6602) <= not(inputs(134)) or (inputs(62));
    layer0_outputs(6603) <= (inputs(47)) and not (inputs(106));
    layer0_outputs(6604) <= (inputs(3)) or (inputs(95));
    layer0_outputs(6605) <= not((inputs(138)) and (inputs(250)));
    layer0_outputs(6606) <= not(inputs(216)) or (inputs(123));
    layer0_outputs(6607) <= not(inputs(131));
    layer0_outputs(6608) <= not((inputs(205)) xor (inputs(124)));
    layer0_outputs(6609) <= inputs(219);
    layer0_outputs(6610) <= not(inputs(25)) or (inputs(188));
    layer0_outputs(6611) <= (inputs(168)) or (inputs(134));
    layer0_outputs(6612) <= not((inputs(170)) or (inputs(46)));
    layer0_outputs(6613) <= not(inputs(217)) or (inputs(113));
    layer0_outputs(6614) <= not((inputs(16)) and (inputs(30)));
    layer0_outputs(6615) <= inputs(71);
    layer0_outputs(6616) <= (inputs(92)) and not (inputs(151));
    layer0_outputs(6617) <= not((inputs(212)) or (inputs(210)));
    layer0_outputs(6618) <= not(inputs(87)) or (inputs(196));
    layer0_outputs(6619) <= not(inputs(92));
    layer0_outputs(6620) <= (inputs(22)) xor (inputs(147));
    layer0_outputs(6621) <= (inputs(146)) and (inputs(76));
    layer0_outputs(6622) <= (inputs(169)) and not (inputs(150));
    layer0_outputs(6623) <= (inputs(90)) and not (inputs(187));
    layer0_outputs(6624) <= inputs(23);
    layer0_outputs(6625) <= inputs(85);
    layer0_outputs(6626) <= (inputs(139)) and (inputs(126));
    layer0_outputs(6627) <= '0';
    layer0_outputs(6628) <= not((inputs(60)) or (inputs(208)));
    layer0_outputs(6629) <= not((inputs(179)) and (inputs(0)));
    layer0_outputs(6630) <= (inputs(121)) or (inputs(208));
    layer0_outputs(6631) <= not(inputs(52)) or (inputs(62));
    layer0_outputs(6632) <= not(inputs(210));
    layer0_outputs(6633) <= inputs(108);
    layer0_outputs(6634) <= not((inputs(247)) and (inputs(172)));
    layer0_outputs(6635) <= '0';
    layer0_outputs(6636) <= (inputs(206)) and not (inputs(213));
    layer0_outputs(6637) <= (inputs(9)) or (inputs(138));
    layer0_outputs(6638) <= not((inputs(126)) or (inputs(213)));
    layer0_outputs(6639) <= inputs(110);
    layer0_outputs(6640) <= '1';
    layer0_outputs(6641) <= (inputs(180)) and not (inputs(96));
    layer0_outputs(6642) <= (inputs(55)) and not (inputs(50));
    layer0_outputs(6643) <= (inputs(75)) or (inputs(31));
    layer0_outputs(6644) <= not(inputs(109));
    layer0_outputs(6645) <= inputs(123);
    layer0_outputs(6646) <= not(inputs(20));
    layer0_outputs(6647) <= (inputs(248)) and (inputs(176));
    layer0_outputs(6648) <= inputs(174);
    layer0_outputs(6649) <= not(inputs(174)) or (inputs(1));
    layer0_outputs(6650) <= not(inputs(114)) or (inputs(202));
    layer0_outputs(6651) <= (inputs(35)) or (inputs(77));
    layer0_outputs(6652) <= inputs(135);
    layer0_outputs(6653) <= (inputs(178)) and not (inputs(40));
    layer0_outputs(6654) <= not(inputs(113)) or (inputs(58));
    layer0_outputs(6655) <= (inputs(187)) and not (inputs(110));
    layer0_outputs(6656) <= not((inputs(151)) or (inputs(181)));
    layer0_outputs(6657) <= inputs(127);
    layer0_outputs(6658) <= inputs(85);
    layer0_outputs(6659) <= inputs(39);
    layer0_outputs(6660) <= not((inputs(127)) and (inputs(55)));
    layer0_outputs(6661) <= (inputs(68)) or (inputs(122));
    layer0_outputs(6662) <= not((inputs(52)) or (inputs(45)));
    layer0_outputs(6663) <= (inputs(35)) or (inputs(205));
    layer0_outputs(6664) <= not(inputs(212));
    layer0_outputs(6665) <= inputs(207);
    layer0_outputs(6666) <= not((inputs(74)) and (inputs(8)));
    layer0_outputs(6667) <= (inputs(154)) or (inputs(220));
    layer0_outputs(6668) <= (inputs(222)) or (inputs(166));
    layer0_outputs(6669) <= inputs(155);
    layer0_outputs(6670) <= inputs(56);
    layer0_outputs(6671) <= '1';
    layer0_outputs(6672) <= not(inputs(151)) or (inputs(202));
    layer0_outputs(6673) <= inputs(73);
    layer0_outputs(6674) <= inputs(212);
    layer0_outputs(6675) <= (inputs(10)) or (inputs(128));
    layer0_outputs(6676) <= (inputs(78)) xor (inputs(165));
    layer0_outputs(6677) <= (inputs(77)) xor (inputs(215));
    layer0_outputs(6678) <= not(inputs(210));
    layer0_outputs(6679) <= (inputs(136)) and not (inputs(76));
    layer0_outputs(6680) <= (inputs(123)) or (inputs(13));
    layer0_outputs(6681) <= not(inputs(127)) or (inputs(103));
    layer0_outputs(6682) <= not((inputs(190)) or (inputs(30)));
    layer0_outputs(6683) <= (inputs(245)) and not (inputs(207));
    layer0_outputs(6684) <= not(inputs(97)) or (inputs(53));
    layer0_outputs(6685) <= not((inputs(183)) and (inputs(52)));
    layer0_outputs(6686) <= not(inputs(145));
    layer0_outputs(6687) <= '0';
    layer0_outputs(6688) <= not(inputs(175));
    layer0_outputs(6689) <= not(inputs(110));
    layer0_outputs(6690) <= inputs(197);
    layer0_outputs(6691) <= (inputs(183)) and (inputs(188));
    layer0_outputs(6692) <= (inputs(59)) and (inputs(148));
    layer0_outputs(6693) <= inputs(168);
    layer0_outputs(6694) <= '0';
    layer0_outputs(6695) <= (inputs(166)) and not (inputs(183));
    layer0_outputs(6696) <= inputs(106);
    layer0_outputs(6697) <= not(inputs(186));
    layer0_outputs(6698) <= '0';
    layer0_outputs(6699) <= (inputs(175)) and (inputs(152));
    layer0_outputs(6700) <= inputs(69);
    layer0_outputs(6701) <= not(inputs(124));
    layer0_outputs(6702) <= not(inputs(10)) or (inputs(2));
    layer0_outputs(6703) <= inputs(84);
    layer0_outputs(6704) <= not(inputs(60)) or (inputs(222));
    layer0_outputs(6705) <= (inputs(69)) and not (inputs(218));
    layer0_outputs(6706) <= not(inputs(4));
    layer0_outputs(6707) <= (inputs(227)) and (inputs(230));
    layer0_outputs(6708) <= (inputs(30)) and not (inputs(226));
    layer0_outputs(6709) <= not((inputs(231)) xor (inputs(142)));
    layer0_outputs(6710) <= inputs(110);
    layer0_outputs(6711) <= not(inputs(219));
    layer0_outputs(6712) <= (inputs(158)) or (inputs(98));
    layer0_outputs(6713) <= not(inputs(113));
    layer0_outputs(6714) <= (inputs(127)) and not (inputs(0));
    layer0_outputs(6715) <= not(inputs(138));
    layer0_outputs(6716) <= not((inputs(134)) or (inputs(122)));
    layer0_outputs(6717) <= (inputs(166)) and not (inputs(110));
    layer0_outputs(6718) <= (inputs(124)) and not (inputs(12));
    layer0_outputs(6719) <= (inputs(63)) or (inputs(79));
    layer0_outputs(6720) <= (inputs(113)) and not (inputs(109));
    layer0_outputs(6721) <= (inputs(230)) or (inputs(2));
    layer0_outputs(6722) <= not(inputs(61));
    layer0_outputs(6723) <= (inputs(228)) and (inputs(162));
    layer0_outputs(6724) <= '0';
    layer0_outputs(6725) <= not(inputs(221));
    layer0_outputs(6726) <= not(inputs(39)) or (inputs(135));
    layer0_outputs(6727) <= (inputs(192)) and not (inputs(172));
    layer0_outputs(6728) <= inputs(52);
    layer0_outputs(6729) <= (inputs(28)) and (inputs(118));
    layer0_outputs(6730) <= not((inputs(223)) and (inputs(31)));
    layer0_outputs(6731) <= not((inputs(171)) xor (inputs(147)));
    layer0_outputs(6732) <= not((inputs(77)) or (inputs(139)));
    layer0_outputs(6733) <= not(inputs(69)) or (inputs(223));
    layer0_outputs(6734) <= (inputs(182)) and not (inputs(40));
    layer0_outputs(6735) <= '1';
    layer0_outputs(6736) <= '1';
    layer0_outputs(6737) <= not((inputs(175)) or (inputs(90)));
    layer0_outputs(6738) <= not(inputs(246)) or (inputs(221));
    layer0_outputs(6739) <= (inputs(82)) xor (inputs(143));
    layer0_outputs(6740) <= not((inputs(164)) or (inputs(150)));
    layer0_outputs(6741) <= inputs(252);
    layer0_outputs(6742) <= inputs(184);
    layer0_outputs(6743) <= not(inputs(189));
    layer0_outputs(6744) <= not(inputs(119));
    layer0_outputs(6745) <= (inputs(158)) and not (inputs(76));
    layer0_outputs(6746) <= (inputs(21)) and not (inputs(245));
    layer0_outputs(6747) <= not(inputs(78));
    layer0_outputs(6748) <= not(inputs(188));
    layer0_outputs(6749) <= not(inputs(244)) or (inputs(201));
    layer0_outputs(6750) <= inputs(100);
    layer0_outputs(6751) <= (inputs(89)) and (inputs(96));
    layer0_outputs(6752) <= not((inputs(137)) or (inputs(51)));
    layer0_outputs(6753) <= not((inputs(135)) or (inputs(164)));
    layer0_outputs(6754) <= not((inputs(79)) or (inputs(5)));
    layer0_outputs(6755) <= inputs(41);
    layer0_outputs(6756) <= not(inputs(69));
    layer0_outputs(6757) <= '0';
    layer0_outputs(6758) <= not(inputs(254));
    layer0_outputs(6759) <= not(inputs(131));
    layer0_outputs(6760) <= not((inputs(101)) or (inputs(31)));
    layer0_outputs(6761) <= not(inputs(13)) or (inputs(102));
    layer0_outputs(6762) <= not(inputs(73));
    layer0_outputs(6763) <= not(inputs(232)) or (inputs(182));
    layer0_outputs(6764) <= (inputs(53)) and not (inputs(48));
    layer0_outputs(6765) <= inputs(234);
    layer0_outputs(6766) <= not(inputs(80)) or (inputs(90));
    layer0_outputs(6767) <= inputs(170);
    layer0_outputs(6768) <= (inputs(145)) or (inputs(156));
    layer0_outputs(6769) <= (inputs(20)) or (inputs(73));
    layer0_outputs(6770) <= '0';
    layer0_outputs(6771) <= (inputs(81)) and not (inputs(232));
    layer0_outputs(6772) <= (inputs(25)) or (inputs(193));
    layer0_outputs(6773) <= not((inputs(213)) or (inputs(228)));
    layer0_outputs(6774) <= not(inputs(190)) or (inputs(165));
    layer0_outputs(6775) <= not((inputs(180)) or (inputs(93)));
    layer0_outputs(6776) <= not(inputs(123)) or (inputs(194));
    layer0_outputs(6777) <= not(inputs(9));
    layer0_outputs(6778) <= (inputs(11)) and (inputs(28));
    layer0_outputs(6779) <= inputs(182);
    layer0_outputs(6780) <= not(inputs(157));
    layer0_outputs(6781) <= (inputs(153)) and not (inputs(23));
    layer0_outputs(6782) <= not((inputs(221)) or (inputs(168)));
    layer0_outputs(6783) <= '0';
    layer0_outputs(6784) <= (inputs(30)) or (inputs(254));
    layer0_outputs(6785) <= '1';
    layer0_outputs(6786) <= not(inputs(67));
    layer0_outputs(6787) <= not(inputs(192)) or (inputs(252));
    layer0_outputs(6788) <= not((inputs(33)) or (inputs(59)));
    layer0_outputs(6789) <= not(inputs(28)) or (inputs(101));
    layer0_outputs(6790) <= inputs(141);
    layer0_outputs(6791) <= not(inputs(42)) or (inputs(161));
    layer0_outputs(6792) <= (inputs(201)) and (inputs(125));
    layer0_outputs(6793) <= inputs(77);
    layer0_outputs(6794) <= not((inputs(67)) or (inputs(254)));
    layer0_outputs(6795) <= (inputs(100)) or (inputs(75));
    layer0_outputs(6796) <= (inputs(139)) or (inputs(154));
    layer0_outputs(6797) <= not((inputs(223)) and (inputs(12)));
    layer0_outputs(6798) <= not(inputs(221));
    layer0_outputs(6799) <= not(inputs(255)) or (inputs(46));
    layer0_outputs(6800) <= not(inputs(235)) or (inputs(148));
    layer0_outputs(6801) <= (inputs(238)) and (inputs(42));
    layer0_outputs(6802) <= (inputs(40)) xor (inputs(8));
    layer0_outputs(6803) <= not(inputs(66));
    layer0_outputs(6804) <= (inputs(160)) xor (inputs(181));
    layer0_outputs(6805) <= (inputs(234)) or (inputs(109));
    layer0_outputs(6806) <= not(inputs(158)) or (inputs(25));
    layer0_outputs(6807) <= not(inputs(193));
    layer0_outputs(6808) <= inputs(187);
    layer0_outputs(6809) <= not((inputs(158)) and (inputs(35)));
    layer0_outputs(6810) <= (inputs(160)) and (inputs(195));
    layer0_outputs(6811) <= (inputs(194)) or (inputs(219));
    layer0_outputs(6812) <= inputs(188);
    layer0_outputs(6813) <= not((inputs(234)) and (inputs(17)));
    layer0_outputs(6814) <= '1';
    layer0_outputs(6815) <= (inputs(111)) or (inputs(75));
    layer0_outputs(6816) <= not(inputs(218));
    layer0_outputs(6817) <= (inputs(227)) and not (inputs(0));
    layer0_outputs(6818) <= '1';
    layer0_outputs(6819) <= inputs(31);
    layer0_outputs(6820) <= (inputs(147)) and not (inputs(119));
    layer0_outputs(6821) <= not(inputs(85));
    layer0_outputs(6822) <= inputs(88);
    layer0_outputs(6823) <= not(inputs(23));
    layer0_outputs(6824) <= not((inputs(80)) or (inputs(212)));
    layer0_outputs(6825) <= (inputs(71)) xor (inputs(85));
    layer0_outputs(6826) <= not((inputs(83)) or (inputs(84)));
    layer0_outputs(6827) <= (inputs(142)) or (inputs(21));
    layer0_outputs(6828) <= (inputs(188)) and not (inputs(140));
    layer0_outputs(6829) <= (inputs(195)) or (inputs(190));
    layer0_outputs(6830) <= not(inputs(7)) or (inputs(227));
    layer0_outputs(6831) <= not((inputs(177)) or (inputs(220)));
    layer0_outputs(6832) <= not((inputs(219)) or (inputs(170)));
    layer0_outputs(6833) <= '1';
    layer0_outputs(6834) <= (inputs(88)) or (inputs(210));
    layer0_outputs(6835) <= inputs(189);
    layer0_outputs(6836) <= (inputs(135)) or (inputs(28));
    layer0_outputs(6837) <= (inputs(229)) and not (inputs(2));
    layer0_outputs(6838) <= (inputs(213)) and not (inputs(46));
    layer0_outputs(6839) <= inputs(95);
    layer0_outputs(6840) <= not((inputs(203)) xor (inputs(252)));
    layer0_outputs(6841) <= not((inputs(123)) and (inputs(40)));
    layer0_outputs(6842) <= not(inputs(217));
    layer0_outputs(6843) <= not(inputs(229));
    layer0_outputs(6844) <= inputs(234);
    layer0_outputs(6845) <= (inputs(224)) and (inputs(130));
    layer0_outputs(6846) <= inputs(136);
    layer0_outputs(6847) <= not((inputs(214)) or (inputs(52)));
    layer0_outputs(6848) <= '1';
    layer0_outputs(6849) <= inputs(27);
    layer0_outputs(6850) <= not((inputs(64)) or (inputs(140)));
    layer0_outputs(6851) <= not(inputs(151));
    layer0_outputs(6852) <= inputs(111);
    layer0_outputs(6853) <= (inputs(230)) and not (inputs(92));
    layer0_outputs(6854) <= (inputs(221)) or (inputs(177));
    layer0_outputs(6855) <= not((inputs(0)) xor (inputs(164)));
    layer0_outputs(6856) <= '1';
    layer0_outputs(6857) <= not((inputs(165)) or (inputs(174)));
    layer0_outputs(6858) <= not((inputs(240)) and (inputs(21)));
    layer0_outputs(6859) <= not(inputs(57)) or (inputs(166));
    layer0_outputs(6860) <= inputs(76);
    layer0_outputs(6861) <= (inputs(131)) or (inputs(95));
    layer0_outputs(6862) <= not(inputs(10));
    layer0_outputs(6863) <= (inputs(60)) or (inputs(227));
    layer0_outputs(6864) <= not(inputs(5));
    layer0_outputs(6865) <= not((inputs(218)) or (inputs(105)));
    layer0_outputs(6866) <= (inputs(252)) or (inputs(148));
    layer0_outputs(6867) <= not(inputs(115));
    layer0_outputs(6868) <= (inputs(56)) or (inputs(33));
    layer0_outputs(6869) <= (inputs(255)) or (inputs(182));
    layer0_outputs(6870) <= (inputs(124)) xor (inputs(4));
    layer0_outputs(6871) <= not((inputs(27)) or (inputs(138)));
    layer0_outputs(6872) <= not(inputs(9));
    layer0_outputs(6873) <= '1';
    layer0_outputs(6874) <= inputs(211);
    layer0_outputs(6875) <= (inputs(53)) and not (inputs(179));
    layer0_outputs(6876) <= not(inputs(213)) or (inputs(243));
    layer0_outputs(6877) <= not(inputs(161)) or (inputs(15));
    layer0_outputs(6878) <= (inputs(44)) xor (inputs(19));
    layer0_outputs(6879) <= '0';
    layer0_outputs(6880) <= inputs(149);
    layer0_outputs(6881) <= (inputs(84)) and (inputs(36));
    layer0_outputs(6882) <= '0';
    layer0_outputs(6883) <= inputs(134);
    layer0_outputs(6884) <= (inputs(241)) and not (inputs(63));
    layer0_outputs(6885) <= (inputs(18)) and (inputs(26));
    layer0_outputs(6886) <= (inputs(145)) and not (inputs(186));
    layer0_outputs(6887) <= (inputs(113)) xor (inputs(114));
    layer0_outputs(6888) <= not(inputs(104));
    layer0_outputs(6889) <= (inputs(252)) or (inputs(81));
    layer0_outputs(6890) <= (inputs(220)) or (inputs(229));
    layer0_outputs(6891) <= not(inputs(28));
    layer0_outputs(6892) <= not(inputs(156)) or (inputs(1));
    layer0_outputs(6893) <= '1';
    layer0_outputs(6894) <= (inputs(235)) and (inputs(153));
    layer0_outputs(6895) <= not(inputs(44)) or (inputs(47));
    layer0_outputs(6896) <= not((inputs(34)) or (inputs(218)));
    layer0_outputs(6897) <= not(inputs(68)) or (inputs(45));
    layer0_outputs(6898) <= not((inputs(85)) and (inputs(200)));
    layer0_outputs(6899) <= (inputs(37)) and not (inputs(207));
    layer0_outputs(6900) <= not(inputs(39));
    layer0_outputs(6901) <= not(inputs(24));
    layer0_outputs(6902) <= (inputs(192)) xor (inputs(243));
    layer0_outputs(6903) <= inputs(30);
    layer0_outputs(6904) <= not(inputs(120)) or (inputs(203));
    layer0_outputs(6905) <= not(inputs(78)) or (inputs(80));
    layer0_outputs(6906) <= not((inputs(247)) or (inputs(188)));
    layer0_outputs(6907) <= not(inputs(98));
    layer0_outputs(6908) <= not((inputs(32)) or (inputs(116)));
    layer0_outputs(6909) <= (inputs(117)) and not (inputs(249));
    layer0_outputs(6910) <= not((inputs(169)) and (inputs(164)));
    layer0_outputs(6911) <= not(inputs(58)) or (inputs(6));
    layer0_outputs(6912) <= not(inputs(54)) or (inputs(149));
    layer0_outputs(6913) <= (inputs(38)) and not (inputs(157));
    layer0_outputs(6914) <= not(inputs(60));
    layer0_outputs(6915) <= not((inputs(94)) or (inputs(244)));
    layer0_outputs(6916) <= (inputs(26)) or (inputs(80));
    layer0_outputs(6917) <= not(inputs(181));
    layer0_outputs(6918) <= not((inputs(55)) and (inputs(54)));
    layer0_outputs(6919) <= not(inputs(6));
    layer0_outputs(6920) <= (inputs(92)) xor (inputs(45));
    layer0_outputs(6921) <= not((inputs(95)) or (inputs(201)));
    layer0_outputs(6922) <= not(inputs(165));
    layer0_outputs(6923) <= (inputs(227)) or (inputs(219));
    layer0_outputs(6924) <= not(inputs(122));
    layer0_outputs(6925) <= not(inputs(234)) or (inputs(63));
    layer0_outputs(6926) <= not(inputs(201));
    layer0_outputs(6927) <= (inputs(101)) and (inputs(82));
    layer0_outputs(6928) <= (inputs(187)) and not (inputs(101));
    layer0_outputs(6929) <= not(inputs(179));
    layer0_outputs(6930) <= (inputs(50)) xor (inputs(20));
    layer0_outputs(6931) <= (inputs(104)) and not (inputs(175));
    layer0_outputs(6932) <= not((inputs(112)) xor (inputs(169)));
    layer0_outputs(6933) <= not((inputs(82)) and (inputs(41)));
    layer0_outputs(6934) <= not(inputs(199));
    layer0_outputs(6935) <= not(inputs(119));
    layer0_outputs(6936) <= not(inputs(196));
    layer0_outputs(6937) <= not(inputs(235)) or (inputs(33));
    layer0_outputs(6938) <= inputs(67);
    layer0_outputs(6939) <= (inputs(166)) and (inputs(123));
    layer0_outputs(6940) <= not(inputs(34));
    layer0_outputs(6941) <= not(inputs(109));
    layer0_outputs(6942) <= not(inputs(218));
    layer0_outputs(6943) <= (inputs(171)) or (inputs(81));
    layer0_outputs(6944) <= not(inputs(24));
    layer0_outputs(6945) <= (inputs(84)) and not (inputs(159));
    layer0_outputs(6946) <= not(inputs(99));
    layer0_outputs(6947) <= not(inputs(217));
    layer0_outputs(6948) <= (inputs(63)) and not (inputs(239));
    layer0_outputs(6949) <= not((inputs(39)) and (inputs(44)));
    layer0_outputs(6950) <= not(inputs(243)) or (inputs(24));
    layer0_outputs(6951) <= (inputs(95)) or (inputs(43));
    layer0_outputs(6952) <= (inputs(70)) xor (inputs(3));
    layer0_outputs(6953) <= inputs(167);
    layer0_outputs(6954) <= not(inputs(106));
    layer0_outputs(6955) <= not((inputs(69)) xor (inputs(49)));
    layer0_outputs(6956) <= (inputs(98)) and not (inputs(170));
    layer0_outputs(6957) <= (inputs(54)) or (inputs(176));
    layer0_outputs(6958) <= (inputs(25)) and (inputs(24));
    layer0_outputs(6959) <= inputs(124);
    layer0_outputs(6960) <= inputs(109);
    layer0_outputs(6961) <= (inputs(122)) or (inputs(246));
    layer0_outputs(6962) <= '1';
    layer0_outputs(6963) <= not(inputs(73)) or (inputs(169));
    layer0_outputs(6964) <= (inputs(249)) and not (inputs(199));
    layer0_outputs(6965) <= (inputs(253)) or (inputs(13));
    layer0_outputs(6966) <= '1';
    layer0_outputs(6967) <= not(inputs(73));
    layer0_outputs(6968) <= not(inputs(45)) or (inputs(87));
    layer0_outputs(6969) <= not((inputs(122)) or (inputs(104)));
    layer0_outputs(6970) <= not(inputs(107)) or (inputs(15));
    layer0_outputs(6971) <= (inputs(97)) and not (inputs(107));
    layer0_outputs(6972) <= not(inputs(74));
    layer0_outputs(6973) <= inputs(58);
    layer0_outputs(6974) <= (inputs(216)) xor (inputs(249));
    layer0_outputs(6975) <= inputs(233);
    layer0_outputs(6976) <= (inputs(45)) and not (inputs(157));
    layer0_outputs(6977) <= (inputs(4)) and (inputs(22));
    layer0_outputs(6978) <= inputs(157);
    layer0_outputs(6979) <= not(inputs(74));
    layer0_outputs(6980) <= not(inputs(8)) or (inputs(84));
    layer0_outputs(6981) <= not(inputs(152)) or (inputs(61));
    layer0_outputs(6982) <= not(inputs(152)) or (inputs(81));
    layer0_outputs(6983) <= inputs(231);
    layer0_outputs(6984) <= (inputs(47)) and not (inputs(174));
    layer0_outputs(6985) <= (inputs(234)) or (inputs(228));
    layer0_outputs(6986) <= '0';
    layer0_outputs(6987) <= '1';
    layer0_outputs(6988) <= (inputs(44)) and (inputs(200));
    layer0_outputs(6989) <= not(inputs(140));
    layer0_outputs(6990) <= (inputs(86)) and not (inputs(49));
    layer0_outputs(6991) <= (inputs(213)) or (inputs(193));
    layer0_outputs(6992) <= (inputs(21)) and (inputs(33));
    layer0_outputs(6993) <= not((inputs(25)) xor (inputs(66)));
    layer0_outputs(6994) <= not(inputs(181));
    layer0_outputs(6995) <= inputs(11);
    layer0_outputs(6996) <= not((inputs(93)) or (inputs(161)));
    layer0_outputs(6997) <= (inputs(115)) and (inputs(124));
    layer0_outputs(6998) <= inputs(104);
    layer0_outputs(6999) <= not(inputs(67)) or (inputs(207));
    layer0_outputs(7000) <= not(inputs(190));
    layer0_outputs(7001) <= not(inputs(21));
    layer0_outputs(7002) <= '0';
    layer0_outputs(7003) <= (inputs(88)) xor (inputs(144));
    layer0_outputs(7004) <= not((inputs(180)) xor (inputs(150)));
    layer0_outputs(7005) <= '0';
    layer0_outputs(7006) <= not(inputs(232));
    layer0_outputs(7007) <= (inputs(151)) xor (inputs(29));
    layer0_outputs(7008) <= not((inputs(56)) xor (inputs(144)));
    layer0_outputs(7009) <= (inputs(255)) xor (inputs(73));
    layer0_outputs(7010) <= not(inputs(179));
    layer0_outputs(7011) <= (inputs(64)) or (inputs(201));
    layer0_outputs(7012) <= (inputs(152)) xor (inputs(88));
    layer0_outputs(7013) <= inputs(222);
    layer0_outputs(7014) <= '0';
    layer0_outputs(7015) <= not(inputs(153));
    layer0_outputs(7016) <= inputs(244);
    layer0_outputs(7017) <= not(inputs(74)) or (inputs(38));
    layer0_outputs(7018) <= not((inputs(50)) or (inputs(198)));
    layer0_outputs(7019) <= not((inputs(123)) or (inputs(145)));
    layer0_outputs(7020) <= '0';
    layer0_outputs(7021) <= (inputs(48)) or (inputs(9));
    layer0_outputs(7022) <= inputs(107);
    layer0_outputs(7023) <= (inputs(140)) or (inputs(176));
    layer0_outputs(7024) <= inputs(32);
    layer0_outputs(7025) <= not(inputs(227));
    layer0_outputs(7026) <= inputs(88);
    layer0_outputs(7027) <= not((inputs(56)) or (inputs(29)));
    layer0_outputs(7028) <= not((inputs(178)) or (inputs(129)));
    layer0_outputs(7029) <= not((inputs(128)) xor (inputs(209)));
    layer0_outputs(7030) <= (inputs(240)) xor (inputs(153));
    layer0_outputs(7031) <= not(inputs(49)) or (inputs(112));
    layer0_outputs(7032) <= (inputs(79)) and not (inputs(174));
    layer0_outputs(7033) <= not(inputs(232));
    layer0_outputs(7034) <= inputs(183);
    layer0_outputs(7035) <= inputs(90);
    layer0_outputs(7036) <= not((inputs(234)) and (inputs(198)));
    layer0_outputs(7037) <= inputs(100);
    layer0_outputs(7038) <= inputs(57);
    layer0_outputs(7039) <= not(inputs(131));
    layer0_outputs(7040) <= not((inputs(157)) or (inputs(172)));
    layer0_outputs(7041) <= not(inputs(137));
    layer0_outputs(7042) <= not(inputs(220)) or (inputs(81));
    layer0_outputs(7043) <= not((inputs(162)) or (inputs(188)));
    layer0_outputs(7044) <= not(inputs(13)) or (inputs(220));
    layer0_outputs(7045) <= inputs(143);
    layer0_outputs(7046) <= not(inputs(133)) or (inputs(203));
    layer0_outputs(7047) <= not((inputs(111)) xor (inputs(115)));
    layer0_outputs(7048) <= inputs(28);
    layer0_outputs(7049) <= '0';
    layer0_outputs(7050) <= inputs(119);
    layer0_outputs(7051) <= not(inputs(112));
    layer0_outputs(7052) <= '0';
    layer0_outputs(7053) <= not(inputs(205)) or (inputs(144));
    layer0_outputs(7054) <= (inputs(203)) and not (inputs(43));
    layer0_outputs(7055) <= '0';
    layer0_outputs(7056) <= not((inputs(98)) or (inputs(7)));
    layer0_outputs(7057) <= not(inputs(247));
    layer0_outputs(7058) <= (inputs(169)) or (inputs(238));
    layer0_outputs(7059) <= inputs(136);
    layer0_outputs(7060) <= not(inputs(2));
    layer0_outputs(7061) <= not((inputs(232)) or (inputs(174)));
    layer0_outputs(7062) <= not(inputs(228));
    layer0_outputs(7063) <= (inputs(92)) xor (inputs(127));
    layer0_outputs(7064) <= not(inputs(129));
    layer0_outputs(7065) <= not(inputs(132));
    layer0_outputs(7066) <= not((inputs(207)) or (inputs(136)));
    layer0_outputs(7067) <= not(inputs(91));
    layer0_outputs(7068) <= not(inputs(2));
    layer0_outputs(7069) <= not((inputs(17)) and (inputs(111)));
    layer0_outputs(7070) <= not((inputs(32)) or (inputs(35)));
    layer0_outputs(7071) <= (inputs(214)) or (inputs(230));
    layer0_outputs(7072) <= not((inputs(123)) and (inputs(138)));
    layer0_outputs(7073) <= '0';
    layer0_outputs(7074) <= (inputs(141)) xor (inputs(189));
    layer0_outputs(7075) <= (inputs(231)) and not (inputs(69));
    layer0_outputs(7076) <= '1';
    layer0_outputs(7077) <= not((inputs(88)) or (inputs(225)));
    layer0_outputs(7078) <= (inputs(66)) xor (inputs(53));
    layer0_outputs(7079) <= not((inputs(92)) and (inputs(72)));
    layer0_outputs(7080) <= (inputs(142)) and not (inputs(26));
    layer0_outputs(7081) <= inputs(145);
    layer0_outputs(7082) <= not(inputs(66)) or (inputs(30));
    layer0_outputs(7083) <= (inputs(109)) and not (inputs(160));
    layer0_outputs(7084) <= not(inputs(117));
    layer0_outputs(7085) <= (inputs(229)) or (inputs(102));
    layer0_outputs(7086) <= not((inputs(229)) xor (inputs(214)));
    layer0_outputs(7087) <= not((inputs(36)) or (inputs(236)));
    layer0_outputs(7088) <= not((inputs(41)) and (inputs(73)));
    layer0_outputs(7089) <= inputs(120);
    layer0_outputs(7090) <= not((inputs(169)) or (inputs(47)));
    layer0_outputs(7091) <= (inputs(61)) xor (inputs(202));
    layer0_outputs(7092) <= '0';
    layer0_outputs(7093) <= inputs(86);
    layer0_outputs(7094) <= not(inputs(106));
    layer0_outputs(7095) <= inputs(150);
    layer0_outputs(7096) <= not(inputs(212)) or (inputs(97));
    layer0_outputs(7097) <= '1';
    layer0_outputs(7098) <= '1';
    layer0_outputs(7099) <= inputs(42);
    layer0_outputs(7100) <= inputs(183);
    layer0_outputs(7101) <= not(inputs(189));
    layer0_outputs(7102) <= not(inputs(255));
    layer0_outputs(7103) <= not(inputs(83)) or (inputs(181));
    layer0_outputs(7104) <= not((inputs(66)) xor (inputs(115)));
    layer0_outputs(7105) <= (inputs(35)) and not (inputs(70));
    layer0_outputs(7106) <= (inputs(225)) and (inputs(100));
    layer0_outputs(7107) <= not((inputs(152)) or (inputs(238)));
    layer0_outputs(7108) <= not(inputs(22)) or (inputs(86));
    layer0_outputs(7109) <= (inputs(229)) or (inputs(7));
    layer0_outputs(7110) <= not((inputs(36)) or (inputs(38)));
    layer0_outputs(7111) <= '1';
    layer0_outputs(7112) <= not(inputs(226)) or (inputs(58));
    layer0_outputs(7113) <= not((inputs(222)) xor (inputs(36)));
    layer0_outputs(7114) <= not(inputs(98)) or (inputs(224));
    layer0_outputs(7115) <= not(inputs(89)) or (inputs(221));
    layer0_outputs(7116) <= inputs(249);
    layer0_outputs(7117) <= (inputs(203)) and not (inputs(223));
    layer0_outputs(7118) <= not((inputs(51)) or (inputs(81)));
    layer0_outputs(7119) <= not(inputs(100)) or (inputs(143));
    layer0_outputs(7120) <= not(inputs(2));
    layer0_outputs(7121) <= not((inputs(83)) or (inputs(188)));
    layer0_outputs(7122) <= not((inputs(242)) and (inputs(236)));
    layer0_outputs(7123) <= not(inputs(69)) or (inputs(20));
    layer0_outputs(7124) <= not(inputs(247)) or (inputs(33));
    layer0_outputs(7125) <= (inputs(224)) or (inputs(202));
    layer0_outputs(7126) <= not(inputs(119));
    layer0_outputs(7127) <= (inputs(222)) or (inputs(55));
    layer0_outputs(7128) <= (inputs(200)) or (inputs(164));
    layer0_outputs(7129) <= not(inputs(99));
    layer0_outputs(7130) <= not(inputs(87));
    layer0_outputs(7131) <= not((inputs(11)) or (inputs(5)));
    layer0_outputs(7132) <= (inputs(224)) and not (inputs(63));
    layer0_outputs(7133) <= not((inputs(200)) or (inputs(253)));
    layer0_outputs(7134) <= not(inputs(114));
    layer0_outputs(7135) <= not(inputs(132));
    layer0_outputs(7136) <= not((inputs(211)) xor (inputs(249)));
    layer0_outputs(7137) <= inputs(40);
    layer0_outputs(7138) <= inputs(77);
    layer0_outputs(7139) <= (inputs(17)) xor (inputs(84));
    layer0_outputs(7140) <= not((inputs(7)) or (inputs(176)));
    layer0_outputs(7141) <= (inputs(226)) and (inputs(62));
    layer0_outputs(7142) <= (inputs(140)) and not (inputs(243));
    layer0_outputs(7143) <= (inputs(241)) and (inputs(238));
    layer0_outputs(7144) <= not(inputs(142)) or (inputs(255));
    layer0_outputs(7145) <= not(inputs(219));
    layer0_outputs(7146) <= '1';
    layer0_outputs(7147) <= (inputs(168)) or (inputs(191));
    layer0_outputs(7148) <= not(inputs(128));
    layer0_outputs(7149) <= (inputs(170)) or (inputs(97));
    layer0_outputs(7150) <= not((inputs(252)) or (inputs(87)));
    layer0_outputs(7151) <= '0';
    layer0_outputs(7152) <= inputs(40);
    layer0_outputs(7153) <= inputs(188);
    layer0_outputs(7154) <= (inputs(13)) and not (inputs(166));
    layer0_outputs(7155) <= '1';
    layer0_outputs(7156) <= (inputs(177)) or (inputs(181));
    layer0_outputs(7157) <= not(inputs(182));
    layer0_outputs(7158) <= not(inputs(172));
    layer0_outputs(7159) <= (inputs(15)) or (inputs(131));
    layer0_outputs(7160) <= not(inputs(167));
    layer0_outputs(7161) <= not(inputs(89));
    layer0_outputs(7162) <= not((inputs(233)) xor (inputs(159)));
    layer0_outputs(7163) <= not((inputs(91)) or (inputs(143)));
    layer0_outputs(7164) <= (inputs(135)) or (inputs(232));
    layer0_outputs(7165) <= (inputs(136)) and (inputs(113));
    layer0_outputs(7166) <= not((inputs(159)) and (inputs(215)));
    layer0_outputs(7167) <= not((inputs(223)) or (inputs(98)));
    layer0_outputs(7168) <= (inputs(51)) or (inputs(127));
    layer0_outputs(7169) <= (inputs(135)) and not (inputs(224));
    layer0_outputs(7170) <= (inputs(60)) or (inputs(210));
    layer0_outputs(7171) <= inputs(237);
    layer0_outputs(7172) <= not((inputs(1)) or (inputs(65)));
    layer0_outputs(7173) <= (inputs(255)) or (inputs(198));
    layer0_outputs(7174) <= (inputs(69)) or (inputs(36));
    layer0_outputs(7175) <= not(inputs(92));
    layer0_outputs(7176) <= not(inputs(90));
    layer0_outputs(7177) <= not(inputs(251)) or (inputs(64));
    layer0_outputs(7178) <= not(inputs(233));
    layer0_outputs(7179) <= (inputs(249)) or (inputs(196));
    layer0_outputs(7180) <= not(inputs(170));
    layer0_outputs(7181) <= (inputs(206)) or (inputs(4));
    layer0_outputs(7182) <= not((inputs(16)) and (inputs(182)));
    layer0_outputs(7183) <= not(inputs(225)) or (inputs(220));
    layer0_outputs(7184) <= not(inputs(12));
    layer0_outputs(7185) <= (inputs(12)) and (inputs(90));
    layer0_outputs(7186) <= not((inputs(76)) or (inputs(201)));
    layer0_outputs(7187) <= (inputs(190)) or (inputs(171));
    layer0_outputs(7188) <= (inputs(129)) or (inputs(211));
    layer0_outputs(7189) <= not(inputs(221));
    layer0_outputs(7190) <= (inputs(25)) and (inputs(27));
    layer0_outputs(7191) <= not(inputs(198)) or (inputs(90));
    layer0_outputs(7192) <= not((inputs(118)) or (inputs(116)));
    layer0_outputs(7193) <= inputs(37);
    layer0_outputs(7194) <= not(inputs(33));
    layer0_outputs(7195) <= (inputs(103)) and not (inputs(47));
    layer0_outputs(7196) <= inputs(177);
    layer0_outputs(7197) <= not(inputs(175)) or (inputs(12));
    layer0_outputs(7198) <= not((inputs(186)) and (inputs(42)));
    layer0_outputs(7199) <= not(inputs(173)) or (inputs(224));
    layer0_outputs(7200) <= (inputs(7)) xor (inputs(77));
    layer0_outputs(7201) <= not(inputs(91));
    layer0_outputs(7202) <= not(inputs(11)) or (inputs(231));
    layer0_outputs(7203) <= '0';
    layer0_outputs(7204) <= (inputs(207)) and (inputs(149));
    layer0_outputs(7205) <= not(inputs(61)) or (inputs(227));
    layer0_outputs(7206) <= '0';
    layer0_outputs(7207) <= '1';
    layer0_outputs(7208) <= (inputs(19)) xor (inputs(52));
    layer0_outputs(7209) <= '1';
    layer0_outputs(7210) <= not(inputs(227)) or (inputs(124));
    layer0_outputs(7211) <= (inputs(203)) xor (inputs(21));
    layer0_outputs(7212) <= not(inputs(81)) or (inputs(176));
    layer0_outputs(7213) <= (inputs(117)) and not (inputs(97));
    layer0_outputs(7214) <= not(inputs(213));
    layer0_outputs(7215) <= not(inputs(84)) or (inputs(33));
    layer0_outputs(7216) <= not(inputs(229)) or (inputs(58));
    layer0_outputs(7217) <= not((inputs(70)) or (inputs(68)));
    layer0_outputs(7218) <= not(inputs(149)) or (inputs(236));
    layer0_outputs(7219) <= '1';
    layer0_outputs(7220) <= (inputs(50)) xor (inputs(4));
    layer0_outputs(7221) <= (inputs(1)) and not (inputs(75));
    layer0_outputs(7222) <= (inputs(136)) and (inputs(74));
    layer0_outputs(7223) <= (inputs(7)) and not (inputs(216));
    layer0_outputs(7224) <= (inputs(166)) and not (inputs(159));
    layer0_outputs(7225) <= (inputs(189)) xor (inputs(102));
    layer0_outputs(7226) <= inputs(116);
    layer0_outputs(7227) <= (inputs(52)) and not (inputs(221));
    layer0_outputs(7228) <= inputs(55);
    layer0_outputs(7229) <= (inputs(178)) and not (inputs(32));
    layer0_outputs(7230) <= not((inputs(173)) and (inputs(72)));
    layer0_outputs(7231) <= (inputs(147)) and not (inputs(2));
    layer0_outputs(7232) <= '1';
    layer0_outputs(7233) <= (inputs(9)) and not (inputs(192));
    layer0_outputs(7234) <= (inputs(242)) and not (inputs(247));
    layer0_outputs(7235) <= (inputs(123)) or (inputs(186));
    layer0_outputs(7236) <= inputs(210);
    layer0_outputs(7237) <= (inputs(26)) or (inputs(112));
    layer0_outputs(7238) <= inputs(25);
    layer0_outputs(7239) <= inputs(161);
    layer0_outputs(7240) <= '0';
    layer0_outputs(7241) <= inputs(5);
    layer0_outputs(7242) <= not(inputs(99));
    layer0_outputs(7243) <= not(inputs(101));
    layer0_outputs(7244) <= (inputs(107)) and (inputs(33));
    layer0_outputs(7245) <= (inputs(67)) and not (inputs(0));
    layer0_outputs(7246) <= inputs(246);
    layer0_outputs(7247) <= not(inputs(104));
    layer0_outputs(7248) <= not(inputs(185)) or (inputs(6));
    layer0_outputs(7249) <= not(inputs(143));
    layer0_outputs(7250) <= (inputs(60)) xor (inputs(30));
    layer0_outputs(7251) <= not(inputs(254));
    layer0_outputs(7252) <= (inputs(233)) and not (inputs(207));
    layer0_outputs(7253) <= '0';
    layer0_outputs(7254) <= (inputs(181)) or (inputs(173));
    layer0_outputs(7255) <= (inputs(207)) and not (inputs(217));
    layer0_outputs(7256) <= inputs(190);
    layer0_outputs(7257) <= not(inputs(118));
    layer0_outputs(7258) <= not((inputs(137)) or (inputs(52)));
    layer0_outputs(7259) <= (inputs(52)) or (inputs(194));
    layer0_outputs(7260) <= (inputs(115)) or (inputs(161));
    layer0_outputs(7261) <= inputs(206);
    layer0_outputs(7262) <= inputs(228);
    layer0_outputs(7263) <= (inputs(11)) or (inputs(21));
    layer0_outputs(7264) <= not(inputs(35));
    layer0_outputs(7265) <= (inputs(109)) or (inputs(33));
    layer0_outputs(7266) <= not(inputs(8)) or (inputs(113));
    layer0_outputs(7267) <= (inputs(233)) and not (inputs(159));
    layer0_outputs(7268) <= (inputs(19)) and not (inputs(224));
    layer0_outputs(7269) <= not(inputs(119)) or (inputs(216));
    layer0_outputs(7270) <= (inputs(185)) and (inputs(28));
    layer0_outputs(7271) <= not((inputs(128)) or (inputs(82)));
    layer0_outputs(7272) <= (inputs(255)) and not (inputs(63));
    layer0_outputs(7273) <= '0';
    layer0_outputs(7274) <= (inputs(132)) and not (inputs(242));
    layer0_outputs(7275) <= (inputs(13)) and not (inputs(153));
    layer0_outputs(7276) <= not(inputs(201));
    layer0_outputs(7277) <= (inputs(160)) or (inputs(245));
    layer0_outputs(7278) <= (inputs(114)) and not (inputs(159));
    layer0_outputs(7279) <= not(inputs(243)) or (inputs(22));
    layer0_outputs(7280) <= '1';
    layer0_outputs(7281) <= not((inputs(153)) or (inputs(119)));
    layer0_outputs(7282) <= not((inputs(131)) or (inputs(141)));
    layer0_outputs(7283) <= not((inputs(207)) or (inputs(164)));
    layer0_outputs(7284) <= not(inputs(12)) or (inputs(140));
    layer0_outputs(7285) <= (inputs(52)) or (inputs(130));
    layer0_outputs(7286) <= (inputs(215)) xor (inputs(246));
    layer0_outputs(7287) <= not(inputs(38));
    layer0_outputs(7288) <= not(inputs(247));
    layer0_outputs(7289) <= (inputs(83)) and not (inputs(55));
    layer0_outputs(7290) <= inputs(88);
    layer0_outputs(7291) <= inputs(189);
    layer0_outputs(7292) <= not(inputs(83));
    layer0_outputs(7293) <= not((inputs(111)) and (inputs(54)));
    layer0_outputs(7294) <= not((inputs(192)) and (inputs(48)));
    layer0_outputs(7295) <= inputs(196);
    layer0_outputs(7296) <= not(inputs(113));
    layer0_outputs(7297) <= (inputs(208)) or (inputs(15));
    layer0_outputs(7298) <= inputs(93);
    layer0_outputs(7299) <= not(inputs(214));
    layer0_outputs(7300) <= (inputs(233)) or (inputs(188));
    layer0_outputs(7301) <= (inputs(26)) and not (inputs(175));
    layer0_outputs(7302) <= (inputs(53)) xor (inputs(24));
    layer0_outputs(7303) <= (inputs(26)) and not (inputs(249));
    layer0_outputs(7304) <= not(inputs(234)) or (inputs(81));
    layer0_outputs(7305) <= '1';
    layer0_outputs(7306) <= not(inputs(217));
    layer0_outputs(7307) <= not((inputs(193)) and (inputs(0)));
    layer0_outputs(7308) <= not((inputs(49)) and (inputs(52)));
    layer0_outputs(7309) <= (inputs(151)) and not (inputs(240));
    layer0_outputs(7310) <= (inputs(188)) and not (inputs(62));
    layer0_outputs(7311) <= '1';
    layer0_outputs(7312) <= not(inputs(20));
    layer0_outputs(7313) <= not((inputs(31)) and (inputs(121)));
    layer0_outputs(7314) <= (inputs(71)) xor (inputs(105));
    layer0_outputs(7315) <= inputs(212);
    layer0_outputs(7316) <= (inputs(232)) and not (inputs(253));
    layer0_outputs(7317) <= not(inputs(75));
    layer0_outputs(7318) <= (inputs(241)) and not (inputs(115));
    layer0_outputs(7319) <= inputs(60);
    layer0_outputs(7320) <= not(inputs(21));
    layer0_outputs(7321) <= not(inputs(147));
    layer0_outputs(7322) <= (inputs(134)) and (inputs(186));
    layer0_outputs(7323) <= (inputs(70)) xor (inputs(99));
    layer0_outputs(7324) <= (inputs(228)) and not (inputs(1));
    layer0_outputs(7325) <= inputs(179);
    layer0_outputs(7326) <= not(inputs(166)) or (inputs(157));
    layer0_outputs(7327) <= inputs(53);
    layer0_outputs(7328) <= inputs(238);
    layer0_outputs(7329) <= (inputs(125)) or (inputs(247));
    layer0_outputs(7330) <= '1';
    layer0_outputs(7331) <= (inputs(242)) xor (inputs(36));
    layer0_outputs(7332) <= inputs(133);
    layer0_outputs(7333) <= '1';
    layer0_outputs(7334) <= not((inputs(237)) or (inputs(167)));
    layer0_outputs(7335) <= not((inputs(199)) or (inputs(73)));
    layer0_outputs(7336) <= not(inputs(72));
    layer0_outputs(7337) <= not(inputs(173)) or (inputs(224));
    layer0_outputs(7338) <= not(inputs(209)) or (inputs(170));
    layer0_outputs(7339) <= not((inputs(164)) or (inputs(111)));
    layer0_outputs(7340) <= (inputs(125)) or (inputs(31));
    layer0_outputs(7341) <= inputs(160);
    layer0_outputs(7342) <= not(inputs(229)) or (inputs(239));
    layer0_outputs(7343) <= not(inputs(199));
    layer0_outputs(7344) <= not((inputs(3)) or (inputs(54)));
    layer0_outputs(7345) <= not((inputs(137)) and (inputs(42)));
    layer0_outputs(7346) <= not(inputs(195)) or (inputs(46));
    layer0_outputs(7347) <= not(inputs(207));
    layer0_outputs(7348) <= inputs(247);
    layer0_outputs(7349) <= not((inputs(56)) xor (inputs(119)));
    layer0_outputs(7350) <= inputs(163);
    layer0_outputs(7351) <= inputs(128);
    layer0_outputs(7352) <= '0';
    layer0_outputs(7353) <= '0';
    layer0_outputs(7354) <= inputs(183);
    layer0_outputs(7355) <= inputs(82);
    layer0_outputs(7356) <= not(inputs(230));
    layer0_outputs(7357) <= not(inputs(82));
    layer0_outputs(7358) <= not(inputs(149)) or (inputs(228));
    layer0_outputs(7359) <= inputs(204);
    layer0_outputs(7360) <= not(inputs(70));
    layer0_outputs(7361) <= (inputs(88)) and (inputs(67));
    layer0_outputs(7362) <= (inputs(45)) or (inputs(166));
    layer0_outputs(7363) <= (inputs(180)) and not (inputs(34));
    layer0_outputs(7364) <= not(inputs(195)) or (inputs(125));
    layer0_outputs(7365) <= inputs(130);
    layer0_outputs(7366) <= (inputs(70)) and not (inputs(60));
    layer0_outputs(7367) <= inputs(91);
    layer0_outputs(7368) <= (inputs(168)) or (inputs(151));
    layer0_outputs(7369) <= not(inputs(179));
    layer0_outputs(7370) <= (inputs(173)) or (inputs(158));
    layer0_outputs(7371) <= not(inputs(12));
    layer0_outputs(7372) <= not(inputs(80)) or (inputs(255));
    layer0_outputs(7373) <= not(inputs(150)) or (inputs(58));
    layer0_outputs(7374) <= (inputs(126)) or (inputs(20));
    layer0_outputs(7375) <= not(inputs(37));
    layer0_outputs(7376) <= not(inputs(175));
    layer0_outputs(7377) <= '1';
    layer0_outputs(7378) <= (inputs(131)) and (inputs(155));
    layer0_outputs(7379) <= not(inputs(27));
    layer0_outputs(7380) <= (inputs(240)) or (inputs(28));
    layer0_outputs(7381) <= (inputs(243)) or (inputs(115));
    layer0_outputs(7382) <= not(inputs(145));
    layer0_outputs(7383) <= (inputs(66)) and not (inputs(106));
    layer0_outputs(7384) <= not(inputs(182));
    layer0_outputs(7385) <= (inputs(80)) and not (inputs(111));
    layer0_outputs(7386) <= (inputs(15)) and not (inputs(236));
    layer0_outputs(7387) <= not(inputs(38)) or (inputs(128));
    layer0_outputs(7388) <= not(inputs(16));
    layer0_outputs(7389) <= (inputs(104)) or (inputs(161));
    layer0_outputs(7390) <= inputs(95);
    layer0_outputs(7391) <= (inputs(151)) or (inputs(32));
    layer0_outputs(7392) <= not((inputs(187)) and (inputs(180)));
    layer0_outputs(7393) <= not(inputs(119));
    layer0_outputs(7394) <= inputs(55);
    layer0_outputs(7395) <= (inputs(153)) and (inputs(84));
    layer0_outputs(7396) <= (inputs(109)) xor (inputs(142));
    layer0_outputs(7397) <= (inputs(165)) or (inputs(126));
    layer0_outputs(7398) <= '0';
    layer0_outputs(7399) <= '1';
    layer0_outputs(7400) <= inputs(84);
    layer0_outputs(7401) <= not((inputs(156)) or (inputs(75)));
    layer0_outputs(7402) <= not((inputs(110)) or (inputs(222)));
    layer0_outputs(7403) <= inputs(248);
    layer0_outputs(7404) <= (inputs(173)) or (inputs(196));
    layer0_outputs(7405) <= not((inputs(99)) or (inputs(56)));
    layer0_outputs(7406) <= not(inputs(186)) or (inputs(76));
    layer0_outputs(7407) <= (inputs(178)) xor (inputs(89));
    layer0_outputs(7408) <= (inputs(172)) or (inputs(219));
    layer0_outputs(7409) <= not(inputs(24)) or (inputs(208));
    layer0_outputs(7410) <= inputs(142);
    layer0_outputs(7411) <= not(inputs(225)) or (inputs(112));
    layer0_outputs(7412) <= not(inputs(70));
    layer0_outputs(7413) <= inputs(171);
    layer0_outputs(7414) <= not((inputs(238)) or (inputs(254)));
    layer0_outputs(7415) <= inputs(226);
    layer0_outputs(7416) <= (inputs(153)) and not (inputs(211));
    layer0_outputs(7417) <= not(inputs(233));
    layer0_outputs(7418) <= (inputs(201)) and (inputs(173));
    layer0_outputs(7419) <= (inputs(168)) and not (inputs(6));
    layer0_outputs(7420) <= (inputs(235)) and not (inputs(142));
    layer0_outputs(7421) <= '0';
    layer0_outputs(7422) <= not(inputs(120)) or (inputs(17));
    layer0_outputs(7423) <= not((inputs(238)) or (inputs(163)));
    layer0_outputs(7424) <= '0';
    layer0_outputs(7425) <= inputs(160);
    layer0_outputs(7426) <= '0';
    layer0_outputs(7427) <= not((inputs(238)) xor (inputs(176)));
    layer0_outputs(7428) <= (inputs(189)) or (inputs(206));
    layer0_outputs(7429) <= not(inputs(57)) or (inputs(15));
    layer0_outputs(7430) <= '0';
    layer0_outputs(7431) <= not(inputs(167)) or (inputs(247));
    layer0_outputs(7432) <= '0';
    layer0_outputs(7433) <= inputs(47);
    layer0_outputs(7434) <= not((inputs(39)) or (inputs(242)));
    layer0_outputs(7435) <= (inputs(187)) and not (inputs(165));
    layer0_outputs(7436) <= (inputs(126)) and not (inputs(195));
    layer0_outputs(7437) <= (inputs(232)) and not (inputs(31));
    layer0_outputs(7438) <= (inputs(80)) and not (inputs(146));
    layer0_outputs(7439) <= not(inputs(13));
    layer0_outputs(7440) <= not(inputs(229)) or (inputs(191));
    layer0_outputs(7441) <= not(inputs(100));
    layer0_outputs(7442) <= (inputs(8)) and (inputs(13));
    layer0_outputs(7443) <= not(inputs(203));
    layer0_outputs(7444) <= not(inputs(254));
    layer0_outputs(7445) <= (inputs(50)) xor (inputs(20));
    layer0_outputs(7446) <= inputs(91);
    layer0_outputs(7447) <= (inputs(19)) and not (inputs(200));
    layer0_outputs(7448) <= inputs(99);
    layer0_outputs(7449) <= (inputs(156)) and (inputs(49));
    layer0_outputs(7450) <= not(inputs(6));
    layer0_outputs(7451) <= inputs(165);
    layer0_outputs(7452) <= not((inputs(31)) and (inputs(125)));
    layer0_outputs(7453) <= not((inputs(15)) or (inputs(130)));
    layer0_outputs(7454) <= not(inputs(142)) or (inputs(5));
    layer0_outputs(7455) <= not((inputs(192)) or (inputs(68)));
    layer0_outputs(7456) <= (inputs(82)) xor (inputs(98));
    layer0_outputs(7457) <= not((inputs(203)) or (inputs(244)));
    layer0_outputs(7458) <= '1';
    layer0_outputs(7459) <= inputs(230);
    layer0_outputs(7460) <= not(inputs(198)) or (inputs(17));
    layer0_outputs(7461) <= inputs(179);
    layer0_outputs(7462) <= not((inputs(141)) xor (inputs(190)));
    layer0_outputs(7463) <= not(inputs(193)) or (inputs(136));
    layer0_outputs(7464) <= not(inputs(71));
    layer0_outputs(7465) <= inputs(200);
    layer0_outputs(7466) <= not(inputs(16)) or (inputs(139));
    layer0_outputs(7467) <= inputs(195);
    layer0_outputs(7468) <= '0';
    layer0_outputs(7469) <= not(inputs(13));
    layer0_outputs(7470) <= (inputs(199)) and not (inputs(156));
    layer0_outputs(7471) <= (inputs(167)) or (inputs(215));
    layer0_outputs(7472) <= '0';
    layer0_outputs(7473) <= not(inputs(206)) or (inputs(175));
    layer0_outputs(7474) <= (inputs(11)) and (inputs(80));
    layer0_outputs(7475) <= not((inputs(226)) and (inputs(0)));
    layer0_outputs(7476) <= '1';
    layer0_outputs(7477) <= not(inputs(138));
    layer0_outputs(7478) <= not(inputs(52));
    layer0_outputs(7479) <= not((inputs(141)) or (inputs(241)));
    layer0_outputs(7480) <= (inputs(207)) and (inputs(49));
    layer0_outputs(7481) <= (inputs(251)) and (inputs(1));
    layer0_outputs(7482) <= (inputs(178)) or (inputs(39));
    layer0_outputs(7483) <= not(inputs(19));
    layer0_outputs(7484) <= not((inputs(22)) xor (inputs(158)));
    layer0_outputs(7485) <= inputs(157);
    layer0_outputs(7486) <= (inputs(168)) and not (inputs(128));
    layer0_outputs(7487) <= not(inputs(159));
    layer0_outputs(7488) <= '0';
    layer0_outputs(7489) <= (inputs(111)) or (inputs(209));
    layer0_outputs(7490) <= (inputs(216)) and (inputs(228));
    layer0_outputs(7491) <= not((inputs(156)) or (inputs(212)));
    layer0_outputs(7492) <= (inputs(243)) and not (inputs(23));
    layer0_outputs(7493) <= not(inputs(208));
    layer0_outputs(7494) <= (inputs(148)) or (inputs(207));
    layer0_outputs(7495) <= not((inputs(65)) or (inputs(9)));
    layer0_outputs(7496) <= not(inputs(196));
    layer0_outputs(7497) <= inputs(194);
    layer0_outputs(7498) <= (inputs(34)) and not (inputs(87));
    layer0_outputs(7499) <= not((inputs(252)) xor (inputs(207)));
    layer0_outputs(7500) <= inputs(104);
    layer0_outputs(7501) <= '0';
    layer0_outputs(7502) <= inputs(58);
    layer0_outputs(7503) <= '0';
    layer0_outputs(7504) <= not(inputs(48));
    layer0_outputs(7505) <= (inputs(132)) and not (inputs(153));
    layer0_outputs(7506) <= '1';
    layer0_outputs(7507) <= (inputs(98)) or (inputs(161));
    layer0_outputs(7508) <= (inputs(76)) and not (inputs(11));
    layer0_outputs(7509) <= not((inputs(140)) and (inputs(127)));
    layer0_outputs(7510) <= '1';
    layer0_outputs(7511) <= not(inputs(170));
    layer0_outputs(7512) <= inputs(137);
    layer0_outputs(7513) <= not(inputs(23));
    layer0_outputs(7514) <= (inputs(31)) and (inputs(161));
    layer0_outputs(7515) <= '0';
    layer0_outputs(7516) <= inputs(249);
    layer0_outputs(7517) <= (inputs(223)) and not (inputs(63));
    layer0_outputs(7518) <= not(inputs(236));
    layer0_outputs(7519) <= not(inputs(72));
    layer0_outputs(7520) <= inputs(84);
    layer0_outputs(7521) <= inputs(59);
    layer0_outputs(7522) <= not(inputs(103)) or (inputs(165));
    layer0_outputs(7523) <= (inputs(167)) or (inputs(166));
    layer0_outputs(7524) <= (inputs(228)) or (inputs(210));
    layer0_outputs(7525) <= not(inputs(164));
    layer0_outputs(7526) <= not(inputs(74)) or (inputs(141));
    layer0_outputs(7527) <= (inputs(189)) or (inputs(163));
    layer0_outputs(7528) <= not(inputs(231));
    layer0_outputs(7529) <= (inputs(194)) and not (inputs(75));
    layer0_outputs(7530) <= not(inputs(172)) or (inputs(215));
    layer0_outputs(7531) <= not((inputs(211)) or (inputs(64)));
    layer0_outputs(7532) <= not((inputs(82)) xor (inputs(68)));
    layer0_outputs(7533) <= not(inputs(51));
    layer0_outputs(7534) <= inputs(220);
    layer0_outputs(7535) <= (inputs(212)) and not (inputs(237));
    layer0_outputs(7536) <= inputs(154);
    layer0_outputs(7537) <= (inputs(126)) xor (inputs(163));
    layer0_outputs(7538) <= not((inputs(71)) xor (inputs(120)));
    layer0_outputs(7539) <= inputs(2);
    layer0_outputs(7540) <= not(inputs(225));
    layer0_outputs(7541) <= inputs(102);
    layer0_outputs(7542) <= (inputs(56)) and (inputs(73));
    layer0_outputs(7543) <= inputs(187);
    layer0_outputs(7544) <= not(inputs(206));
    layer0_outputs(7545) <= inputs(200);
    layer0_outputs(7546) <= inputs(42);
    layer0_outputs(7547) <= inputs(114);
    layer0_outputs(7548) <= not(inputs(82));
    layer0_outputs(7549) <= inputs(7);
    layer0_outputs(7550) <= not((inputs(252)) or (inputs(191)));
    layer0_outputs(7551) <= (inputs(9)) and (inputs(102));
    layer0_outputs(7552) <= inputs(229);
    layer0_outputs(7553) <= (inputs(148)) and not (inputs(11));
    layer0_outputs(7554) <= inputs(230);
    layer0_outputs(7555) <= (inputs(182)) and not (inputs(217));
    layer0_outputs(7556) <= (inputs(170)) or (inputs(152));
    layer0_outputs(7557) <= not(inputs(105));
    layer0_outputs(7558) <= not(inputs(241)) or (inputs(46));
    layer0_outputs(7559) <= not(inputs(26)) or (inputs(208));
    layer0_outputs(7560) <= (inputs(78)) or (inputs(190));
    layer0_outputs(7561) <= not(inputs(100)) or (inputs(224));
    layer0_outputs(7562) <= not((inputs(185)) and (inputs(249)));
    layer0_outputs(7563) <= inputs(24);
    layer0_outputs(7564) <= (inputs(227)) xor (inputs(53));
    layer0_outputs(7565) <= not((inputs(81)) and (inputs(145)));
    layer0_outputs(7566) <= not((inputs(70)) or (inputs(243)));
    layer0_outputs(7567) <= '0';
    layer0_outputs(7568) <= (inputs(34)) xor (inputs(62));
    layer0_outputs(7569) <= '0';
    layer0_outputs(7570) <= (inputs(98)) or (inputs(96));
    layer0_outputs(7571) <= '1';
    layer0_outputs(7572) <= inputs(104);
    layer0_outputs(7573) <= inputs(190);
    layer0_outputs(7574) <= (inputs(59)) and not (inputs(126));
    layer0_outputs(7575) <= not(inputs(22));
    layer0_outputs(7576) <= inputs(171);
    layer0_outputs(7577) <= (inputs(174)) or (inputs(28));
    layer0_outputs(7578) <= inputs(0);
    layer0_outputs(7579) <= (inputs(34)) xor (inputs(135));
    layer0_outputs(7580) <= not(inputs(97));
    layer0_outputs(7581) <= (inputs(54)) and not (inputs(218));
    layer0_outputs(7582) <= (inputs(53)) and (inputs(207));
    layer0_outputs(7583) <= not(inputs(77));
    layer0_outputs(7584) <= inputs(64);
    layer0_outputs(7585) <= inputs(74);
    layer0_outputs(7586) <= not((inputs(118)) or (inputs(241)));
    layer0_outputs(7587) <= (inputs(63)) and not (inputs(207));
    layer0_outputs(7588) <= not((inputs(58)) xor (inputs(46)));
    layer0_outputs(7589) <= inputs(115);
    layer0_outputs(7590) <= (inputs(108)) and not (inputs(4));
    layer0_outputs(7591) <= '1';
    layer0_outputs(7592) <= not(inputs(34));
    layer0_outputs(7593) <= not((inputs(76)) xor (inputs(195)));
    layer0_outputs(7594) <= not((inputs(33)) and (inputs(220)));
    layer0_outputs(7595) <= not(inputs(194));
    layer0_outputs(7596) <= not(inputs(232));
    layer0_outputs(7597) <= inputs(238);
    layer0_outputs(7598) <= '1';
    layer0_outputs(7599) <= (inputs(216)) or (inputs(159));
    layer0_outputs(7600) <= '0';
    layer0_outputs(7601) <= not((inputs(8)) or (inputs(203)));
    layer0_outputs(7602) <= not((inputs(94)) or (inputs(253)));
    layer0_outputs(7603) <= not((inputs(163)) or (inputs(223)));
    layer0_outputs(7604) <= inputs(103);
    layer0_outputs(7605) <= not(inputs(33));
    layer0_outputs(7606) <= (inputs(219)) and not (inputs(185));
    layer0_outputs(7607) <= (inputs(101)) and not (inputs(88));
    layer0_outputs(7608) <= not(inputs(241));
    layer0_outputs(7609) <= '1';
    layer0_outputs(7610) <= not(inputs(212));
    layer0_outputs(7611) <= not((inputs(65)) and (inputs(17)));
    layer0_outputs(7612) <= inputs(86);
    layer0_outputs(7613) <= not(inputs(128));
    layer0_outputs(7614) <= (inputs(211)) and not (inputs(104));
    layer0_outputs(7615) <= not(inputs(185));
    layer0_outputs(7616) <= not(inputs(8));
    layer0_outputs(7617) <= inputs(4);
    layer0_outputs(7618) <= (inputs(60)) xor (inputs(237));
    layer0_outputs(7619) <= '0';
    layer0_outputs(7620) <= inputs(16);
    layer0_outputs(7621) <= inputs(132);
    layer0_outputs(7622) <= not((inputs(201)) or (inputs(221)));
    layer0_outputs(7623) <= (inputs(25)) and not (inputs(157));
    layer0_outputs(7624) <= not((inputs(217)) or (inputs(232)));
    layer0_outputs(7625) <= (inputs(243)) or (inputs(192));
    layer0_outputs(7626) <= not(inputs(194)) or (inputs(146));
    layer0_outputs(7627) <= not(inputs(234)) or (inputs(85));
    layer0_outputs(7628) <= not(inputs(151)) or (inputs(14));
    layer0_outputs(7629) <= not(inputs(54));
    layer0_outputs(7630) <= (inputs(31)) and (inputs(68));
    layer0_outputs(7631) <= not((inputs(56)) and (inputs(46)));
    layer0_outputs(7632) <= not((inputs(189)) or (inputs(69)));
    layer0_outputs(7633) <= not((inputs(248)) xor (inputs(186)));
    layer0_outputs(7634) <= not((inputs(3)) or (inputs(34)));
    layer0_outputs(7635) <= not(inputs(86)) or (inputs(225));
    layer0_outputs(7636) <= inputs(21);
    layer0_outputs(7637) <= (inputs(212)) or (inputs(44));
    layer0_outputs(7638) <= inputs(113);
    layer0_outputs(7639) <= not((inputs(23)) or (inputs(22)));
    layer0_outputs(7640) <= not((inputs(43)) xor (inputs(40)));
    layer0_outputs(7641) <= '1';
    layer0_outputs(7642) <= (inputs(39)) and not (inputs(174));
    layer0_outputs(7643) <= (inputs(233)) and not (inputs(209));
    layer0_outputs(7644) <= '0';
    layer0_outputs(7645) <= not((inputs(145)) and (inputs(151)));
    layer0_outputs(7646) <= inputs(136);
    layer0_outputs(7647) <= not(inputs(202));
    layer0_outputs(7648) <= (inputs(81)) or (inputs(197));
    layer0_outputs(7649) <= inputs(27);
    layer0_outputs(7650) <= inputs(90);
    layer0_outputs(7651) <= inputs(18);
    layer0_outputs(7652) <= inputs(43);
    layer0_outputs(7653) <= not(inputs(151));
    layer0_outputs(7654) <= (inputs(234)) or (inputs(193));
    layer0_outputs(7655) <= (inputs(68)) or (inputs(209));
    layer0_outputs(7656) <= inputs(125);
    layer0_outputs(7657) <= not(inputs(71)) or (inputs(250));
    layer0_outputs(7658) <= not(inputs(77));
    layer0_outputs(7659) <= (inputs(142)) xor (inputs(190));
    layer0_outputs(7660) <= not(inputs(144)) or (inputs(243));
    layer0_outputs(7661) <= inputs(123);
    layer0_outputs(7662) <= inputs(228);
    layer0_outputs(7663) <= not(inputs(199)) or (inputs(129));
    layer0_outputs(7664) <= (inputs(48)) and not (inputs(9));
    layer0_outputs(7665) <= (inputs(237)) xor (inputs(161));
    layer0_outputs(7666) <= inputs(101);
    layer0_outputs(7667) <= '1';
    layer0_outputs(7668) <= not((inputs(205)) or (inputs(180)));
    layer0_outputs(7669) <= '0';
    layer0_outputs(7670) <= inputs(168);
    layer0_outputs(7671) <= (inputs(199)) and (inputs(156));
    layer0_outputs(7672) <= (inputs(1)) xor (inputs(136));
    layer0_outputs(7673) <= inputs(127);
    layer0_outputs(7674) <= not(inputs(155));
    layer0_outputs(7675) <= inputs(202);
    layer0_outputs(7676) <= not((inputs(224)) xor (inputs(31)));
    layer0_outputs(7677) <= (inputs(60)) and not (inputs(186));
    layer0_outputs(7678) <= not((inputs(50)) or (inputs(169)));
    layer0_outputs(7679) <= '0';
    layer1_outputs(0) <= '0';
    layer1_outputs(1) <= layer0_outputs(7247);
    layer1_outputs(2) <= (layer0_outputs(3254)) or (layer0_outputs(291));
    layer1_outputs(3) <= not((layer0_outputs(3170)) and (layer0_outputs(5887)));
    layer1_outputs(4) <= not(layer0_outputs(6607));
    layer1_outputs(5) <= layer0_outputs(81);
    layer1_outputs(6) <= (layer0_outputs(515)) and not (layer0_outputs(1546));
    layer1_outputs(7) <= '0';
    layer1_outputs(8) <= not(layer0_outputs(6508));
    layer1_outputs(9) <= not(layer0_outputs(2225));
    layer1_outputs(10) <= not((layer0_outputs(5429)) and (layer0_outputs(624)));
    layer1_outputs(11) <= (layer0_outputs(1601)) or (layer0_outputs(6657));
    layer1_outputs(12) <= layer0_outputs(4250);
    layer1_outputs(13) <= (layer0_outputs(662)) and (layer0_outputs(7507));
    layer1_outputs(14) <= (layer0_outputs(3881)) and (layer0_outputs(793));
    layer1_outputs(15) <= '0';
    layer1_outputs(16) <= (layer0_outputs(353)) and not (layer0_outputs(6237));
    layer1_outputs(17) <= '1';
    layer1_outputs(18) <= not(layer0_outputs(2764));
    layer1_outputs(19) <= not(layer0_outputs(629));
    layer1_outputs(20) <= not((layer0_outputs(2730)) and (layer0_outputs(937)));
    layer1_outputs(21) <= not(layer0_outputs(1724)) or (layer0_outputs(2760));
    layer1_outputs(22) <= not((layer0_outputs(712)) and (layer0_outputs(5569)));
    layer1_outputs(23) <= layer0_outputs(4350);
    layer1_outputs(24) <= not((layer0_outputs(4603)) and (layer0_outputs(3164)));
    layer1_outputs(25) <= not(layer0_outputs(2283));
    layer1_outputs(26) <= layer0_outputs(2657);
    layer1_outputs(27) <= not(layer0_outputs(2848)) or (layer0_outputs(6216));
    layer1_outputs(28) <= layer0_outputs(169);
    layer1_outputs(29) <= layer0_outputs(1827);
    layer1_outputs(30) <= (layer0_outputs(6394)) or (layer0_outputs(4005));
    layer1_outputs(31) <= not(layer0_outputs(2929)) or (layer0_outputs(3291));
    layer1_outputs(32) <= not((layer0_outputs(3736)) or (layer0_outputs(2655)));
    layer1_outputs(33) <= layer0_outputs(3626);
    layer1_outputs(34) <= not(layer0_outputs(6127));
    layer1_outputs(35) <= (layer0_outputs(5727)) and not (layer0_outputs(557));
    layer1_outputs(36) <= not(layer0_outputs(6413)) or (layer0_outputs(2884));
    layer1_outputs(37) <= layer0_outputs(697);
    layer1_outputs(38) <= not((layer0_outputs(5388)) and (layer0_outputs(7605)));
    layer1_outputs(39) <= (layer0_outputs(6451)) or (layer0_outputs(7567));
    layer1_outputs(40) <= not(layer0_outputs(1238));
    layer1_outputs(41) <= (layer0_outputs(839)) and not (layer0_outputs(4054));
    layer1_outputs(42) <= not((layer0_outputs(6055)) xor (layer0_outputs(3324)));
    layer1_outputs(43) <= not(layer0_outputs(3641)) or (layer0_outputs(4149));
    layer1_outputs(44) <= (layer0_outputs(4446)) and not (layer0_outputs(4758));
    layer1_outputs(45) <= not(layer0_outputs(6285));
    layer1_outputs(46) <= not(layer0_outputs(138)) or (layer0_outputs(6065));
    layer1_outputs(47) <= not(layer0_outputs(1487));
    layer1_outputs(48) <= (layer0_outputs(447)) and (layer0_outputs(4104));
    layer1_outputs(49) <= not(layer0_outputs(2382)) or (layer0_outputs(6032));
    layer1_outputs(50) <= not(layer0_outputs(7236));
    layer1_outputs(51) <= layer0_outputs(6507);
    layer1_outputs(52) <= (layer0_outputs(2183)) and not (layer0_outputs(6825));
    layer1_outputs(53) <= not(layer0_outputs(3847));
    layer1_outputs(54) <= layer0_outputs(4884);
    layer1_outputs(55) <= layer0_outputs(7208);
    layer1_outputs(56) <= (layer0_outputs(6909)) or (layer0_outputs(3178));
    layer1_outputs(57) <= layer0_outputs(993);
    layer1_outputs(58) <= not(layer0_outputs(2789));
    layer1_outputs(59) <= not(layer0_outputs(5748));
    layer1_outputs(60) <= not(layer0_outputs(6558));
    layer1_outputs(61) <= (layer0_outputs(1617)) and (layer0_outputs(3389));
    layer1_outputs(62) <= layer0_outputs(1421);
    layer1_outputs(63) <= (layer0_outputs(3387)) and not (layer0_outputs(396));
    layer1_outputs(64) <= '1';
    layer1_outputs(65) <= not(layer0_outputs(4464)) or (layer0_outputs(2562));
    layer1_outputs(66) <= not((layer0_outputs(4545)) or (layer0_outputs(195)));
    layer1_outputs(67) <= not(layer0_outputs(7398));
    layer1_outputs(68) <= not((layer0_outputs(1285)) xor (layer0_outputs(5975)));
    layer1_outputs(69) <= layer0_outputs(7422);
    layer1_outputs(70) <= not(layer0_outputs(3887)) or (layer0_outputs(1026));
    layer1_outputs(71) <= (layer0_outputs(4039)) and (layer0_outputs(2881));
    layer1_outputs(72) <= layer0_outputs(7661);
    layer1_outputs(73) <= not(layer0_outputs(4400));
    layer1_outputs(74) <= layer0_outputs(5230);
    layer1_outputs(75) <= (layer0_outputs(736)) and not (layer0_outputs(1831));
    layer1_outputs(76) <= (layer0_outputs(3988)) xor (layer0_outputs(2321));
    layer1_outputs(77) <= layer0_outputs(4049);
    layer1_outputs(78) <= '0';
    layer1_outputs(79) <= layer0_outputs(19);
    layer1_outputs(80) <= (layer0_outputs(6043)) or (layer0_outputs(6593));
    layer1_outputs(81) <= not(layer0_outputs(5670));
    layer1_outputs(82) <= not(layer0_outputs(2296));
    layer1_outputs(83) <= (layer0_outputs(4346)) and (layer0_outputs(4617));
    layer1_outputs(84) <= not(layer0_outputs(3621));
    layer1_outputs(85) <= (layer0_outputs(2757)) or (layer0_outputs(7679));
    layer1_outputs(86) <= (layer0_outputs(268)) or (layer0_outputs(5915));
    layer1_outputs(87) <= not(layer0_outputs(6806)) or (layer0_outputs(6336));
    layer1_outputs(88) <= '1';
    layer1_outputs(89) <= layer0_outputs(377);
    layer1_outputs(90) <= '1';
    layer1_outputs(91) <= (layer0_outputs(6943)) and not (layer0_outputs(2306));
    layer1_outputs(92) <= not(layer0_outputs(1645));
    layer1_outputs(93) <= (layer0_outputs(3310)) or (layer0_outputs(4813));
    layer1_outputs(94) <= not(layer0_outputs(2682)) or (layer0_outputs(4186));
    layer1_outputs(95) <= '1';
    layer1_outputs(96) <= layer0_outputs(2875);
    layer1_outputs(97) <= not((layer0_outputs(6323)) xor (layer0_outputs(6708)));
    layer1_outputs(98) <= not(layer0_outputs(6557));
    layer1_outputs(99) <= not((layer0_outputs(2242)) or (layer0_outputs(6058)));
    layer1_outputs(100) <= not((layer0_outputs(4614)) and (layer0_outputs(7102)));
    layer1_outputs(101) <= (layer0_outputs(66)) and not (layer0_outputs(5951));
    layer1_outputs(102) <= '0';
    layer1_outputs(103) <= not(layer0_outputs(1971));
    layer1_outputs(104) <= not((layer0_outputs(3206)) xor (layer0_outputs(7279)));
    layer1_outputs(105) <= (layer0_outputs(1241)) or (layer0_outputs(882));
    layer1_outputs(106) <= '1';
    layer1_outputs(107) <= '1';
    layer1_outputs(108) <= (layer0_outputs(5261)) and (layer0_outputs(5550));
    layer1_outputs(109) <= not(layer0_outputs(2162)) or (layer0_outputs(1957));
    layer1_outputs(110) <= (layer0_outputs(1763)) or (layer0_outputs(6373));
    layer1_outputs(111) <= (layer0_outputs(4711)) and (layer0_outputs(1649));
    layer1_outputs(112) <= (layer0_outputs(4634)) and not (layer0_outputs(5991));
    layer1_outputs(113) <= not(layer0_outputs(377));
    layer1_outputs(114) <= (layer0_outputs(4948)) and not (layer0_outputs(1638));
    layer1_outputs(115) <= not(layer0_outputs(3789)) or (layer0_outputs(436));
    layer1_outputs(116) <= not(layer0_outputs(2405)) or (layer0_outputs(910));
    layer1_outputs(117) <= '1';
    layer1_outputs(118) <= not(layer0_outputs(6139));
    layer1_outputs(119) <= not((layer0_outputs(6343)) or (layer0_outputs(2577)));
    layer1_outputs(120) <= (layer0_outputs(7180)) and not (layer0_outputs(6252));
    layer1_outputs(121) <= (layer0_outputs(293)) and not (layer0_outputs(4570));
    layer1_outputs(122) <= layer0_outputs(2172);
    layer1_outputs(123) <= layer0_outputs(3511);
    layer1_outputs(124) <= not(layer0_outputs(3541));
    layer1_outputs(125) <= layer0_outputs(1530);
    layer1_outputs(126) <= not(layer0_outputs(1680));
    layer1_outputs(127) <= (layer0_outputs(4906)) and (layer0_outputs(674));
    layer1_outputs(128) <= layer0_outputs(4495);
    layer1_outputs(129) <= not((layer0_outputs(4279)) xor (layer0_outputs(1771)));
    layer1_outputs(130) <= not(layer0_outputs(2543));
    layer1_outputs(131) <= not(layer0_outputs(6859)) or (layer0_outputs(6675));
    layer1_outputs(132) <= not(layer0_outputs(3152));
    layer1_outputs(133) <= (layer0_outputs(2927)) xor (layer0_outputs(4918));
    layer1_outputs(134) <= '0';
    layer1_outputs(135) <= '0';
    layer1_outputs(136) <= (layer0_outputs(5694)) xor (layer0_outputs(7539));
    layer1_outputs(137) <= not((layer0_outputs(6690)) and (layer0_outputs(6776)));
    layer1_outputs(138) <= (layer0_outputs(1289)) and not (layer0_outputs(4536));
    layer1_outputs(139) <= not((layer0_outputs(1128)) xor (layer0_outputs(7090)));
    layer1_outputs(140) <= '1';
    layer1_outputs(141) <= layer0_outputs(6584);
    layer1_outputs(142) <= layer0_outputs(5792);
    layer1_outputs(143) <= not(layer0_outputs(3702)) or (layer0_outputs(1041));
    layer1_outputs(144) <= not(layer0_outputs(7435));
    layer1_outputs(145) <= layer0_outputs(6515);
    layer1_outputs(146) <= '0';
    layer1_outputs(147) <= '0';
    layer1_outputs(148) <= layer0_outputs(147);
    layer1_outputs(149) <= not((layer0_outputs(6276)) and (layer0_outputs(6813)));
    layer1_outputs(150) <= not((layer0_outputs(3481)) xor (layer0_outputs(2460)));
    layer1_outputs(151) <= (layer0_outputs(1976)) and (layer0_outputs(4946));
    layer1_outputs(152) <= (layer0_outputs(2600)) and not (layer0_outputs(961));
    layer1_outputs(153) <= not((layer0_outputs(1775)) or (layer0_outputs(638)));
    layer1_outputs(154) <= not(layer0_outputs(3266)) or (layer0_outputs(1286));
    layer1_outputs(155) <= layer0_outputs(1829);
    layer1_outputs(156) <= layer0_outputs(4468);
    layer1_outputs(157) <= not((layer0_outputs(3913)) or (layer0_outputs(358)));
    layer1_outputs(158) <= (layer0_outputs(7602)) xor (layer0_outputs(3916));
    layer1_outputs(159) <= not((layer0_outputs(2898)) and (layer0_outputs(1674)));
    layer1_outputs(160) <= (layer0_outputs(384)) xor (layer0_outputs(4213));
    layer1_outputs(161) <= '1';
    layer1_outputs(162) <= not((layer0_outputs(6383)) xor (layer0_outputs(2136)));
    layer1_outputs(163) <= not(layer0_outputs(4587));
    layer1_outputs(164) <= not(layer0_outputs(5493));
    layer1_outputs(165) <= not(layer0_outputs(6988)) or (layer0_outputs(2108));
    layer1_outputs(166) <= (layer0_outputs(5644)) and not (layer0_outputs(2272));
    layer1_outputs(167) <= (layer0_outputs(4568)) and not (layer0_outputs(4393));
    layer1_outputs(168) <= '1';
    layer1_outputs(169) <= (layer0_outputs(2971)) and not (layer0_outputs(4445));
    layer1_outputs(170) <= (layer0_outputs(5277)) and not (layer0_outputs(5262));
    layer1_outputs(171) <= not(layer0_outputs(7298));
    layer1_outputs(172) <= not(layer0_outputs(266)) or (layer0_outputs(2792));
    layer1_outputs(173) <= layer0_outputs(456);
    layer1_outputs(174) <= '1';
    layer1_outputs(175) <= layer0_outputs(4955);
    layer1_outputs(176) <= (layer0_outputs(2120)) and not (layer0_outputs(5672));
    layer1_outputs(177) <= (layer0_outputs(2640)) or (layer0_outputs(7018));
    layer1_outputs(178) <= not((layer0_outputs(1682)) and (layer0_outputs(6307)));
    layer1_outputs(179) <= layer0_outputs(2752);
    layer1_outputs(180) <= not(layer0_outputs(1545));
    layer1_outputs(181) <= not(layer0_outputs(7432)) or (layer0_outputs(4386));
    layer1_outputs(182) <= (layer0_outputs(6034)) xor (layer0_outputs(5759));
    layer1_outputs(183) <= not(layer0_outputs(5754));
    layer1_outputs(184) <= layer0_outputs(6375);
    layer1_outputs(185) <= layer0_outputs(1270);
    layer1_outputs(186) <= (layer0_outputs(2586)) or (layer0_outputs(1159));
    layer1_outputs(187) <= not((layer0_outputs(7272)) and (layer0_outputs(3394)));
    layer1_outputs(188) <= (layer0_outputs(367)) and not (layer0_outputs(5909));
    layer1_outputs(189) <= '0';
    layer1_outputs(190) <= layer0_outputs(3336);
    layer1_outputs(191) <= layer0_outputs(1214);
    layer1_outputs(192) <= layer0_outputs(1189);
    layer1_outputs(193) <= not((layer0_outputs(914)) and (layer0_outputs(4690)));
    layer1_outputs(194) <= '0';
    layer1_outputs(195) <= not((layer0_outputs(5328)) and (layer0_outputs(3900)));
    layer1_outputs(196) <= not(layer0_outputs(1653)) or (layer0_outputs(2829));
    layer1_outputs(197) <= not(layer0_outputs(1800));
    layer1_outputs(198) <= not((layer0_outputs(6822)) or (layer0_outputs(2908)));
    layer1_outputs(199) <= (layer0_outputs(773)) or (layer0_outputs(7195));
    layer1_outputs(200) <= not((layer0_outputs(1253)) and (layer0_outputs(7317)));
    layer1_outputs(201) <= (layer0_outputs(4374)) or (layer0_outputs(4598));
    layer1_outputs(202) <= not((layer0_outputs(4977)) or (layer0_outputs(3643)));
    layer1_outputs(203) <= not((layer0_outputs(5675)) or (layer0_outputs(2713)));
    layer1_outputs(204) <= (layer0_outputs(5247)) and not (layer0_outputs(3066));
    layer1_outputs(205) <= not(layer0_outputs(5006));
    layer1_outputs(206) <= not(layer0_outputs(4361));
    layer1_outputs(207) <= not(layer0_outputs(5317));
    layer1_outputs(208) <= '1';
    layer1_outputs(209) <= not(layer0_outputs(7372));
    layer1_outputs(210) <= layer0_outputs(51);
    layer1_outputs(211) <= layer0_outputs(98);
    layer1_outputs(212) <= '1';
    layer1_outputs(213) <= '0';
    layer1_outputs(214) <= (layer0_outputs(4296)) or (layer0_outputs(473));
    layer1_outputs(215) <= (layer0_outputs(1189)) and (layer0_outputs(305));
    layer1_outputs(216) <= not((layer0_outputs(1032)) xor (layer0_outputs(221)));
    layer1_outputs(217) <= '0';
    layer1_outputs(218) <= layer0_outputs(2275);
    layer1_outputs(219) <= not(layer0_outputs(4676));
    layer1_outputs(220) <= '0';
    layer1_outputs(221) <= not(layer0_outputs(3260));
    layer1_outputs(222) <= (layer0_outputs(6673)) and (layer0_outputs(1095));
    layer1_outputs(223) <= not((layer0_outputs(6347)) and (layer0_outputs(2667)));
    layer1_outputs(224) <= not(layer0_outputs(6973));
    layer1_outputs(225) <= not(layer0_outputs(3453));
    layer1_outputs(226) <= not(layer0_outputs(3217));
    layer1_outputs(227) <= (layer0_outputs(6910)) or (layer0_outputs(5467));
    layer1_outputs(228) <= layer0_outputs(6072);
    layer1_outputs(229) <= (layer0_outputs(192)) and not (layer0_outputs(5854));
    layer1_outputs(230) <= layer0_outputs(7331);
    layer1_outputs(231) <= layer0_outputs(453);
    layer1_outputs(232) <= not(layer0_outputs(4828)) or (layer0_outputs(6366));
    layer1_outputs(233) <= not(layer0_outputs(1993));
    layer1_outputs(234) <= not(layer0_outputs(1120));
    layer1_outputs(235) <= not((layer0_outputs(4247)) and (layer0_outputs(6665)));
    layer1_outputs(236) <= not((layer0_outputs(2014)) or (layer0_outputs(6793)));
    layer1_outputs(237) <= not((layer0_outputs(3283)) and (layer0_outputs(3305)));
    layer1_outputs(238) <= layer0_outputs(2070);
    layer1_outputs(239) <= not(layer0_outputs(2846));
    layer1_outputs(240) <= layer0_outputs(7011);
    layer1_outputs(241) <= not((layer0_outputs(5907)) or (layer0_outputs(7284)));
    layer1_outputs(242) <= (layer0_outputs(7480)) or (layer0_outputs(3275));
    layer1_outputs(243) <= not((layer0_outputs(2498)) or (layer0_outputs(2125)));
    layer1_outputs(244) <= not((layer0_outputs(6433)) or (layer0_outputs(4589)));
    layer1_outputs(245) <= not(layer0_outputs(3888));
    layer1_outputs(246) <= (layer0_outputs(3927)) xor (layer0_outputs(1648));
    layer1_outputs(247) <= (layer0_outputs(3418)) or (layer0_outputs(7022));
    layer1_outputs(248) <= (layer0_outputs(1402)) and not (layer0_outputs(1745));
    layer1_outputs(249) <= (layer0_outputs(2926)) and (layer0_outputs(2958));
    layer1_outputs(250) <= not(layer0_outputs(2033));
    layer1_outputs(251) <= (layer0_outputs(7158)) and not (layer0_outputs(7023));
    layer1_outputs(252) <= layer0_outputs(1009);
    layer1_outputs(253) <= (layer0_outputs(461)) and not (layer0_outputs(4732));
    layer1_outputs(254) <= layer0_outputs(3432);
    layer1_outputs(255) <= layer0_outputs(2121);
    layer1_outputs(256) <= not(layer0_outputs(391)) or (layer0_outputs(6766));
    layer1_outputs(257) <= (layer0_outputs(4752)) and (layer0_outputs(1106));
    layer1_outputs(258) <= not(layer0_outputs(3225)) or (layer0_outputs(2685));
    layer1_outputs(259) <= (layer0_outputs(982)) and (layer0_outputs(3739));
    layer1_outputs(260) <= (layer0_outputs(4055)) or (layer0_outputs(7500));
    layer1_outputs(261) <= '0';
    layer1_outputs(262) <= not(layer0_outputs(2262));
    layer1_outputs(263) <= (layer0_outputs(1231)) and not (layer0_outputs(4058));
    layer1_outputs(264) <= (layer0_outputs(7551)) and not (layer0_outputs(4488));
    layer1_outputs(265) <= not(layer0_outputs(3326)) or (layer0_outputs(1686));
    layer1_outputs(266) <= not(layer0_outputs(60));
    layer1_outputs(267) <= not(layer0_outputs(2959));
    layer1_outputs(268) <= not(layer0_outputs(2641));
    layer1_outputs(269) <= not((layer0_outputs(7446)) and (layer0_outputs(4292)));
    layer1_outputs(270) <= (layer0_outputs(7045)) and not (layer0_outputs(3373));
    layer1_outputs(271) <= (layer0_outputs(5206)) and (layer0_outputs(7024));
    layer1_outputs(272) <= not(layer0_outputs(6121)) or (layer0_outputs(6145));
    layer1_outputs(273) <= (layer0_outputs(7186)) or (layer0_outputs(3847));
    layer1_outputs(274) <= (layer0_outputs(4886)) or (layer0_outputs(7157));
    layer1_outputs(275) <= layer0_outputs(5135);
    layer1_outputs(276) <= not((layer0_outputs(4418)) and (layer0_outputs(7417)));
    layer1_outputs(277) <= not(layer0_outputs(1204));
    layer1_outputs(278) <= '1';
    layer1_outputs(279) <= not((layer0_outputs(936)) or (layer0_outputs(182)));
    layer1_outputs(280) <= (layer0_outputs(6247)) or (layer0_outputs(2624));
    layer1_outputs(281) <= (layer0_outputs(6569)) or (layer0_outputs(3118));
    layer1_outputs(282) <= not(layer0_outputs(2963)) or (layer0_outputs(6296));
    layer1_outputs(283) <= layer0_outputs(3209);
    layer1_outputs(284) <= layer0_outputs(4683);
    layer1_outputs(285) <= (layer0_outputs(4458)) or (layer0_outputs(6442));
    layer1_outputs(286) <= layer0_outputs(2259);
    layer1_outputs(287) <= not((layer0_outputs(6799)) or (layer0_outputs(234)));
    layer1_outputs(288) <= (layer0_outputs(6461)) and not (layer0_outputs(6827));
    layer1_outputs(289) <= not(layer0_outputs(1088));
    layer1_outputs(290) <= not(layer0_outputs(7583));
    layer1_outputs(291) <= layer0_outputs(4485);
    layer1_outputs(292) <= not((layer0_outputs(6759)) and (layer0_outputs(7197)));
    layer1_outputs(293) <= (layer0_outputs(4604)) or (layer0_outputs(7581));
    layer1_outputs(294) <= not(layer0_outputs(1270));
    layer1_outputs(295) <= (layer0_outputs(277)) and not (layer0_outputs(1673));
    layer1_outputs(296) <= layer0_outputs(3581);
    layer1_outputs(297) <= (layer0_outputs(5793)) xor (layer0_outputs(1906));
    layer1_outputs(298) <= not((layer0_outputs(4435)) and (layer0_outputs(4980)));
    layer1_outputs(299) <= not(layer0_outputs(4769));
    layer1_outputs(300) <= layer0_outputs(2205);
    layer1_outputs(301) <= (layer0_outputs(970)) or (layer0_outputs(1572));
    layer1_outputs(302) <= not(layer0_outputs(551));
    layer1_outputs(303) <= not(layer0_outputs(4647));
    layer1_outputs(304) <= layer0_outputs(800);
    layer1_outputs(305) <= (layer0_outputs(6997)) xor (layer0_outputs(3352));
    layer1_outputs(306) <= not(layer0_outputs(2319)) or (layer0_outputs(7224));
    layer1_outputs(307) <= '0';
    layer1_outputs(308) <= (layer0_outputs(7503)) and (layer0_outputs(2776));
    layer1_outputs(309) <= not(layer0_outputs(2639));
    layer1_outputs(310) <= (layer0_outputs(5905)) or (layer0_outputs(6869));
    layer1_outputs(311) <= (layer0_outputs(115)) or (layer0_outputs(6530));
    layer1_outputs(312) <= (layer0_outputs(6211)) and (layer0_outputs(7320));
    layer1_outputs(313) <= not(layer0_outputs(4059));
    layer1_outputs(314) <= not(layer0_outputs(5982));
    layer1_outputs(315) <= not((layer0_outputs(5105)) or (layer0_outputs(2905)));
    layer1_outputs(316) <= layer0_outputs(1183);
    layer1_outputs(317) <= not(layer0_outputs(6982));
    layer1_outputs(318) <= not(layer0_outputs(5044)) or (layer0_outputs(0));
    layer1_outputs(319) <= layer0_outputs(148);
    layer1_outputs(320) <= layer0_outputs(5994);
    layer1_outputs(321) <= not(layer0_outputs(7465)) or (layer0_outputs(2690));
    layer1_outputs(322) <= layer0_outputs(4631);
    layer1_outputs(323) <= not(layer0_outputs(3594));
    layer1_outputs(324) <= not((layer0_outputs(4153)) xor (layer0_outputs(7559)));
    layer1_outputs(325) <= (layer0_outputs(3451)) or (layer0_outputs(2196));
    layer1_outputs(326) <= not(layer0_outputs(2204));
    layer1_outputs(327) <= not(layer0_outputs(5435));
    layer1_outputs(328) <= (layer0_outputs(585)) and not (layer0_outputs(17));
    layer1_outputs(329) <= not((layer0_outputs(1434)) xor (layer0_outputs(6931)));
    layer1_outputs(330) <= (layer0_outputs(3425)) xor (layer0_outputs(4958));
    layer1_outputs(331) <= not(layer0_outputs(4721));
    layer1_outputs(332) <= '1';
    layer1_outputs(333) <= (layer0_outputs(151)) or (layer0_outputs(4415));
    layer1_outputs(334) <= not((layer0_outputs(1220)) xor (layer0_outputs(1986)));
    layer1_outputs(335) <= not((layer0_outputs(205)) and (layer0_outputs(2232)));
    layer1_outputs(336) <= (layer0_outputs(5995)) and (layer0_outputs(1516));
    layer1_outputs(337) <= (layer0_outputs(136)) and (layer0_outputs(2326));
    layer1_outputs(338) <= (layer0_outputs(6897)) and not (layer0_outputs(4429));
    layer1_outputs(339) <= not(layer0_outputs(5369));
    layer1_outputs(340) <= not(layer0_outputs(766)) or (layer0_outputs(3740));
    layer1_outputs(341) <= not(layer0_outputs(1654));
    layer1_outputs(342) <= (layer0_outputs(4059)) and (layer0_outputs(3223));
    layer1_outputs(343) <= layer0_outputs(5264);
    layer1_outputs(344) <= not(layer0_outputs(1087));
    layer1_outputs(345) <= layer0_outputs(988);
    layer1_outputs(346) <= '1';
    layer1_outputs(347) <= (layer0_outputs(6599)) or (layer0_outputs(2723));
    layer1_outputs(348) <= not((layer0_outputs(6750)) or (layer0_outputs(2419)));
    layer1_outputs(349) <= not((layer0_outputs(4966)) and (layer0_outputs(1550)));
    layer1_outputs(350) <= '1';
    layer1_outputs(351) <= '1';
    layer1_outputs(352) <= (layer0_outputs(2276)) and (layer0_outputs(3300));
    layer1_outputs(353) <= not(layer0_outputs(4526));
    layer1_outputs(354) <= not(layer0_outputs(6420));
    layer1_outputs(355) <= (layer0_outputs(1983)) or (layer0_outputs(4000));
    layer1_outputs(356) <= not(layer0_outputs(3379)) or (layer0_outputs(322));
    layer1_outputs(357) <= not(layer0_outputs(2991));
    layer1_outputs(358) <= '0';
    layer1_outputs(359) <= layer0_outputs(990);
    layer1_outputs(360) <= not(layer0_outputs(5243));
    layer1_outputs(361) <= '1';
    layer1_outputs(362) <= layer0_outputs(6619);
    layer1_outputs(363) <= (layer0_outputs(5801)) or (layer0_outputs(6280));
    layer1_outputs(364) <= not((layer0_outputs(1025)) or (layer0_outputs(5439)));
    layer1_outputs(365) <= not(layer0_outputs(5443));
    layer1_outputs(366) <= (layer0_outputs(7028)) and not (layer0_outputs(1741));
    layer1_outputs(367) <= (layer0_outputs(1215)) and not (layer0_outputs(3019));
    layer1_outputs(368) <= not(layer0_outputs(3747));
    layer1_outputs(369) <= not(layer0_outputs(2445)) or (layer0_outputs(5980));
    layer1_outputs(370) <= not(layer0_outputs(1360));
    layer1_outputs(371) <= layer0_outputs(1814);
    layer1_outputs(372) <= not(layer0_outputs(705)) or (layer0_outputs(800));
    layer1_outputs(373) <= not(layer0_outputs(5546)) or (layer0_outputs(2682));
    layer1_outputs(374) <= not(layer0_outputs(2868)) or (layer0_outputs(2711));
    layer1_outputs(375) <= (layer0_outputs(5568)) and not (layer0_outputs(2141));
    layer1_outputs(376) <= (layer0_outputs(2982)) and not (layer0_outputs(4746));
    layer1_outputs(377) <= (layer0_outputs(4708)) and (layer0_outputs(848));
    layer1_outputs(378) <= not(layer0_outputs(5616));
    layer1_outputs(379) <= not((layer0_outputs(7643)) and (layer0_outputs(4455)));
    layer1_outputs(380) <= layer0_outputs(6810);
    layer1_outputs(381) <= not(layer0_outputs(6029));
    layer1_outputs(382) <= (layer0_outputs(2699)) and (layer0_outputs(5237));
    layer1_outputs(383) <= (layer0_outputs(1229)) and not (layer0_outputs(1979));
    layer1_outputs(384) <= (layer0_outputs(4249)) xor (layer0_outputs(1207));
    layer1_outputs(385) <= layer0_outputs(5588);
    layer1_outputs(386) <= (layer0_outputs(5137)) or (layer0_outputs(1391));
    layer1_outputs(387) <= not((layer0_outputs(854)) and (layer0_outputs(4870)));
    layer1_outputs(388) <= not(layer0_outputs(2582)) or (layer0_outputs(4430));
    layer1_outputs(389) <= not(layer0_outputs(2988));
    layer1_outputs(390) <= layer0_outputs(3336);
    layer1_outputs(391) <= not((layer0_outputs(1758)) or (layer0_outputs(3030)));
    layer1_outputs(392) <= not(layer0_outputs(3818)) or (layer0_outputs(3924));
    layer1_outputs(393) <= (layer0_outputs(4318)) and not (layer0_outputs(3906));
    layer1_outputs(394) <= (layer0_outputs(5004)) and not (layer0_outputs(2492));
    layer1_outputs(395) <= layer0_outputs(3139);
    layer1_outputs(396) <= layer0_outputs(864);
    layer1_outputs(397) <= not(layer0_outputs(3303)) or (layer0_outputs(5654));
    layer1_outputs(398) <= (layer0_outputs(7451)) or (layer0_outputs(7035));
    layer1_outputs(399) <= (layer0_outputs(4701)) and not (layer0_outputs(1037));
    layer1_outputs(400) <= not((layer0_outputs(7577)) and (layer0_outputs(3197)));
    layer1_outputs(401) <= (layer0_outputs(6443)) and not (layer0_outputs(4468));
    layer1_outputs(402) <= '0';
    layer1_outputs(403) <= not(layer0_outputs(3156));
    layer1_outputs(404) <= (layer0_outputs(3086)) or (layer0_outputs(72));
    layer1_outputs(405) <= (layer0_outputs(5478)) and not (layer0_outputs(980));
    layer1_outputs(406) <= layer0_outputs(351);
    layer1_outputs(407) <= (layer0_outputs(3626)) and not (layer0_outputs(1797));
    layer1_outputs(408) <= '1';
    layer1_outputs(409) <= not((layer0_outputs(5364)) or (layer0_outputs(7166)));
    layer1_outputs(410) <= not(layer0_outputs(5645));
    layer1_outputs(411) <= (layer0_outputs(220)) and not (layer0_outputs(5988));
    layer1_outputs(412) <= layer0_outputs(7528);
    layer1_outputs(413) <= not(layer0_outputs(900));
    layer1_outputs(414) <= not(layer0_outputs(4605));
    layer1_outputs(415) <= '1';
    layer1_outputs(416) <= layer0_outputs(4055);
    layer1_outputs(417) <= '0';
    layer1_outputs(418) <= not((layer0_outputs(2129)) or (layer0_outputs(2517)));
    layer1_outputs(419) <= not((layer0_outputs(1406)) and (layer0_outputs(3591)));
    layer1_outputs(420) <= '0';
    layer1_outputs(421) <= layer0_outputs(501);
    layer1_outputs(422) <= (layer0_outputs(7191)) and not (layer0_outputs(3865));
    layer1_outputs(423) <= (layer0_outputs(1275)) and not (layer0_outputs(2605));
    layer1_outputs(424) <= '0';
    layer1_outputs(425) <= not(layer0_outputs(3485)) or (layer0_outputs(7009));
    layer1_outputs(426) <= '1';
    layer1_outputs(427) <= layer0_outputs(3819);
    layer1_outputs(428) <= not(layer0_outputs(6106));
    layer1_outputs(429) <= (layer0_outputs(1716)) xor (layer0_outputs(2044));
    layer1_outputs(430) <= (layer0_outputs(724)) and not (layer0_outputs(2096));
    layer1_outputs(431) <= layer0_outputs(6737);
    layer1_outputs(432) <= (layer0_outputs(4914)) and not (layer0_outputs(7303));
    layer1_outputs(433) <= not(layer0_outputs(4424));
    layer1_outputs(434) <= not(layer0_outputs(1738)) or (layer0_outputs(684));
    layer1_outputs(435) <= (layer0_outputs(3844)) and not (layer0_outputs(7465));
    layer1_outputs(436) <= not(layer0_outputs(4576));
    layer1_outputs(437) <= not((layer0_outputs(2902)) and (layer0_outputs(98)));
    layer1_outputs(438) <= (layer0_outputs(6075)) xor (layer0_outputs(4447));
    layer1_outputs(439) <= not(layer0_outputs(4559));
    layer1_outputs(440) <= '1';
    layer1_outputs(441) <= not(layer0_outputs(2294));
    layer1_outputs(442) <= layer0_outputs(2500);
    layer1_outputs(443) <= not((layer0_outputs(2629)) or (layer0_outputs(5236)));
    layer1_outputs(444) <= layer0_outputs(4938);
    layer1_outputs(445) <= not(layer0_outputs(2409));
    layer1_outputs(446) <= '1';
    layer1_outputs(447) <= not(layer0_outputs(6679)) or (layer0_outputs(423));
    layer1_outputs(448) <= (layer0_outputs(6604)) and not (layer0_outputs(3393));
    layer1_outputs(449) <= (layer0_outputs(4220)) and not (layer0_outputs(1356));
    layer1_outputs(450) <= (layer0_outputs(920)) xor (layer0_outputs(6538));
    layer1_outputs(451) <= not(layer0_outputs(3368));
    layer1_outputs(452) <= not(layer0_outputs(7540));
    layer1_outputs(453) <= (layer0_outputs(5114)) or (layer0_outputs(7362));
    layer1_outputs(454) <= (layer0_outputs(4625)) xor (layer0_outputs(6091));
    layer1_outputs(455) <= (layer0_outputs(1854)) or (layer0_outputs(6165));
    layer1_outputs(456) <= layer0_outputs(7047);
    layer1_outputs(457) <= layer0_outputs(1372);
    layer1_outputs(458) <= (layer0_outputs(813)) xor (layer0_outputs(5823));
    layer1_outputs(459) <= not(layer0_outputs(1531)) or (layer0_outputs(4041));
    layer1_outputs(460) <= not(layer0_outputs(4588)) or (layer0_outputs(2697));
    layer1_outputs(461) <= not(layer0_outputs(292));
    layer1_outputs(462) <= not((layer0_outputs(1465)) or (layer0_outputs(5816)));
    layer1_outputs(463) <= '1';
    layer1_outputs(464) <= layer0_outputs(859);
    layer1_outputs(465) <= (layer0_outputs(2484)) and not (layer0_outputs(2902));
    layer1_outputs(466) <= (layer0_outputs(2660)) and not (layer0_outputs(6281));
    layer1_outputs(467) <= '1';
    layer1_outputs(468) <= not(layer0_outputs(7518));
    layer1_outputs(469) <= layer0_outputs(4470);
    layer1_outputs(470) <= not(layer0_outputs(4076));
    layer1_outputs(471) <= not((layer0_outputs(5165)) or (layer0_outputs(1670)));
    layer1_outputs(472) <= (layer0_outputs(1620)) and not (layer0_outputs(3430));
    layer1_outputs(473) <= not(layer0_outputs(7041)) or (layer0_outputs(7670));
    layer1_outputs(474) <= (layer0_outputs(1173)) and (layer0_outputs(4709));
    layer1_outputs(475) <= (layer0_outputs(189)) xor (layer0_outputs(2374));
    layer1_outputs(476) <= (layer0_outputs(7618)) and not (layer0_outputs(2462));
    layer1_outputs(477) <= not(layer0_outputs(2269));
    layer1_outputs(478) <= layer0_outputs(1914);
    layer1_outputs(479) <= not(layer0_outputs(2689)) or (layer0_outputs(6250));
    layer1_outputs(480) <= not(layer0_outputs(6760));
    layer1_outputs(481) <= (layer0_outputs(978)) or (layer0_outputs(997));
    layer1_outputs(482) <= layer0_outputs(2257);
    layer1_outputs(483) <= not(layer0_outputs(2236));
    layer1_outputs(484) <= (layer0_outputs(2677)) or (layer0_outputs(2857));
    layer1_outputs(485) <= not(layer0_outputs(4922));
    layer1_outputs(486) <= not(layer0_outputs(2901));
    layer1_outputs(487) <= not(layer0_outputs(849));
    layer1_outputs(488) <= '0';
    layer1_outputs(489) <= not((layer0_outputs(4773)) and (layer0_outputs(3443)));
    layer1_outputs(490) <= '0';
    layer1_outputs(491) <= not(layer0_outputs(836));
    layer1_outputs(492) <= (layer0_outputs(1560)) xor (layer0_outputs(83));
    layer1_outputs(493) <= not(layer0_outputs(3528));
    layer1_outputs(494) <= not(layer0_outputs(4690)) or (layer0_outputs(3181));
    layer1_outputs(495) <= not((layer0_outputs(4275)) and (layer0_outputs(2082)));
    layer1_outputs(496) <= (layer0_outputs(3154)) and not (layer0_outputs(7548));
    layer1_outputs(497) <= not(layer0_outputs(6689));
    layer1_outputs(498) <= '1';
    layer1_outputs(499) <= (layer0_outputs(3588)) and not (layer0_outputs(7534));
    layer1_outputs(500) <= layer0_outputs(1875);
    layer1_outputs(501) <= not((layer0_outputs(4313)) xor (layer0_outputs(4174)));
    layer1_outputs(502) <= not(layer0_outputs(3788));
    layer1_outputs(503) <= not((layer0_outputs(817)) or (layer0_outputs(1085)));
    layer1_outputs(504) <= not(layer0_outputs(127));
    layer1_outputs(505) <= layer0_outputs(3081);
    layer1_outputs(506) <= not(layer0_outputs(3301));
    layer1_outputs(507) <= not((layer0_outputs(3330)) and (layer0_outputs(2532)));
    layer1_outputs(508) <= not(layer0_outputs(2922));
    layer1_outputs(509) <= (layer0_outputs(6540)) and (layer0_outputs(4618));
    layer1_outputs(510) <= not((layer0_outputs(735)) and (layer0_outputs(6220)));
    layer1_outputs(511) <= (layer0_outputs(1853)) or (layer0_outputs(1476));
    layer1_outputs(512) <= not(layer0_outputs(498));
    layer1_outputs(513) <= not(layer0_outputs(506));
    layer1_outputs(514) <= (layer0_outputs(7660)) and not (layer0_outputs(3921));
    layer1_outputs(515) <= not((layer0_outputs(7298)) and (layer0_outputs(2093)));
    layer1_outputs(516) <= (layer0_outputs(5116)) and not (layer0_outputs(3276));
    layer1_outputs(517) <= layer0_outputs(1495);
    layer1_outputs(518) <= not(layer0_outputs(4319));
    layer1_outputs(519) <= (layer0_outputs(4708)) or (layer0_outputs(4373));
    layer1_outputs(520) <= not((layer0_outputs(1375)) xor (layer0_outputs(4248)));
    layer1_outputs(521) <= not(layer0_outputs(2005));
    layer1_outputs(522) <= '0';
    layer1_outputs(523) <= layer0_outputs(6884);
    layer1_outputs(524) <= not(layer0_outputs(5428));
    layer1_outputs(525) <= layer0_outputs(4147);
    layer1_outputs(526) <= '0';
    layer1_outputs(527) <= not((layer0_outputs(6685)) xor (layer0_outputs(4962)));
    layer1_outputs(528) <= not(layer0_outputs(3713)) or (layer0_outputs(4298));
    layer1_outputs(529) <= '1';
    layer1_outputs(530) <= not(layer0_outputs(6179));
    layer1_outputs(531) <= layer0_outputs(3205);
    layer1_outputs(532) <= not(layer0_outputs(1565)) or (layer0_outputs(519));
    layer1_outputs(533) <= (layer0_outputs(6403)) and not (layer0_outputs(6157));
    layer1_outputs(534) <= (layer0_outputs(3518)) and not (layer0_outputs(5127));
    layer1_outputs(535) <= layer0_outputs(6594);
    layer1_outputs(536) <= not(layer0_outputs(3832));
    layer1_outputs(537) <= '0';
    layer1_outputs(538) <= (layer0_outputs(6257)) or (layer0_outputs(3821));
    layer1_outputs(539) <= not(layer0_outputs(3584)) or (layer0_outputs(7323));
    layer1_outputs(540) <= (layer0_outputs(4163)) or (layer0_outputs(4199));
    layer1_outputs(541) <= '0';
    layer1_outputs(542) <= not(layer0_outputs(1340)) or (layer0_outputs(2371));
    layer1_outputs(543) <= layer0_outputs(4368);
    layer1_outputs(544) <= (layer0_outputs(3331)) and not (layer0_outputs(6244));
    layer1_outputs(545) <= not(layer0_outputs(2006));
    layer1_outputs(546) <= not(layer0_outputs(4910));
    layer1_outputs(547) <= layer0_outputs(928);
    layer1_outputs(548) <= (layer0_outputs(2654)) and not (layer0_outputs(4222));
    layer1_outputs(549) <= '1';
    layer1_outputs(550) <= (layer0_outputs(6125)) or (layer0_outputs(2640));
    layer1_outputs(551) <= not(layer0_outputs(2233));
    layer1_outputs(552) <= '1';
    layer1_outputs(553) <= not(layer0_outputs(1086));
    layer1_outputs(554) <= not((layer0_outputs(5633)) and (layer0_outputs(832)));
    layer1_outputs(555) <= layer0_outputs(995);
    layer1_outputs(556) <= not(layer0_outputs(7435)) or (layer0_outputs(7555));
    layer1_outputs(557) <= layer0_outputs(3091);
    layer1_outputs(558) <= layer0_outputs(3326);
    layer1_outputs(559) <= not(layer0_outputs(7511)) or (layer0_outputs(1029));
    layer1_outputs(560) <= layer0_outputs(1194);
    layer1_outputs(561) <= not((layer0_outputs(6528)) and (layer0_outputs(7019)));
    layer1_outputs(562) <= layer0_outputs(4483);
    layer1_outputs(563) <= layer0_outputs(1989);
    layer1_outputs(564) <= not(layer0_outputs(6843));
    layer1_outputs(565) <= layer0_outputs(1918);
    layer1_outputs(566) <= not(layer0_outputs(6440));
    layer1_outputs(567) <= '1';
    layer1_outputs(568) <= not((layer0_outputs(86)) xor (layer0_outputs(1774)));
    layer1_outputs(569) <= (layer0_outputs(5327)) or (layer0_outputs(336));
    layer1_outputs(570) <= '1';
    layer1_outputs(571) <= (layer0_outputs(4647)) or (layer0_outputs(68));
    layer1_outputs(572) <= not(layer0_outputs(5359));
    layer1_outputs(573) <= (layer0_outputs(1366)) xor (layer0_outputs(4272));
    layer1_outputs(574) <= not(layer0_outputs(5105));
    layer1_outputs(575) <= not(layer0_outputs(3994));
    layer1_outputs(576) <= not((layer0_outputs(526)) xor (layer0_outputs(2581)));
    layer1_outputs(577) <= not(layer0_outputs(70));
    layer1_outputs(578) <= layer0_outputs(1791);
    layer1_outputs(579) <= layer0_outputs(1483);
    layer1_outputs(580) <= not(layer0_outputs(3762)) or (layer0_outputs(5264));
    layer1_outputs(581) <= not(layer0_outputs(7051));
    layer1_outputs(582) <= (layer0_outputs(5767)) or (layer0_outputs(126));
    layer1_outputs(583) <= layer0_outputs(2123);
    layer1_outputs(584) <= not((layer0_outputs(10)) or (layer0_outputs(3698)));
    layer1_outputs(585) <= '1';
    layer1_outputs(586) <= not(layer0_outputs(6934));
    layer1_outputs(587) <= (layer0_outputs(1469)) and not (layer0_outputs(6835));
    layer1_outputs(588) <= '0';
    layer1_outputs(589) <= not((layer0_outputs(3278)) and (layer0_outputs(2234)));
    layer1_outputs(590) <= '1';
    layer1_outputs(591) <= '0';
    layer1_outputs(592) <= not(layer0_outputs(5055));
    layer1_outputs(593) <= not(layer0_outputs(1801));
    layer1_outputs(594) <= not(layer0_outputs(7046)) or (layer0_outputs(7593));
    layer1_outputs(595) <= layer0_outputs(3943);
    layer1_outputs(596) <= (layer0_outputs(1664)) and (layer0_outputs(2022));
    layer1_outputs(597) <= (layer0_outputs(3392)) and (layer0_outputs(5116));
    layer1_outputs(598) <= not((layer0_outputs(4313)) or (layer0_outputs(6492)));
    layer1_outputs(599) <= '0';
    layer1_outputs(600) <= '1';
    layer1_outputs(601) <= not(layer0_outputs(6707)) or (layer0_outputs(887));
    layer1_outputs(602) <= not((layer0_outputs(888)) or (layer0_outputs(562)));
    layer1_outputs(603) <= not(layer0_outputs(5255));
    layer1_outputs(604) <= '0';
    layer1_outputs(605) <= '0';
    layer1_outputs(606) <= not(layer0_outputs(1595)) or (layer0_outputs(4830));
    layer1_outputs(607) <= layer0_outputs(4737);
    layer1_outputs(608) <= not(layer0_outputs(4204)) or (layer0_outputs(7192));
    layer1_outputs(609) <= layer0_outputs(3579);
    layer1_outputs(610) <= not(layer0_outputs(7166)) or (layer0_outputs(78));
    layer1_outputs(611) <= not(layer0_outputs(4988));
    layer1_outputs(612) <= (layer0_outputs(6711)) and not (layer0_outputs(3074));
    layer1_outputs(613) <= not(layer0_outputs(3891));
    layer1_outputs(614) <= not(layer0_outputs(2469)) or (layer0_outputs(5475));
    layer1_outputs(615) <= not((layer0_outputs(6939)) or (layer0_outputs(2791)));
    layer1_outputs(616) <= '1';
    layer1_outputs(617) <= not(layer0_outputs(4356)) or (layer0_outputs(6013));
    layer1_outputs(618) <= not((layer0_outputs(1712)) xor (layer0_outputs(233)));
    layer1_outputs(619) <= not((layer0_outputs(3822)) or (layer0_outputs(4654)));
    layer1_outputs(620) <= not((layer0_outputs(5312)) or (layer0_outputs(2755)));
    layer1_outputs(621) <= layer0_outputs(625);
    layer1_outputs(622) <= not(layer0_outputs(1735)) or (layer0_outputs(5464));
    layer1_outputs(623) <= '0';
    layer1_outputs(624) <= '1';
    layer1_outputs(625) <= not(layer0_outputs(5106));
    layer1_outputs(626) <= not(layer0_outputs(169));
    layer1_outputs(627) <= not(layer0_outputs(6274));
    layer1_outputs(628) <= (layer0_outputs(5954)) or (layer0_outputs(6987));
    layer1_outputs(629) <= '1';
    layer1_outputs(630) <= not(layer0_outputs(5521));
    layer1_outputs(631) <= (layer0_outputs(1947)) and not (layer0_outputs(441));
    layer1_outputs(632) <= '1';
    layer1_outputs(633) <= (layer0_outputs(939)) and not (layer0_outputs(7646));
    layer1_outputs(634) <= (layer0_outputs(2810)) or (layer0_outputs(2352));
    layer1_outputs(635) <= not((layer0_outputs(1463)) or (layer0_outputs(157)));
    layer1_outputs(636) <= not((layer0_outputs(987)) or (layer0_outputs(7355)));
    layer1_outputs(637) <= not(layer0_outputs(3639));
    layer1_outputs(638) <= layer0_outputs(253);
    layer1_outputs(639) <= layer0_outputs(5238);
    layer1_outputs(640) <= (layer0_outputs(3506)) and not (layer0_outputs(2619));
    layer1_outputs(641) <= not((layer0_outputs(5266)) or (layer0_outputs(31)));
    layer1_outputs(642) <= not((layer0_outputs(3586)) and (layer0_outputs(3753)));
    layer1_outputs(643) <= (layer0_outputs(4349)) and not (layer0_outputs(7500));
    layer1_outputs(644) <= layer0_outputs(5182);
    layer1_outputs(645) <= not(layer0_outputs(5088));
    layer1_outputs(646) <= (layer0_outputs(383)) or (layer0_outputs(7116));
    layer1_outputs(647) <= '0';
    layer1_outputs(648) <= not((layer0_outputs(2495)) and (layer0_outputs(3601)));
    layer1_outputs(649) <= not(layer0_outputs(6228));
    layer1_outputs(650) <= not((layer0_outputs(4308)) or (layer0_outputs(1610)));
    layer1_outputs(651) <= not(layer0_outputs(2160)) or (layer0_outputs(6687));
    layer1_outputs(652) <= not((layer0_outputs(3243)) xor (layer0_outputs(7219)));
    layer1_outputs(653) <= not(layer0_outputs(3167)) or (layer0_outputs(1640));
    layer1_outputs(654) <= not(layer0_outputs(7387));
    layer1_outputs(655) <= (layer0_outputs(2816)) and not (layer0_outputs(1666));
    layer1_outputs(656) <= not(layer0_outputs(6969));
    layer1_outputs(657) <= not((layer0_outputs(6522)) or (layer0_outputs(3995)));
    layer1_outputs(658) <= not(layer0_outputs(6398)) or (layer0_outputs(2070));
    layer1_outputs(659) <= layer0_outputs(5984);
    layer1_outputs(660) <= layer0_outputs(6800);
    layer1_outputs(661) <= (layer0_outputs(5727)) and not (layer0_outputs(2071));
    layer1_outputs(662) <= not(layer0_outputs(2937));
    layer1_outputs(663) <= '0';
    layer1_outputs(664) <= '0';
    layer1_outputs(665) <= (layer0_outputs(3059)) and (layer0_outputs(3094));
    layer1_outputs(666) <= not(layer0_outputs(6802)) or (layer0_outputs(4017));
    layer1_outputs(667) <= (layer0_outputs(2291)) or (layer0_outputs(1290));
    layer1_outputs(668) <= layer0_outputs(559);
    layer1_outputs(669) <= (layer0_outputs(4080)) or (layer0_outputs(4437));
    layer1_outputs(670) <= layer0_outputs(4337);
    layer1_outputs(671) <= layer0_outputs(3907);
    layer1_outputs(672) <= not(layer0_outputs(4922));
    layer1_outputs(673) <= not(layer0_outputs(5510)) or (layer0_outputs(2620));
    layer1_outputs(674) <= not(layer0_outputs(6750));
    layer1_outputs(675) <= not(layer0_outputs(6208)) or (layer0_outputs(330));
    layer1_outputs(676) <= not((layer0_outputs(6111)) xor (layer0_outputs(4338)));
    layer1_outputs(677) <= not(layer0_outputs(7036));
    layer1_outputs(678) <= '0';
    layer1_outputs(679) <= not(layer0_outputs(7537));
    layer1_outputs(680) <= (layer0_outputs(7245)) xor (layer0_outputs(6689));
    layer1_outputs(681) <= not(layer0_outputs(1435)) or (layer0_outputs(589));
    layer1_outputs(682) <= not((layer0_outputs(2485)) and (layer0_outputs(5757)));
    layer1_outputs(683) <= (layer0_outputs(6795)) and not (layer0_outputs(4084));
    layer1_outputs(684) <= not(layer0_outputs(1088));
    layer1_outputs(685) <= not(layer0_outputs(2096));
    layer1_outputs(686) <= (layer0_outputs(4377)) or (layer0_outputs(840));
    layer1_outputs(687) <= not(layer0_outputs(7119));
    layer1_outputs(688) <= layer0_outputs(1213);
    layer1_outputs(689) <= (layer0_outputs(349)) and (layer0_outputs(313));
    layer1_outputs(690) <= not((layer0_outputs(3410)) or (layer0_outputs(5018)));
    layer1_outputs(691) <= layer0_outputs(6743);
    layer1_outputs(692) <= layer0_outputs(6787);
    layer1_outputs(693) <= (layer0_outputs(3004)) and not (layer0_outputs(2117));
    layer1_outputs(694) <= layer0_outputs(6486);
    layer1_outputs(695) <= '0';
    layer1_outputs(696) <= not(layer0_outputs(7188)) or (layer0_outputs(363));
    layer1_outputs(697) <= '1';
    layer1_outputs(698) <= not(layer0_outputs(3637));
    layer1_outputs(699) <= not((layer0_outputs(7024)) and (layer0_outputs(4522)));
    layer1_outputs(700) <= (layer0_outputs(1689)) and (layer0_outputs(4310));
    layer1_outputs(701) <= not(layer0_outputs(363));
    layer1_outputs(702) <= '1';
    layer1_outputs(703) <= (layer0_outputs(2531)) and not (layer0_outputs(4125));
    layer1_outputs(704) <= not(layer0_outputs(1352));
    layer1_outputs(705) <= (layer0_outputs(3941)) and not (layer0_outputs(2677));
    layer1_outputs(706) <= not(layer0_outputs(514));
    layer1_outputs(707) <= '0';
    layer1_outputs(708) <= not(layer0_outputs(1448));
    layer1_outputs(709) <= (layer0_outputs(2059)) or (layer0_outputs(1224));
    layer1_outputs(710) <= not(layer0_outputs(6432)) or (layer0_outputs(7492));
    layer1_outputs(711) <= layer0_outputs(4091);
    layer1_outputs(712) <= not((layer0_outputs(6098)) and (layer0_outputs(6940)));
    layer1_outputs(713) <= not(layer0_outputs(7393));
    layer1_outputs(714) <= layer0_outputs(3251);
    layer1_outputs(715) <= not(layer0_outputs(4624));
    layer1_outputs(716) <= not(layer0_outputs(7275));
    layer1_outputs(717) <= not((layer0_outputs(6556)) and (layer0_outputs(3133)));
    layer1_outputs(718) <= (layer0_outputs(4875)) and not (layer0_outputs(3903));
    layer1_outputs(719) <= (layer0_outputs(7604)) and not (layer0_outputs(1031));
    layer1_outputs(720) <= (layer0_outputs(3286)) and not (layer0_outputs(814));
    layer1_outputs(721) <= (layer0_outputs(3746)) and (layer0_outputs(979));
    layer1_outputs(722) <= layer0_outputs(7572);
    layer1_outputs(723) <= layer0_outputs(5886);
    layer1_outputs(724) <= not((layer0_outputs(6170)) and (layer0_outputs(575)));
    layer1_outputs(725) <= layer0_outputs(5404);
    layer1_outputs(726) <= not(layer0_outputs(645)) or (layer0_outputs(6146));
    layer1_outputs(727) <= layer0_outputs(4911);
    layer1_outputs(728) <= (layer0_outputs(468)) and not (layer0_outputs(4817));
    layer1_outputs(729) <= not(layer0_outputs(5575));
    layer1_outputs(730) <= not((layer0_outputs(7415)) or (layer0_outputs(1696)));
    layer1_outputs(731) <= '1';
    layer1_outputs(732) <= not(layer0_outputs(345));
    layer1_outputs(733) <= not(layer0_outputs(4688)) or (layer0_outputs(3604));
    layer1_outputs(734) <= layer0_outputs(3856);
    layer1_outputs(735) <= (layer0_outputs(824)) and not (layer0_outputs(6923));
    layer1_outputs(736) <= (layer0_outputs(4444)) and not (layer0_outputs(5278));
    layer1_outputs(737) <= (layer0_outputs(2742)) and not (layer0_outputs(6758));
    layer1_outputs(738) <= not(layer0_outputs(7662));
    layer1_outputs(739) <= not(layer0_outputs(729)) or (layer0_outputs(546));
    layer1_outputs(740) <= not(layer0_outputs(1476));
    layer1_outputs(741) <= not((layer0_outputs(6338)) or (layer0_outputs(2545)));
    layer1_outputs(742) <= not(layer0_outputs(7455)) or (layer0_outputs(567));
    layer1_outputs(743) <= not(layer0_outputs(281)) or (layer0_outputs(5504));
    layer1_outputs(744) <= '0';
    layer1_outputs(745) <= not((layer0_outputs(7521)) and (layer0_outputs(1534)));
    layer1_outputs(746) <= not(layer0_outputs(6221));
    layer1_outputs(747) <= not(layer0_outputs(4465));
    layer1_outputs(748) <= (layer0_outputs(6190)) or (layer0_outputs(4335));
    layer1_outputs(749) <= layer0_outputs(7121);
    layer1_outputs(750) <= '1';
    layer1_outputs(751) <= '1';
    layer1_outputs(752) <= not((layer0_outputs(5711)) and (layer0_outputs(22)));
    layer1_outputs(753) <= layer0_outputs(1330);
    layer1_outputs(754) <= not(layer0_outputs(2257));
    layer1_outputs(755) <= layer0_outputs(2802);
    layer1_outputs(756) <= not(layer0_outputs(4835)) or (layer0_outputs(578));
    layer1_outputs(757) <= '0';
    layer1_outputs(758) <= not(layer0_outputs(6978));
    layer1_outputs(759) <= not((layer0_outputs(215)) or (layer0_outputs(7265)));
    layer1_outputs(760) <= layer0_outputs(2951);
    layer1_outputs(761) <= layer0_outputs(1436);
    layer1_outputs(762) <= not(layer0_outputs(3803)) or (layer0_outputs(2407));
    layer1_outputs(763) <= (layer0_outputs(1719)) and not (layer0_outputs(5295));
    layer1_outputs(764) <= (layer0_outputs(1781)) and (layer0_outputs(7300));
    layer1_outputs(765) <= not(layer0_outputs(1626));
    layer1_outputs(766) <= (layer0_outputs(3089)) and not (layer0_outputs(1307));
    layer1_outputs(767) <= not((layer0_outputs(791)) and (layer0_outputs(6509)));
    layer1_outputs(768) <= (layer0_outputs(7275)) and not (layer0_outputs(3114));
    layer1_outputs(769) <= (layer0_outputs(3501)) or (layer0_outputs(7289));
    layer1_outputs(770) <= not(layer0_outputs(2592));
    layer1_outputs(771) <= (layer0_outputs(2477)) and (layer0_outputs(6916));
    layer1_outputs(772) <= not((layer0_outputs(879)) and (layer0_outputs(2393)));
    layer1_outputs(773) <= layer0_outputs(1570);
    layer1_outputs(774) <= '0';
    layer1_outputs(775) <= not(layer0_outputs(3923)) or (layer0_outputs(5873));
    layer1_outputs(776) <= not((layer0_outputs(4291)) or (layer0_outputs(5331)));
    layer1_outputs(777) <= (layer0_outputs(7070)) and (layer0_outputs(5985));
    layer1_outputs(778) <= not(layer0_outputs(6591));
    layer1_outputs(779) <= (layer0_outputs(3464)) or (layer0_outputs(5349));
    layer1_outputs(780) <= not((layer0_outputs(7026)) xor (layer0_outputs(2473)));
    layer1_outputs(781) <= (layer0_outputs(5686)) and not (layer0_outputs(5476));
    layer1_outputs(782) <= '0';
    layer1_outputs(783) <= '0';
    layer1_outputs(784) <= not(layer0_outputs(2795));
    layer1_outputs(785) <= '1';
    layer1_outputs(786) <= (layer0_outputs(1109)) or (layer0_outputs(958));
    layer1_outputs(787) <= not(layer0_outputs(5109));
    layer1_outputs(788) <= '0';
    layer1_outputs(789) <= (layer0_outputs(4307)) or (layer0_outputs(5902));
    layer1_outputs(790) <= layer0_outputs(4474);
    layer1_outputs(791) <= (layer0_outputs(3281)) or (layer0_outputs(5925));
    layer1_outputs(792) <= not(layer0_outputs(4840));
    layer1_outputs(793) <= not((layer0_outputs(1016)) or (layer0_outputs(4182)));
    layer1_outputs(794) <= not(layer0_outputs(6902));
    layer1_outputs(795) <= (layer0_outputs(6927)) and not (layer0_outputs(5729));
    layer1_outputs(796) <= not(layer0_outputs(818)) or (layer0_outputs(4172));
    layer1_outputs(797) <= not((layer0_outputs(5258)) xor (layer0_outputs(7519)));
    layer1_outputs(798) <= not((layer0_outputs(3669)) or (layer0_outputs(4373)));
    layer1_outputs(799) <= layer0_outputs(7663);
    layer1_outputs(800) <= layer0_outputs(6124);
    layer1_outputs(801) <= not((layer0_outputs(4992)) or (layer0_outputs(527)));
    layer1_outputs(802) <= (layer0_outputs(953)) and not (layer0_outputs(7467));
    layer1_outputs(803) <= not((layer0_outputs(382)) or (layer0_outputs(2428)));
    layer1_outputs(804) <= not(layer0_outputs(5855));
    layer1_outputs(805) <= not(layer0_outputs(7262));
    layer1_outputs(806) <= (layer0_outputs(54)) or (layer0_outputs(1340));
    layer1_outputs(807) <= '1';
    layer1_outputs(808) <= '0';
    layer1_outputs(809) <= '0';
    layer1_outputs(810) <= '1';
    layer1_outputs(811) <= not((layer0_outputs(7423)) xor (layer0_outputs(7499)));
    layer1_outputs(812) <= not((layer0_outputs(699)) and (layer0_outputs(1048)));
    layer1_outputs(813) <= layer0_outputs(2387);
    layer1_outputs(814) <= not(layer0_outputs(6555));
    layer1_outputs(815) <= (layer0_outputs(380)) and not (layer0_outputs(295));
    layer1_outputs(816) <= not(layer0_outputs(5060));
    layer1_outputs(817) <= layer0_outputs(7129);
    layer1_outputs(818) <= not(layer0_outputs(5152));
    layer1_outputs(819) <= (layer0_outputs(739)) and not (layer0_outputs(7415));
    layer1_outputs(820) <= not(layer0_outputs(7484));
    layer1_outputs(821) <= (layer0_outputs(647)) or (layer0_outputs(5768));
    layer1_outputs(822) <= layer0_outputs(3650);
    layer1_outputs(823) <= not(layer0_outputs(5913));
    layer1_outputs(824) <= layer0_outputs(325);
    layer1_outputs(825) <= not(layer0_outputs(2006));
    layer1_outputs(826) <= (layer0_outputs(6916)) and not (layer0_outputs(2148));
    layer1_outputs(827) <= not((layer0_outputs(3939)) xor (layer0_outputs(5207)));
    layer1_outputs(828) <= layer0_outputs(6164);
    layer1_outputs(829) <= layer0_outputs(4194);
    layer1_outputs(830) <= not((layer0_outputs(4335)) or (layer0_outputs(5417)));
    layer1_outputs(831) <= (layer0_outputs(5932)) or (layer0_outputs(5242));
    layer1_outputs(832) <= not(layer0_outputs(4130));
    layer1_outputs(833) <= (layer0_outputs(7118)) and not (layer0_outputs(6672));
    layer1_outputs(834) <= layer0_outputs(1374);
    layer1_outputs(835) <= layer0_outputs(471);
    layer1_outputs(836) <= (layer0_outputs(4539)) and not (layer0_outputs(6842));
    layer1_outputs(837) <= not(layer0_outputs(1706));
    layer1_outputs(838) <= '1';
    layer1_outputs(839) <= (layer0_outputs(3501)) or (layer0_outputs(5090));
    layer1_outputs(840) <= not((layer0_outputs(3679)) or (layer0_outputs(5292)));
    layer1_outputs(841) <= (layer0_outputs(2002)) and not (layer0_outputs(5068));
    layer1_outputs(842) <= layer0_outputs(663);
    layer1_outputs(843) <= not(layer0_outputs(4069));
    layer1_outputs(844) <= not((layer0_outputs(1225)) and (layer0_outputs(958)));
    layer1_outputs(845) <= layer0_outputs(6018);
    layer1_outputs(846) <= (layer0_outputs(6639)) or (layer0_outputs(3064));
    layer1_outputs(847) <= not(layer0_outputs(28)) or (layer0_outputs(4934));
    layer1_outputs(848) <= not(layer0_outputs(5318)) or (layer0_outputs(5344));
    layer1_outputs(849) <= not((layer0_outputs(2282)) or (layer0_outputs(3372)));
    layer1_outputs(850) <= (layer0_outputs(617)) or (layer0_outputs(5365));
    layer1_outputs(851) <= '1';
    layer1_outputs(852) <= (layer0_outputs(1174)) and not (layer0_outputs(55));
    layer1_outputs(853) <= layer0_outputs(850);
    layer1_outputs(854) <= not(layer0_outputs(5226));
    layer1_outputs(855) <= (layer0_outputs(4859)) and (layer0_outputs(6933));
    layer1_outputs(856) <= (layer0_outputs(239)) and not (layer0_outputs(308));
    layer1_outputs(857) <= layer0_outputs(4435);
    layer1_outputs(858) <= not(layer0_outputs(3462));
    layer1_outputs(859) <= not(layer0_outputs(7523));
    layer1_outputs(860) <= not((layer0_outputs(301)) or (layer0_outputs(1543)));
    layer1_outputs(861) <= (layer0_outputs(4900)) and (layer0_outputs(3602));
    layer1_outputs(862) <= not((layer0_outputs(6181)) or (layer0_outputs(5029)));
    layer1_outputs(863) <= not((layer0_outputs(3780)) xor (layer0_outputs(2922)));
    layer1_outputs(864) <= not(layer0_outputs(7615));
    layer1_outputs(865) <= not((layer0_outputs(5185)) and (layer0_outputs(556)));
    layer1_outputs(866) <= (layer0_outputs(1750)) and (layer0_outputs(1306));
    layer1_outputs(867) <= not(layer0_outputs(209));
    layer1_outputs(868) <= (layer0_outputs(2287)) and not (layer0_outputs(6779));
    layer1_outputs(869) <= not(layer0_outputs(4266));
    layer1_outputs(870) <= not(layer0_outputs(3905));
    layer1_outputs(871) <= not(layer0_outputs(1050));
    layer1_outputs(872) <= '0';
    layer1_outputs(873) <= (layer0_outputs(7263)) and not (layer0_outputs(2817));
    layer1_outputs(874) <= not(layer0_outputs(1464));
    layer1_outputs(875) <= layer0_outputs(465);
    layer1_outputs(876) <= not((layer0_outputs(3713)) xor (layer0_outputs(5372)));
    layer1_outputs(877) <= (layer0_outputs(256)) or (layer0_outputs(4951));
    layer1_outputs(878) <= (layer0_outputs(1719)) or (layer0_outputs(3820));
    layer1_outputs(879) <= not(layer0_outputs(7434));
    layer1_outputs(880) <= (layer0_outputs(2893)) and (layer0_outputs(2949));
    layer1_outputs(881) <= layer0_outputs(303);
    layer1_outputs(882) <= not(layer0_outputs(4677));
    layer1_outputs(883) <= not(layer0_outputs(3551)) or (layer0_outputs(1449));
    layer1_outputs(884) <= (layer0_outputs(7000)) or (layer0_outputs(140));
    layer1_outputs(885) <= not((layer0_outputs(3784)) and (layer0_outputs(6332)));
    layer1_outputs(886) <= not(layer0_outputs(2369)) or (layer0_outputs(5218));
    layer1_outputs(887) <= not((layer0_outputs(3766)) or (layer0_outputs(3129)));
    layer1_outputs(888) <= (layer0_outputs(1291)) xor (layer0_outputs(6331));
    layer1_outputs(889) <= not((layer0_outputs(5979)) xor (layer0_outputs(6730)));
    layer1_outputs(890) <= layer0_outputs(2019);
    layer1_outputs(891) <= (layer0_outputs(6123)) and not (layer0_outputs(5095));
    layer1_outputs(892) <= layer0_outputs(4729);
    layer1_outputs(893) <= '0';
    layer1_outputs(894) <= layer0_outputs(2911);
    layer1_outputs(895) <= layer0_outputs(3053);
    layer1_outputs(896) <= not(layer0_outputs(2293));
    layer1_outputs(897) <= not(layer0_outputs(2991));
    layer1_outputs(898) <= (layer0_outputs(1369)) and not (layer0_outputs(76));
    layer1_outputs(899) <= not(layer0_outputs(4607)) or (layer0_outputs(163));
    layer1_outputs(900) <= (layer0_outputs(7030)) xor (layer0_outputs(1561));
    layer1_outputs(901) <= (layer0_outputs(546)) xor (layer0_outputs(5296));
    layer1_outputs(902) <= '1';
    layer1_outputs(903) <= layer0_outputs(727);
    layer1_outputs(904) <= layer0_outputs(1786);
    layer1_outputs(905) <= (layer0_outputs(3474)) or (layer0_outputs(5019));
    layer1_outputs(906) <= not(layer0_outputs(2278));
    layer1_outputs(907) <= layer0_outputs(827);
    layer1_outputs(908) <= layer0_outputs(265);
    layer1_outputs(909) <= '1';
    layer1_outputs(910) <= '1';
    layer1_outputs(911) <= layer0_outputs(3355);
    layer1_outputs(912) <= not(layer0_outputs(2206));
    layer1_outputs(913) <= not(layer0_outputs(5063)) or (layer0_outputs(6597));
    layer1_outputs(914) <= not(layer0_outputs(2646)) or (layer0_outputs(940));
    layer1_outputs(915) <= '0';
    layer1_outputs(916) <= layer0_outputs(3873);
    layer1_outputs(917) <= not(layer0_outputs(3918)) or (layer0_outputs(5705));
    layer1_outputs(918) <= '0';
    layer1_outputs(919) <= not(layer0_outputs(6991));
    layer1_outputs(920) <= not(layer0_outputs(5244));
    layer1_outputs(921) <= '1';
    layer1_outputs(922) <= layer0_outputs(4331);
    layer1_outputs(923) <= (layer0_outputs(6532)) or (layer0_outputs(7258));
    layer1_outputs(924) <= not((layer0_outputs(6990)) xor (layer0_outputs(1371)));
    layer1_outputs(925) <= layer0_outputs(6493);
    layer1_outputs(926) <= (layer0_outputs(3569)) and (layer0_outputs(4519));
    layer1_outputs(927) <= (layer0_outputs(185)) and (layer0_outputs(1081));
    layer1_outputs(928) <= not(layer0_outputs(6317)) or (layer0_outputs(3789));
    layer1_outputs(929) <= not(layer0_outputs(4757)) or (layer0_outputs(6446));
    layer1_outputs(930) <= not((layer0_outputs(3092)) or (layer0_outputs(4628)));
    layer1_outputs(931) <= not(layer0_outputs(7198));
    layer1_outputs(932) <= not(layer0_outputs(314));
    layer1_outputs(933) <= '1';
    layer1_outputs(934) <= layer0_outputs(5085);
    layer1_outputs(935) <= layer0_outputs(3253);
    layer1_outputs(936) <= (layer0_outputs(4937)) and not (layer0_outputs(1272));
    layer1_outputs(937) <= (layer0_outputs(4795)) and (layer0_outputs(32));
    layer1_outputs(938) <= not(layer0_outputs(481));
    layer1_outputs(939) <= not((layer0_outputs(4606)) and (layer0_outputs(5181)));
    layer1_outputs(940) <= not(layer0_outputs(541)) or (layer0_outputs(560));
    layer1_outputs(941) <= (layer0_outputs(1756)) and not (layer0_outputs(5290));
    layer1_outputs(942) <= layer0_outputs(1318);
    layer1_outputs(943) <= not((layer0_outputs(2167)) and (layer0_outputs(17)));
    layer1_outputs(944) <= (layer0_outputs(4535)) and (layer0_outputs(5889));
    layer1_outputs(945) <= layer0_outputs(4881);
    layer1_outputs(946) <= layer0_outputs(4848);
    layer1_outputs(947) <= (layer0_outputs(1924)) or (layer0_outputs(2249));
    layer1_outputs(948) <= not(layer0_outputs(974)) or (layer0_outputs(3199));
    layer1_outputs(949) <= '1';
    layer1_outputs(950) <= (layer0_outputs(1666)) and (layer0_outputs(6911));
    layer1_outputs(951) <= (layer0_outputs(3264)) and (layer0_outputs(5662));
    layer1_outputs(952) <= not(layer0_outputs(3733)) or (layer0_outputs(407));
    layer1_outputs(953) <= '1';
    layer1_outputs(954) <= not(layer0_outputs(4869));
    layer1_outputs(955) <= not((layer0_outputs(4560)) or (layer0_outputs(4751)));
    layer1_outputs(956) <= layer0_outputs(4327);
    layer1_outputs(957) <= not((layer0_outputs(5495)) and (layer0_outputs(1689)));
    layer1_outputs(958) <= not((layer0_outputs(5535)) or (layer0_outputs(584)));
    layer1_outputs(959) <= not(layer0_outputs(1364)) or (layer0_outputs(6524));
    layer1_outputs(960) <= not(layer0_outputs(2519)) or (layer0_outputs(3745));
    layer1_outputs(961) <= (layer0_outputs(6251)) and not (layer0_outputs(4358));
    layer1_outputs(962) <= layer0_outputs(2159);
    layer1_outputs(963) <= not(layer0_outputs(1252)) or (layer0_outputs(7477));
    layer1_outputs(964) <= not((layer0_outputs(7546)) and (layer0_outputs(6466)));
    layer1_outputs(965) <= (layer0_outputs(3076)) and not (layer0_outputs(7182));
    layer1_outputs(966) <= not(layer0_outputs(3570)) or (layer0_outputs(1355));
    layer1_outputs(967) <= not(layer0_outputs(3175));
    layer1_outputs(968) <= not((layer0_outputs(6237)) or (layer0_outputs(3930)));
    layer1_outputs(969) <= not(layer0_outputs(2438));
    layer1_outputs(970) <= (layer0_outputs(6159)) and not (layer0_outputs(2948));
    layer1_outputs(971) <= not(layer0_outputs(202)) or (layer0_outputs(1397));
    layer1_outputs(972) <= not((layer0_outputs(2526)) and (layer0_outputs(5439)));
    layer1_outputs(973) <= layer0_outputs(3419);
    layer1_outputs(974) <= not((layer0_outputs(1465)) and (layer0_outputs(3837)));
    layer1_outputs(975) <= layer0_outputs(4847);
    layer1_outputs(976) <= (layer0_outputs(3693)) or (layer0_outputs(3425));
    layer1_outputs(977) <= (layer0_outputs(5744)) and not (layer0_outputs(6100));
    layer1_outputs(978) <= '0';
    layer1_outputs(979) <= not(layer0_outputs(2867));
    layer1_outputs(980) <= not((layer0_outputs(7252)) and (layer0_outputs(6972)));
    layer1_outputs(981) <= (layer0_outputs(5963)) and (layer0_outputs(5313));
    layer1_outputs(982) <= layer0_outputs(5289);
    layer1_outputs(983) <= '0';
    layer1_outputs(984) <= (layer0_outputs(191)) or (layer0_outputs(1093));
    layer1_outputs(985) <= not(layer0_outputs(495)) or (layer0_outputs(3262));
    layer1_outputs(986) <= (layer0_outputs(1325)) or (layer0_outputs(630));
    layer1_outputs(987) <= not(layer0_outputs(3252));
    layer1_outputs(988) <= not((layer0_outputs(5588)) or (layer0_outputs(5536)));
    layer1_outputs(989) <= not(layer0_outputs(5926));
    layer1_outputs(990) <= layer0_outputs(2749);
    layer1_outputs(991) <= layer0_outputs(1363);
    layer1_outputs(992) <= (layer0_outputs(5028)) and (layer0_outputs(1821));
    layer1_outputs(993) <= (layer0_outputs(5117)) and not (layer0_outputs(1905));
    layer1_outputs(994) <= layer0_outputs(2065);
    layer1_outputs(995) <= not(layer0_outputs(3118)) or (layer0_outputs(5104));
    layer1_outputs(996) <= layer0_outputs(1214);
    layer1_outputs(997) <= (layer0_outputs(5881)) xor (layer0_outputs(429));
    layer1_outputs(998) <= '0';
    layer1_outputs(999) <= (layer0_outputs(2141)) or (layer0_outputs(5436));
    layer1_outputs(1000) <= '0';
    layer1_outputs(1001) <= not(layer0_outputs(24)) or (layer0_outputs(5233));
    layer1_outputs(1002) <= not(layer0_outputs(5846)) or (layer0_outputs(6938));
    layer1_outputs(1003) <= not(layer0_outputs(6005));
    layer1_outputs(1004) <= not(layer0_outputs(7635));
    layer1_outputs(1005) <= (layer0_outputs(1764)) and (layer0_outputs(6754));
    layer1_outputs(1006) <= layer0_outputs(442);
    layer1_outputs(1007) <= layer0_outputs(6017);
    layer1_outputs(1008) <= not((layer0_outputs(7255)) or (layer0_outputs(1863)));
    layer1_outputs(1009) <= (layer0_outputs(5494)) and (layer0_outputs(2899));
    layer1_outputs(1010) <= not((layer0_outputs(6010)) xor (layer0_outputs(229)));
    layer1_outputs(1011) <= (layer0_outputs(2084)) xor (layer0_outputs(871));
    layer1_outputs(1012) <= (layer0_outputs(3988)) and not (layer0_outputs(3673));
    layer1_outputs(1013) <= '1';
    layer1_outputs(1014) <= not(layer0_outputs(1378)) or (layer0_outputs(5270));
    layer1_outputs(1015) <= not((layer0_outputs(1566)) or (layer0_outputs(6324)));
    layer1_outputs(1016) <= not(layer0_outputs(4829)) or (layer0_outputs(631));
    layer1_outputs(1017) <= not((layer0_outputs(3040)) xor (layer0_outputs(6583)));
    layer1_outputs(1018) <= layer0_outputs(4882);
    layer1_outputs(1019) <= layer0_outputs(3802);
    layer1_outputs(1020) <= (layer0_outputs(5628)) and (layer0_outputs(3850));
    layer1_outputs(1021) <= not(layer0_outputs(4806));
    layer1_outputs(1022) <= not(layer0_outputs(3672)) or (layer0_outputs(5393));
    layer1_outputs(1023) <= not((layer0_outputs(4763)) or (layer0_outputs(6269)));
    layer1_outputs(1024) <= not((layer0_outputs(877)) xor (layer0_outputs(7167)));
    layer1_outputs(1025) <= layer0_outputs(7554);
    layer1_outputs(1026) <= (layer0_outputs(743)) and not (layer0_outputs(3890));
    layer1_outputs(1027) <= not(layer0_outputs(346));
    layer1_outputs(1028) <= layer0_outputs(4549);
    layer1_outputs(1029) <= (layer0_outputs(3570)) and (layer0_outputs(5425));
    layer1_outputs(1030) <= not(layer0_outputs(6728));
    layer1_outputs(1031) <= not(layer0_outputs(4651)) or (layer0_outputs(1765));
    layer1_outputs(1032) <= not(layer0_outputs(5203));
    layer1_outputs(1033) <= layer0_outputs(3356);
    layer1_outputs(1034) <= (layer0_outputs(4025)) or (layer0_outputs(3961));
    layer1_outputs(1035) <= (layer0_outputs(2942)) and not (layer0_outputs(6771));
    layer1_outputs(1036) <= not((layer0_outputs(3979)) or (layer0_outputs(1780)));
    layer1_outputs(1037) <= (layer0_outputs(3874)) or (layer0_outputs(4821));
    layer1_outputs(1038) <= layer0_outputs(5195);
    layer1_outputs(1039) <= not(layer0_outputs(5960));
    layer1_outputs(1040) <= not(layer0_outputs(2637)) or (layer0_outputs(170));
    layer1_outputs(1041) <= not(layer0_outputs(1927)) or (layer0_outputs(5973));
    layer1_outputs(1042) <= not(layer0_outputs(928));
    layer1_outputs(1043) <= not(layer0_outputs(3096));
    layer1_outputs(1044) <= (layer0_outputs(269)) or (layer0_outputs(152));
    layer1_outputs(1045) <= '1';
    layer1_outputs(1046) <= layer0_outputs(1977);
    layer1_outputs(1047) <= not(layer0_outputs(3585));
    layer1_outputs(1048) <= '1';
    layer1_outputs(1049) <= (layer0_outputs(2385)) and (layer0_outputs(3352));
    layer1_outputs(1050) <= not(layer0_outputs(1736));
    layer1_outputs(1051) <= layer0_outputs(7077);
    layer1_outputs(1052) <= layer0_outputs(1810);
    layer1_outputs(1053) <= layer0_outputs(2293);
    layer1_outputs(1054) <= layer0_outputs(6944);
    layer1_outputs(1055) <= layer0_outputs(4393);
    layer1_outputs(1056) <= (layer0_outputs(554)) and not (layer0_outputs(4510));
    layer1_outputs(1057) <= (layer0_outputs(4501)) or (layer0_outputs(2165));
    layer1_outputs(1058) <= not((layer0_outputs(276)) or (layer0_outputs(1005)));
    layer1_outputs(1059) <= layer0_outputs(2352);
    layer1_outputs(1060) <= not(layer0_outputs(3623));
    layer1_outputs(1061) <= (layer0_outputs(4820)) or (layer0_outputs(7293));
    layer1_outputs(1062) <= layer0_outputs(3652);
    layer1_outputs(1063) <= not(layer0_outputs(2180));
    layer1_outputs(1064) <= (layer0_outputs(6087)) and (layer0_outputs(3117));
    layer1_outputs(1065) <= not((layer0_outputs(502)) and (layer0_outputs(3869)));
    layer1_outputs(1066) <= layer0_outputs(7521);
    layer1_outputs(1067) <= (layer0_outputs(2950)) and not (layer0_outputs(5325));
    layer1_outputs(1068) <= not(layer0_outputs(2997));
    layer1_outputs(1069) <= layer0_outputs(478);
    layer1_outputs(1070) <= (layer0_outputs(4795)) and not (layer0_outputs(3162));
    layer1_outputs(1071) <= not(layer0_outputs(5944)) or (layer0_outputs(2222));
    layer1_outputs(1072) <= not(layer0_outputs(914)) or (layer0_outputs(4290));
    layer1_outputs(1073) <= layer0_outputs(1651);
    layer1_outputs(1074) <= not((layer0_outputs(1343)) and (layer0_outputs(986)));
    layer1_outputs(1075) <= '0';
    layer1_outputs(1076) <= not((layer0_outputs(2619)) and (layer0_outputs(1533)));
    layer1_outputs(1077) <= (layer0_outputs(2254)) and not (layer0_outputs(5208));
    layer1_outputs(1078) <= (layer0_outputs(7639)) and (layer0_outputs(1426));
    layer1_outputs(1079) <= not(layer0_outputs(919));
    layer1_outputs(1080) <= (layer0_outputs(3016)) and (layer0_outputs(2875));
    layer1_outputs(1081) <= (layer0_outputs(6361)) and not (layer0_outputs(6732));
    layer1_outputs(1082) <= layer0_outputs(6386);
    layer1_outputs(1083) <= not(layer0_outputs(518));
    layer1_outputs(1084) <= (layer0_outputs(2729)) or (layer0_outputs(3529));
    layer1_outputs(1085) <= layer0_outputs(4726);
    layer1_outputs(1086) <= (layer0_outputs(6637)) or (layer0_outputs(5276));
    layer1_outputs(1087) <= not(layer0_outputs(743));
    layer1_outputs(1088) <= (layer0_outputs(6206)) or (layer0_outputs(7109));
    layer1_outputs(1089) <= not(layer0_outputs(6505)) or (layer0_outputs(4683));
    layer1_outputs(1090) <= not(layer0_outputs(7575));
    layer1_outputs(1091) <= (layer0_outputs(347)) and (layer0_outputs(3940));
    layer1_outputs(1092) <= not(layer0_outputs(1296));
    layer1_outputs(1093) <= not(layer0_outputs(811));
    layer1_outputs(1094) <= not(layer0_outputs(1433)) or (layer0_outputs(5266));
    layer1_outputs(1095) <= not(layer0_outputs(3087));
    layer1_outputs(1096) <= '0';
    layer1_outputs(1097) <= layer0_outputs(3686);
    layer1_outputs(1098) <= not((layer0_outputs(3860)) or (layer0_outputs(1438)));
    layer1_outputs(1099) <= not((layer0_outputs(2538)) or (layer0_outputs(20)));
    layer1_outputs(1100) <= not((layer0_outputs(2027)) or (layer0_outputs(4054)));
    layer1_outputs(1101) <= not((layer0_outputs(3984)) xor (layer0_outputs(7429)));
    layer1_outputs(1102) <= (layer0_outputs(692)) and not (layer0_outputs(3248));
    layer1_outputs(1103) <= not((layer0_outputs(7111)) xor (layer0_outputs(6951)));
    layer1_outputs(1104) <= (layer0_outputs(3460)) and not (layer0_outputs(342));
    layer1_outputs(1105) <= layer0_outputs(4682);
    layer1_outputs(1106) <= (layer0_outputs(6993)) and (layer0_outputs(7085));
    layer1_outputs(1107) <= not(layer0_outputs(1651));
    layer1_outputs(1108) <= (layer0_outputs(3632)) or (layer0_outputs(6531));
    layer1_outputs(1109) <= not(layer0_outputs(2471));
    layer1_outputs(1110) <= not(layer0_outputs(2012)) or (layer0_outputs(5440));
    layer1_outputs(1111) <= not(layer0_outputs(4224));
    layer1_outputs(1112) <= (layer0_outputs(1752)) and not (layer0_outputs(247));
    layer1_outputs(1113) <= not((layer0_outputs(2980)) xor (layer0_outputs(7283)));
    layer1_outputs(1114) <= not((layer0_outputs(2475)) and (layer0_outputs(4537)));
    layer1_outputs(1115) <= not(layer0_outputs(5138)) or (layer0_outputs(497));
    layer1_outputs(1116) <= not(layer0_outputs(6489));
    layer1_outputs(1117) <= not((layer0_outputs(7069)) or (layer0_outputs(4466)));
    layer1_outputs(1118) <= not(layer0_outputs(3395)) or (layer0_outputs(31));
    layer1_outputs(1119) <= layer0_outputs(6566);
    layer1_outputs(1120) <= layer0_outputs(2534);
    layer1_outputs(1121) <= not(layer0_outputs(5392));
    layer1_outputs(1122) <= not((layer0_outputs(4623)) and (layer0_outputs(2966)));
    layer1_outputs(1123) <= layer0_outputs(172);
    layer1_outputs(1124) <= not(layer0_outputs(2137));
    layer1_outputs(1125) <= not(layer0_outputs(2224));
    layer1_outputs(1126) <= '1';
    layer1_outputs(1127) <= not((layer0_outputs(3163)) and (layer0_outputs(1772)));
    layer1_outputs(1128) <= not(layer0_outputs(662));
    layer1_outputs(1129) <= not(layer0_outputs(387)) or (layer0_outputs(5722));
    layer1_outputs(1130) <= not(layer0_outputs(2113));
    layer1_outputs(1131) <= layer0_outputs(7594);
    layer1_outputs(1132) <= (layer0_outputs(6818)) and (layer0_outputs(684));
    layer1_outputs(1133) <= (layer0_outputs(6628)) or (layer0_outputs(2428));
    layer1_outputs(1134) <= not(layer0_outputs(7463));
    layer1_outputs(1135) <= '0';
    layer1_outputs(1136) <= not(layer0_outputs(5916));
    layer1_outputs(1137) <= layer0_outputs(7136);
    layer1_outputs(1138) <= not(layer0_outputs(1779)) or (layer0_outputs(2935));
    layer1_outputs(1139) <= (layer0_outputs(5689)) xor (layer0_outputs(3344));
    layer1_outputs(1140) <= not(layer0_outputs(6321)) or (layer0_outputs(4400));
    layer1_outputs(1141) <= (layer0_outputs(1846)) and not (layer0_outputs(2775));
    layer1_outputs(1142) <= not(layer0_outputs(1866));
    layer1_outputs(1143) <= (layer0_outputs(4880)) and not (layer0_outputs(3527));
    layer1_outputs(1144) <= (layer0_outputs(6391)) and (layer0_outputs(1386));
    layer1_outputs(1145) <= not(layer0_outputs(2365)) or (layer0_outputs(5022));
    layer1_outputs(1146) <= not((layer0_outputs(1437)) and (layer0_outputs(7346)));
    layer1_outputs(1147) <= not((layer0_outputs(603)) and (layer0_outputs(5481)));
    layer1_outputs(1148) <= not((layer0_outputs(4772)) xor (layer0_outputs(5801)));
    layer1_outputs(1149) <= not((layer0_outputs(6904)) or (layer0_outputs(6710)));
    layer1_outputs(1150) <= not(layer0_outputs(4740));
    layer1_outputs(1151) <= (layer0_outputs(7471)) or (layer0_outputs(1130));
    layer1_outputs(1152) <= '1';
    layer1_outputs(1153) <= '0';
    layer1_outputs(1154) <= layer0_outputs(3198);
    layer1_outputs(1155) <= (layer0_outputs(2401)) and not (layer0_outputs(6369));
    layer1_outputs(1156) <= (layer0_outputs(3308)) xor (layer0_outputs(1660));
    layer1_outputs(1157) <= not(layer0_outputs(5596)) or (layer0_outputs(1301));
    layer1_outputs(1158) <= not(layer0_outputs(6251));
    layer1_outputs(1159) <= layer0_outputs(4785);
    layer1_outputs(1160) <= (layer0_outputs(7157)) or (layer0_outputs(2908));
    layer1_outputs(1161) <= (layer0_outputs(3520)) xor (layer0_outputs(4241));
    layer1_outputs(1162) <= (layer0_outputs(1912)) and not (layer0_outputs(5450));
    layer1_outputs(1163) <= (layer0_outputs(654)) or (layer0_outputs(294));
    layer1_outputs(1164) <= (layer0_outputs(2442)) and not (layer0_outputs(6306));
    layer1_outputs(1165) <= layer0_outputs(6354);
    layer1_outputs(1166) <= not(layer0_outputs(4794));
    layer1_outputs(1167) <= not(layer0_outputs(6104));
    layer1_outputs(1168) <= (layer0_outputs(5924)) and (layer0_outputs(2854));
    layer1_outputs(1169) <= not(layer0_outputs(2135));
    layer1_outputs(1170) <= layer0_outputs(6544);
    layer1_outputs(1171) <= not(layer0_outputs(3992));
    layer1_outputs(1172) <= '1';
    layer1_outputs(1173) <= (layer0_outputs(4987)) and (layer0_outputs(4257));
    layer1_outputs(1174) <= '0';
    layer1_outputs(1175) <= not(layer0_outputs(2758)) or (layer0_outputs(1475));
    layer1_outputs(1176) <= not((layer0_outputs(2443)) or (layer0_outputs(6267)));
    layer1_outputs(1177) <= (layer0_outputs(1850)) xor (layer0_outputs(4070));
    layer1_outputs(1178) <= not((layer0_outputs(2990)) or (layer0_outputs(3825)));
    layer1_outputs(1179) <= (layer0_outputs(3666)) or (layer0_outputs(2886));
    layer1_outputs(1180) <= (layer0_outputs(4546)) and not (layer0_outputs(1919));
    layer1_outputs(1181) <= (layer0_outputs(105)) and (layer0_outputs(2199));
    layer1_outputs(1182) <= not(layer0_outputs(4981)) or (layer0_outputs(867));
    layer1_outputs(1183) <= (layer0_outputs(6151)) and not (layer0_outputs(6003));
    layer1_outputs(1184) <= not(layer0_outputs(6724)) or (layer0_outputs(622));
    layer1_outputs(1185) <= not(layer0_outputs(3620));
    layer1_outputs(1186) <= (layer0_outputs(1894)) and not (layer0_outputs(1063));
    layer1_outputs(1187) <= (layer0_outputs(7497)) or (layer0_outputs(2903));
    layer1_outputs(1188) <= not(layer0_outputs(5584)) or (layer0_outputs(4546));
    layer1_outputs(1189) <= (layer0_outputs(117)) and not (layer0_outputs(5337));
    layer1_outputs(1190) <= not((layer0_outputs(155)) and (layer0_outputs(2445)));
    layer1_outputs(1191) <= layer0_outputs(6156);
    layer1_outputs(1192) <= layer0_outputs(3876);
    layer1_outputs(1193) <= not((layer0_outputs(3374)) and (layer0_outputs(3448)));
    layer1_outputs(1194) <= not(layer0_outputs(2267));
    layer1_outputs(1195) <= not((layer0_outputs(5898)) or (layer0_outputs(2706)));
    layer1_outputs(1196) <= (layer0_outputs(6693)) and not (layer0_outputs(106));
    layer1_outputs(1197) <= not((layer0_outputs(1401)) or (layer0_outputs(4894)));
    layer1_outputs(1198) <= not(layer0_outputs(5594)) or (layer0_outputs(3914));
    layer1_outputs(1199) <= not(layer0_outputs(2337)) or (layer0_outputs(4816));
    layer1_outputs(1200) <= not(layer0_outputs(6347)) or (layer0_outputs(3608));
    layer1_outputs(1201) <= '1';
    layer1_outputs(1202) <= not((layer0_outputs(881)) and (layer0_outputs(6415)));
    layer1_outputs(1203) <= not(layer0_outputs(5535));
    layer1_outputs(1204) <= not((layer0_outputs(2574)) and (layer0_outputs(7073)));
    layer1_outputs(1205) <= not((layer0_outputs(5039)) and (layer0_outputs(2038)));
    layer1_outputs(1206) <= not(layer0_outputs(2670));
    layer1_outputs(1207) <= not(layer0_outputs(4734)) or (layer0_outputs(428));
    layer1_outputs(1208) <= layer0_outputs(2896);
    layer1_outputs(1209) <= '0';
    layer1_outputs(1210) <= not(layer0_outputs(7625));
    layer1_outputs(1211) <= layer0_outputs(496);
    layer1_outputs(1212) <= not(layer0_outputs(6449)) or (layer0_outputs(6388));
    layer1_outputs(1213) <= layer0_outputs(1636);
    layer1_outputs(1214) <= layer0_outputs(2082);
    layer1_outputs(1215) <= layer0_outputs(2357);
    layer1_outputs(1216) <= not(layer0_outputs(3880));
    layer1_outputs(1217) <= layer0_outputs(5164);
    layer1_outputs(1218) <= not(layer0_outputs(5554));
    layer1_outputs(1219) <= not(layer0_outputs(1029)) or (layer0_outputs(6519));
    layer1_outputs(1220) <= layer0_outputs(655);
    layer1_outputs(1221) <= (layer0_outputs(5317)) and not (layer0_outputs(7651));
    layer1_outputs(1222) <= not(layer0_outputs(6414));
    layer1_outputs(1223) <= layer0_outputs(4287);
    layer1_outputs(1224) <= (layer0_outputs(55)) or (layer0_outputs(1036));
    layer1_outputs(1225) <= (layer0_outputs(6893)) or (layer0_outputs(5119));
    layer1_outputs(1226) <= not((layer0_outputs(6644)) and (layer0_outputs(4691)));
    layer1_outputs(1227) <= not((layer0_outputs(7003)) or (layer0_outputs(2697)));
    layer1_outputs(1228) <= layer0_outputs(1921);
    layer1_outputs(1229) <= (layer0_outputs(1269)) and not (layer0_outputs(4923));
    layer1_outputs(1230) <= not(layer0_outputs(1390)) or (layer0_outputs(823));
    layer1_outputs(1231) <= (layer0_outputs(1592)) and not (layer0_outputs(6946));
    layer1_outputs(1232) <= '0';
    layer1_outputs(1233) <= (layer0_outputs(147)) xor (layer0_outputs(6025));
    layer1_outputs(1234) <= not(layer0_outputs(7464));
    layer1_outputs(1235) <= (layer0_outputs(1432)) and (layer0_outputs(4818));
    layer1_outputs(1236) <= '1';
    layer1_outputs(1237) <= not(layer0_outputs(5788));
    layer1_outputs(1238) <= '0';
    layer1_outputs(1239) <= not((layer0_outputs(5303)) or (layer0_outputs(1916)));
    layer1_outputs(1240) <= not(layer0_outputs(1710));
    layer1_outputs(1241) <= not((layer0_outputs(1735)) and (layer0_outputs(3217)));
    layer1_outputs(1242) <= not((layer0_outputs(2781)) and (layer0_outputs(3931)));
    layer1_outputs(1243) <= not(layer0_outputs(2430)) or (layer0_outputs(4351));
    layer1_outputs(1244) <= not((layer0_outputs(4131)) or (layer0_outputs(1944)));
    layer1_outputs(1245) <= '0';
    layer1_outputs(1246) <= not((layer0_outputs(4339)) and (layer0_outputs(7318)));
    layer1_outputs(1247) <= '1';
    layer1_outputs(1248) <= not(layer0_outputs(5059)) or (layer0_outputs(3122));
    layer1_outputs(1249) <= not(layer0_outputs(4195));
    layer1_outputs(1250) <= layer0_outputs(189);
    layer1_outputs(1251) <= not(layer0_outputs(7269));
    layer1_outputs(1252) <= (layer0_outputs(738)) and (layer0_outputs(3654));
    layer1_outputs(1253) <= not((layer0_outputs(6085)) and (layer0_outputs(6202)));
    layer1_outputs(1254) <= (layer0_outputs(5950)) and (layer0_outputs(5771));
    layer1_outputs(1255) <= not(layer0_outputs(7016));
    layer1_outputs(1256) <= layer0_outputs(2492);
    layer1_outputs(1257) <= layer0_outputs(1493);
    layer1_outputs(1258) <= '1';
    layer1_outputs(1259) <= not(layer0_outputs(3567)) or (layer0_outputs(458));
    layer1_outputs(1260) <= (layer0_outputs(4029)) or (layer0_outputs(238));
    layer1_outputs(1261) <= not((layer0_outputs(323)) or (layer0_outputs(6182)));
    layer1_outputs(1262) <= (layer0_outputs(6603)) and not (layer0_outputs(4885));
    layer1_outputs(1263) <= '0';
    layer1_outputs(1264) <= (layer0_outputs(2986)) and not (layer0_outputs(6304));
    layer1_outputs(1265) <= layer0_outputs(7235);
    layer1_outputs(1266) <= layer0_outputs(5884);
    layer1_outputs(1267) <= not(layer0_outputs(1607));
    layer1_outputs(1268) <= (layer0_outputs(2661)) or (layer0_outputs(5666));
    layer1_outputs(1269) <= '1';
    layer1_outputs(1270) <= not(layer0_outputs(7647));
    layer1_outputs(1271) <= '1';
    layer1_outputs(1272) <= layer0_outputs(3649);
    layer1_outputs(1273) <= not((layer0_outputs(6920)) xor (layer0_outputs(4131)));
    layer1_outputs(1274) <= not(layer0_outputs(5326));
    layer1_outputs(1275) <= not(layer0_outputs(5540));
    layer1_outputs(1276) <= layer0_outputs(3731);
    layer1_outputs(1277) <= '1';
    layer1_outputs(1278) <= (layer0_outputs(4137)) or (layer0_outputs(5763));
    layer1_outputs(1279) <= not((layer0_outputs(2694)) and (layer0_outputs(4553)));
    layer1_outputs(1280) <= (layer0_outputs(846)) and (layer0_outputs(907));
    layer1_outputs(1281) <= not(layer0_outputs(58)) or (layer0_outputs(2135));
    layer1_outputs(1282) <= (layer0_outputs(1122)) and (layer0_outputs(6879));
    layer1_outputs(1283) <= not((layer0_outputs(3858)) and (layer0_outputs(4602)));
    layer1_outputs(1284) <= not(layer0_outputs(3039)) or (layer0_outputs(3999));
    layer1_outputs(1285) <= layer0_outputs(131);
    layer1_outputs(1286) <= not(layer0_outputs(3149));
    layer1_outputs(1287) <= '1';
    layer1_outputs(1288) <= (layer0_outputs(6674)) or (layer0_outputs(2658));
    layer1_outputs(1289) <= not((layer0_outputs(4867)) and (layer0_outputs(2446)));
    layer1_outputs(1290) <= not(layer0_outputs(5159)) or (layer0_outputs(3356));
    layer1_outputs(1291) <= '0';
    layer1_outputs(1292) <= (layer0_outputs(2392)) and not (layer0_outputs(602));
    layer1_outputs(1293) <= not(layer0_outputs(2448));
    layer1_outputs(1294) <= (layer0_outputs(5161)) and not (layer0_outputs(3414));
    layer1_outputs(1295) <= not(layer0_outputs(3115)) or (layer0_outputs(6485));
    layer1_outputs(1296) <= (layer0_outputs(4554)) or (layer0_outputs(4633));
    layer1_outputs(1297) <= layer0_outputs(6258);
    layer1_outputs(1298) <= not(layer0_outputs(7432));
    layer1_outputs(1299) <= not((layer0_outputs(829)) xor (layer0_outputs(7316)));
    layer1_outputs(1300) <= (layer0_outputs(573)) and not (layer0_outputs(7592));
    layer1_outputs(1301) <= layer0_outputs(3546);
    layer1_outputs(1302) <= '0';
    layer1_outputs(1303) <= not(layer0_outputs(46));
    layer1_outputs(1304) <= not(layer0_outputs(4610)) or (layer0_outputs(1675));
    layer1_outputs(1305) <= not(layer0_outputs(2529)) or (layer0_outputs(2885));
    layer1_outputs(1306) <= not((layer0_outputs(782)) or (layer0_outputs(3733)));
    layer1_outputs(1307) <= not(layer0_outputs(7199));
    layer1_outputs(1308) <= (layer0_outputs(6854)) and (layer0_outputs(6297));
    layer1_outputs(1309) <= not((layer0_outputs(3105)) or (layer0_outputs(6881)));
    layer1_outputs(1310) <= layer0_outputs(6135);
    layer1_outputs(1311) <= layer0_outputs(4072);
    layer1_outputs(1312) <= (layer0_outputs(1621)) and not (layer0_outputs(1217));
    layer1_outputs(1313) <= not(layer0_outputs(2281)) or (layer0_outputs(3910));
    layer1_outputs(1314) <= layer0_outputs(6487);
    layer1_outputs(1315) <= layer0_outputs(394);
    layer1_outputs(1316) <= '1';
    layer1_outputs(1317) <= not(layer0_outputs(6365)) or (layer0_outputs(4518));
    layer1_outputs(1318) <= not((layer0_outputs(2808)) and (layer0_outputs(3315)));
    layer1_outputs(1319) <= layer0_outputs(5067);
    layer1_outputs(1320) <= (layer0_outputs(1035)) and not (layer0_outputs(3616));
    layer1_outputs(1321) <= (layer0_outputs(1911)) and not (layer0_outputs(1186));
    layer1_outputs(1322) <= not((layer0_outputs(5296)) xor (layer0_outputs(3153)));
    layer1_outputs(1323) <= not(layer0_outputs(2034));
    layer1_outputs(1324) <= not((layer0_outputs(6712)) or (layer0_outputs(1686)));
    layer1_outputs(1325) <= (layer0_outputs(4210)) and (layer0_outputs(784));
    layer1_outputs(1326) <= (layer0_outputs(6093)) and not (layer0_outputs(2233));
    layer1_outputs(1327) <= not(layer0_outputs(3271));
    layer1_outputs(1328) <= (layer0_outputs(3431)) and (layer0_outputs(3855));
    layer1_outputs(1329) <= (layer0_outputs(6012)) and not (layer0_outputs(1668));
    layer1_outputs(1330) <= not((layer0_outputs(1742)) or (layer0_outputs(3183)));
    layer1_outputs(1331) <= (layer0_outputs(5246)) and not (layer0_outputs(417));
    layer1_outputs(1332) <= '0';
    layer1_outputs(1333) <= (layer0_outputs(6489)) or (layer0_outputs(3098));
    layer1_outputs(1334) <= not(layer0_outputs(3630)) or (layer0_outputs(4574));
    layer1_outputs(1335) <= '0';
    layer1_outputs(1336) <= (layer0_outputs(5825)) and (layer0_outputs(3010));
    layer1_outputs(1337) <= '0';
    layer1_outputs(1338) <= not(layer0_outputs(2268)) or (layer0_outputs(7113));
    layer1_outputs(1339) <= (layer0_outputs(2606)) and (layer0_outputs(4246));
    layer1_outputs(1340) <= layer0_outputs(10);
    layer1_outputs(1341) <= (layer0_outputs(3048)) and not (layer0_outputs(1037));
    layer1_outputs(1342) <= not(layer0_outputs(4655));
    layer1_outputs(1343) <= not(layer0_outputs(3211));
    layer1_outputs(1344) <= not(layer0_outputs(2833));
    layer1_outputs(1345) <= layer0_outputs(7343);
    layer1_outputs(1346) <= not(layer0_outputs(4145));
    layer1_outputs(1347) <= layer0_outputs(1040);
    layer1_outputs(1348) <= (layer0_outputs(4541)) or (layer0_outputs(4095));
    layer1_outputs(1349) <= '0';
    layer1_outputs(1350) <= not(layer0_outputs(4534));
    layer1_outputs(1351) <= not(layer0_outputs(2800));
    layer1_outputs(1352) <= not(layer0_outputs(1206)) or (layer0_outputs(2996));
    layer1_outputs(1353) <= (layer0_outputs(701)) and not (layer0_outputs(4720));
    layer1_outputs(1354) <= not(layer0_outputs(6571)) or (layer0_outputs(5812));
    layer1_outputs(1355) <= not(layer0_outputs(5587)) or (layer0_outputs(3505));
    layer1_outputs(1356) <= (layer0_outputs(534)) and (layer0_outputs(6365));
    layer1_outputs(1357) <= not(layer0_outputs(6851));
    layer1_outputs(1358) <= not(layer0_outputs(880)) or (layer0_outputs(7425));
    layer1_outputs(1359) <= not(layer0_outputs(4843));
    layer1_outputs(1360) <= not(layer0_outputs(5250)) or (layer0_outputs(5113));
    layer1_outputs(1361) <= (layer0_outputs(7402)) xor (layer0_outputs(3389));
    layer1_outputs(1362) <= (layer0_outputs(7277)) xor (layer0_outputs(2344));
    layer1_outputs(1363) <= not(layer0_outputs(3976));
    layer1_outputs(1364) <= not((layer0_outputs(3967)) and (layer0_outputs(3848)));
    layer1_outputs(1365) <= not(layer0_outputs(4608)) or (layer0_outputs(2322));
    layer1_outputs(1366) <= (layer0_outputs(775)) or (layer0_outputs(1384));
    layer1_outputs(1367) <= layer0_outputs(7518);
    layer1_outputs(1368) <= (layer0_outputs(7114)) or (layer0_outputs(1207));
    layer1_outputs(1369) <= not((layer0_outputs(6337)) and (layer0_outputs(6560)));
    layer1_outputs(1370) <= not(layer0_outputs(3745));
    layer1_outputs(1371) <= (layer0_outputs(1617)) and not (layer0_outputs(1501));
    layer1_outputs(1372) <= not((layer0_outputs(6860)) and (layer0_outputs(7270)));
    layer1_outputs(1373) <= not(layer0_outputs(7130));
    layer1_outputs(1374) <= not(layer0_outputs(3880));
    layer1_outputs(1375) <= (layer0_outputs(20)) and not (layer0_outputs(5104));
    layer1_outputs(1376) <= '0';
    layer1_outputs(1377) <= not(layer0_outputs(833)) or (layer0_outputs(4417));
    layer1_outputs(1378) <= layer0_outputs(2037);
    layer1_outputs(1379) <= not(layer0_outputs(2705));
    layer1_outputs(1380) <= (layer0_outputs(1985)) and not (layer0_outputs(6855));
    layer1_outputs(1381) <= not(layer0_outputs(5081));
    layer1_outputs(1382) <= not(layer0_outputs(1358));
    layer1_outputs(1383) <= '1';
    layer1_outputs(1384) <= not((layer0_outputs(7492)) and (layer0_outputs(3742)));
    layer1_outputs(1385) <= (layer0_outputs(3981)) or (layer0_outputs(2954));
    layer1_outputs(1386) <= (layer0_outputs(2590)) and not (layer0_outputs(7035));
    layer1_outputs(1387) <= '0';
    layer1_outputs(1388) <= not(layer0_outputs(6014));
    layer1_outputs(1389) <= layer0_outputs(2672);
    layer1_outputs(1390) <= (layer0_outputs(1631)) and not (layer0_outputs(3470));
    layer1_outputs(1391) <= (layer0_outputs(1118)) and not (layer0_outputs(5821));
    layer1_outputs(1392) <= (layer0_outputs(6026)) or (layer0_outputs(4251));
    layer1_outputs(1393) <= layer0_outputs(2181);
    layer1_outputs(1394) <= not((layer0_outputs(6790)) or (layer0_outputs(288)));
    layer1_outputs(1395) <= not((layer0_outputs(3046)) or (layer0_outputs(5509)));
    layer1_outputs(1396) <= (layer0_outputs(7224)) or (layer0_outputs(235));
    layer1_outputs(1397) <= (layer0_outputs(4064)) and (layer0_outputs(5219));
    layer1_outputs(1398) <= not(layer0_outputs(3839)) or (layer0_outputs(5335));
    layer1_outputs(1399) <= (layer0_outputs(2414)) and not (layer0_outputs(586));
    layer1_outputs(1400) <= layer0_outputs(911);
    layer1_outputs(1401) <= '0';
    layer1_outputs(1402) <= not((layer0_outputs(701)) xor (layer0_outputs(1082)));
    layer1_outputs(1403) <= not(layer0_outputs(5872)) or (layer0_outputs(6394));
    layer1_outputs(1404) <= not((layer0_outputs(383)) or (layer0_outputs(4369)));
    layer1_outputs(1405) <= not((layer0_outputs(2839)) or (layer0_outputs(3996)));
    layer1_outputs(1406) <= not(layer0_outputs(1150));
    layer1_outputs(1407) <= not(layer0_outputs(3892)) or (layer0_outputs(367));
    layer1_outputs(1408) <= layer0_outputs(1936);
    layer1_outputs(1409) <= (layer0_outputs(5507)) and not (layer0_outputs(7295));
    layer1_outputs(1410) <= layer0_outputs(1263);
    layer1_outputs(1411) <= not(layer0_outputs(4205));
    layer1_outputs(1412) <= not(layer0_outputs(3685));
    layer1_outputs(1413) <= (layer0_outputs(5865)) and not (layer0_outputs(5404));
    layer1_outputs(1414) <= not((layer0_outputs(7440)) or (layer0_outputs(5490)));
    layer1_outputs(1415) <= not((layer0_outputs(1099)) and (layer0_outputs(3224)));
    layer1_outputs(1416) <= '1';
    layer1_outputs(1417) <= not(layer0_outputs(5168)) or (layer0_outputs(4902));
    layer1_outputs(1418) <= layer0_outputs(6007);
    layer1_outputs(1419) <= (layer0_outputs(7056)) or (layer0_outputs(3264));
    layer1_outputs(1420) <= not((layer0_outputs(3534)) and (layer0_outputs(6524)));
    layer1_outputs(1421) <= not(layer0_outputs(337)) or (layer0_outputs(5381));
    layer1_outputs(1422) <= (layer0_outputs(2559)) and not (layer0_outputs(704));
    layer1_outputs(1423) <= (layer0_outputs(4757)) and not (layer0_outputs(7381));
    layer1_outputs(1424) <= not((layer0_outputs(6400)) and (layer0_outputs(2408)));
    layer1_outputs(1425) <= layer0_outputs(3671);
    layer1_outputs(1426) <= not((layer0_outputs(1755)) and (layer0_outputs(5606)));
    layer1_outputs(1427) <= layer0_outputs(2685);
    layer1_outputs(1428) <= layer0_outputs(5982);
    layer1_outputs(1429) <= '1';
    layer1_outputs(1430) <= not(layer0_outputs(5809));
    layer1_outputs(1431) <= (layer0_outputs(7261)) or (layer0_outputs(2665));
    layer1_outputs(1432) <= (layer0_outputs(6301)) and not (layer0_outputs(3526));
    layer1_outputs(1433) <= not(layer0_outputs(2416));
    layer1_outputs(1434) <= not((layer0_outputs(5472)) xor (layer0_outputs(1298)));
    layer1_outputs(1435) <= layer0_outputs(6700);
    layer1_outputs(1436) <= (layer0_outputs(5845)) or (layer0_outputs(7519));
    layer1_outputs(1437) <= layer0_outputs(4836);
    layer1_outputs(1438) <= layer0_outputs(4592);
    layer1_outputs(1439) <= (layer0_outputs(3102)) or (layer0_outputs(4143));
    layer1_outputs(1440) <= layer0_outputs(2466);
    layer1_outputs(1441) <= not((layer0_outputs(2392)) and (layer0_outputs(5159)));
    layer1_outputs(1442) <= layer0_outputs(4595);
    layer1_outputs(1443) <= not((layer0_outputs(4068)) and (layer0_outputs(237)));
    layer1_outputs(1444) <= layer0_outputs(7373);
    layer1_outputs(1445) <= (layer0_outputs(4456)) and not (layer0_outputs(132));
    layer1_outputs(1446) <= (layer0_outputs(4037)) and (layer0_outputs(6765));
    layer1_outputs(1447) <= '1';
    layer1_outputs(1448) <= not(layer0_outputs(3611)) or (layer0_outputs(5949));
    layer1_outputs(1449) <= (layer0_outputs(621)) xor (layer0_outputs(5078));
    layer1_outputs(1450) <= layer0_outputs(3324);
    layer1_outputs(1451) <= not((layer0_outputs(1511)) and (layer0_outputs(4421)));
    layer1_outputs(1452) <= not(layer0_outputs(373)) or (layer0_outputs(666));
    layer1_outputs(1453) <= not(layer0_outputs(5777)) or (layer0_outputs(1077));
    layer1_outputs(1454) <= not(layer0_outputs(4590)) or (layer0_outputs(955));
    layer1_outputs(1455) <= '1';
    layer1_outputs(1456) <= (layer0_outputs(1111)) or (layer0_outputs(5288));
    layer1_outputs(1457) <= layer0_outputs(3587);
    layer1_outputs(1458) <= layer0_outputs(2507);
    layer1_outputs(1459) <= not(layer0_outputs(4235)) or (layer0_outputs(6701));
    layer1_outputs(1460) <= not(layer0_outputs(2842)) or (layer0_outputs(3595));
    layer1_outputs(1461) <= not(layer0_outputs(2522)) or (layer0_outputs(4562));
    layer1_outputs(1462) <= (layer0_outputs(5763)) or (layer0_outputs(5936));
    layer1_outputs(1463) <= '0';
    layer1_outputs(1464) <= not(layer0_outputs(5983));
    layer1_outputs(1465) <= '1';
    layer1_outputs(1466) <= layer0_outputs(2742);
    layer1_outputs(1467) <= not(layer0_outputs(6839)) or (layer0_outputs(5653));
    layer1_outputs(1468) <= not((layer0_outputs(3416)) or (layer0_outputs(2365)));
    layer1_outputs(1469) <= '1';
    layer1_outputs(1470) <= '1';
    layer1_outputs(1471) <= not((layer0_outputs(2844)) or (layer0_outputs(571)));
    layer1_outputs(1472) <= not(layer0_outputs(5598));
    layer1_outputs(1473) <= not(layer0_outputs(2591)) or (layer0_outputs(6559));
    layer1_outputs(1474) <= not(layer0_outputs(5845)) or (layer0_outputs(6611));
    layer1_outputs(1475) <= not(layer0_outputs(5534));
    layer1_outputs(1476) <= '1';
    layer1_outputs(1477) <= (layer0_outputs(888)) and not (layer0_outputs(2849));
    layer1_outputs(1478) <= (layer0_outputs(4176)) and not (layer0_outputs(4377));
    layer1_outputs(1479) <= not(layer0_outputs(176));
    layer1_outputs(1480) <= not(layer0_outputs(2836));
    layer1_outputs(1481) <= (layer0_outputs(3615)) and not (layer0_outputs(7260));
    layer1_outputs(1482) <= (layer0_outputs(6702)) and (layer0_outputs(7616));
    layer1_outputs(1483) <= not((layer0_outputs(5294)) xor (layer0_outputs(5213)));
    layer1_outputs(1484) <= not(layer0_outputs(6135));
    layer1_outputs(1485) <= not((layer0_outputs(2956)) and (layer0_outputs(6110)));
    layer1_outputs(1486) <= (layer0_outputs(7675)) and not (layer0_outputs(1261));
    layer1_outputs(1487) <= '0';
    layer1_outputs(1488) <= (layer0_outputs(6196)) or (layer0_outputs(7074));
    layer1_outputs(1489) <= (layer0_outputs(5463)) and (layer0_outputs(5066));
    layer1_outputs(1490) <= not(layer0_outputs(3445));
    layer1_outputs(1491) <= (layer0_outputs(4206)) and not (layer0_outputs(5423));
    layer1_outputs(1492) <= (layer0_outputs(1402)) and not (layer0_outputs(2730));
    layer1_outputs(1493) <= layer0_outputs(6901);
    layer1_outputs(1494) <= (layer0_outputs(2514)) and not (layer0_outputs(5070));
    layer1_outputs(1495) <= (layer0_outputs(4974)) and not (layer0_outputs(4838));
    layer1_outputs(1496) <= (layer0_outputs(2031)) and not (layer0_outputs(6129));
    layer1_outputs(1497) <= (layer0_outputs(5657)) and not (layer0_outputs(2367));
    layer1_outputs(1498) <= not(layer0_outputs(3536));
    layer1_outputs(1499) <= not(layer0_outputs(6945));
    layer1_outputs(1500) <= not(layer0_outputs(385)) or (layer0_outputs(2874));
    layer1_outputs(1501) <= layer0_outputs(1639);
    layer1_outputs(1502) <= layer0_outputs(7384);
    layer1_outputs(1503) <= not((layer0_outputs(1795)) and (layer0_outputs(3368)));
    layer1_outputs(1504) <= not((layer0_outputs(4594)) xor (layer0_outputs(6460)));
    layer1_outputs(1505) <= '0';
    layer1_outputs(1506) <= (layer0_outputs(7668)) and not (layer0_outputs(413));
    layer1_outputs(1507) <= not(layer0_outputs(6980)) or (layer0_outputs(5581));
    layer1_outputs(1508) <= layer0_outputs(3617);
    layer1_outputs(1509) <= layer0_outputs(1532);
    layer1_outputs(1510) <= not(layer0_outputs(3991));
    layer1_outputs(1511) <= not(layer0_outputs(3444));
    layer1_outputs(1512) <= (layer0_outputs(3294)) and not (layer0_outputs(1473));
    layer1_outputs(1513) <= '0';
    layer1_outputs(1514) <= (layer0_outputs(4642)) and not (layer0_outputs(1457));
    layer1_outputs(1515) <= not(layer0_outputs(3550)) or (layer0_outputs(2261));
    layer1_outputs(1516) <= not(layer0_outputs(1633));
    layer1_outputs(1517) <= (layer0_outputs(1334)) and not (layer0_outputs(981));
    layer1_outputs(1518) <= not((layer0_outputs(6096)) and (layer0_outputs(5539)));
    layer1_outputs(1519) <= '1';
    layer1_outputs(1520) <= '1';
    layer1_outputs(1521) <= not(layer0_outputs(5087));
    layer1_outputs(1522) <= not(layer0_outputs(2882));
    layer1_outputs(1523) <= not(layer0_outputs(4010)) or (layer0_outputs(2729));
    layer1_outputs(1524) <= layer0_outputs(956);
    layer1_outputs(1525) <= not(layer0_outputs(765));
    layer1_outputs(1526) <= not((layer0_outputs(3589)) and (layer0_outputs(398)));
    layer1_outputs(1527) <= not((layer0_outputs(7382)) and (layer0_outputs(3683)));
    layer1_outputs(1528) <= not(layer0_outputs(7049)) or (layer0_outputs(6284));
    layer1_outputs(1529) <= (layer0_outputs(1196)) and not (layer0_outputs(6180));
    layer1_outputs(1530) <= '0';
    layer1_outputs(1531) <= layer0_outputs(4803);
    layer1_outputs(1532) <= (layer0_outputs(3060)) and not (layer0_outputs(4798));
    layer1_outputs(1533) <= not(layer0_outputs(6226));
    layer1_outputs(1534) <= not(layer0_outputs(7261));
    layer1_outputs(1535) <= not((layer0_outputs(4852)) and (layer0_outputs(5536)));
    layer1_outputs(1536) <= not((layer0_outputs(142)) and (layer0_outputs(4867)));
    layer1_outputs(1537) <= not(layer0_outputs(1510));
    layer1_outputs(1538) <= not((layer0_outputs(3543)) and (layer0_outputs(5169)));
    layer1_outputs(1539) <= not((layer0_outputs(5471)) or (layer0_outputs(7219)));
    layer1_outputs(1540) <= not(layer0_outputs(1999));
    layer1_outputs(1541) <= not(layer0_outputs(3826)) or (layer0_outputs(5735));
    layer1_outputs(1542) <= (layer0_outputs(6883)) and not (layer0_outputs(2713));
    layer1_outputs(1543) <= (layer0_outputs(4165)) xor (layer0_outputs(6917));
    layer1_outputs(1544) <= layer0_outputs(5881);
    layer1_outputs(1545) <= not(layer0_outputs(511));
    layer1_outputs(1546) <= (layer0_outputs(3112)) and not (layer0_outputs(34));
    layer1_outputs(1547) <= not(layer0_outputs(2900));
    layer1_outputs(1548) <= not(layer0_outputs(1591));
    layer1_outputs(1549) <= (layer0_outputs(1748)) or (layer0_outputs(3461));
    layer1_outputs(1550) <= not(layer0_outputs(2243)) or (layer0_outputs(4622));
    layer1_outputs(1551) <= (layer0_outputs(934)) or (layer0_outputs(2091));
    layer1_outputs(1552) <= (layer0_outputs(5241)) and not (layer0_outputs(6203));
    layer1_outputs(1553) <= (layer0_outputs(2797)) and not (layer0_outputs(348));
    layer1_outputs(1554) <= (layer0_outputs(5908)) and not (layer0_outputs(4659));
    layer1_outputs(1555) <= not(layer0_outputs(3514));
    layer1_outputs(1556) <= not(layer0_outputs(7433));
    layer1_outputs(1557) <= not(layer0_outputs(1101)) or (layer0_outputs(1838));
    layer1_outputs(1558) <= not(layer0_outputs(3848));
    layer1_outputs(1559) <= (layer0_outputs(5287)) and not (layer0_outputs(6415));
    layer1_outputs(1560) <= (layer0_outputs(5773)) and not (layer0_outputs(2569));
    layer1_outputs(1561) <= not((layer0_outputs(4278)) and (layer0_outputs(3541)));
    layer1_outputs(1562) <= (layer0_outputs(5126)) or (layer0_outputs(4265));
    layer1_outputs(1563) <= (layer0_outputs(3293)) and not (layer0_outputs(4189));
    layer1_outputs(1564) <= '1';
    layer1_outputs(1565) <= layer0_outputs(2262);
    layer1_outputs(1566) <= (layer0_outputs(6368)) or (layer0_outputs(6650));
    layer1_outputs(1567) <= layer0_outputs(5652);
    layer1_outputs(1568) <= not(layer0_outputs(4379));
    layer1_outputs(1569) <= (layer0_outputs(3338)) and not (layer0_outputs(4216));
    layer1_outputs(1570) <= (layer0_outputs(7421)) and (layer0_outputs(1922));
    layer1_outputs(1571) <= not(layer0_outputs(4264)) or (layer0_outputs(6528));
    layer1_outputs(1572) <= layer0_outputs(4260);
    layer1_outputs(1573) <= (layer0_outputs(756)) and not (layer0_outputs(6081));
    layer1_outputs(1574) <= not(layer0_outputs(3108)) or (layer0_outputs(4873));
    layer1_outputs(1575) <= not(layer0_outputs(3804)) or (layer0_outputs(6597));
    layer1_outputs(1576) <= layer0_outputs(4632);
    layer1_outputs(1577) <= layer0_outputs(1272);
    layer1_outputs(1578) <= '1';
    layer1_outputs(1579) <= '0';
    layer1_outputs(1580) <= '0';
    layer1_outputs(1581) <= layer0_outputs(5039);
    layer1_outputs(1582) <= not(layer0_outputs(2390));
    layer1_outputs(1583) <= (layer0_outputs(4909)) and (layer0_outputs(2404));
    layer1_outputs(1584) <= not(layer0_outputs(3608));
    layer1_outputs(1585) <= layer0_outputs(6385);
    layer1_outputs(1586) <= layer0_outputs(4599);
    layer1_outputs(1587) <= '1';
    layer1_outputs(1588) <= not(layer0_outputs(5020));
    layer1_outputs(1589) <= layer0_outputs(6452);
    layer1_outputs(1590) <= '1';
    layer1_outputs(1591) <= not(layer0_outputs(4405));
    layer1_outputs(1592) <= not(layer0_outputs(728)) or (layer0_outputs(2069));
    layer1_outputs(1593) <= not(layer0_outputs(1498));
    layer1_outputs(1594) <= (layer0_outputs(4357)) xor (layer0_outputs(938));
    layer1_outputs(1595) <= (layer0_outputs(1114)) or (layer0_outputs(4882));
    layer1_outputs(1596) <= layer0_outputs(7286);
    layer1_outputs(1597) <= '1';
    layer1_outputs(1598) <= '0';
    layer1_outputs(1599) <= (layer0_outputs(1046)) or (layer0_outputs(7283));
    layer1_outputs(1600) <= (layer0_outputs(5256)) or (layer0_outputs(3680));
    layer1_outputs(1601) <= (layer0_outputs(3346)) and not (layer0_outputs(229));
    layer1_outputs(1602) <= (layer0_outputs(678)) and (layer0_outputs(4038));
    layer1_outputs(1603) <= not(layer0_outputs(3079)) or (layer0_outputs(6912));
    layer1_outputs(1604) <= not((layer0_outputs(3655)) or (layer0_outputs(788)));
    layer1_outputs(1605) <= not(layer0_outputs(137));
    layer1_outputs(1606) <= layer0_outputs(171);
    layer1_outputs(1607) <= not(layer0_outputs(6439));
    layer1_outputs(1608) <= (layer0_outputs(6015)) and not (layer0_outputs(4565));
    layer1_outputs(1609) <= not(layer0_outputs(2509));
    layer1_outputs(1610) <= layer0_outputs(7005);
    layer1_outputs(1611) <= not((layer0_outputs(2820)) and (layer0_outputs(5851)));
    layer1_outputs(1612) <= (layer0_outputs(3123)) and not (layer0_outputs(6640));
    layer1_outputs(1613) <= (layer0_outputs(2894)) xor (layer0_outputs(6532));
    layer1_outputs(1614) <= not((layer0_outputs(5511)) and (layer0_outputs(5441)));
    layer1_outputs(1615) <= not((layer0_outputs(5976)) and (layer0_outputs(3870)));
    layer1_outputs(1616) <= not(layer0_outputs(5687));
    layer1_outputs(1617) <= (layer0_outputs(3204)) and not (layer0_outputs(6364));
    layer1_outputs(1618) <= not((layer0_outputs(3218)) or (layer0_outputs(5687)));
    layer1_outputs(1619) <= (layer0_outputs(1629)) and (layer0_outputs(7478));
    layer1_outputs(1620) <= not(layer0_outputs(4949)) or (layer0_outputs(3247));
    layer1_outputs(1621) <= layer0_outputs(2062);
    layer1_outputs(1622) <= not((layer0_outputs(1314)) and (layer0_outputs(5731)));
    layer1_outputs(1623) <= (layer0_outputs(6978)) and not (layer0_outputs(5993));
    layer1_outputs(1624) <= (layer0_outputs(7140)) and not (layer0_outputs(7385));
    layer1_outputs(1625) <= not(layer0_outputs(6346));
    layer1_outputs(1626) <= (layer0_outputs(6212)) and not (layer0_outputs(6919));
    layer1_outputs(1627) <= not(layer0_outputs(3401)) or (layer0_outputs(3990));
    layer1_outputs(1628) <= not((layer0_outputs(4791)) and (layer0_outputs(1109)));
    layer1_outputs(1629) <= not((layer0_outputs(1355)) or (layer0_outputs(6289)));
    layer1_outputs(1630) <= not(layer0_outputs(6918)) or (layer0_outputs(7127));
    layer1_outputs(1631) <= (layer0_outputs(726)) or (layer0_outputs(3129));
    layer1_outputs(1632) <= not(layer0_outputs(381));
    layer1_outputs(1633) <= not((layer0_outputs(6809)) or (layer0_outputs(1429)));
    layer1_outputs(1634) <= not((layer0_outputs(5099)) or (layer0_outputs(4371)));
    layer1_outputs(1635) <= layer0_outputs(4818);
    layer1_outputs(1636) <= (layer0_outputs(7302)) and (layer0_outputs(7082));
    layer1_outputs(1637) <= layer0_outputs(2941);
    layer1_outputs(1638) <= not(layer0_outputs(4951));
    layer1_outputs(1639) <= not(layer0_outputs(6658));
    layer1_outputs(1640) <= (layer0_outputs(1134)) and not (layer0_outputs(3358));
    layer1_outputs(1641) <= (layer0_outputs(4314)) and (layer0_outputs(7460));
    layer1_outputs(1642) <= '1';
    layer1_outputs(1643) <= layer0_outputs(1045);
    layer1_outputs(1644) <= not(layer0_outputs(6961)) or (layer0_outputs(1201));
    layer1_outputs(1645) <= (layer0_outputs(5991)) or (layer0_outputs(5285));
    layer1_outputs(1646) <= layer0_outputs(3053);
    layer1_outputs(1647) <= layer0_outputs(470);
    layer1_outputs(1648) <= (layer0_outputs(6501)) and not (layer0_outputs(7370));
    layer1_outputs(1649) <= layer0_outputs(6595);
    layer1_outputs(1650) <= (layer0_outputs(6300)) and not (layer0_outputs(5717));
    layer1_outputs(1651) <= '0';
    layer1_outputs(1652) <= layer0_outputs(5082);
    layer1_outputs(1653) <= (layer0_outputs(4281)) and not (layer0_outputs(7407));
    layer1_outputs(1654) <= (layer0_outputs(3268)) and (layer0_outputs(1421));
    layer1_outputs(1655) <= not((layer0_outputs(2767)) and (layer0_outputs(2710)));
    layer1_outputs(1656) <= not((layer0_outputs(4361)) and (layer0_outputs(4512)));
    layer1_outputs(1657) <= not(layer0_outputs(1974));
    layer1_outputs(1658) <= (layer0_outputs(2822)) or (layer0_outputs(5770));
    layer1_outputs(1659) <= (layer0_outputs(5364)) or (layer0_outputs(7181));
    layer1_outputs(1660) <= not(layer0_outputs(1221));
    layer1_outputs(1661) <= '0';
    layer1_outputs(1662) <= layer0_outputs(4968);
    layer1_outputs(1663) <= not((layer0_outputs(2273)) or (layer0_outputs(3990)));
    layer1_outputs(1664) <= not(layer0_outputs(3565));
    layer1_outputs(1665) <= (layer0_outputs(1131)) xor (layer0_outputs(484));
    layer1_outputs(1666) <= (layer0_outputs(2203)) and not (layer0_outputs(5443));
    layer1_outputs(1667) <= not(layer0_outputs(1821)) or (layer0_outputs(5210));
    layer1_outputs(1668) <= (layer0_outputs(1462)) and (layer0_outputs(1368));
    layer1_outputs(1669) <= layer0_outputs(1853);
    layer1_outputs(1670) <= not((layer0_outputs(7591)) and (layer0_outputs(4844)));
    layer1_outputs(1671) <= (layer0_outputs(2720)) and not (layer0_outputs(5758));
    layer1_outputs(1672) <= not((layer0_outputs(5538)) or (layer0_outputs(2360)));
    layer1_outputs(1673) <= layer0_outputs(2749);
    layer1_outputs(1674) <= (layer0_outputs(507)) or (layer0_outputs(3337));
    layer1_outputs(1675) <= layer0_outputs(7062);
    layer1_outputs(1676) <= not(layer0_outputs(3084)) or (layer0_outputs(694));
    layer1_outputs(1677) <= not(layer0_outputs(5229));
    layer1_outputs(1678) <= layer0_outputs(2120);
    layer1_outputs(1679) <= layer0_outputs(2972);
    layer1_outputs(1680) <= not(layer0_outputs(3054));
    layer1_outputs(1681) <= not((layer0_outputs(2852)) xor (layer0_outputs(6070)));
    layer1_outputs(1682) <= layer0_outputs(6506);
    layer1_outputs(1683) <= not(layer0_outputs(4088));
    layer1_outputs(1684) <= layer0_outputs(7497);
    layer1_outputs(1685) <= not((layer0_outputs(1031)) and (layer0_outputs(4563)));
    layer1_outputs(1686) <= not((layer0_outputs(7105)) or (layer0_outputs(5123)));
    layer1_outputs(1687) <= layer0_outputs(2263);
    layer1_outputs(1688) <= layer0_outputs(1695);
    layer1_outputs(1689) <= not(layer0_outputs(1909));
    layer1_outputs(1690) <= not(layer0_outputs(489)) or (layer0_outputs(702));
    layer1_outputs(1691) <= not((layer0_outputs(3284)) xor (layer0_outputs(6392)));
    layer1_outputs(1692) <= not(layer0_outputs(2080));
    layer1_outputs(1693) <= not((layer0_outputs(3404)) or (layer0_outputs(4049)));
    layer1_outputs(1694) <= '0';
    layer1_outputs(1695) <= (layer0_outputs(2972)) and not (layer0_outputs(2238));
    layer1_outputs(1696) <= (layer0_outputs(7139)) and (layer0_outputs(1961));
    layer1_outputs(1697) <= layer0_outputs(5354);
    layer1_outputs(1698) <= (layer0_outputs(3034)) and not (layer0_outputs(3769));
    layer1_outputs(1699) <= (layer0_outputs(122)) or (layer0_outputs(4557));
    layer1_outputs(1700) <= '0';
    layer1_outputs(1701) <= (layer0_outputs(4928)) xor (layer0_outputs(5744));
    layer1_outputs(1702) <= (layer0_outputs(6235)) and (layer0_outputs(402));
    layer1_outputs(1703) <= not(layer0_outputs(6887));
    layer1_outputs(1704) <= not((layer0_outputs(4112)) and (layer0_outputs(6570)));
    layer1_outputs(1705) <= not(layer0_outputs(7658)) or (layer0_outputs(5501));
    layer1_outputs(1706) <= not((layer0_outputs(3355)) or (layer0_outputs(4425)));
    layer1_outputs(1707) <= layer0_outputs(2219);
    layer1_outputs(1708) <= not(layer0_outputs(6352));
    layer1_outputs(1709) <= '0';
    layer1_outputs(1710) <= (layer0_outputs(6419)) and not (layer0_outputs(7149));
    layer1_outputs(1711) <= not(layer0_outputs(4784));
    layer1_outputs(1712) <= '0';
    layer1_outputs(1713) <= not(layer0_outputs(125));
    layer1_outputs(1714) <= (layer0_outputs(6729)) or (layer0_outputs(7267));
    layer1_outputs(1715) <= not((layer0_outputs(3933)) and (layer0_outputs(2172)));
    layer1_outputs(1716) <= '1';
    layer1_outputs(1717) <= not(layer0_outputs(7205)) or (layer0_outputs(4129));
    layer1_outputs(1718) <= not(layer0_outputs(4529)) or (layer0_outputs(2472));
    layer1_outputs(1719) <= not((layer0_outputs(2379)) or (layer0_outputs(1151)));
    layer1_outputs(1720) <= not(layer0_outputs(148));
    layer1_outputs(1721) <= not((layer0_outputs(5835)) or (layer0_outputs(2163)));
    layer1_outputs(1722) <= not(layer0_outputs(2873)) or (layer0_outputs(7105));
    layer1_outputs(1723) <= not(layer0_outputs(7532));
    layer1_outputs(1724) <= not(layer0_outputs(465));
    layer1_outputs(1725) <= not(layer0_outputs(2883)) or (layer0_outputs(6609));
    layer1_outputs(1726) <= not((layer0_outputs(709)) and (layer0_outputs(2543)));
    layer1_outputs(1727) <= not(layer0_outputs(3948)) or (layer0_outputs(5330));
    layer1_outputs(1728) <= not(layer0_outputs(577));
    layer1_outputs(1729) <= (layer0_outputs(174)) and (layer0_outputs(195));
    layer1_outputs(1730) <= not(layer0_outputs(1965));
    layer1_outputs(1731) <= (layer0_outputs(1969)) and not (layer0_outputs(6854));
    layer1_outputs(1732) <= (layer0_outputs(6652)) and not (layer0_outputs(6246));
    layer1_outputs(1733) <= not((layer0_outputs(5670)) and (layer0_outputs(6423)));
    layer1_outputs(1734) <= not((layer0_outputs(5992)) and (layer0_outputs(28)));
    layer1_outputs(1735) <= (layer0_outputs(3148)) and not (layer0_outputs(3471));
    layer1_outputs(1736) <= '0';
    layer1_outputs(1737) <= (layer0_outputs(5831)) and not (layer0_outputs(6870));
    layer1_outputs(1738) <= (layer0_outputs(3048)) and not (layer0_outputs(4090));
    layer1_outputs(1739) <= not((layer0_outputs(143)) and (layer0_outputs(5230)));
    layer1_outputs(1740) <= (layer0_outputs(1692)) or (layer0_outputs(2745));
    layer1_outputs(1741) <= (layer0_outputs(2131)) or (layer0_outputs(3924));
    layer1_outputs(1742) <= (layer0_outputs(6126)) and not (layer0_outputs(2502));
    layer1_outputs(1743) <= not(layer0_outputs(4347)) or (layer0_outputs(6441));
    layer1_outputs(1744) <= layer0_outputs(6294);
    layer1_outputs(1745) <= not(layer0_outputs(5036));
    layer1_outputs(1746) <= not(layer0_outputs(990));
    layer1_outputs(1747) <= layer0_outputs(2269);
    layer1_outputs(1748) <= not(layer0_outputs(6026));
    layer1_outputs(1749) <= (layer0_outputs(6467)) or (layer0_outputs(871));
    layer1_outputs(1750) <= not(layer0_outputs(4012)) or (layer0_outputs(2528));
    layer1_outputs(1751) <= (layer0_outputs(6256)) and (layer0_outputs(7159));
    layer1_outputs(1752) <= (layer0_outputs(5862)) and not (layer0_outputs(7330));
    layer1_outputs(1753) <= (layer0_outputs(7169)) and (layer0_outputs(6132));
    layer1_outputs(1754) <= not(layer0_outputs(2728));
    layer1_outputs(1755) <= not(layer0_outputs(3519)) or (layer0_outputs(1901));
    layer1_outputs(1756) <= '1';
    layer1_outputs(1757) <= not((layer0_outputs(4986)) or (layer0_outputs(1902)));
    layer1_outputs(1758) <= not(layer0_outputs(2312)) or (layer0_outputs(6512));
    layer1_outputs(1759) <= (layer0_outputs(6686)) xor (layer0_outputs(1789));
    layer1_outputs(1760) <= not(layer0_outputs(897));
    layer1_outputs(1761) <= '1';
    layer1_outputs(1762) <= not(layer0_outputs(2703));
    layer1_outputs(1763) <= '1';
    layer1_outputs(1764) <= not((layer0_outputs(3124)) or (layer0_outputs(6763)));
    layer1_outputs(1765) <= not((layer0_outputs(2572)) or (layer0_outputs(4192)));
    layer1_outputs(1766) <= (layer0_outputs(3793)) or (layer0_outputs(4913));
    layer1_outputs(1767) <= not(layer0_outputs(2212)) or (layer0_outputs(2568));
    layer1_outputs(1768) <= not(layer0_outputs(613));
    layer1_outputs(1769) <= layer0_outputs(6896);
    layer1_outputs(1770) <= (layer0_outputs(5733)) xor (layer0_outputs(3582));
    layer1_outputs(1771) <= not(layer0_outputs(2996)) or (layer0_outputs(6518));
    layer1_outputs(1772) <= layer0_outputs(6968);
    layer1_outputs(1773) <= not((layer0_outputs(6573)) and (layer0_outputs(5802)));
    layer1_outputs(1774) <= (layer0_outputs(1451)) and not (layer0_outputs(2731));
    layer1_outputs(1775) <= not(layer0_outputs(6583));
    layer1_outputs(1776) <= not((layer0_outputs(1580)) xor (layer0_outputs(3665)));
    layer1_outputs(1777) <= not(layer0_outputs(2099));
    layer1_outputs(1778) <= not(layer0_outputs(1479));
    layer1_outputs(1779) <= not(layer0_outputs(6755));
    layer1_outputs(1780) <= (layer0_outputs(5679)) and (layer0_outputs(4723));
    layer1_outputs(1781) <= not(layer0_outputs(186));
    layer1_outputs(1782) <= not((layer0_outputs(1597)) xor (layer0_outputs(4431)));
    layer1_outputs(1783) <= not(layer0_outputs(2072)) or (layer0_outputs(2156));
    layer1_outputs(1784) <= layer0_outputs(543);
    layer1_outputs(1785) <= not((layer0_outputs(7273)) or (layer0_outputs(7409)));
    layer1_outputs(1786) <= not((layer0_outputs(3814)) or (layer0_outputs(1919)));
    layer1_outputs(1787) <= layer0_outputs(5456);
    layer1_outputs(1788) <= (layer0_outputs(2106)) and not (layer0_outputs(2841));
    layer1_outputs(1789) <= not(layer0_outputs(3850));
    layer1_outputs(1790) <= '1';
    layer1_outputs(1791) <= not(layer0_outputs(633));
    layer1_outputs(1792) <= not(layer0_outputs(7315)) or (layer0_outputs(7570));
    layer1_outputs(1793) <= not(layer0_outputs(1271));
    layer1_outputs(1794) <= not((layer0_outputs(7138)) or (layer0_outputs(2504)));
    layer1_outputs(1795) <= (layer0_outputs(4635)) or (layer0_outputs(6218));
    layer1_outputs(1796) <= not(layer0_outputs(2235));
    layer1_outputs(1797) <= not(layer0_outputs(5373));
    layer1_outputs(1798) <= not(layer0_outputs(5167));
    layer1_outputs(1799) <= layer0_outputs(3319);
    layer1_outputs(1800) <= not(layer0_outputs(5854));
    layer1_outputs(1801) <= not(layer0_outputs(185)) or (layer0_outputs(3885));
    layer1_outputs(1802) <= (layer0_outputs(6868)) and not (layer0_outputs(3134));
    layer1_outputs(1803) <= '1';
    layer1_outputs(1804) <= not(layer0_outputs(4629)) or (layer0_outputs(5648));
    layer1_outputs(1805) <= (layer0_outputs(7446)) and not (layer0_outputs(1081));
    layer1_outputs(1806) <= layer0_outputs(2218);
    layer1_outputs(1807) <= not(layer0_outputs(1966)) or (layer0_outputs(708));
    layer1_outputs(1808) <= layer0_outputs(848);
    layer1_outputs(1809) <= not(layer0_outputs(4887));
    layer1_outputs(1810) <= not(layer0_outputs(764));
    layer1_outputs(1811) <= (layer0_outputs(1153)) or (layer0_outputs(5424));
    layer1_outputs(1812) <= (layer0_outputs(6266)) or (layer0_outputs(2956));
    layer1_outputs(1813) <= not(layer0_outputs(6678));
    layer1_outputs(1814) <= (layer0_outputs(6069)) and (layer0_outputs(542));
    layer1_outputs(1815) <= (layer0_outputs(1833)) xor (layer0_outputs(5086));
    layer1_outputs(1816) <= '1';
    layer1_outputs(1817) <= (layer0_outputs(7152)) and (layer0_outputs(3652));
    layer1_outputs(1818) <= not(layer0_outputs(4567)) or (layer0_outputs(783));
    layer1_outputs(1819) <= (layer0_outputs(5933)) or (layer0_outputs(369));
    layer1_outputs(1820) <= not(layer0_outputs(3315)) or (layer0_outputs(3899));
    layer1_outputs(1821) <= not((layer0_outputs(1268)) and (layer0_outputs(3307)));
    layer1_outputs(1822) <= (layer0_outputs(1893)) xor (layer0_outputs(1477));
    layer1_outputs(1823) <= '1';
    layer1_outputs(1824) <= layer0_outputs(3576);
    layer1_outputs(1825) <= (layer0_outputs(4123)) and (layer0_outputs(7212));
    layer1_outputs(1826) <= (layer0_outputs(42)) and (layer0_outputs(2580));
    layer1_outputs(1827) <= (layer0_outputs(1275)) and not (layer0_outputs(2332));
    layer1_outputs(1828) <= (layer0_outputs(1298)) and not (layer0_outputs(4200));
    layer1_outputs(1829) <= '0';
    layer1_outputs(1830) <= (layer0_outputs(6320)) and (layer0_outputs(4177));
    layer1_outputs(1831) <= (layer0_outputs(6684)) or (layer0_outputs(111));
    layer1_outputs(1832) <= (layer0_outputs(1858)) and not (layer0_outputs(4245));
    layer1_outputs(1833) <= layer0_outputs(6143);
    layer1_outputs(1834) <= not((layer0_outputs(2238)) xor (layer0_outputs(5949)));
    layer1_outputs(1835) <= not(layer0_outputs(5293));
    layer1_outputs(1836) <= '0';
    layer1_outputs(1837) <= '0';
    layer1_outputs(1838) <= '0';
    layer1_outputs(1839) <= not(layer0_outputs(5422));
    layer1_outputs(1840) <= layer0_outputs(992);
    layer1_outputs(1841) <= '1';
    layer1_outputs(1842) <= (layer0_outputs(3338)) and not (layer0_outputs(4410));
    layer1_outputs(1843) <= (layer0_outputs(1797)) and not (layer0_outputs(1292));
    layer1_outputs(1844) <= not((layer0_outputs(852)) or (layer0_outputs(1731)));
    layer1_outputs(1845) <= not(layer0_outputs(3912));
    layer1_outputs(1846) <= (layer0_outputs(6073)) and (layer0_outputs(3719));
    layer1_outputs(1847) <= (layer0_outputs(7354)) and not (layer0_outputs(5025));
    layer1_outputs(1848) <= not(layer0_outputs(3891));
    layer1_outputs(1849) <= '1';
    layer1_outputs(1850) <= layer0_outputs(7013);
    layer1_outputs(1851) <= (layer0_outputs(4659)) or (layer0_outputs(650));
    layer1_outputs(1852) <= not(layer0_outputs(1574));
    layer1_outputs(1853) <= not(layer0_outputs(3668));
    layer1_outputs(1854) <= not(layer0_outputs(611)) or (layer0_outputs(3299));
    layer1_outputs(1855) <= not(layer0_outputs(2388));
    layer1_outputs(1856) <= (layer0_outputs(3144)) and not (layer0_outputs(4191));
    layer1_outputs(1857) <= not(layer0_outputs(1650)) or (layer0_outputs(3893));
    layer1_outputs(1858) <= (layer0_outputs(3413)) and not (layer0_outputs(6887));
    layer1_outputs(1859) <= not((layer0_outputs(553)) xor (layer0_outputs(6636)));
    layer1_outputs(1860) <= (layer0_outputs(5562)) and not (layer0_outputs(6270));
    layer1_outputs(1861) <= '0';
    layer1_outputs(1862) <= not(layer0_outputs(5918)) or (layer0_outputs(6925));
    layer1_outputs(1863) <= (layer0_outputs(5842)) and not (layer0_outputs(1287));
    layer1_outputs(1864) <= not(layer0_outputs(6051)) or (layer0_outputs(1113));
    layer1_outputs(1865) <= not(layer0_outputs(4021));
    layer1_outputs(1866) <= layer0_outputs(4183);
    layer1_outputs(1867) <= not((layer0_outputs(1093)) xor (layer0_outputs(6481)));
    layer1_outputs(1868) <= not(layer0_outputs(1440)) or (layer0_outputs(1705));
    layer1_outputs(1869) <= (layer0_outputs(4925)) and not (layer0_outputs(7050));
    layer1_outputs(1870) <= not((layer0_outputs(3554)) or (layer0_outputs(4514)));
    layer1_outputs(1871) <= not(layer0_outputs(3295));
    layer1_outputs(1872) <= not(layer0_outputs(6131)) or (layer0_outputs(5147));
    layer1_outputs(1873) <= not(layer0_outputs(673));
    layer1_outputs(1874) <= not((layer0_outputs(7560)) or (layer0_outputs(3948)));
    layer1_outputs(1875) <= not(layer0_outputs(476));
    layer1_outputs(1876) <= layer0_outputs(5893);
    layer1_outputs(1877) <= not(layer0_outputs(5996));
    layer1_outputs(1878) <= (layer0_outputs(3827)) xor (layer0_outputs(5663));
    layer1_outputs(1879) <= not(layer0_outputs(4797)) or (layer0_outputs(4277));
    layer1_outputs(1880) <= (layer0_outputs(355)) and (layer0_outputs(1139));
    layer1_outputs(1881) <= not(layer0_outputs(3212)) or (layer0_outputs(298));
    layer1_outputs(1882) <= not((layer0_outputs(5120)) xor (layer0_outputs(4611)));
    layer1_outputs(1883) <= (layer0_outputs(7349)) and not (layer0_outputs(3734));
    layer1_outputs(1884) <= not(layer0_outputs(5133)) or (layer0_outputs(5030));
    layer1_outputs(1885) <= not(layer0_outputs(5776));
    layer1_outputs(1886) <= not(layer0_outputs(6190)) or (layer0_outputs(7048));
    layer1_outputs(1887) <= (layer0_outputs(4771)) xor (layer0_outputs(4982));
    layer1_outputs(1888) <= not(layer0_outputs(1541));
    layer1_outputs(1889) <= not(layer0_outputs(7556)) or (layer0_outputs(1552));
    layer1_outputs(1890) <= (layer0_outputs(3831)) and (layer0_outputs(1625));
    layer1_outputs(1891) <= not(layer0_outputs(901)) or (layer0_outputs(6559));
    layer1_outputs(1892) <= not(layer0_outputs(7001)) or (layer0_outputs(4621));
    layer1_outputs(1893) <= layer0_outputs(2074);
    layer1_outputs(1894) <= layer0_outputs(977);
    layer1_outputs(1895) <= (layer0_outputs(5758)) and not (layer0_outputs(6278));
    layer1_outputs(1896) <= not((layer0_outputs(4358)) xor (layer0_outputs(7272)));
    layer1_outputs(1897) <= (layer0_outputs(844)) and (layer0_outputs(3507));
    layer1_outputs(1898) <= (layer0_outputs(7650)) or (layer0_outputs(434));
    layer1_outputs(1899) <= not(layer0_outputs(850));
    layer1_outputs(1900) <= layer0_outputs(3119);
    layer1_outputs(1901) <= not(layer0_outputs(1273)) or (layer0_outputs(5533));
    layer1_outputs(1902) <= not((layer0_outputs(16)) or (layer0_outputs(6048)));
    layer1_outputs(1903) <= layer0_outputs(3405);
    layer1_outputs(1904) <= (layer0_outputs(240)) and not (layer0_outputs(7558));
    layer1_outputs(1905) <= (layer0_outputs(2202)) and (layer0_outputs(7457));
    layer1_outputs(1906) <= '0';
    layer1_outputs(1907) <= not(layer0_outputs(6214));
    layer1_outputs(1908) <= not((layer0_outputs(508)) or (layer0_outputs(3982)));
    layer1_outputs(1909) <= not(layer0_outputs(3014));
    layer1_outputs(1910) <= layer0_outputs(3099);
    layer1_outputs(1911) <= layer0_outputs(3364);
    layer1_outputs(1912) <= '0';
    layer1_outputs(1913) <= (layer0_outputs(6206)) and not (layer0_outputs(5895));
    layer1_outputs(1914) <= not(layer0_outputs(1205));
    layer1_outputs(1915) <= not(layer0_outputs(5627));
    layer1_outputs(1916) <= not((layer0_outputs(2468)) and (layer0_outputs(7629)));
    layer1_outputs(1917) <= not((layer0_outputs(4670)) or (layer0_outputs(1346)));
    layer1_outputs(1918) <= (layer0_outputs(842)) and not (layer0_outputs(7634));
    layer1_outputs(1919) <= layer0_outputs(2974);
    layer1_outputs(1920) <= (layer0_outputs(3872)) and (layer0_outputs(4213));
    layer1_outputs(1921) <= '0';
    layer1_outputs(1922) <= not((layer0_outputs(964)) and (layer0_outputs(5791)));
    layer1_outputs(1923) <= (layer0_outputs(5501)) or (layer0_outputs(4511));
    layer1_outputs(1924) <= not(layer0_outputs(1458));
    layer1_outputs(1925) <= (layer0_outputs(5190)) or (layer0_outputs(7620));
    layer1_outputs(1926) <= not(layer0_outputs(3628));
    layer1_outputs(1927) <= layer0_outputs(1285);
    layer1_outputs(1928) <= not(layer0_outputs(5065)) or (layer0_outputs(4424));
    layer1_outputs(1929) <= layer0_outputs(4443);
    layer1_outputs(1930) <= not(layer0_outputs(3838)) or (layer0_outputs(6817));
    layer1_outputs(1931) <= not((layer0_outputs(119)) or (layer0_outputs(7040)));
    layer1_outputs(1932) <= not((layer0_outputs(3096)) xor (layer0_outputs(6626)));
    layer1_outputs(1933) <= (layer0_outputs(6419)) and (layer0_outputs(202));
    layer1_outputs(1934) <= (layer0_outputs(6352)) or (layer0_outputs(3438));
    layer1_outputs(1935) <= not(layer0_outputs(4534));
    layer1_outputs(1936) <= not(layer0_outputs(2564));
    layer1_outputs(1937) <= not((layer0_outputs(3589)) or (layer0_outputs(7490)));
    layer1_outputs(1938) <= (layer0_outputs(5066)) and not (layer0_outputs(5482));
    layer1_outputs(1939) <= '1';
    layer1_outputs(1940) <= not(layer0_outputs(4908));
    layer1_outputs(1941) <= not(layer0_outputs(3080)) or (layer0_outputs(7015));
    layer1_outputs(1942) <= (layer0_outputs(561)) or (layer0_outputs(2931));
    layer1_outputs(1943) <= layer0_outputs(6975);
    layer1_outputs(1944) <= (layer0_outputs(3011)) and not (layer0_outputs(5064));
    layer1_outputs(1945) <= (layer0_outputs(1201)) or (layer0_outputs(5586));
    layer1_outputs(1946) <= (layer0_outputs(1633)) and not (layer0_outputs(26));
    layer1_outputs(1947) <= not((layer0_outputs(393)) or (layer0_outputs(2152)));
    layer1_outputs(1948) <= not((layer0_outputs(2315)) or (layer0_outputs(5442)));
    layer1_outputs(1949) <= (layer0_outputs(4593)) and not (layer0_outputs(1468));
    layer1_outputs(1950) <= not(layer0_outputs(1815));
    layer1_outputs(1951) <= not(layer0_outputs(7619)) or (layer0_outputs(7506));
    layer1_outputs(1952) <= not((layer0_outputs(2934)) and (layer0_outputs(1321)));
    layer1_outputs(1953) <= not(layer0_outputs(5780));
    layer1_outputs(1954) <= '0';
    layer1_outputs(1955) <= not((layer0_outputs(4862)) or (layer0_outputs(7269)));
    layer1_outputs(1956) <= (layer0_outputs(7081)) or (layer0_outputs(2859));
    layer1_outputs(1957) <= layer0_outputs(2575);
    layer1_outputs(1958) <= not(layer0_outputs(4469));
    layer1_outputs(1959) <= (layer0_outputs(2498)) and not (layer0_outputs(2912));
    layer1_outputs(1960) <= (layer0_outputs(4422)) and not (layer0_outputs(6253));
    layer1_outputs(1961) <= not(layer0_outputs(4787));
    layer1_outputs(1962) <= not(layer0_outputs(1056));
    layer1_outputs(1963) <= not(layer0_outputs(838));
    layer1_outputs(1964) <= not(layer0_outputs(1202));
    layer1_outputs(1965) <= layer0_outputs(2414);
    layer1_outputs(1966) <= layer0_outputs(2512);
    layer1_outputs(1967) <= (layer0_outputs(1536)) and not (layer0_outputs(4953));
    layer1_outputs(1968) <= not((layer0_outputs(5305)) and (layer0_outputs(6101)));
    layer1_outputs(1969) <= not(layer0_outputs(2030)) or (layer0_outputs(1337));
    layer1_outputs(1970) <= not(layer0_outputs(5769)) or (layer0_outputs(5098));
    layer1_outputs(1971) <= not((layer0_outputs(845)) and (layer0_outputs(179)));
    layer1_outputs(1972) <= (layer0_outputs(1026)) and not (layer0_outputs(1001));
    layer1_outputs(1973) <= not(layer0_outputs(414)) or (layer0_outputs(5860));
    layer1_outputs(1974) <= layer0_outputs(6386);
    layer1_outputs(1975) <= not((layer0_outputs(956)) and (layer0_outputs(5107)));
    layer1_outputs(1976) <= not((layer0_outputs(1822)) or (layer0_outputs(7564)));
    layer1_outputs(1977) <= not((layer0_outputs(3248)) or (layer0_outputs(6163)));
    layer1_outputs(1978) <= layer0_outputs(6162);
    layer1_outputs(1979) <= '1';
    layer1_outputs(1980) <= not((layer0_outputs(3379)) and (layer0_outputs(1879)));
    layer1_outputs(1981) <= not(layer0_outputs(4606)) or (layer0_outputs(418));
    layer1_outputs(1982) <= not(layer0_outputs(7358));
    layer1_outputs(1983) <= (layer0_outputs(3985)) and (layer0_outputs(3274));
    layer1_outputs(1984) <= layer0_outputs(5417);
    layer1_outputs(1985) <= not((layer0_outputs(4873)) and (layer0_outputs(4258)));
    layer1_outputs(1986) <= not(layer0_outputs(4727));
    layer1_outputs(1987) <= (layer0_outputs(2277)) xor (layer0_outputs(2488));
    layer1_outputs(1988) <= (layer0_outputs(6460)) or (layer0_outputs(1422));
    layer1_outputs(1989) <= (layer0_outputs(3844)) and not (layer0_outputs(5542));
    layer1_outputs(1990) <= not(layer0_outputs(7307)) or (layer0_outputs(4494));
    layer1_outputs(1991) <= not(layer0_outputs(5731)) or (layer0_outputs(1425));
    layer1_outputs(1992) <= '0';
    layer1_outputs(1993) <= (layer0_outputs(6455)) and not (layer0_outputs(894));
    layer1_outputs(1994) <= (layer0_outputs(2437)) and not (layer0_outputs(7477));
    layer1_outputs(1995) <= not((layer0_outputs(5474)) and (layer0_outputs(5937)));
    layer1_outputs(1996) <= not(layer0_outputs(1363)) or (layer0_outputs(2370));
    layer1_outputs(1997) <= not(layer0_outputs(1125)) or (layer0_outputs(2636));
    layer1_outputs(1998) <= (layer0_outputs(3197)) and not (layer0_outputs(1179));
    layer1_outputs(1999) <= '1';
    layer1_outputs(2000) <= '0';
    layer1_outputs(2001) <= layer0_outputs(4805);
    layer1_outputs(2002) <= layer0_outputs(7360);
    layer1_outputs(2003) <= not((layer0_outputs(102)) or (layer0_outputs(841)));
    layer1_outputs(2004) <= not((layer0_outputs(4001)) and (layer0_outputs(6940)));
    layer1_outputs(2005) <= (layer0_outputs(3653)) and (layer0_outputs(6322));
    layer1_outputs(2006) <= (layer0_outputs(3082)) and not (layer0_outputs(5563));
    layer1_outputs(2007) <= (layer0_outputs(3794)) and not (layer0_outputs(3018));
    layer1_outputs(2008) <= not((layer0_outputs(259)) and (layer0_outputs(7399)));
    layer1_outputs(2009) <= not(layer0_outputs(5290));
    layer1_outputs(2010) <= not(layer0_outputs(2909));
    layer1_outputs(2011) <= '0';
    layer1_outputs(2012) <= (layer0_outputs(4339)) and (layer0_outputs(2229));
    layer1_outputs(2013) <= not(layer0_outputs(4903));
    layer1_outputs(2014) <= (layer0_outputs(7420)) or (layer0_outputs(745));
    layer1_outputs(2015) <= (layer0_outputs(2383)) and (layer0_outputs(765));
    layer1_outputs(2016) <= layer0_outputs(4954);
    layer1_outputs(2017) <= not((layer0_outputs(2935)) and (layer0_outputs(6389)));
    layer1_outputs(2018) <= not(layer0_outputs(2087)) or (layer0_outputs(4274));
    layer1_outputs(2019) <= not((layer0_outputs(2338)) xor (layer0_outputs(4042)));
    layer1_outputs(2020) <= not((layer0_outputs(6006)) xor (layer0_outputs(7163)));
    layer1_outputs(2021) <= (layer0_outputs(1768)) and not (layer0_outputs(184));
    layer1_outputs(2022) <= not(layer0_outputs(178));
    layer1_outputs(2023) <= layer0_outputs(2616);
    layer1_outputs(2024) <= (layer0_outputs(5177)) xor (layer0_outputs(6688));
    layer1_outputs(2025) <= not((layer0_outputs(1750)) and (layer0_outputs(6264)));
    layer1_outputs(2026) <= (layer0_outputs(7483)) and not (layer0_outputs(786));
    layer1_outputs(2027) <= layer0_outputs(5725);
    layer1_outputs(2028) <= layer0_outputs(6362);
    layer1_outputs(2029) <= (layer0_outputs(5260)) and (layer0_outputs(3953));
    layer1_outputs(2030) <= not(layer0_outputs(6484)) or (layer0_outputs(6781));
    layer1_outputs(2031) <= not(layer0_outputs(1949)) or (layer0_outputs(2124));
    layer1_outputs(2032) <= not(layer0_outputs(7309));
    layer1_outputs(2033) <= layer0_outputs(3658);
    layer1_outputs(2034) <= not((layer0_outputs(1145)) or (layer0_outputs(4579)));
    layer1_outputs(2035) <= (layer0_outputs(6225)) and not (layer0_outputs(2984));
    layer1_outputs(2036) <= layer0_outputs(6619);
    layer1_outputs(2037) <= '0';
    layer1_outputs(2038) <= not((layer0_outputs(5061)) and (layer0_outputs(4094)));
    layer1_outputs(2039) <= not((layer0_outputs(1997)) or (layer0_outputs(1349)));
    layer1_outputs(2040) <= (layer0_outputs(1790)) and not (layer0_outputs(3165));
    layer1_outputs(2041) <= '0';
    layer1_outputs(2042) <= layer0_outputs(6120);
    layer1_outputs(2043) <= not(layer0_outputs(7078));
    layer1_outputs(2044) <= not((layer0_outputs(6646)) xor (layer0_outputs(6539)));
    layer1_outputs(2045) <= '1';
    layer1_outputs(2046) <= not((layer0_outputs(5048)) and (layer0_outputs(3401)));
    layer1_outputs(2047) <= layer0_outputs(6);
    layer1_outputs(2048) <= layer0_outputs(1895);
    layer1_outputs(2049) <= (layer0_outputs(6654)) or (layer0_outputs(5736));
    layer1_outputs(2050) <= '0';
    layer1_outputs(2051) <= (layer0_outputs(2542)) or (layer0_outputs(7452));
    layer1_outputs(2052) <= not(layer0_outputs(2227)) or (layer0_outputs(852));
    layer1_outputs(2053) <= '0';
    layer1_outputs(2054) <= not(layer0_outputs(7312)) or (layer0_outputs(5765));
    layer1_outputs(2055) <= layer0_outputs(5358);
    layer1_outputs(2056) <= (layer0_outputs(587)) and not (layer0_outputs(2351));
    layer1_outputs(2057) <= not(layer0_outputs(7495));
    layer1_outputs(2058) <= not(layer0_outputs(797)) or (layer0_outputs(2725));
    layer1_outputs(2059) <= layer0_outputs(7635);
    layer1_outputs(2060) <= layer0_outputs(4626);
    layer1_outputs(2061) <= '0';
    layer1_outputs(2062) <= layer0_outputs(3657);
    layer1_outputs(2063) <= not((layer0_outputs(5800)) or (layer0_outputs(1396)));
    layer1_outputs(2064) <= not(layer0_outputs(1274));
    layer1_outputs(2065) <= layer0_outputs(5095);
    layer1_outputs(2066) <= layer0_outputs(1488);
    layer1_outputs(2067) <= '0';
    layer1_outputs(2068) <= layer0_outputs(4849);
    layer1_outputs(2069) <= not(layer0_outputs(5795)) or (layer0_outputs(5166));
    layer1_outputs(2070) <= '1';
    layer1_outputs(2071) <= (layer0_outputs(1499)) and not (layer0_outputs(1766));
    layer1_outputs(2072) <= not(layer0_outputs(4767));
    layer1_outputs(2073) <= not(layer0_outputs(5969));
    layer1_outputs(2074) <= layer0_outputs(5038);
    layer1_outputs(2075) <= not((layer0_outputs(4755)) and (layer0_outputs(913)));
    layer1_outputs(2076) <= layer0_outputs(592);
    layer1_outputs(2077) <= not(layer0_outputs(7229));
    layer1_outputs(2078) <= (layer0_outputs(3617)) and not (layer0_outputs(2408));
    layer1_outputs(2079) <= not(layer0_outputs(6146)) or (layer0_outputs(3398));
    layer1_outputs(2080) <= '1';
    layer1_outputs(2081) <= layer0_outputs(1018);
    layer1_outputs(2082) <= not(layer0_outputs(1954)) or (layer0_outputs(2164));
    layer1_outputs(2083) <= '1';
    layer1_outputs(2084) <= '1';
    layer1_outputs(2085) <= layer0_outputs(3593);
    layer1_outputs(2086) <= layer0_outputs(4626);
    layer1_outputs(2087) <= not((layer0_outputs(2598)) and (layer0_outputs(4618)));
    layer1_outputs(2088) <= not(layer0_outputs(2103)) or (layer0_outputs(4100));
    layer1_outputs(2089) <= not(layer0_outputs(4582));
    layer1_outputs(2090) <= not(layer0_outputs(943));
    layer1_outputs(2091) <= layer0_outputs(5669);
    layer1_outputs(2092) <= not(layer0_outputs(6188));
    layer1_outputs(2093) <= (layer0_outputs(4267)) and (layer0_outputs(3049));
    layer1_outputs(2094) <= not(layer0_outputs(6147));
    layer1_outputs(2095) <= not(layer0_outputs(5704));
    layer1_outputs(2096) <= '0';
    layer1_outputs(2097) <= not((layer0_outputs(5978)) or (layer0_outputs(368)));
    layer1_outputs(2098) <= not(layer0_outputs(6539));
    layer1_outputs(2099) <= not(layer0_outputs(4392));
    layer1_outputs(2100) <= (layer0_outputs(2807)) and not (layer0_outputs(1415));
    layer1_outputs(2101) <= not((layer0_outputs(6322)) or (layer0_outputs(6182)));
    layer1_outputs(2102) <= '1';
    layer1_outputs(2103) <= (layer0_outputs(1362)) and (layer0_outputs(4293));
    layer1_outputs(2104) <= not(layer0_outputs(774)) or (layer0_outputs(6494));
    layer1_outputs(2105) <= not(layer0_outputs(7530)) or (layer0_outputs(4547));
    layer1_outputs(2106) <= not((layer0_outputs(1939)) and (layer0_outputs(688)));
    layer1_outputs(2107) <= layer0_outputs(1636);
    layer1_outputs(2108) <= not(layer0_outputs(1525));
    layer1_outputs(2109) <= not((layer0_outputs(6287)) and (layer0_outputs(1923)));
    layer1_outputs(2110) <= not(layer0_outputs(3911));
    layer1_outputs(2111) <= layer0_outputs(6592);
    layer1_outputs(2112) <= not((layer0_outputs(2351)) and (layer0_outputs(3132)));
    layer1_outputs(2113) <= '0';
    layer1_outputs(2114) <= not((layer0_outputs(4027)) and (layer0_outputs(5368)));
    layer1_outputs(2115) <= not(layer0_outputs(2178));
    layer1_outputs(2116) <= not(layer0_outputs(1622));
    layer1_outputs(2117) <= '1';
    layer1_outputs(2118) <= layer0_outputs(582);
    layer1_outputs(2119) <= '1';
    layer1_outputs(2120) <= not((layer0_outputs(979)) xor (layer0_outputs(7146)));
    layer1_outputs(2121) <= not((layer0_outputs(5456)) and (layer0_outputs(3627)));
    layer1_outputs(2122) <= (layer0_outputs(6713)) xor (layer0_outputs(5997));
    layer1_outputs(2123) <= not((layer0_outputs(1060)) or (layer0_outputs(6804)));
    layer1_outputs(2124) <= not(layer0_outputs(646)) or (layer0_outputs(5922));
    layer1_outputs(2125) <= (layer0_outputs(1316)) and not (layer0_outputs(1571));
    layer1_outputs(2126) <= not((layer0_outputs(1970)) or (layer0_outputs(307)));
    layer1_outputs(2127) <= '0';
    layer1_outputs(2128) <= layer0_outputs(11);
    layer1_outputs(2129) <= not((layer0_outputs(6806)) and (layer0_outputs(2328)));
    layer1_outputs(2130) <= not(layer0_outputs(866)) or (layer0_outputs(3718));
    layer1_outputs(2131) <= not(layer0_outputs(6282));
    layer1_outputs(2132) <= not((layer0_outputs(4152)) and (layer0_outputs(4658)));
    layer1_outputs(2133) <= not(layer0_outputs(1518)) or (layer0_outputs(6710));
    layer1_outputs(2134) <= (layer0_outputs(5087)) and not (layer0_outputs(6350));
    layer1_outputs(2135) <= not(layer0_outputs(4069)) or (layer0_outputs(7116));
    layer1_outputs(2136) <= not(layer0_outputs(2736));
    layer1_outputs(2137) <= (layer0_outputs(6869)) or (layer0_outputs(1613));
    layer1_outputs(2138) <= not(layer0_outputs(4976)) or (layer0_outputs(2693));
    layer1_outputs(2139) <= not((layer0_outputs(5927)) or (layer0_outputs(4797)));
    layer1_outputs(2140) <= (layer0_outputs(4078)) or (layer0_outputs(6078));
    layer1_outputs(2141) <= not((layer0_outputs(3868)) and (layer0_outputs(5864)));
    layer1_outputs(2142) <= not(layer0_outputs(5148));
    layer1_outputs(2143) <= (layer0_outputs(5794)) xor (layer0_outputs(3768));
    layer1_outputs(2144) <= (layer0_outputs(426)) and not (layer0_outputs(5756));
    layer1_outputs(2145) <= not((layer0_outputs(2106)) or (layer0_outputs(4812)));
    layer1_outputs(2146) <= not(layer0_outputs(4315)) or (layer0_outputs(7403));
    layer1_outputs(2147) <= (layer0_outputs(6587)) and not (layer0_outputs(6655));
    layer1_outputs(2148) <= layer0_outputs(5455);
    layer1_outputs(2149) <= layer0_outputs(1404);
    layer1_outputs(2150) <= (layer0_outputs(496)) or (layer0_outputs(5850));
    layer1_outputs(2151) <= not(layer0_outputs(2130));
    layer1_outputs(2152) <= not((layer0_outputs(1444)) or (layer0_outputs(4877)));
    layer1_outputs(2153) <= '0';
    layer1_outputs(2154) <= layer0_outputs(3603);
    layer1_outputs(2155) <= (layer0_outputs(2189)) and (layer0_outputs(2803));
    layer1_outputs(2156) <= (layer0_outputs(4045)) and not (layer0_outputs(3280));
    layer1_outputs(2157) <= not(layer0_outputs(7148));
    layer1_outputs(2158) <= not(layer0_outputs(4363)) or (layer0_outputs(833));
    layer1_outputs(2159) <= not(layer0_outputs(1264));
    layer1_outputs(2160) <= not(layer0_outputs(5520)) or (layer0_outputs(2594));
    layer1_outputs(2161) <= (layer0_outputs(5985)) and (layer0_outputs(4965));
    layer1_outputs(2162) <= (layer0_outputs(5168)) or (layer0_outputs(1731));
    layer1_outputs(2163) <= (layer0_outputs(6732)) and not (layer0_outputs(1801));
    layer1_outputs(2164) <= not(layer0_outputs(3168));
    layer1_outputs(2165) <= not((layer0_outputs(1181)) or (layer0_outputs(4842)));
    layer1_outputs(2166) <= layer0_outputs(7230);
    layer1_outputs(2167) <= (layer0_outputs(458)) or (layer0_outputs(2460));
    layer1_outputs(2168) <= (layer0_outputs(3402)) and not (layer0_outputs(3659));
    layer1_outputs(2169) <= not(layer0_outputs(5688));
    layer1_outputs(2170) <= layer0_outputs(5863);
    layer1_outputs(2171) <= not((layer0_outputs(4596)) and (layer0_outputs(4748)));
    layer1_outputs(2172) <= not(layer0_outputs(3663));
    layer1_outputs(2173) <= (layer0_outputs(2126)) and not (layer0_outputs(1757));
    layer1_outputs(2174) <= layer0_outputs(5820);
    layer1_outputs(2175) <= (layer0_outputs(1802)) and not (layer0_outputs(5698));
    layer1_outputs(2176) <= '1';
    layer1_outputs(2177) <= not(layer0_outputs(359)) or (layer0_outputs(5837));
    layer1_outputs(2178) <= (layer0_outputs(3371)) or (layer0_outputs(4943));
    layer1_outputs(2179) <= layer0_outputs(1054);
    layer1_outputs(2180) <= layer0_outputs(1561);
    layer1_outputs(2181) <= layer0_outputs(3200);
    layer1_outputs(2182) <= not((layer0_outputs(952)) xor (layer0_outputs(7437)));
    layer1_outputs(2183) <= not(layer0_outputs(82));
    layer1_outputs(2184) <= (layer0_outputs(1302)) xor (layer0_outputs(874));
    layer1_outputs(2185) <= layer0_outputs(5339);
    layer1_outputs(2186) <= layer0_outputs(939);
    layer1_outputs(2187) <= not(layer0_outputs(1950)) or (layer0_outputs(3447));
    layer1_outputs(2188) <= (layer0_outputs(7232)) and not (layer0_outputs(4440));
    layer1_outputs(2189) <= not((layer0_outputs(802)) and (layer0_outputs(6846)));
    layer1_outputs(2190) <= (layer0_outputs(5662)) and (layer0_outputs(7114));
    layer1_outputs(2191) <= not((layer0_outputs(3088)) or (layer0_outputs(2290)));
    layer1_outputs(2192) <= '1';
    layer1_outputs(2193) <= '0';
    layer1_outputs(2194) <= layer0_outputs(6204);
    layer1_outputs(2195) <= not(layer0_outputs(1643)) or (layer0_outputs(2538));
    layer1_outputs(2196) <= not((layer0_outputs(4110)) and (layer0_outputs(4900)));
    layer1_outputs(2197) <= not((layer0_outputs(2626)) and (layer0_outputs(2213)));
    layer1_outputs(2198) <= '1';
    layer1_outputs(2199) <= (layer0_outputs(4497)) and not (layer0_outputs(5086));
    layer1_outputs(2200) <= layer0_outputs(128);
    layer1_outputs(2201) <= (layer0_outputs(4638)) and not (layer0_outputs(1555));
    layer1_outputs(2202) <= (layer0_outputs(6894)) and not (layer0_outputs(2229));
    layer1_outputs(2203) <= not((layer0_outputs(660)) and (layer0_outputs(7010)));
    layer1_outputs(2204) <= not(layer0_outputs(2940));
    layer1_outputs(2205) <= not(layer0_outputs(412)) or (layer0_outputs(7537));
    layer1_outputs(2206) <= (layer0_outputs(3944)) and (layer0_outputs(4219));
    layer1_outputs(2207) <= not(layer0_outputs(4395));
    layer1_outputs(2208) <= not(layer0_outputs(3761));
    layer1_outputs(2209) <= not((layer0_outputs(6083)) or (layer0_outputs(7576)));
    layer1_outputs(2210) <= (layer0_outputs(4362)) or (layer0_outputs(2487));
    layer1_outputs(2211) <= layer0_outputs(998);
    layer1_outputs(2212) <= layer0_outputs(467);
    layer1_outputs(2213) <= layer0_outputs(1506);
    layer1_outputs(2214) <= not(layer0_outputs(3000)) or (layer0_outputs(4603));
    layer1_outputs(2215) <= not(layer0_outputs(7230)) or (layer0_outputs(1306));
    layer1_outputs(2216) <= not((layer0_outputs(163)) or (layer0_outputs(3960)));
    layer1_outputs(2217) <= (layer0_outputs(3597)) xor (layer0_outputs(101));
    layer1_outputs(2218) <= not((layer0_outputs(1856)) and (layer0_outputs(7573)));
    layer1_outputs(2219) <= layer0_outputs(6504);
    layer1_outputs(2220) <= layer0_outputs(7485);
    layer1_outputs(2221) <= not(layer0_outputs(365)) or (layer0_outputs(408));
    layer1_outputs(2222) <= not((layer0_outputs(7361)) and (layer0_outputs(4417)));
    layer1_outputs(2223) <= '0';
    layer1_outputs(2224) <= not((layer0_outputs(1168)) or (layer0_outputs(2845)));
    layer1_outputs(2225) <= '0';
    layer1_outputs(2226) <= '1';
    layer1_outputs(2227) <= layer0_outputs(2855);
    layer1_outputs(2228) <= not((layer0_outputs(2537)) and (layer0_outputs(1946)));
    layer1_outputs(2229) <= (layer0_outputs(7244)) and (layer0_outputs(7125));
    layer1_outputs(2230) <= (layer0_outputs(3611)) and (layer0_outputs(6370));
    layer1_outputs(2231) <= layer0_outputs(1844);
    layer1_outputs(2232) <= layer0_outputs(6342);
    layer1_outputs(2233) <= not((layer0_outputs(7119)) and (layer0_outputs(6759)));
    layer1_outputs(2234) <= not(layer0_outputs(5714)) or (layer0_outputs(3965));
    layer1_outputs(2235) <= layer0_outputs(5473);
    layer1_outputs(2236) <= not(layer0_outputs(2654));
    layer1_outputs(2237) <= not(layer0_outputs(4717)) or (layer0_outputs(2663));
    layer1_outputs(2238) <= '0';
    layer1_outputs(2239) <= (layer0_outputs(3915)) and not (layer0_outputs(6194));
    layer1_outputs(2240) <= layer0_outputs(7009);
    layer1_outputs(2241) <= not(layer0_outputs(2720));
    layer1_outputs(2242) <= (layer0_outputs(7331)) and not (layer0_outputs(2183));
    layer1_outputs(2243) <= not((layer0_outputs(39)) or (layer0_outputs(1324)));
    layer1_outputs(2244) <= not(layer0_outputs(2885));
    layer1_outputs(2245) <= layer0_outputs(3281);
    layer1_outputs(2246) <= not(layer0_outputs(3216)) or (layer0_outputs(4433));
    layer1_outputs(2247) <= (layer0_outputs(1937)) xor (layer0_outputs(7366));
    layer1_outputs(2248) <= not(layer0_outputs(4858));
    layer1_outputs(2249) <= not((layer0_outputs(1612)) xor (layer0_outputs(2653)));
    layer1_outputs(2250) <= not(layer0_outputs(5192)) or (layer0_outputs(996));
    layer1_outputs(2251) <= layer0_outputs(1054);
    layer1_outputs(2252) <= (layer0_outputs(5859)) xor (layer0_outputs(7511));
    layer1_outputs(2253) <= (layer0_outputs(292)) and (layer0_outputs(5355));
    layer1_outputs(2254) <= (layer0_outputs(250)) or (layer0_outputs(6812));
    layer1_outputs(2255) <= (layer0_outputs(7531)) and not (layer0_outputs(1052));
    layer1_outputs(2256) <= '1';
    layer1_outputs(2257) <= (layer0_outputs(715)) and not (layer0_outputs(3827));
    layer1_outputs(2258) <= (layer0_outputs(3427)) and not (layer0_outputs(4121));
    layer1_outputs(2259) <= not(layer0_outputs(6114)) or (layer0_outputs(4380));
    layer1_outputs(2260) <= (layer0_outputs(6837)) or (layer0_outputs(2429));
    layer1_outputs(2261) <= (layer0_outputs(4621)) and (layer0_outputs(7359));
    layer1_outputs(2262) <= layer0_outputs(938);
    layer1_outputs(2263) <= not(layer0_outputs(3297)) or (layer0_outputs(6286));
    layer1_outputs(2264) <= not(layer0_outputs(7310)) or (layer0_outputs(6480));
    layer1_outputs(2265) <= (layer0_outputs(3100)) and not (layer0_outputs(902));
    layer1_outputs(2266) <= '1';
    layer1_outputs(2267) <= layer0_outputs(779);
    layer1_outputs(2268) <= not(layer0_outputs(6185));
    layer1_outputs(2269) <= not(layer0_outputs(3782)) or (layer0_outputs(6138));
    layer1_outputs(2270) <= '0';
    layer1_outputs(2271) <= not(layer0_outputs(1247)) or (layer0_outputs(4376));
    layer1_outputs(2272) <= not(layer0_outputs(7514)) or (layer0_outputs(3553));
    layer1_outputs(2273) <= not(layer0_outputs(6802));
    layer1_outputs(2274) <= not(layer0_outputs(4076));
    layer1_outputs(2275) <= not((layer0_outputs(235)) or (layer0_outputs(5657)));
    layer1_outputs(2276) <= (layer0_outputs(6283)) and not (layer0_outputs(5338));
    layer1_outputs(2277) <= not(layer0_outputs(4731));
    layer1_outputs(2278) <= (layer0_outputs(6198)) and (layer0_outputs(1669));
    layer1_outputs(2279) <= not((layer0_outputs(4639)) or (layer0_outputs(4782)));
    layer1_outputs(2280) <= not(layer0_outputs(4551));
    layer1_outputs(2281) <= layer0_outputs(6516);
    layer1_outputs(2282) <= not(layer0_outputs(4500)) or (layer0_outputs(2380));
    layer1_outputs(2283) <= (layer0_outputs(3075)) or (layer0_outputs(1906));
    layer1_outputs(2284) <= not((layer0_outputs(3578)) and (layer0_outputs(1744)));
    layer1_outputs(2285) <= '0';
    layer1_outputs(2286) <= layer0_outputs(4032);
    layer1_outputs(2287) <= not(layer0_outputs(2057)) or (layer0_outputs(1229));
    layer1_outputs(2288) <= not(layer0_outputs(6946));
    layer1_outputs(2289) <= not(layer0_outputs(2824));
    layer1_outputs(2290) <= not(layer0_outputs(7374));
    layer1_outputs(2291) <= (layer0_outputs(7678)) and (layer0_outputs(23));
    layer1_outputs(2292) <= '1';
    layer1_outputs(2293) <= (layer0_outputs(4564)) and (layer0_outputs(4678));
    layer1_outputs(2294) <= layer0_outputs(6354);
    layer1_outputs(2295) <= '1';
    layer1_outputs(2296) <= (layer0_outputs(5554)) and not (layer0_outputs(7266));
    layer1_outputs(2297) <= not((layer0_outputs(3790)) or (layer0_outputs(1010)));
    layer1_outputs(2298) <= not(layer0_outputs(6343)) or (layer0_outputs(4481));
    layer1_outputs(2299) <= layer0_outputs(3384);
    layer1_outputs(2300) <= layer0_outputs(1542);
    layer1_outputs(2301) <= (layer0_outputs(3313)) and not (layer0_outputs(945));
    layer1_outputs(2302) <= layer0_outputs(3741);
    layer1_outputs(2303) <= not(layer0_outputs(7058));
    layer1_outputs(2304) <= (layer0_outputs(7184)) and (layer0_outputs(6563));
    layer1_outputs(2305) <= (layer0_outputs(2503)) or (layer0_outputs(4145));
    layer1_outputs(2306) <= not(layer0_outputs(7504));
    layer1_outputs(2307) <= layer0_outputs(4301);
    layer1_outputs(2308) <= layer0_outputs(2813);
    layer1_outputs(2309) <= not((layer0_outputs(1942)) and (layer0_outputs(5774)));
    layer1_outputs(2310) <= layer0_outputs(4227);
    layer1_outputs(2311) <= layer0_outputs(5383);
    layer1_outputs(2312) <= (layer0_outputs(1808)) and not (layer0_outputs(2571));
    layer1_outputs(2313) <= (layer0_outputs(5597)) and not (layer0_outputs(6795));
    layer1_outputs(2314) <= not(layer0_outputs(102));
    layer1_outputs(2315) <= (layer0_outputs(5489)) or (layer0_outputs(740));
    layer1_outputs(2316) <= not(layer0_outputs(7107)) or (layer0_outputs(1489));
    layer1_outputs(2317) <= (layer0_outputs(6911)) and not (layer0_outputs(4003));
    layer1_outputs(2318) <= '0';
    layer1_outputs(2319) <= not((layer0_outputs(3846)) and (layer0_outputs(4676)));
    layer1_outputs(2320) <= (layer0_outputs(2075)) and not (layer0_outputs(6677));
    layer1_outputs(2321) <= (layer0_outputs(1942)) and not (layer0_outputs(4704));
    layer1_outputs(2322) <= not(layer0_outputs(7470)) or (layer0_outputs(6578));
    layer1_outputs(2323) <= not(layer0_outputs(212));
    layer1_outputs(2324) <= layer0_outputs(3058);
    layer1_outputs(2325) <= layer0_outputs(4175);
    layer1_outputs(2326) <= not(layer0_outputs(357));
    layer1_outputs(2327) <= layer0_outputs(9);
    layer1_outputs(2328) <= not((layer0_outputs(5252)) and (layer0_outputs(431)));
    layer1_outputs(2329) <= not(layer0_outputs(6379)) or (layer0_outputs(5762));
    layer1_outputs(2330) <= (layer0_outputs(3304)) or (layer0_outputs(2217));
    layer1_outputs(2331) <= layer0_outputs(1399);
    layer1_outputs(2332) <= not(layer0_outputs(6963)) or (layer0_outputs(2983));
    layer1_outputs(2333) <= layer0_outputs(6116);
    layer1_outputs(2334) <= not(layer0_outputs(2645));
    layer1_outputs(2335) <= layer0_outputs(5149);
    layer1_outputs(2336) <= not(layer0_outputs(6172));
    layer1_outputs(2337) <= (layer0_outputs(3267)) or (layer0_outputs(4550));
    layer1_outputs(2338) <= not(layer0_outputs(3656)) or (layer0_outputs(7401));
    layer1_outputs(2339) <= (layer0_outputs(4411)) xor (layer0_outputs(2622));
    layer1_outputs(2340) <= layer0_outputs(7238);
    layer1_outputs(2341) <= not((layer0_outputs(564)) or (layer0_outputs(5377)));
    layer1_outputs(2342) <= (layer0_outputs(6803)) and not (layer0_outputs(3535));
    layer1_outputs(2343) <= layer0_outputs(7321);
    layer1_outputs(2344) <= layer0_outputs(6880);
    layer1_outputs(2345) <= not((layer0_outputs(410)) or (layer0_outputs(7064)));
    layer1_outputs(2346) <= not(layer0_outputs(2181));
    layer1_outputs(2347) <= layer0_outputs(6773);
    layer1_outputs(2348) <= not((layer0_outputs(1023)) or (layer0_outputs(6142)));
    layer1_outputs(2349) <= not(layer0_outputs(3664));
    layer1_outputs(2350) <= '0';
    layer1_outputs(2351) <= (layer0_outputs(5867)) and (layer0_outputs(2341));
    layer1_outputs(2352) <= not(layer0_outputs(5747));
    layer1_outputs(2353) <= '1';
    layer1_outputs(2354) <= not((layer0_outputs(3071)) or (layer0_outputs(2479)));
    layer1_outputs(2355) <= not(layer0_outputs(2920));
    layer1_outputs(2356) <= (layer0_outputs(4167)) xor (layer0_outputs(3632));
    layer1_outputs(2357) <= not(layer0_outputs(5408)) or (layer0_outputs(1837));
    layer1_outputs(2358) <= not(layer0_outputs(7648)) or (layer0_outputs(42));
    layer1_outputs(2359) <= (layer0_outputs(7192)) and not (layer0_outputs(2660));
    layer1_outputs(2360) <= not((layer0_outputs(1713)) or (layer0_outputs(5786)));
    layer1_outputs(2361) <= not(layer0_outputs(5015));
    layer1_outputs(2362) <= (layer0_outputs(1217)) and not (layer0_outputs(4470));
    layer1_outputs(2363) <= not((layer0_outputs(6964)) xor (layer0_outputs(7058)));
    layer1_outputs(2364) <= '0';
    layer1_outputs(2365) <= (layer0_outputs(4478)) or (layer0_outputs(3852));
    layer1_outputs(2366) <= not(layer0_outputs(1059));
    layer1_outputs(2367) <= not(layer0_outputs(62));
    layer1_outputs(2368) <= not(layer0_outputs(5400));
    layer1_outputs(2369) <= not((layer0_outputs(3070)) and (layer0_outputs(3279)));
    layer1_outputs(2370) <= (layer0_outputs(6840)) or (layer0_outputs(3300));
    layer1_outputs(2371) <= (layer0_outputs(1317)) and (layer0_outputs(7031));
    layer1_outputs(2372) <= not((layer0_outputs(1522)) and (layer0_outputs(6679)));
    layer1_outputs(2373) <= not(layer0_outputs(3806));
    layer1_outputs(2374) <= not(layer0_outputs(62));
    layer1_outputs(2375) <= '0';
    layer1_outputs(2376) <= (layer0_outputs(6778)) and not (layer0_outputs(1878));
    layer1_outputs(2377) <= not(layer0_outputs(3207)) or (layer0_outputs(2289));
    layer1_outputs(2378) <= (layer0_outputs(1635)) and not (layer0_outputs(6069));
    layer1_outputs(2379) <= (layer0_outputs(2549)) and not (layer0_outputs(4613));
    layer1_outputs(2380) <= layer0_outputs(5118);
    layer1_outputs(2381) <= layer0_outputs(6571);
    layer1_outputs(2382) <= not((layer0_outputs(5547)) and (layer0_outputs(6929)));
    layer1_outputs(2383) <= not((layer0_outputs(826)) or (layer0_outputs(775)));
    layer1_outputs(2384) <= not((layer0_outputs(3242)) or (layer0_outputs(5145)));
    layer1_outputs(2385) <= not(layer0_outputs(2647)) or (layer0_outputs(776));
    layer1_outputs(2386) <= (layer0_outputs(3456)) or (layer0_outputs(912));
    layer1_outputs(2387) <= '0';
    layer1_outputs(2388) <= not(layer0_outputs(5006));
    layer1_outputs(2389) <= not(layer0_outputs(6794)) or (layer0_outputs(4053));
    layer1_outputs(2390) <= layer0_outputs(6041);
    layer1_outputs(2391) <= '1';
    layer1_outputs(2392) <= not(layer0_outputs(2503));
    layer1_outputs(2393) <= not((layer0_outputs(6970)) and (layer0_outputs(1144)));
    layer1_outputs(2394) <= (layer0_outputs(7206)) and not (layer0_outputs(6299));
    layer1_outputs(2395) <= not(layer0_outputs(999)) or (layer0_outputs(7566));
    layer1_outputs(2396) <= '0';
    layer1_outputs(2397) <= not(layer0_outputs(123));
    layer1_outputs(2398) <= '0';
    layer1_outputs(2399) <= layer0_outputs(137);
    layer1_outputs(2400) <= (layer0_outputs(6329)) and (layer0_outputs(5630));
    layer1_outputs(2401) <= not(layer0_outputs(3179));
    layer1_outputs(2402) <= not(layer0_outputs(5749));
    layer1_outputs(2403) <= layer0_outputs(6938);
    layer1_outputs(2404) <= not(layer0_outputs(895));
    layer1_outputs(2405) <= (layer0_outputs(703)) and (layer0_outputs(1115));
    layer1_outputs(2406) <= (layer0_outputs(176)) and not (layer0_outputs(1442));
    layer1_outputs(2407) <= not(layer0_outputs(982));
    layer1_outputs(2408) <= (layer0_outputs(4616)) and not (layer0_outputs(4367));
    layer1_outputs(2409) <= not(layer0_outputs(6048));
    layer1_outputs(2410) <= layer0_outputs(438);
    layer1_outputs(2411) <= not(layer0_outputs(916)) or (layer0_outputs(3817));
    layer1_outputs(2412) <= (layer0_outputs(197)) or (layer0_outputs(5632));
    layer1_outputs(2413) <= layer0_outputs(452);
    layer1_outputs(2414) <= (layer0_outputs(933)) and (layer0_outputs(5460));
    layer1_outputs(2415) <= (layer0_outputs(6965)) and not (layer0_outputs(4050));
    layer1_outputs(2416) <= not(layer0_outputs(2865));
    layer1_outputs(2417) <= (layer0_outputs(6820)) and not (layer0_outputs(2869));
    layer1_outputs(2418) <= (layer0_outputs(3809)) and not (layer0_outputs(2));
    layer1_outputs(2419) <= not(layer0_outputs(576));
    layer1_outputs(2420) <= not(layer0_outputs(4029));
    layer1_outputs(2421) <= not((layer0_outputs(6734)) xor (layer0_outputs(6341)));
    layer1_outputs(2422) <= (layer0_outputs(5379)) or (layer0_outputs(6131));
    layer1_outputs(2423) <= not(layer0_outputs(3110)) or (layer0_outputs(4765));
    layer1_outputs(2424) <= not(layer0_outputs(1216));
    layer1_outputs(2425) <= not(layer0_outputs(6315));
    layer1_outputs(2426) <= not((layer0_outputs(6783)) and (layer0_outputs(4523)));
    layer1_outputs(2427) <= layer0_outputs(5809);
    layer1_outputs(2428) <= not((layer0_outputs(3104)) or (layer0_outputs(6593)));
    layer1_outputs(2429) <= '1';
    layer1_outputs(2430) <= (layer0_outputs(6567)) and not (layer0_outputs(1744));
    layer1_outputs(2431) <= (layer0_outputs(2431)) and not (layer0_outputs(7330));
    layer1_outputs(2432) <= '1';
    layer1_outputs(2433) <= (layer0_outputs(3615)) and (layer0_outputs(4482));
    layer1_outputs(2434) <= '0';
    layer1_outputs(2435) <= not(layer0_outputs(6865));
    layer1_outputs(2436) <= not(layer0_outputs(1341));
    layer1_outputs(2437) <= not(layer0_outputs(5555));
    layer1_outputs(2438) <= not(layer0_outputs(296)) or (layer0_outputs(5840));
    layer1_outputs(2439) <= not(layer0_outputs(3697));
    layer1_outputs(2440) <= (layer0_outputs(4380)) and (layer0_outputs(5865));
    layer1_outputs(2441) <= layer0_outputs(2102);
    layer1_outputs(2442) <= not((layer0_outputs(5852)) or (layer0_outputs(6599)));
    layer1_outputs(2443) <= not(layer0_outputs(5406)) or (layer0_outputs(4375));
    layer1_outputs(2444) <= layer0_outputs(1414);
    layer1_outputs(2445) <= layer0_outputs(4238);
    layer1_outputs(2446) <= not(layer0_outputs(5558));
    layer1_outputs(2447) <= not(layer0_outputs(6907));
    layer1_outputs(2448) <= not((layer0_outputs(4100)) and (layer0_outputs(1014)));
    layer1_outputs(2449) <= not((layer0_outputs(1728)) and (layer0_outputs(7025)));
    layer1_outputs(2450) <= layer0_outputs(1376);
    layer1_outputs(2451) <= layer0_outputs(1053);
    layer1_outputs(2452) <= layer0_outputs(726);
    layer1_outputs(2453) <= not(layer0_outputs(4487));
    layer1_outputs(2454) <= '0';
    layer1_outputs(2455) <= (layer0_outputs(7573)) and not (layer0_outputs(2586));
    layer1_outputs(2456) <= '0';
    layer1_outputs(2457) <= (layer0_outputs(2042)) and not (layer0_outputs(1676));
    layer1_outputs(2458) <= (layer0_outputs(7228)) and not (layer0_outputs(6552));
    layer1_outputs(2459) <= (layer0_outputs(3779)) and not (layer0_outputs(343));
    layer1_outputs(2460) <= not(layer0_outputs(3857));
    layer1_outputs(2461) <= layer0_outputs(1367);
    layer1_outputs(2462) <= not((layer0_outputs(5734)) or (layer0_outputs(5081)));
    layer1_outputs(2463) <= (layer0_outputs(6577)) and not (layer0_outputs(5614));
    layer1_outputs(2464) <= not((layer0_outputs(2698)) or (layer0_outputs(1793)));
    layer1_outputs(2465) <= not(layer0_outputs(3920));
    layer1_outputs(2466) <= (layer0_outputs(294)) and not (layer0_outputs(4369));
    layer1_outputs(2467) <= layer0_outputs(7675);
    layer1_outputs(2468) <= layer0_outputs(1784);
    layer1_outputs(2469) <= (layer0_outputs(3556)) and (layer0_outputs(2708));
    layer1_outputs(2470) <= layer0_outputs(4195);
    layer1_outputs(2471) <= not((layer0_outputs(6192)) and (layer0_outputs(4517)));
    layer1_outputs(2472) <= layer0_outputs(759);
    layer1_outputs(2473) <= '0';
    layer1_outputs(2474) <= '1';
    layer1_outputs(2475) <= (layer0_outputs(3323)) or (layer0_outputs(4257));
    layer1_outputs(2476) <= not((layer0_outputs(5635)) or (layer0_outputs(3480)));
    layer1_outputs(2477) <= '0';
    layer1_outputs(2478) <= (layer0_outputs(6796)) and not (layer0_outputs(6622));
    layer1_outputs(2479) <= '1';
    layer1_outputs(2480) <= not((layer0_outputs(4211)) and (layer0_outputs(419)));
    layer1_outputs(2481) <= layer0_outputs(5642);
    layer1_outputs(2482) <= not(layer0_outputs(7150));
    layer1_outputs(2483) <= not((layer0_outputs(3744)) and (layer0_outputs(5690)));
    layer1_outputs(2484) <= not((layer0_outputs(3533)) and (layer0_outputs(1250)));
    layer1_outputs(2485) <= (layer0_outputs(452)) and not (layer0_outputs(2536));
    layer1_outputs(2486) <= (layer0_outputs(1897)) and not (layer0_outputs(661));
    layer1_outputs(2487) <= not((layer0_outputs(5880)) or (layer0_outputs(5143)));
    layer1_outputs(2488) <= (layer0_outputs(1294)) xor (layer0_outputs(1003));
    layer1_outputs(2489) <= (layer0_outputs(6464)) and not (layer0_outputs(675));
    layer1_outputs(2490) <= not(layer0_outputs(3523));
    layer1_outputs(2491) <= '1';
    layer1_outputs(2492) <= (layer0_outputs(6423)) and not (layer0_outputs(5193));
    layer1_outputs(2493) <= not(layer0_outputs(1690));
    layer1_outputs(2494) <= layer0_outputs(1233);
    layer1_outputs(2495) <= not((layer0_outputs(206)) or (layer0_outputs(4020)));
    layer1_outputs(2496) <= not(layer0_outputs(399));
    layer1_outputs(2497) <= not(layer0_outputs(2105)) or (layer0_outputs(2060));
    layer1_outputs(2498) <= not(layer0_outputs(7112)) or (layer0_outputs(1828));
    layer1_outputs(2499) <= not((layer0_outputs(6576)) and (layer0_outputs(707)));
    layer1_outputs(2500) <= (layer0_outputs(1598)) and not (layer0_outputs(13));
    layer1_outputs(2501) <= not((layer0_outputs(3397)) xor (layer0_outputs(7213)));
    layer1_outputs(2502) <= '0';
    layer1_outputs(2503) <= not((layer0_outputs(4011)) and (layer0_outputs(538)));
    layer1_outputs(2504) <= (layer0_outputs(6169)) and (layer0_outputs(1276));
    layer1_outputs(2505) <= not(layer0_outputs(3067));
    layer1_outputs(2506) <= not(layer0_outputs(4295));
    layer1_outputs(2507) <= layer0_outputs(1477);
    layer1_outputs(2508) <= (layer0_outputs(3221)) and not (layer0_outputs(984));
    layer1_outputs(2509) <= not(layer0_outputs(7040));
    layer1_outputs(2510) <= (layer0_outputs(616)) or (layer0_outputs(1508));
    layer1_outputs(2511) <= layer0_outputs(5620);
    layer1_outputs(2512) <= not(layer0_outputs(861));
    layer1_outputs(2513) <= not((layer0_outputs(6606)) and (layer0_outputs(497)));
    layer1_outputs(2514) <= (layer0_outputs(5368)) and not (layer0_outputs(2632));
    layer1_outputs(2515) <= '0';
    layer1_outputs(2516) <= not(layer0_outputs(5824)) or (layer0_outputs(5726));
    layer1_outputs(2517) <= (layer0_outputs(2192)) and not (layer0_outputs(3812));
    layer1_outputs(2518) <= not(layer0_outputs(5284)) or (layer0_outputs(2236));
    layer1_outputs(2519) <= not(layer0_outputs(1044)) or (layer0_outputs(539));
    layer1_outputs(2520) <= (layer0_outputs(4598)) and not (layer0_outputs(796));
    layer1_outputs(2521) <= '0';
    layer1_outputs(2522) <= (layer0_outputs(4103)) and not (layer0_outputs(6226));
    layer1_outputs(2523) <= not((layer0_outputs(3246)) or (layer0_outputs(3244)));
    layer1_outputs(2524) <= (layer0_outputs(4985)) and not (layer0_outputs(5497));
    layer1_outputs(2525) <= (layer0_outputs(2725)) and (layer0_outputs(7110));
    layer1_outputs(2526) <= (layer0_outputs(6936)) and not (layer0_outputs(1499));
    layer1_outputs(2527) <= not(layer0_outputs(7026)) or (layer0_outputs(2402));
    layer1_outputs(2528) <= (layer0_outputs(3644)) and not (layer0_outputs(5321));
    layer1_outputs(2529) <= layer0_outputs(5170);
    layer1_outputs(2530) <= not((layer0_outputs(835)) or (layer0_outputs(1755)));
    layer1_outputs(2531) <= '0';
    layer1_outputs(2532) <= not((layer0_outputs(1753)) or (layer0_outputs(6734)));
    layer1_outputs(2533) <= not((layer0_outputs(7461)) or (layer0_outputs(7617)));
    layer1_outputs(2534) <= (layer0_outputs(7410)) and not (layer0_outputs(3759));
    layer1_outputs(2535) <= (layer0_outputs(2491)) and not (layer0_outputs(4074));
    layer1_outputs(2536) <= layer0_outputs(1478);
    layer1_outputs(2537) <= layer0_outputs(180);
    layer1_outputs(2538) <= layer0_outputs(7371);
    layer1_outputs(2539) <= (layer0_outputs(51)) xor (layer0_outputs(6625));
    layer1_outputs(2540) <= layer0_outputs(2516);
    layer1_outputs(2541) <= '0';
    layer1_outputs(2542) <= (layer0_outputs(4565)) and (layer0_outputs(6537));
    layer1_outputs(2543) <= (layer0_outputs(7282)) and not (layer0_outputs(6648));
    layer1_outputs(2544) <= not((layer0_outputs(4981)) or (layer0_outputs(2127)));
    layer1_outputs(2545) <= (layer0_outputs(6834)) or (layer0_outputs(2));
    layer1_outputs(2546) <= '0';
    layer1_outputs(2547) <= (layer0_outputs(1385)) and (layer0_outputs(3413));
    layer1_outputs(2548) <= not(layer0_outputs(635));
    layer1_outputs(2549) <= not(layer0_outputs(341)) or (layer0_outputs(7274));
    layer1_outputs(2550) <= '0';
    layer1_outputs(2551) <= (layer0_outputs(3993)) and not (layer0_outputs(7023));
    layer1_outputs(2552) <= not(layer0_outputs(1543));
    layer1_outputs(2553) <= (layer0_outputs(7044)) and not (layer0_outputs(1073));
    layer1_outputs(2554) <= (layer0_outputs(6864)) and not (layer0_outputs(6739));
    layer1_outputs(2555) <= not(layer0_outputs(6037)) or (layer0_outputs(5533));
    layer1_outputs(2556) <= not(layer0_outputs(6693));
    layer1_outputs(2557) <= (layer0_outputs(5455)) and (layer0_outputs(2324));
    layer1_outputs(2558) <= not(layer0_outputs(6141));
    layer1_outputs(2559) <= (layer0_outputs(3711)) or (layer0_outputs(6853));
    layer1_outputs(2560) <= layer0_outputs(3622);
    layer1_outputs(2561) <= (layer0_outputs(4190)) and not (layer0_outputs(2587));
    layer1_outputs(2562) <= not(layer0_outputs(3347)) or (layer0_outputs(6954));
    layer1_outputs(2563) <= not(layer0_outputs(2555)) or (layer0_outputs(5201));
    layer1_outputs(2564) <= '0';
    layer1_outputs(2565) <= not(layer0_outputs(2083)) or (layer0_outputs(1136));
    layer1_outputs(2566) <= layer0_outputs(1903);
    layer1_outputs(2567) <= (layer0_outputs(647)) and not (layer0_outputs(2138));
    layer1_outputs(2568) <= (layer0_outputs(1794)) or (layer0_outputs(6603));
    layer1_outputs(2569) <= (layer0_outputs(7436)) or (layer0_outputs(2053));
    layer1_outputs(2570) <= '1';
    layer1_outputs(2571) <= (layer0_outputs(6272)) xor (layer0_outputs(3811));
    layer1_outputs(2572) <= (layer0_outputs(2415)) and not (layer0_outputs(4090));
    layer1_outputs(2573) <= (layer0_outputs(6762)) and not (layer0_outputs(7038));
    layer1_outputs(2574) <= not(layer0_outputs(280)) or (layer0_outputs(3436));
    layer1_outputs(2575) <= (layer0_outputs(874)) and (layer0_outputs(7610));
    layer1_outputs(2576) <= not(layer0_outputs(6838));
    layer1_outputs(2577) <= not(layer0_outputs(2201)) or (layer0_outputs(2726));
    layer1_outputs(2578) <= not(layer0_outputs(4146)) or (layer0_outputs(264));
    layer1_outputs(2579) <= (layer0_outputs(6222)) and not (layer0_outputs(7268));
    layer1_outputs(2580) <= not(layer0_outputs(2069)) or (layer0_outputs(4091));
    layer1_outputs(2581) <= (layer0_outputs(2754)) xor (layer0_outputs(3128));
    layer1_outputs(2582) <= not(layer0_outputs(1724)) or (layer0_outputs(5974));
    layer1_outputs(2583) <= not(layer0_outputs(4005));
    layer1_outputs(2584) <= (layer0_outputs(50)) and not (layer0_outputs(6410));
    layer1_outputs(2585) <= not(layer0_outputs(403)) or (layer0_outputs(7063));
    layer1_outputs(2586) <= layer0_outputs(6995);
    layer1_outputs(2587) <= (layer0_outputs(4403)) and not (layer0_outputs(1512));
    layer1_outputs(2588) <= not((layer0_outputs(5294)) or (layer0_outputs(1142)));
    layer1_outputs(2589) <= (layer0_outputs(2381)) and not (layer0_outputs(2883));
    layer1_outputs(2590) <= not((layer0_outputs(5613)) and (layer0_outputs(3670)));
    layer1_outputs(2591) <= not(layer0_outputs(3289)) or (layer0_outputs(4064));
    layer1_outputs(2592) <= not(layer0_outputs(1058));
    layer1_outputs(2593) <= not(layer0_outputs(7640)) or (layer0_outputs(446));
    layer1_outputs(2594) <= '0';
    layer1_outputs(2595) <= (layer0_outputs(5200)) xor (layer0_outputs(4537));
    layer1_outputs(2596) <= not(layer0_outputs(6411));
    layer1_outputs(2597) <= layer0_outputs(6847);
    layer1_outputs(2598) <= not(layer0_outputs(1460)) or (layer0_outputs(6853));
    layer1_outputs(2599) <= layer0_outputs(3968);
    layer1_outputs(2600) <= layer0_outputs(2634);
    layer1_outputs(2601) <= (layer0_outputs(4600)) and not (layer0_outputs(7042));
    layer1_outputs(2602) <= not((layer0_outputs(3380)) or (layer0_outputs(5212)));
    layer1_outputs(2603) <= not(layer0_outputs(7360)) or (layer0_outputs(4698));
    layer1_outputs(2604) <= '1';
    layer1_outputs(2605) <= (layer0_outputs(6984)) and (layer0_outputs(6543));
    layer1_outputs(2606) <= not(layer0_outputs(2580)) or (layer0_outputs(565));
    layer1_outputs(2607) <= (layer0_outputs(4320)) and not (layer0_outputs(4207));
    layer1_outputs(2608) <= (layer0_outputs(1697)) and not (layer0_outputs(7536));
    layer1_outputs(2609) <= (layer0_outputs(6823)) and not (layer0_outputs(1089));
    layer1_outputs(2610) <= (layer0_outputs(3210)) xor (layer0_outputs(2589));
    layer1_outputs(2611) <= (layer0_outputs(1166)) xor (layer0_outputs(4019));
    layer1_outputs(2612) <= (layer0_outputs(3214)) and not (layer0_outputs(3760));
    layer1_outputs(2613) <= not((layer0_outputs(6330)) xor (layer0_outputs(432)));
    layer1_outputs(2614) <= layer0_outputs(4759);
    layer1_outputs(2615) <= layer0_outputs(3312);
    layer1_outputs(2616) <= not(layer0_outputs(3687));
    layer1_outputs(2617) <= not(layer0_outputs(1441));
    layer1_outputs(2618) <= not(layer0_outputs(4098)) or (layer0_outputs(614));
    layer1_outputs(2619) <= '0';
    layer1_outputs(2620) <= '0';
    layer1_outputs(2621) <= layer0_outputs(1644);
    layer1_outputs(2622) <= (layer0_outputs(5647)) and (layer0_outputs(2539));
    layer1_outputs(2623) <= not(layer0_outputs(4769)) or (layer0_outputs(3037));
    layer1_outputs(2624) <= not(layer0_outputs(7214)) or (layer0_outputs(6043));
    layer1_outputs(2625) <= layer0_outputs(6482);
    layer1_outputs(2626) <= (layer0_outputs(4947)) and not (layer0_outputs(3534));
    layer1_outputs(2627) <= (layer0_outputs(1200)) or (layer0_outputs(5272));
    layer1_outputs(2628) <= '1';
    layer1_outputs(2629) <= not(layer0_outputs(1000));
    layer1_outputs(2630) <= not(layer0_outputs(6044));
    layer1_outputs(2631) <= layer0_outputs(4420);
    layer1_outputs(2632) <= not(layer0_outputs(3576));
    layer1_outputs(2633) <= (layer0_outputs(2659)) or (layer0_outputs(3011));
    layer1_outputs(2634) <= layer0_outputs(5470);
    layer1_outputs(2635) <= (layer0_outputs(5211)) xor (layer0_outputs(6277));
    layer1_outputs(2636) <= (layer0_outputs(7200)) and not (layer0_outputs(1915));
    layer1_outputs(2637) <= not(layer0_outputs(4237));
    layer1_outputs(2638) <= (layer0_outputs(5414)) and not (layer0_outputs(709));
    layer1_outputs(2639) <= layer0_outputs(1859);
    layer1_outputs(2640) <= '1';
    layer1_outputs(2641) <= not(layer0_outputs(355)) or (layer0_outputs(4547));
    layer1_outputs(2642) <= not((layer0_outputs(1368)) and (layer0_outputs(5626)));
    layer1_outputs(2643) <= (layer0_outputs(6462)) xor (layer0_outputs(3482));
    layer1_outputs(2644) <= not(layer0_outputs(1335)) or (layer0_outputs(5304));
    layer1_outputs(2645) <= not(layer0_outputs(7231));
    layer1_outputs(2646) <= layer0_outputs(5023);
    layer1_outputs(2647) <= '1';
    layer1_outputs(2648) <= not(layer0_outputs(4326));
    layer1_outputs(2649) <= '1';
    layer1_outputs(2650) <= not(layer0_outputs(3104)) or (layer0_outputs(7243));
    layer1_outputs(2651) <= (layer0_outputs(156)) and (layer0_outputs(3792));
    layer1_outputs(2652) <= not(layer0_outputs(7481));
    layer1_outputs(2653) <= not((layer0_outputs(4816)) and (layer0_outputs(2401)));
    layer1_outputs(2654) <= not((layer0_outputs(3220)) and (layer0_outputs(4007)));
    layer1_outputs(2655) <= not((layer0_outputs(5570)) or (layer0_outputs(2596)));
    layer1_outputs(2656) <= layer0_outputs(6349);
    layer1_outputs(2657) <= not(layer0_outputs(3824));
    layer1_outputs(2658) <= (layer0_outputs(274)) and (layer0_outputs(715));
    layer1_outputs(2659) <= layer0_outputs(1496);
    layer1_outputs(2660) <= '1';
    layer1_outputs(2661) <= '1';
    layer1_outputs(2662) <= (layer0_outputs(710)) and (layer0_outputs(3944));
    layer1_outputs(2663) <= layer0_outputs(5559);
    layer1_outputs(2664) <= not(layer0_outputs(5075)) or (layer0_outputs(671));
    layer1_outputs(2665) <= not((layer0_outputs(5428)) and (layer0_outputs(6622)));
    layer1_outputs(2666) <= not(layer0_outputs(6817));
    layer1_outputs(2667) <= not((layer0_outputs(1861)) and (layer0_outputs(4396)));
    layer1_outputs(2668) <= not((layer0_outputs(5145)) or (layer0_outputs(2656)));
    layer1_outputs(2669) <= (layer0_outputs(1445)) and (layer0_outputs(6260));
    layer1_outputs(2670) <= layer0_outputs(7607);
    layer1_outputs(2671) <= layer0_outputs(2004);
    layer1_outputs(2672) <= layer0_outputs(5117);
    layer1_outputs(2673) <= not(layer0_outputs(4103));
    layer1_outputs(2674) <= not(layer0_outputs(4767));
    layer1_outputs(2675) <= layer0_outputs(2975);
    layer1_outputs(2676) <= not(layer0_outputs(2221));
    layer1_outputs(2677) <= '1';
    layer1_outputs(2678) <= not((layer0_outputs(5072)) xor (layer0_outputs(4444)));
    layer1_outputs(2679) <= '0';
    layer1_outputs(2680) <= (layer0_outputs(2030)) and (layer0_outputs(5722));
    layer1_outputs(2681) <= '0';
    layer1_outputs(2682) <= '1';
    layer1_outputs(2683) <= not(layer0_outputs(4761));
    layer1_outputs(2684) <= not(layer0_outputs(5451));
    layer1_outputs(2685) <= (layer0_outputs(3465)) or (layer0_outputs(4685));
    layer1_outputs(2686) <= not(layer0_outputs(4276)) or (layer0_outputs(2032));
    layer1_outputs(2687) <= not(layer0_outputs(3509)) or (layer0_outputs(7386));
    layer1_outputs(2688) <= (layer0_outputs(2188)) or (layer0_outputs(2433));
    layer1_outputs(2689) <= layer0_outputs(1596);
    layer1_outputs(2690) <= not(layer0_outputs(4274));
    layer1_outputs(2691) <= not(layer0_outputs(4555));
    layer1_outputs(2692) <= not(layer0_outputs(3594));
    layer1_outputs(2693) <= '0';
    layer1_outputs(2694) <= layer0_outputs(5552);
    layer1_outputs(2695) <= not(layer0_outputs(1920)) or (layer0_outputs(5205));
    layer1_outputs(2696) <= not((layer0_outputs(6635)) or (layer0_outputs(3227)));
    layer1_outputs(2697) <= layer0_outputs(6601);
    layer1_outputs(2698) <= layer0_outputs(2803);
    layer1_outputs(2699) <= not(layer0_outputs(5029));
    layer1_outputs(2700) <= not(layer0_outputs(3751));
    layer1_outputs(2701) <= not(layer0_outputs(658));
    layer1_outputs(2702) <= (layer0_outputs(3399)) and (layer0_outputs(331));
    layer1_outputs(2703) <= '1';
    layer1_outputs(2704) <= '1';
    layer1_outputs(2705) <= layer0_outputs(1418);
    layer1_outputs(2706) <= '0';
    layer1_outputs(2707) <= not(layer0_outputs(6496)) or (layer0_outputs(2194));
    layer1_outputs(2708) <= not(layer0_outputs(3351)) or (layer0_outputs(5126));
    layer1_outputs(2709) <= (layer0_outputs(5868)) and (layer0_outputs(4724));
    layer1_outputs(2710) <= layer0_outputs(7531);
    layer1_outputs(2711) <= layer0_outputs(336);
    layer1_outputs(2712) <= not(layer0_outputs(4236));
    layer1_outputs(2713) <= not(layer0_outputs(6900));
    layer1_outputs(2714) <= '1';
    layer1_outputs(2715) <= not((layer0_outputs(680)) or (layer0_outputs(1967)));
    layer1_outputs(2716) <= (layer0_outputs(4329)) and not (layer0_outputs(7404));
    layer1_outputs(2717) <= not((layer0_outputs(1990)) or (layer0_outputs(5058)));
    layer1_outputs(2718) <= not(layer0_outputs(714)) or (layer0_outputs(2148));
    layer1_outputs(2719) <= '0';
    layer1_outputs(2720) <= layer0_outputs(1157);
    layer1_outputs(2721) <= not(layer0_outputs(544));
    layer1_outputs(2722) <= layer0_outputs(3761);
    layer1_outputs(2723) <= (layer0_outputs(283)) or (layer0_outputs(7442));
    layer1_outputs(2724) <= not(layer0_outputs(492));
    layer1_outputs(2725) <= not(layer0_outputs(1203));
    layer1_outputs(2726) <= '1';
    layer1_outputs(2727) <= (layer0_outputs(3583)) and not (layer0_outputs(2215));
    layer1_outputs(2728) <= not(layer0_outputs(1108)) or (layer0_outputs(3008));
    layer1_outputs(2729) <= (layer0_outputs(1132)) and not (layer0_outputs(2436));
    layer1_outputs(2730) <= (layer0_outputs(859)) and not (layer0_outputs(375));
    layer1_outputs(2731) <= not(layer0_outputs(1169)) or (layer0_outputs(1056));
    layer1_outputs(2732) <= not(layer0_outputs(6238));
    layer1_outputs(2733) <= not((layer0_outputs(809)) or (layer0_outputs(4807)));
    layer1_outputs(2734) <= '0';
    layer1_outputs(2735) <= '0';
    layer1_outputs(2736) <= not(layer0_outputs(7412));
    layer1_outputs(2737) <= (layer0_outputs(4303)) and (layer0_outputs(6360));
    layer1_outputs(2738) <= layer0_outputs(5804);
    layer1_outputs(2739) <= layer0_outputs(5204);
    layer1_outputs(2740) <= (layer0_outputs(4294)) and (layer0_outputs(4687));
    layer1_outputs(2741) <= not(layer0_outputs(2296));
    layer1_outputs(2742) <= (layer0_outputs(7652)) and not (layer0_outputs(104));
    layer1_outputs(2743) <= (layer0_outputs(3286)) and (layer0_outputs(7541));
    layer1_outputs(2744) <= not((layer0_outputs(769)) or (layer0_outputs(1980)));
    layer1_outputs(2745) <= not(layer0_outputs(5721));
    layer1_outputs(2746) <= not(layer0_outputs(910)) or (layer0_outputs(7552));
    layer1_outputs(2747) <= layer0_outputs(588);
    layer1_outputs(2748) <= (layer0_outputs(3957)) xor (layer0_outputs(3559));
    layer1_outputs(2749) <= (layer0_outputs(4857)) and not (layer0_outputs(6848));
    layer1_outputs(2750) <= (layer0_outputs(3749)) xor (layer0_outputs(2334));
    layer1_outputs(2751) <= not(layer0_outputs(4193));
    layer1_outputs(2752) <= not(layer0_outputs(5514)) or (layer0_outputs(6691));
    layer1_outputs(2753) <= (layer0_outputs(2692)) and not (layer0_outputs(3819));
    layer1_outputs(2754) <= (layer0_outputs(1303)) and not (layer0_outputs(4270));
    layer1_outputs(2755) <= not(layer0_outputs(5237)) or (layer0_outputs(1440));
    layer1_outputs(2756) <= layer0_outputs(4551);
    layer1_outputs(2757) <= not((layer0_outputs(4524)) or (layer0_outputs(2288)));
    layer1_outputs(2758) <= (layer0_outputs(2853)) or (layer0_outputs(3852));
    layer1_outputs(2759) <= '0';
    layer1_outputs(2760) <= not(layer0_outputs(5891));
    layer1_outputs(2761) <= layer0_outputs(6033);
    layer1_outputs(2762) <= not(layer0_outputs(5195));
    layer1_outputs(2763) <= '0';
    layer1_outputs(2764) <= not(layer0_outputs(808));
    layer1_outputs(2765) <= not(layer0_outputs(1155)) or (layer0_outputs(4142));
    layer1_outputs(2766) <= not((layer0_outputs(6704)) or (layer0_outputs(1089)));
    layer1_outputs(2767) <= (layer0_outputs(1502)) and (layer0_outputs(1630));
    layer1_outputs(2768) <= not(layer0_outputs(985)) or (layer0_outputs(1098));
    layer1_outputs(2769) <= (layer0_outputs(5161)) and (layer0_outputs(3949));
    layer1_outputs(2770) <= (layer0_outputs(7502)) or (layer0_outputs(6753));
    layer1_outputs(2771) <= layer0_outputs(5821);
    layer1_outputs(2772) <= not(layer0_outputs(6659));
    layer1_outputs(2773) <= '0';
    layer1_outputs(2774) <= layer0_outputs(4706);
    layer1_outputs(2775) <= not(layer0_outputs(2801)) or (layer0_outputs(3978));
    layer1_outputs(2776) <= (layer0_outputs(2987)) or (layer0_outputs(1721));
    layer1_outputs(2777) <= not((layer0_outputs(7087)) xor (layer0_outputs(3875)));
    layer1_outputs(2778) <= not(layer0_outputs(2077)) or (layer0_outputs(3786));
    layer1_outputs(2779) <= layer0_outputs(412);
    layer1_outputs(2780) <= layer0_outputs(1841);
    layer1_outputs(2781) <= (layer0_outputs(3562)) and (layer0_outputs(3397));
    layer1_outputs(2782) <= (layer0_outputs(4829)) and not (layer0_outputs(1581));
    layer1_outputs(2783) <= not(layer0_outputs(2458));
    layer1_outputs(2784) <= layer0_outputs(1769);
    layer1_outputs(2785) <= '1';
    layer1_outputs(2786) <= not(layer0_outputs(1932));
    layer1_outputs(2787) <= not(layer0_outputs(637)) or (layer0_outputs(1743));
    layer1_outputs(2788) <= (layer0_outputs(891)) or (layer0_outputs(1024));
    layer1_outputs(2789) <= (layer0_outputs(2058)) or (layer0_outputs(880));
    layer1_outputs(2790) <= not(layer0_outputs(2304));
    layer1_outputs(2791) <= (layer0_outputs(4146)) and (layer0_outputs(6814));
    layer1_outputs(2792) <= (layer0_outputs(6815)) and not (layer0_outputs(6779));
    layer1_outputs(2793) <= not((layer0_outputs(3883)) or (layer0_outputs(2734)));
    layer1_outputs(2794) <= layer0_outputs(2973);
    layer1_outputs(2795) <= layer0_outputs(4649);
    layer1_outputs(2796) <= (layer0_outputs(1116)) and not (layer0_outputs(3141));
    layer1_outputs(2797) <= not(layer0_outputs(3052)) or (layer0_outputs(2627));
    layer1_outputs(2798) <= not(layer0_outputs(4413)) or (layer0_outputs(2164));
    layer1_outputs(2799) <= layer0_outputs(4451);
    layer1_outputs(2800) <= layer0_outputs(1810);
    layer1_outputs(2801) <= not(layer0_outputs(550)) or (layer0_outputs(6316));
    layer1_outputs(2802) <= (layer0_outputs(1258)) and not (layer0_outputs(7335));
    layer1_outputs(2803) <= not(layer0_outputs(1749)) or (layer0_outputs(1838));
    layer1_outputs(2804) <= layer0_outputs(1451);
    layer1_outputs(2805) <= not((layer0_outputs(626)) or (layer0_outputs(5078)));
    layer1_outputs(2806) <= not(layer0_outputs(1365)) or (layer0_outputs(1585));
    layer1_outputs(2807) <= not((layer0_outputs(2825)) and (layer0_outputs(590)));
    layer1_outputs(2808) <= not(layer0_outputs(2794));
    layer1_outputs(2809) <= not(layer0_outputs(2539));
    layer1_outputs(2810) <= (layer0_outputs(2612)) and not (layer0_outputs(4934));
    layer1_outputs(2811) <= not((layer0_outputs(2943)) or (layer0_outputs(7490)));
    layer1_outputs(2812) <= not((layer0_outputs(3797)) and (layer0_outputs(6049)));
    layer1_outputs(2813) <= (layer0_outputs(7101)) and not (layer0_outputs(1862));
    layer1_outputs(2814) <= not((layer0_outputs(1410)) or (layer0_outputs(7610)));
    layer1_outputs(2815) <= not((layer0_outputs(5815)) or (layer0_outputs(1212)));
    layer1_outputs(2816) <= layer0_outputs(6257);
    layer1_outputs(2817) <= '0';
    layer1_outputs(2818) <= (layer0_outputs(4558)) and (layer0_outputs(1041));
    layer1_outputs(2819) <= not(layer0_outputs(6472)) or (layer0_outputs(6963));
    layer1_outputs(2820) <= layer0_outputs(4871);
    layer1_outputs(2821) <= layer0_outputs(7313);
    layer1_outputs(2822) <= (layer0_outputs(7190)) or (layer0_outputs(2646));
    layer1_outputs(2823) <= (layer0_outputs(3499)) or (layer0_outputs(3375));
    layer1_outputs(2824) <= not((layer0_outputs(3878)) or (layer0_outputs(5785)));
    layer1_outputs(2825) <= not(layer0_outputs(6918));
    layer1_outputs(2826) <= not(layer0_outputs(1155));
    layer1_outputs(2827) <= '0';
    layer1_outputs(2828) <= layer0_outputs(3410);
    layer1_outputs(2829) <= '0';
    layer1_outputs(2830) <= not(layer0_outputs(4150)) or (layer0_outputs(396));
    layer1_outputs(2831) <= not(layer0_outputs(6050));
    layer1_outputs(2832) <= layer0_outputs(6977);
    layer1_outputs(2833) <= not(layer0_outputs(7131)) or (layer0_outputs(3115));
    layer1_outputs(2834) <= '1';
    layer1_outputs(2835) <= (layer0_outputs(4748)) and not (layer0_outputs(2577));
    layer1_outputs(2836) <= (layer0_outputs(5817)) and not (layer0_outputs(5969));
    layer1_outputs(2837) <= layer0_outputs(2993);
    layer1_outputs(2838) <= layer0_outputs(6046);
    layer1_outputs(2839) <= not(layer0_outputs(1137));
    layer1_outputs(2840) <= layer0_outputs(3943);
    layer1_outputs(2841) <= layer0_outputs(607);
    layer1_outputs(2842) <= '0';
    layer1_outputs(2843) <= (layer0_outputs(6564)) and (layer0_outputs(7346));
    layer1_outputs(2844) <= not(layer0_outputs(1276));
    layer1_outputs(2845) <= layer0_outputs(4729);
    layer1_outputs(2846) <= not(layer0_outputs(5716)) or (layer0_outputs(6047));
    layer1_outputs(2847) <= (layer0_outputs(455)) and not (layer0_outputs(5775));
    layer1_outputs(2848) <= not((layer0_outputs(479)) or (layer0_outputs(901)));
    layer1_outputs(2849) <= not(layer0_outputs(3269));
    layer1_outputs(2850) <= layer0_outputs(7332);
    layer1_outputs(2851) <= (layer0_outputs(3634)) and not (layer0_outputs(5236));
    layer1_outputs(2852) <= not(layer0_outputs(5016));
    layer1_outputs(2853) <= not(layer0_outputs(4345));
    layer1_outputs(2854) <= not(layer0_outputs(6888));
    layer1_outputs(2855) <= (layer0_outputs(4650)) and not (layer0_outputs(3884));
    layer1_outputs(2856) <= (layer0_outputs(3721)) or (layer0_outputs(2410));
    layer1_outputs(2857) <= (layer0_outputs(7524)) or (layer0_outputs(779));
    layer1_outputs(2858) <= (layer0_outputs(4367)) and not (layer0_outputs(1152));
    layer1_outputs(2859) <= (layer0_outputs(6867)) or (layer0_outputs(2475));
    layer1_outputs(2860) <= not((layer0_outputs(1509)) and (layer0_outputs(863)));
    layer1_outputs(2861) <= not((layer0_outputs(3235)) or (layer0_outputs(4253)));
    layer1_outputs(2862) <= (layer0_outputs(1955)) or (layer0_outputs(6794));
    layer1_outputs(2863) <= (layer0_outputs(5271)) and not (layer0_outputs(2656));
    layer1_outputs(2864) <= (layer0_outputs(4845)) and (layer0_outputs(1431));
    layer1_outputs(2865) <= (layer0_outputs(5080)) and not (layer0_outputs(7220));
    layer1_outputs(2866) <= '1';
    layer1_outputs(2867) <= '0';
    layer1_outputs(2868) <= layer0_outputs(1565);
    layer1_outputs(2869) <= not(layer0_outputs(2967));
    layer1_outputs(2870) <= not(layer0_outputs(574)) or (layer0_outputs(1310));
    layer1_outputs(2871) <= (layer0_outputs(885)) and not (layer0_outputs(5748));
    layer1_outputs(2872) <= not((layer0_outputs(2089)) and (layer0_outputs(3322)));
    layer1_outputs(2873) <= (layer0_outputs(1670)) xor (layer0_outputs(4021));
    layer1_outputs(2874) <= '0';
    layer1_outputs(2875) <= (layer0_outputs(4111)) and not (layer0_outputs(6861));
    layer1_outputs(2876) <= not(layer0_outputs(3385));
    layer1_outputs(2877) <= '1';
    layer1_outputs(2878) <= not(layer0_outputs(3461));
    layer1_outputs(2879) <= not(layer0_outputs(444));
    layer1_outputs(2880) <= not(layer0_outputs(6288));
    layer1_outputs(2881) <= (layer0_outputs(812)) or (layer0_outputs(7136));
    layer1_outputs(2882) <= layer0_outputs(2200);
    layer1_outputs(2883) <= layer0_outputs(1206);
    layer1_outputs(2884) <= layer0_outputs(2015);
    layer1_outputs(2885) <= not(layer0_outputs(6461));
    layer1_outputs(2886) <= not((layer0_outputs(5102)) and (layer0_outputs(1017)));
    layer1_outputs(2887) <= '0';
    layer1_outputs(2888) <= (layer0_outputs(2450)) and not (layer0_outputs(1566));
    layer1_outputs(2889) <= (layer0_outputs(3280)) and (layer0_outputs(6389));
    layer1_outputs(2890) <= '1';
    layer1_outputs(2891) <= (layer0_outputs(4855)) or (layer0_outputs(3580));
    layer1_outputs(2892) <= layer0_outputs(3006);
    layer1_outputs(2893) <= (layer0_outputs(6845)) or (layer0_outputs(3646));
    layer1_outputs(2894) <= (layer0_outputs(5199)) and not (layer0_outputs(7177));
    layer1_outputs(2895) <= not(layer0_outputs(1767));
    layer1_outputs(2896) <= not(layer0_outputs(1283)) or (layer0_outputs(1129));
    layer1_outputs(2897) <= not(layer0_outputs(5144));
    layer1_outputs(2898) <= not(layer0_outputs(3989)) or (layer0_outputs(1726));
    layer1_outputs(2899) <= not(layer0_outputs(4279));
    layer1_outputs(2900) <= not(layer0_outputs(1240)) or (layer0_outputs(3640));
    layer1_outputs(2901) <= not((layer0_outputs(3142)) or (layer0_outputs(3077)));
    layer1_outputs(2902) <= '0';
    layer1_outputs(2903) <= layer0_outputs(1405);
    layer1_outputs(2904) <= (layer0_outputs(5676)) and not (layer0_outputs(1492));
    layer1_outputs(2905) <= not(layer0_outputs(2899));
    layer1_outputs(2906) <= '1';
    layer1_outputs(2907) <= not(layer0_outputs(6025)) or (layer0_outputs(7115));
    layer1_outputs(2908) <= (layer0_outputs(503)) and (layer0_outputs(5638));
    layer1_outputs(2909) <= not(layer0_outputs(721)) or (layer0_outputs(4788));
    layer1_outputs(2910) <= '0';
    layer1_outputs(2911) <= layer0_outputs(2053);
    layer1_outputs(2912) <= not(layer0_outputs(1829)) or (layer0_outputs(6683));
    layer1_outputs(2913) <= (layer0_outputs(6608)) and not (layer0_outputs(86));
    layer1_outputs(2914) <= not((layer0_outputs(3159)) or (layer0_outputs(2620)));
    layer1_outputs(2915) <= (layer0_outputs(2721)) and (layer0_outputs(5857));
    layer1_outputs(2916) <= '1';
    layer1_outputs(2917) <= not(layer0_outputs(3195)) or (layer0_outputs(5540));
    layer1_outputs(2918) <= (layer0_outputs(4741)) and not (layer0_outputs(4171));
    layer1_outputs(2919) <= (layer0_outputs(4695)) or (layer0_outputs(7423));
    layer1_outputs(2920) <= not((layer0_outputs(5469)) and (layer0_outputs(6375)));
    layer1_outputs(2921) <= layer0_outputs(4409);
    layer1_outputs(2922) <= not(layer0_outputs(5943)) or (layer0_outputs(7564));
    layer1_outputs(2923) <= not(layer0_outputs(4149)) or (layer0_outputs(6641));
    layer1_outputs(2924) <= (layer0_outputs(4703)) and not (layer0_outputs(6516));
    layer1_outputs(2925) <= not((layer0_outputs(271)) and (layer0_outputs(203)));
    layer1_outputs(2926) <= not(layer0_outputs(3555)) or (layer0_outputs(1753));
    layer1_outputs(2927) <= (layer0_outputs(1160)) and (layer0_outputs(3027));
    layer1_outputs(2928) <= (layer0_outputs(925)) and not (layer0_outputs(3483));
    layer1_outputs(2929) <= (layer0_outputs(2154)) and not (layer0_outputs(6985));
    layer1_outputs(2930) <= not(layer0_outputs(1909)) or (layer0_outputs(6890));
    layer1_outputs(2931) <= not(layer0_outputs(376));
    layer1_outputs(2932) <= '1';
    layer1_outputs(2933) <= (layer0_outputs(362)) and not (layer0_outputs(2766));
    layer1_outputs(2934) <= not(layer0_outputs(2584)) or (layer0_outputs(4428));
    layer1_outputs(2935) <= not(layer0_outputs(5707)) or (layer0_outputs(5448));
    layer1_outputs(2936) <= (layer0_outputs(1166)) and (layer0_outputs(2020));
    layer1_outputs(2937) <= not(layer0_outputs(314));
    layer1_outputs(2938) <= not(layer0_outputs(793));
    layer1_outputs(2939) <= not((layer0_outputs(3720)) or (layer0_outputs(3699)));
    layer1_outputs(2940) <= layer0_outputs(5154);
    layer1_outputs(2941) <= layer0_outputs(2671);
    layer1_outputs(2942) <= (layer0_outputs(3370)) and not (layer0_outputs(5747));
    layer1_outputs(2943) <= not(layer0_outputs(7222));
    layer1_outputs(2944) <= (layer0_outputs(7054)) or (layer0_outputs(7621));
    layer1_outputs(2945) <= '1';
    layer1_outputs(2946) <= not(layer0_outputs(725)) or (layer0_outputs(4986));
    layer1_outputs(2947) <= not(layer0_outputs(3908));
    layer1_outputs(2948) <= (layer0_outputs(2050)) and not (layer0_outputs(3067));
    layer1_outputs(2949) <= not((layer0_outputs(7305)) or (layer0_outputs(4232)));
    layer1_outputs(2950) <= not((layer0_outputs(4933)) or (layer0_outputs(7133)));
    layer1_outputs(2951) <= not(layer0_outputs(510)) or (layer0_outputs(2887));
    layer1_outputs(2952) <= not(layer0_outputs(2783));
    layer1_outputs(2953) <= (layer0_outputs(171)) and (layer0_outputs(2094));
    layer1_outputs(2954) <= (layer0_outputs(1570)) and (layer0_outputs(4411));
    layer1_outputs(2955) <= not((layer0_outputs(2467)) or (layer0_outputs(6252)));
    layer1_outputs(2956) <= (layer0_outputs(2452)) and not (layer0_outputs(4325));
    layer1_outputs(2957) <= (layer0_outputs(870)) and (layer0_outputs(3748));
    layer1_outputs(2958) <= (layer0_outputs(201)) or (layer0_outputs(3561));
    layer1_outputs(2959) <= (layer0_outputs(488)) and (layer0_outputs(5397));
    layer1_outputs(2960) <= (layer0_outputs(2168)) and (layer0_outputs(4556));
    layer1_outputs(2961) <= not(layer0_outputs(1032));
    layer1_outputs(2962) <= layer0_outputs(7538);
    layer1_outputs(2963) <= layer0_outputs(6930);
    layer1_outputs(2964) <= (layer0_outputs(4963)) and (layer0_outputs(693));
    layer1_outputs(2965) <= not((layer0_outputs(529)) and (layer0_outputs(500)));
    layer1_outputs(2966) <= layer0_outputs(7544);
    layer1_outputs(2967) <= not(layer0_outputs(1568));
    layer1_outputs(2968) <= not(layer0_outputs(723)) or (layer0_outputs(1610));
    layer1_outputs(2969) <= not((layer0_outputs(5023)) or (layer0_outputs(4060)));
    layer1_outputs(2970) <= (layer0_outputs(4511)) and (layer0_outputs(1659));
    layer1_outputs(2971) <= layer0_outputs(5461);
    layer1_outputs(2972) <= '1';
    layer1_outputs(2973) <= '0';
    layer1_outputs(2974) <= layer0_outputs(45);
    layer1_outputs(2975) <= not(layer0_outputs(2231)) or (layer0_outputs(7048));
    layer1_outputs(2976) <= not((layer0_outputs(3406)) and (layer0_outputs(2634)));
    layer1_outputs(2977) <= (layer0_outputs(2486)) and (layer0_outputs(6589));
    layer1_outputs(2978) <= not(layer0_outputs(5506)) or (layer0_outputs(2130));
    layer1_outputs(2979) <= layer0_outputs(15);
    layer1_outputs(2980) <= not((layer0_outputs(298)) and (layer0_outputs(6328)));
    layer1_outputs(2981) <= not((layer0_outputs(5532)) and (layer0_outputs(1873)));
    layer1_outputs(2982) <= not(layer0_outputs(1123));
    layer1_outputs(2983) <= (layer0_outputs(4531)) and not (layer0_outputs(2843));
    layer1_outputs(2984) <= not((layer0_outputs(2277)) xor (layer0_outputs(1231)));
    layer1_outputs(2985) <= (layer0_outputs(5128)) and not (layer0_outputs(2424));
    layer1_outputs(2986) <= (layer0_outputs(4814)) or (layer0_outputs(7051));
    layer1_outputs(2987) <= not((layer0_outputs(3471)) and (layer0_outputs(2801)));
    layer1_outputs(2988) <= layer0_outputs(4056);
    layer1_outputs(2989) <= '1';
    layer1_outputs(2990) <= not(layer0_outputs(4794)) or (layer0_outputs(127));
    layer1_outputs(2991) <= not((layer0_outputs(6991)) or (layer0_outputs(1480)));
    layer1_outputs(2992) <= (layer0_outputs(35)) and not (layer0_outputs(6623));
    layer1_outputs(2993) <= (layer0_outputs(3592)) or (layer0_outputs(1003));
    layer1_outputs(2994) <= not(layer0_outputs(6072));
    layer1_outputs(2995) <= not(layer0_outputs(4521));
    layer1_outputs(2996) <= '1';
    layer1_outputs(2997) <= not((layer0_outputs(4641)) or (layer0_outputs(5091)));
    layer1_outputs(2998) <= not(layer0_outputs(5054));
    layer1_outputs(2999) <= (layer0_outputs(4407)) and not (layer0_outputs(2879));
    layer1_outputs(3000) <= (layer0_outputs(6899)) and not (layer0_outputs(3309));
    layer1_outputs(3001) <= not(layer0_outputs(533));
    layer1_outputs(3002) <= not((layer0_outputs(1698)) and (layer0_outputs(6313)));
    layer1_outputs(3003) <= layer0_outputs(7338);
    layer1_outputs(3004) <= not(layer0_outputs(400)) or (layer0_outputs(3070));
    layer1_outputs(3005) <= not(layer0_outputs(4099));
    layer1_outputs(3006) <= not((layer0_outputs(3629)) or (layer0_outputs(6782)));
    layer1_outputs(3007) <= layer0_outputs(5931);
    layer1_outputs(3008) <= layer0_outputs(2966);
    layer1_outputs(3009) <= layer0_outputs(3228);
    layer1_outputs(3010) <= not(layer0_outputs(1606));
    layer1_outputs(3011) <= not(layer0_outputs(4790)) or (layer0_outputs(1460));
    layer1_outputs(3012) <= (layer0_outputs(1725)) and (layer0_outputs(3613));
    layer1_outputs(3013) <= '0';
    layer1_outputs(3014) <= (layer0_outputs(4110)) or (layer0_outputs(360));
    layer1_outputs(3015) <= not(layer0_outputs(3052));
    layer1_outputs(3016) <= layer0_outputs(1538);
    layer1_outputs(3017) <= (layer0_outputs(5837)) and not (layer0_outputs(2638));
    layer1_outputs(3018) <= not(layer0_outputs(7094));
    layer1_outputs(3019) <= not((layer0_outputs(5307)) or (layer0_outputs(998)));
    layer1_outputs(3020) <= not(layer0_outputs(749)) or (layer0_outputs(2964));
    layer1_outputs(3021) <= (layer0_outputs(1904)) and not (layer0_outputs(1634));
    layer1_outputs(3022) <= not(layer0_outputs(1366));
    layer1_outputs(3023) <= layer0_outputs(690);
    layer1_outputs(3024) <= '1';
    layer1_outputs(3025) <= not(layer0_outputs(4036));
    layer1_outputs(3026) <= layer0_outputs(7335);
    layer1_outputs(3027) <= not(layer0_outputs(6216)) or (layer0_outputs(5344));
    layer1_outputs(3028) <= (layer0_outputs(3366)) and not (layer0_outputs(7376));
    layer1_outputs(3029) <= '1';
    layer1_outputs(3030) <= (layer0_outputs(3455)) and not (layer0_outputs(2140));
    layer1_outputs(3031) <= not(layer0_outputs(716));
    layer1_outputs(3032) <= not(layer0_outputs(3035)) or (layer0_outputs(4671));
    layer1_outputs(3033) <= not(layer0_outputs(6443));
    layer1_outputs(3034) <= not(layer0_outputs(3590)) or (layer0_outputs(368));
    layer1_outputs(3035) <= layer0_outputs(4989);
    layer1_outputs(3036) <= (layer0_outputs(2226)) or (layer0_outputs(4485));
    layer1_outputs(3037) <= not(layer0_outputs(43)) or (layer0_outputs(3073));
    layer1_outputs(3038) <= (layer0_outputs(2828)) and not (layer0_outputs(4566));
    layer1_outputs(3039) <= (layer0_outputs(5122)) and not (layer0_outputs(2792));
    layer1_outputs(3040) <= not((layer0_outputs(543)) or (layer0_outputs(3748)));
    layer1_outputs(3041) <= '1';
    layer1_outputs(3042) <= not(layer0_outputs(1226)) or (layer0_outputs(6488));
    layer1_outputs(3043) <= (layer0_outputs(686)) and not (layer0_outputs(3845));
    layer1_outputs(3044) <= (layer0_outputs(1677)) and not (layer0_outputs(5840));
    layer1_outputs(3045) <= not((layer0_outputs(2117)) or (layer0_outputs(5213)));
    layer1_outputs(3046) <= not(layer0_outputs(5356));
    layer1_outputs(3047) <= not((layer0_outputs(1413)) and (layer0_outputs(4942)));
    layer1_outputs(3048) <= (layer0_outputs(6819)) and not (layer0_outputs(3446));
    layer1_outputs(3049) <= not(layer0_outputs(4097)) or (layer0_outputs(4808));
    layer1_outputs(3050) <= layer0_outputs(1035);
    layer1_outputs(3051) <= not(layer0_outputs(2576));
    layer1_outputs(3052) <= not(layer0_outputs(989)) or (layer0_outputs(361));
    layer1_outputs(3053) <= not(layer0_outputs(6474));
    layer1_outputs(3054) <= (layer0_outputs(1107)) and not (layer0_outputs(3296));
    layer1_outputs(3055) <= not(layer0_outputs(4770));
    layer1_outputs(3056) <= (layer0_outputs(3303)) and not (layer0_outputs(6898));
    layer1_outputs(3057) <= not(layer0_outputs(4375));
    layer1_outputs(3058) <= not(layer0_outputs(5409)) or (layer0_outputs(570));
    layer1_outputs(3059) <= '1';
    layer1_outputs(3060) <= not((layer0_outputs(3479)) or (layer0_outputs(1730)));
    layer1_outputs(3061) <= layer0_outputs(3040);
    layer1_outputs(3062) <= not((layer0_outputs(5941)) or (layer0_outputs(778)));
    layer1_outputs(3063) <= layer0_outputs(3517);
    layer1_outputs(3064) <= (layer0_outputs(3185)) and not (layer0_outputs(1747));
    layer1_outputs(3065) <= layer0_outputs(6493);
    layer1_outputs(3066) <= not(layer0_outputs(1030));
    layer1_outputs(3067) <= layer0_outputs(4724);
    layer1_outputs(3068) <= layer0_outputs(7603);
    layer1_outputs(3069) <= not(layer0_outputs(142));
    layer1_outputs(3070) <= layer0_outputs(5557);
    layer1_outputs(3071) <= (layer0_outputs(7376)) and not (layer0_outputs(2835));
    layer1_outputs(3072) <= (layer0_outputs(2563)) and not (layer0_outputs(6785));
    layer1_outputs(3073) <= layer0_outputs(7144);
    layer1_outputs(3074) <= (layer0_outputs(7088)) and not (layer0_outputs(2301));
    layer1_outputs(3075) <= (layer0_outputs(5607)) xor (layer0_outputs(144));
    layer1_outputs(3076) <= not(layer0_outputs(44)) or (layer0_outputs(613));
    layer1_outputs(3077) <= (layer0_outputs(7108)) and (layer0_outputs(80));
    layer1_outputs(3078) <= not(layer0_outputs(2861));
    layer1_outputs(3079) <= not(layer0_outputs(4203)) or (layer0_outputs(1338));
    layer1_outputs(3080) <= not(layer0_outputs(5));
    layer1_outputs(3081) <= layer0_outputs(5599);
    layer1_outputs(3082) <= (layer0_outputs(4028)) or (layer0_outputs(1890));
    layer1_outputs(3083) <= not(layer0_outputs(3790)) or (layer0_outputs(2092));
    layer1_outputs(3084) <= not((layer0_outputs(2125)) or (layer0_outputs(6810)));
    layer1_outputs(3085) <= (layer0_outputs(474)) and not (layer0_outputs(7568));
    layer1_outputs(3086) <= not((layer0_outputs(5811)) xor (layer0_outputs(1551)));
    layer1_outputs(3087) <= (layer0_outputs(6642)) and not (layer0_outputs(2404));
    layer1_outputs(3088) <= not(layer0_outputs(4372));
    layer1_outputs(3089) <= '0';
    layer1_outputs(3090) <= layer0_outputs(2826);
    layer1_outputs(3091) <= layer0_outputs(3911);
    layer1_outputs(3092) <= not((layer0_outputs(1532)) and (layer0_outputs(1475)));
    layer1_outputs(3093) <= '0';
    layer1_outputs(3094) <= not(layer0_outputs(6740));
    layer1_outputs(3095) <= not(layer0_outputs(6839)) or (layer0_outputs(891));
    layer1_outputs(3096) <= not(layer0_outputs(2895));
    layer1_outputs(3097) <= not(layer0_outputs(3353));
    layer1_outputs(3098) <= layer0_outputs(4918);
    layer1_outputs(3099) <= (layer0_outputs(5186)) or (layer0_outputs(3804));
    layer1_outputs(3100) <= not(layer0_outputs(4154));
    layer1_outputs(3101) <= not(layer0_outputs(4065));
    layer1_outputs(3102) <= not(layer0_outputs(6054)) or (layer0_outputs(2828));
    layer1_outputs(3103) <= (layer0_outputs(5813)) and not (layer0_outputs(5885));
    layer1_outputs(3104) <= not(layer0_outputs(5055)) or (layer0_outputs(5767));
    layer1_outputs(3105) <= '1';
    layer1_outputs(3106) <= '1';
    layer1_outputs(3107) <= (layer0_outputs(1419)) and not (layer0_outputs(4128));
    layer1_outputs(3108) <= layer0_outputs(528);
    layer1_outputs(3109) <= not(layer0_outputs(6175)) or (layer0_outputs(6922));
    layer1_outputs(3110) <= (layer0_outputs(5784)) xor (layer0_outputs(4921));
    layer1_outputs(3111) <= not((layer0_outputs(1249)) or (layer0_outputs(7582)));
    layer1_outputs(3112) <= (layer0_outputs(3481)) and (layer0_outputs(6116));
    layer1_outputs(3113) <= layer0_outputs(3783);
    layer1_outputs(3114) <= not(layer0_outputs(7093)) or (layer0_outputs(6380));
    layer1_outputs(3115) <= '0';
    layer1_outputs(3116) <= '1';
    layer1_outputs(3117) <= (layer0_outputs(2239)) or (layer0_outputs(1096));
    layer1_outputs(3118) <= '1';
    layer1_outputs(3119) <= layer0_outputs(2769);
    layer1_outputs(3120) <= not((layer0_outputs(6289)) and (layer0_outputs(7326)));
    layer1_outputs(3121) <= not(layer0_outputs(1172));
    layer1_outputs(3122) <= layer0_outputs(2878);
    layer1_outputs(3123) <= not(layer0_outputs(2714));
    layer1_outputs(3124) <= not(layer0_outputs(59));
    layer1_outputs(3125) <= (layer0_outputs(6136)) xor (layer0_outputs(1479));
    layer1_outputs(3126) <= (layer0_outputs(6067)) and not (layer0_outputs(5681));
    layer1_outputs(3127) <= not((layer0_outputs(6805)) xor (layer0_outputs(4139)));
    layer1_outputs(3128) <= not(layer0_outputs(1179));
    layer1_outputs(3129) <= (layer0_outputs(5999)) xor (layer0_outputs(821));
    layer1_outputs(3130) <= '0';
    layer1_outputs(3131) <= (layer0_outputs(2076)) and (layer0_outputs(6434));
    layer1_outputs(3132) <= not(layer0_outputs(82)) or (layer0_outputs(403));
    layer1_outputs(3133) <= not((layer0_outputs(4893)) or (layer0_outputs(3025)));
    layer1_outputs(3134) <= layer0_outputs(5322);
    layer1_outputs(3135) <= not(layer0_outputs(915)) or (layer0_outputs(3431));
    layer1_outputs(3136) <= not(layer0_outputs(6436)) or (layer0_outputs(4084));
    layer1_outputs(3137) <= layer0_outputs(2602);
    layer1_outputs(3138) <= not(layer0_outputs(5360));
    layer1_outputs(3139) <= layer0_outputs(139);
    layer1_outputs(3140) <= not(layer0_outputs(4895));
    layer1_outputs(3141) <= (layer0_outputs(5893)) or (layer0_outputs(338));
    layer1_outputs(3142) <= (layer0_outputs(5076)) and (layer0_outputs(214));
    layer1_outputs(3143) <= (layer0_outputs(7426)) and not (layer0_outputs(4272));
    layer1_outputs(3144) <= (layer0_outputs(4917)) and (layer0_outputs(4549));
    layer1_outputs(3145) <= not(layer0_outputs(5838)) or (layer0_outputs(1103));
    layer1_outputs(3146) <= '1';
    layer1_outputs(3147) <= (layer0_outputs(2021)) xor (layer0_outputs(1388));
    layer1_outputs(3148) <= (layer0_outputs(7008)) and not (layer0_outputs(5491));
    layer1_outputs(3149) <= not(layer0_outputs(4403)) or (layer0_outputs(224));
    layer1_outputs(3150) <= '1';
    layer1_outputs(3151) <= '0';
    layer1_outputs(3152) <= (layer0_outputs(7099)) and not (layer0_outputs(1972));
    layer1_outputs(3153) <= (layer0_outputs(4726)) or (layer0_outputs(2894));
    layer1_outputs(3154) <= not(layer0_outputs(4940)) or (layer0_outputs(5438));
    layer1_outputs(3155) <= (layer0_outputs(425)) and not (layer0_outputs(4967));
    layer1_outputs(3156) <= (layer0_outputs(4990)) and (layer0_outputs(6148));
    layer1_outputs(3157) <= (layer0_outputs(3994)) and not (layer0_outputs(6526));
    layer1_outputs(3158) <= layer0_outputs(1637);
    layer1_outputs(3159) <= not(layer0_outputs(5741));
    layer1_outputs(3160) <= not((layer0_outputs(4930)) and (layer0_outputs(7317)));
    layer1_outputs(3161) <= not(layer0_outputs(420)) or (layer0_outputs(1638));
    layer1_outputs(3162) <= not(layer0_outputs(5602));
    layer1_outputs(3163) <= not((layer0_outputs(4689)) or (layer0_outputs(3055)));
    layer1_outputs(3164) <= (layer0_outputs(5336)) or (layer0_outputs(3334));
    layer1_outputs(3165) <= not(layer0_outputs(173));
    layer1_outputs(3166) <= not(layer0_outputs(3562));
    layer1_outputs(3167) <= layer0_outputs(4460);
    layer1_outputs(3168) <= (layer0_outputs(6764)) or (layer0_outputs(7591));
    layer1_outputs(3169) <= not(layer0_outputs(6123));
    layer1_outputs(3170) <= not(layer0_outputs(3262));
    layer1_outputs(3171) <= (layer0_outputs(153)) and not (layer0_outputs(4892));
    layer1_outputs(3172) <= layer0_outputs(2434);
    layer1_outputs(3173) <= not((layer0_outputs(2002)) or (layer0_outputs(3127)));
    layer1_outputs(3174) <= (layer0_outputs(7622)) and not (layer0_outputs(1138));
    layer1_outputs(3175) <= not(layer0_outputs(5345));
    layer1_outputs(3176) <= not(layer0_outputs(3833));
    layer1_outputs(3177) <= (layer0_outputs(963)) or (layer0_outputs(1682));
    layer1_outputs(3178) <= (layer0_outputs(484)) xor (layer0_outputs(4287));
    layer1_outputs(3179) <= (layer0_outputs(4520)) xor (layer0_outputs(300));
    layer1_outputs(3180) <= '1';
    layer1_outputs(3181) <= not(layer0_outputs(3955));
    layer1_outputs(3182) <= (layer0_outputs(556)) and not (layer0_outputs(7418));
    layer1_outputs(3183) <= '0';
    layer1_outputs(3184) <= layer0_outputs(4136);
    layer1_outputs(3185) <= (layer0_outputs(3723)) and not (layer0_outputs(3119));
    layer1_outputs(3186) <= not(layer0_outputs(2545)) or (layer0_outputs(1459));
    layer1_outputs(3187) <= layer0_outputs(1266);
    layer1_outputs(3188) <= (layer0_outputs(6113)) and not (layer0_outputs(2298));
    layer1_outputs(3189) <= layer0_outputs(1419);
    layer1_outputs(3190) <= (layer0_outputs(2155)) or (layer0_outputs(4117));
    layer1_outputs(3191) <= (layer0_outputs(6956)) or (layer0_outputs(6967));
    layer1_outputs(3192) <= '0';
    layer1_outputs(3193) <= (layer0_outputs(2938)) and not (layer0_outputs(2595));
    layer1_outputs(3194) <= (layer0_outputs(4807)) or (layer0_outputs(29));
    layer1_outputs(3195) <= not(layer0_outputs(1935));
    layer1_outputs(3196) <= (layer0_outputs(3229)) and (layer0_outputs(4214));
    layer1_outputs(3197) <= layer0_outputs(3679);
    layer1_outputs(3198) <= not(layer0_outputs(4654));
    layer1_outputs(3199) <= layer0_outputs(2747);
    layer1_outputs(3200) <= (layer0_outputs(973)) and not (layer0_outputs(959));
    layer1_outputs(3201) <= not((layer0_outputs(6843)) and (layer0_outputs(3063)));
    layer1_outputs(3202) <= (layer0_outputs(5977)) xor (layer0_outputs(7332));
    layer1_outputs(3203) <= not(layer0_outputs(1831));
    layer1_outputs(3204) <= '1';
    layer1_outputs(3205) <= '0';
    layer1_outputs(3206) <= not((layer0_outputs(3729)) and (layer0_outputs(3822)));
    layer1_outputs(3207) <= not(layer0_outputs(560)) or (layer0_outputs(7080));
    layer1_outputs(3208) <= layer0_outputs(2909);
    layer1_outputs(3209) <= layer0_outputs(4909);
    layer1_outputs(3210) <= (layer0_outputs(3926)) or (layer0_outputs(4499));
    layer1_outputs(3211) <= not(layer0_outputs(3408));
    layer1_outputs(3212) <= not(layer0_outputs(995));
    layer1_outputs(3213) <= layer0_outputs(2771);
    layer1_outputs(3214) <= not((layer0_outputs(6326)) and (layer0_outputs(5470)));
    layer1_outputs(3215) <= (layer0_outputs(6221)) and (layer0_outputs(5782));
    layer1_outputs(3216) <= (layer0_outputs(2613)) and not (layer0_outputs(745));
    layer1_outputs(3217) <= '1';
    layer1_outputs(3218) <= (layer0_outputs(3820)) or (layer0_outputs(2413));
    layer1_outputs(3219) <= not(layer0_outputs(1676));
    layer1_outputs(3220) <= not((layer0_outputs(1563)) and (layer0_outputs(3524)));
    layer1_outputs(3221) <= '1';
    layer1_outputs(3222) <= (layer0_outputs(1062)) and (layer0_outputs(4811));
    layer1_outputs(3223) <= not(layer0_outputs(6536)) or (layer0_outputs(5216));
    layer1_outputs(3224) <= not((layer0_outputs(2363)) and (layer0_outputs(6809)));
    layer1_outputs(3225) <= not((layer0_outputs(1010)) and (layer0_outputs(6459)));
    layer1_outputs(3226) <= not(layer0_outputs(5906)) or (layer0_outputs(4971));
    layer1_outputs(3227) <= not(layer0_outputs(5305));
    layer1_outputs(3228) <= not(layer0_outputs(2366)) or (layer0_outputs(1057));
    layer1_outputs(3229) <= layer0_outputs(5079);
    layer1_outputs(3230) <= not(layer0_outputs(2618));
    layer1_outputs(3231) <= not(layer0_outputs(2511));
    layer1_outputs(3232) <= not(layer0_outputs(5643)) or (layer0_outputs(794));
    layer1_outputs(3233) <= layer0_outputs(1104);
    layer1_outputs(3234) <= not((layer0_outputs(4353)) xor (layer0_outputs(6682)));
    layer1_outputs(3235) <= (layer0_outputs(6664)) and not (layer0_outputs(3112));
    layer1_outputs(3236) <= not(layer0_outputs(6044));
    layer1_outputs(3237) <= (layer0_outputs(3558)) xor (layer0_outputs(5600));
    layer1_outputs(3238) <= not(layer0_outputs(4648)) or (layer0_outputs(4356));
    layer1_outputs(3239) <= '0';
    layer1_outputs(3240) <= not(layer0_outputs(2025)) or (layer0_outputs(5297));
    layer1_outputs(3241) <= not(layer0_outputs(7665)) or (layer0_outputs(464));
    layer1_outputs(3242) <= (layer0_outputs(1553)) and (layer0_outputs(46));
    layer1_outputs(3243) <= not(layer0_outputs(5967)) or (layer0_outputs(402));
    layer1_outputs(3244) <= not(layer0_outputs(6540));
    layer1_outputs(3245) <= not(layer0_outputs(7217)) or (layer0_outputs(6340));
    layer1_outputs(3246) <= (layer0_outputs(2701)) and not (layer0_outputs(3301));
    layer1_outputs(3247) <= layer0_outputs(473);
    layer1_outputs(3248) <= not(layer0_outputs(1351)) or (layer0_outputs(5580));
    layer1_outputs(3249) <= (layer0_outputs(3605)) or (layer0_outputs(2275));
    layer1_outputs(3250) <= not((layer0_outputs(1939)) xor (layer0_outputs(4073)));
    layer1_outputs(3251) <= '0';
    layer1_outputs(3252) <= not(layer0_outputs(4919)) or (layer0_outputs(3226));
    layer1_outputs(3253) <= not(layer0_outputs(4391));
    layer1_outputs(3254) <= not(layer0_outputs(2738));
    layer1_outputs(3255) <= (layer0_outputs(6039)) and not (layer0_outputs(2515));
    layer1_outputs(3256) <= not(layer0_outputs(6013)) or (layer0_outputs(7179));
    layer1_outputs(3257) <= (layer0_outputs(2647)) and not (layer0_outputs(7258));
    layer1_outputs(3258) <= not(layer0_outputs(1377));
    layer1_outputs(3259) <= layer0_outputs(1161);
    layer1_outputs(3260) <= not(layer0_outputs(5050)) or (layer0_outputs(6714));
    layer1_outputs(3261) <= (layer0_outputs(5308)) and (layer0_outputs(3928));
    layer1_outputs(3262) <= (layer0_outputs(187)) or (layer0_outputs(3969));
    layer1_outputs(3263) <= (layer0_outputs(1647)) and not (layer0_outputs(1737));
    layer1_outputs(3264) <= layer0_outputs(676);
    layer1_outputs(3265) <= not(layer0_outputs(5367));
    layer1_outputs(3266) <= (layer0_outputs(2901)) and not (layer0_outputs(6067));
    layer1_outputs(3267) <= not(layer0_outputs(6219));
    layer1_outputs(3268) <= layer0_outputs(4018);
    layer1_outputs(3269) <= not(layer0_outputs(64)) or (layer0_outputs(2412));
    layer1_outputs(3270) <= (layer0_outputs(4364)) or (layer0_outputs(5200));
    layer1_outputs(3271) <= '0';
    layer1_outputs(3272) <= layer0_outputs(2075);
    layer1_outputs(3273) <= layer0_outputs(3667);
    layer1_outputs(3274) <= not((layer0_outputs(4253)) and (layer0_outputs(6650)));
    layer1_outputs(3275) <= not((layer0_outputs(7410)) and (layer0_outputs(1184)));
    layer1_outputs(3276) <= not(layer0_outputs(4336));
    layer1_outputs(3277) <= '1';
    layer1_outputs(3278) <= (layer0_outputs(2180)) or (layer0_outputs(533));
    layer1_outputs(3279) <= '0';
    layer1_outputs(3280) <= not(layer0_outputs(6143)) or (layer0_outputs(5021));
    layer1_outputs(3281) <= layer0_outputs(1312);
    layer1_outputs(3282) <= (layer0_outputs(2079)) and not (layer0_outputs(5964));
    layer1_outputs(3283) <= (layer0_outputs(3333)) and (layer0_outputs(1237));
    layer1_outputs(3284) <= not(layer0_outputs(5124));
    layer1_outputs(3285) <= layer0_outputs(7078);
    layer1_outputs(3286) <= (layer0_outputs(1307)) and (layer0_outputs(5617));
    layer1_outputs(3287) <= not((layer0_outputs(2639)) or (layer0_outputs(4662)));
    layer1_outputs(3288) <= (layer0_outputs(4745)) and not (layer0_outputs(333));
    layer1_outputs(3289) <= not((layer0_outputs(5987)) xor (layer0_outputs(3370)));
    layer1_outputs(3290) <= (layer0_outputs(5083)) and not (layer0_outputs(5218));
    layer1_outputs(3291) <= '1';
    layer1_outputs(3292) <= (layer0_outputs(3065)) and (layer0_outputs(4413));
    layer1_outputs(3293) <= layer0_outputs(5591);
    layer1_outputs(3294) <= (layer0_outputs(1466)) xor (layer0_outputs(4510));
    layer1_outputs(3295) <= (layer0_outputs(4584)) and not (layer0_outputs(7188));
    layer1_outputs(3296) <= not((layer0_outputs(1359)) or (layer0_outputs(1948)));
    layer1_outputs(3297) <= not(layer0_outputs(2349));
    layer1_outputs(3298) <= not((layer0_outputs(6633)) or (layer0_outputs(6059)));
    layer1_outputs(3299) <= layer0_outputs(225);
    layer1_outputs(3300) <= not(layer0_outputs(2641));
    layer1_outputs(3301) <= not((layer0_outputs(3066)) or (layer0_outputs(5473)));
    layer1_outputs(3302) <= not((layer0_outputs(1025)) or (layer0_outputs(3959)));
    layer1_outputs(3303) <= layer0_outputs(2531);
    layer1_outputs(3304) <= (layer0_outputs(5014)) xor (layer0_outputs(5024));
    layer1_outputs(3305) <= not((layer0_outputs(6999)) or (layer0_outputs(2487)));
    layer1_outputs(3306) <= (layer0_outputs(5964)) and not (layer0_outputs(2448));
    layer1_outputs(3307) <= not(layer0_outputs(7229));
    layer1_outputs(3308) <= not((layer0_outputs(4223)) or (layer0_outputs(6202)));
    layer1_outputs(3309) <= layer0_outputs(7301);
    layer1_outputs(3310) <= not((layer0_outputs(7580)) and (layer0_outputs(1456)));
    layer1_outputs(3311) <= (layer0_outputs(675)) and (layer0_outputs(227));
    layer1_outputs(3312) <= layer0_outputs(4132);
    layer1_outputs(3313) <= not((layer0_outputs(4841)) or (layer0_outputs(4196)));
    layer1_outputs(3314) <= not((layer0_outputs(2811)) and (layer0_outputs(3260)));
    layer1_outputs(3315) <= (layer0_outputs(1347)) and (layer0_outputs(1438));
    layer1_outputs(3316) <= layer0_outputs(6112);
    layer1_outputs(3317) <= not(layer0_outputs(1069));
    layer1_outputs(3318) <= not((layer0_outputs(5971)) and (layer0_outputs(2830)));
    layer1_outputs(3319) <= not(layer0_outputs(1696)) or (layer0_outputs(4481));
    layer1_outputs(3320) <= not((layer0_outputs(38)) and (layer0_outputs(4712)));
    layer1_outputs(3321) <= layer0_outputs(3178);
    layer1_outputs(3322) <= not(layer0_outputs(4936));
    layer1_outputs(3323) <= not(layer0_outputs(2128)) or (layer0_outputs(7620));
    layer1_outputs(3324) <= not(layer0_outputs(4516)) or (layer0_outputs(7065));
    layer1_outputs(3325) <= not(layer0_outputs(3208)) or (layer0_outputs(1683));
    layer1_outputs(3326) <= not((layer0_outputs(2173)) or (layer0_outputs(6004)));
    layer1_outputs(3327) <= not((layer0_outputs(872)) and (layer0_outputs(1897)));
    layer1_outputs(3328) <= layer0_outputs(1319);
    layer1_outputs(3329) <= not(layer0_outputs(4068));
    layer1_outputs(3330) <= (layer0_outputs(6481)) and not (layer0_outputs(7494));
    layer1_outputs(3331) <= not(layer0_outputs(2161)) or (layer0_outputs(1061));
    layer1_outputs(3332) <= not(layer0_outputs(890)) or (layer0_outputs(2484));
    layer1_outputs(3333) <= not((layer0_outputs(3012)) or (layer0_outputs(577)));
    layer1_outputs(3334) <= not((layer0_outputs(1126)) and (layer0_outputs(6313)));
    layer1_outputs(3335) <= not(layer0_outputs(7314)) or (layer0_outputs(6704));
    layer1_outputs(3336) <= layer0_outputs(4970);
    layer1_outputs(3337) <= not(layer0_outputs(4899)) or (layer0_outputs(5073));
    layer1_outputs(3338) <= (layer0_outputs(4234)) xor (layer0_outputs(3426));
    layer1_outputs(3339) <= not((layer0_outputs(6403)) or (layer0_outputs(4903)));
    layer1_outputs(3340) <= layer0_outputs(5629);
    layer1_outputs(3341) <= (layer0_outputs(1182)) and not (layer0_outputs(4719));
    layer1_outputs(3342) <= (layer0_outputs(5017)) and not (layer0_outputs(3144));
    layer1_outputs(3343) <= not(layer0_outputs(5577));
    layer1_outputs(3344) <= not(layer0_outputs(7049)) or (layer0_outputs(999));
    layer1_outputs(3345) <= layer0_outputs(5383);
    layer1_outputs(3346) <= (layer0_outputs(6778)) and (layer0_outputs(2799));
    layer1_outputs(3347) <= not(layer0_outputs(1839));
    layer1_outputs(3348) <= not(layer0_outputs(6038));
    layer1_outputs(3349) <= not((layer0_outputs(3878)) or (layer0_outputs(799)));
    layer1_outputs(3350) <= (layer0_outputs(5135)) or (layer0_outputs(7654));
    layer1_outputs(3351) <= '0';
    layer1_outputs(3352) <= (layer0_outputs(7001)) and not (layer0_outputs(2732));
    layer1_outputs(3353) <= (layer0_outputs(2108)) and not (layer0_outputs(2450));
    layer1_outputs(3354) <= not(layer0_outputs(3568));
    layer1_outputs(3355) <= not(layer0_outputs(6273));
    layer1_outputs(3356) <= not(layer0_outputs(3618));
    layer1_outputs(3357) <= not(layer0_outputs(3033)) or (layer0_outputs(7459));
    layer1_outputs(3358) <= (layer0_outputs(4057)) and not (layer0_outputs(568));
    layer1_outputs(3359) <= not(layer0_outputs(969)) or (layer0_outputs(3983));
    layer1_outputs(3360) <= (layer0_outputs(6009)) and not (layer0_outputs(814));
    layer1_outputs(3361) <= layer0_outputs(479);
    layer1_outputs(3362) <= not((layer0_outputs(306)) and (layer0_outputs(3021)));
    layer1_outputs(3363) <= '0';
    layer1_outputs(3364) <= (layer0_outputs(5561)) and not (layer0_outputs(4738));
    layer1_outputs(3365) <= not((layer0_outputs(2965)) or (layer0_outputs(4035)));
    layer1_outputs(3366) <= not(layer0_outputs(6630));
    layer1_outputs(3367) <= not((layer0_outputs(5150)) and (layer0_outputs(4298)));
    layer1_outputs(3368) <= layer0_outputs(5703);
    layer1_outputs(3369) <= not(layer0_outputs(2695)) or (layer0_outputs(607));
    layer1_outputs(3370) <= not((layer0_outputs(87)) or (layer0_outputs(5590)));
    layer1_outputs(3371) <= not(layer0_outputs(2495));
    layer1_outputs(3372) <= not(layer0_outputs(7647));
    layer1_outputs(3373) <= not(layer0_outputs(2788)) or (layer0_outputs(4074));
    layer1_outputs(3374) <= not(layer0_outputs(7065)) or (layer0_outputs(175));
    layer1_outputs(3375) <= layer0_outputs(2054);
    layer1_outputs(3376) <= not((layer0_outputs(2387)) and (layer0_outputs(3478)));
    layer1_outputs(3377) <= not((layer0_outputs(5545)) or (layer0_outputs(1811)));
    layer1_outputs(3378) <= not(layer0_outputs(4538));
    layer1_outputs(3379) <= layer0_outputs(2407);
    layer1_outputs(3380) <= not(layer0_outputs(1131)) or (layer0_outputs(5052));
    layer1_outputs(3381) <= not((layer0_outputs(4548)) or (layer0_outputs(5700)));
    layer1_outputs(3382) <= (layer0_outputs(6826)) or (layer0_outputs(6040));
    layer1_outputs(3383) <= not(layer0_outputs(3131));
    layer1_outputs(3384) <= (layer0_outputs(6187)) and not (layer0_outputs(3573));
    layer1_outputs(3385) <= (layer0_outputs(5585)) or (layer0_outputs(3704));
    layer1_outputs(3386) <= not(layer0_outputs(1245));
    layer1_outputs(3387) <= (layer0_outputs(1259)) and (layer0_outputs(5295));
    layer1_outputs(3388) <= not(layer0_outputs(7304));
    layer1_outputs(3389) <= not(layer0_outputs(3500)) or (layer0_outputs(125));
    layer1_outputs(3390) <= layer0_outputs(976);
    layer1_outputs(3391) <= not((layer0_outputs(2362)) and (layer0_outputs(5778)));
    layer1_outputs(3392) <= not(layer0_outputs(4946)) or (layer0_outputs(2521));
    layer1_outputs(3393) <= '0';
    layer1_outputs(3394) <= layer0_outputs(6);
    layer1_outputs(3395) <= not((layer0_outputs(2536)) or (layer0_outputs(2061)));
    layer1_outputs(3396) <= (layer0_outputs(1864)) and not (layer0_outputs(5118));
    layer1_outputs(3397) <= not((layer0_outputs(5990)) or (layer0_outputs(7669)));
    layer1_outputs(3398) <= not(layer0_outputs(1348));
    layer1_outputs(3399) <= (layer0_outputs(4378)) and not (layer0_outputs(632));
    layer1_outputs(3400) <= (layer0_outputs(1571)) or (layer0_outputs(7636));
    layer1_outputs(3401) <= not((layer0_outputs(2361)) xor (layer0_outputs(1339)));
    layer1_outputs(3402) <= (layer0_outputs(7336)) and (layer0_outputs(2675));
    layer1_outputs(3403) <= not((layer0_outputs(7232)) xor (layer0_outputs(4746)));
    layer1_outputs(3404) <= not(layer0_outputs(2232));
    layer1_outputs(3405) <= layer0_outputs(1908);
    layer1_outputs(3406) <= '1';
    layer1_outputs(3407) <= not(layer0_outputs(1007)) or (layer0_outputs(1642));
    layer1_outputs(3408) <= (layer0_outputs(4111)) xor (layer0_outputs(4688));
    layer1_outputs(3409) <= not(layer0_outputs(5381));
    layer1_outputs(3410) <= not((layer0_outputs(1392)) and (layer0_outputs(4269)));
    layer1_outputs(3411) <= not(layer0_outputs(3219));
    layer1_outputs(3412) <= not(layer0_outputs(6039));
    layer1_outputs(3413) <= (layer0_outputs(5683)) and not (layer0_outputs(6706));
    layer1_outputs(3414) <= not((layer0_outputs(7123)) and (layer0_outputs(6132)));
    layer1_outputs(3415) <= layer0_outputs(2162);
    layer1_outputs(3416) <= not((layer0_outputs(4062)) and (layer0_outputs(79)));
    layer1_outputs(3417) <= (layer0_outputs(6318)) or (layer0_outputs(4741));
    layer1_outputs(3418) <= not(layer0_outputs(4897));
    layer1_outputs(3419) <= (layer0_outputs(4333)) or (layer0_outputs(1924));
    layer1_outputs(3420) <= not(layer0_outputs(1135));
    layer1_outputs(3421) <= layer0_outputs(5395);
    layer1_outputs(3422) <= not((layer0_outputs(2435)) or (layer0_outputs(2933)));
    layer1_outputs(3423) <= not((layer0_outputs(1004)) or (layer0_outputs(6000)));
    layer1_outputs(3424) <= layer0_outputs(4171);
    layer1_outputs(3425) <= layer0_outputs(417);
    layer1_outputs(3426) <= (layer0_outputs(1090)) and not (layer0_outputs(5348));
    layer1_outputs(3427) <= layer0_outputs(1870);
    layer1_outputs(3428) <= not(layer0_outputs(5889)) or (layer0_outputs(6388));
    layer1_outputs(3429) <= not((layer0_outputs(324)) xor (layer0_outputs(6876)));
    layer1_outputs(3430) <= layer0_outputs(6922);
    layer1_outputs(3431) <= (layer0_outputs(3237)) and not (layer0_outputs(5979));
    layer1_outputs(3432) <= (layer0_outputs(7549)) xor (layer0_outputs(977));
    layer1_outputs(3433) <= '0';
    layer1_outputs(3434) <= (layer0_outputs(3204)) and (layer0_outputs(3676));
    layer1_outputs(3435) <= layer0_outputs(7590);
    layer1_outputs(3436) <= layer0_outputs(4526);
    layer1_outputs(3437) <= layer0_outputs(2474);
    layer1_outputs(3438) <= not(layer0_outputs(7075));
    layer1_outputs(3439) <= not(layer0_outputs(528)) or (layer0_outputs(588));
    layer1_outputs(3440) <= '0';
    layer1_outputs(3441) <= not(layer0_outputs(4180));
    layer1_outputs(3442) <= (layer0_outputs(415)) and (layer0_outputs(160));
    layer1_outputs(3443) <= not(layer0_outputs(2773)) or (layer0_outputs(1045));
    layer1_outputs(3444) <= (layer0_outputs(2089)) or (layer0_outputs(111));
    layer1_outputs(3445) <= not(layer0_outputs(454));
    layer1_outputs(3446) <= not((layer0_outputs(5586)) and (layer0_outputs(1192)));
    layer1_outputs(3447) <= not((layer0_outputs(676)) and (layer0_outputs(5998)));
    layer1_outputs(3448) <= not((layer0_outputs(6103)) and (layer0_outputs(3404)));
    layer1_outputs(3449) <= layer0_outputs(2480);
    layer1_outputs(3450) <= (layer0_outputs(5830)) and not (layer0_outputs(4105));
    layer1_outputs(3451) <= layer0_outputs(1855);
    layer1_outputs(3452) <= '1';
    layer1_outputs(3453) <= not((layer0_outputs(3391)) and (layer0_outputs(4039)));
    layer1_outputs(3454) <= not((layer0_outputs(4824)) and (layer0_outputs(5254)));
    layer1_outputs(3455) <= layer0_outputs(5046);
    layer1_outputs(3456) <= not((layer0_outputs(6234)) xor (layer0_outputs(7362)));
    layer1_outputs(3457) <= not(layer0_outputs(6613)) or (layer0_outputs(7461));
    layer1_outputs(3458) <= not((layer0_outputs(6748)) or (layer0_outputs(6954)));
    layer1_outputs(3459) <= (layer0_outputs(6788)) and not (layer0_outputs(3718));
    layer1_outputs(3460) <= not(layer0_outputs(7322));
    layer1_outputs(3461) <= not((layer0_outputs(6345)) and (layer0_outputs(4552)));
    layer1_outputs(3462) <= not(layer0_outputs(3409));
    layer1_outputs(3463) <= '1';
    layer1_outputs(3464) <= (layer0_outputs(3767)) and not (layer0_outputs(835));
    layer1_outputs(3465) <= not(layer0_outputs(5756)) or (layer0_outputs(1151));
    layer1_outputs(3466) <= not(layer0_outputs(6742)) or (layer0_outputs(6230));
    layer1_outputs(3467) <= (layer0_outputs(945)) and not (layer0_outputs(1657));
    layer1_outputs(3468) <= layer0_outputs(4561);
    layer1_outputs(3469) <= not(layer0_outputs(5499)) or (layer0_outputs(1240));
    layer1_outputs(3470) <= (layer0_outputs(1344)) and not (layer0_outputs(2515));
    layer1_outputs(3471) <= not(layer0_outputs(6575));
    layer1_outputs(3472) <= not(layer0_outputs(4396));
    layer1_outputs(3473) <= not((layer0_outputs(4416)) and (layer0_outputs(1524)));
    layer1_outputs(3474) <= not(layer0_outputs(2525)) or (layer0_outputs(4969));
    layer1_outputs(3475) <= '0';
    layer1_outputs(3476) <= (layer0_outputs(327)) or (layer0_outputs(1762));
    layer1_outputs(3477) <= layer0_outputs(7160);
    layer1_outputs(3478) <= layer0_outputs(3369);
    layer1_outputs(3479) <= layer0_outputs(4505);
    layer1_outputs(3480) <= layer0_outputs(5067);
    layer1_outputs(3481) <= (layer0_outputs(2932)) and not (layer0_outputs(598));
    layer1_outputs(3482) <= (layer0_outputs(4521)) and not (layer0_outputs(6224));
    layer1_outputs(3483) <= '1';
    layer1_outputs(3484) <= (layer0_outputs(1227)) and not (layer0_outputs(3546));
    layer1_outputs(3485) <= (layer0_outputs(3783)) or (layer0_outputs(6632));
    layer1_outputs(3486) <= not(layer0_outputs(5913)) or (layer0_outputs(4147));
    layer1_outputs(3487) <= not((layer0_outputs(110)) or (layer0_outputs(2644)));
    layer1_outputs(3488) <= not(layer0_outputs(708)) or (layer0_outputs(3801));
    layer1_outputs(3489) <= '1';
    layer1_outputs(3490) <= (layer0_outputs(3851)) or (layer0_outputs(6844));
    layer1_outputs(3491) <= not(layer0_outputs(4043));
    layer1_outputs(3492) <= layer0_outputs(1074);
    layer1_outputs(3493) <= layer0_outputs(7496);
    layer1_outputs(3494) <= not(layer0_outputs(1618));
    layer1_outputs(3495) <= layer0_outputs(7443);
    layer1_outputs(3496) <= not(layer0_outputs(7152));
    layer1_outputs(3497) <= not(layer0_outputs(2066));
    layer1_outputs(3498) <= (layer0_outputs(4282)) and not (layer0_outputs(1326));
    layer1_outputs(3499) <= (layer0_outputs(3147)) and not (layer0_outputs(7291));
    layer1_outputs(3500) <= layer0_outputs(285);
    layer1_outputs(3501) <= not(layer0_outputs(7520));
    layer1_outputs(3502) <= layer0_outputs(2160);
    layer1_outputs(3503) <= not((layer0_outputs(4694)) and (layer0_outputs(7140)));
    layer1_outputs(3504) <= layer0_outputs(4989);
    layer1_outputs(3505) <= not((layer0_outputs(4449)) or (layer0_outputs(3830)));
    layer1_outputs(3506) <= not(layer0_outputs(6431));
    layer1_outputs(3507) <= not((layer0_outputs(1734)) and (layer0_outputs(409)));
    layer1_outputs(3508) <= (layer0_outputs(5923)) and (layer0_outputs(3565));
    layer1_outputs(3509) <= (layer0_outputs(3173)) or (layer0_outputs(1138));
    layer1_outputs(3510) <= (layer0_outputs(4503)) and (layer0_outputs(5818));
    layer1_outputs(3511) <= layer0_outputs(5032);
    layer1_outputs(3512) <= not(layer0_outputs(4607));
    layer1_outputs(3513) <= (layer0_outputs(7472)) or (layer0_outputs(3676));
    layer1_outputs(3514) <= (layer0_outputs(7168)) and not (layer0_outputs(689));
    layer1_outputs(3515) <= not(layer0_outputs(3505));
    layer1_outputs(3516) <= layer0_outputs(965);
    layer1_outputs(3517) <= '1';
    layer1_outputs(3518) <= '0';
    layer1_outputs(3519) <= not((layer0_outputs(3760)) and (layer0_outputs(6472)));
    layer1_outputs(3520) <= layer0_outputs(3450);
    layer1_outputs(3521) <= (layer0_outputs(1445)) and not (layer0_outputs(4211));
    layer1_outputs(3522) <= (layer0_outputs(3986)) and (layer0_outputs(7451));
    layer1_outputs(3523) <= not(layer0_outputs(6215)) or (layer0_outputs(1818));
    layer1_outputs(3524) <= layer0_outputs(2626);
    layer1_outputs(3525) <= not(layer0_outputs(4083)) or (layer0_outputs(5259));
    layer1_outputs(3526) <= (layer0_outputs(6341)) and not (layer0_outputs(1395));
    layer1_outputs(3527) <= not(layer0_outputs(5806));
    layer1_outputs(3528) <= layer0_outputs(5910);
    layer1_outputs(3529) <= (layer0_outputs(4899)) and not (layer0_outputs(6741));
    layer1_outputs(3530) <= (layer0_outputs(6205)) and not (layer0_outputs(440));
    layer1_outputs(3531) <= layer0_outputs(3415);
    layer1_outputs(3532) <= layer0_outputs(2611);
    layer1_outputs(3533) <= not(layer0_outputs(1567));
    layer1_outputs(3534) <= layer0_outputs(3853);
    layer1_outputs(3535) <= (layer0_outputs(6120)) and not (layer0_outputs(4462));
    layer1_outputs(3536) <= not(layer0_outputs(7030));
    layer1_outputs(3537) <= (layer0_outputs(4223)) or (layer0_outputs(2886));
    layer1_outputs(3538) <= (layer0_outputs(4079)) and not (layer0_outputs(1336));
    layer1_outputs(3539) <= layer0_outputs(130);
    layer1_outputs(3540) <= (layer0_outputs(1533)) or (layer0_outputs(3908));
    layer1_outputs(3541) <= (layer0_outputs(2274)) and not (layer0_outputs(6903));
    layer1_outputs(3542) <= (layer0_outputs(2051)) and (layer0_outputs(6358));
    layer1_outputs(3543) <= not(layer0_outputs(1877));
    layer1_outputs(3544) <= not((layer0_outputs(783)) and (layer0_outputs(1647)));
    layer1_outputs(3545) <= (layer0_outputs(5093)) and (layer0_outputs(3624));
    layer1_outputs(3546) <= not(layer0_outputs(6004));
    layer1_outputs(3547) <= '1';
    layer1_outputs(3548) <= not(layer0_outputs(3102));
    layer1_outputs(3549) <= layer0_outputs(6682);
    layer1_outputs(3550) <= not((layer0_outputs(822)) xor (layer0_outputs(5062)));
    layer1_outputs(3551) <= not(layer0_outputs(3564));
    layer1_outputs(3552) <= layer0_outputs(4866);
    layer1_outputs(3553) <= layer0_outputs(1060);
    layer1_outputs(3554) <= (layer0_outputs(3872)) and not (layer0_outputs(7124));
    layer1_outputs(3555) <= (layer0_outputs(5980)) or (layer0_outputs(4701));
    layer1_outputs(3556) <= (layer0_outputs(4571)) and (layer0_outputs(3886));
    layer1_outputs(3557) <= not(layer0_outputs(4581)) or (layer0_outputs(6355));
    layer1_outputs(3558) <= layer0_outputs(2480);
    layer1_outputs(3559) <= not((layer0_outputs(78)) or (layer0_outputs(2552)));
    layer1_outputs(3560) <= (layer0_outputs(1808)) and (layer0_outputs(4429));
    layer1_outputs(3561) <= not((layer0_outputs(1732)) or (layer0_outputs(3145)));
    layer1_outputs(3562) <= not((layer0_outputs(993)) xor (layer0_outputs(3928)));
    layer1_outputs(3563) <= (layer0_outputs(1669)) and (layer0_outputs(5179));
    layer1_outputs(3564) <= not(layer0_outputs(1619));
    layer1_outputs(3565) <= '1';
    layer1_outputs(3566) <= '0';
    layer1_outputs(3567) <= (layer0_outputs(3846)) xor (layer0_outputs(2546));
    layer1_outputs(3568) <= '1';
    layer1_outputs(3569) <= not(layer0_outputs(3253)) or (layer0_outputs(3205));
    layer1_outputs(3570) <= (layer0_outputs(289)) and not (layer0_outputs(401));
    layer1_outputs(3571) <= not((layer0_outputs(967)) and (layer0_outputs(1211)));
    layer1_outputs(3572) <= not(layer0_outputs(876));
    layer1_outputs(3573) <= not(layer0_outputs(2621));
    layer1_outputs(3574) <= layer0_outputs(6486);
    layer1_outputs(3575) <= layer0_outputs(4181);
    layer1_outputs(3576) <= (layer0_outputs(1788)) xor (layer0_outputs(955));
    layer1_outputs(3577) <= not(layer0_outputs(7489));
    layer1_outputs(3578) <= not(layer0_outputs(2239)) or (layer0_outputs(1733));
    layer1_outputs(3579) <= layer0_outputs(2288);
    layer1_outputs(3580) <= not(layer0_outputs(7025)) or (layer0_outputs(141));
    layer1_outputs(3581) <= not(layer0_outputs(3561)) or (layer0_outputs(4800));
    layer1_outputs(3582) <= (layer0_outputs(3532)) xor (layer0_outputs(6640));
    layer1_outputs(3583) <= not((layer0_outputs(3114)) xor (layer0_outputs(2168)));
    layer1_outputs(3584) <= (layer0_outputs(3493)) xor (layer0_outputs(5027));
    layer1_outputs(3585) <= layer0_outputs(2304);
    layer1_outputs(3586) <= not(layer0_outputs(3391)) or (layer0_outputs(3302));
    layer1_outputs(3587) <= not(layer0_outputs(6974));
    layer1_outputs(3588) <= (layer0_outputs(2088)) and (layer0_outputs(6906));
    layer1_outputs(3589) <= (layer0_outputs(7084)) and (layer0_outputs(4116));
    layer1_outputs(3590) <= not(layer0_outputs(4221)) or (layer0_outputs(1830));
    layer1_outputs(3591) <= (layer0_outputs(4744)) or (layer0_outputs(6421));
    layer1_outputs(3592) <= '1';
    layer1_outputs(3593) <= not(layer0_outputs(3700)) or (layer0_outputs(6378));
    layer1_outputs(3594) <= layer0_outputs(1423);
    layer1_outputs(3595) <= not((layer0_outputs(1537)) or (layer0_outputs(5100)));
    layer1_outputs(3596) <= not(layer0_outputs(2712));
    layer1_outputs(3597) <= (layer0_outputs(2147)) or (layer0_outputs(5492));
    layer1_outputs(3598) <= not(layer0_outputs(4806));
    layer1_outputs(3599) <= '0';
    layer1_outputs(3600) <= not(layer0_outputs(4119));
    layer1_outputs(3601) <= '1';
    layer1_outputs(3602) <= (layer0_outputs(6752)) and (layer0_outputs(3454));
    layer1_outputs(3603) <= '0';
    layer1_outputs(3604) <= '0';
    layer1_outputs(3605) <= (layer0_outputs(3140)) and not (layer0_outputs(4895));
    layer1_outputs(3606) <= layer0_outputs(2955);
    layer1_outputs(3607) <= not(layer0_outputs(3441)) or (layer0_outputs(1614));
    layer1_outputs(3608) <= not(layer0_outputs(4646));
    layer1_outputs(3609) <= layer0_outputs(393);
    layer1_outputs(3610) <= not(layer0_outputs(1986));
    layer1_outputs(3611) <= '1';
    layer1_outputs(3612) <= not(layer0_outputs(3322)) or (layer0_outputs(2513));
    layer1_outputs(3613) <= (layer0_outputs(802)) and (layer0_outputs(4372));
    layer1_outputs(3614) <= '0';
    layer1_outputs(3615) <= layer0_outputs(3969);
    layer1_outputs(3616) <= (layer0_outputs(6606)) and not (layer0_outputs(3459));
    layer1_outputs(3617) <= (layer0_outputs(1783)) and (layer0_outputs(7154));
    layer1_outputs(3618) <= not((layer0_outputs(310)) xor (layer0_outputs(954)));
    layer1_outputs(3619) <= not(layer0_outputs(1883));
    layer1_outputs(3620) <= not(layer0_outputs(3642));
    layer1_outputs(3621) <= layer0_outputs(4862);
    layer1_outputs(3622) <= not(layer0_outputs(4426));
    layer1_outputs(3623) <= not(layer0_outputs(7015)) or (layer0_outputs(5427));
    layer1_outputs(3624) <= not((layer0_outputs(4863)) and (layer0_outputs(827)));
    layer1_outputs(3625) <= '0';
    layer1_outputs(3626) <= (layer0_outputs(1389)) and (layer0_outputs(5684));
    layer1_outputs(3627) <= (layer0_outputs(3109)) and (layer0_outputs(3952));
    layer1_outputs(3628) <= not(layer0_outputs(1868));
    layer1_outputs(3629) <= not(layer0_outputs(5974));
    layer1_outputs(3630) <= '1';
    layer1_outputs(3631) <= '0';
    layer1_outputs(3632) <= layer0_outputs(6883);
    layer1_outputs(3633) <= layer0_outputs(1772);
    layer1_outputs(3634) <= (layer0_outputs(7575)) or (layer0_outputs(172));
    layer1_outputs(3635) <= (layer0_outputs(3044)) and not (layer0_outputs(1158));
    layer1_outputs(3636) <= layer0_outputs(2237);
    layer1_outputs(3637) <= layer0_outputs(6703);
    layer1_outputs(3638) <= '1';
    layer1_outputs(3639) <= not(layer0_outputs(5669));
    layer1_outputs(3640) <= not(layer0_outputs(4089)) or (layer0_outputs(5567));
    layer1_outputs(3641) <= (layer0_outputs(3590)) or (layer0_outputs(5841));
    layer1_outputs(3642) <= not(layer0_outputs(2761));
    layer1_outputs(3643) <= (layer0_outputs(1884)) and not (layer0_outputs(4387));
    layer1_outputs(3644) <= layer0_outputs(3641);
    layer1_outputs(3645) <= (layer0_outputs(1575)) and (layer0_outputs(5346));
    layer1_outputs(3646) <= not((layer0_outputs(1526)) and (layer0_outputs(414)));
    layer1_outputs(3647) <= not((layer0_outputs(5225)) and (layer0_outputs(7581)));
    layer1_outputs(3648) <= not((layer0_outputs(2315)) and (layer0_outputs(1635)));
    layer1_outputs(3649) <= not((layer0_outputs(3320)) or (layer0_outputs(1594)));
    layer1_outputs(3650) <= not(layer0_outputs(7522));
    layer1_outputs(3651) <= not(layer0_outputs(4581));
    layer1_outputs(3652) <= '0';
    layer1_outputs(3653) <= (layer0_outputs(4186)) and (layer0_outputs(2688));
    layer1_outputs(3654) <= not(layer0_outputs(7196)) or (layer0_outputs(2047));
    layer1_outputs(3655) <= not((layer0_outputs(1960)) xor (layer0_outputs(2953)));
    layer1_outputs(3656) <= not(layer0_outputs(7542));
    layer1_outputs(3657) <= not(layer0_outputs(6996));
    layer1_outputs(3658) <= (layer0_outputs(6447)) and (layer0_outputs(2707));
    layer1_outputs(3659) <= layer0_outputs(1952);
    layer1_outputs(3660) <= (layer0_outputs(5413)) and not (layer0_outputs(2981));
    layer1_outputs(3661) <= (layer0_outputs(7171)) or (layer0_outputs(309));
    layer1_outputs(3662) <= not(layer0_outputs(317));
    layer1_outputs(3663) <= (layer0_outputs(6060)) and not (layer0_outputs(1485));
    layer1_outputs(3664) <= not(layer0_outputs(499)) or (layer0_outputs(2553));
    layer1_outputs(3665) <= not((layer0_outputs(3032)) xor (layer0_outputs(1490)));
    layer1_outputs(3666) <= '1';
    layer1_outputs(3667) <= not((layer0_outputs(2623)) and (layer0_outputs(1629)));
    layer1_outputs(3668) <= (layer0_outputs(58)) and (layer0_outputs(4368));
    layer1_outputs(3669) <= not(layer0_outputs(3090));
    layer1_outputs(3670) <= not((layer0_outputs(994)) or (layer0_outputs(7474)));
    layer1_outputs(3671) <= layer0_outputs(430);
    layer1_outputs(3672) <= not(layer0_outputs(1129));
    layer1_outputs(3673) <= not(layer0_outputs(1119));
    layer1_outputs(3674) <= not(layer0_outputs(6232));
    layer1_outputs(3675) <= layer0_outputs(7279);
    layer1_outputs(3676) <= layer0_outputs(7185);
    layer1_outputs(3677) <= not((layer0_outputs(1915)) xor (layer0_outputs(6374)));
    layer1_outputs(3678) <= not((layer0_outputs(4528)) or (layer0_outputs(5818)));
    layer1_outputs(3679) <= not((layer0_outputs(1679)) and (layer0_outputs(6823)));
    layer1_outputs(3680) <= layer0_outputs(4365);
    layer1_outputs(3681) <= not(layer0_outputs(5937)) or (layer0_outputs(5304));
    layer1_outputs(3682) <= not(layer0_outputs(7499));
    layer1_outputs(3683) <= not(layer0_outputs(6502)) or (layer0_outputs(7053));
    layer1_outputs(3684) <= not((layer0_outputs(6077)) or (layer0_outputs(3374)));
    layer1_outputs(3685) <= (layer0_outputs(5003)) and not (layer0_outputs(5490));
    layer1_outputs(3686) <= (layer0_outputs(6596)) and (layer0_outputs(1640));
    layer1_outputs(3687) <= (layer0_outputs(6589)) and (layer0_outputs(2551));
    layer1_outputs(3688) <= (layer0_outputs(7628)) and (layer0_outputs(6961));
    layer1_outputs(3689) <= (layer0_outputs(6717)) and (layer0_outputs(4788));
    layer1_outputs(3690) <= layer0_outputs(5582);
    layer1_outputs(3691) <= (layer0_outputs(4955)) and (layer0_outputs(7513));
    layer1_outputs(3692) <= '1';
    layer1_outputs(3693) <= layer0_outputs(3130);
    layer1_outputs(3694) <= layer0_outputs(4968);
    layer1_outputs(3695) <= (layer0_outputs(5435)) and (layer0_outputs(7561));
    layer1_outputs(3696) <= not(layer0_outputs(2110)) or (layer0_outputs(1834));
    layer1_outputs(3697) <= layer0_outputs(6789);
    layer1_outputs(3698) <= not(layer0_outputs(1357));
    layer1_outputs(3699) <= not(layer0_outputs(7208));
    layer1_outputs(3700) <= (layer0_outputs(291)) and not (layer0_outputs(4185));
    layer1_outputs(3701) <= (layer0_outputs(842)) or (layer0_outputs(5644));
    layer1_outputs(3702) <= not((layer0_outputs(362)) xor (layer0_outputs(7167)));
    layer1_outputs(3703) <= (layer0_outputs(5487)) or (layer0_outputs(5370));
    layer1_outputs(3704) <= not((layer0_outputs(2333)) or (layer0_outputs(2578)));
    layer1_outputs(3705) <= '1';
    layer1_outputs(3706) <= layer0_outputs(4988);
    layer1_outputs(3707) <= not(layer0_outputs(5198)) or (layer0_outputs(7658));
    layer1_outputs(3708) <= not(layer0_outputs(2945));
    layer1_outputs(3709) <= (layer0_outputs(5387)) and not (layer0_outputs(135));
    layer1_outputs(3710) <= (layer0_outputs(374)) and not (layer0_outputs(4630));
    layer1_outputs(3711) <= not(layer0_outputs(1547));
    layer1_outputs(3712) <= '1';
    layer1_outputs(3713) <= (layer0_outputs(7594)) and (layer0_outputs(7378));
    layer1_outputs(3714) <= layer0_outputs(6282);
    layer1_outputs(3715) <= '1';
    layer1_outputs(3716) <= not((layer0_outputs(3597)) or (layer0_outputs(7409)));
    layer1_outputs(3717) <= not((layer0_outputs(2252)) and (layer0_outputs(627)));
    layer1_outputs(3718) <= not((layer0_outputs(5572)) and (layer0_outputs(1505)));
    layer1_outputs(3719) <= not(layer0_outputs(6811)) or (layer0_outputs(1589));
    layer1_outputs(3720) <= not(layer0_outputs(1414)) or (layer0_outputs(4830));
    layer1_outputs(3721) <= not(layer0_outputs(1065)) or (layer0_outputs(3520));
    layer1_outputs(3722) <= (layer0_outputs(2375)) xor (layer0_outputs(6053));
    layer1_outputs(3723) <= (layer0_outputs(238)) xor (layer0_outputs(7467));
    layer1_outputs(3724) <= layer0_outputs(6189);
    layer1_outputs(3725) <= (layer0_outputs(7237)) or (layer0_outputs(4692));
    layer1_outputs(3726) <= (layer0_outputs(4739)) and not (layer0_outputs(5701));
    layer1_outputs(3727) <= '0';
    layer1_outputs(3728) <= (layer0_outputs(159)) and (layer0_outputs(1835));
    layer1_outputs(3729) <= layer0_outputs(7309);
    layer1_outputs(3730) <= (layer0_outputs(203)) and not (layer0_outputs(2772));
    layer1_outputs(3731) <= not(layer0_outputs(4994));
    layer1_outputs(3732) <= not(layer0_outputs(1027));
    layer1_outputs(3733) <= not(layer0_outputs(7650));
    layer1_outputs(3734) <= layer0_outputs(4433);
    layer1_outputs(3735) <= not((layer0_outputs(2550)) or (layer0_outputs(2228)));
    layer1_outputs(3736) <= not(layer0_outputs(2077)) or (layer0_outputs(451));
    layer1_outputs(3737) <= layer0_outputs(7164);
    layer1_outputs(3738) <= not(layer0_outputs(3786)) or (layer0_outputs(2559));
    layer1_outputs(3739) <= '0';
    layer1_outputs(3740) <= not((layer0_outputs(1899)) or (layer0_outputs(354)));
    layer1_outputs(3741) <= (layer0_outputs(5815)) and not (layer0_outputs(1572));
    layer1_outputs(3742) <= not(layer0_outputs(3082));
    layer1_outputs(3743) <= not(layer0_outputs(1342));
    layer1_outputs(3744) <= not(layer0_outputs(2056));
    layer1_outputs(3745) <= not((layer0_outputs(962)) or (layer0_outputs(1758)));
    layer1_outputs(3746) <= not(layer0_outputs(2890)) or (layer0_outputs(6908));
    layer1_outputs(3747) <= (layer0_outputs(3473)) and (layer0_outputs(6057));
    layer1_outputs(3748) <= not((layer0_outputs(2017)) and (layer0_outputs(4127)));
    layer1_outputs(3749) <= not(layer0_outputs(2439));
    layer1_outputs(3750) <= not(layer0_outputs(3693));
    layer1_outputs(3751) <= (layer0_outputs(4273)) xor (layer0_outputs(3792));
    layer1_outputs(3752) <= (layer0_outputs(1220)) and not (layer0_outputs(6852));
    layer1_outputs(3753) <= not(layer0_outputs(1583));
    layer1_outputs(3754) <= (layer0_outputs(6628)) and not (layer0_outputs(36));
    layer1_outputs(3755) <= not(layer0_outputs(1917)) or (layer0_outputs(1427));
    layer1_outputs(3756) <= not(layer0_outputs(3703)) or (layer0_outputs(7615));
    layer1_outputs(3757) <= '1';
    layer1_outputs(3758) <= (layer0_outputs(6738)) and not (layer0_outputs(3077));
    layer1_outputs(3759) <= layer0_outputs(1888);
    layer1_outputs(3760) <= not(layer0_outputs(713));
    layer1_outputs(3761) <= layer0_outputs(4267);
    layer1_outputs(3762) <= layer0_outputs(1721);
    layer1_outputs(3763) <= not(layer0_outputs(2692));
    layer1_outputs(3764) <= not((layer0_outputs(5996)) and (layer0_outputs(2904)));
    layer1_outputs(3765) <= not(layer0_outputs(4452));
    layer1_outputs(3766) <= (layer0_outputs(6213)) and not (layer0_outputs(1425));
    layer1_outputs(3767) <= layer0_outputs(4627);
    layer1_outputs(3768) <= layer0_outputs(512);
    layer1_outputs(3769) <= not((layer0_outputs(2643)) and (layer0_outputs(3171)));
    layer1_outputs(3770) <= not(layer0_outputs(5537));
    layer1_outputs(3771) <= (layer0_outputs(254)) and not (layer0_outputs(2201));
    layer1_outputs(3772) <= not(layer0_outputs(3922)) or (layer0_outputs(7125));
    layer1_outputs(3773) <= (layer0_outputs(4)) and not (layer0_outputs(1546));
    layer1_outputs(3774) <= (layer0_outputs(5676)) and (layer0_outputs(4727));
    layer1_outputs(3775) <= '1';
    layer1_outputs(3776) <= not((layer0_outputs(4405)) or (layer0_outputs(6688)));
    layer1_outputs(3777) <= '0';
    layer1_outputs(3778) <= not((layer0_outputs(2804)) or (layer0_outputs(2090)));
    layer1_outputs(3779) <= not((layer0_outputs(5612)) or (layer0_outputs(124)));
    layer1_outputs(3780) <= not(layer0_outputs(7678)) or (layer0_outputs(898));
    layer1_outputs(3781) <= not(layer0_outputs(174));
    layer1_outputs(3782) <= not(layer0_outputs(919));
    layer1_outputs(3783) <= '0';
    layer1_outputs(3784) <= not(layer0_outputs(935));
    layer1_outputs(3785) <= not(layer0_outputs(5903));
    layer1_outputs(3786) <= not(layer0_outputs(4913));
    layer1_outputs(3787) <= (layer0_outputs(4141)) and (layer0_outputs(3377));
    layer1_outputs(3788) <= not(layer0_outputs(1707));
    layer1_outputs(3789) <= (layer0_outputs(2847)) and not (layer0_outputs(3317));
    layer1_outputs(3790) <= (layer0_outputs(3653)) and not (layer0_outputs(2565));
    layer1_outputs(3791) <= (layer0_outputs(4128)) or (layer0_outputs(7419));
    layer1_outputs(3792) <= layer0_outputs(3755);
    layer1_outputs(3793) <= not(layer0_outputs(2878));
    layer1_outputs(3794) <= (layer0_outputs(7276)) and (layer0_outputs(6612));
    layer1_outputs(3795) <= not((layer0_outputs(1121)) or (layer0_outputs(2265)));
    layer1_outputs(3796) <= '0';
    layer1_outputs(3797) <= (layer0_outputs(6299)) and not (layer0_outputs(7440));
    layer1_outputs(3798) <= not(layer0_outputs(7588)) or (layer0_outputs(1411));
    layer1_outputs(3799) <= '1';
    layer1_outputs(3800) <= layer0_outputs(5591);
    layer1_outputs(3801) <= not(layer0_outputs(657));
    layer1_outputs(3802) <= layer0_outputs(447);
    layer1_outputs(3803) <= not((layer0_outputs(4256)) xor (layer0_outputs(4766)));
    layer1_outputs(3804) <= not(layer0_outputs(953));
    layer1_outputs(3805) <= (layer0_outputs(7094)) or (layer0_outputs(3357));
    layer1_outputs(3806) <= not(layer0_outputs(4133));
    layer1_outputs(3807) <= layer0_outputs(4706);
    layer1_outputs(3808) <= not((layer0_outputs(4158)) or (layer0_outputs(2132)));
    layer1_outputs(3809) <= not(layer0_outputs(4144));
    layer1_outputs(3810) <= layer0_outputs(6314);
    layer1_outputs(3811) <= layer0_outputs(2668);
    layer1_outputs(3812) <= '0';
    layer1_outputs(3813) <= layer0_outputs(4301);
    layer1_outputs(3814) <= (layer0_outputs(5787)) or (layer0_outputs(1975));
    layer1_outputs(3815) <= '1';
    layer1_outputs(3816) <= layer0_outputs(1061);
    layer1_outputs(3817) <= layer0_outputs(6611);
    layer1_outputs(3818) <= (layer0_outputs(5184)) and (layer0_outputs(5659));
    layer1_outputs(3819) <= not(layer0_outputs(4502));
    layer1_outputs(3820) <= not(layer0_outputs(1639));
    layer1_outputs(3821) <= (layer0_outputs(3980)) or (layer0_outputs(2526));
    layer1_outputs(3822) <= '1';
    layer1_outputs(3823) <= not(layer0_outputs(1398)) or (layer0_outputs(3614));
    layer1_outputs(3824) <= not((layer0_outputs(1514)) xor (layer0_outputs(3774)));
    layer1_outputs(3825) <= '0';
    layer1_outputs(3826) <= not(layer0_outputs(1447)) or (layer0_outputs(2723));
    layer1_outputs(3827) <= (layer0_outputs(1930)) or (layer0_outputs(60));
    layer1_outputs(3828) <= (layer0_outputs(3302)) and (layer0_outputs(435));
    layer1_outputs(3829) <= layer0_outputs(847);
    layer1_outputs(3830) <= layer0_outputs(836);
    layer1_outputs(3831) <= (layer0_outputs(2400)) or (layer0_outputs(6109));
    layer1_outputs(3832) <= layer0_outputs(1609);
    layer1_outputs(3833) <= not((layer0_outputs(2507)) and (layer0_outputs(1218)));
    layer1_outputs(3834) <= not(layer0_outputs(2215));
    layer1_outputs(3835) <= not(layer0_outputs(5958));
    layer1_outputs(3836) <= (layer0_outputs(1331)) and not (layer0_outputs(6980));
    layer1_outputs(3837) <= not(layer0_outputs(3664)) or (layer0_outputs(210));
    layer1_outputs(3838) <= not(layer0_outputs(6642)) or (layer0_outputs(6931));
    layer1_outputs(3839) <= not((layer0_outputs(1289)) and (layer0_outputs(4620)));
    layer1_outputs(3840) <= (layer0_outputs(6926)) and not (layer0_outputs(460));
    layer1_outputs(3841) <= '1';
    layer1_outputs(3842) <= not(layer0_outputs(4138)) or (layer0_outputs(5920));
    layer1_outputs(3843) <= not((layer0_outputs(7180)) xor (layer0_outputs(116)));
    layer1_outputs(3844) <= '0';
    layer1_outputs(3845) <= layer0_outputs(6125);
    layer1_outputs(3846) <= (layer0_outputs(7169)) and not (layer0_outputs(3798));
    layer1_outputs(3847) <= not((layer0_outputs(744)) and (layer0_outputs(4760)));
    layer1_outputs(3848) <= (layer0_outputs(4406)) and (layer0_outputs(5411));
    layer1_outputs(3849) <= not((layer0_outputs(2918)) and (layer0_outputs(2673)));
    layer1_outputs(3850) <= (layer0_outputs(6003)) and (layer0_outputs(3542));
    layer1_outputs(3851) <= layer0_outputs(3348);
    layer1_outputs(3852) <= not((layer0_outputs(3670)) or (layer0_outputs(6076)));
    layer1_outputs(3853) <= not(layer0_outputs(6807)) or (layer0_outputs(3648));
    layer1_outputs(3854) <= not((layer0_outputs(2432)) xor (layer0_outputs(2585)));
    layer1_outputs(3855) <= (layer0_outputs(7535)) and (layer0_outputs(2031));
    layer1_outputs(3856) <= (layer0_outputs(655)) or (layer0_outputs(2508));
    layer1_outputs(3857) <= layer0_outputs(1173);
    layer1_outputs(3858) <= (layer0_outputs(7478)) or (layer0_outputs(3689));
    layer1_outputs(3859) <= '0';
    layer1_outputs(3860) <= not((layer0_outputs(3609)) or (layer0_outputs(2420)));
    layer1_outputs(3861) <= layer0_outputs(289);
    layer1_outputs(3862) <= not(layer0_outputs(2563));
    layer1_outputs(3863) <= not(layer0_outputs(4780)) or (layer0_outputs(6797));
    layer1_outputs(3864) <= not(layer0_outputs(2255)) or (layer0_outputs(7289));
    layer1_outputs(3865) <= (layer0_outputs(1200)) and not (layer0_outputs(1427));
    layer1_outputs(3866) <= not(layer0_outputs(5139));
    layer1_outputs(3867) <= not((layer0_outputs(3843)) xor (layer0_outputs(1556)));
    layer1_outputs(3868) <= (layer0_outputs(4583)) or (layer0_outputs(7448));
    layer1_outputs(3869) <= not((layer0_outputs(5539)) or (layer0_outputs(5677)));
    layer1_outputs(3870) <= layer0_outputs(7579);
    layer1_outputs(3871) <= not(layer0_outputs(6981)) or (layer0_outputs(5564));
    layer1_outputs(3872) <= (layer0_outputs(242)) and (layer0_outputs(5241));
    layer1_outputs(3873) <= (layer0_outputs(2397)) and not (layer0_outputs(4652));
    layer1_outputs(3874) <= not(layer0_outputs(240)) or (layer0_outputs(7239));
    layer1_outputs(3875) <= not((layer0_outputs(4660)) and (layer0_outputs(1760)));
    layer1_outputs(3876) <= (layer0_outputs(5866)) and not (layer0_outputs(6107));
    layer1_outputs(3877) <= not(layer0_outputs(1265));
    layer1_outputs(3878) <= not(layer0_outputs(4889));
    layer1_outputs(3879) <= layer0_outputs(674);
    layer1_outputs(3880) <= not(layer0_outputs(3691));
    layer1_outputs(3881) <= not(layer0_outputs(4939));
    layer1_outputs(3882) <= (layer0_outputs(7337)) and not (layer0_outputs(6604));
    layer1_outputs(3883) <= (layer0_outputs(7460)) and not (layer0_outputs(7252));
    layer1_outputs(3884) <= not(layer0_outputs(763)) or (layer0_outputs(6941));
    layer1_outputs(3885) <= not((layer0_outputs(4821)) and (layer0_outputs(4666)));
    layer1_outputs(3886) <= not(layer0_outputs(2011));
    layer1_outputs(3887) <= (layer0_outputs(3717)) or (layer0_outputs(7318));
    layer1_outputs(3888) <= layer0_outputs(5142);
    layer1_outputs(3889) <= not((layer0_outputs(6917)) and (layer0_outputs(4866)));
    layer1_outputs(3890) <= not(layer0_outputs(3354)) or (layer0_outputs(2384));
    layer1_outputs(3891) <= layer0_outputs(4854);
    layer1_outputs(3892) <= layer0_outputs(4684);
    layer1_outputs(3893) <= not(layer0_outputs(453)) or (layer0_outputs(2671));
    layer1_outputs(3894) <= not(layer0_outputs(2813)) or (layer0_outputs(5341));
    layer1_outputs(3895) <= layer0_outputs(1762);
    layer1_outputs(3896) <= (layer0_outputs(754)) and not (layer0_outputs(2600));
    layer1_outputs(3897) <= layer0_outputs(3730);
    layer1_outputs(3898) <= layer0_outputs(5426);
    layer1_outputs(3899) <= not((layer0_outputs(3937)) or (layer0_outputs(1181)));
    layer1_outputs(3900) <= (layer0_outputs(275)) and not (layer0_outputs(4193));
    layer1_outputs(3901) <= not((layer0_outputs(7173)) and (layer0_outputs(3189)));
    layer1_outputs(3902) <= layer0_outputs(4875);
    layer1_outputs(3903) <= '0';
    layer1_outputs(3904) <= not(layer0_outputs(7288));
    layer1_outputs(3905) <= (layer0_outputs(5429)) and not (layer0_outputs(4442));
    layer1_outputs(3906) <= (layer0_outputs(653)) and not (layer0_outputs(7462));
    layer1_outputs(3907) <= not(layer0_outputs(4480)) or (layer0_outputs(7495));
    layer1_outputs(3908) <= layer0_outputs(5178);
    layer1_outputs(3909) <= not(layer0_outputs(3917));
    layer1_outputs(3910) <= not(layer0_outputs(5605)) or (layer0_outputs(3192));
    layer1_outputs(3911) <= (layer0_outputs(392)) and (layer0_outputs(4594));
    layer1_outputs(3912) <= not((layer0_outputs(6385)) or (layer0_outputs(6610)));
    layer1_outputs(3913) <= not(layer0_outputs(3136));
    layer1_outputs(3914) <= not(layer0_outputs(1655));
    layer1_outputs(3915) <= layer0_outputs(6288);
    layer1_outputs(3916) <= not((layer0_outputs(6832)) xor (layer0_outputs(2528)));
    layer1_outputs(3917) <= '1';
    layer1_outputs(3918) <= not((layer0_outputs(720)) xor (layer0_outputs(4965)));
    layer1_outputs(3919) <= not((layer0_outputs(3271)) and (layer0_outputs(4783)));
    layer1_outputs(3920) <= not((layer0_outputs(4041)) or (layer0_outputs(7631)));
    layer1_outputs(3921) <= not(layer0_outputs(1342)) or (layer0_outputs(1170));
    layer1_outputs(3922) <= not(layer0_outputs(4242));
    layer1_outputs(3923) <= layer0_outputs(7124);
    layer1_outputs(3924) <= layer0_outputs(5660);
    layer1_outputs(3925) <= (layer0_outputs(6892)) and (layer0_outputs(4126));
    layer1_outputs(3926) <= layer0_outputs(5931);
    layer1_outputs(3927) <= not(layer0_outputs(7303));
    layer1_outputs(3928) <= not(layer0_outputs(2292)) or (layer0_outputs(3221));
    layer1_outputs(3929) <= not(layer0_outputs(7153));
    layer1_outputs(3930) <= layer0_outputs(6501);
    layer1_outputs(3931) <= not(layer0_outputs(2808));
    layer1_outputs(3932) <= not(layer0_outputs(4434)) or (layer0_outputs(7246));
    layer1_outputs(3933) <= not(layer0_outputs(7274));
    layer1_outputs(3934) <= (layer0_outputs(2827)) or (layer0_outputs(3947));
    layer1_outputs(3935) <= layer0_outputs(5665);
    layer1_outputs(3936) <= not((layer0_outputs(1690)) or (layer0_outputs(7396)));
    layer1_outputs(3937) <= layer0_outputs(3290);
    layer1_outputs(3938) <= not((layer0_outputs(2785)) or (layer0_outputs(5073)));
    layer1_outputs(3939) <= (layer0_outputs(3071)) or (layer0_outputs(669));
    layer1_outputs(3940) <= not(layer0_outputs(751)) or (layer0_outputs(359));
    layer1_outputs(3941) <= (layer0_outputs(7629)) and not (layer0_outputs(4140));
    layer1_outputs(3942) <= (layer0_outputs(5174)) or (layer0_outputs(5445));
    layer1_outputs(3943) <= (layer0_outputs(6161)) and not (layer0_outputs(4208));
    layer1_outputs(3944) <= layer0_outputs(4848);
    layer1_outputs(3945) <= layer0_outputs(7672);
    layer1_outputs(3946) <= (layer0_outputs(2142)) and (layer0_outputs(4525));
    layer1_outputs(3947) <= not(layer0_outputs(1167));
    layer1_outputs(3948) <= layer0_outputs(3016);
    layer1_outputs(3949) <= not((layer0_outputs(6719)) or (layer0_outputs(6031)));
    layer1_outputs(3950) <= layer0_outputs(1382);
    layer1_outputs(3951) <= not((layer0_outputs(3521)) or (layer0_outputs(5171)));
    layer1_outputs(3952) <= not(layer0_outputs(281));
    layer1_outputs(3953) <= not(layer0_outputs(5311));
    layer1_outputs(3954) <= layer0_outputs(3586);
    layer1_outputs(3955) <= not(layer0_outputs(2975)) or (layer0_outputs(4486));
    layer1_outputs(3956) <= (layer0_outputs(5153)) and (layer0_outputs(5593));
    layer1_outputs(3957) <= not(layer0_outputs(4167)) or (layer0_outputs(6245));
    layer1_outputs(3958) <= not(layer0_outputs(6638)) or (layer0_outputs(2306));
    layer1_outputs(3959) <= (layer0_outputs(2436)) and (layer0_outputs(3407));
    layer1_outputs(3960) <= layer0_outputs(4215);
    layer1_outputs(3961) <= (layer0_outputs(491)) and not (layer0_outputs(482));
    layer1_outputs(3962) <= layer0_outputs(1422);
    layer1_outputs(3963) <= layer0_outputs(2147);
    layer1_outputs(3964) <= '1';
    layer1_outputs(3965) <= not(layer0_outputs(2755)) or (layer0_outputs(5797));
    layer1_outputs(3966) <= not(layer0_outputs(6016));
    layer1_outputs(3967) <= (layer0_outputs(2299)) and (layer0_outputs(997));
    layer1_outputs(3968) <= layer0_outputs(348);
    layer1_outputs(3969) <= not(layer0_outputs(4702)) or (layer0_outputs(5496));
    layer1_outputs(3970) <= not(layer0_outputs(5740));
    layer1_outputs(3971) <= not(layer0_outputs(2704));
    layer1_outputs(3972) <= (layer0_outputs(3808)) and (layer0_outputs(6427));
    layer1_outputs(3973) <= not((layer0_outputs(5169)) and (layer0_outputs(4225)));
    layer1_outputs(3974) <= not((layer0_outputs(3232)) or (layer0_outputs(1665)));
    layer1_outputs(3975) <= not(layer0_outputs(2313));
    layer1_outputs(3976) <= (layer0_outputs(564)) or (layer0_outputs(6535));
    layer1_outputs(3977) <= layer0_outputs(2137);
    layer1_outputs(3978) <= (layer0_outputs(7486)) and not (layer0_outputs(4543));
    layer1_outputs(3979) <= (layer0_outputs(7212)) or (layer0_outputs(7239));
    layer1_outputs(3980) <= layer0_outputs(438);
    layer1_outputs(3981) <= (layer0_outputs(6090)) and not (layer0_outputs(2320));
    layer1_outputs(3982) <= (layer0_outputs(4451)) and not (layer0_outputs(2063));
    layer1_outputs(3983) <= (layer0_outputs(4978)) and not (layer0_outputs(6255));
    layer1_outputs(3984) <= '0';
    layer1_outputs(3985) <= (layer0_outputs(3258)) and not (layer0_outputs(6479));
    layer1_outputs(3986) <= not((layer0_outputs(3563)) and (layer0_outputs(1742)));
    layer1_outputs(3987) <= not(layer0_outputs(1247));
    layer1_outputs(3988) <= not(layer0_outputs(4226)) or (layer0_outputs(4617));
    layer1_outputs(3989) <= (layer0_outputs(4455)) and not (layer0_outputs(6820));
    layer1_outputs(3990) <= layer0_outputs(2518);
    layer1_outputs(3991) <= layer0_outputs(2845);
    layer1_outputs(3992) <= not(layer0_outputs(2737));
    layer1_outputs(3993) <= not((layer0_outputs(68)) or (layer0_outputs(6217)));
    layer1_outputs(3994) <= (layer0_outputs(4673)) xor (layer0_outputs(5611));
    layer1_outputs(3995) <= (layer0_outputs(1663)) xor (layer0_outputs(2026));
    layer1_outputs(3996) <= not(layer0_outputs(3292));
    layer1_outputs(3997) <= not(layer0_outputs(1766));
    layer1_outputs(3998) <= (layer0_outputs(7031)) and (layer0_outputs(3600));
    layer1_outputs(3999) <= (layer0_outputs(4410)) and (layer0_outputs(2317));
    layer1_outputs(4000) <= layer0_outputs(4896);
    layer1_outputs(4001) <= layer0_outputs(7235);
    layer1_outputs(4002) <= not(layer0_outputs(978)) or (layer0_outputs(5878));
    layer1_outputs(4003) <= (layer0_outputs(5382)) and not (layer0_outputs(2217));
    layer1_outputs(4004) <= not(layer0_outputs(4217));
    layer1_outputs(4005) <= not(layer0_outputs(5795));
    layer1_outputs(4006) <= not(layer0_outputs(2144)) or (layer0_outputs(1462));
    layer1_outputs(4007) <= not(layer0_outputs(4520));
    layer1_outputs(4008) <= '1';
    layer1_outputs(4009) <= (layer0_outputs(7321)) and (layer0_outputs(7391));
    layer1_outputs(4010) <= (layer0_outputs(4326)) xor (layer0_outputs(7574));
    layer1_outputs(4011) <= (layer0_outputs(2390)) and (layer0_outputs(2174));
    layer1_outputs(4012) <= not((layer0_outputs(1973)) and (layer0_outputs(75)));
    layer1_outputs(4013) <= (layer0_outputs(7172)) and not (layer0_outputs(3554));
    layer1_outputs(4014) <= (layer0_outputs(3325)) and not (layer0_outputs(1043));
    layer1_outputs(4015) <= '0';
    layer1_outputs(4016) <= (layer0_outputs(1587)) and (layer0_outputs(3157));
    layer1_outputs(4017) <= (layer0_outputs(877)) or (layer0_outputs(7659));
    layer1_outputs(4018) <= layer0_outputs(6949);
    layer1_outputs(4019) <= (layer0_outputs(1331)) and (layer0_outputs(331));
    layer1_outputs(4020) <= not(layer0_outputs(7265));
    layer1_outputs(4021) <= (layer0_outputs(5905)) and not (layer0_outputs(2437));
    layer1_outputs(4022) <= layer0_outputs(4878);
    layer1_outputs(4023) <= (layer0_outputs(1576)) and not (layer0_outputs(2744));
    layer1_outputs(4024) <= (layer0_outputs(2000)) or (layer0_outputs(6919));
    layer1_outputs(4025) <= not(layer0_outputs(7047)) or (layer0_outputs(2990));
    layer1_outputs(4026) <= not(layer0_outputs(278)) or (layer0_outputs(2230));
    layer1_outputs(4027) <= not((layer0_outputs(4355)) and (layer0_outputs(5740)));
    layer1_outputs(4028) <= layer0_outputs(7445);
    layer1_outputs(4029) <= (layer0_outputs(3449)) and (layer0_outputs(3855));
    layer1_outputs(4030) <= not((layer0_outputs(5248)) and (layer0_outputs(7079)));
    layer1_outputs(4031) <= (layer0_outputs(1615)) and (layer0_outputs(1258));
    layer1_outputs(4032) <= (layer0_outputs(3223)) or (layer0_outputs(6064));
    layer1_outputs(4033) <= not(layer0_outputs(4768));
    layer1_outputs(4034) <= not(layer0_outputs(2260));
    layer1_outputs(4035) <= (layer0_outputs(3553)) and not (layer0_outputs(2394));
    layer1_outputs(4036) <= (layer0_outputs(973)) and not (layer0_outputs(2687));
    layer1_outputs(4037) <= not(layer0_outputs(6096));
    layer1_outputs(4038) <= (layer0_outputs(7299)) and not (layer0_outputs(1059));
    layer1_outputs(4039) <= layer0_outputs(5563);
    layer1_outputs(4040) <= not(layer0_outputs(5221));
    layer1_outputs(4041) <= '0';
    layer1_outputs(4042) <= not(layer0_outputs(6905)) or (layer0_outputs(3475));
    layer1_outputs(4043) <= (layer0_outputs(6497)) and not (layer0_outputs(7156));
    layer1_outputs(4044) <= (layer0_outputs(1929)) and not (layer0_outputs(5720));
    layer1_outputs(4045) <= '1';
    layer1_outputs(4046) <= layer0_outputs(5398);
    layer1_outputs(4047) <= (layer0_outputs(2540)) or (layer0_outputs(5204));
    layer1_outputs(4048) <= (layer0_outputs(6169)) or (layer0_outputs(4070));
    layer1_outputs(4049) <= layer0_outputs(6298);
    layer1_outputs(4050) <= layer0_outputs(4658);
    layer1_outputs(4051) <= layer0_outputs(204);
    layer1_outputs(4052) <= (layer0_outputs(1112)) or (layer0_outputs(6935));
    layer1_outputs(4053) <= '1';
    layer1_outputs(4054) <= (layer0_outputs(6747)) or (layer0_outputs(2757));
    layer1_outputs(4055) <= not(layer0_outputs(3512)) or (layer0_outputs(6908));
    layer1_outputs(4056) <= (layer0_outputs(3423)) and not (layer0_outputs(1246));
    layer1_outputs(4057) <= '0';
    layer1_outputs(4058) <= layer0_outputs(4736);
    layer1_outputs(4059) <= layer0_outputs(1515);
    layer1_outputs(4060) <= not(layer0_outputs(866));
    layer1_outputs(4061) <= (layer0_outputs(6542)) and not (layer0_outputs(6949));
    layer1_outputs(4062) <= not((layer0_outputs(5867)) or (layer0_outputs(388)));
    layer1_outputs(4063) <= layer0_outputs(1169);
    layer1_outputs(4064) <= not(layer0_outputs(5123));
    layer1_outputs(4065) <= not((layer0_outputs(2483)) or (layer0_outputs(1042)));
    layer1_outputs(4066) <= (layer0_outputs(6150)) and not (layer0_outputs(1446));
    layer1_outputs(4067) <= layer0_outputs(4259);
    layer1_outputs(4068) <= not(layer0_outputs(6233)) or (layer0_outputs(2396));
    layer1_outputs(4069) <= layer0_outputs(1195);
    layer1_outputs(4070) <= (layer0_outputs(2699)) and (layer0_outputs(5804));
    layer1_outputs(4071) <= layer0_outputs(6054);
    layer1_outputs(4072) <= not(layer0_outputs(4749)) or (layer0_outputs(5203));
    layer1_outputs(4073) <= not(layer0_outputs(4704)) or (layer0_outputs(5026));
    layer1_outputs(4074) <= (layer0_outputs(1563)) and not (layer0_outputs(1426));
    layer1_outputs(4075) <= (layer0_outputs(149)) and (layer0_outputs(5148));
    layer1_outputs(4076) <= not(layer0_outputs(4745));
    layer1_outputs(4077) <= '1';
    layer1_outputs(4078) <= layer0_outputs(3603);
    layer1_outputs(4079) <= (layer0_outputs(4063)) or (layer0_outputs(5163));
    layer1_outputs(4080) <= '1';
    layer1_outputs(4081) <= not(layer0_outputs(4441));
    layer1_outputs(4082) <= not((layer0_outputs(1393)) and (layer0_outputs(4288)));
    layer1_outputs(4083) <= (layer0_outputs(3777)) and not (layer0_outputs(6395));
    layer1_outputs(4084) <= '1';
    layer1_outputs(4085) <= '0';
    layer1_outputs(4086) <= '1';
    layer1_outputs(4087) <= not((layer0_outputs(1267)) xor (layer0_outputs(4178)));
    layer1_outputs(4088) <= '0';
    layer1_outputs(4089) <= not(layer0_outputs(5351)) or (layer0_outputs(1337));
    layer1_outputs(4090) <= not(layer0_outputs(4331)) or (layer0_outputs(6160));
    layer1_outputs(4091) <= layer0_outputs(3918);
    layer1_outputs(4092) <= not(layer0_outputs(2678));
    layer1_outputs(4093) <= layer0_outputs(2080);
    layer1_outputs(4094) <= (layer0_outputs(7430)) and (layer0_outputs(1854));
    layer1_outputs(4095) <= (layer0_outputs(3304)) or (layer0_outputs(4850));
    layer1_outputs(4096) <= (layer0_outputs(1329)) and not (layer0_outputs(2880));
    layer1_outputs(4097) <= layer0_outputs(3703);
    layer1_outputs(4098) <= not((layer0_outputs(4408)) or (layer0_outputs(1608)));
    layer1_outputs(4099) <= layer0_outputs(2045);
    layer1_outputs(4100) <= (layer0_outputs(554)) and (layer0_outputs(1149));
    layer1_outputs(4101) <= not(layer0_outputs(7674));
    layer1_outputs(4102) <= not(layer0_outputs(6027));
    layer1_outputs(4103) <= not(layer0_outputs(5952));
    layer1_outputs(4104) <= (layer0_outputs(3751)) or (layer0_outputs(3981));
    layer1_outputs(4105) <= not(layer0_outputs(7447)) or (layer0_outputs(3638));
    layer1_outputs(4106) <= not((layer0_outputs(3007)) and (layer0_outputs(6616)));
    layer1_outputs(4107) <= not((layer0_outputs(4118)) and (layer0_outputs(1446)));
    layer1_outputs(4108) <= (layer0_outputs(883)) and not (layer0_outputs(4756));
    layer1_outputs(4109) <= not((layer0_outputs(3776)) and (layer0_outputs(3042)));
    layer1_outputs(4110) <= '1';
    layer1_outputs(4111) <= not(layer0_outputs(6977));
    layer1_outputs(4112) <= '1';
    layer1_outputs(4113) <= not((layer0_outputs(5955)) and (layer0_outputs(1857)));
    layer1_outputs(4114) <= not((layer0_outputs(7117)) and (layer0_outputs(3330)));
    layer1_outputs(4115) <= not(layer0_outputs(4342)) or (layer0_outputs(4177));
    layer1_outputs(4116) <= not(layer0_outputs(3341)) or (layer0_outputs(7367));
    layer1_outputs(4117) <= not(layer0_outputs(90));
    layer1_outputs(4118) <= not(layer0_outputs(2411)) or (layer0_outputs(7512));
    layer1_outputs(4119) <= (layer0_outputs(2533)) or (layer0_outputs(4048));
    layer1_outputs(4120) <= (layer0_outputs(7371)) or (layer0_outputs(4148));
    layer1_outputs(4121) <= not((layer0_outputs(5836)) xor (layer0_outputs(216)));
    layer1_outputs(4122) <= not(layer0_outputs(5138));
    layer1_outputs(4123) <= (layer0_outputs(1929)) xor (layer0_outputs(206));
    layer1_outputs(4124) <= layer0_outputs(1594);
    layer1_outputs(4125) <= layer0_outputs(419);
    layer1_outputs(4126) <= '1';
    layer1_outputs(4127) <= (layer0_outputs(6269)) and not (layer0_outputs(6819));
    layer1_outputs(4128) <= layer0_outputs(3180);
    layer1_outputs(4129) <= not(layer0_outputs(5507));
    layer1_outputs(4130) <= not((layer0_outputs(7170)) or (layer0_outputs(6094)));
    layer1_outputs(4131) <= layer0_outputs(1079);
    layer1_outputs(4132) <= (layer0_outputs(6602)) and (layer0_outputs(2588));
    layer1_outputs(4133) <= (layer0_outputs(951)) and not (layer0_outputs(4528));
    layer1_outputs(4134) <= (layer0_outputs(4847)) and (layer0_outputs(5146));
    layer1_outputs(4135) <= not((layer0_outputs(5525)) xor (layer0_outputs(4323)));
    layer1_outputs(4136) <= '0';
    layer1_outputs(4137) <= not(layer0_outputs(7327));
    layer1_outputs(4138) <= not(layer0_outputs(1456));
    layer1_outputs(4139) <= not(layer0_outputs(5096));
    layer1_outputs(4140) <= not((layer0_outputs(3955)) and (layer0_outputs(6942)));
    layer1_outputs(4141) <= '1';
    layer1_outputs(4142) <= layer0_outputs(6129);
    layer1_outputs(4143) <= not(layer0_outputs(2992));
    layer1_outputs(4144) <= (layer0_outputs(7648)) and not (layer0_outputs(629));
    layer1_outputs(4145) <= (layer0_outputs(3417)) and not (layer0_outputs(7165));
    layer1_outputs(4146) <= not((layer0_outputs(6615)) xor (layer0_outputs(5771)));
    layer1_outputs(4147) <= layer0_outputs(5556);
    layer1_outputs(4148) <= not((layer0_outputs(2244)) and (layer0_outputs(899)));
    layer1_outputs(4149) <= (layer0_outputs(305)) or (layer0_outputs(5702));
    layer1_outputs(4150) <= not(layer0_outputs(728));
    layer1_outputs(4151) <= (layer0_outputs(1621)) or (layer0_outputs(69));
    layer1_outputs(4152) <= not((layer0_outputs(4114)) and (layer0_outputs(263)));
    layer1_outputs(4153) <= layer0_outputs(2893);
    layer1_outputs(4154) <= not(layer0_outputs(2411)) or (layer0_outputs(177));
    layer1_outputs(4155) <= not(layer0_outputs(7210)) or (layer0_outputs(35));
    layer1_outputs(4156) <= (layer0_outputs(91)) and not (layer0_outputs(6316));
    layer1_outputs(4157) <= not(layer0_outputs(1299)) or (layer0_outputs(687));
    layer1_outputs(4158) <= not(layer0_outputs(2560));
    layer1_outputs(4159) <= (layer0_outputs(198)) and (layer0_outputs(1051));
    layer1_outputs(4160) <= (layer0_outputs(3598)) and not (layer0_outputs(949));
    layer1_outputs(4161) <= not(layer0_outputs(4919)) or (layer0_outputs(1046));
    layer1_outputs(4162) <= layer0_outputs(3510);
    layer1_outputs(4163) <= not(layer0_outputs(3061));
    layer1_outputs(4164) <= not((layer0_outputs(3467)) or (layer0_outputs(4366)));
    layer1_outputs(4165) <= (layer0_outputs(6668)) and not (layer0_outputs(5043));
    layer1_outputs(4166) <= (layer0_outputs(2100)) and (layer0_outputs(4923));
    layer1_outputs(4167) <= not(layer0_outputs(4505));
    layer1_outputs(4168) <= not(layer0_outputs(1387)) or (layer0_outputs(6805));
    layer1_outputs(4169) <= not(layer0_outputs(4426)) or (layer0_outputs(339));
    layer1_outputs(4170) <= layer0_outputs(1227);
    layer1_outputs(4171) <= (layer0_outputs(1960)) or (layer0_outputs(2131));
    layer1_outputs(4172) <= not(layer0_outputs(608));
    layer1_outputs(4173) <= layer0_outputs(2010);
    layer1_outputs(4174) <= not(layer0_outputs(5494)) or (layer0_outputs(2617));
    layer1_outputs(4175) <= not(layer0_outputs(5306));
    layer1_outputs(4176) <= not(layer0_outputs(3634));
    layer1_outputs(4177) <= not((layer0_outputs(6784)) and (layer0_outputs(3544)));
    layer1_outputs(4178) <= not((layer0_outputs(3658)) or (layer0_outputs(1509)));
    layer1_outputs(4179) <= layer0_outputs(3113);
    layer1_outputs(4180) <= not(layer0_outputs(7557));
    layer1_outputs(4181) <= not(layer0_outputs(4465)) or (layer0_outputs(7404));
    layer1_outputs(4182) <= not(layer0_outputs(1693));
    layer1_outputs(4183) <= not((layer0_outputs(7055)) and (layer0_outputs(2056)));
    layer1_outputs(4184) <= layer0_outputs(7135);
    layer1_outputs(4185) <= '1';
    layer1_outputs(4186) <= not((layer0_outputs(3957)) or (layer0_outputs(1581)));
    layer1_outputs(4187) <= layer0_outputs(5498);
    layer1_outputs(4188) <= (layer0_outputs(3888)) and not (layer0_outputs(5667));
    layer1_outputs(4189) <= not(layer0_outputs(6397)) or (layer0_outputs(1573));
    layer1_outputs(4190) <= not((layer0_outputs(5385)) and (layer0_outputs(5064)));
    layer1_outputs(4191) <= (layer0_outputs(7260)) and not (layer0_outputs(4115));
    layer1_outputs(4192) <= '1';
    layer1_outputs(4193) <= '0';
    layer1_outputs(4194) <= not(layer0_outputs(1044)) or (layer0_outputs(7018));
    layer1_outputs(4195) <= not((layer0_outputs(3974)) or (layer0_outputs(5312)));
    layer1_outputs(4196) <= '0';
    layer1_outputs(4197) <= layer0_outputs(6769);
    layer1_outputs(4198) <= not(layer0_outputs(2579)) or (layer0_outputs(7292));
    layer1_outputs(4199) <= not(layer0_outputs(6998)) or (layer0_outputs(4953));
    layer1_outputs(4200) <= layer0_outputs(904);
    layer1_outputs(4201) <= not(layer0_outputs(347)) or (layer0_outputs(678));
    layer1_outputs(4202) <= layer0_outputs(6651);
    layer1_outputs(4203) <= (layer0_outputs(3476)) or (layer0_outputs(5208));
    layer1_outputs(4204) <= layer0_outputs(5387);
    layer1_outputs(4205) <= (layer0_outputs(5516)) and not (layer0_outputs(722));
    layer1_outputs(4206) <= layer0_outputs(1642);
    layer1_outputs(4207) <= not(layer0_outputs(4344)) or (layer0_outputs(3120));
    layer1_outputs(4208) <= (layer0_outputs(5361)) and (layer0_outputs(6029));
    layer1_outputs(4209) <= (layer0_outputs(2693)) or (layer0_outputs(6063));
    layer1_outputs(4210) <= (layer0_outputs(6260)) and not (layer0_outputs(7487));
    layer1_outputs(4211) <= '0';
    layer1_outputs(4212) <= not((layer0_outputs(3411)) and (layer0_outputs(1428)));
    layer1_outputs(4213) <= (layer0_outputs(3836)) or (layer0_outputs(2962));
    layer1_outputs(4214) <= (layer0_outputs(1175)) and not (layer0_outputs(7533));
    layer1_outputs(4215) <= not(layer0_outputs(3470)) or (layer0_outputs(5861));
    layer1_outputs(4216) <= not(layer0_outputs(2326)) or (layer0_outputs(839));
    layer1_outputs(4217) <= (layer0_outputs(7367)) xor (layer0_outputs(6193));
    layer1_outputs(4218) <= (layer0_outputs(1373)) and not (layer0_outputs(5816));
    layer1_outputs(4219) <= '1';
    layer1_outputs(4220) <= (layer0_outputs(5452)) and not (layer0_outputs(4450));
    layer1_outputs(4221) <= layer0_outputs(3917);
    layer1_outputs(4222) <= '0';
    layer1_outputs(4223) <= layer0_outputs(5714);
    layer1_outputs(4224) <= (layer0_outputs(2770)) and (layer0_outputs(1948));
    layer1_outputs(4225) <= (layer0_outputs(7380)) and not (layer0_outputs(5407));
    layer1_outputs(4226) <= layer0_outputs(581);
    layer1_outputs(4227) <= layer0_outputs(7250);
    layer1_outputs(4228) <= not((layer0_outputs(3415)) and (layer0_outputs(63)));
    layer1_outputs(4229) <= (layer0_outputs(1314)) or (layer0_outputs(567));
    layer1_outputs(4230) <= '1';
    layer1_outputs(4231) <= (layer0_outputs(3272)) and not (layer0_outputs(1176));
    layer1_outputs(4232) <= (layer0_outputs(1995)) and not (layer0_outputs(4860));
    layer1_outputs(4233) <= (layer0_outputs(5697)) and not (layer0_outputs(3970));
    layer1_outputs(4234) <= not((layer0_outputs(1662)) and (layer0_outputs(4916)));
    layer1_outputs(4235) <= layer0_outputs(1620);
    layer1_outputs(4236) <= '1';
    layer1_outputs(4237) <= not(layer0_outputs(5720));
    layer1_outputs(4238) <= not((layer0_outputs(1177)) or (layer0_outputs(1415)));
    layer1_outputs(4239) <= (layer0_outputs(3350)) and not (layer0_outputs(5573));
    layer1_outputs(4240) <= not((layer0_outputs(2384)) xor (layer0_outputs(1196)));
    layer1_outputs(4241) <= not(layer0_outputs(4644));
    layer1_outputs(4242) <= not(layer0_outputs(3074));
    layer1_outputs(4243) <= not(layer0_outputs(1518));
    layer1_outputs(4244) <= (layer0_outputs(12)) xor (layer0_outputs(486));
    layer1_outputs(4245) <= not(layer0_outputs(868));
    layer1_outputs(4246) <= layer0_outputs(838);
    layer1_outputs(4247) <= layer0_outputs(5051);
    layer1_outputs(4248) <= (layer0_outputs(2227)) and (layer0_outputs(3989));
    layer1_outputs(4249) <= layer0_outputs(75);
    layer1_outputs(4250) <= '0';
    layer1_outputs(4251) <= (layer0_outputs(6236)) xor (layer0_outputs(2958));
    layer1_outputs(4252) <= (layer0_outputs(7388)) and (layer0_outputs(2994));
    layer1_outputs(4253) <= (layer0_outputs(4716)) and (layer0_outputs(6669));
    layer1_outputs(4254) <= '1';
    layer1_outputs(4255) <= (layer0_outputs(1790)) or (layer0_outputs(4926));
    layer1_outputs(4256) <= (layer0_outputs(5917)) or (layer0_outputs(388));
    layer1_outputs(4257) <= (layer0_outputs(2115)) and not (layer0_outputs(5010));
    layer1_outputs(4258) <= layer0_outputs(4228);
    layer1_outputs(4259) <= layer0_outputs(477);
    layer1_outputs(4260) <= (layer0_outputs(3815)) and not (layer0_outputs(6381));
    layer1_outputs(4261) <= (layer0_outputs(1996)) and (layer0_outputs(1625));
    layer1_outputs(4262) <= not(layer0_outputs(541));
    layer1_outputs(4263) <= '1';
    layer1_outputs(4264) <= not(layer0_outputs(1820)) or (layer0_outputs(1124));
    layer1_outputs(4265) <= not(layer0_outputs(2931)) or (layer0_outputs(2057));
    layer1_outputs(4266) <= (layer0_outputs(7221)) and not (layer0_outputs(7644));
    layer1_outputs(4267) <= (layer0_outputs(5346)) and not (layer0_outputs(5215));
    layer1_outputs(4268) <= not(layer0_outputs(6948)) or (layer0_outputs(5327));
    layer1_outputs(4269) <= '1';
    layer1_outputs(4270) <= (layer0_outputs(4382)) or (layer0_outputs(2179));
    layer1_outputs(4271) <= '1';
    layer1_outputs(4272) <= layer0_outputs(6090);
    layer1_outputs(4273) <= not((layer0_outputs(7479)) or (layer0_outputs(4378)));
    layer1_outputs(4274) <= not(layer0_outputs(4275)) or (layer0_outputs(228));
    layer1_outputs(4275) <= not(layer0_outputs(3135));
    layer1_outputs(4276) <= (layer0_outputs(3813)) or (layer0_outputs(4902));
    layer1_outputs(4277) <= '1';
    layer1_outputs(4278) <= layer0_outputs(791);
    layer1_outputs(4279) <= not(layer0_outputs(3956));
    layer1_outputs(4280) <= layer0_outputs(2917);
    layer1_outputs(4281) <= layer0_outputs(4943);
    layer1_outputs(4282) <= layer0_outputs(2710);
    layer1_outputs(4283) <= (layer0_outputs(4292)) and not (layer0_outputs(1697));
    layer1_outputs(4284) <= (layer0_outputs(6609)) and not (layer0_outputs(4648));
    layer1_outputs(4285) <= '0';
    layer1_outputs(4286) <= '0';
    layer1_outputs(4287) <= layer0_outputs(7191);
    layer1_outputs(4288) <= not(layer0_outputs(3027));
    layer1_outputs(4289) <= layer0_outputs(2918);
    layer1_outputs(4290) <= (layer0_outputs(7391)) and not (layer0_outputs(1628));
    layer1_outputs(4291) <= (layer0_outputs(7334)) and (layer0_outputs(5733));
    layer1_outputs(4292) <= not((layer0_outputs(109)) and (layer0_outputs(1615)));
    layer1_outputs(4293) <= not(layer0_outputs(6402)) or (layer0_outputs(502));
    layer1_outputs(4294) <= (layer0_outputs(6236)) xor (layer0_outputs(7102));
    layer1_outputs(4295) <= not(layer0_outputs(5981));
    layer1_outputs(4296) <= not(layer0_outputs(3448)) or (layer0_outputs(5053));
    layer1_outputs(4297) <= (layer0_outputs(4535)) and not (layer0_outputs(2038));
    layer1_outputs(4298) <= (layer0_outputs(7223)) and (layer0_outputs(4490));
    layer1_outputs(4299) <= not(layer0_outputs(972)) or (layer0_outputs(3763));
    layer1_outputs(4300) <= layer0_outputs(491);
    layer1_outputs(4301) <= '1';
    layer1_outputs(4302) <= layer0_outputs(4538);
    layer1_outputs(4303) <= not(layer0_outputs(1632)) or (layer0_outputs(6572));
    layer1_outputs(4304) <= layer0_outputs(2107);
    layer1_outputs(4305) <= '0';
    layer1_outputs(4306) <= layer0_outputs(6268);
    layer1_outputs(4307) <= not(layer0_outputs(2683)) or (layer0_outputs(4506));
    layer1_outputs(4308) <= (layer0_outputs(1274)) and (layer0_outputs(1752));
    layer1_outputs(4309) <= not((layer0_outputs(3087)) and (layer0_outputs(3645)));
    layer1_outputs(4310) <= (layer0_outputs(5520)) or (layer0_outputs(2910));
    layer1_outputs(4311) <= layer0_outputs(409);
    layer1_outputs(4312) <= (layer0_outputs(1847)) and not (layer0_outputs(6040));
    layer1_outputs(4313) <= layer0_outputs(3828);
    layer1_outputs(4314) <= (layer0_outputs(5760)) and (layer0_outputs(7213));
    layer1_outputs(4315) <= not(layer0_outputs(1362));
    layer1_outputs(4316) <= layer0_outputs(483);
    layer1_outputs(4317) <= layer0_outputs(2952);
    layer1_outputs(4318) <= not((layer0_outputs(1001)) and (layer0_outputs(3500)));
    layer1_outputs(4319) <= layer0_outputs(6421);
    layer1_outputs(4320) <= not((layer0_outputs(1242)) or (layer0_outputs(5187)));
    layer1_outputs(4321) <= not((layer0_outputs(4620)) or (layer0_outputs(7)));
    layer1_outputs(4322) <= (layer0_outputs(3929)) or (layer0_outputs(1168));
    layer1_outputs(4323) <= not((layer0_outputs(5694)) and (layer0_outputs(6108)));
    layer1_outputs(4324) <= not(layer0_outputs(3898));
    layer1_outputs(4325) <= not(layer0_outputs(1495));
    layer1_outputs(4326) <= not(layer0_outputs(1434)) or (layer0_outputs(5465));
    layer1_outputs(4327) <= not(layer0_outputs(459));
    layer1_outputs(4328) <= (layer0_outputs(3487)) or (layer0_outputs(52));
    layer1_outputs(4329) <= not(layer0_outputs(3743));
    layer1_outputs(4330) <= not(layer0_outputs(1600)) or (layer0_outputs(3245));
    layer1_outputs(4331) <= not(layer0_outputs(4660));
    layer1_outputs(4332) <= (layer0_outputs(781)) xor (layer0_outputs(6222));
    layer1_outputs(4333) <= not((layer0_outputs(2650)) and (layer0_outputs(2796)));
    layer1_outputs(4334) <= (layer0_outputs(7597)) and not (layer0_outputs(8));
    layer1_outputs(4335) <= not((layer0_outputs(3937)) xor (layer0_outputs(6408)));
    layer1_outputs(4336) <= not(layer0_outputs(54));
    layer1_outputs(4337) <= (layer0_outputs(4305)) and not (layer0_outputs(4486));
    layer1_outputs(4338) <= not(layer0_outputs(4280));
    layer1_outputs(4339) <= (layer0_outputs(4031)) xor (layer0_outputs(4002));
    layer1_outputs(4340) <= not(layer0_outputs(614)) or (layer0_outputs(11));
    layer1_outputs(4341) <= not((layer0_outputs(3265)) xor (layer0_outputs(2382)));
    layer1_outputs(4342) <= not((layer0_outputs(1082)) and (layer0_outputs(5424)));
    layer1_outputs(4343) <= (layer0_outputs(7211)) or (layer0_outputs(5205));
    layer1_outputs(4344) <= '1';
    layer1_outputs(4345) <= not(layer0_outputs(5557));
    layer1_outputs(4346) <= layer0_outputs(372);
    layer1_outputs(4347) <= not((layer0_outputs(4179)) and (layer0_outputs(4227)));
    layer1_outputs(4348) <= '1';
    layer1_outputs(4349) <= (layer0_outputs(1875)) or (layer0_outputs(5430));
    layer1_outputs(4350) <= not(layer0_outputs(887));
    layer1_outputs(4351) <= (layer0_outputs(7553)) and not (layer0_outputs(5677));
    layer1_outputs(4352) <= (layer0_outputs(3841)) or (layer0_outputs(1584));
    layer1_outputs(4353) <= not(layer0_outputs(4401));
    layer1_outputs(4354) <= not(layer0_outputs(4575)) or (layer0_outputs(2198));
    layer1_outputs(4355) <= '0';
    layer1_outputs(4356) <= not(layer0_outputs(3241));
    layer1_outputs(4357) <= not(layer0_outputs(3477));
    layer1_outputs(4358) <= layer0_outputs(7226);
    layer1_outputs(4359) <= not(layer0_outputs(6509)) or (layer0_outputs(3068));
    layer1_outputs(4360) <= layer0_outputs(6366);
    layer1_outputs(4361) <= layer0_outputs(3489);
    layer1_outputs(4362) <= not((layer0_outputs(5637)) or (layer0_outputs(4956)));
    layer1_outputs(4363) <= not(layer0_outputs(3638)) or (layer0_outputs(1297));
    layer1_outputs(4364) <= (layer0_outputs(4472)) and (layer0_outputs(636));
    layer1_outputs(4365) <= not(layer0_outputs(3834));
    layer1_outputs(4366) <= not(layer0_outputs(4463));
    layer1_outputs(4367) <= not((layer0_outputs(4703)) xor (layer0_outputs(332)));
    layer1_outputs(4368) <= layer0_outputs(6176);
    layer1_outputs(4369) <= not(layer0_outputs(5137));
    layer1_outputs(4370) <= not(layer0_outputs(677));
    layer1_outputs(4371) <= layer0_outputs(2889);
    layer1_outputs(4372) <= (layer0_outputs(713)) or (layer0_outputs(950));
    layer1_outputs(4373) <= not(layer0_outputs(4586)) or (layer0_outputs(4719));
    layer1_outputs(4374) <= (layer0_outputs(2920)) xor (layer0_outputs(4599));
    layer1_outputs(4375) <= not(layer0_outputs(1770)) or (layer0_outputs(308));
    layer1_outputs(4376) <= layer0_outputs(3543);
    layer1_outputs(4377) <= not(layer0_outputs(1334)) or (layer0_outputs(1073));
    layer1_outputs(4378) <= not(layer0_outputs(566)) or (layer0_outputs(1104));
    layer1_outputs(4379) <= not(layer0_outputs(1378)) or (layer0_outputs(6155));
    layer1_outputs(4380) <= not(layer0_outputs(1552)) or (layer0_outputs(3023));
    layer1_outputs(4381) <= '1';
    layer1_outputs(4382) <= '1';
    layer1_outputs(4383) <= '0';
    layer1_outputs(4384) <= not(layer0_outputs(3764)) or (layer0_outputs(6632));
    layer1_outputs(4385) <= not(layer0_outputs(5273));
    layer1_outputs(4386) <= not((layer0_outputs(3365)) or (layer0_outputs(2939)));
    layer1_outputs(4387) <= (layer0_outputs(5870)) xor (layer0_outputs(5031));
    layer1_outputs(4388) <= not(layer0_outputs(5210));
    layer1_outputs(4389) <= not(layer0_outputs(4941));
    layer1_outputs(4390) <= '0';
    layer1_outputs(4391) <= not(layer0_outputs(841)) or (layer0_outputs(1705));
    layer1_outputs(4392) <= '0';
    layer1_outputs(4393) <= not(layer0_outputs(785)) or (layer0_outputs(4123));
    layer1_outputs(4394) <= (layer0_outputs(4230)) and not (layer0_outputs(1236));
    layer1_outputs(4395) <= not(layer0_outputs(418));
    layer1_outputs(4396) <= '0';
    layer1_outputs(4397) <= not(layer0_outputs(5445));
    layer1_outputs(4398) <= not(layer0_outputs(4894));
    layer1_outputs(4399) <= layer0_outputs(3678);
    layer1_outputs(4400) <= layer0_outputs(2506);
    layer1_outputs(4401) <= layer0_outputs(7433);
    layer1_outputs(4402) <= not(layer0_outputs(6675)) or (layer0_outputs(1174));
    layer1_outputs(4403) <= (layer0_outputs(876)) and not (layer0_outputs(5711));
    layer1_outputs(4404) <= not(layer0_outputs(2046)) or (layer0_outputs(7248));
    layer1_outputs(4405) <= layer0_outputs(7424);
    layer1_outputs(4406) <= not(layer0_outputs(3138));
    layer1_outputs(4407) <= not(layer0_outputs(2313));
    layer1_outputs(4408) <= layer0_outputs(208);
    layer1_outputs(4409) <= '0';
    layer1_outputs(4410) <= (layer0_outputs(5103)) and not (layer0_outputs(725));
    layer1_outputs(4411) <= (layer0_outputs(5265)) and not (layer0_outputs(7107));
    layer1_outputs(4412) <= layer0_outputs(2529);
    layer1_outputs(4413) <= layer0_outputs(3392);
    layer1_outputs(4414) <= (layer0_outputs(7547)) or (layer0_outputs(1579));
    layer1_outputs(4415) <= '0';
    layer1_outputs(4416) <= (layer0_outputs(5321)) or (layer0_outputs(7578));
    layer1_outputs(4417) <= (layer0_outputs(947)) and not (layer0_outputs(5992));
    layer1_outputs(4418) <= layer0_outputs(740);
    layer1_outputs(4419) <= not(layer0_outputs(5033));
    layer1_outputs(4420) <= not((layer0_outputs(3306)) or (layer0_outputs(6670)));
    layer1_outputs(4421) <= layer0_outputs(782);
    layer1_outputs(4422) <= not(layer0_outputs(334));
    layer1_outputs(4423) <= (layer0_outputs(4823)) and (layer0_outputs(4804));
    layer1_outputs(4424) <= not(layer0_outputs(2957));
    layer1_outputs(4425) <= (layer0_outputs(5056)) and (layer0_outputs(7117));
    layer1_outputs(4426) <= not(layer0_outputs(5088));
    layer1_outputs(4427) <= (layer0_outputs(5914)) or (layer0_outputs(2727));
    layer1_outputs(4428) <= not(layer0_outputs(3015));
    layer1_outputs(4429) <= not(layer0_outputs(571)) or (layer0_outputs(7324));
    layer1_outputs(4430) <= '1';
    layer1_outputs(4431) <= not((layer0_outputs(4854)) and (layer0_outputs(3236)));
    layer1_outputs(4432) <= layer0_outputs(5951);
    layer1_outputs(4433) <= (layer0_outputs(1641)) and (layer0_outputs(5510));
    layer1_outputs(4434) <= not(layer0_outputs(6483));
    layer1_outputs(4435) <= not(layer0_outputs(4597));
    layer1_outputs(4436) <= (layer0_outputs(7585)) or (layer0_outputs(627));
    layer1_outputs(4437) <= layer0_outputs(909);
    layer1_outputs(4438) <= not(layer0_outputs(730));
    layer1_outputs(4439) <= not((layer0_outputs(2264)) or (layer0_outputs(272)));
    layer1_outputs(4440) <= (layer0_outputs(5119)) and not (layer0_outputs(3099));
    layer1_outputs(4441) <= not(layer0_outputs(757)) or (layer0_outputs(6530));
    layer1_outputs(4442) <= not(layer0_outputs(7287));
    layer1_outputs(4443) <= not(layer0_outputs(2736));
    layer1_outputs(4444) <= layer0_outputs(7120);
    layer1_outputs(4445) <= not(layer0_outputs(6735)) or (layer0_outputs(5561));
    layer1_outputs(4446) <= (layer0_outputs(145)) and not (layer0_outputs(2368));
    layer1_outputs(4447) <= layer0_outputs(7201);
    layer1_outputs(4448) <= not(layer0_outputs(7448));
    layer1_outputs(4449) <= layer0_outputs(3289);
    layer1_outputs(4450) <= (layer0_outputs(5408)) and not (layer0_outputs(3877));
    layer1_outputs(4451) <= '1';
    layer1_outputs(4452) <= (layer0_outputs(4758)) and not (layer0_outputs(107));
    layer1_outputs(4453) <= not((layer0_outputs(7233)) and (layer0_outputs(4786)));
    layer1_outputs(4454) <= (layer0_outputs(4914)) and (layer0_outputs(5002));
    layer1_outputs(4455) <= not(layer0_outputs(5940)) or (layer0_outputs(3706));
    layer1_outputs(4456) <= (layer0_outputs(2118)) and (layer0_outputs(7397));
    layer1_outputs(4457) <= not((layer0_outputs(4239)) or (layer0_outputs(5717)));
    layer1_outputs(4458) <= not((layer0_outputs(212)) and (layer0_outputs(326)));
    layer1_outputs(4459) <= not((layer0_outputs(7528)) and (layer0_outputs(158)));
    layer1_outputs(4460) <= layer0_outputs(2182);
    layer1_outputs(4461) <= not(layer0_outputs(940));
    layer1_outputs(4462) <= not(layer0_outputs(6878)) or (layer0_outputs(3682));
    layer1_outputs(4463) <= '1';
    layer1_outputs(4464) <= not(layer0_outputs(1569)) or (layer0_outputs(4646));
    layer1_outputs(4465) <= layer0_outputs(4152);
    layer1_outputs(4466) <= not((layer0_outputs(5691)) and (layer0_outputs(6223)));
    layer1_outputs(4467) <= (layer0_outputs(2042)) and not (layer0_outputs(679));
    layer1_outputs(4468) <= '1';
    layer1_outputs(4469) <= not(layer0_outputs(5901)) or (layer0_outputs(3902));
    layer1_outputs(4470) <= not(layer0_outputs(1591));
    layer1_outputs(4471) <= not((layer0_outputs(6283)) and (layer0_outputs(2058)));
    layer1_outputs(4472) <= not((layer0_outputs(5658)) and (layer0_outputs(606)));
    layer1_outputs(4473) <= layer0_outputs(4898);
    layer1_outputs(4474) <= not((layer0_outputs(5891)) xor (layer0_outputs(2331)));
    layer1_outputs(4475) <= (layer0_outputs(2642)) and not (layer0_outputs(7641));
    layer1_outputs(4476) <= '0';
    layer1_outputs(4477) <= '1';
    layer1_outputs(4478) <= not(layer0_outputs(2000)) or (layer0_outputs(2998));
    layer1_outputs(4479) <= not(layer0_outputs(3383));
    layer1_outputs(4480) <= (layer0_outputs(968)) and (layer0_outputs(6545));
    layer1_outputs(4481) <= not(layer0_outputs(4209));
    layer1_outputs(4482) <= (layer0_outputs(5610)) and not (layer0_outputs(2508));
    layer1_outputs(4483) <= layer0_outputs(4691);
    layer1_outputs(4484) <= (layer0_outputs(1528)) and not (layer0_outputs(118));
    layer1_outputs(4485) <= not(layer0_outputs(1520));
    layer1_outputs(4486) <= not(layer0_outputs(5743)) or (layer0_outputs(3906));
    layer1_outputs(4487) <= '1';
    layer1_outputs(4488) <= not(layer0_outputs(4489)) or (layer0_outputs(2044));
    layer1_outputs(4489) <= '0';
    layer1_outputs(4490) <= not(layer0_outputs(1194)) or (layer0_outputs(3377));
    layer1_outputs(4491) <= not(layer0_outputs(1508));
    layer1_outputs(4492) <= (layer0_outputs(3442)) and (layer0_outputs(2177));
    layer1_outputs(4493) <= layer0_outputs(215);
    layer1_outputs(4494) <= not(layer0_outputs(2242));
    layer1_outputs(4495) <= layer0_outputs(318);
    layer1_outputs(4496) <= '1';
    layer1_outputs(4497) <= not((layer0_outputs(2728)) and (layer0_outputs(7387)));
    layer1_outputs(4498) <= (layer0_outputs(4354)) or (layer0_outputs(3826));
    layer1_outputs(4499) <= layer0_outputs(67);
    layer1_outputs(4500) <= not((layer0_outputs(796)) or (layer0_outputs(3646)));
    layer1_outputs(4501) <= (layer0_outputs(2300)) xor (layer0_outputs(249));
    layer1_outputs(4502) <= (layer0_outputs(2364)) and not (layer0_outputs(5629));
    layer1_outputs(4503) <= not(layer0_outputs(2116)) or (layer0_outputs(1892));
    layer1_outputs(4504) <= layer0_outputs(804);
    layer1_outputs(4505) <= '1';
    layer1_outputs(4506) <= not(layer0_outputs(5664)) or (layer0_outputs(513));
    layer1_outputs(4507) <= (layer0_outputs(7079)) and not (layer0_outputs(7668));
    layer1_outputs(4508) <= layer0_outputs(2890);
    layer1_outputs(4509) <= layer0_outputs(1235);
    layer1_outputs(4510) <= (layer0_outputs(6741)) and (layer0_outputs(7454));
    layer1_outputs(4511) <= not(layer0_outputs(486));
    layer1_outputs(4512) <= not(layer0_outputs(2936)) or (layer0_outputs(3696));
    layer1_outputs(4513) <= not(layer0_outputs(5636)) or (layer0_outputs(5841));
    layer1_outputs(4514) <= not((layer0_outputs(6965)) and (layer0_outputs(3041)));
    layer1_outputs(4515) <= not((layer0_outputs(2914)) or (layer0_outputs(6868)));
    layer1_outputs(4516) <= not(layer0_outputs(2142));
    layer1_outputs(4517) <= '0';
    layer1_outputs(4518) <= (layer0_outputs(420)) and not (layer0_outputs(5692));
    layer1_outputs(4519) <= (layer0_outputs(5842)) xor (layer0_outputs(3063));
    layer1_outputs(4520) <= (layer0_outputs(3950)) and not (layer0_outputs(3619));
    layer1_outputs(4521) <= (layer0_outputs(2139)) and (layer0_outputs(3132));
    layer1_outputs(4522) <= (layer0_outputs(328)) xor (layer0_outputs(5324));
    layer1_outputs(4523) <= not(layer0_outputs(7215)) or (layer0_outputs(2584));
    layer1_outputs(4524) <= layer0_outputs(1103);
    layer1_outputs(4525) <= layer0_outputs(3309);
    layer1_outputs(4526) <= not((layer0_outputs(255)) or (layer0_outputs(4681)));
    layer1_outputs(4527) <= not(layer0_outputs(316)) or (layer0_outputs(6406));
    layer1_outputs(4528) <= (layer0_outputs(4519)) and not (layer0_outputs(7559));
    layer1_outputs(4529) <= layer0_outputs(716);
    layer1_outputs(4530) <= not(layer0_outputs(1471)) or (layer0_outputs(3732));
    layer1_outputs(4531) <= not(layer0_outputs(537)) or (layer0_outputs(6137));
    layer1_outputs(4532) <= (layer0_outputs(7263)) and (layer0_outputs(2948));
    layer1_outputs(4533) <= '1';
    layer1_outputs(4534) <= not(layer0_outputs(1940));
    layer1_outputs(4535) <= not((layer0_outputs(4884)) xor (layer0_outputs(2927)));
    layer1_outputs(4536) <= not(layer0_outputs(406)) or (layer0_outputs(1143));
    layer1_outputs(4537) <= not((layer0_outputs(3962)) and (layer0_outputs(4490)));
    layer1_outputs(4538) <= layer0_outputs(3861);
    layer1_outputs(4539) <= not(layer0_outputs(6296)) or (layer0_outputs(3524));
    layer1_outputs(4540) <= '1';
    layer1_outputs(4541) <= '0';
    layer1_outputs(4542) <= not(layer0_outputs(264));
    layer1_outputs(4543) <= layer0_outputs(3714);
    layer1_outputs(4544) <= (layer0_outputs(3147)) and not (layer0_outputs(5553));
    layer1_outputs(4545) <= (layer0_outputs(3596)) and not (layer0_outputs(1230));
    layer1_outputs(4546) <= not(layer0_outputs(7308)) or (layer0_outputs(4784));
    layer1_outputs(4547) <= (layer0_outputs(1184)) and not (layer0_outputs(6186));
    layer1_outputs(4548) <= (layer0_outputs(5111)) and (layer0_outputs(353));
    layer1_outputs(4549) <= layer0_outputs(4874);
    layer1_outputs(4550) <= (layer0_outputs(2824)) and not (layer0_outputs(1058));
    layer1_outputs(4551) <= (layer0_outputs(4343)) and not (layer0_outputs(3987));
    layer1_outputs(4552) <= '0';
    layer1_outputs(4553) <= not((layer0_outputs(6130)) or (layer0_outputs(6830)));
    layer1_outputs(4554) <= not((layer0_outputs(222)) and (layer0_outputs(3901)));
    layer1_outputs(4555) <= not(layer0_outputs(2305));
    layer1_outputs(4556) <= not((layer0_outputs(6692)) or (layer0_outputs(7139)));
    layer1_outputs(4557) <= (layer0_outputs(5737)) or (layer0_outputs(3842));
    layer1_outputs(4558) <= not(layer0_outputs(398)) or (layer0_outputs(1588));
    layer1_outputs(4559) <= not(layer0_outputs(6712));
    layer1_outputs(4560) <= not(layer0_outputs(4428)) or (layer0_outputs(6610));
    layer1_outputs(4561) <= not(layer0_outputs(4157)) or (layer0_outputs(1951));
    layer1_outputs(4562) <= not(layer0_outputs(3660)) or (layer0_outputs(1840));
    layer1_outputs(4563) <= not(layer0_outputs(7194));
    layer1_outputs(4564) <= (layer0_outputs(2926)) xor (layer0_outputs(5037));
    layer1_outputs(4565) <= not(layer0_outputs(4121));
    layer1_outputs(4566) <= (layer0_outputs(3492)) and not (layer0_outputs(1925));
    layer1_outputs(4567) <= (layer0_outputs(1379)) and not (layer0_outputs(6371));
    layer1_outputs(4568) <= (layer0_outputs(5000)) and not (layer0_outputs(1251));
    layer1_outputs(4569) <= not(layer0_outputs(3395));
    layer1_outputs(4570) <= (layer0_outputs(1078)) and (layer0_outputs(7227));
    layer1_outputs(4571) <= (layer0_outputs(9)) and not (layer0_outputs(7590));
    layer1_outputs(4572) <= not(layer0_outputs(4593));
    layer1_outputs(4573) <= (layer0_outputs(4809)) or (layer0_outputs(6005));
    layer1_outputs(4574) <= '0';
    layer1_outputs(4575) <= layer0_outputs(5839);
    layer1_outputs(4576) <= not(layer0_outputs(1504));
    layer1_outputs(4577) <= layer0_outputs(6425);
    layer1_outputs(4578) <= '1';
    layer1_outputs(4579) <= (layer0_outputs(1315)) and (layer0_outputs(665));
    layer1_outputs(4580) <= (layer0_outputs(5194)) xor (layer0_outputs(2839));
    layer1_outputs(4581) <= (layer0_outputs(449)) and not (layer0_outputs(4889));
    layer1_outputs(4582) <= '1';
    layer1_outputs(4583) <= not(layer0_outputs(5485));
    layer1_outputs(4584) <= layer0_outputs(5806);
    layer1_outputs(4585) <= not(layer0_outputs(5121));
    layer1_outputs(4586) <= not(layer0_outputs(5054)) or (layer0_outputs(1383));
    layer1_outputs(4587) <= layer0_outputs(7226);
    layer1_outputs(4588) <= (layer0_outputs(1886)) or (layer0_outputs(3097));
    layer1_outputs(4589) <= not(layer0_outputs(2591));
    layer1_outputs(4590) <= not((layer0_outputs(1466)) xor (layer0_outputs(6263)));
    layer1_outputs(4591) <= layer0_outputs(3177);
    layer1_outputs(4592) <= layer0_outputs(3202);
    layer1_outputs(4593) <= not(layer0_outputs(698)) or (layer0_outputs(3244));
    layer1_outputs(4594) <= '0';
    layer1_outputs(4595) <= '0';
    layer1_outputs(4596) <= (layer0_outputs(5939)) or (layer0_outputs(6174));
    layer1_outputs(4597) <= not(layer0_outputs(6334));
    layer1_outputs(4598) <= (layer0_outputs(3367)) or (layer0_outputs(7592));
    layer1_outputs(4599) <= (layer0_outputs(677)) and (layer0_outputs(5474));
    layer1_outputs(4600) <= not(layer0_outputs(6831)) or (layer0_outputs(6707));
    layer1_outputs(4601) <= layer0_outputs(6775);
    layer1_outputs(4602) <= '0';
    layer1_outputs(4603) <= not(layer0_outputs(1018));
    layer1_outputs(4604) <= layer0_outputs(5196);
    layer1_outputs(4605) <= not((layer0_outputs(1488)) and (layer0_outputs(6822)));
    layer1_outputs(4606) <= not(layer0_outputs(3772));
    layer1_outputs(4607) <= layer0_outputs(5125);
    layer1_outputs(4608) <= layer0_outputs(3871);
    layer1_outputs(4609) <= (layer0_outputs(2985)) and not (layer0_outputs(6248));
    layer1_outputs(4610) <= layer0_outputs(584);
    layer1_outputs(4611) <= (layer0_outputs(1940)) or (layer0_outputs(648));
    layer1_outputs(4612) <= not((layer0_outputs(4624)) and (layer0_outputs(213)));
    layer1_outputs(4613) <= not(layer0_outputs(6936)) or (layer0_outputs(7089));
    layer1_outputs(4614) <= not((layer0_outputs(5660)) and (layer0_outputs(3311)));
    layer1_outputs(4615) <= (layer0_outputs(7296)) and not (layer0_outputs(2454));
    layer1_outputs(4616) <= (layer0_outputs(507)) or (layer0_outputs(5887));
    layer1_outputs(4617) <= not((layer0_outputs(6232)) or (layer0_outputs(5257)));
    layer1_outputs(4618) <= (layer0_outputs(5899)) and not (layer0_outputs(2606));
    layer1_outputs(4619) <= (layer0_outputs(1269)) and not (layer0_outputs(4792));
    layer1_outputs(4620) <= not(layer0_outputs(7416));
    layer1_outputs(4621) <= not(layer0_outputs(2406));
    layer1_outputs(4622) <= layer0_outputs(4509);
    layer1_outputs(4623) <= layer0_outputs(1914);
    layer1_outputs(4624) <= (layer0_outputs(3958)) and not (layer0_outputs(1870));
    layer1_outputs(4625) <= (layer0_outputs(2001)) and (layer0_outputs(2862));
    layer1_outputs(4626) <= (layer0_outputs(6681)) xor (layer0_outputs(7532));
    layer1_outputs(4627) <= layer0_outputs(6912);
    layer1_outputs(4628) <= (layer0_outputs(3539)) or (layer0_outputs(3195));
    layer1_outputs(4629) <= not(layer0_outputs(4502));
    layer1_outputs(4630) <= not(layer0_outputs(2688)) or (layer0_outputs(4907));
    layer1_outputs(4631) <= (layer0_outputs(707)) and not (layer0_outputs(831));
    layer1_outputs(4632) <= not(layer0_outputs(463));
    layer1_outputs(4633) <= not(layer0_outputs(5581)) or (layer0_outputs(5549));
    layer1_outputs(4634) <= not(layer0_outputs(3800)) or (layer0_outputs(6095));
    layer1_outputs(4635) <= (layer0_outputs(7037)) xor (layer0_outputs(5603));
    layer1_outputs(4636) <= (layer0_outputs(161)) and not (layer0_outputs(5829));
    layer1_outputs(4637) <= (layer0_outputs(4479)) and not (layer0_outputs(6878));
    layer1_outputs(4638) <= layer0_outputs(7354);
    layer1_outputs(4639) <= '1';
    layer1_outputs(4640) <= (layer0_outputs(6621)) and not (layer0_outputs(6989));
    layer1_outputs(4641) <= layer0_outputs(2322);
    layer1_outputs(4642) <= '0';
    layer1_outputs(4643) <= not(layer0_outputs(3175)) or (layer0_outputs(6469));
    layer1_outputs(4644) <= '1';
    layer1_outputs(4645) <= not(layer0_outputs(1347));
    layer1_outputs(4646) <= (layer0_outputs(5315)) and not (layer0_outputs(426));
    layer1_outputs(4647) <= (layer0_outputs(6873)) and (layer0_outputs(632));
    layer1_outputs(4648) <= '0';
    layer1_outputs(4649) <= '1';
    layer1_outputs(4650) <= (layer0_outputs(1261)) and (layer0_outputs(5051));
    layer1_outputs(4651) <= (layer0_outputs(7081)) or (layer0_outputs(423));
    layer1_outputs(4652) <= layer0_outputs(5112);
    layer1_outputs(4653) <= (layer0_outputs(6450)) or (layer0_outputs(2929));
    layer1_outputs(4654) <= (layer0_outputs(787)) and not (layer0_outputs(4744));
    layer1_outputs(4655) <= layer0_outputs(806);
    layer1_outputs(4656) <= layer0_outputs(120);
    layer1_outputs(4657) <= (layer0_outputs(3998)) and not (layer0_outputs(7329));
    layer1_outputs(4658) <= not(layer0_outputs(2520)) or (layer0_outputs(3263));
    layer1_outputs(4659) <= (layer0_outputs(2350)) and not (layer0_outputs(2189));
    layer1_outputs(4660) <= not(layer0_outputs(668));
    layer1_outputs(4661) <= not(layer0_outputs(5130));
    layer1_outputs(4662) <= not(layer0_outputs(1880));
    layer1_outputs(4663) <= not(layer0_outputs(4668)) or (layer0_outputs(6340));
    layer1_outputs(4664) <= not(layer0_outputs(2253));
    layer1_outputs(4665) <= not((layer0_outputs(6697)) and (layer0_outputs(3773)));
    layer1_outputs(4666) <= not(layer0_outputs(7282));
    layer1_outputs(4667) <= (layer0_outputs(312)) and (layer0_outputs(5573));
    layer1_outputs(4668) <= '0';
    layer1_outputs(4669) <= (layer0_outputs(6455)) and (layer0_outputs(6771));
    layer1_outputs(4670) <= not(layer0_outputs(379)) or (layer0_outputs(2974));
    layer1_outputs(4671) <= layer0_outputs(1096);
    layer1_outputs(4672) <= layer0_outputs(2776);
    layer1_outputs(4673) <= not((layer0_outputs(5825)) or (layer0_outputs(2867)));
    layer1_outputs(4674) <= not((layer0_outputs(5794)) or (layer0_outputs(7327)));
    layer1_outputs(4675) <= layer0_outputs(2426);
    layer1_outputs(4676) <= (layer0_outputs(2336)) or (layer0_outputs(3631));
    layer1_outputs(4677) <= not(layer0_outputs(2154)) or (layer0_outputs(4234));
    layer1_outputs(4678) <= (layer0_outputs(4026)) or (layer0_outputs(1681));
    layer1_outputs(4679) <= layer0_outputs(3999);
    layer1_outputs(4680) <= (layer0_outputs(7351)) and not (layer0_outputs(1147));
    layer1_outputs(4681) <= not(layer0_outputs(3742));
    layer1_outputs(4682) <= not(layer0_outputs(6506));
    layer1_outputs(4683) <= not(layer0_outputs(4288));
    layer1_outputs(4684) <= layer0_outputs(1845);
    layer1_outputs(4685) <= layer0_outputs(4187);
    layer1_outputs(4686) <= not(layer0_outputs(6925));
    layer1_outputs(4687) <= layer0_outputs(319);
    layer1_outputs(4688) <= not(layer0_outputs(2231));
    layer1_outputs(4689) <= layer0_outputs(6972);
    layer1_outputs(4690) <= (layer0_outputs(1567)) and not (layer0_outputs(114));
    layer1_outputs(4691) <= layer0_outputs(4423);
    layer1_outputs(4692) <= layer0_outputs(6850);
    layer1_outputs(4693) <= not(layer0_outputs(1019)) or (layer0_outputs(643));
    layer1_outputs(4694) <= not(layer0_outputs(1557));
    layer1_outputs(4695) <= not(layer0_outputs(177));
    layer1_outputs(4696) <= not((layer0_outputs(3298)) or (layer0_outputs(4026)));
    layer1_outputs(4697) <= not(layer0_outputs(5289));
    layer1_outputs(4698) <= not(layer0_outputs(6551)) or (layer0_outputs(6076));
    layer1_outputs(4699) <= not(layer0_outputs(5943)) or (layer0_outputs(1497));
    layer1_outputs(4700) <= not(layer0_outputs(1297));
    layer1_outputs(4701) <= (layer0_outputs(6351)) and not (layer0_outputs(3001));
    layer1_outputs(4702) <= (layer0_outputs(6555)) and not (layer0_outputs(2850));
    layer1_outputs(4703) <= not(layer0_outputs(1407)) or (layer0_outputs(6649));
    layer1_outputs(4704) <= not(layer0_outputs(6428));
    layer1_outputs(4705) <= (layer0_outputs(4920)) or (layer0_outputs(3193));
    layer1_outputs(4706) <= (layer0_outputs(5077)) and not (layer0_outputs(2739));
    layer1_outputs(4707) <= layer0_outputs(2951);
    layer1_outputs(4708) <= layer0_outputs(490);
    layer1_outputs(4709) <= not(layer0_outputs(3058)) or (layer0_outputs(7120));
    layer1_outputs(4710) <= not(layer0_outputs(3272));
    layer1_outputs(4711) <= layer0_outputs(5156);
    layer1_outputs(4712) <= not((layer0_outputs(6239)) xor (layer0_outputs(3522)));
    layer1_outputs(4713) <= layer0_outputs(794);
    layer1_outputs(4714) <= not(layer0_outputs(5477)) or (layer0_outputs(7517));
    layer1_outputs(4715) <= not(layer0_outputs(792)) or (layer0_outputs(6803));
    layer1_outputs(4716) <= not(layer0_outputs(4938));
    layer1_outputs(4717) <= not(layer0_outputs(4612));
    layer1_outputs(4718) <= not(layer0_outputs(1006));
    layer1_outputs(4719) <= not(layer0_outputs(5141));
    layer1_outputs(4720) <= not(layer0_outputs(7471)) or (layer0_outputs(7222));
    layer1_outputs(4721) <= not(layer0_outputs(3213));
    layer1_outputs(4722) <= layer0_outputs(6378);
    layer1_outputs(4723) <= not((layer0_outputs(6151)) or (layer0_outputs(1580)));
    layer1_outputs(4724) <= not(layer0_outputs(7441)) or (layer0_outputs(6333));
    layer1_outputs(4725) <= not(layer0_outputs(7096));
    layer1_outputs(4726) <= not((layer0_outputs(934)) and (layer0_outputs(5910)));
    layer1_outputs(4727) <= not(layer0_outputs(7254));
    layer1_outputs(4728) <= layer0_outputs(3794);
    layer1_outputs(4729) <= layer0_outputs(1071);
    layer1_outputs(4730) <= (layer0_outputs(7422)) or (layer0_outputs(7159));
    layer1_outputs(4731) <= (layer0_outputs(7074)) and not (layer0_outputs(1536));
    layer1_outputs(4732) <= layer0_outputs(927);
    layer1_outputs(4733) <= not(layer0_outputs(5334));
    layer1_outputs(4734) <= (layer0_outputs(284)) xor (layer0_outputs(576));
    layer1_outputs(4735) <= not((layer0_outputs(1067)) or (layer0_outputs(7578)));
    layer1_outputs(4736) <= not(layer0_outputs(1852)) or (layer0_outputs(4578));
    layer1_outputs(4737) <= layer0_outputs(225);
    layer1_outputs(4738) <= not((layer0_outputs(6971)) and (layer0_outputs(2176)));
    layer1_outputs(4739) <= not(layer0_outputs(4231));
    layer1_outputs(4740) <= (layer0_outputs(7453)) and (layer0_outputs(6867));
    layer1_outputs(4741) <= (layer0_outputs(5552)) and not (layer0_outputs(628));
    layer1_outputs(4742) <= layer0_outputs(1584);
    layer1_outputs(4743) <= not((layer0_outputs(1164)) or (layer0_outputs(996)));
    layer1_outputs(4744) <= not((layer0_outputs(787)) or (layer0_outputs(5360)));
    layer1_outputs(4745) <= (layer0_outputs(5930)) xor (layer0_outputs(6012));
    layer1_outputs(4746) <= (layer0_outputs(1528)) or (layer0_outputs(1404));
    layer1_outputs(4747) <= layer0_outputs(4226);
    layer1_outputs(4748) <= not(layer0_outputs(1141)) or (layer0_outputs(2719));
    layer1_outputs(4749) <= (layer0_outputs(2768)) and not (layer0_outputs(1450));
    layer1_outputs(4750) <= not(layer0_outputs(7010));
    layer1_outputs(4751) <= not((layer0_outputs(3973)) and (layer0_outputs(5042)));
    layer1_outputs(4752) <= not(layer0_outputs(5967)) or (layer0_outputs(1076));
    layer1_outputs(4753) <= layer0_outputs(644);
    layer1_outputs(4754) <= not(layer0_outputs(849)) or (layer0_outputs(5885));
    layer1_outputs(4755) <= not(layer0_outputs(682)) or (layer0_outputs(1711));
    layer1_outputs(4756) <= not((layer0_outputs(4436)) or (layer0_outputs(1144)));
    layer1_outputs(4757) <= '1';
    layer1_outputs(4758) <= (layer0_outputs(2937)) and (layer0_outputs(4341));
    layer1_outputs(4759) <= not((layer0_outputs(1834)) and (layer0_outputs(6471)));
    layer1_outputs(4760) <= not(layer0_outputs(5942)) or (layer0_outputs(109));
    layer1_outputs(4761) <= (layer0_outputs(7083)) and not (layer0_outputs(5128));
    layer1_outputs(4762) <= not(layer0_outputs(2034));
    layer1_outputs(4763) <= layer0_outputs(6286);
    layer1_outputs(4764) <= not(layer0_outputs(970));
    layer1_outputs(4765) <= not(layer0_outputs(6727)) or (layer0_outputs(3769));
    layer1_outputs(4766) <= (layer0_outputs(7221)) and not (layer0_outputs(4697));
    layer1_outputs(4767) <= not(layer0_outputs(2882)) or (layer0_outputs(1470));
    layer1_outputs(4768) <= (layer0_outputs(3749)) and not (layer0_outputs(5709));
    layer1_outputs(4769) <= not(layer0_outputs(1090)) or (layer0_outputs(2041));
    layer1_outputs(4770) <= layer0_outputs(1099);
    layer1_outputs(4771) <= layer0_outputs(6700);
    layer1_outputs(4772) <= not((layer0_outputs(7233)) and (layer0_outputs(1855)));
    layer1_outputs(4773) <= '0';
    layer1_outputs(4774) <= (layer0_outputs(6261)) and not (layer0_outputs(4340));
    layer1_outputs(4775) <= not(layer0_outputs(936)) or (layer0_outputs(7244));
    layer1_outputs(4776) <= not(layer0_outputs(6886));
    layer1_outputs(4777) <= not(layer0_outputs(3862)) or (layer0_outputs(5612));
    layer1_outputs(4778) <= not(layer0_outputs(593));
    layer1_outputs(4779) <= layer0_outputs(1809);
    layer1_outputs(4780) <= (layer0_outputs(5877)) and (layer0_outputs(3869));
    layer1_outputs(4781) <= not((layer0_outputs(5375)) and (layer0_outputs(705)));
    layer1_outputs(4782) <= layer0_outputs(5462);
    layer1_outputs(4783) <= not((layer0_outputs(4108)) or (layer0_outputs(5827)));
    layer1_outputs(4784) <= (layer0_outputs(516)) and (layer0_outputs(4507));
    layer1_outputs(4785) <= not(layer0_outputs(6264));
    layer1_outputs(4786) <= '1';
    layer1_outputs(4787) <= not(layer0_outputs(6312));
    layer1_outputs(4788) <= not(layer0_outputs(3284));
    layer1_outputs(4789) <= (layer0_outputs(5038)) and not (layer0_outputs(4466));
    layer1_outputs(4790) <= not(layer0_outputs(3484));
    layer1_outputs(4791) <= not(layer0_outputs(385));
    layer1_outputs(4792) <= (layer0_outputs(4569)) and (layer0_outputs(896));
    layer1_outputs(4793) <= not(layer0_outputs(4300));
    layer1_outputs(4794) <= layer0_outputs(741);
    layer1_outputs(4795) <= not((layer0_outputs(6914)) and (layer0_outputs(6891)));
    layer1_outputs(4796) <= not((layer0_outputs(4799)) or (layer0_outputs(6446)));
    layer1_outputs(4797) <= not(layer0_outputs(797)) or (layer0_outputs(6184));
    layer1_outputs(4798) <= not(layer0_outputs(719)) or (layer0_outputs(1551));
    layer1_outputs(4799) <= layer0_outputs(3474);
    layer1_outputs(4800) <= not(layer0_outputs(6279)) or (layer0_outputs(2963));
    layer1_outputs(4801) <= not(layer0_outputs(2910));
    layer1_outputs(4802) <= (layer0_outputs(4983)) and not (layer0_outputs(7154));
    layer1_outputs(4803) <= (layer0_outputs(6529)) or (layer0_outputs(5927));
    layer1_outputs(4804) <= not(layer0_outputs(1303)) or (layer0_outputs(5853));
    layer1_outputs(4805) <= not(layer0_outputs(569));
    layer1_outputs(4806) <= layer0_outputs(1931);
    layer1_outputs(4807) <= (layer0_outputs(1798)) or (layer0_outputs(2005));
    layer1_outputs(4808) <= layer0_outputs(92);
    layer1_outputs(4809) <= not((layer0_outputs(2216)) xor (layer0_outputs(2683)));
    layer1_outputs(4810) <= layer0_outputs(4040);
    layer1_outputs(4811) <= not(layer0_outputs(7372)) or (layer0_outputs(7381));
    layer1_outputs(4812) <= not(layer0_outputs(3308));
    layer1_outputs(4813) <= layer0_outputs(7091);
    layer1_outputs(4814) <= '0';
    layer1_outputs(4815) <= not((layer0_outputs(1643)) xor (layer0_outputs(4798)));
    layer1_outputs(4816) <= not(layer0_outputs(1467));
    layer1_outputs(4817) <= layer0_outputs(5522);
    layer1_outputs(4818) <= layer0_outputs(1922);
    layer1_outputs(4819) <= not((layer0_outputs(468)) or (layer0_outputs(1219)));
    layer1_outputs(4820) <= not(layer0_outputs(557));
    layer1_outputs(4821) <= (layer0_outputs(2175)) and not (layer0_outputs(2074));
    layer1_outputs(4822) <= layer0_outputs(6500);
    layer1_outputs(4823) <= (layer0_outputs(364)) and (layer0_outputs(5357));
    layer1_outputs(4824) <= not(layer0_outputs(7584)) or (layer0_outputs(2485));
    layer1_outputs(4825) <= layer0_outputs(6086);
    layer1_outputs(4826) <= (layer0_outputs(2941)) and not (layer0_outputs(5345));
    layer1_outputs(4827) <= '1';
    layer1_outputs(4828) <= (layer0_outputs(295)) and not (layer0_outputs(5772));
    layer1_outputs(4829) <= (layer0_outputs(4048)) and (layer0_outputs(4187));
    layer1_outputs(4830) <= layer0_outputs(6756);
    layer1_outputs(4831) <= not(layer0_outputs(5811));
    layer1_outputs(4832) <= '1';
    layer1_outputs(4833) <= not(layer0_outputs(6068));
    layer1_outputs(4834) <= layer0_outputs(1233);
    layer1_outputs(4835) <= not((layer0_outputs(2268)) and (layer0_outputs(6523)));
    layer1_outputs(4836) <= '1';
    layer1_outputs(4837) <= (layer0_outputs(2197)) and (layer0_outputs(4268));
    layer1_outputs(4838) <= (layer0_outputs(925)) and not (layer0_outputs(3136));
    layer1_outputs(4839) <= (layer0_outputs(5562)) and not (layer0_outputs(4969));
    layer1_outputs(4840) <= layer0_outputs(1503);
    layer1_outputs(4841) <= layer0_outputs(4793);
    layer1_outputs(4842) <= '0';
    layer1_outputs(4843) <= not(layer0_outputs(586));
    layer1_outputs(4844) <= (layer0_outputs(3966)) and not (layer0_outputs(2609));
    layer1_outputs(4845) <= (layer0_outputs(5723)) and not (layer0_outputs(2607));
    layer1_outputs(4846) <= layer0_outputs(7242);
    layer1_outputs(4847) <= '1';
    layer1_outputs(4848) <= not((layer0_outputs(2059)) and (layer0_outputs(3145)));
    layer1_outputs(4849) <= '1';
    layer1_outputs(4850) <= (layer0_outputs(1357)) and not (layer0_outputs(773));
    layer1_outputs(4851) <= (layer0_outputs(4550)) and not (layer0_outputs(2455));
    layer1_outputs(4852) <= (layer0_outputs(6651)) and (layer0_outputs(3032));
    layer1_outputs(4853) <= not(layer0_outputs(3694)) or (layer0_outputs(3497));
    layer1_outputs(4854) <= '1';
    layer1_outputs(4855) <= (layer0_outputs(3946)) and (layer0_outputs(4097));
    layer1_outputs(4856) <= (layer0_outputs(3523)) and not (layer0_outputs(3674));
    layer1_outputs(4857) <= '0';
    layer1_outputs(4858) <= not(layer0_outputs(4508));
    layer1_outputs(4859) <= (layer0_outputs(6242)) and not (layer0_outputs(4945));
    layer1_outputs(4860) <= not((layer0_outputs(3970)) and (layer0_outputs(3708)));
    layer1_outputs(4861) <= not(layer0_outputs(2897));
    layer1_outputs(4862) <= not(layer0_outputs(7562));
    layer1_outputs(4863) <= not(layer0_outputs(3251)) or (layer0_outputs(1176));
    layer1_outputs(4864) <= '0';
    layer1_outputs(4865) <= not((layer0_outputs(4663)) xor (layer0_outputs(3228)));
    layer1_outputs(4866) <= layer0_outputs(5678);
    layer1_outputs(4867) <= not(layer0_outputs(4612));
    layer1_outputs(4868) <= '1';
    layer1_outputs(4869) <= (layer0_outputs(2496)) and (layer0_outputs(7071));
    layer1_outputs(4870) <= '1';
    layer1_outputs(4871) <= (layer0_outputs(1684)) or (layer0_outputs(889));
    layer1_outputs(4872) <= not(layer0_outputs(2611));
    layer1_outputs(4873) <= not(layer0_outputs(6208)) or (layer0_outputs(5314));
    layer1_outputs(4874) <= (layer0_outputs(2273)) and (layer0_outputs(3134));
    layer1_outputs(4875) <= layer0_outputs(6862);
    layer1_outputs(4876) <= layer0_outputs(5188);
    layer1_outputs(4877) <= layer0_outputs(2247);
    layer1_outputs(4878) <= not(layer0_outputs(2367));
    layer1_outputs(4879) <= (layer0_outputs(231)) and not (layer0_outputs(5750));
    layer1_outputs(4880) <= not(layer0_outputs(2043));
    layer1_outputs(4881) <= not(layer0_outputs(2605));
    layer1_outputs(4882) <= '1';
    layer1_outputs(4883) <= layer0_outputs(4945);
    layer1_outputs(4884) <= not(layer0_outputs(4215)) or (layer0_outputs(6930));
    layer1_outputs(4885) <= not(layer0_outputs(3967)) or (layer0_outputs(7350));
    layer1_outputs(4886) <= (layer0_outputs(5975)) and not (layer0_outputs(7665));
    layer1_outputs(4887) <= not(layer0_outputs(3526));
    layer1_outputs(4888) <= (layer0_outputs(4319)) and not (layer0_outputs(5736));
    layer1_outputs(4889) <= not((layer0_outputs(3936)) or (layer0_outputs(4516)));
    layer1_outputs(4890) <= not((layer0_outputs(4057)) and (layer0_outputs(475)));
    layer1_outputs(4891) <= not(layer0_outputs(6242));
    layer1_outputs(4892) <= layer0_outputs(1674);
    layer1_outputs(4893) <= not(layer0_outputs(3414));
    layer1_outputs(4894) <= not(layer0_outputs(7340));
    layer1_outputs(4895) <= '1';
    layer1_outputs(4896) <= not((layer0_outputs(2465)) and (layer0_outputs(2871)));
    layer1_outputs(4897) <= not((layer0_outputs(4321)) and (layer0_outputs(1517)));
    layer1_outputs(4898) <= not(layer0_outputs(3860));
    layer1_outputs(4899) <= not(layer0_outputs(6105));
    layer1_outputs(4900) <= layer0_outputs(2818);
    layer1_outputs(4901) <= not((layer0_outputs(522)) or (layer0_outputs(2919)));
    layer1_outputs(4902) <= layer0_outputs(4206);
    layer1_outputs(4903) <= not((layer0_outputs(6944)) and (layer0_outputs(3029)));
    layer1_outputs(4904) <= not(layer0_outputs(5930));
    layer1_outputs(4905) <= '1';
    layer1_outputs(4906) <= not(layer0_outputs(4942));
    layer1_outputs(4907) <= (layer0_outputs(4675)) and (layer0_outputs(664));
    layer1_outputs(4908) <= not((layer0_outputs(3731)) or (layer0_outputs(4661)));
    layer1_outputs(4909) <= not(layer0_outputs(2830));
    layer1_outputs(4910) <= (layer0_outputs(6874)) and not (layer0_outputs(1856));
    layer1_outputs(4911) <= not((layer0_outputs(3799)) or (layer0_outputs(7016)));
    layer1_outputs(4912) <= layer0_outputs(6356);
    layer1_outputs(4913) <= layer0_outputs(4176);
    layer1_outputs(4914) <= layer0_outputs(4438);
    layer1_outputs(4915) <= '1';
    layer1_outputs(4916) <= '0';
    layer1_outputs(4917) <= (layer0_outputs(2346)) xor (layer0_outputs(3171));
    layer1_outputs(4918) <= not((layer0_outputs(6507)) and (layer0_outputs(3625)));
    layer1_outputs(4919) <= (layer0_outputs(3584)) and (layer0_outputs(815));
    layer1_outputs(4920) <= (layer0_outputs(2815)) and not (layer0_outputs(373));
    layer1_outputs(4921) <= (layer0_outputs(1548)) and not (layer0_outputs(6062));
    layer1_outputs(4922) <= (layer0_outputs(6457)) and not (layer0_outputs(4086));
    layer1_outputs(4923) <= (layer0_outputs(5604)) and not (layer0_outputs(5492));
    layer1_outputs(4924) <= not(layer0_outputs(2451));
    layer1_outputs(4925) <= (layer0_outputs(525)) and not (layer0_outputs(2872));
    layer1_outputs(4926) <= (layer0_outputs(2190)) and not (layer0_outputs(1147));
    layer1_outputs(4927) <= layer0_outputs(2092);
    layer1_outputs(4928) <= not((layer0_outputs(2588)) or (layer0_outputs(7626)));
    layer1_outputs(4929) <= layer0_outputs(6751);
    layer1_outputs(4930) <= (layer0_outputs(4619)) and not (layer0_outputs(153));
    layer1_outputs(4931) <= layer0_outputs(7007);
    layer1_outputs(4932) <= not(layer0_outputs(5388));
    layer1_outputs(4933) <= not(layer0_outputs(1680));
    layer1_outputs(4934) <= '0';
    layer1_outputs(4935) <= (layer0_outputs(5729)) and not (layer0_outputs(7091));
    layer1_outputs(4936) <= (layer0_outputs(321)) or (layer0_outputs(2571));
    layer1_outputs(4937) <= layer0_outputs(2013);
    layer1_outputs(4938) <= (layer0_outputs(6111)) or (layer0_outputs(599));
    layer1_outputs(4939) <= '1';
    layer1_outputs(4940) <= (layer0_outputs(4692)) and not (layer0_outputs(5320));
    layer1_outputs(4941) <= (layer0_outputs(6061)) and (layer0_outputs(4268));
    layer1_outputs(4942) <= layer0_outputs(1784);
    layer1_outputs(4943) <= (layer0_outputs(5347)) or (layer0_outputs(5384));
    layer1_outputs(4944) <= layer0_outputs(4881);
    layer1_outputs(4945) <= '1';
    layer1_outputs(4946) <= (layer0_outputs(1864)) or (layer0_outputs(6071));
    layer1_outputs(4947) <= (layer0_outputs(4126)) and not (layer0_outputs(6198));
    layer1_outputs(4948) <= (layer0_outputs(7344)) and not (layer0_outputs(5579));
    layer1_outputs(4949) <= not((layer0_outputs(7412)) or (layer0_outputs(3238)));
    layer1_outputs(4950) <= (layer0_outputs(5718)) or (layer0_outputs(199));
    layer1_outputs(4951) <= layer0_outputs(7672);
    layer1_outputs(4952) <= layer0_outputs(809);
    layer1_outputs(4953) <= (layer0_outputs(2334)) and (layer0_outputs(6879));
    layer1_outputs(4954) <= not(layer0_outputs(3125));
    layer1_outputs(4955) <= layer0_outputs(3154);
    layer1_outputs(4956) <= not(layer0_outputs(5454));
    layer1_outputs(4957) <= (layer0_outputs(3497)) and (layer0_outputs(5618));
    layer1_outputs(4958) <= (layer0_outputs(4166)) and not (layer0_outputs(7088));
    layer1_outputs(4959) <= not((layer0_outputs(1941)) or (layer0_outputs(2398)));
    layer1_outputs(4960) <= not((layer0_outputs(4890)) or (layer0_outputs(1328)));
    layer1_outputs(4961) <= not(layer0_outputs(6582)) or (layer0_outputs(1887));
    layer1_outputs(4962) <= not(layer0_outputs(6023));
    layer1_outputs(4963) <= not((layer0_outputs(7504)) and (layer0_outputs(3061)));
    layer1_outputs(4964) <= layer0_outputs(636);
    layer1_outputs(4965) <= (layer0_outputs(3494)) and not (layer0_outputs(4575));
    layer1_outputs(4966) <= not(layer0_outputs(1979));
    layer1_outputs(4967) <= layer0_outputs(2145);
    layer1_outputs(4968) <= layer0_outputs(5704);
    layer1_outputs(4969) <= layer0_outputs(3490);
    layer1_outputs(4970) <= not((layer0_outputs(2323)) and (layer0_outputs(897)));
    layer1_outputs(4971) <= not(layer0_outputs(5032));
    layer1_outputs(4972) <= not((layer0_outputs(2249)) and (layer0_outputs(5968)));
    layer1_outputs(4973) <= not((layer0_outputs(7509)) and (layer0_outputs(1213)));
    layer1_outputs(4974) <= (layer0_outputs(5251)) or (layer0_outputs(5015));
    layer1_outputs(4975) <= (layer0_outputs(3361)) or (layer0_outputs(247));
    layer1_outputs(4976) <= not(layer0_outputs(4864));
    layer1_outputs(4977) <= (layer0_outputs(1068)) or (layer0_outputs(2903));
    layer1_outputs(4978) <= '1';
    layer1_outputs(4979) <= not(layer0_outputs(7482));
    layer1_outputs(4980) <= (layer0_outputs(4255)) and not (layer0_outputs(6326));
    layer1_outputs(4981) <= not(layer0_outputs(1556)) or (layer0_outputs(2483));
    layer1_outputs(4982) <= not(layer0_outputs(1910));
    layer1_outputs(4983) <= (layer0_outputs(2821)) and not (layer0_outputs(3785));
    layer1_outputs(4984) <= (layer0_outputs(4864)) and not (layer0_outputs(7168));
    layer1_outputs(4985) <= not((layer0_outputs(6436)) or (layer0_outputs(4901)));
    layer1_outputs(4986) <= not((layer0_outputs(444)) xor (layer0_outputs(4318)));
    layer1_outputs(4987) <= layer0_outputs(1256);
    layer1_outputs(4988) <= (layer0_outputs(358)) or (layer0_outputs(6776));
    layer1_outputs(4989) <= layer0_outputs(5249);
    layer1_outputs(4990) <= not(layer0_outputs(771)) or (layer0_outputs(6162));
    layer1_outputs(4991) <= (layer0_outputs(3256)) or (layer0_outputs(6046));
    layer1_outputs(4992) <= not(layer0_outputs(6910));
    layer1_outputs(4993) <= (layer0_outputs(3366)) and not (layer0_outputs(4995));
    layer1_outputs(4994) <= (layer0_outputs(4699)) and not (layer0_outputs(5019));
    layer1_outputs(4995) <= not(layer0_outputs(6348));
    layer1_outputs(4996) <= not(layer0_outputs(4695)) or (layer0_outputs(2645));
    layer1_outputs(4997) <= not((layer0_outputs(4208)) xor (layer0_outputs(266)));
    layer1_outputs(4998) <= layer0_outputs(5998);
    layer1_outputs(4999) <= (layer0_outputs(4431)) or (layer0_outputs(868));
    layer1_outputs(5000) <= not((layer0_outputs(6567)) or (layer0_outputs(668)));
    layer1_outputs(5001) <= not((layer0_outputs(6694)) and (layer0_outputs(91)));
    layer1_outputs(5002) <= not(layer0_outputs(7611)) or (layer0_outputs(5952));
    layer1_outputs(5003) <= layer0_outputs(3386);
    layer1_outputs(5004) <= not((layer0_outputs(2684)) xor (layer0_outputs(7073)));
    layer1_outputs(5005) <= (layer0_outputs(4082)) xor (layer0_outputs(139));
    layer1_outputs(5006) <= (layer0_outputs(3243)) and not (layer0_outputs(1656));
    layer1_outputs(5007) <= not(layer0_outputs(5275));
    layer1_outputs(5008) <= not((layer0_outputs(5940)) and (layer0_outputs(2635)));
    layer1_outputs(5009) <= not(layer0_outputs(4743));
    layer1_outputs(5010) <= layer0_outputs(3364);
    layer1_outputs(5011) <= (layer0_outputs(7027)) or (layer0_outputs(3327));
    layer1_outputs(5012) <= not((layer0_outputs(5527)) or (layer0_outputs(7083)));
    layer1_outputs(5013) <= not(layer0_outputs(695)) or (layer0_outputs(1718));
    layer1_outputs(5014) <= (layer0_outputs(3866)) and (layer0_outputs(3513));
    layer1_outputs(5015) <= not((layer0_outputs(1593)) or (layer0_outputs(7656)));
    layer1_outputs(5016) <= (layer0_outputs(2659)) and not (layer0_outputs(7066));
    layer1_outputs(5017) <= '0';
    layer1_outputs(5018) <= layer0_outputs(5069);
    layer1_outputs(5019) <= layer0_outputs(517);
    layer1_outputs(5020) <= '0';
    layer1_outputs(5021) <= not(layer0_outputs(4651)) or (layer0_outputs(318));
    layer1_outputs(5022) <= (layer0_outputs(2988)) and (layer0_outputs(4843));
    layer1_outputs(5023) <= '1';
    layer1_outputs(5024) <= not(layer0_outputs(2925)) or (layer0_outputs(5862));
    layer1_outputs(5025) <= (layer0_outputs(5735)) and (layer0_outputs(1963));
    layer1_outputs(5026) <= '1';
    layer1_outputs(5027) <= layer0_outputs(6731);
    layer1_outputs(5028) <= (layer0_outputs(2570)) and (layer0_outputs(2567));
    layer1_outputs(5029) <= (layer0_outputs(5291)) or (layer0_outputs(433));
    layer1_outputs(5030) <= (layer0_outputs(2542)) and not (layer0_outputs(4810));
    layer1_outputs(5031) <= not((layer0_outputs(7657)) and (layer0_outputs(7093)));
    layer1_outputs(5032) <= not(layer0_outputs(3327));
    layer1_outputs(5033) <= not(layer0_outputs(2225));
    layer1_outputs(5034) <= not(layer0_outputs(1554));
    layer1_outputs(5035) <= layer0_outputs(123);
    layer1_outputs(5036) <= (layer0_outputs(61)) or (layer0_outputs(5753));
    layer1_outputs(5037) <= (layer0_outputs(2090)) and not (layer0_outputs(5750));
    layer1_outputs(5038) <= (layer0_outputs(5227)) or (layer0_outputs(2866));
    layer1_outputs(5039) <= '1';
    layer1_outputs(5040) <= (layer0_outputs(4667)) and not (layer0_outputs(243));
    layer1_outputs(5041) <= (layer0_outputs(6024)) or (layer0_outputs(4450));
    layer1_outputs(5042) <= (layer0_outputs(3047)) and not (layer0_outputs(4876));
    layer1_outputs(5043) <= '1';
    layer1_outputs(5044) <= layer0_outputs(3173);
    layer1_outputs(5045) <= not((layer0_outputs(1390)) and (layer0_outputs(7466)));
    layer1_outputs(5046) <= layer0_outputs(1954);
    layer1_outputs(5047) <= layer0_outputs(2095);
    layer1_outputs(5048) <= not((layer0_outputs(2900)) xor (layer0_outputs(4441)));
    layer1_outputs(5049) <= not(layer0_outputs(6082)) or (layer0_outputs(7342));
    layer1_outputs(5050) <= (layer0_outputs(2702)) xor (layer0_outputs(2812));
    layer1_outputs(5051) <= not((layer0_outputs(5688)) or (layer0_outputs(7314)));
    layer1_outputs(5052) <= not(layer0_outputs(1163)) or (layer0_outputs(6568));
    layer1_outputs(5053) <= not((layer0_outputs(5074)) or (layer0_outputs(446)));
    layer1_outputs(5054) <= layer0_outputs(4099);
    layer1_outputs(5055) <= not((layer0_outputs(4135)) or (layer0_outputs(1902)));
    layer1_outputs(5056) <= not(layer0_outputs(30)) or (layer0_outputs(1749));
    layer1_outputs(5057) <= (layer0_outputs(5683)) and not (layer0_outputs(5547));
    layer1_outputs(5058) <= '1';
    layer1_outputs(5059) <= not(layer0_outputs(7162)) or (layer0_outputs(6680));
    layer1_outputs(5060) <= layer0_outputs(5008);
    layer1_outputs(5061) <= not(layer0_outputs(3172));
    layer1_outputs(5062) <= not(layer0_outputs(1777)) or (layer0_outputs(884));
    layer1_outputs(5063) <= (layer0_outputs(3635)) and (layer0_outputs(6303));
    layer1_outputs(5064) <= not(layer0_outputs(1889));
    layer1_outputs(5065) <= '1';
    layer1_outputs(5066) <= not(layer0_outputs(4209));
    layer1_outputs(5067) <= not((layer0_outputs(1599)) and (layer0_outputs(4712)));
    layer1_outputs(5068) <= not(layer0_outputs(3054)) or (layer0_outputs(2869));
    layer1_outputs(5069) <= not((layer0_outputs(241)) or (layer0_outputs(5013)));
    layer1_outputs(5070) <= layer0_outputs(2389);
    layer1_outputs(5071) <= not(layer0_outputs(1420));
    layer1_outputs(5072) <= (layer0_outputs(7508)) and not (layer0_outputs(777));
    layer1_outputs(5073) <= not(layer0_outputs(7174));
    layer1_outputs(5074) <= not((layer0_outputs(5603)) or (layer0_outputs(3312)));
    layer1_outputs(5075) <= (layer0_outputs(6189)) and not (layer0_outputs(1083));
    layer1_outputs(5076) <= (layer0_outputs(213)) and not (layer0_outputs(2743));
    layer1_outputs(5077) <= layer0_outputs(2746);
    layer1_outputs(5078) <= not((layer0_outputs(4574)) or (layer0_outputs(5894)));
    layer1_outputs(5079) <= (layer0_outputs(2417)) or (layer0_outputs(4761));
    layer1_outputs(5080) <= not(layer0_outputs(6860));
    layer1_outputs(5081) <= not(layer0_outputs(2983));
    layer1_outputs(5082) <= layer0_outputs(3100);
    layer1_outputs(5083) <= not(layer0_outputs(7013)) or (layer0_outputs(2246));
    layer1_outputs(5084) <= '0';
    layer1_outputs(5085) <= '1';
    layer1_outputs(5086) <= not(layer0_outputs(7475)) or (layer0_outputs(7251));
    layer1_outputs(5087) <= not(layer0_outputs(1021));
    layer1_outputs(5088) <= not((layer0_outputs(6605)) and (layer0_outputs(5457)));
    layer1_outputs(5089) <= not((layer0_outputs(3146)) or (layer0_outputs(2127)));
    layer1_outputs(5090) <= layer0_outputs(2093);
    layer1_outputs(5091) <= (layer0_outputs(6618)) and (layer0_outputs(2327));
    layer1_outputs(5092) <= not(layer0_outputs(1284)) or (layer0_outputs(1888));
    layer1_outputs(5093) <= layer0_outputs(3929);
    layer1_outputs(5094) <= not(layer0_outputs(6372));
    layer1_outputs(5095) <= not(layer0_outputs(1094)) or (layer0_outputs(6416));
    layer1_outputs(5096) <= not(layer0_outputs(5760));
    layer1_outputs(5097) <= not(layer0_outputs(6786));
    layer1_outputs(5098) <= not(layer0_outputs(4453)) or (layer0_outputs(2633));
    layer1_outputs(5099) <= not(layer0_outputs(4155)) or (layer0_outputs(7060));
    layer1_outputs(5100) <= not(layer0_outputs(4144));
    layer1_outputs(5101) <= not(layer0_outputs(6830));
    layer1_outputs(5102) <= '1';
    layer1_outputs(5103) <= not(layer0_outputs(3403));
    layer1_outputs(5104) <= not(layer0_outputs(2836)) or (layer0_outputs(1277));
    layer1_outputs(5105) <= layer0_outputs(4787);
    layer1_outputs(5106) <= not((layer0_outputs(37)) and (layer0_outputs(635)));
    layer1_outputs(5107) <= not(layer0_outputs(599)) or (layer0_outputs(166));
    layer1_outputs(5108) <= (layer0_outputs(3465)) and (layer0_outputs(1760));
    layer1_outputs(5109) <= not(layer0_outputs(1468));
    layer1_outputs(5110) <= not(layer0_outputs(2488));
    layer1_outputs(5111) <= not(layer0_outputs(3728));
    layer1_outputs(5112) <= not((layer0_outputs(3538)) and (layer0_outputs(770)));
    layer1_outputs(5113) <= (layer0_outputs(7565)) and not (layer0_outputs(2906));
    layer1_outputs(5114) <= (layer0_outputs(3616)) and not (layer0_outputs(94));
    layer1_outputs(5115) <= not((layer0_outputs(6144)) xor (layer0_outputs(5097)));
    layer1_outputs(5116) <= not(layer0_outputs(6053)) or (layer0_outputs(315));
    layer1_outputs(5117) <= '1';
    layer1_outputs(5118) <= layer0_outputs(1497);
    layer1_outputs(5119) <= not(layer0_outputs(3075)) or (layer0_outputs(5873));
    layer1_outputs(5120) <= (layer0_outputs(3187)) and not (layer0_outputs(5115));
    layer1_outputs(5121) <= not(layer0_outputs(3663)) or (layer0_outputs(6661));
    layer1_outputs(5122) <= not(layer0_outputs(270)) or (layer0_outputs(4541));
    layer1_outputs(5123) <= layer0_outputs(574);
    layer1_outputs(5124) <= layer0_outputs(1882);
    layer1_outputs(5125) <= not(layer0_outputs(1356));
    layer1_outputs(5126) <= not(layer0_outputs(2027));
    layer1_outputs(5127) <= layer0_outputs(5308);
    layer1_outputs(5128) <= not(layer0_outputs(3376));
    layer1_outputs(5129) <= not(layer0_outputs(6722));
    layer1_outputs(5130) <= not(layer0_outputs(7144));
    layer1_outputs(5131) <= '1';
    layer1_outputs(5132) <= not(layer0_outputs(5918));
    layer1_outputs(5133) <= not(layer0_outputs(2425));
    layer1_outputs(5134) <= '0';
    layer1_outputs(5135) <= (layer0_outputs(5422)) or (layer0_outputs(2674));
    layer1_outputs(5136) <= not((layer0_outputs(3985)) or (layer0_outputs(3476)));
    layer1_outputs(5137) <= (layer0_outputs(3849)) and not (layer0_outputs(823));
    layer1_outputs(5138) <= '1';
    layer1_outputs(5139) <= '1';
    layer1_outputs(5140) <= not(layer0_outputs(3128)) or (layer0_outputs(617));
    layer1_outputs(5141) <= (layer0_outputs(4959)) and not (layer0_outputs(3184));
    layer1_outputs(5142) <= not(layer0_outputs(3275)) or (layer0_outputs(6895));
    layer1_outputs(5143) <= (layer0_outputs(3575)) and (layer0_outputs(7067));
    layer1_outputs(5144) <= layer0_outputs(4927);
    layer1_outputs(5145) <= not((layer0_outputs(2429)) or (layer0_outputs(2523)));
    layer1_outputs(5146) <= layer0_outputs(4452);
    layer1_outputs(5147) <= (layer0_outputs(6554)) or (layer0_outputs(3577));
    layer1_outputs(5148) <= not(layer0_outputs(5874));
    layer1_outputs(5149) <= not((layer0_outputs(5112)) xor (layer0_outputs(2361)));
    layer1_outputs(5150) <= (layer0_outputs(6099)) and (layer0_outputs(5508));
    layer1_outputs(5151) <= (layer0_outputs(2532)) and (layer0_outputs(5280));
    layer1_outputs(5152) <= layer0_outputs(4382);
    layer1_outputs(5153) <= not(layer0_outputs(7227));
    layer1_outputs(5154) <= (layer0_outputs(2980)) and (layer0_outputs(1098));
    layer1_outputs(5155) <= (layer0_outputs(2840)) and not (layer0_outputs(6770));
    layer1_outputs(5156) <= not(layer0_outputs(4779));
    layer1_outputs(5157) <= not((layer0_outputs(1597)) and (layer0_outputs(4404)));
    layer1_outputs(5158) <= (layer0_outputs(3842)) and (layer0_outputs(7407));
    layer1_outputs(5159) <= layer0_outputs(7134);
    layer1_outputs(5160) <= layer0_outputs(4359);
    layer1_outputs(5161) <= not(layer0_outputs(4832));
    layer1_outputs(5162) <= (layer0_outputs(4686)) and (layer0_outputs(4800));
    layer1_outputs(5163) <= (layer0_outputs(2230)) and not (layer0_outputs(7225));
    layer1_outputs(5164) <= not(layer0_outputs(4342));
    layer1_outputs(5165) <= not((layer0_outputs(7589)) xor (layer0_outputs(5239)));
    layer1_outputs(5166) <= not(layer0_outputs(6798)) or (layer0_outputs(4643));
    layer1_outputs(5167) <= (layer0_outputs(7178)) and (layer0_outputs(5420));
    layer1_outputs(5168) <= layer0_outputs(5415);
    layer1_outputs(5169) <= (layer0_outputs(549)) and not (layer0_outputs(1786));
    layer1_outputs(5170) <= not(layer0_outputs(165));
    layer1_outputs(5171) <= not(layer0_outputs(4173));
    layer1_outputs(5172) <= '0';
    layer1_outputs(5173) <= not(layer0_outputs(2907));
    layer1_outputs(5174) <= not(layer0_outputs(3429)) or (layer0_outputs(7017));
    layer1_outputs(5175) <= not(layer0_outputs(3756));
    layer1_outputs(5176) <= layer0_outputs(2197);
    layer1_outputs(5177) <= not(layer0_outputs(918)) or (layer0_outputs(3273));
    layer1_outputs(5178) <= (layer0_outputs(3083)) xor (layer0_outputs(7365));
    layer1_outputs(5179) <= layer0_outputs(6520);
    layer1_outputs(5180) <= (layer0_outputs(333)) or (layer0_outputs(6808));
    layer1_outputs(5181) <= not(layer0_outputs(1372));
    layer1_outputs(5182) <= layer0_outputs(1133);
    layer1_outputs(5183) <= not((layer0_outputs(1873)) and (layer0_outputs(1033)));
    layer1_outputs(5184) <= layer0_outputs(2354);
    layer1_outputs(5185) <= not((layer0_outputs(2793)) xor (layer0_outputs(5476)));
    layer1_outputs(5186) <= (layer0_outputs(3269)) or (layer0_outputs(558));
    layer1_outputs(5187) <= not((layer0_outputs(7242)) and (layer0_outputs(805)));
    layer1_outputs(5188) <= (layer0_outputs(4324)) and not (layer0_outputs(2169));
    layer1_outputs(5189) <= layer0_outputs(3318);
    layer1_outputs(5190) <= not((layer0_outputs(3098)) or (layer0_outputs(4542)));
    layer1_outputs(5191) <= (layer0_outputs(2055)) and not (layer0_outputs(7655));
    layer1_outputs(5192) <= (layer0_outputs(5860)) or (layer0_outputs(992));
    layer1_outputs(5193) <= not((layer0_outputs(3380)) and (layer0_outputs(4140)));
    layer1_outputs(5194) <= not(layer0_outputs(539)) or (layer0_outputs(7411));
    layer1_outputs(5195) <= layer0_outputs(6349);
    layer1_outputs(5196) <= layer0_outputs(924);
    layer1_outputs(5197) <= (layer0_outputs(1606)) and (layer0_outputs(920));
    layer1_outputs(5198) <= (layer0_outputs(748)) and not (layer0_outputs(2451));
    layer1_outputs(5199) <= not((layer0_outputs(3504)) or (layer0_outputs(1952)));
    layer1_outputs(5200) <= layer0_outputs(1806);
    layer1_outputs(5201) <= (layer0_outputs(2649)) and (layer0_outputs(2802));
    layer1_outputs(5202) <= (layer0_outputs(1311)) and (layer0_outputs(906));
    layer1_outputs(5203) <= not((layer0_outputs(6523)) xor (layer0_outputs(2653)));
    layer1_outputs(5204) <= (layer0_outputs(656)) and not (layer0_outputs(2597));
    layer1_outputs(5205) <= (layer0_outputs(408)) and not (layer0_outputs(3572));
    layer1_outputs(5206) <= layer0_outputs(1798);
    layer1_outputs(5207) <= not(layer0_outputs(3138));
    layer1_outputs(5208) <= layer0_outputs(1759);
    layer1_outputs(5209) <= not(layer0_outputs(3062));
    layer1_outputs(5210) <= (layer0_outputs(7285)) or (layer0_outputs(540));
    layer1_outputs(5211) <= (layer0_outputs(4354)) and (layer0_outputs(2705));
    layer1_outputs(5212) <= not((layer0_outputs(5338)) or (layer0_outputs(1112)));
    layer1_outputs(5213) <= not(layer0_outputs(3440)) or (layer0_outputs(4379));
    layer1_outputs(5214) <= (layer0_outputs(1740)) or (layer0_outputs(4289));
    layer1_outputs(5215) <= layer0_outputs(7308);
    layer1_outputs(5216) <= layer0_outputs(2747);
    layer1_outputs(5217) <= not(layer0_outputs(6482));
    layer1_outputs(5218) <= not(layer0_outputs(4122));
    layer1_outputs(5219) <= layer0_outputs(7515);
    layer1_outputs(5220) <= (layer0_outputs(257)) and (layer0_outputs(7632));
    layer1_outputs(5221) <= '1';
    layer1_outputs(5222) <= (layer0_outputs(2565)) xor (layer0_outputs(3233));
    layer1_outputs(5223) <= (layer0_outputs(5214)) or (layer0_outputs(83));
    layer1_outputs(5224) <= (layer0_outputs(737)) and not (layer0_outputs(4856));
    layer1_outputs(5225) <= not(layer0_outputs(4457));
    layer1_outputs(5226) <= layer0_outputs(463);
    layer1_outputs(5227) <= not(layer0_outputs(5363));
    layer1_outputs(5228) <= not(layer0_outputs(7640));
    layer1_outputs(5229) <= not(layer0_outputs(829));
    layer1_outputs(5230) <= not(layer0_outputs(5310));
    layer1_outputs(5231) <= layer0_outputs(926);
    layer1_outputs(5232) <= layer0_outputs(4609);
    layer1_outputs(5233) <= not(layer0_outputs(2245));
    layer1_outputs(5234) <= layer0_outputs(7414);
    layer1_outputs(5235) <= not((layer0_outputs(4317)) and (layer0_outputs(1118)));
    layer1_outputs(5236) <= '1';
    layer1_outputs(5237) <= not(layer0_outputs(4023)) or (layer0_outputs(4771));
    layer1_outputs(5238) <= not((layer0_outputs(2294)) and (layer0_outputs(1573)));
    layer1_outputs(5239) <= not(layer0_outputs(490)) or (layer0_outputs(2568));
    layer1_outputs(5240) <= not(layer0_outputs(5149));
    layer1_outputs(5241) <= '0';
    layer1_outputs(5242) <= (layer0_outputs(7042)) and not (layer0_outputs(781));
    layer1_outputs(5243) <= '1';
    layer1_outputs(5244) <= not(layer0_outputs(7491));
    layer1_outputs(5245) <= '1';
    layer1_outputs(5246) <= layer0_outputs(2932);
    layer1_outputs(5247) <= '0';
    layer1_outputs(5248) <= layer0_outputs(935);
    layer1_outputs(5249) <= (layer0_outputs(2593)) or (layer0_outputs(5814));
    layer1_outputs(5250) <= layer0_outputs(4523);
    layer1_outputs(5251) <= layer0_outputs(3252);
    layer1_outputs(5252) <= not((layer0_outputs(3966)) and (layer0_outputs(5849)));
    layer1_outputs(5253) <= (layer0_outputs(6958)) and (layer0_outputs(3484));
    layer1_outputs(5254) <= layer0_outputs(663);
    layer1_outputs(5255) <= not((layer0_outputs(5156)) and (layer0_outputs(1284)));
    layer1_outputs(5256) <= layer0_outputs(130);
    layer1_outputs(5257) <= (layer0_outputs(3349)) and (layer0_outputs(3960));
    layer1_outputs(5258) <= not(layer0_outputs(33));
    layer1_outputs(5259) <= (layer0_outputs(4322)) or (layer0_outputs(1953));
    layer1_outputs(5260) <= (layer0_outputs(356)) or (layer0_outputs(6447));
    layer1_outputs(5261) <= (layer0_outputs(6662)) and not (layer0_outputs(4238));
    layer1_outputs(5262) <= layer0_outputs(6773);
    layer1_outputs(5263) <= not(layer0_outputs(692)) or (layer0_outputs(6404));
    layer1_outputs(5264) <= not(layer0_outputs(4644));
    layer1_outputs(5265) <= (layer0_outputs(4536)) and (layer0_outputs(7306));
    layer1_outputs(5266) <= not((layer0_outputs(5527)) xor (layer0_outputs(5734)));
    layer1_outputs(5267) <= not((layer0_outputs(7296)) or (layer0_outputs(5071)));
    layer1_outputs(5268) <= (layer0_outputs(646)) and not (layer0_outputs(4096));
    layer1_outputs(5269) <= not(layer0_outputs(1484)) or (layer0_outputs(7155));
    layer1_outputs(5270) <= layer0_outputs(4159);
    layer1_outputs(5271) <= layer0_outputs(4143);
    layer1_outputs(5272) <= not((layer0_outputs(4385)) and (layer0_outputs(2608)));
    layer1_outputs(5273) <= not(layer0_outputs(5454));
    layer1_outputs(5274) <= not(layer0_outputs(1754));
    layer1_outputs(5275) <= (layer0_outputs(652)) or (layer0_outputs(3));
    layer1_outputs(5276) <= (layer0_outputs(6947)) and (layer0_outputs(1424));
    layer1_outputs(5277) <= (layer0_outputs(3257)) and (layer0_outputs(5044));
    layer1_outputs(5278) <= layer0_outputs(2779);
    layer1_outputs(5279) <= not(layer0_outputs(4964));
    layer1_outputs(5280) <= not(layer0_outputs(3464)) or (layer0_outputs(3235));
    layer1_outputs(5281) <= (layer0_outputs(1211)) and not (layer0_outputs(1804));
    layer1_outputs(5282) <= layer0_outputs(149);
    layer1_outputs(5283) <= not(layer0_outputs(5363)) or (layer0_outputs(260));
    layer1_outputs(5284) <= not(layer0_outputs(2377));
    layer1_outputs(5285) <= not(layer0_outputs(4027)) or (layer0_outputs(3454));
    layer1_outputs(5286) <= (layer0_outputs(860)) and not (layer0_outputs(7457));
    layer1_outputs(5287) <= not(layer0_outputs(7527)) or (layer0_outputs(2624));
    layer1_outputs(5288) <= not(layer0_outputs(3578));
    layer1_outputs(5289) <= not(layer0_outputs(1047)) or (layer0_outputs(3867));
    layer1_outputs(5290) <= '0';
    layer1_outputs(5291) <= not((layer0_outputs(2582)) xor (layer0_outputs(756)));
    layer1_outputs(5292) <= (layer0_outputs(6517)) or (layer0_outputs(493));
    layer1_outputs(5293) <= layer0_outputs(4270);
    layer1_outputs(5294) <= '0';
    layer1_outputs(5295) <= '0';
    layer1_outputs(5296) <= (layer0_outputs(5689)) and (layer0_outputs(3825));
    layer1_outputs(5297) <= layer0_outputs(5121);
    layer1_outputs(5298) <= layer0_outputs(2430);
    layer1_outputs(5299) <= (layer0_outputs(7203)) and (layer0_outputs(4912));
    layer1_outputs(5300) <= layer0_outputs(962);
    layer1_outputs(5301) <= not((layer0_outputs(3832)) and (layer0_outputs(2025)));
    layer1_outputs(5302) <= not(layer0_outputs(5352));
    layer1_outputs(5303) <= not(layer0_outputs(2769)) or (layer0_outputs(4783));
    layer1_outputs(5304) <= layer0_outputs(768);
    layer1_outputs(5305) <= (layer0_outputs(5318)) xor (layer0_outputs(1863));
    layer1_outputs(5306) <= (layer0_outputs(4812)) and not (layer0_outputs(3643));
    layer1_outputs(5307) <= not(layer0_outputs(6028));
    layer1_outputs(5308) <= not((layer0_outputs(2013)) and (layer0_outputs(1249)));
    layer1_outputs(5309) <= (layer0_outputs(5661)) xor (layer0_outputs(5453));
    layer1_outputs(5310) <= (layer0_outputs(3137)) and not (layer0_outputs(3238));
    layer1_outputs(5311) <= not(layer0_outputs(7214));
    layer1_outputs(5312) <= not(layer0_outputs(1827));
    layer1_outputs(5313) <= not(layer0_outputs(4827));
    layer1_outputs(5314) <= layer0_outputs(597);
    layer1_outputs(5315) <= not(layer0_outputs(268));
    layer1_outputs(5316) <= '0';
    layer1_outputs(5317) <= not(layer0_outputs(3150));
    layer1_outputs(5318) <= not((layer0_outputs(2638)) and (layer0_outputs(2798)));
    layer1_outputs(5319) <= (layer0_outputs(6088)) and not (layer0_outputs(7380));
    layer1_outputs(5320) <= (layer0_outputs(2762)) and (layer0_outputs(3105));
    layer1_outputs(5321) <= (layer0_outputs(4904)) and not (layer0_outputs(694));
    layer1_outputs(5322) <= '1';
    layer1_outputs(5323) <= layer0_outputs(767);
    layer1_outputs(5324) <= layer0_outputs(6663);
    layer1_outputs(5325) <= (layer0_outputs(6761)) and (layer0_outputs(3206));
    layer1_outputs(5326) <= not(layer0_outputs(48));
    layer1_outputs(5327) <= not((layer0_outputs(1210)) and (layer0_outputs(702)));
    layer1_outputs(5328) <= not(layer0_outputs(3707)) or (layer0_outputs(2128));
    layer1_outputs(5329) <= (layer0_outputs(3758)) and (layer0_outputs(3560));
    layer1_outputs(5330) <= not(layer0_outputs(5166));
    layer1_outputs(5331) <= (layer0_outputs(376)) and (layer0_outputs(1208));
    layer1_outputs(5332) <= not((layer0_outputs(3525)) or (layer0_outputs(1869)));
    layer1_outputs(5333) <= not((layer0_outputs(384)) xor (layer0_outputs(2800)));
    layer1_outputs(5334) <= not(layer0_outputs(4188));
    layer1_outputs(5335) <= (layer0_outputs(4714)) and (layer0_outputs(5246));
    layer1_outputs(5336) <= not((layer0_outputs(2827)) xor (layer0_outputs(1471)));
    layer1_outputs(5337) <= layer0_outputs(1727);
    layer1_outputs(5338) <= layer0_outputs(4585);
    layer1_outputs(5339) <= layer0_outputs(6772);
    layer1_outputs(5340) <= (layer0_outputs(6238)) and not (layer0_outputs(3796));
    layer1_outputs(5341) <= not(layer0_outputs(1983));
    layer1_outputs(5342) <= not(layer0_outputs(469));
    layer1_outputs(5343) <= (layer0_outputs(6627)) or (layer0_outputs(4861));
    layer1_outputs(5344) <= not(layer0_outputs(145)) or (layer0_outputs(1164));
    layer1_outputs(5345) <= layer0_outputs(4738);
    layer1_outputs(5346) <= not(layer0_outputs(1882));
    layer1_outputs(5347) <= layer0_outputs(2489);
    layer1_outputs(5348) <= not(layer0_outputs(7637));
    layer1_outputs(5349) <= not(layer0_outputs(768));
    layer1_outputs(5350) <= layer0_outputs(6456);
    layer1_outputs(5351) <= '1';
    layer1_outputs(5352) <= layer0_outputs(6828);
    layer1_outputs(5353) <= not((layer0_outputs(4013)) or (layer0_outputs(2364)));
    layer1_outputs(5354) <= layer0_outputs(3288);
    layer1_outputs(5355) <= not(layer0_outputs(3339));
    layer1_outputs(5356) <= (layer0_outputs(7462)) and not (layer0_outputs(6706));
    layer1_outputs(5357) <= (layer0_outputs(1336)) or (layer0_outputs(6199));
    layer1_outputs(5358) <= not(layer0_outputs(2353));
    layer1_outputs(5359) <= (layer0_outputs(6420)) and not (layer0_outputs(5234));
    layer1_outputs(5360) <= (layer0_outputs(6401)) and not (layer0_outputs(4975));
    layer1_outputs(5361) <= not(layer0_outputs(1992));
    layer1_outputs(5362) <= layer0_outputs(4602);
    layer1_outputs(5363) <= '0';
    layer1_outputs(5364) <= (layer0_outputs(6656)) and not (layer0_outputs(4640));
    layer1_outputs(5365) <= (layer0_outputs(7614)) and not (layer0_outputs(1913));
    layer1_outputs(5366) <= layer0_outputs(6775);
    layer1_outputs(5367) <= layer0_outputs(2522);
    layer1_outputs(5368) <= (layer0_outputs(6324)) and (layer0_outputs(563));
    layer1_outputs(5369) <= not(layer0_outputs(2258)) or (layer0_outputs(6728));
    layer1_outputs(5370) <= (layer0_outputs(1071)) and (layer0_outputs(3889));
    layer1_outputs(5371) <= layer0_outputs(5521);
    layer1_outputs(5372) <= '0';
    layer1_outputs(5373) <= not(layer0_outputs(2525));
    layer1_outputs(5374) <= '1';
    layer1_outputs(5375) <= not(layer0_outputs(3180)) or (layer0_outputs(7604));
    layer1_outputs(5376) <= layer0_outputs(5017);
    layer1_outputs(5377) <= (layer0_outputs(5089)) and not (layer0_outputs(4112));
    layer1_outputs(5378) <= layer0_outputs(5430);
    layer1_outputs(5379) <= not((layer0_outputs(3452)) or (layer0_outputs(6601)));
    layer1_outputs(5380) <= (layer0_outputs(4034)) and (layer0_outputs(4302));
    layer1_outputs(5381) <= (layer0_outputs(509)) and not (layer0_outputs(4851));
    layer1_outputs(5382) <= (layer0_outputs(5516)) xor (layer0_outputs(595));
    layer1_outputs(5383) <= not(layer0_outputs(1713)) or (layer0_outputs(4343));
    layer1_outputs(5384) <= not((layer0_outputs(326)) or (layer0_outputs(277)));
    layer1_outputs(5385) <= not(layer0_outputs(5011));
    layer1_outputs(5386) <= not(layer0_outputs(1064)) or (layer0_outputs(6989));
    layer1_outputs(5387) <= '1';
    layer1_outputs(5388) <= not(layer0_outputs(5655));
    layer1_outputs(5389) <= '1';
    layer1_outputs(5390) <= layer0_outputs(5433);
    layer1_outputs(5391) <= (layer0_outputs(3342)) xor (layer0_outputs(4297));
    layer1_outputs(5392) <= (layer0_outputs(6426)) and not (layer0_outputs(1257));
    layer1_outputs(5393) <= not(layer0_outputs(544));
    layer1_outputs(5394) <= (layer0_outputs(5371)) or (layer0_outputs(110));
    layer1_outputs(5395) <= (layer0_outputs(2510)) and (layer0_outputs(4868));
    layer1_outputs(5396) <= not((layer0_outputs(178)) or (layer0_outputs(2674)));
    layer1_outputs(5397) <= '1';
    layer1_outputs(5398) <= layer0_outputs(3212);
    layer1_outputs(5399) <= (layer0_outputs(5919)) and not (layer0_outputs(4789));
    layer1_outputs(5400) <= '1';
    layer1_outputs(5401) <= layer0_outputs(93);
    layer1_outputs(5402) <= layer0_outputs(3599);
    layer1_outputs(5403) <= not(layer0_outputs(6831)) or (layer0_outputs(780));
    layer1_outputs(5404) <= not((layer0_outputs(3896)) and (layer0_outputs(4567)));
    layer1_outputs(5405) <= (layer0_outputs(2599)) xor (layer0_outputs(7022));
    layer1_outputs(5406) <= (layer0_outputs(5250)) and not (layer0_outputs(1905));
    layer1_outputs(5407) <= layer0_outputs(3150);
    layer1_outputs(5408) <= (layer0_outputs(5966)) and (layer0_outputs(6792));
    layer1_outputs(5409) <= (layer0_outputs(6268)) or (layer0_outputs(7286));
    layer1_outputs(5410) <= not(layer0_outputs(2738));
    layer1_outputs(5411) <= not(layer0_outputs(2003)) or (layer0_outputs(5833));
    layer1_outputs(5412) <= (layer0_outputs(1084)) and not (layer0_outputs(5043));
    layer1_outputs(5413) <= not(layer0_outputs(3341));
    layer1_outputs(5414) <= not(layer0_outputs(1350)) or (layer0_outputs(5745));
    layer1_outputs(5415) <= '1';
    layer1_outputs(5416) <= '1';
    layer1_outputs(5417) <= (layer0_outputs(2047)) and not (layer0_outputs(6453));
    layer1_outputs(5418) <= (layer0_outputs(7639)) xor (layer0_outputs(6277));
    layer1_outputs(5419) <= layer0_outputs(5129);
    layer1_outputs(5420) <= not(layer0_outputs(2345)) or (layer0_outputs(4248));
    layer1_outputs(5421) <= layer0_outputs(624);
    layer1_outputs(5422) <= (layer0_outputs(4627)) and not (layer0_outputs(6546));
    layer1_outputs(5423) <= layer0_outputs(2652);
    layer1_outputs(5424) <= not(layer0_outputs(2138)) or (layer0_outputs(4905));
    layer1_outputs(5425) <= (layer0_outputs(2220)) and (layer0_outputs(4482));
    layer1_outputs(5426) <= not(layer0_outputs(3240));
    layer1_outputs(5427) <= (layer0_outputs(81)) and (layer0_outputs(1787));
    layer1_outputs(5428) <= (layer0_outputs(7406)) and not (layer0_outputs(6230));
    layer1_outputs(5429) <= '1';
    layer1_outputs(5430) <= not(layer0_outputs(1975));
    layer1_outputs(5431) <= not(layer0_outputs(6859)) or (layer0_outputs(2631));
    layer1_outputs(5432) <= not(layer0_outputs(405));
    layer1_outputs(5433) <= not((layer0_outputs(932)) or (layer0_outputs(7311)));
    layer1_outputs(5434) <= '1';
    layer1_outputs(5435) <= '0';
    layer1_outputs(5436) <= not(layer0_outputs(5609)) or (layer0_outputs(1900));
    layer1_outputs(5437) <= '0';
    layer1_outputs(5438) <= (layer0_outputs(7484)) and not (layer0_outputs(6849));
    layer1_outputs(5439) <= layer0_outputs(4475);
    layer1_outputs(5440) <= not((layer0_outputs(1746)) and (layer0_outputs(1185)));
    layer1_outputs(5441) <= layer0_outputs(2664);
    layer1_outputs(5442) <= not((layer0_outputs(233)) xor (layer0_outputs(2737)));
    layer1_outputs(5443) <= '0';
    layer1_outputs(5444) <= not(layer0_outputs(5808));
    layer1_outputs(5445) <= (layer0_outputs(509)) and (layer0_outputs(5685));
    layer1_outputs(5446) <= layer0_outputs(3552);
    layer1_outputs(5447) <= not(layer0_outputs(3163));
    layer1_outputs(5448) <= not((layer0_outputs(6115)) and (layer0_outputs(6690)));
    layer1_outputs(5449) <= not(layer0_outputs(5373));
    layer1_outputs(5450) <= not((layer0_outputs(7616)) and (layer0_outputs(1354)));
    layer1_outputs(5451) <= not(layer0_outputs(4573));
    layer1_outputs(5452) <= (layer0_outputs(6902)) and not (layer0_outputs(4350));
    layer1_outputs(5453) <= not(layer0_outputs(538)) or (layer0_outputs(2395));
    layer1_outputs(5454) <= not(layer0_outputs(2104));
    layer1_outputs(5455) <= not((layer0_outputs(7393)) xor (layer0_outputs(6240)));
    layer1_outputs(5456) <= layer0_outputs(7066);
    layer1_outputs(5457) <= not(layer0_outputs(6128));
    layer1_outputs(5458) <= not(layer0_outputs(3660));
    layer1_outputs(5459) <= not(layer0_outputs(5850));
    layer1_outputs(5460) <= not(layer0_outputs(7645)) or (layer0_outputs(4984));
    layer1_outputs(5461) <= (layer0_outputs(5226)) and not (layer0_outputs(5000));
    layer1_outputs(5462) <= layer0_outputs(59);
    layer1_outputs(5463) <= (layer0_outputs(4650)) or (layer0_outputs(4094));
    layer1_outputs(5464) <= layer0_outputs(5188);
    layer1_outputs(5465) <= (layer0_outputs(5488)) or (layer0_outputs(5392));
    layer1_outputs(5466) <= not((layer0_outputs(1159)) and (layer0_outputs(1526)));
    layer1_outputs(5467) <= not((layer0_outputs(685)) or (layer0_outputs(1158)));
    layer1_outputs(5468) <= (layer0_outputs(6798)) and not (layer0_outputs(6078));
    layer1_outputs(5469) <= layer0_outputs(5907);
    layer1_outputs(5470) <= not(layer0_outputs(6309));
    layer1_outputs(5471) <= not(layer0_outputs(2049)) or (layer0_outputs(2566));
    layer1_outputs(5472) <= (layer0_outputs(2806)) and (layer0_outputs(5425));
    layer1_outputs(5473) <= layer0_outputs(6666);
    layer1_outputs(5474) <= not(layer0_outputs(2942));
    layer1_outputs(5475) <= (layer0_outputs(7473)) and (layer0_outputs(6924));
    layer1_outputs(5476) <= not(layer0_outputs(5165));
    layer1_outputs(5477) <= layer0_outputs(7468);
    layer1_outputs(5478) <= not((layer0_outputs(18)) or (layer0_outputs(7027)));
    layer1_outputs(5479) <= layer0_outputs(1126);
    layer1_outputs(5480) <= (layer0_outputs(2185)) and (layer0_outputs(5329));
    layer1_outputs(5481) <= (layer0_outputs(2340)) and not (layer0_outputs(3143));
    layer1_outputs(5482) <= not((layer0_outputs(3199)) or (layer0_outputs(869)));
    layer1_outputs(5483) <= (layer0_outputs(4579)) and not (layer0_outputs(4401));
    layer1_outputs(5484) <= not((layer0_outputs(6557)) or (layer0_outputs(4398)));
    layer1_outputs(5485) <= not((layer0_outputs(1592)) or (layer0_outputs(181)));
    layer1_outputs(5486) <= (layer0_outputs(7505)) or (layer0_outputs(1764));
    layer1_outputs(5487) <= (layer0_outputs(4420)) and not (layer0_outputs(3768));
    layer1_outputs(5488) <= layer0_outputs(563);
    layer1_outputs(5489) <= (layer0_outputs(693)) xor (layer0_outputs(6094));
    layer1_outputs(5490) <= not(layer0_outputs(1507)) or (layer0_outputs(6170));
    layer1_outputs(5491) <= layer0_outputs(4418);
    layer1_outputs(5492) <= (layer0_outputs(3680)) and not (layer0_outputs(4390));
    layer1_outputs(5493) <= '1';
    layer1_outputs(5494) <= not((layer0_outputs(984)) and (layer0_outputs(5396)));
    layer1_outputs(5495) <= layer0_outputs(4122);
    layer1_outputs(5496) <= not((layer0_outputs(2035)) and (layer0_outputs(1345)));
    layer1_outputs(5497) <= not(layer0_outputs(5929));
    layer1_outputs(5498) <= (layer0_outputs(4904)) and not (layer0_outputs(6149));
    layer1_outputs(5499) <= not((layer0_outputs(926)) or (layer0_outputs(2084)));
    layer1_outputs(5500) <= (layer0_outputs(952)) and not (layer0_outputs(5045));
    layer1_outputs(5501) <= not(layer0_outputs(885)) or (layer0_outputs(5935));
    layer1_outputs(5502) <= '1';
    layer1_outputs(5503) <= '1';
    layer1_outputs(5504) <= not(layer0_outputs(7130));
    layer1_outputs(5505) <= not(layer0_outputs(5901)) or (layer0_outputs(2366));
    layer1_outputs(5506) <= layer0_outputs(7276);
    layer1_outputs(5507) <= '1';
    layer1_outputs(5508) <= (layer0_outputs(4932)) xor (layer0_outputs(535));
    layer1_outputs(5509) <= (layer0_outputs(3231)) and not (layer0_outputs(5384));
    layer1_outputs(5510) <= not(layer0_outputs(3600));
    layer1_outputs(5511) <= not((layer0_outputs(1370)) or (layer0_outputs(445)));
    layer1_outputs(5512) <= layer0_outputs(7476);
    layer1_outputs(5513) <= layer0_outputs(6406);
    layer1_outputs(5514) <= not(layer0_outputs(3926));
    layer1_outputs(5515) <= '0';
    layer1_outputs(5516) <= (layer0_outputs(1850)) and not (layer0_outputs(1717));
    layer1_outputs(5517) <= not((layer0_outputs(1678)) or (layer0_outputs(6740)));
    layer1_outputs(5518) <= not(layer0_outputs(3716));
    layer1_outputs(5519) <= not(layer0_outputs(2759));
    layer1_outputs(5520) <= not(layer0_outputs(2213)) or (layer0_outputs(4674));
    layer1_outputs(5521) <= not(layer0_outputs(351));
    layer1_outputs(5522) <= layer0_outputs(4072);
    layer1_outputs(5523) <= not(layer0_outputs(4115));
    layer1_outputs(5524) <= '1';
    layer1_outputs(5525) <= (layer0_outputs(5619)) and not (layer0_outputs(2339));
    layer1_outputs(5526) <= not(layer0_outputs(6527));
    layer1_outputs(5527) <= (layer0_outputs(4629)) and (layer0_outputs(1280));
    layer1_outputs(5528) <= not(layer0_outputs(6780)) or (layer0_outputs(65));
    layer1_outputs(5529) <= not((layer0_outputs(4320)) or (layer0_outputs(3569)));
    layer1_outputs(5530) <= '1';
    layer1_outputs(5531) <= not(layer0_outputs(4051));
    layer1_outputs(5532) <= not(layer0_outputs(4515)) or (layer0_outputs(3525));
    layer1_outputs(5533) <= not(layer0_outputs(5939));
    layer1_outputs(5534) <= (layer0_outputs(6703)) and not (layer0_outputs(7348));
    layer1_outputs(5535) <= layer0_outputs(1074);
    layer1_outputs(5536) <= not((layer0_outputs(3824)) and (layer0_outputs(4713)));
    layer1_outputs(5537) <= not((layer0_outputs(7297)) and (layer0_outputs(190)));
    layer1_outputs(5538) <= not(layer0_outputs(1776));
    layer1_outputs(5539) <= not(layer0_outputs(6133)) or (layer0_outputs(4762));
    layer1_outputs(5540) <= not((layer0_outputs(37)) or (layer0_outputs(5544)));
    layer1_outputs(5541) <= '0';
    layer1_outputs(5542) <= (layer0_outputs(2144)) and not (layer0_outputs(6615));
    layer1_outputs(5543) <= not(layer0_outputs(1359));
    layer1_outputs(5544) <= not(layer0_outputs(3155)) or (layer0_outputs(4479));
    layer1_outputs(5545) <= not(layer0_outputs(6760));
    layer1_outputs(5546) <= '0';
    layer1_outputs(5547) <= not(layer0_outputs(4793));
    layer1_outputs(5548) <= not(layer0_outputs(4619));
    layer1_outputs(5549) <= layer0_outputs(190);
    layer1_outputs(5550) <= not((layer0_outputs(7593)) and (layer0_outputs(5347)));
    layer1_outputs(5551) <= '0';
    layer1_outputs(5552) <= not(layer0_outputs(2207));
    layer1_outputs(5553) <= layer0_outputs(6363);
    layer1_outputs(5554) <= layer0_outputs(2281);
    layer1_outputs(5555) <= not(layer0_outputs(3472));
    layer1_outputs(5556) <= (layer0_outputs(7290)) and not (layer0_outputs(1956));
    layer1_outputs(5557) <= (layer0_outputs(3622)) and not (layer0_outputs(4493));
    layer1_outputs(5558) <= '1';
    layer1_outputs(5559) <= layer0_outputs(3339);
    layer1_outputs(5560) <= layer0_outputs(7285);
    layer1_outputs(5561) <= '0';
    layer1_outputs(5562) <= layer0_outputs(5196);
    layer1_outputs(5563) <= '0';
    layer1_outputs(5564) <= (layer0_outputs(5244)) and not (layer0_outputs(3354));
    layer1_outputs(5565) <= (layer0_outputs(1816)) and not (layer0_outputs(2314));
    layer1_outputs(5566) <= not(layer0_outputs(5269));
    layer1_outputs(5567) <= not(layer0_outputs(5486));
    layer1_outputs(5568) <= not(layer0_outputs(5730));
    layer1_outputs(5569) <= (layer0_outputs(338)) and (layer0_outputs(3486));
    layer1_outputs(5570) <= not(layer0_outputs(2880));
    layer1_outputs(5571) <= (layer0_outputs(4823)) and not (layer0_outputs(1310));
    layer1_outputs(5572) <= layer0_outputs(370);
    layer1_outputs(5573) <= layer0_outputs(845);
    layer1_outputs(5574) <= not((layer0_outputs(1653)) and (layer0_outputs(4118)));
    layer1_outputs(5575) <= layer0_outputs(7034);
    layer1_outputs(5576) <= not(layer0_outputs(3479));
    layer1_outputs(5577) <= layer0_outputs(3458);
    layer1_outputs(5578) <= not(layer0_outputs(4398));
    layer1_outputs(5579) <= layer0_outputs(6297);
    layer1_outputs(5580) <= not((layer0_outputs(5576)) and (layer0_outputs(3065)));
    layer1_outputs(5581) <= '0';
    layer1_outputs(5582) <= '0';
    layer1_outputs(5583) <= layer0_outputs(1008);
    layer1_outputs(5584) <= not(layer0_outputs(1110));
    layer1_outputs(5585) <= not(layer0_outputs(531)) or (layer0_outputs(3536));
    layer1_outputs(5586) <= (layer0_outputs(5836)) and not (layer0_outputs(4258));
    layer1_outputs(5587) <= layer0_outputs(4762);
    layer1_outputs(5588) <= (layer0_outputs(3453)) or (layer0_outputs(7574));
    layer1_outputs(5589) <= layer0_outputs(6525);
    layer1_outputs(5590) <= not(layer0_outputs(2134));
    layer1_outputs(5591) <= not(layer0_outputs(4837)) or (layer0_outputs(3884));
    layer1_outputs(5592) <= (layer0_outputs(5594)) xor (layer0_outputs(2982));
    layer1_outputs(5593) <= not((layer0_outputs(7315)) or (layer0_outputs(5746)));
    layer1_outputs(5594) <= (layer0_outputs(7097)) and not (layer0_outputs(4548));
    layer1_outputs(5595) <= not(layer0_outputs(2557));
    layer1_outputs(5596) <= layer0_outputs(1157);
    layer1_outputs(5597) <= (layer0_outputs(4355)) and not (layer0_outputs(3605));
    layer1_outputs(5598) <= (layer0_outputs(3821)) and not (layer0_outputs(3005));
    layer1_outputs(5599) <= '1';
    layer1_outputs(5600) <= layer0_outputs(7340);
    layer1_outputs(5601) <= '0';
    layer1_outputs(5602) <= layer0_outputs(2815);
    layer1_outputs(5603) <= (layer0_outputs(4458)) and not (layer0_outputs(5503));
    layer1_outputs(5604) <= not((layer0_outputs(2037)) or (layer0_outputs(688)));
    layer1_outputs(5605) <= not(layer0_outputs(6983));
    layer1_outputs(5606) <= not(layer0_outputs(4160));
    layer1_outputs(5607) <= not(layer0_outputs(4340));
    layer1_outputs(5608) <= not(layer0_outputs(6520));
    layer1_outputs(5609) <= '0';
    layer1_outputs(5610) <= layer0_outputs(5016);
    layer1_outputs(5611) <= layer0_outputs(1280);
    layer1_outputs(5612) <= not(layer0_outputs(6749));
    layer1_outputs(5613) <= layer0_outputs(4636);
    layer1_outputs(5614) <= not(layer0_outputs(2081));
    layer1_outputs(5615) <= (layer0_outputs(4089)) or (layer0_outputs(6020));
    layer1_outputs(5616) <= not((layer0_outputs(6163)) or (layer0_outputs(1077)));
    layer1_outputs(5617) <= not(layer0_outputs(2149)) or (layer0_outputs(1339));
    layer1_outputs(5618) <= '0';
    layer1_outputs(5619) <= '1';
    layer1_outputs(5620) <= (layer0_outputs(1405)) or (layer0_outputs(7352));
    layer1_outputs(5621) <= not(layer0_outputs(3702));
    layer1_outputs(5622) <= not((layer0_outputs(3691)) or (layer0_outputs(1704)));
    layer1_outputs(5623) <= not(layer0_outputs(4416));
    layer1_outputs(5624) <= layer0_outputs(19);
    layer1_outputs(5625) <= not(layer0_outputs(3571)) or (layer0_outputs(5007));
    layer1_outputs(5626) <= '1';
    layer1_outputs(5627) <= (layer0_outputs(899)) and (layer0_outputs(2086));
    layer1_outputs(5628) <= '1';
    layer1_outputs(5629) <= layer0_outputs(1178);
    layer1_outputs(5630) <= (layer0_outputs(4202)) and not (layer0_outputs(5635));
    layer1_outputs(5631) <= layer0_outputs(311);
    layer1_outputs(5632) <= '0';
    layer1_outputs(5633) <= (layer0_outputs(6536)) and (layer0_outputs(1860));
    layer1_outputs(5634) <= '0';
    layer1_outputs(5635) <= layer0_outputs(2891);
    layer1_outputs(5636) <= not((layer0_outputs(6373)) and (layer0_outputs(7413)));
    layer1_outputs(5637) <= not(layer0_outputs(2405));
    layer1_outputs(5638) <= not(layer0_outputs(3557));
    layer1_outputs(5639) <= (layer0_outputs(5789)) and not (layer0_outputs(3045));
    layer1_outputs(5640) <= not((layer0_outputs(1896)) or (layer0_outputs(3239)));
    layer1_outputs(5641) <= '1';
    layer1_outputs(5642) <= not(layer0_outputs(3421));
    layer1_outputs(5643) <= '0';
    layer1_outputs(5644) <= (layer0_outputs(7611)) or (layer0_outputs(164));
    layer1_outputs(5645) <= not(layer0_outputs(5895));
    layer1_outputs(5646) <= not(layer0_outputs(4151)) or (layer0_outputs(219));
    layer1_outputs(5647) <= layer0_outputs(2171);
    layer1_outputs(5648) <= not((layer0_outputs(4034)) and (layer0_outputs(6889)));
    layer1_outputs(5649) <= layer0_outputs(5879);
    layer1_outputs(5650) <= layer0_outputs(2123);
    layer1_outputs(5651) <= layer0_outputs(4016);
    layer1_outputs(5652) <= layer0_outputs(4570);
    layer1_outputs(5653) <= not(layer0_outputs(4868)) or (layer0_outputs(2101));
    layer1_outputs(5654) <= not((layer0_outputs(2924)) xor (layer0_outputs(2234)));
    layer1_outputs(5655) <= layer0_outputs(5151);
    layer1_outputs(5656) <= (layer0_outputs(6950)) or (layer0_outputs(106));
    layer1_outputs(5657) <= '1';
    layer1_outputs(5658) <= '0';
    layer1_outputs(5659) <= not(layer0_outputs(5254));
    layer1_outputs(5660) <= not(layer0_outputs(1496));
    layer1_outputs(5661) <= not((layer0_outputs(4846)) and (layer0_outputs(3)));
    layer1_outputs(5662) <= not(layer0_outputs(5458)) or (layer0_outputs(199));
    layer1_outputs(5663) <= not(layer0_outputs(6661)) or (layer0_outputs(6503));
    layer1_outputs(5664) <= not(layer0_outputs(4633));
    layer1_outputs(5665) <= not(layer0_outputs(2454));
    layer1_outputs(5666) <= (layer0_outputs(4015)) and not (layer0_outputs(2022));
    layer1_outputs(5667) <= '1';
    layer1_outputs(5668) <= not(layer0_outputs(4935));
    layer1_outputs(5669) <= layer0_outputs(6469);
    layer1_outputs(5670) <= (layer0_outputs(1243)) and not (layer0_outputs(284));
    layer1_outputs(5671) <= layer0_outputs(2119);
    layer1_outputs(5672) <= not((layer0_outputs(6440)) xor (layer0_outputs(322)));
    layer1_outputs(5673) <= layer0_outputs(3991);
    layer1_outputs(5674) <= (layer0_outputs(889)) and (layer0_outputs(7251));
    layer1_outputs(5675) <= (layer0_outputs(5880)) and not (layer0_outputs(6510));
    layer1_outputs(5676) <= layer0_outputs(2447);
    layer1_outputs(5677) <= (layer0_outputs(1770)) or (layer0_outputs(6660));
    layer1_outputs(5678) <= not(layer0_outputs(2603)) or (layer0_outputs(154));
    layer1_outputs(5679) <= layer0_outputs(7536);
    layer1_outputs(5680) <= not(layer0_outputs(7241)) or (layer0_outputs(5496));
    layer1_outputs(5681) <= (layer0_outputs(3270)) and not (layer0_outputs(3987));
    layer1_outputs(5682) <= not(layer0_outputs(7649));
    layer1_outputs(5683) <= (layer0_outputs(7494)) xor (layer0_outputs(746));
    layer1_outputs(5684) <= not(layer0_outputs(466));
    layer1_outputs(5685) <= '1';
    layer1_outputs(5686) <= '1';
    layer1_outputs(5687) <= (layer0_outputs(712)) or (layer0_outputs(7082));
    layer1_outputs(5688) <= (layer0_outputs(1803)) and not (layer0_outputs(2889));
    layer1_outputs(5689) <= not(layer0_outputs(3287)) or (layer0_outputs(166));
    layer1_outputs(5690) <= '0';
    layer1_outputs(5691) <= not(layer0_outputs(6424)) or (layer0_outputs(4507));
    layer1_outputs(5692) <= layer0_outputs(1111);
    layer1_outputs(5693) <= not(layer0_outputs(1990)) or (layer0_outputs(5457));
    layer1_outputs(5694) <= not(layer0_outputs(6445)) or (layer0_outputs(6148));
    layer1_outputs(5695) <= not(layer0_outputs(4929));
    layer1_outputs(5696) <= layer0_outputs(2046);
    layer1_outputs(5697) <= not(layer0_outputs(2024));
    layer1_outputs(5698) <= not(layer0_outputs(6066)) or (layer0_outputs(2343));
    layer1_outputs(5699) <= layer0_outputs(6114);
    layer1_outputs(5700) <= not((layer0_outputs(817)) and (layer0_outputs(7636)));
    layer1_outputs(5701) <= layer0_outputs(2662);
    layer1_outputs(5702) <= not((layer0_outputs(7183)) xor (layer0_outputs(825)));
    layer1_outputs(5703) <= not(layer0_outputs(6490)) or (layer0_outputs(2789));
    layer1_outputs(5704) <= not((layer0_outputs(5732)) or (layer0_outputs(3013)));
    layer1_outputs(5705) <= not(layer0_outputs(7077));
    layer1_outputs(5706) <= not(layer0_outputs(1675));
    layer1_outputs(5707) <= (layer0_outputs(3437)) or (layer0_outputs(7621));
    layer1_outputs(5708) <= (layer0_outputs(2018)) and not (layer0_outputs(1999));
    layer1_outputs(5709) <= (layer0_outputs(769)) and not (layer0_outputs(6639));
    layer1_outputs(5710) <= not(layer0_outputs(5170));
    layer1_outputs(5711) <= not(layer0_outputs(4637));
    layer1_outputs(5712) <= not(layer0_outputs(5079));
    layer1_outputs(5713) <= not((layer0_outputs(5823)) or (layer0_outputs(5012)));
    layer1_outputs(5714) <= not(layer0_outputs(1222));
    layer1_outputs(5715) <= not((layer0_outputs(2668)) and (layer0_outputs(3222)));
    layer1_outputs(5716) <= not(layer0_outputs(5446));
    layer1_outputs(5717) <= (layer0_outputs(5278)) and not (layer0_outputs(4674));
    layer1_outputs(5718) <= not(layer0_outputs(2898)) or (layer0_outputs(6191));
    layer1_outputs(5719) <= '1';
    layer1_outputs(5720) <= (layer0_outputs(2449)) and (layer0_outputs(5070));
    layer1_outputs(5721) <= not((layer0_outputs(5499)) and (layer0_outputs(6495)));
    layer1_outputs(5722) <= (layer0_outputs(3120)) or (layer0_outputs(2570));
    layer1_outputs(5723) <= (layer0_outputs(6435)) and not (layer0_outputs(2589));
    layer1_outputs(5724) <= '0';
    layer1_outputs(5725) <= (layer0_outputs(1244)) or (layer0_outputs(3936));
    layer1_outputs(5726) <= (layer0_outputs(6200)) and not (layer0_outputs(2372));
    layer1_outputs(5727) <= (layer0_outputs(2156)) and not (layer0_outputs(6422));
    layer1_outputs(5728) <= layer0_outputs(3623);
    layer1_outputs(5729) <= not(layer0_outputs(3018)) or (layer0_outputs(5868));
    layer1_outputs(5730) <= not((layer0_outputs(1055)) xor (layer0_outputs(2833)));
    layer1_outputs(5731) <= not((layer0_outputs(3349)) and (layer0_outputs(5071)));
    layer1_outputs(5732) <= (layer0_outputs(3161)) and not (layer0_outputs(7673));
    layer1_outputs(5733) <= not(layer0_outputs(6311));
    layer1_outputs(5734) <= (layer0_outputs(5888)) and (layer0_outputs(4879));
    layer1_outputs(5735) <= (layer0_outputs(1480)) xor (layer0_outputs(1443));
    layer1_outputs(5736) <= not(layer0_outputs(5928)) or (layer0_outputs(3956));
    layer1_outputs(5737) <= layer0_outputs(4063);
    layer1_outputs(5738) <= (layer0_outputs(1710)) and not (layer0_outputs(6448));
    layer1_outputs(5739) <= not(layer0_outputs(6294));
    layer1_outputs(5740) <= not(layer0_outputs(1034)) or (layer0_outputs(422));
    layer1_outputs(5741) <= not((layer0_outputs(5932)) and (layer0_outputs(6017)));
    layer1_outputs(5742) <= (layer0_outputs(857)) and not (layer0_outputs(6903));
    layer1_outputs(5743) <= layer0_outputs(642);
    layer1_outputs(5744) <= (layer0_outputs(321)) and not (layer0_outputs(6904));
    layer1_outputs(5745) <= (layer0_outputs(5389)) and (layer0_outputs(2740));
    layer1_outputs(5746) <= '1';
    layer1_outputs(5747) <= not(layer0_outputs(5451)) or (layer0_outputs(4109));
    layer1_outputs(5748) <= not(layer0_outputs(4972));
    layer1_outputs(5749) <= '0';
    layer1_outputs(5750) <= not((layer0_outputs(1626)) and (layer0_outputs(7150)));
    layer1_outputs(5751) <= '0';
    layer1_outputs(5752) <= '1';
    layer1_outputs(5753) <= (layer0_outputs(858)) and (layer0_outputs(2840));
    layer1_outputs(5754) <= layer0_outputs(7614);
    layer1_outputs(5755) <= (layer0_outputs(435)) and not (layer0_outputs(2079));
    layer1_outputs(5756) <= not(layer0_outputs(5187));
    layer1_outputs(5757) <= (layer0_outputs(6849)) or (layer0_outputs(6068));
    layer1_outputs(5758) <= layer0_outputs(4038);
    layer1_outputs(5759) <= layer0_outputs(610);
    layer1_outputs(5760) <= not((layer0_outputs(1309)) and (layer0_outputs(7194)));
    layer1_outputs(5761) <= not(layer0_outputs(5906));
    layer1_outputs(5762) <= (layer0_outputs(7544)) xor (layer0_outputs(6177));
    layer1_outputs(5763) <= not((layer0_outputs(696)) xor (layer0_outputs(3028)));
    layer1_outputs(5764) <= not(layer0_outputs(84));
    layer1_outputs(5765) <= (layer0_outputs(7326)) and (layer0_outputs(3791));
    layer1_outputs(5766) <= not(layer0_outputs(3181));
    layer1_outputs(5767) <= not(layer0_outputs(1947)) or (layer0_outputs(1588));
    layer1_outputs(5768) <= layer0_outputs(5966);
    layer1_outputs(5769) <= '0';
    layer1_outputs(5770) <= '0';
    layer1_outputs(5771) <= (layer0_outputs(948)) and not (layer0_outputs(4710));
    layer1_outputs(5772) <= not(layer0_outputs(4962)) or (layer0_outputs(898));
    layer1_outputs(5773) <= (layer0_outputs(917)) and (layer0_outputs(555));
    layer1_outputs(5774) <= (layer0_outputs(6028)) and (layer0_outputs(4328));
    layer1_outputs(5775) <= (layer0_outputs(5972)) and not (layer0_outputs(1309));
    layer1_outputs(5776) <= '0';
    layer1_outputs(5777) <= not(layer0_outputs(424)) or (layer0_outputs(6723));
    layer1_outputs(5778) <= (layer0_outputs(1991)) and (layer0_outputs(697));
    layer1_outputs(5779) <= not((layer0_outputs(5526)) or (layer0_outputs(7143)));
    layer1_outputs(5780) <= not(layer0_outputs(1011)) or (layer0_outputs(1934));
    layer1_outputs(5781) <= (layer0_outputs(7540)) and (layer0_outputs(6014));
    layer1_outputs(5782) <= not(layer0_outputs(2604));
    layer1_outputs(5783) <= (layer0_outputs(2623)) and (layer0_outputs(1389));
    layer1_outputs(5784) <= not((layer0_outputs(3106)) and (layer0_outputs(3992)));
    layer1_outputs(5785) <= '1';
    layer1_outputs(5786) <= (layer0_outputs(4235)) and not (layer0_outputs(2700));
    layer1_outputs(5787) <= not(layer0_outputs(3363));
    layer1_outputs(5788) <= not(layer0_outputs(2481));
    layer1_outputs(5789) <= not(layer0_outputs(2115));
    layer1_outputs(5790) <= not((layer0_outputs(2551)) xor (layer0_outputs(6020)));
    layer1_outputs(5791) <= (layer0_outputs(5883)) or (layer0_outputs(4779));
    layer1_outputs(5792) <= (layer0_outputs(641)) or (layer0_outputs(6431));
    layer1_outputs(5793) <= not((layer0_outputs(2309)) xor (layer0_outputs(4169)));
    layer1_outputs(5794) <= layer0_outputs(1102);
    layer1_outputs(5795) <= not(layer0_outputs(2302)) or (layer0_outputs(5198));
    layer1_outputs(5796) <= layer0_outputs(2746);
    layer1_outputs(5797) <= not((layer0_outputs(3022)) and (layer0_outputs(404)));
    layer1_outputs(5798) <= (layer0_outputs(4664)) or (layer0_outputs(76));
    layer1_outputs(5799) <= layer0_outputs(2610);
    layer1_outputs(5800) <= (layer0_outputs(4684)) or (layer0_outputs(6270));
    layer1_outputs(5801) <= (layer0_outputs(4391)) and (layer0_outputs(3155));
    layer1_outputs(5802) <= '0';
    layer1_outputs(5803) <= not(layer0_outputs(95)) or (layer0_outputs(1932));
    layer1_outputs(5804) <= '0';
    layer1_outputs(5805) <= not((layer0_outputs(1976)) xor (layer0_outputs(6022)));
    layer1_outputs(5806) <= (layer0_outputs(747)) and (layer0_outputs(2993));
    layer1_outputs(5807) <= layer0_outputs(6376);
    layer1_outputs(5808) <= '0';
    layer1_outputs(5809) <= not((layer0_outputs(4972)) and (layer0_outputs(1185)));
    layer1_outputs(5810) <= layer0_outputs(6957);
    layer1_outputs(5811) <= not(layer0_outputs(4009)) or (layer0_outputs(1341));
    layer1_outputs(5812) <= layer0_outputs(1918);
    layer1_outputs(5813) <= layer0_outputs(2169);
    layer1_outputs(5814) <= not(layer0_outputs(4636));
    layer1_outputs(5815) <= not(layer0_outputs(3557)) or (layer0_outputs(216));
    layer1_outputs(5816) <= layer0_outputs(2549);
    layer1_outputs(5817) <= not(layer0_outputs(5724)) or (layer0_outputs(5706));
    layer1_outputs(5818) <= (layer0_outputs(3510)) and (layer0_outputs(6846));
    layer1_outputs(5819) <= layer0_outputs(136);
    layer1_outputs(5820) <= '1';
    layer1_outputs(5821) <= (layer0_outputs(6166)) and not (layer0_outputs(1587));
    layer1_outputs(5822) <= not(layer0_outputs(5319)) or (layer0_outputs(6768));
    layer1_outputs(5823) <= not((layer0_outputs(2717)) and (layer0_outputs(1867)));
    layer1_outputs(5824) <= layer0_outputs(3111);
    layer1_outputs(5825) <= '1';
    layer1_outputs(5826) <= not((layer0_outputs(122)) and (layer0_outputs(1232)));
    layer1_outputs(5827) <= (layer0_outputs(2977)) and not (layer0_outputs(1614));
    layer1_outputs(5828) <= (layer0_outputs(236)) and not (layer0_outputs(1938));
    layer1_outputs(5829) <= (layer0_outputs(1407)) or (layer0_outputs(2174));
    layer1_outputs(5830) <= '0';
    layer1_outputs(5831) <= (layer0_outputs(7100)) and (layer0_outputs(7137));
    layer1_outputs(5832) <= not(layer0_outputs(1782));
    layer1_outputs(5833) <= (layer0_outputs(2583)) xor (layer0_outputs(6319));
    layer1_outputs(5834) <= not((layer0_outputs(1880)) and (layer0_outputs(4774)));
    layer1_outputs(5835) <= not(layer0_outputs(7408)) or (layer0_outputs(2583));
    layer1_outputs(5836) <= '1';
    layer1_outputs(5837) <= layer0_outputs(2199);
    layer1_outputs(5838) <= not(layer0_outputs(7400));
    layer1_outputs(5839) <= (layer0_outputs(7388)) or (layer0_outputs(283));
    layer1_outputs(5840) <= not(layer0_outputs(3126));
    layer1_outputs(5841) <= (layer0_outputs(3935)) and not (layer0_outputs(7193));
    layer1_outputs(5842) <= not(layer0_outputs(4192));
    layer1_outputs(5843) <= (layer0_outputs(2098)) or (layer0_outputs(5410));
    layer1_outputs(5844) <= layer0_outputs(304);
    layer1_outputs(5845) <= not((layer0_outputs(7384)) and (layer0_outputs(5769)));
    layer1_outputs(5846) <= layer0_outputs(457);
    layer1_outputs(5847) <= (layer0_outputs(4469)) and (layer0_outputs(5526));
    layer1_outputs(5848) <= not(layer0_outputs(6124));
    layer1_outputs(5849) <= not(layer0_outputs(3787)) or (layer0_outputs(2272));
    layer1_outputs(5850) <= (layer0_outputs(2009)) xor (layer0_outputs(3182));
    layer1_outputs(5851) <= not((layer0_outputs(6711)) xor (layer0_outputs(4184)));
    layer1_outputs(5852) <= (layer0_outputs(6896)) and (layer0_outputs(2979));
    layer1_outputs(5853) <= not((layer0_outputs(1819)) or (layer0_outputs(3673)));
    layer1_outputs(5854) <= layer0_outputs(2391);
    layer1_outputs(5855) <= (layer0_outputs(3292)) or (layer0_outputs(1703));
    layer1_outputs(5856) <= not(layer0_outputs(1555)) or (layer0_outputs(2735));
    layer1_outputs(5857) <= not(layer0_outputs(7259)) or (layer0_outputs(1824));
    layer1_outputs(5858) <= not(layer0_outputs(6191)) or (layer0_outputs(6118));
    layer1_outputs(5859) <= layer0_outputs(471);
    layer1_outputs(5860) <= not(layer0_outputs(2416)) or (layer0_outputs(3237));
    layer1_outputs(5861) <= (layer0_outputs(7543)) and not (layer0_outputs(7325));
    layer1_outputs(5862) <= layer0_outputs(7638);
    layer1_outputs(5863) <= (layer0_outputs(7223)) or (layer0_outputs(3813));
    layer1_outputs(5864) <= layer0_outputs(97);
    layer1_outputs(5865) <= not(layer0_outputs(3559));
    layer1_outputs(5866) <= not(layer0_outputs(4459));
    layer1_outputs(5867) <= not(layer0_outputs(6716));
    layer1_outputs(5868) <= not((layer0_outputs(948)) or (layer0_outputs(7085)));
    layer1_outputs(5869) <= not((layer0_outputs(7132)) or (layer0_outputs(1925)));
    layer1_outputs(5870) <= layer0_outputs(2823);
    layer1_outputs(5871) <= layer0_outputs(6498);
    layer1_outputs(5872) <= '1';
    layer1_outputs(5873) <= (layer0_outputs(5229)) xor (layer0_outputs(374));
    layer1_outputs(5874) <= not(layer0_outputs(3877));
    layer1_outputs(5875) <= '0';
    layer1_outputs(5876) <= '1';
    layer1_outputs(5877) <= '0';
    layer1_outputs(5878) <= not((layer0_outputs(3549)) and (layer0_outputs(3502)));
    layer1_outputs(5879) <= not(layer0_outputs(7543)) or (layer0_outputs(7498));
    layer1_outputs(5880) <= not((layer0_outputs(6184)) and (layer0_outputs(6665)));
    layer1_outputs(5881) <= '1';
    layer1_outputs(5882) <= (layer0_outputs(6399)) and not (layer0_outputs(3009));
    layer1_outputs(5883) <= not(layer0_outputs(3435)) or (layer0_outputs(2477));
    layer1_outputs(5884) <= '1';
    layer1_outputs(5885) <= '1';
    layer1_outputs(5886) <= layer0_outputs(1142);
    layer1_outputs(5887) <= layer0_outputs(1203);
    layer1_outputs(5888) <= not((layer0_outputs(3220)) or (layer0_outputs(1886)));
    layer1_outputs(5889) <= not(layer0_outputs(1898));
    layer1_outputs(5890) <= layer0_outputs(6371);
    layer1_outputs(5891) <= layer0_outputs(3542);
    layer1_outputs(5892) <= (layer0_outputs(1767)) xor (layer0_outputs(310));
    layer1_outputs(5893) <= layer0_outputs(6586);
    layer1_outputs(5894) <= not(layer0_outputs(2146)) or (layer0_outputs(4736));
    layer1_outputs(5895) <= not(layer0_outputs(3473));
    layer1_outputs(5896) <= not((layer0_outputs(7271)) xor (layer0_outputs(761)));
    layer1_outputs(5897) <= (layer0_outputs(3765)) or (layer0_outputs(1394));
    layer1_outputs(5898) <= not((layer0_outputs(4586)) and (layer0_outputs(6836)));
    layer1_outputs(5899) <= not((layer0_outputs(4073)) and (layer0_outputs(2490)));
    layer1_outputs(5900) <= (layer0_outputs(4360)) and not (layer0_outputs(4872));
    layer1_outputs(5901) <= (layer0_outputs(3057)) and not (layer0_outputs(40));
    layer1_outputs(5902) <= layer0_outputs(1154);
    layer1_outputs(5903) <= not((layer0_outputs(4484)) xor (layer0_outputs(3254)));
    layer1_outputs(5904) <= not(layer0_outputs(4432)) or (layer0_outputs(439));
    layer1_outputs(5905) <= (layer0_outputs(3879)) xor (layer0_outputs(2191));
    layer1_outputs(5906) <= not(layer0_outputs(4181)) or (layer0_outputs(6572));
    layer1_outputs(5907) <= not((layer0_outputs(3607)) or (layer0_outputs(1323)));
    layer1_outputs(5908) <= not(layer0_outputs(7542));
    layer1_outputs(5909) <= layer0_outputs(1926);
    layer1_outputs(5910) <= not((layer0_outputs(3755)) and (layer0_outputs(7121)));
    layer1_outputs(5911) <= (layer0_outputs(3738)) and not (layer0_outputs(6952));
    layer1_outputs(5912) <= (layer0_outputs(7584)) and not (layer0_outputs(6011));
    layer1_outputs(5913) <= '0';
    layer1_outputs(5914) <= not((layer0_outputs(3348)) or (layer0_outputs(6660)));
    layer1_outputs(5915) <= layer0_outputs(273);
    layer1_outputs(5916) <= layer0_outputs(6789);
    layer1_outputs(5917) <= '1';
    layer1_outputs(5918) <= not((layer0_outputs(6783)) or (layer0_outputs(100)));
    layer1_outputs(5919) <= not((layer0_outputs(4178)) and (layer0_outputs(2007)));
    layer1_outputs(5920) <= '0';
    layer1_outputs(5921) <= not(layer0_outputs(6346)) or (layer0_outputs(4092));
    layer1_outputs(5922) <= (layer0_outputs(4709)) and not (layer0_outputs(1973));
    layer1_outputs(5923) <= layer0_outputs(3582);
    layer1_outputs(5924) <= '1';
    layer1_outputs(5925) <= not((layer0_outputs(2425)) xor (layer0_outputs(5618)));
    layer1_outputs(5926) <= (layer0_outputs(5593)) and not (layer0_outputs(1659));
    layer1_outputs(5927) <= layer0_outputs(6517);
    layer1_outputs(5928) <= not(layer0_outputs(820));
    layer1_outputs(5929) <= '1';
    layer1_outputs(5930) <= '1';
    layer1_outputs(5931) <= '1';
    layer1_outputs(5932) <= not((layer0_outputs(448)) and (layer0_outputs(472)));
    layer1_outputs(5933) <= not((layer0_outputs(5886)) or (layer0_outputs(2474)));
    layer1_outputs(5934) <= not((layer0_outputs(805)) and (layer0_outputs(5625)));
    layer1_outputs(5935) <= (layer0_outputs(5191)) and (layer0_outputs(4831));
    layer1_outputs(5936) <= not(layer0_outputs(7122));
    layer1_outputs(5937) <= not((layer0_outputs(659)) and (layer0_outputs(6685)));
    layer1_outputs(5938) <= not(layer0_outputs(4419)) or (layer0_outputs(6412));
    layer1_outputs(5939) <= not(layer0_outputs(7071));
    layer1_outputs(5940) <= not((layer0_outputs(1491)) or (layer0_outputs(5377)));
    layer1_outputs(5941) <= not(layer0_outputs(4028)) or (layer0_outputs(2336));
    layer1_outputs(5942) <= not(layer0_outputs(5353));
    layer1_outputs(5943) <= (layer0_outputs(4251)) or (layer0_outputs(6513));
    layer1_outputs(5944) <= not(layer0_outputs(3567)) or (layer0_outputs(3647));
    layer1_outputs(5945) <= not(layer0_outputs(2734)) or (layer0_outputs(5352));
    layer1_outputs(5946) <= not(layer0_outputs(6338));
    layer1_outputs(5947) <= '1';
    layer1_outputs(5948) <= (layer0_outputs(3915)) and not (layer0_outputs(3607));
    layer1_outputs(5949) <= (layer0_outputs(5638)) xor (layer0_outputs(1083));
    layer1_outputs(5950) <= not(layer0_outputs(5097));
    layer1_outputs(5951) <= (layer0_outputs(3993)) and not (layer0_outputs(1478));
    layer1_outputs(5952) <= not(layer0_outputs(3642));
    layer1_outputs(5953) <= (layer0_outputs(3659)) and not (layer0_outputs(3566));
    layer1_outputs(5954) <= (layer0_outputs(3090)) and not (layer0_outputs(6084));
    layer1_outputs(5955) <= not(layer0_outputs(6748)) or (layer0_outputs(4645));
    layer1_outputs(5956) <= (layer0_outputs(4492)) xor (layer0_outputs(5279));
    layer1_outputs(5957) <= not(layer0_outputs(3176)) or (layer0_outputs(6772));
    layer1_outputs(5958) <= not(layer0_outputs(2347)) or (layer0_outputs(1125));
    layer1_outputs(5959) <= layer0_outputs(6404);
    layer1_outputs(5960) <= '1';
    layer1_outputs(5961) <= layer0_outputs(2721);
    layer1_outputs(5962) <= (layer0_outputs(2439)) and not (layer0_outputs(2246));
    layer1_outputs(5963) <= layer0_outputs(2040);
    layer1_outputs(5964) <= not((layer0_outputs(1349)) and (layer0_outputs(5994)));
    layer1_outputs(5965) <= layer0_outputs(4887);
    layer1_outputs(5966) <= not(layer0_outputs(7447)) or (layer0_outputs(7548));
    layer1_outputs(5967) <= layer0_outputs(5350);
    layer1_outputs(5968) <= not(layer0_outputs(1969));
    layer1_outputs(5969) <= (layer0_outputs(3026)) and not (layer0_outputs(2604));
    layer1_outputs(5970) <= (layer0_outputs(315)) and not (layer0_outputs(4925));
    layer1_outputs(5971) <= (layer0_outputs(3433)) and (layer0_outputs(6941));
    layer1_outputs(5972) <= not(layer0_outputs(2858)) or (layer0_outputs(1318));
    layer1_outputs(5973) <= (layer0_outputs(2862)) and not (layer0_outputs(785));
    layer1_outputs(5974) <= layer0_outputs(5057);
    layer1_outputs(5975) <= (layer0_outputs(200)) xor (layer0_outputs(5058));
    layer1_outputs(5976) <= layer0_outputs(33);
    layer1_outputs(5977) <= not(layer0_outputs(5353)) or (layer0_outputs(825));
    layer1_outputs(5978) <= not(layer0_outputs(47));
    layer1_outputs(5979) <= layer0_outputs(3503);
    layer1_outputs(5980) <= layer0_outputs(3889);
    layer1_outputs(5981) <= layer0_outputs(530);
    layer1_outputs(5982) <= not(layer0_outputs(618));
    layer1_outputs(5983) <= layer0_outputs(3935);
    layer1_outputs(5984) <= (layer0_outputs(4667)) and not (layer0_outputs(731));
    layer1_outputs(5985) <= not(layer0_outputs(5031)) or (layer0_outputs(7292));
    layer1_outputs(5986) <= '0';
    layer1_outputs(5987) <= not((layer0_outputs(7211)) and (layer0_outputs(5027)));
    layer1_outputs(5988) <= not((layer0_outputs(6451)) and (layer0_outputs(6099)));
    layer1_outputs(5989) <= layer0_outputs(7586);
    layer1_outputs(5990) <= (layer0_outputs(5394)) and (layer0_outputs(254));
    layer1_outputs(5991) <= not((layer0_outputs(29)) and (layer0_outputs(6429)));
    layer1_outputs(5992) <= (layer0_outputs(589)) and (layer0_outputs(5235));
    layer1_outputs(5993) <= (layer0_outputs(6484)) and not (layer0_outputs(6374));
    layer1_outputs(5994) <= layer0_outputs(5822);
    layer1_outputs(5995) <= not((layer0_outputs(1817)) and (layer0_outputs(5810)));
    layer1_outputs(5996) <= '1';
    layer1_outputs(5997) <= (layer0_outputs(5656)) and not (layer0_outputs(5464));
    layer1_outputs(5998) <= (layer0_outputs(1263)) and not (layer0_outputs(1549));
    layer1_outputs(5999) <= (layer0_outputs(5959)) or (layer0_outputs(4102));
    layer1_outputs(6000) <= (layer0_outputs(3764)) xor (layer0_outputs(4384));
    layer1_outputs(6001) <= (layer0_outputs(2453)) and not (layer0_outputs(3069));
    layer1_outputs(6002) <= not((layer0_outputs(1650)) or (layer0_outputs(2892)));
    layer1_outputs(6003) <= not((layer0_outputs(1761)) or (layer0_outputs(3359)));
    layer1_outputs(6004) <= not(layer0_outputs(3516));
    layer1_outputs(6005) <= (layer0_outputs(6414)) and (layer0_outputs(2290));
    layer1_outputs(6006) <= layer0_outputs(2809);
    layer1_outputs(6007) <= '0';
    layer1_outputs(6008) <= layer0_outputs(1282);
    layer1_outputs(6009) <= (layer0_outputs(3383)) xor (layer0_outputs(5475));
    layer1_outputs(6010) <= not((layer0_outputs(3771)) or (layer0_outputs(7243)));
    layer1_outputs(6011) <= not(layer0_outputs(3900));
    layer1_outputs(6012) <= not(layer0_outputs(5194));
    layer1_outputs(6013) <= (layer0_outputs(1253)) and not (layer0_outputs(4682));
    layer1_outputs(6014) <= layer0_outputs(7400);
    layer1_outputs(6015) <= not((layer0_outputs(5589)) or (layer0_outputs(1254)));
    layer1_outputs(6016) <= layer0_outputs(7405);
    layer1_outputs(6017) <= not(layer0_outputs(3921));
    layer1_outputs(6018) <= not(layer0_outputs(3669)) or (layer0_outputs(7205));
    layer1_outputs(6019) <= '1';
    layer1_outputs(6020) <= (layer0_outputs(6405)) and not (layer0_outputs(1048));
    layer1_outputs(6021) <= layer0_outputs(3905);
    layer1_outputs(6022) <= layer0_outputs(7539);
    layer1_outputs(6023) <= not(layer0_outputs(5770));
    layer1_outputs(6024) <= (layer0_outputs(2060)) and not (layer0_outputs(4422));
    layer1_outputs(6025) <= (layer0_outputs(4457)) or (layer0_outputs(5800));
    layer1_outputs(6026) <= not((layer0_outputs(6171)) or (layer0_outputs(1703)));
    layer1_outputs(6027) <= not(layer0_outputs(4717)) or (layer0_outputs(3712));
    layer1_outputs(6028) <= (layer0_outputs(2716)) and not (layer0_outputs(652));
    layer1_outputs(6029) <= (layer0_outputs(700)) and not (layer0_outputs(7657));
    layer1_outputs(6030) <= layer0_outputs(4861);
    layer1_outputs(6031) <= '0';
    layer1_outputs(6032) <= '1';
    layer1_outputs(6033) <= (layer0_outputs(4415)) and not (layer0_outputs(961));
    layer1_outputs(6034) <= not(layer0_outputs(7627));
    layer1_outputs(6035) <= not(layer0_outputs(5776)) or (layer0_outputs(2316));
    layer1_outputs(6036) <= layer0_outputs(7339);
    layer1_outputs(6037) <= not(layer0_outputs(1123));
    layer1_outputs(6038) <= not(layer0_outputs(5724));
    layer1_outputs(6039) <= layer0_outputs(4501);
    layer1_outputs(6040) <= not((layer0_outputs(6030)) and (layer0_outputs(4835)));
    layer1_outputs(6041) <= layer0_outputs(3856);
    layer1_outputs(6042) <= not(layer0_outputs(1521));
    layer1_outputs(6043) <= not(layer0_outputs(278));
    layer1_outputs(6044) <= layer0_outputs(3437);
    layer1_outputs(6045) <= not(layer0_outputs(6454));
    layer1_outputs(6046) <= '1';
    layer1_outputs(6047) <= layer0_outputs(2386);
    layer1_outputs(6048) <= (layer0_outputs(5340)) and not (layer0_outputs(959));
    layer1_outputs(6049) <= (layer0_outputs(2043)) and not (layer0_outputs(1700));
    layer1_outputs(6050) <= not(layer0_outputs(667));
    layer1_outputs(6051) <= layer0_outputs(1501);
    layer1_outputs(6052) <= not((layer0_outputs(3106)) and (layer0_outputs(5709)));
    layer1_outputs(6053) <= layer0_outputs(3419);
    layer1_outputs(6054) <= (layer0_outputs(3750)) or (layer0_outputs(443));
    layer1_outputs(6055) <= not(layer0_outputs(2112)) or (layer0_outputs(3116));
    layer1_outputs(6056) <= (layer0_outputs(2533)) and not (layer0_outputs(1783));
    layer1_outputs(6057) <= not(layer0_outputs(4637));
    layer1_outputs(6058) <= not((layer0_outputs(4040)) or (layer0_outputs(6478)));
    layer1_outputs(6059) <= not(layer0_outputs(3654));
    layer1_outputs(6060) <= (layer0_outputs(6641)) xor (layer0_outputs(2614));
    layer1_outputs(6061) <= not(layer0_outputs(4730)) or (layer0_outputs(4476));
    layer1_outputs(6062) <= not(layer0_outputs(3954)) or (layer0_outputs(6721));
    layer1_outputs(6063) <= not((layer0_outputs(3201)) and (layer0_outputs(548)));
    layer1_outputs(6064) <= not(layer0_outputs(3386)) or (layer0_outputs(2385));
    layer1_outputs(6065) <= not(layer0_outputs(2295));
    layer1_outputs(6066) <= layer0_outputs(3946);
    layer1_outputs(6067) <= not((layer0_outputs(1221)) and (layer0_outputs(6186)));
    layer1_outputs(6068) <= not((layer0_outputs(5134)) and (layer0_outputs(2858)));
    layer1_outputs(6069) <= not(layer0_outputs(6527));
    layer1_outputs(6070) <= '0';
    layer1_outputs(6071) <= layer0_outputs(2863);
    layer1_outputs(6072) <= layer0_outputs(299);
    layer1_outputs(6073) <= not(layer0_outputs(4033));
    layer1_outputs(6074) <= not(layer0_outputs(5712)) or (layer0_outputs(3186));
    layer1_outputs(6075) <= layer0_outputs(3188);
    layer1_outputs(6076) <= (layer0_outputs(4491)) and not (layer0_outputs(2240));
    layer1_outputs(6077) <= not(layer0_outputs(7264));
    layer1_outputs(6078) <= not(layer0_outputs(5723));
    layer1_outputs(6079) <= (layer0_outputs(4185)) or (layer0_outputs(4190));
    layer1_outputs(6080) <= not((layer0_outputs(3823)) and (layer0_outputs(1461)));
    layer1_outputs(6081) <= layer0_outputs(4921);
    layer1_outputs(6082) <= not(layer0_outputs(520));
    layer1_outputs(6083) <= layer0_outputs(2329);
    layer1_outputs(6084) <= layer0_outputs(7450);
    layer1_outputs(6085) <= '0';
    layer1_outputs(6086) <= not(layer0_outputs(804));
    layer1_outputs(6087) <= not((layer0_outputs(2212)) or (layer0_outputs(3290)));
    layer1_outputs(6088) <= (layer0_outputs(1865)) and not (layer0_outputs(2957));
    layer1_outputs(6089) <= (layer0_outputs(4834)) or (layer0_outputs(4993));
    layer1_outputs(6090) <= (layer0_outputs(4772)) and not (layer0_outputs(1598));
    layer1_outputs(6091) <= not(layer0_outputs(1375)) or (layer0_outputs(73));
    layer1_outputs(6092) <= (layer0_outputs(1699)) and not (layer0_outputs(1920));
    layer1_outputs(6093) <= '0';
    layer1_outputs(6094) <= '1';
    layer1_outputs(6095) <= not(layer0_outputs(5047));
    layer1_outputs(6096) <= layer0_outputs(2039);
    layer1_outputs(6097) <= layer0_outputs(1568);
    layer1_outputs(6098) <= not((layer0_outputs(5519)) and (layer0_outputs(6901)));
    layer1_outputs(6099) <= layer0_outputs(3279);
    layer1_outputs(6100) <= (layer0_outputs(6671)) and not (layer0_outputs(389));
    layer1_outputs(6101) <= not(layer0_outputs(5524)) or (layer0_outputs(2314));
    layer1_outputs(6102) <= (layer0_outputs(3092)) and not (layer0_outputs(6743));
    layer1_outputs(6103) <= (layer0_outputs(1688)) and not (layer0_outputs(5960));
    layer1_outputs(6104) <= not(layer0_outputs(3242));
    layer1_outputs(6105) <= (layer0_outputs(3028)) or (layer0_outputs(5929));
    layer1_outputs(6106) <= not(layer0_outputs(2214));
    layer1_outputs(6107) <= not(layer0_outputs(4394)) or (layer0_outputs(748));
    layer1_outputs(6108) <= not(layer0_outputs(5331));
    layer1_outputs(6109) <= layer0_outputs(510);
    layer1_outputs(6110) <= (layer0_outputs(448)) and not (layer0_outputs(532));
    layer1_outputs(6111) <= layer0_outputs(1376);
    layer1_outputs(6112) <= not(layer0_outputs(6937));
    layer1_outputs(6113) <= (layer0_outputs(4543)) xor (layer0_outputs(7587));
    layer1_outputs(6114) <= '0';
    layer1_outputs(6115) <= '1';
    layer1_outputs(6116) <= not(layer0_outputs(6247));
    layer1_outputs(6117) <= not(layer0_outputs(4720)) or (layer0_outputs(7524));
    layer1_outputs(6118) <= (layer0_outputs(1618)) and not (layer0_outputs(5936));
    layer1_outputs(6119) <= not((layer0_outputs(4580)) and (layer0_outputs(2187)));
    layer1_outputs(6120) <= '1';
    layer1_outputs(6121) <= not(layer0_outputs(941)) or (layer0_outputs(6801));
    layer1_outputs(6122) <= not(layer0_outputs(16));
    layer1_outputs(6123) <= not((layer0_outputs(6312)) or (layer0_outputs(6107)));
    layer1_outputs(6124) <= layer0_outputs(4513);
    layer1_outputs(6125) <= (layer0_outputs(593)) and not (layer0_outputs(5337));
    layer1_outputs(6126) <= not(layer0_outputs(2928)) or (layer0_outputs(4957));
    layer1_outputs(6127) <= layer0_outputs(2357);
    layer1_outputs(6128) <= not((layer0_outputs(7455)) or (layer0_outputs(439)));
    layer1_outputs(6129) <= not(layer0_outputs(4877));
    layer1_outputs(6130) <= (layer0_outputs(1013)) and not (layer0_outputs(5653));
    layer1_outputs(6131) <= not(layer0_outputs(1401));
    layer1_outputs(6132) <= '1';
    layer1_outputs(6133) <= (layer0_outputs(3012)) or (layer0_outputs(6726));
    layer1_outputs(6134) <= not((layer0_outputs(6926)) and (layer0_outputs(5566)));
    layer1_outputs(6135) <= '1';
    layer1_outputs(6136) <= (layer0_outputs(1148)) and not (layer0_outputs(6994));
    layer1_outputs(6137) <= not((layer0_outputs(2863)) or (layer0_outputs(587)));
    layer1_outputs(6138) <= (layer0_outputs(2805)) and not (layer0_outputs(2768));
    layer1_outputs(6139) <= (layer0_outputs(1996)) or (layer0_outputs(3056));
    layer1_outputs(6140) <= (layer0_outputs(706)) and not (layer0_outputs(865));
    layer1_outputs(6141) <= (layer0_outputs(6764)) and not (layer0_outputs(7617));
    layer1_outputs(6142) <= (layer0_outputs(4338)) and not (layer0_outputs(3023));
    layer1_outputs(6143) <= not(layer0_outputs(5002)) or (layer0_outputs(5558));
    layer1_outputs(6144) <= layer0_outputs(4489);
    layer1_outputs(6145) <= layer0_outputs(5814);
    layer1_outputs(6146) <= not(layer0_outputs(957));
    layer1_outputs(6147) <= layer0_outputs(2465);
    layer1_outputs(6148) <= layer0_outputs(2762);
    layer1_outputs(6149) <= layer0_outputs(1264);
    layer1_outputs(6150) <= not((layer0_outputs(5190)) and (layer0_outputs(6292)));
    layer1_outputs(6151) <= '1';
    layer1_outputs(6152) <= (layer0_outputs(6254)) and not (layer0_outputs(4096));
    layer1_outputs(6153) <= layer0_outputs(96);
    layer1_outputs(6154) <= layer0_outputs(6696);
    layer1_outputs(6155) <= (layer0_outputs(6504)) and not (layer0_outputs(7450));
    layer1_outputs(6156) <= layer0_outputs(3767);
    layer1_outputs(6157) <= not(layer0_outputs(382)) or (layer0_outputs(3037));
    layer1_outputs(6158) <= (layer0_outputs(6492)) xor (layer0_outputs(5878));
    layer1_outputs(6159) <= (layer0_outputs(3800)) xor (layer0_outputs(290));
    layer1_outputs(6160) <= not(layer0_outputs(931));
    layer1_outputs(6161) <= not((layer0_outputs(6731)) xor (layer0_outputs(5434)));
    layer1_outputs(6162) <= not((layer0_outputs(6468)) and (layer0_outputs(3980)));
    layer1_outputs(6163) <= (layer0_outputs(5523)) and not (layer0_outputs(2700));
    layer1_outputs(6164) <= not((layer0_outputs(5757)) or (layer0_outputs(6668)));
    layer1_outputs(6165) <= not(layer0_outputs(527));
    layer1_outputs(6166) <= not((layer0_outputs(2255)) or (layer0_outputs(1417)));
    layer1_outputs(6167) <= layer0_outputs(1722);
    layer1_outputs(6168) <= not(layer0_outputs(5866)) or (layer0_outputs(3808));
    layer1_outputs(6169) <= layer0_outputs(5680);
    layer1_outputs(6170) <= not(layer0_outputs(2673));
    layer1_outputs(6171) <= not(layer0_outputs(2718));
    layer1_outputs(6172) <= not(layer0_outputs(288)) or (layer0_outputs(1481));
    layer1_outputs(6173) <= (layer0_outputs(5472)) and not (layer0_outputs(2518));
    layer1_outputs(6174) <= '0';
    layer1_outputs(6175) <= not(layer0_outputs(941));
    layer1_outputs(6176) <= layer0_outputs(3113);
    layer1_outputs(6177) <= '0';
    layer1_outputs(6178) <= not(layer0_outputs(6274));
    layer1_outputs(6179) <= not(layer0_outputs(6231)) or (layer0_outputs(4306));
    layer1_outputs(6180) <= not((layer0_outputs(1070)) xor (layer0_outputs(4023)));
    layer1_outputs(6181) <= not((layer0_outputs(7374)) or (layer0_outputs(272)));
    layer1_outputs(6182) <= not(layer0_outputs(2419));
    layer1_outputs(6183) <= (layer0_outputs(1644)) xor (layer0_outputs(2782));
    layer1_outputs(6184) <= not((layer0_outputs(5538)) xor (layer0_outputs(942)));
    layer1_outputs(6185) <= layer0_outputs(2462);
    layer1_outputs(6186) <= layer0_outputs(4033);
    layer1_outputs(6187) <= not((layer0_outputs(480)) and (layer0_outputs(6011)));
    layer1_outputs(6188) <= (layer0_outputs(5578)) or (layer0_outputs(4239));
    layer1_outputs(6189) <= '0';
    layer1_outputs(6190) <= not((layer0_outputs(217)) or (layer0_outputs(204)));
    layer1_outputs(6191) <= layer0_outputs(3381);
    layer1_outputs(6192) <= not(layer0_outputs(1987));
    layer1_outputs(6193) <= not((layer0_outputs(578)) and (layer0_outputs(3648)));
    layer1_outputs(6194) <= not(layer0_outputs(7456)) or (layer0_outputs(3435));
    layer1_outputs(6195) <= (layer0_outputs(4504)) and not (layer0_outputs(2243));
    layer1_outputs(6196) <= not(layer0_outputs(3320)) or (layer0_outputs(1813));
    layer1_outputs(6197) <= not((layer0_outputs(639)) and (layer0_outputs(6473)));
    layer1_outputs(6198) <= not((layer0_outputs(3123)) and (layer0_outputs(3371)));
    layer1_outputs(6199) <= not(layer0_outputs(4929));
    layer1_outputs(6200) <= not((layer0_outputs(5798)) and (layer0_outputs(4725)));
    layer1_outputs(6201) <= '1';
    layer1_outputs(6202) <= (layer0_outputs(6568)) xor (layer0_outputs(7328));
    layer1_outputs(6203) <= not((layer0_outputs(7439)) and (layer0_outputs(6276)));
    layer1_outputs(6204) <= not(layer0_outputs(6428)) or (layer0_outputs(3863));
    layer1_outputs(6205) <= not(layer0_outputs(3273));
    layer1_outputs(6206) <= '1';
    layer1_outputs(6207) <= not((layer0_outputs(3746)) and (layer0_outputs(1967)));
    layer1_outputs(6208) <= layer0_outputs(4348);
    layer1_outputs(6209) <= layer0_outputs(7007);
    layer1_outputs(6210) <= (layer0_outputs(6512)) and not (layer0_outputs(3752));
    layer1_outputs(6211) <= '1';
    layer1_outputs(6212) <= layer0_outputs(7425);
    layer1_outputs(6213) <= layer0_outputs(2622);
    layer1_outputs(6214) <= not(layer0_outputs(3697)) or (layer0_outputs(4025));
    layer1_outputs(6215) <= (layer0_outputs(2513)) and not (layer0_outputs(2976));
    layer1_outputs(6216) <= (layer0_outputs(5040)) xor (layer0_outputs(323));
    layer1_outputs(6217) <= not(layer0_outputs(6390));
    layer1_outputs(6218) <= not(layer0_outputs(3744)) or (layer0_outputs(3942));
    layer1_outputs(6219) <= layer0_outputs(5024);
    layer1_outputs(6220) <= layer0_outputs(6118);
    layer1_outputs(6221) <= (layer0_outputs(4328)) and not (layer0_outputs(5431));
    layer1_outputs(6222) <= not(layer0_outputs(2917)) or (layer0_outputs(7316));
    layer1_outputs(6223) <= '1';
    layer1_outputs(6224) <= layer0_outputs(5280);
    layer1_outputs(6225) <= not(layer0_outputs(2086));
    layer1_outputs(6226) <= layer0_outputs(124);
    layer1_outputs(6227) <= layer0_outputs(6325);
    layer1_outputs(6228) <= not(layer0_outputs(3141));
    layer1_outputs(6229) <= not(layer0_outputs(3930));
    layer1_outputs(6230) <= layer0_outputs(1860);
    layer1_outputs(6231) <= not((layer0_outputs(4991)) and (layer0_outputs(7355)));
    layer1_outputs(6232) <= not((layer0_outputs(2270)) and (layer0_outputs(2362)));
    layer1_outputs(6233) <= '1';
    layer1_outputs(6234) <= (layer0_outputs(1370)) or (layer0_outputs(6409));
    layer1_outputs(6235) <= not(layer0_outputs(6180));
    layer1_outputs(6236) <= not((layer0_outputs(7161)) and (layer0_outputs(7454)));
    layer1_outputs(6237) <= '1';
    layer1_outputs(6238) <= layer0_outputs(6863);
    layer1_outputs(6239) <= not(layer0_outputs(735)) or (layer0_outputs(5469));
    layer1_outputs(6240) <= (layer0_outputs(6307)) and (layer0_outputs(2976));
    layer1_outputs(6241) <= (layer0_outputs(6990)) xor (layer0_outputs(4256));
    layer1_outputs(6242) <= (layer0_outputs(4327)) and not (layer0_outputs(7493));
    layer1_outputs(6243) <= '1';
    layer1_outputs(6244) <= (layer0_outputs(4839)) and not (layer0_outputs(3801));
    layer1_outputs(6245) <= '0';
    layer1_outputs(6246) <= not(layer0_outputs(3211));
    layer1_outputs(6247) <= (layer0_outputs(3328)) and (layer0_outputs(6648));
    layer1_outputs(6248) <= layer0_outputs(1701);
    layer1_outputs(6249) <= layer0_outputs(1350);
    layer1_outputs(6250) <= not(layer0_outputs(3588)) or (layer0_outputs(208));
    layer1_outputs(6251) <= layer0_outputs(1070);
    layer1_outputs(6252) <= (layer0_outputs(2625)) or (layer0_outputs(7627));
    layer1_outputs(6253) <= not(layer0_outputs(610));
    layer1_outputs(6254) <= not(layer0_outputs(242)) or (layer0_outputs(5436));
    layer1_outputs(6255) <= '0';
    layer1_outputs(6256) <= not(layer0_outputs(5556)) or (layer0_outputs(6541));
    layer1_outputs(6257) <= not((layer0_outputs(5849)) or (layer0_outputs(3859)));
    layer1_outputs(6258) <= (layer0_outputs(7613)) and not (layer0_outputs(391));
    layer1_outputs(6259) <= (layer0_outputs(6629)) and not (layer0_outputs(2337));
    layer1_outputs(6260) <= not((layer0_outputs(1238)) xor (layer0_outputs(7383)));
    layer1_outputs(6261) <= layer0_outputs(3879);
    layer1_outputs(6262) <= layer0_outputs(6168);
    layer1_outputs(6263) <= not(layer0_outputs(4698)) or (layer0_outputs(3162));
    layer1_outputs(6264) <= not(layer0_outputs(6585));
    layer1_outputs(6265) <= (layer0_outputs(5150)) and not (layer0_outputs(4180));
    layer1_outputs(6266) <= not(layer0_outputs(1751));
    layer1_outputs(6267) <= (layer0_outputs(3089)) and not (layer0_outputs(2386));
    layer1_outputs(6268) <= not(layer0_outputs(6154));
    layer1_outputs(6269) <= not((layer0_outputs(2892)) xor (layer0_outputs(3631)));
    layer1_outputs(6270) <= not(layer0_outputs(7141)) or (layer0_outputs(2844));
    layer1_outputs(6271) <= not(layer0_outputs(6142)) or (layer0_outputs(1700));
    layer1_outputs(6272) <= (layer0_outputs(2369)) and (layer0_outputs(7019));
    layer1_outputs(6273) <= not((layer0_outputs(256)) and (layer0_outputs(615)));
    layer1_outputs(6274) <= not(layer0_outputs(1723)) or (layer0_outputs(3722));
    layer1_outputs(6275) <= not(layer0_outputs(1288));
    layer1_outputs(6276) <= (layer0_outputs(1819)) and not (layer0_outputs(4998));
    layer1_outputs(6277) <= (layer0_outputs(1162)) xor (layer0_outputs(6085));
    layer1_outputs(6278) <= (layer0_outputs(3705)) and not (layer0_outputs(7633));
    layer1_outputs(6279) <= (layer0_outputs(2016)) and not (layer0_outputs(6271));
    layer1_outputs(6280) <= '1';
    layer1_outputs(6281) <= (layer0_outputs(6152)) and not (layer0_outputs(3743));
    layer1_outputs(6282) <= '0';
    layer1_outputs(6283) <= not(layer0_outputs(6695));
    layer1_outputs(6284) <= layer0_outputs(4737);
    layer1_outputs(6285) <= not((layer0_outputs(3508)) and (layer0_outputs(6671)));
    layer1_outputs(6286) <= not(layer0_outputs(5848));
    layer1_outputs(6287) <= '0';
    layer1_outputs(6288) <= not((layer0_outputs(7443)) xor (layer0_outputs(1)));
    layer1_outputs(6289) <= not(layer0_outputs(7633));
    layer1_outputs(6290) <= layer0_outputs(3540);
    layer1_outputs(6291) <= (layer0_outputs(6681)) and not (layer0_outputs(1197));
    layer1_outputs(6292) <= (layer0_outputs(1293)) and not (layer0_outputs(4713));
    layer1_outputs(6293) <= not(layer0_outputs(3558));
    layer1_outputs(6294) <= not((layer0_outputs(2953)) xor (layer0_outputs(5796)));
    layer1_outputs(6295) <= not(layer0_outputs(5624)) or (layer0_outputs(2820));
    layer1_outputs(6296) <= '1';
    layer1_outputs(6297) <= (layer0_outputs(1012)) or (layer0_outputs(6137));
    layer1_outputs(6298) <= not(layer0_outputs(5950)) or (layer0_outputs(5755));
    layer1_outputs(6299) <= (layer0_outputs(4639)) or (layer0_outputs(7599));
    layer1_outputs(6300) <= layer0_outputs(1122);
    layer1_outputs(6301) <= (layer0_outputs(6412)) and not (layer0_outputs(4657));
    layer1_outputs(6302) <= layer0_outputs(601);
    layer1_outputs(6303) <= (layer0_outputs(7607)) and not (layer0_outputs(7012));
    layer1_outputs(6304) <= layer0_outputs(4271);
    layer1_outputs(6305) <= (layer0_outputs(5542)) or (layer0_outputs(5157));
    layer1_outputs(6306) <= not(layer0_outputs(5248)) or (layer0_outputs(4346));
    layer1_outputs(6307) <= (layer0_outputs(5094)) or (layer0_outputs(2778));
    layer1_outputs(6308) <= (layer0_outputs(3489)) and (layer0_outputs(3875));
    layer1_outputs(6309) <= not(layer0_outputs(3736)) or (layer0_outputs(3335));
    layer1_outputs(6310) <= not((layer0_outputs(3068)) and (layer0_outputs(1412)));
    layer1_outputs(6311) <= not(layer0_outputs(2501));
    layer1_outputs(6312) <= '0';
    layer1_outputs(6313) <= '1';
    layer1_outputs(6314) <= not((layer0_outputs(700)) or (layer0_outputs(4604)));
    layer1_outputs(6315) <= not(layer0_outputs(1290));
    layer1_outputs(6316) <= '0';
    layer1_outputs(6317) <= not(layer0_outputs(5458));
    layer1_outputs(6318) <= not(layer0_outputs(4796));
    layer1_outputs(6319) <= not(layer0_outputs(2179));
    layer1_outputs(6320) <= not((layer0_outputs(5847)) and (layer0_outputs(2547)));
    layer1_outputs(6321) <= not((layer0_outputs(1858)) or (layer0_outputs(732)));
    layer1_outputs(6322) <= (layer0_outputs(2560)) or (layer0_outputs(6971));
    layer1_outputs(6323) <= not(layer0_outputs(3983));
    layer1_outputs(6324) <= layer0_outputs(3422);
    layer1_outputs(6325) <= layer0_outputs(5276);
    layer1_outputs(6326) <= not((layer0_outputs(5574)) or (layer0_outputs(2774)));
    layer1_outputs(6327) <= not((layer0_outputs(3941)) or (layer0_outputs(300)));
    layer1_outputs(6328) <= not(layer0_outputs(1630));
    layer1_outputs(6329) <= not(layer0_outputs(4053));
    layer1_outputs(6330) <= layer0_outputs(52);
    layer1_outputs(6331) <= not(layer0_outputs(7109));
    layer1_outputs(6332) <= layer0_outputs(3159);
    layer1_outputs(6333) <= (layer0_outputs(5546)) and not (layer0_outputs(820));
    layer1_outputs(6334) <= (layer0_outputs(2940)) and (layer0_outputs(255));
    layer1_outputs(6335) <= not((layer0_outputs(1040)) and (layer0_outputs(2767)));
    layer1_outputs(6336) <= not((layer0_outputs(5035)) and (layer0_outputs(7171)));
    layer1_outputs(6337) <= (layer0_outputs(279)) or (layer0_outputs(4056));
    layer1_outputs(6338) <= layer0_outputs(2684);
    layer1_outputs(6339) <= (layer0_outputs(5566)) and (layer0_outputs(7106));
    layer1_outputs(6340) <= (layer0_outputs(2399)) and (layer0_outputs(5782));
    layer1_outputs(6341) <= layer0_outputs(1847);
    layer1_outputs(6342) <= '0';
    layer1_outputs(6343) <= layer0_outputs(4198);
    layer1_outputs(6344) <= (layer0_outputs(5500)) and not (layer0_outputs(5412));
    layer1_outputs(6345) <= layer0_outputs(1995);
    layer1_outputs(6346) <= not(layer0_outputs(313));
    layer1_outputs(6347) <= (layer0_outputs(4381)) and not (layer0_outputs(515));
    layer1_outputs(6348) <= (layer0_outputs(5500)) and not (layer0_outputs(4306));
    layer1_outputs(6349) <= (layer0_outputs(7095)) xor (layer0_outputs(3259));
    layer1_outputs(6350) <= layer0_outputs(7324);
    layer1_outputs(6351) <= layer0_outputs(5919);
    layer1_outputs(6352) <= not(layer0_outputs(972));
    layer1_outputs(6353) <= not((layer0_outputs(3169)) and (layer0_outputs(232)));
    layer1_outputs(6354) <= not((layer0_outputs(7395)) and (layer0_outputs(6967)));
    layer1_outputs(6355) <= layer0_outputs(2195);
    layer1_outputs(6356) <= not(layer0_outputs(155));
    layer1_outputs(6357) <= '0';
    layer1_outputs(6358) <= (layer0_outputs(4833)) or (layer0_outputs(3158));
    layer1_outputs(6359) <= '0';
    layer1_outputs(6360) <= '0';
    layer1_outputs(6361) <= '0';
    layer1_outputs(6362) <= (layer0_outputs(2698)) and not (layer0_outputs(1403));
    layer1_outputs(6363) <= layer0_outputs(5898);
    layer1_outputs(6364) <= not((layer0_outputs(1560)) or (layer0_outputs(3124)));
    layer1_outputs(6365) <= not(layer0_outputs(6996)) or (layer0_outputs(4739));
    layer1_outputs(6366) <= (layer0_outputs(6255)) or (layer0_outputs(7567));
    layer1_outputs(6367) <= '0';
    layer1_outputs(6368) <= layer0_outputs(2610);
    layer1_outputs(6369) <= '0';
    layer1_outputs(6370) <= (layer0_outputs(5915)) and not (layer0_outputs(1605));
    layer1_outputs(6371) <= not(layer0_outputs(3722)) or (layer0_outputs(4132));
    layer1_outputs(6372) <= not(layer0_outputs(349)) or (layer0_outputs(6995));
    layer1_outputs(6373) <= '0';
    layer1_outputs(6374) <= not((layer0_outputs(1292)) or (layer0_outputs(695)));
    layer1_outputs(6375) <= not((layer0_outputs(6458)) and (layer0_outputs(6308)));
    layer1_outputs(6376) <= not(layer0_outputs(245)) or (layer0_outputs(5432));
    layer1_outputs(6377) <= '0';
    layer1_outputs(6378) <= layer0_outputs(3003);
    layer1_outputs(6379) <= layer0_outputs(6000);
    layer1_outputs(6380) <= not(layer0_outputs(5981));
    layer1_outputs(6381) <= not(layer0_outputs(4173));
    layer1_outputs(6382) <= (layer0_outputs(2535)) and (layer0_outputs(3530));
    layer1_outputs(6383) <= not(layer0_outputs(7445));
    layer1_outputs(6384) <= (layer0_outputs(2062)) and (layer0_outputs(5839));
    layer1_outputs(6385) <= layer0_outputs(5061);
    layer1_outputs(6386) <= (layer0_outputs(5471)) and not (layer0_outputs(2014));
    layer1_outputs(6387) <= (layer0_outputs(5342)) and not (layer0_outputs(6331));
    layer1_outputs(6388) <= not((layer0_outputs(3393)) or (layer0_outputs(2984)));
    layer1_outputs(6389) <= '1';
    layer1_outputs(6390) <= not((layer0_outputs(1396)) and (layer0_outputs(7379)));
    layer1_outputs(6391) <= not((layer0_outputs(1814)) and (layer0_outputs(2192)));
    layer1_outputs(6392) <= not((layer0_outputs(752)) xor (layer0_outputs(4299)));
    layer1_outputs(6393) <= not(layer0_outputs(1793));
    layer1_outputs(6394) <= not((layer0_outputs(4789)) or (layer0_outputs(6007)));
    layer1_outputs(6395) <= not(layer0_outputs(2494));
    layer1_outputs(6396) <= (layer0_outputs(4961)) and (layer0_outputs(3867));
    layer1_outputs(6397) <= not(layer0_outputs(4174)) or (layer0_outputs(3511));
    layer1_outputs(6398) <= (layer0_outputs(7111)) and not (layer0_outputs(7588));
    layer1_outputs(6399) <= (layer0_outputs(6101)) and not (layer0_outputs(4777));
    layer1_outputs(6400) <= not((layer0_outputs(2278)) or (layer0_outputs(711)));
    layer1_outputs(6401) <= not(layer0_outputs(6976));
    layer1_outputs(6402) <= not(layer0_outputs(7563));
    layer1_outputs(6403) <= (layer0_outputs(3035)) xor (layer0_outputs(1777));
    layer1_outputs(6404) <= not(layer0_outputs(7266));
    layer1_outputs(6405) <= layer0_outputs(4681);
    layer1_outputs(6406) <= not(layer0_outputs(1097));
    layer1_outputs(6407) <= layer0_outputs(115);
    layer1_outputs(6408) <= (layer0_outputs(4686)) and (layer0_outputs(1985));
    layer1_outputs(6409) <= not(layer0_outputs(3717));
    layer1_outputs(6410) <= (layer0_outputs(3986)) or (layer0_outputs(4478));
    layer1_outputs(6411) <= (layer0_outputs(4199)) or (layer0_outputs(6223));
    layer1_outputs(6412) <= not(layer0_outputs(1885));
    layer1_outputs(6413) <= (layer0_outputs(4571)) and not (layer0_outputs(5820));
    layer1_outputs(6414) <= layer0_outputs(2751);
    layer1_outputs(6415) <= '0';
    layer1_outputs(6416) <= (layer0_outputs(4819)) and not (layer0_outputs(2433));
    layer1_outputs(6417) <= (layer0_outputs(3362)) or (layer0_outputs(5282));
    layer1_outputs(6418) <= not(layer0_outputs(4423));
    layer1_outputs(6419) <= (layer0_outputs(2285)) and (layer0_outputs(4082));
    layer1_outputs(6420) <= not((layer0_outputs(5624)) or (layer0_outputs(2325)));
    layer1_outputs(6421) <= not(layer0_outputs(3895)) or (layer0_outputs(4491));
    layer1_outputs(6422) <= not(layer0_outputs(1672));
    layer1_outputs(6423) <= not(layer0_outputs(746));
    layer1_outputs(6424) <= '1';
    layer1_outputs(6425) <= (layer0_outputs(1232)) and not (layer0_outputs(1706));
    layer1_outputs(6426) <= (layer0_outputs(513)) and (layer0_outputs(683));
    layer1_outputs(6427) <= layer0_outputs(3961);
    layer1_outputs(6428) <= (layer0_outputs(2193)) xor (layer0_outputs(6543));
    layer1_outputs(6429) <= not(layer0_outputs(4891));
    layer1_outputs(6430) <= '0';
    layer1_outputs(6431) <= not((layer0_outputs(3975)) or (layer0_outputs(25)));
    layer1_outputs(6432) <= (layer0_outputs(7414)) and not (layer0_outputs(7062));
    layer1_outputs(6433) <= not(layer0_outputs(3085));
    layer1_outputs(6434) <= layer0_outputs(5668);
    layer1_outputs(6435) <= layer0_outputs(670);
    layer1_outputs(6436) <= (layer0_outputs(2777)) or (layer0_outputs(6733));
    layer1_outputs(6437) <= layer0_outputs(483);
    layer1_outputs(6438) <= not(layer0_outputs(5131));
    layer1_outputs(6439) <= not(layer0_outputs(3938)) or (layer0_outputs(2303));
    layer1_outputs(6440) <= layer0_outputs(4002);
    layer1_outputs(6441) <= not(layer0_outputs(7257));
    layer1_outputs(6442) <= not(layer0_outputs(5259));
    layer1_outputs(6443) <= (layer0_outputs(7098)) or (layer0_outputs(5057));
    layer1_outputs(6444) <= not(layer0_outputs(7067));
    layer1_outputs(6445) <= (layer0_outputs(7189)) and not (layer0_outputs(2838));
    layer1_outputs(6446) <= not(layer0_outputs(12));
    layer1_outputs(6447) <= not(layer0_outputs(2403));
    layer1_outputs(6448) <= not(layer0_outputs(5703)) or (layer0_outputs(535));
    layer1_outputs(6449) <= (layer0_outputs(7045)) xor (layer0_outputs(1564));
    layer1_outputs(6450) <= not(layer0_outputs(6106));
    layer1_outputs(6451) <= not((layer0_outputs(5775)) and (layer0_outputs(5693)));
    layer1_outputs(6452) <= layer0_outputs(6807);
    layer1_outputs(6453) <= (layer0_outputs(3491)) and not (layer0_outputs(6399));
    layer1_outputs(6454) <= (layer0_outputs(5461)) or (layer0_outputs(1820));
    layer1_outputs(6455) <= (layer0_outputs(4058)) and not (layer0_outputs(3725));
    layer1_outputs(6456) <= not((layer0_outputs(2664)) and (layer0_outputs(4289)));
    layer1_outputs(6457) <= (layer0_outputs(7420)) and not (layer0_outputs(964));
    layer1_outputs(6458) <= layer0_outputs(3430);
    layer1_outputs(6459) <= not((layer0_outputs(1525)) or (layer0_outputs(900)));
    layer1_outputs(6460) <= not((layer0_outputs(6209)) or (layer0_outputs(4168)));
    layer1_outputs(6461) <= not(layer0_outputs(319));
    layer1_outputs(6462) <= not(layer0_outputs(7104));
    layer1_outputs(6463) <= (layer0_outputs(2023)) or (layer0_outputs(4774));
    layer1_outputs(6464) <= layer0_outputs(1877);
    layer1_outputs(6465) <= not(layer0_outputs(6285));
    layer1_outputs(6466) <= not(layer0_outputs(5350));
    layer1_outputs(6467) <= (layer0_outputs(4508)) or (layer0_outputs(6784));
    layer1_outputs(6468) <= layer0_outputs(3343);
    layer1_outputs(6469) <= layer0_outputs(1795);
    layer1_outputs(6470) <= not(layer0_outputs(864));
    layer1_outputs(6471) <= (layer0_outputs(3776)) and (layer0_outputs(4728));
    layer1_outputs(6472) <= not(layer0_outputs(4370));
    layer1_outputs(6473) <= '1';
    layer1_outputs(6474) <= '1';
    layer1_outputs(6475) <= not(layer0_outputs(6774)) or (layer0_outputs(5427));
    layer1_outputs(6476) <= not(layer0_outputs(6279));
    layer1_outputs(6477) <= layer0_outputs(3925);
    layer1_outputs(6478) <= '0';
    layer1_outputs(6479) <= layer0_outputs(6826);
    layer1_outputs(6480) <= not((layer0_outputs(3402)) and (layer0_outputs(704)));
    layer1_outputs(6481) <= (layer0_outputs(4018)) and (layer0_outputs(7148));
    layer1_outputs(6482) <= '0';
    layer1_outputs(6483) <= not(layer0_outputs(7101));
    layer1_outputs(6484) <= not(layer0_outputs(4044));
    layer1_outputs(6485) <= not(layer0_outputs(5743));
    layer1_outputs(6486) <= (layer0_outputs(2440)) and not (layer0_outputs(5970));
    layer1_outputs(6487) <= layer0_outputs(3424);
    layer1_outputs(6488) <= not(layer0_outputs(152));
    layer1_outputs(6489) <= (layer0_outputs(3977)) and (layer0_outputs(3190));
    layer1_outputs(6490) <= not(layer0_outputs(2977));
    layer1_outputs(6491) <= layer0_outputs(2194);
    layer1_outputs(6492) <= '1';
    layer1_outputs(6493) <= not(layer0_outputs(441));
    layer1_outputs(6494) <= layer0_outputs(7147);
    layer1_outputs(6495) <= (layer0_outputs(267)) and not (layer0_outputs(3793));
    layer1_outputs(6496) <= '0';
    layer1_outputs(6497) <= (layer0_outputs(395)) and not (layer0_outputs(2159));
    layer1_outputs(6498) <= (layer0_outputs(854)) and not (layer0_outputs(2461));
    layer1_outputs(6499) <= not((layer0_outputs(4576)) or (layer0_outputs(2151)));
    layer1_outputs(6500) <= (layer0_outputs(5007)) and not (layer0_outputs(4052));
    layer1_outputs(6501) <= not(layer0_outputs(7577)) or (layer0_outputs(77));
    layer1_outputs(6502) <= not(layer0_outputs(1004));
    layer1_outputs(6503) <= '1';
    layer1_outputs(6504) <= layer0_outputs(2527);
    layer1_outputs(6505) <= not(layer0_outputs(2088));
    layer1_outputs(6506) <= not((layer0_outputs(2546)) or (layer0_outputs(5874)));
    layer1_outputs(6507) <= layer0_outputs(2799);
    layer1_outputs(6508) <= not((layer0_outputs(450)) or (layer0_outputs(5608)));
    layer1_outputs(6509) <= not(layer0_outputs(3897));
    layer1_outputs(6510) <= '1';
    layer1_outputs(6511) <= not(layer0_outputs(7459));
    layer1_outputs(6512) <= layer0_outputs(6617);
    layer1_outputs(6513) <= not(layer0_outputs(3798));
    layer1_outputs(6514) <= not(layer0_outputs(3026)) or (layer0_outputs(1430));
    layer1_outputs(6515) <= (layer0_outputs(1053)) and not (layer0_outputs(6842));
    layer1_outputs(6516) <= (layer0_outputs(798)) or (layer0_outputs(2394));
    layer1_outputs(6517) <= not(layer0_outputs(5607));
    layer1_outputs(6518) <= (layer0_outputs(69)) and not (layer0_outputs(3047));
    layer1_outputs(6519) <= (layer0_outputs(2759)) and not (layer0_outputs(5072));
    layer1_outputs(6520) <= not(layer0_outputs(2191)) or (layer0_outputs(3650));
    layer1_outputs(6521) <= not(layer0_outputs(244)) or (layer0_outputs(6548));
    layer1_outputs(6522) <= not(layer0_outputs(1544)) or (layer0_outputs(43));
    layer1_outputs(6523) <= not(layer0_outputs(6262));
    layer1_outputs(6524) <= not(layer0_outputs(6713));
    layer1_outputs(6525) <= not(layer0_outputs(703)) or (layer0_outputs(3868));
    layer1_outputs(6526) <= layer0_outputs(512);
    layer1_outputs(6527) <= not(layer0_outputs(3198)) or (layer0_outputs(1494));
    layer1_outputs(6528) <= not((layer0_outputs(4845)) or (layer0_outputs(893)));
    layer1_outputs(6529) <= layer0_outputs(4067);
    layer1_outputs(6530) <= not(layer0_outputs(6265));
    layer1_outputs(6531) <= not((layer0_outputs(3828)) xor (layer0_outputs(320)));
    layer1_outputs(6532) <= not(layer0_outputs(2464)) or (layer0_outputs(1959));
    layer1_outputs(6533) <= (layer0_outputs(462)) and not (layer0_outputs(2786));
    layer1_outputs(6534) <= not(layer0_outputs(5884));
    layer1_outputs(6535) <= layer0_outputs(685);
    layer1_outputs(6536) <= (layer0_outputs(4255)) or (layer0_outputs(6503));
    layer1_outputs(6537) <= not((layer0_outputs(5920)) or (layer0_outputs(4540)));
    layer1_outputs(6538) <= '1';
    layer1_outputs(6539) <= not((layer0_outputs(2558)) and (layer0_outputs(2556)));
    layer1_outputs(6540) <= (layer0_outputs(1295)) or (layer0_outputs(6441));
    layer1_outputs(6541) <= (layer0_outputs(1739)) and not (layer0_outputs(6694));
    layer1_outputs(6542) <= not(layer0_outputs(3388));
    layer1_outputs(6543) <= not(layer0_outputs(493)) or (layer0_outputs(3805));
    layer1_outputs(6544) <= not(layer0_outputs(2456));
    layer1_outputs(6545) <= not(layer0_outputs(2457));
    layer1_outputs(6546) <= (layer0_outputs(3072)) or (layer0_outputs(3485));
    layer1_outputs(6547) <= not((layer0_outputs(3881)) and (layer0_outputs(4750)));
    layer1_outputs(6548) <= not((layer0_outputs(7375)) and (layer0_outputs(4352)));
    layer1_outputs(6549) <= not(layer0_outputs(4086));
    layer1_outputs(6550) <= (layer0_outputs(562)) and not (layer0_outputs(719));
    layer1_outputs(6551) <= not(layer0_outputs(3107));
    layer1_outputs(6552) <= '0';
    layer1_outputs(6553) <= not(layer0_outputs(3775));
    layer1_outputs(6554) <= not(layer0_outputs(4001));
    layer1_outputs(6555) <= (layer0_outputs(4290)) and not (layer0_outputs(5651));
    layer1_outputs(6556) <= layer0_outputs(1893);
    layer1_outputs(6557) <= not(layer0_outputs(2743));
    layer1_outputs(6558) <= not(layer0_outputs(3509));
    layer1_outputs(6559) <= (layer0_outputs(5448)) and not (layer0_outputs(2960));
    layer1_outputs(6560) <= '1';
    layer1_outputs(6561) <= layer0_outputs(5334);
    layer1_outputs(6562) <= not(layer0_outputs(3345));
    layer1_outputs(6563) <= not(layer0_outputs(7084));
    layer1_outputs(6564) <= (layer0_outputs(6465)) and (layer0_outputs(5719));
    layer1_outputs(6565) <= not((layer0_outputs(7305)) or (layer0_outputs(1286)));
    layer1_outputs(6566) <= not((layer0_outputs(7172)) and (layer0_outputs(4011)));
    layer1_outputs(6567) <= not(layer0_outputs(7161));
    layer1_outputs(6568) <= layer0_outputs(2321);
    layer1_outputs(6569) <= (layer0_outputs(6052)) and not (layer0_outputs(5253));
    layer1_outputs(6570) <= layer0_outputs(2756);
    layer1_outputs(6571) <= not((layer0_outputs(4003)) or (layer0_outputs(4893)));
    layer1_outputs(6572) <= not(layer0_outputs(5240));
    layer1_outputs(6573) <= (layer0_outputs(1677)) and not (layer0_outputs(1857));
    layer1_outputs(6574) <= not((layer0_outputs(5797)) and (layer0_outputs(7006)));
    layer1_outputs(6575) <= (layer0_outputs(366)) and (layer0_outputs(2770));
    layer1_outputs(6576) <= not(layer0_outputs(5403));
    layer1_outputs(6577) <= not((layer0_outputs(4811)) or (layer0_outputs(4500)));
    layer1_outputs(6578) <= not((layer0_outputs(3714)) and (layer0_outputs(6953)));
    layer1_outputs(6579) <= not((layer0_outputs(4127)) or (layer0_outputs(1332)));
    layer1_outputs(6580) <= (layer0_outputs(4826)) or (layer0_outputs(3003));
    layer1_outputs(6581) <= not(layer0_outputs(2614));
    layer1_outputs(6582) <= not(layer0_outputs(5844));
    layer1_outputs(6583) <= not((layer0_outputs(4804)) and (layer0_outputs(3153)));
    layer1_outputs(6584) <= layer0_outputs(6248);
    layer1_outputs(6585) <= '1';
    layer1_outputs(6586) <= layer0_outputs(921);
    layer1_outputs(6587) <= layer0_outputs(3072);
    layer1_outputs(6588) <= (layer0_outputs(6134)) and not (layer0_outputs(366));
    layer1_outputs(6589) <= (layer0_outputs(5053)) and not (layer0_outputs(1416));
    layer1_outputs(6590) <= not((layer0_outputs(3039)) xor (layer0_outputs(3579)));
    layer1_outputs(6591) <= layer0_outputs(6841);
    layer1_outputs(6592) <= '0';
    layer1_outputs(6593) <= (layer0_outputs(6400)) or (layer0_outputs(5946));
    layer1_outputs(6594) <= not((layer0_outputs(3170)) or (layer0_outputs(1987)));
    layer1_outputs(6595) <= (layer0_outputs(5784)) and (layer0_outputs(2350));
    layer1_outputs(6596) <= '0';
    layer1_outputs(6597) <= (layer0_outputs(5888)) and not (layer0_outputs(7231));
    layer1_outputs(6598) <= not((layer0_outputs(5037)) and (layer0_outputs(7329)));
    layer1_outputs(6599) <= (layer0_outputs(4763)) and not (layer0_outputs(2969));
    layer1_outputs(6600) <= layer0_outputs(7100);
    layer1_outputs(6601) <= not(layer0_outputs(342));
    layer1_outputs(6602) <= not((layer0_outputs(1322)) and (layer0_outputs(2214)));
    layer1_outputs(6603) <= not(layer0_outputs(651));
    layer1_outputs(6604) <= not((layer0_outputs(2780)) and (layer0_outputs(6466)));
    layer1_outputs(6605) <= (layer0_outputs(6511)) and not (layer0_outputs(6224));
    layer1_outputs(6606) <= (layer0_outputs(2870)) or (layer0_outputs(6487));
    layer1_outputs(6607) <= layer0_outputs(7427);
    layer1_outputs(6608) <= (layer0_outputs(6976)) and (layer0_outputs(6115));
    layer1_outputs(6609) <= not(layer0_outputs(5832)) or (layer0_outputs(1110));
    layer1_outputs(6610) <= layer0_outputs(6586);
    layer1_outputs(6611) <= layer0_outputs(4265);
    layer1_outputs(6612) <= (layer0_outputs(2036)) and (layer0_outputs(5972));
    layer1_outputs(6613) <= (layer0_outputs(532)) and not (layer0_outputs(7216));
    layer1_outputs(6614) <= (layer0_outputs(5314)) and (layer0_outputs(3901));
    layer1_outputs(6615) <= layer0_outputs(4264);
    layer1_outputs(6616) <= layer0_outputs(7259);
    layer1_outputs(6617) <= layer0_outputs(1868);
    layer1_outputs(6618) <= not((layer0_outputs(1282)) and (layer0_outputs(1988)));
    layer1_outputs(6619) <= (layer0_outputs(1319)) or (layer0_outputs(53));
    layer1_outputs(6620) <= (layer0_outputs(1020)) and not (layer0_outputs(6361));
    layer1_outputs(6621) <= layer0_outputs(7086);
    layer1_outputs(6622) <= not(layer0_outputs(6840)) or (layer0_outputs(6047));
    layer1_outputs(6623) <= (layer0_outputs(6411)) and not (layer0_outputs(6256));
    layer1_outputs(6624) <= not(layer0_outputs(1511));
    layer1_outputs(6625) <= (layer0_outputs(4217)) and not (layer0_outputs(6702));
    layer1_outputs(6626) <= layer0_outputs(1889);
    layer1_outputs(6627) <= not((layer0_outputs(5214)) and (layer0_outputs(6708)));
    layer1_outputs(6628) <= (layer0_outputs(5506)) and not (layer0_outputs(335));
    layer1_outputs(6629) <= not((layer0_outputs(7530)) xor (layer0_outputs(5426)));
    layer1_outputs(6630) <= layer0_outputs(3022);
    layer1_outputs(6631) <= not(layer0_outputs(71));
    layer1_outputs(6632) <= (layer0_outputs(5370)) and not (layer0_outputs(723));
    layer1_outputs(6633) <= not(layer0_outputs(4205));
    layer1_outputs(6634) <= (layer0_outputs(2486)) and (layer0_outputs(6036));
    layer1_outputs(6635) <= (layer0_outputs(4569)) xor (layer0_outputs(4075));
    layer1_outputs(6636) <= not((layer0_outputs(7491)) and (layer0_outputs(6391)));
    layer1_outputs(6637) <= not(layer0_outputs(2068)) or (layer0_outputs(1934));
    layer1_outputs(6638) <= '1';
    layer1_outputs(6639) <= layer0_outputs(4454);
    layer1_outputs(6640) <= (layer0_outputs(7428)) and not (layer0_outputs(339));
    layer1_outputs(6641) <= not((layer0_outputs(3215)) xor (layer0_outputs(2139)));
    layer1_outputs(6642) <= layer0_outputs(2184);
    layer1_outputs(6643) <= (layer0_outputs(6181)) and (layer0_outputs(3411));
    layer1_outputs(6644) <= '0';
    layer1_outputs(6645) <= not((layer0_outputs(6709)) and (layer0_outputs(4242)));
    layer1_outputs(6646) <= layer0_outputs(6733);
    layer1_outputs(6647) <= not(layer0_outputs(679)) or (layer0_outputs(1411));
    layer1_outputs(6648) <= '0';
    layer1_outputs(6649) <= not(layer0_outputs(4582));
    layer1_outputs(6650) <= not((layer0_outputs(3466)) and (layer0_outputs(806)));
    layer1_outputs(6651) <= not((layer0_outputs(5223)) and (layer0_outputs(7586)));
    layer1_outputs(6652) <= not(layer0_outputs(989)) or (layer0_outputs(2400));
    layer1_outputs(6653) <= (layer0_outputs(2208)) and not (layer0_outputs(7596));
    layer1_outputs(6654) <= not((layer0_outputs(7043)) and (layer0_outputs(6612)));
    layer1_outputs(6655) <= not(layer0_outputs(3385)) or (layer0_outputs(5449));
    layer1_outputs(6656) <= (layer0_outputs(3234)) and not (layer0_outputs(2701));
    layer1_outputs(6657) <= (layer0_outputs(565)) and not (layer0_outputs(5008));
    layer1_outputs(6658) <= not(layer0_outputs(5176));
    layer1_outputs(6659) <= not(layer0_outputs(4407)) or (layer0_outputs(118));
    layer1_outputs(6660) <= '1';
    layer1_outputs(6661) <= layer0_outputs(4188);
    layer1_outputs(6662) <= not(layer0_outputs(5153));
    layer1_outputs(6663) <= not((layer0_outputs(1904)) or (layer0_outputs(5631)));
    layer1_outputs(6664) <= not(layer0_outputs(57));
    layer1_outputs(6665) <= not(layer0_outputs(1732));
    layer1_outputs(6666) <= (layer0_outputs(4824)) and not (layer0_outputs(6083));
    layer1_outputs(6667) <= '0';
    layer1_outputs(6668) <= not(layer0_outputs(3219));
    layer1_outputs(6669) <= not(layer0_outputs(4261));
    layer1_outputs(6670) <= (layer0_outputs(4950)) and not (layer0_outputs(5790));
    layer1_outputs(6671) <= not(layer0_outputs(6016));
    layer1_outputs(6672) <= not(layer0_outputs(4159)) or (layer0_outputs(2308));
    layer1_outputs(6673) <= not((layer0_outputs(5702)) or (layer0_outputs(7277)));
    layer1_outputs(6674) <= '1';
    layer1_outputs(6675) <= (layer0_outputs(6519)) and not (layer0_outputs(304));
    layer1_outputs(6676) <= (layer0_outputs(5541)) and not (layer0_outputs(7280));
    layer1_outputs(6677) <= not(layer0_outputs(1844)) or (layer0_outputs(6174));
    layer1_outputs(6678) <= (layer0_outputs(6444)) and (layer0_outputs(1787));
    layer1_outputs(6679) <= layer0_outputs(4668);
    layer1_outputs(6680) <= not(layer0_outputs(661));
    layer1_outputs(6681) <= layer0_outputs(5433);
    layer1_outputs(6682) <= layer0_outputs(6308);
    layer1_outputs(6683) <= not((layer0_outputs(406)) and (layer0_outputs(6514)));
    layer1_outputs(6684) <= not(layer0_outputs(6533)) or (layer0_outputs(6956));
    layer1_outputs(6685) <= not(layer0_outputs(5659)) or (layer0_outputs(6432));
    layer1_outputs(6686) <= (layer0_outputs(1535)) or (layer0_outputs(2254));
    layer1_outputs(6687) <= layer0_outputs(1332);
    layer1_outputs(6688) <= '1';
    layer1_outputs(6689) <= (layer0_outputs(1691)) or (layer0_outputs(4456));
    layer1_outputs(6690) <= '1';
    layer1_outputs(6691) <= '1';
    layer1_outputs(6692) <= (layer0_outputs(1578)) or (layer0_outputs(2251));
    layer1_outputs(6693) <= not(layer0_outputs(487));
    layer1_outputs(6694) <= not(layer0_outputs(2500)) or (layer0_outputs(7562));
    layer1_outputs(6695) <= (layer0_outputs(1961)) or (layer0_outputs(7302));
    layer1_outputs(6696) <= (layer0_outputs(7075)) and not (layer0_outputs(2087));
    layer1_outputs(6697) <= layer0_outputs(1482);
    layer1_outputs(6698) <= not(layer0_outputs(4776)) or (layer0_outputs(6727));
    layer1_outputs(6699) <= (layer0_outputs(7061)) and not (layer0_outputs(6015));
    layer1_outputs(6700) <= (layer0_outputs(226)) and not (layer0_outputs(5251));
    layer1_outputs(6701) <= not((layer0_outputs(4130)) and (layer0_outputs(5667)));
    layer1_outputs(6702) <= layer0_outputs(2171);
    layer1_outputs(6703) <= not(layer0_outputs(5622));
    layer1_outputs(6704) <= not(layer0_outputs(2923));
    layer1_outputs(6705) <= not(layer0_outputs(5300)) or (layer0_outputs(1364));
    layer1_outputs(6706) <= (layer0_outputs(6662)) xor (layer0_outputs(5523));
    layer1_outputs(6707) <= '0';
    layer1_outputs(6708) <= not(layer0_outputs(1100));
    layer1_outputs(6709) <= not(layer0_outputs(5869)) or (layer0_outputs(5634));
    layer1_outputs(6710) <= layer0_outputs(1761);
    layer1_outputs(6711) <= '0';
    layer1_outputs(6712) <= layer0_outputs(3831);
    layer1_outputs(6713) <= (layer0_outputs(6720)) and not (layer0_outputs(7418));
    layer1_outputs(6714) <= (layer0_outputs(3775)) and not (layer0_outputs(73));
    layer1_outputs(6715) <= (layer0_outputs(1395)) xor (layer0_outputs(6234));
    layer1_outputs(6716) <= not(layer0_outputs(4796));
    layer1_outputs(6717) <= (layer0_outputs(5415)) xor (layer0_outputs(2271));
    layer1_outputs(6718) <= '0';
    layer1_outputs(6719) <= (layer0_outputs(6998)) and not (layer0_outputs(3887));
    layer1_outputs(6720) <= (layer0_outputs(6834)) or (layer0_outputs(4517));
    layer1_outputs(6721) <= '1';
    layer1_outputs(6722) <= not((layer0_outputs(3187)) or (layer0_outputs(101)));
    layer1_outputs(6723) <= not(layer0_outputs(1901));
    layer1_outputs(6724) <= (layer0_outputs(5313)) and not (layer0_outputs(837));
    layer1_outputs(6725) <= not(layer0_outputs(1652));
    layer1_outputs(6726) <= (layer0_outputs(6427)) and (layer0_outputs(5938));
    layer1_outputs(6727) <= (layer0_outputs(3782)) xor (layer0_outputs(22));
    layer1_outputs(6728) <= (layer0_outputs(4383)) and not (layer0_outputs(234));
    layer1_outputs(6729) <= '0';
    layer1_outputs(6730) <= not(layer0_outputs(2829));
    layer1_outputs(6731) <= not(layer0_outputs(286));
    layer1_outputs(6732) <= (layer0_outputs(2921)) and not (layer0_outputs(686));
    layer1_outputs(6733) <= '0';
    layer1_outputs(6734) <= not(layer0_outputs(4584)) or (layer0_outputs(3628));
    layer1_outputs(6735) <= not((layer0_outputs(7228)) and (layer0_outputs(3684)));
    layer1_outputs(6736) <= (layer0_outputs(6547)) and not (layer0_outputs(7512));
    layer1_outputs(6737) <= '0';
    layer1_outputs(6738) <= not((layer0_outputs(2355)) and (layer0_outputs(7489)));
    layer1_outputs(6739) <= not((layer0_outputs(4087)) and (layer0_outputs(6598)));
    layer1_outputs(6740) <= not(layer0_outputs(1709));
    layer1_outputs(6741) <= (layer0_outputs(1602)) or (layer0_outputs(4136));
    layer1_outputs(6742) <= '0';
    layer1_outputs(6743) <= layer0_outputs(5211);
    layer1_outputs(6744) <= not(layer0_outputs(5803)) or (layer0_outputs(3724));
    layer1_outputs(6745) <= (layer0_outputs(5393)) or (layer0_outputs(1452));
    layer1_outputs(6746) <= layer0_outputs(5987);
    layer1_outputs(6747) <= not(layer0_outputs(2510));
    layer1_outputs(6748) <= not(layer0_outputs(3440)) or (layer0_outputs(2915));
    layer1_outputs(6749) <= (layer0_outputs(2310)) or (layer0_outputs(6636));
    layer1_outputs(6750) <= not((layer0_outputs(6476)) xor (layer0_outputs(5234)));
    layer1_outputs(6751) <= layer0_outputs(851);
    layer1_outputs(6752) <= not((layer0_outputs(6367)) xor (layer0_outputs(50)));
    layer1_outputs(6753) <= not((layer0_outputs(6866)) or (layer0_outputs(4477)));
    layer1_outputs(6754) <= '0';
    layer1_outputs(6755) <= layer0_outputs(6905);
    layer1_outputs(6756) <= not(layer0_outputs(1900));
    layer1_outputs(6757) <= (layer0_outputs(585)) xor (layer0_outputs(1163));
    layer1_outputs(6758) <= (layer0_outputs(6790)) and not (layer0_outputs(1133));
    layer1_outputs(6759) <= not(layer0_outputs(6001));
    layer1_outputs(6760) <= not(layer0_outputs(2741)) or (layer0_outputs(680));
    layer1_outputs(6761) <= '1';
    layer1_outputs(6762) <= not(layer0_outputs(7525));
    layer1_outputs(6763) <= not(layer0_outputs(6738)) or (layer0_outputs(6045));
    layer1_outputs(6764) <= not((layer0_outputs(3424)) and (layer0_outputs(4164)));
    layer1_outputs(6765) <= not(layer0_outputs(4908));
    layer1_outputs(6766) <= layer0_outputs(3196);
    layer1_outputs(6767) <= not(layer0_outputs(1582));
    layer1_outputs(6768) <= (layer0_outputs(4628)) and (layer0_outputs(1223));
    layer1_outputs(6769) <= not((layer0_outputs(1991)) or (layer0_outputs(1409)));
    layer1_outputs(6770) <= layer0_outputs(6796);
    layer1_outputs(6771) <= not(layer0_outputs(5164));
    layer1_outputs(6772) <= not(layer0_outputs(6565));
    layer1_outputs(6773) <= not(layer0_outputs(1741)) or (layer0_outputs(5608));
    layer1_outputs(6774) <= (layer0_outputs(5189)) and not (layer0_outputs(2102));
    layer1_outputs(6775) <= (layer0_outputs(5989)) xor (layer0_outputs(4284));
    layer1_outputs(6776) <= not(layer0_outputs(1452));
    layer1_outputs(6777) <= not(layer0_outputs(5569));
    layer1_outputs(6778) <= not(layer0_outputs(6144));
    layer1_outputs(6779) <= not((layer0_outputs(1016)) xor (layer0_outputs(94)));
    layer1_outputs(6780) <= not((layer0_outputs(2091)) and (layer0_outputs(6195)));
    layer1_outputs(6781) <= (layer0_outputs(7550)) xor (layer0_outputs(3954));
    layer1_outputs(6782) <= (layer0_outputs(3591)) and (layer0_outputs(2345));
    layer1_outputs(6783) <= (layer0_outputs(3149)) xor (layer0_outputs(230));
    layer1_outputs(6784) <= '1';
    layer1_outputs(6785) <= not((layer0_outputs(1582)) and (layer0_outputs(5511)));
    layer1_outputs(6786) <= layer0_outputs(4399);
    layer1_outputs(6787) <= (layer0_outputs(7099)) and (layer0_outputs(2794));
    layer1_outputs(6788) <= (layer0_outputs(1281)) and not (layer0_outputs(5339));
    layer1_outputs(6789) <= (layer0_outputs(186)) and not (layer0_outputs(7295));
    layer1_outputs(6790) <= layer0_outputs(4387);
    layer1_outputs(6791) <= (layer0_outputs(5328)) and not (layer0_outputs(1024));
    layer1_outputs(6792) <= (layer0_outputs(2302)) or (layer0_outputs(7163));
    layer1_outputs(6793) <= layer0_outputs(5094);
    layer1_outputs(6794) <= not(layer0_outputs(4334));
    layer1_outputs(6795) <= not((layer0_outputs(7631)) and (layer0_outputs(3932)));
    layer1_outputs(6796) <= (layer0_outputs(7132)) or (layer0_outputs(4672));
    layer1_outputs(6797) <= layer0_outputs(6397);
    layer1_outputs(6798) <= '1';
    layer1_outputs(6799) <= (layer0_outputs(2190)) and (layer0_outputs(5068));
    layer1_outputs(6800) <= layer0_outputs(87);
    layer1_outputs(6801) <= not(layer0_outputs(6113));
    layer1_outputs(6802) <= not((layer0_outputs(6439)) and (layer0_outputs(2353)));
    layer1_outputs(6803) <= (layer0_outputs(2788)) or (layer0_outputs(4362));
    layer1_outputs(6804) <= layer0_outputs(5531);
    layer1_outputs(6805) <= '1';
    layer1_outputs(6806) <= layer0_outputs(6566);
    layer1_outputs(6807) <= layer0_outputs(4677);
    layer1_outputs(6808) <= layer0_outputs(160);
    layer1_outputs(6809) <= (layer0_outputs(6812)) and (layer0_outputs(4778));
    layer1_outputs(6810) <= (layer0_outputs(5759)) and (layer0_outputs(6696));
    layer1_outputs(6811) <= layer0_outputs(7534);
    layer1_outputs(6812) <= (layer0_outputs(1602)) and not (layer0_outputs(1330));
    layer1_outputs(6813) <= not((layer0_outputs(1191)) or (layer0_outputs(2099)));
    layer1_outputs(6814) <= (layer0_outputs(6598)) and not (layer0_outputs(2359));
    layer1_outputs(6815) <= (layer0_outputs(4680)) and not (layer0_outputs(5502));
    layer1_outputs(6816) <= (layer0_outputs(2753)) and (layer0_outputs(1305));
    layer1_outputs(6817) <= not((layer0_outputs(1013)) xor (layer0_outputs(2777)));
    layer1_outputs(6818) <= (layer0_outputs(1611)) and not (layer0_outputs(1047));
    layer1_outputs(6819) <= not(layer0_outputs(5309)) or (layer0_outputs(1259));
    layer1_outputs(6820) <= (layer0_outputs(6791)) or (layer0_outputs(810));
    layer1_outputs(6821) <= layer0_outputs(3962);
    layer1_outputs(6822) <= not(layer0_outputs(2817));
    layer1_outputs(6823) <= '0';
    layer1_outputs(6824) <= layer0_outputs(7552);
    layer1_outputs(6825) <= (layer0_outputs(459)) and not (layer0_outputs(1603));
    layer1_outputs(6826) <= not(layer0_outputs(2750));
    layer1_outputs(6827) <= (layer0_outputs(4201)) and not (layer0_outputs(1140));
    layer1_outputs(6828) <= (layer0_outputs(5781)) and not (layer0_outputs(6717));
    layer1_outputs(6829) <= not(layer0_outputs(3976));
    layer1_outputs(6830) <= (layer0_outputs(1623)) and not (layer0_outputs(449));
    layer1_outputs(6831) <= not((layer0_outputs(1756)) and (layer0_outputs(7236)));
    layer1_outputs(6832) <= not(layer0_outputs(4240)) or (layer0_outputs(4530));
    layer1_outputs(6833) <= not(layer0_outputs(5583)) or (layer0_outputs(7545));
    layer1_outputs(6834) <= (layer0_outputs(1527)) and (layer0_outputs(5355));
    layer1_outputs(6835) <= '1';
    layer1_outputs(6836) <= '1';
    layer1_outputs(6837) <= not(layer0_outputs(5788));
    layer1_outputs(6838) <= (layer0_outputs(7249)) and not (layer0_outputs(1));
    layer1_outputs(6839) <= layer0_outputs(6767);
    layer1_outputs(6840) <= '1';
    layer1_outputs(6841) <= not(layer0_outputs(1523));
    layer1_outputs(6842) <= (layer0_outputs(2648)) and (layer0_outputs(4310));
    layer1_outputs(6843) <= layer0_outputs(2395);
    layer1_outputs(6844) <= not((layer0_outputs(2967)) or (layer0_outputs(1373)));
    layer1_outputs(6845) <= (layer0_outputs(1439)) and not (layer0_outputs(2417));
    layer1_outputs(6846) <= not(layer0_outputs(1649));
    layer1_outputs(6847) <= layer0_outputs(2832);
    layer1_outputs(6848) <= not(layer0_outputs(7637));
    layer1_outputs(6849) <= not(layer0_outputs(1723)) or (layer0_outputs(4294));
    layer1_outputs(6850) <= not((layer0_outputs(5332)) and (layer0_outputs(4170)));
    layer1_outputs(6851) <= (layer0_outputs(4822)) and not (layer0_outputs(1691));
    layer1_outputs(6852) <= (layer0_outputs(5142)) xor (layer0_outputs(1609));
    layer1_outputs(6853) <= not(layer0_outputs(2028)) or (layer0_outputs(5754));
    layer1_outputs(6854) <= layer0_outputs(5668);
    layer1_outputs(6855) <= layer0_outputs(2204);
    layer1_outputs(6856) <= '1';
    layer1_outputs(6857) <= layer0_outputs(5935);
    layer1_outputs(6858) <= not(layer0_outputs(4060));
    layer1_outputs(6859) <= not(layer0_outputs(5871));
    layer1_outputs(6860) <= not((layer0_outputs(5227)) and (layer0_outputs(6627)));
    layer1_outputs(6861) <= '0';
    layer1_outputs(6862) <= layer0_outputs(7281);
    layer1_outputs(6863) <= not((layer0_outputs(1388)) xor (layer0_outputs(3311)));
    layer1_outputs(6864) <= not(layer0_outputs(1535));
    layer1_outputs(6865) <= not(layer0_outputs(595));
    layer1_outputs(6866) <= not(layer0_outputs(4077));
    layer1_outputs(6867) <= not(layer0_outputs(6295));
    layer1_outputs(6868) <= layer0_outputs(770);
    layer1_outputs(6869) <= not(layer0_outputs(2534)) or (layer0_outputs(1832));
    layer1_outputs(6870) <= (layer0_outputs(3107)) or (layer0_outputs(923));
    layer1_outputs(6871) <= layer0_outputs(625);
    layer1_outputs(6872) <= (layer0_outputs(2707)) and not (layer0_outputs(4540));
    layer1_outputs(6873) <= layer0_outputs(5215);
    layer1_outputs(6874) <= not(layer0_outputs(7417));
    layer1_outputs(6875) <= not((layer0_outputs(7369)) or (layer0_outputs(903)));
    layer1_outputs(6876) <= (layer0_outputs(2793)) and not (layer0_outputs(2107));
    layer1_outputs(6877) <= not(layer0_outputs(6777));
    layer1_outputs(6878) <= (layer0_outputs(2669)) and not (layer0_outputs(4473));
    layer1_outputs(6879) <= not(layer0_outputs(6474)) or (layer0_outputs(3388));
    layer1_outputs(6880) <= layer0_outputs(4588);
    layer1_outputs(6881) <= not((layer0_outputs(4825)) xor (layer0_outputs(3895)));
    layer1_outputs(6882) <= not(layer0_outputs(175));
    layer1_outputs(6883) <= not(layer0_outputs(3017)) or (layer0_outputs(5934));
    layer1_outputs(6884) <= (layer0_outputs(1869)) or (layer0_outputs(6960));
    layer1_outputs(6885) <= not(layer0_outputs(6767));
    layer1_outputs(6886) <= not(layer0_outputs(3949)) or (layer0_outputs(605));
    layer1_outputs(6887) <= '1';
    layer1_outputs(6888) <= not(layer0_outputs(5870)) or (layer0_outputs(5240));
    layer1_outputs(6889) <= '0';
    layer1_outputs(6890) <= not(layer0_outputs(5783)) or (layer0_outputs(7029));
    layer1_outputs(6891) <= (layer0_outputs(6031)) or (layer0_outputs(612));
    layer1_outputs(6892) <= layer0_outputs(6204);
    layer1_outputs(6893) <= (layer0_outputs(2575)) and not (layer0_outputs(5108));
    layer1_outputs(6894) <= not(layer0_outputs(287)) or (layer0_outputs(2914));
    layer1_outputs(6895) <= (layer0_outputs(3537)) or (layer0_outputs(4032));
    layer1_outputs(6896) <= '1';
    layer1_outputs(6897) <= (layer0_outputs(5710)) or (layer0_outputs(4260));
    layer1_outputs(6898) <= '0';
    layer1_outputs(6899) <= not(layer0_outputs(7288));
    layer1_outputs(6900) <= layer0_outputs(6533);
    layer1_outputs(6901) <= not(layer0_outputs(878));
    layer1_outputs(6902) <= not(layer0_outputs(2745)) or (layer0_outputs(983));
    layer1_outputs(6903) <= not((layer0_outputs(5851)) and (layer0_outputs(6526)));
    layer1_outputs(6904) <= '0';
    layer1_outputs(6905) <= layer0_outputs(5397);
    layer1_outputs(6906) <= layer0_outputs(2078);
    layer1_outputs(6907) <= not(layer0_outputs(6126)) or (layer0_outputs(2331));
    layer1_outputs(6908) <= (layer0_outputs(4133)) xor (layer0_outputs(170));
    layer1_outputs(6909) <= not((layer0_outputs(1799)) and (layer0_outputs(6756)));
    layer1_outputs(6910) <= layer0_outputs(3724);
    layer1_outputs(6911) <= layer0_outputs(878);
    layer1_outputs(6912) <= (layer0_outputs(6754)) or (layer0_outputs(3062));
    layer1_outputs(6913) <= not(layer0_outputs(3444)) or (layer0_outputs(282));
    layer1_outputs(6914) <= not(layer0_outputs(5674)) or (layer0_outputs(3580));
    layer1_outputs(6915) <= not(layer0_outputs(5856)) or (layer0_outputs(3817));
    layer1_outputs(6916) <= not((layer0_outputs(5326)) and (layer0_outputs(7394)));
    layer1_outputs(6917) <= not(layer0_outputs(1851));
    layer1_outputs(6918) <= layer0_outputs(21);
    layer1_outputs(6919) <= layer0_outputs(2078);
    layer1_outputs(6920) <= (layer0_outputs(2100)) and not (layer0_outputs(4898));
    layer1_outputs(6921) <= '1';
    layer1_outputs(6922) <= (layer0_outputs(4740)) and not (layer0_outputs(1156));
    layer1_outputs(6923) <= not(layer0_outputs(1736));
    layer1_outputs(6924) <= (layer0_outputs(6744)) or (layer0_outputs(5611));
    layer1_outputs(6925) <= (layer0_outputs(2423)) and (layer0_outputs(5332));
    layer1_outputs(6926) <= layer0_outputs(5202);
    layer1_outputs(6927) <= layer0_outputs(2716);
    layer1_outputs(6928) <= not(layer0_outputs(6165)) or (layer0_outputs(4182));
    layer1_outputs(6929) <= layer0_outputs(5810);
    layer1_outputs(6930) <= not((layer0_outputs(3709)) or (layer0_outputs(7671)));
    layer1_outputs(6931) <= (layer0_outputs(3818)) or (layer0_outputs(1871));
    layer1_outputs(6932) <= (layer0_outputs(2567)) or (layer0_outputs(7359));
    layer1_outputs(6933) <= '1';
    layer1_outputs(6934) <= layer0_outputs(4341);
    layer1_outputs(6935) <= '0';
    layer1_outputs(6936) <= not(layer0_outputs(5807));
    layer1_outputs(6937) <= layer0_outputs(340);
    layer1_outputs(6938) <= not((layer0_outputs(5602)) or (layer0_outputs(3913)));
    layer1_outputs(6939) <= not(layer0_outputs(4671));
    layer1_outputs(6940) <= not(layer0_outputs(5493));
    layer1_outputs(6941) <= not(layer0_outputs(6290)) or (layer0_outputs(5180));
    layer1_outputs(6942) <= not((layer0_outputs(6320)) xor (layer0_outputs(7569)));
    layer1_outputs(6943) <= '1';
    layer1_outputs(6944) <= layer0_outputs(467);
    layer1_outputs(6945) <= not((layer0_outputs(6213)) or (layer0_outputs(7195)));
    layer1_outputs(6946) <= not(layer0_outputs(4263));
    layer1_outputs(6947) <= not(layer0_outputs(5129)) or (layer0_outputs(3996));
    layer1_outputs(6948) <= not((layer0_outputs(5565)) and (layer0_outputs(6880)));
    layer1_outputs(6949) <= not(layer0_outputs(2561));
    layer1_outputs(6950) <= not(layer0_outputs(7444)) or (layer0_outputs(7625));
    layer1_outputs(6951) <= not(layer0_outputs(2338));
    layer1_outputs(6952) <= not(layer0_outputs(6877)) or (layer0_outputs(5333));
    layer1_outputs(6953) <= not(layer0_outputs(232));
    layer1_outputs(6954) <= '1';
    layer1_outputs(6955) <= layer0_outputs(4827);
    layer1_outputs(6956) <= not((layer0_outputs(727)) and (layer0_outputs(3451)));
    layer1_outputs(6957) <= (layer0_outputs(472)) and not (layer0_outputs(1113));
    layer1_outputs(6958) <= '1';
    layer1_outputs(6959) <= not(layer0_outputs(741));
    layer1_outputs(6960) <= (layer0_outputs(1687)) or (layer0_outputs(1459));
    layer1_outputs(6961) <= (layer0_outputs(7383)) or (layer0_outputs(6382));
    layer1_outputs(6962) <= (layer0_outputs(6932)) xor (layer0_outputs(5768));
    layer1_outputs(6963) <= layer0_outputs(1800);
    layer1_outputs(6964) <= (layer0_outputs(4557)) xor (layer0_outputs(5491));
    layer1_outputs(6965) <= (layer0_outputs(3672)) and not (layer0_outputs(2950));
    layer1_outputs(6966) <= (layer0_outputs(2751)) and not (layer0_outputs(689));
    layer1_outputs(6967) <= (layer0_outputs(6515)) and (layer0_outputs(2468));
    layer1_outputs(6968) <= (layer0_outputs(2068)) xor (layer0_outputs(4814));
    layer1_outputs(6969) <= layer0_outputs(6467);
    layer1_outputs(6970) <= layer0_outputs(1569);
    layer1_outputs(6971) <= (layer0_outputs(3715)) or (layer0_outputs(3225));
    layer1_outputs(6972) <= (layer0_outputs(6102)) or (layer0_outputs(3995));
    layer1_outputs(6973) <= not((layer0_outputs(2681)) or (layer0_outputs(196)));
    layer1_outputs(6974) <= '0';
    layer1_outputs(6975) <= not(layer0_outputs(7674));
    layer1_outputs(6976) <= (layer0_outputs(3457)) xor (layer0_outputs(5323));
    layer1_outputs(6977) <= (layer0_outputs(3690)) and not (layer0_outputs(6275));
    layer1_outputs(6978) <= not(layer0_outputs(2224)) or (layer0_outputs(410));
    layer1_outputs(6979) <= not(layer0_outputs(6923));
    layer1_outputs(6980) <= (layer0_outputs(4224)) and (layer0_outputs(3428));
    layer1_outputs(6981) <= not(layer0_outputs(722));
    layer1_outputs(6982) <= not(layer0_outputs(5479));
    layer1_outputs(6983) <= layer0_outputs(1619);
    layer1_outputs(6984) <= not((layer0_outputs(5592)) or (layer0_outputs(5376)));
    layer1_outputs(6985) <= (layer0_outputs(884)) or (layer0_outputs(2143));
    layer1_outputs(6986) <= (layer0_outputs(1193)) or (layer0_outputs(7126));
    layer1_outputs(6987) <= layer0_outputs(6192);
    layer1_outputs(6988) <= layer0_outputs(105);
    layer1_outputs(6989) <= (layer0_outputs(3277)) and not (layer0_outputs(1529));
    layer1_outputs(6990) <= (layer0_outputs(3447)) and (layer0_outputs(7036));
    layer1_outputs(6991) <= (layer0_outputs(630)) or (layer0_outputs(4281));
    layer1_outputs(6992) <= layer0_outputs(7032);
    layer1_outputs(6993) <= layer0_outputs(371);
    layer1_outputs(6994) <= '0';
    layer1_outputs(6995) <= not(layer0_outputs(4580)) or (layer0_outputs(5567));
    layer1_outputs(6996) <= '1';
    layer1_outputs(6997) <= not(layer0_outputs(4052)) or (layer0_outputs(909));
    layer1_outputs(6998) <= not(layer0_outputs(2670));
    layer1_outputs(6999) <= not(layer0_outputs(6920)) or (layer0_outputs(5480));
    layer1_outputs(7000) <= layer0_outputs(2548);
    layer1_outputs(7001) <= (layer0_outputs(3581)) xor (layer0_outputs(5877));
    layer1_outputs(7002) <= layer0_outputs(1038);
    layer1_outputs(7003) <= (layer0_outputs(1544)) and (layer0_outputs(6465));
    layer1_outputs(7004) <= not(layer0_outputs(6051)) or (layer0_outputs(1981));
    layer1_outputs(7005) <= not(layer0_outputs(1848)) or (layer0_outputs(2438));
    layer1_outputs(7006) <= '1';
    layer1_outputs(7007) <= layer0_outputs(5544);
    layer1_outputs(7008) <= not(layer0_outputs(1198));
    layer1_outputs(7009) <= (layer0_outputs(681)) or (layer0_outputs(6595));
    layer1_outputs(7010) <= (layer0_outputs(1457)) and not (layer0_outputs(7378));
    layer1_outputs(7011) <= not(layer0_outputs(1458));
    layer1_outputs(7012) <= (layer0_outputs(2897)) or (layer0_outputs(7595));
    layer1_outputs(7013) <= not(layer0_outputs(4927));
    layer1_outputs(7014) <= (layer0_outputs(2048)) and not (layer0_outputs(5341));
    layer1_outputs(7015) <= not(layer0_outputs(4148)) or (layer0_outputs(2962));
    layer1_outputs(7016) <= not((layer0_outputs(3042)) or (layer0_outputs(1899)));
    layer1_outputs(7017) <= not(layer0_outputs(580)) or (layer0_outputs(2136));
    layer1_outputs(7018) <= layer0_outputs(4915);
    layer1_outputs(7019) <= layer0_outputs(6983);
    layer1_outputs(7020) <= (layer0_outputs(667)) and not (layer0_outputs(4347));
    layer1_outputs(7021) <= layer0_outputs(2287);
    layer1_outputs(7022) <= (layer0_outputs(4865)) and not (layer0_outputs(3417));
    layer1_outputs(7023) <= (layer0_outputs(4782)) and not (layer0_outputs(2219));
    layer1_outputs(7024) <= not(layer0_outputs(3953)) or (layer0_outputs(6122));
    layer1_outputs(7025) <= layer0_outputs(198);
    layer1_outputs(7026) <= layer0_outputs(1825);
    layer1_outputs(7027) <= not(layer0_outputs(2422));
    layer1_outputs(7028) <= (layer0_outputs(5033)) and (layer0_outputs(5876));
    layer1_outputs(7029) <= '0';
    layer1_outputs(7030) <= not(layer0_outputs(4045));
    layer1_outputs(7031) <= not(layer0_outputs(2854)) or (layer0_outputs(2719));
    layer1_outputs(7032) <= layer0_outputs(7661);
    layer1_outputs(7033) <= layer0_outputs(1423);
    layer1_outputs(7034) <= not((layer0_outputs(4931)) and (layer0_outputs(1320)));
    layer1_outputs(7035) <= (layer0_outputs(1964)) and not (layer0_outputs(4522));
    layer1_outputs(7036) <= (layer0_outputs(2339)) and (layer0_outputs(2065));
    layer1_outputs(7037) <= (layer0_outputs(4975)) and not (layer0_outputs(930));
    layer1_outputs(7038) <= not((layer0_outputs(1484)) or (layer0_outputs(3527)));
    layer1_outputs(7039) <= not(layer0_outputs(2324));
    layer1_outputs(7040) <= not(layer0_outputs(3343));
    layer1_outputs(7041) <= (layer0_outputs(7187)) or (layer0_outputs(2446));
    layer1_outputs(7042) <= not(layer0_outputs(132)) or (layer0_outputs(619));
    layer1_outputs(7043) <= not(layer0_outputs(2787));
    layer1_outputs(7044) <= layer0_outputs(6220);
    layer1_outputs(7045) <= (layer0_outputs(4225)) or (layer0_outputs(4999));
    layer1_outputs(7046) <= (layer0_outputs(840)) and (layer0_outputs(7466));
    layer1_outputs(7047) <= layer0_outputs(683);
    layer1_outputs(7048) <= (layer0_outputs(5172)) and (layer0_outputs(4337));
    layer1_outputs(7049) <= not(layer0_outputs(604));
    layer1_outputs(7050) <= (layer0_outputs(1663)) and (layer0_outputs(1198));
    layer1_outputs(7051) <= (layer0_outputs(4219)) and not (layer0_outputs(894));
    layer1_outputs(7052) <= layer0_outputs(6722);
    layer1_outputs(7053) <= layer0_outputs(4254);
    layer1_outputs(7054) <= not(layer0_outputs(7291));
    layer1_outputs(7055) <= layer0_outputs(2969);
    layer1_outputs(7056) <= '0';
    layer1_outputs(7057) <= layer0_outputs(6497);
    layer1_outputs(7058) <= not((layer0_outputs(660)) or (layer0_outputs(619)));
    layer1_outputs(7059) <= (layer0_outputs(7597)) or (layer0_outputs(3432));
    layer1_outputs(7060) <= (layer0_outputs(3619)) and (layer0_outputs(784));
    layer1_outputs(7061) <= not((layer0_outputs(551)) and (layer0_outputs(1646)));
    layer1_outputs(7062) <= not(layer0_outputs(742)) or (layer0_outputs(3117));
    layer1_outputs(7063) <= (layer0_outputs(648)) or (layer0_outputs(4822));
    layer1_outputs(7064) <= layer0_outputs(6590);
    layer1_outputs(7065) <= layer0_outputs(690);
    layer1_outputs(7066) <= not(layer0_outputs(7369));
    layer1_outputs(7067) <= (layer0_outputs(7287)) and (layer0_outputs(6339));
    layer1_outputs(7068) <= not((layer0_outputs(4625)) and (layer0_outputs(7392)));
    layer1_outputs(7069) <= not(layer0_outputs(1486));
    layer1_outputs(7070) <= not(layer0_outputs(2804)) or (layer0_outputs(2727));
    layer1_outputs(7071) <= (layer0_outputs(1538)) and (layer0_outputs(5896));
    layer1_outputs(7072) <= not(layer0_outputs(5755));
    layer1_outputs(7073) <= not(layer0_outputs(4645)) or (layer0_outputs(5101));
    layer1_outputs(7074) <= not((layer0_outputs(2722)) and (layer0_outputs(5700)));
    layer1_outputs(7075) <= not(layer0_outputs(4539));
    layer1_outputs(7076) <= (layer0_outputs(4370)) and (layer0_outputs(1482));
    layer1_outputs(7077) <= layer0_outputs(4399);
    layer1_outputs(7078) <= not((layer0_outputs(7000)) or (layer0_outputs(324)));
    layer1_outputs(7079) <= not(layer0_outputs(2121));
    layer1_outputs(7080) <= not((layer0_outputs(1933)) and (layer0_outputs(1894)));
    layer1_outputs(7081) <= (layer0_outputs(7421)) or (layer0_outputs(3862));
    layer1_outputs(7082) <= layer0_outputs(7175);
    layer1_outputs(7083) <= not(layer0_outputs(7254));
    layer1_outputs(7084) <= layer0_outputs(6227);
    layer1_outputs(7085) <= not(layer0_outputs(488)) or (layer0_outputs(3568));
    layer1_outputs(7086) <= (layer0_outputs(2017)) and (layer0_outputs(7033));
    layer1_outputs(7087) <= (layer0_outputs(5348)) and (layer0_outputs(4802));
    layer1_outputs(7088) <= (layer0_outputs(4151)) and not (layer0_outputs(4860));
    layer1_outputs(7089) <= (layer0_outputs(980)) and not (layer0_outputs(7510));
    layer1_outputs(7090) <= (layer0_outputs(1729)) and (layer0_outputs(6058));
    layer1_outputs(7091) <= not(layer0_outputs(7601));
    layer1_outputs(7092) <= layer0_outputs(1768);
    layer1_outputs(7093) <= layer0_outputs(6811);
    layer1_outputs(7094) <= (layer0_outputs(623)) and not (layer0_outputs(121));
    layer1_outputs(7095) <= not((layer0_outputs(1779)) and (layer0_outputs(1492)));
    layer1_outputs(7096) <= layer0_outputs(6709);
    layer1_outputs(7097) <= not(layer0_outputs(1034));
    layer1_outputs(7098) <= not(layer0_outputs(3420));
    layer1_outputs(7099) <= (layer0_outputs(6899)) or (layer0_outputs(7278));
    layer1_outputs(7100) <= layer0_outputs(1601);
    layer1_outputs(7101) <= layer0_outputs(7486);
    layer1_outputs(7102) <= not((layer0_outputs(7197)) or (layer0_outputs(7307)));
    layer1_outputs(7103) <= (layer0_outputs(5682)) and (layer0_outputs(5102));
    layer1_outputs(7104) <= (layer0_outputs(521)) and not (layer0_outputs(5617));
    layer1_outputs(7105) <= not((layer0_outputs(2389)) or (layer0_outputs(3157)));
    layer1_outputs(7106) <= not((layer0_outputs(7653)) or (layer0_outputs(3874)));
    layer1_outputs(7107) <= not(layer0_outputs(550));
    layer1_outputs(7108) <= '1';
    layer1_outputs(7109) <= not(layer0_outputs(1963));
    layer1_outputs(7110) <= (layer0_outputs(6581)) or (layer0_outputs(1038));
    layer1_outputs(7111) <= not((layer0_outputs(5690)) or (layer0_outputs(5658)));
    layer1_outputs(7112) <= layer0_outputs(6829);
    layer1_outputs(7113) <= (layer0_outputs(6241)) and (layer0_outputs(3876));
    layer1_outputs(7114) <= layer0_outputs(7458);
    layer1_outputs(7115) <= (layer0_outputs(2023)) or (layer0_outputs(6219));
    layer1_outputs(7116) <= '1';
    layer1_outputs(7117) <= '1';
    layer1_outputs(7118) <= layer0_outputs(3093);
    layer1_outputs(7119) <= (layer0_outputs(7356)) and not (layer0_outputs(392));
    layer1_outputs(7120) <= (layer0_outputs(7217)) xor (layer0_outputs(121));
    layer1_outputs(7121) <= (layer0_outputs(2835)) and not (layer0_outputs(3232));
    layer1_outputs(7122) <= layer0_outputs(5708);
    layer1_outputs(7123) <= not((layer0_outputs(1288)) or (layer0_outputs(4979)));
    layer1_outputs(7124) <= '1';
    layer1_outputs(7125) <= layer0_outputs(1080);
    layer1_outputs(7126) <= '1';
    layer1_outputs(7127) <= not((layer0_outputs(7368)) and (layer0_outputs(5990)));
    layer1_outputs(7128) <= not(layer0_outputs(1994));
    layer1_outputs(7129) <= not((layer0_outputs(5401)) or (layer0_outputs(691)));
    layer1_outputs(7130) <= not(layer0_outputs(2855)) or (layer0_outputs(4221));
    layer1_outputs(7131) <= '0';
    layer1_outputs(7132) <= layer0_outputs(4949);
    layer1_outputs(7133) <= not(layer0_outputs(2944)) or (layer0_outputs(2888));
    layer1_outputs(7134) <= not(layer0_outputs(7112)) or (layer0_outputs(1950));
    layer1_outputs(7135) <= not(layer0_outputs(6766));
    layer1_outputs(7136) <= not(layer0_outputs(1982));
    layer1_outputs(7137) <= (layer0_outputs(4135)) or (layer0_outputs(7474));
    layer1_outputs(7138) <= not(layer0_outputs(2001));
    layer1_outputs(7139) <= (layer0_outputs(293)) and not (layer0_outputs(6233));
    layer1_outputs(7140) <= (layer0_outputs(5127)) and not (layer0_outputs(6737));
    layer1_outputs(7141) <= layer0_outputs(6570);
    layer1_outputs(7142) <= not(layer0_outputs(3894));
    layer1_outputs(7143) <= not((layer0_outputs(4303)) and (layer0_outputs(5560)));
    layer1_outputs(7144) <= (layer0_outputs(95)) or (layer0_outputs(2530));
    layer1_outputs(7145) <= layer0_outputs(6456);
    layer1_outputs(7146) <= layer0_outputs(7483);
    layer1_outputs(7147) <= not((layer0_outputs(1153)) or (layer0_outputs(3835)));
    layer1_outputs(7148) <= not(layer0_outputs(2470));
    layer1_outputs(7149) <= layer0_outputs(3795);
    layer1_outputs(7150) <= (layer0_outputs(4678)) and not (layer0_outputs(3972));
    layer1_outputs(7151) <= not((layer0_outputs(1066)) and (layer0_outputs(3704)));
    layer1_outputs(7152) <= not((layer0_outputs(3871)) and (layer0_outputs(895)));
    layer1_outputs(7153) <= (layer0_outputs(4752)) and (layer0_outputs(2258));
    layer1_outputs(7154) <= not(layer0_outputs(2856)) or (layer0_outputs(6850));
    layer1_outputs(7155) <= not(layer0_outputs(4114)) or (layer0_outputs(3041));
    layer1_outputs(7156) <= not(layer0_outputs(290));
    layer1_outputs(7157) <= (layer0_outputs(4008)) and not (layer0_outputs(6576));
    layer1_outputs(7158) <= not(layer0_outputs(621));
    layer1_outputs(7159) <= not(layer0_outputs(6133)) or (layer0_outputs(3564));
    layer1_outputs(7160) <= (layer0_outputs(3614)) or (layer0_outputs(4006));
    layer1_outputs(7161) <= layer0_outputs(2572);
    layer1_outputs(7162) <= (layer0_outputs(2548)) and not (layer0_outputs(3861));
    layer1_outputs(7163) <= not(layer0_outputs(5319));
    layer1_outputs(7164) <= not((layer0_outputs(2140)) and (layer0_outputs(6002)));
    layer1_outputs(7165) <= not((layer0_outputs(1360)) or (layer0_outputs(7396)));
    layer1_outputs(7166) <= not(layer0_outputs(494)) or (layer0_outputs(4446));
    layer1_outputs(7167) <= (layer0_outputs(7189)) and (layer0_outputs(2868));
    layer1_outputs(7168) <= not(layer0_outputs(505)) or (layer0_outputs(4995));
    layer1_outputs(7169) <= not(layer0_outputs(246)) or (layer0_outputs(6281));
    layer1_outputs(7170) <= layer0_outputs(7089);
    layer1_outputs(7171) <= not(layer0_outputs(7218));
    layer1_outputs(7172) <= '1';
    layer1_outputs(7173) <= layer0_outputs(4231);
    layer1_outputs(7174) <= layer0_outputs(6417);
    layer1_outputs(7175) <= (layer0_outputs(6272)) and not (layer0_outputs(3572));
    layer1_outputs(7176) <= '0';
    layer1_outputs(7177) <= layer0_outputs(1343);
    layer1_outputs(7178) <= (layer0_outputs(3169)) and not (layer0_outputs(4545));
    layer1_outputs(7179) <= layer0_outputs(4515);
    layer1_outputs(7180) <= '0';
    layer1_outputs(7181) <= layer0_outputs(2995);
    layer1_outputs(7182) <= layer0_outputs(1403);
    layer1_outputs(7183) <= not((layer0_outputs(411)) or (layer0_outputs(4643)));
    layer1_outputs(7184) <= layer0_outputs(7612);
    layer1_outputs(7185) <= (layer0_outputs(3468)) or (layer0_outputs(2202));
    layer1_outputs(7186) <= (layer0_outputs(747)) and not (layer0_outputs(3958));
    layer1_outputs(7187) <= '0';
    layer1_outputs(7188) <= not(layer0_outputs(6993));
    layer1_outputs(7189) <= layer0_outputs(3007);
    layer1_outputs(7190) <= (layer0_outputs(1410)) and not (layer0_outputs(7278));
    layer1_outputs(7191) <= not((layer0_outputs(7178)) and (layer0_outputs(7319)));
    layer1_outputs(7192) <= not(layer0_outputs(167));
    layer1_outputs(7193) <= (layer0_outputs(6103)) and not (layer0_outputs(2343));
    layer1_outputs(7194) <= (layer0_outputs(1600)) or (layer0_outputs(5861));
    layer1_outputs(7195) <= layer0_outputs(1453);
    layer1_outputs(7196) <= layer0_outputs(5049);
    layer1_outputs(7197) <= layer0_outputs(7204);
    layer1_outputs(7198) <= not(layer0_outputs(2261));
    layer1_outputs(7199) <= not((layer0_outputs(5928)) xor (layer0_outputs(2341)));
    layer1_outputs(7200) <= not((layer0_outputs(6618)) or (layer0_outputs(2864)));
    layer1_outputs(7201) <= not((layer0_outputs(3116)) and (layer0_outputs(2511)));
    layer1_outputs(7202) <= '0';
    layer1_outputs(7203) <= not(layer0_outputs(6964));
    layer1_outputs(7204) <= (layer0_outputs(3340)) or (layer0_outputs(3427));
    layer1_outputs(7205) <= layer0_outputs(89);
    layer1_outputs(7206) <= not(layer0_outputs(4874));
    layer1_outputs(7207) <= not(layer0_outputs(7623)) or (layer0_outputs(3899));
    layer1_outputs(7208) <= (layer0_outputs(1807)) and (layer0_outputs(6577));
    layer1_outputs(7209) <= not((layer0_outputs(3229)) or (layer0_outputs(1072)));
    layer1_outputs(7210) <= layer0_outputs(923);
    layer1_outputs(7211) <= not(layer0_outputs(5420));
    layer1_outputs(7212) <= (layer0_outputs(3384)) or (layer0_outputs(2422));
    layer1_outputs(7213) <= '0';
    layer1_outputs(7214) <= not(layer0_outputs(2964)) or (layer0_outputs(2098));
    layer1_outputs(7215) <= (layer0_outputs(1685)) xor (layer0_outputs(5843));
    layer1_outputs(7216) <= (layer0_outputs(1595)) and not (layer0_outputs(801));
    layer1_outputs(7217) <= not(layer0_outputs(1872));
    layer1_outputs(7218) <= not(layer0_outputs(2444));
    layer1_outputs(7219) <= layer0_outputs(173);
    layer1_outputs(7220) <= (layer0_outputs(3151)) or (layer0_outputs(3784));
    layer1_outputs(7221) <= not(layer0_outputs(7426));
    layer1_outputs(7222) <= not(layer0_outputs(1896));
    layer1_outputs(7223) <= (layer0_outputs(1320)) and (layer0_outputs(3285));
    layer1_outputs(7224) <= not((layer0_outputs(6975)) or (layer0_outputs(5263)));
    layer1_outputs(7225) <= not(layer0_outputs(5779)) or (layer0_outputs(5160));
    layer1_outputs(7226) <= not((layer0_outputs(2617)) or (layer0_outputs(1377)));
    layer1_outputs(7227) <= layer0_outputs(3353);
    layer1_outputs(7228) <= layer0_outputs(3020);
    layer1_outputs(7229) <= not(layer0_outputs(2008)) or (layer0_outputs(2915));
    layer1_outputs(7230) <= not((layer0_outputs(5791)) or (layer0_outputs(6958)));
    layer1_outputs(7231) <= (layer0_outputs(4853)) and not (layer0_outputs(3239));
    layer1_outputs(7232) <= not((layer0_outputs(2906)) or (layer0_outputs(4312)));
    layer1_outputs(7233) <= layer0_outputs(2319);
    layer1_outputs(7234) <= layer0_outputs(6188);
    layer1_outputs(7235) <= not((layer0_outputs(4483)) xor (layer0_outputs(489)));
    layer1_outputs(7236) <= (layer0_outputs(4309)) or (layer0_outputs(644));
    layer1_outputs(7237) <= (layer0_outputs(5130)) or (layer0_outputs(5085));
    layer1_outputs(7238) <= layer0_outputs(6607);
    layer1_outputs(7239) <= '0';
    layer1_outputs(7240) <= not(layer0_outputs(7525));
    layer1_outputs(7241) <= (layer0_outputs(2374)) or (layer0_outputs(317));
    layer1_outputs(7242) <= not(layer0_outputs(2393)) or (layer0_outputs(7342));
    layer1_outputs(7243) <= (layer0_outputs(2052)) and (layer0_outputs(1982));
    layer1_outputs(7244) <= not(layer0_outputs(2170)) or (layer0_outputs(7368));
    layer1_outputs(7245) <= (layer0_outputs(100)) and (layer0_outputs(2860));
    layer1_outputs(7246) <= layer0_outputs(5578);
    layer1_outputs(7247) <= layer0_outputs(659);
    layer1_outputs(7248) <= not(layer0_outputs(5300)) or (layer0_outputs(6881));
    layer1_outputs(7249) <= (layer0_outputs(6430)) and not (layer0_outputs(5018));
    layer1_outputs(7250) <= '0';
    layer1_outputs(7251) <= not(layer0_outputs(2722));
    layer1_outputs(7252) <= (layer0_outputs(2592)) or (layer0_outputs(4657));
    layer1_outputs(7253) <= layer0_outputs(4710);
    layer1_outputs(7254) <= not(layer0_outputs(5664)) or (layer0_outputs(4013));
    layer1_outputs(7255) <= not(layer0_outputs(5399)) or (layer0_outputs(4871));
    layer1_outputs(7256) <= not((layer0_outputs(4436)) xor (layer0_outputs(3816)));
    layer1_outputs(7257) <= (layer0_outputs(1075)) and not (layer0_outputs(4753));
    layer1_outputs(7258) <= (layer0_outputs(93)) or (layer0_outputs(3125));
    layer1_outputs(7259) <= not(layer0_outputs(6278));
    layer1_outputs(7260) <= '1';
    layer1_outputs(7261) <= (layer0_outputs(5605)) and not (layer0_outputs(5948));
    layer1_outputs(7262) <= (layer0_outputs(5001)) and (layer0_outputs(7653));
    layer1_outputs(7263) <= layer0_outputs(4061);
    layer1_outputs(7264) <= not(layer0_outputs(2388)) or (layer0_outputs(5515));
    layer1_outputs(7265) <= not(layer0_outputs(3449));
    layer1_outputs(7266) <= (layer0_outputs(7238)) or (layer0_outputs(5628));
    layer1_outputs(7267) <= (layer0_outputs(114)) and not (layer0_outputs(3780));
    layer1_outputs(7268) <= not((layer0_outputs(150)) and (layer0_outputs(2524)));
    layer1_outputs(7269) <= (layer0_outputs(650)) and not (layer0_outputs(916));
    layer1_outputs(7270) <= not(layer0_outputs(2676)) or (layer0_outputs(2616));
    layer1_outputs(7271) <= layer0_outputs(3639);
    layer1_outputs(7272) <= not(layer0_outputs(3492)) or (layer0_outputs(2021));
    layer1_outputs(7273) <= not(layer0_outputs(5778));
    layer1_outputs(7274) <= layer0_outputs(1022);
    layer1_outputs(7275) <= (layer0_outputs(1117)) or (layer0_outputs(5110));
    layer1_outputs(7276) <= layer0_outputs(7204);
    layer1_outputs(7277) <= not(layer0_outputs(4562));
    layer1_outputs(7278) <= (layer0_outputs(6491)) and (layer0_outputs(1622));
    layer1_outputs(7279) <= (layer0_outputs(1346)) and not (layer0_outputs(7363));
    layer1_outputs(7280) <= (layer0_outputs(3084)) and not (layer0_outputs(4015));
    layer1_outputs(7281) <= not((layer0_outputs(931)) or (layer0_outputs(2632)));
    layer1_outputs(7282) <= not((layer0_outputs(1672)) or (layer0_outputs(2328)));
    layer1_outputs(7283) <= not((layer0_outputs(6207)) and (layer0_outputs(4721)));
    layer1_outputs(7284) <= not((layer0_outputs(2223)) xor (layer0_outputs(6561)));
    layer1_outputs(7285) <= not((layer0_outputs(6705)) xor (layer0_outputs(1523)));
    layer1_outputs(7286) <= (layer0_outputs(4315)) or (layer0_outputs(301));
    layer1_outputs(7287) <= not(layer0_outputs(2317)) or (layer0_outputs(1845));
    layer1_outputs(7288) <= '1';
    layer1_outputs(7289) <= (layer0_outputs(469)) and not (layer0_outputs(2691));
    layer1_outputs(7290) <= not(layer0_outputs(179)) or (layer0_outputs(7165));
    layer1_outputs(7291) <= (layer0_outputs(5267)) or (layer0_outputs(4831));
    layer1_outputs(7292) <= not(layer0_outputs(2033));
    layer1_outputs(7293) <= (layer0_outputs(2329)) and not (layer0_outputs(6653));
    layer1_outputs(7294) <= (layer0_outputs(279)) or (layer0_outputs(1959));
    layer1_outputs(7295) <= not((layer0_outputs(1491)) and (layer0_outputs(3627)));
    layer1_outputs(7296) <= layer0_outputs(5925);
    layer1_outputs(7297) <= (layer0_outputs(3347)) and not (layer0_outputs(3103));
    layer1_outputs(7298) <= (layer0_outputs(5819)) or (layer0_outputs(7193));
    layer1_outputs(7299) <= not((layer0_outputs(1418)) and (layer0_outputs(2318)));
    layer1_outputs(7300) <= '1';
    layer1_outputs(7301) <= layer0_outputs(1852);
    layer1_outputs(7302) <= not(layer0_outputs(6747));
    layer1_outputs(7303) <= not(layer0_outputs(766));
    layer1_outputs(7304) <= (layer0_outputs(3612)) or (layer0_outputs(84));
    layer1_outputs(7305) <= not((layer0_outputs(4747)) and (layer0_outputs(6301)));
    layer1_outputs(7306) <= (layer0_outputs(6872)) and not (layer0_outputs(2256));
    layer1_outputs(7307) <= (layer0_outputs(3297)) and not (layer0_outputs(3620));
    layer1_outputs(7308) <= not((layer0_outputs(5322)) and (layer0_outputs(3381)));
    layer1_outputs(7309) <= not((layer0_outputs(5489)) and (layer0_outputs(3886)));
    layer1_outputs(7310) <= not(layer0_outputs(2026));
    layer1_outputs(7311) <= not((layer0_outputs(1127)) and (layer0_outputs(2132)));
    layer1_outputs(7312) <= '0';
    layer1_outputs(7313) <= layer0_outputs(3747);
    layer1_outputs(7314) <= not(layer0_outputs(6141));
    layer1_outputs(7315) <= layer0_outputs(2323);
    layer1_outputs(7316) <= (layer0_outputs(3241)) and not (layer0_outputs(3904));
    layer1_outputs(7317) <= '1';
    layer1_outputs(7318) <= not(layer0_outputs(5306));
    layer1_outputs(7319) <= (layer0_outputs(579)) and not (layer0_outputs(3268));
    layer1_outputs(7320) <= not(layer0_outputs(1171));
    layer1_outputs(7321) <= not(layer0_outputs(1325));
    layer1_outputs(7322) <= (layer0_outputs(4083)) and not (layer0_outputs(1192));
    layer1_outputs(7323) <= not((layer0_outputs(1734)) and (layer0_outputs(6321)));
    layer1_outputs(7324) <= not(layer0_outputs(2558));
    layer1_outputs(7325) <= '0';
    layer1_outputs(7326) <= (layer0_outputs(2806)) or (layer0_outputs(2555));
    layer1_outputs(7327) <= layer0_outputs(2718);
    layer1_outputs(7328) <= (layer0_outputs(3213)) or (layer0_outputs(18));
    layer1_outputs(7329) <= layer0_outputs(2780);
    layer1_outputs(7330) <= not(layer0_outputs(856));
    layer1_outputs(7331) <= (layer0_outputs(4819)) and not (layer0_outputs(2297));
    layer1_outputs(7332) <= not((layer0_outputs(5513)) xor (layer0_outputs(5369)));
    layer1_outputs(7333) <= (layer0_outputs(3408)) and not (layer0_outputs(4960));
    layer1_outputs(7334) <= not((layer0_outputs(4728)) and (layer0_outputs(197)));
    layer1_outputs(7335) <= not((layer0_outputs(7449)) and (layer0_outputs(4707)));
    layer1_outputs(7336) <= not(layer0_outputs(4722));
    layer1_outputs(7337) <= layer0_outputs(7021);
    layer1_outputs(7338) <= not((layer0_outputs(6929)) and (layer0_outputs(3080)));
    layer1_outputs(7339) <= not(layer0_outputs(1304)) or (layer0_outputs(3771));
    layer1_outputs(7340) <= (layer0_outputs(306)) and not (layer0_outputs(807));
    layer1_outputs(7341) <= layer0_outputs(1791);
    layer1_outputs(7342) <= layer0_outputs(6835);
    layer1_outputs(7343) <= (layer0_outputs(14)) and (layer0_outputs(7364));
    layer1_outputs(7344) <= (layer0_outputs(5708)) or (layer0_outputs(6804));
    layer1_outputs(7345) <= (layer0_outputs(7613)) and not (layer0_outputs(1707));
    layer1_outputs(7346) <= (layer0_outputs(4437)) or (layer0_outputs(2133));
    layer1_outputs(7347) <= (layer0_outputs(6450)) and not (layer0_outputs(905));
    layer1_outputs(7348) <= layer0_outputs(6302);
    layer1_outputs(7349) <= '1';
    layer1_outputs(7350) <= not((layer0_outputs(2061)) or (layer0_outputs(1849)));
    layer1_outputs(7351) <= not(layer0_outputs(6865)) or (layer0_outputs(6229));
    layer1_outputs(7352) <= (layer0_outputs(5385)) and (layer0_outputs(4971));
    layer1_outputs(7353) <= not(layer0_outputs(4322));
    layer1_outputs(7354) <= (layer0_outputs(3692)) and not (layer0_outputs(6553));
    layer1_outputs(7355) <= not((layer0_outputs(506)) xor (layer0_outputs(7301)));
    layer1_outputs(7356) <= '0';
    layer1_outputs(7357) <= layer0_outputs(4042);
    layer1_outputs(7358) <= (layer0_outputs(1413)) or (layer0_outputs(860));
    layer1_outputs(7359) <= not((layer0_outputs(1453)) or (layer0_outputs(4296)));
    layer1_outputs(7360) <= layer0_outputs(5382);
    layer1_outputs(7361) <= '1';
    layer1_outputs(7362) <= not(layer0_outputs(6424));
    layer1_outputs(7363) <= layer0_outputs(3314);
    layer1_outputs(7364) <= not(layer0_outputs(4815));
    layer1_outputs(7365) <= not(layer0_outputs(3291)) or (layer0_outputs(7642));
    layer1_outputs(7366) <= (layer0_outputs(2036)) and not (layer0_outputs(6418));
    layer1_outputs(7367) <= layer0_outputs(2864);
    layer1_outputs(7368) <= (layer0_outputs(2735)) and not (layer0_outputs(4533));
    layer1_outputs(7369) <= (layer0_outputs(1516)) and (layer0_outputs(2071));
    layer1_outputs(7370) <= not((layer0_outputs(1774)) and (layer0_outputs(4813)));
    layer1_outputs(7371) <= layer0_outputs(3934);
    layer1_outputs(7372) <= not(layer0_outputs(3496));
    layer1_outputs(7373) <= not(layer0_outputs(6953));
    layer1_outputs(7374) <= (layer0_outputs(4384)) or (layer0_outputs(1519));
    layer1_outputs(7375) <= not(layer0_outputs(7437));
    layer1_outputs(7376) <= (layer0_outputs(2775)) and (layer0_outputs(4568));
    layer1_outputs(7377) <= (layer0_outputs(1725)) and not (layer0_outputs(5114));
    layer1_outputs(7378) <= (layer0_outputs(3547)) or (layer0_outputs(2520));
    layer1_outputs(7379) <= not(layer0_outputs(5162)) or (layer0_outputs(5026));
    layer1_outputs(7380) <= not((layer0_outputs(7294)) and (layer0_outputs(2375)));
    layer1_outputs(7381) <= not((layer0_outputs(6600)) and (layer0_outputs(5957)));
    layer1_outputs(7382) <= not(layer0_outputs(4707));
    layer1_outputs(7383) <= '1';
    layer1_outputs(7384) <= not((layer0_outputs(2377)) and (layer0_outputs(1547)));
    layer1_outputs(7385) <= not(layer0_outputs(5681)) or (layer0_outputs(1260));
    layer1_outputs(7386) <= (layer0_outputs(5550)) or (layer0_outputs(280));
    layer1_outputs(7387) <= '1';
    layer1_outputs(7388) <= layer0_outputs(2657);
    layer1_outputs(7389) <= (layer0_outputs(6075)) or (layer0_outputs(3522));
    layer1_outputs(7390) <= not((layer0_outputs(3596)) and (layer0_outputs(3682)));
    layer1_outputs(7391) <= (layer0_outputs(6200)) and not (layer0_outputs(2866));
    layer1_outputs(7392) <= not(layer0_outputs(1818)) or (layer0_outputs(7535));
    layer1_outputs(7393) <= (layer0_outputs(4853)) or (layer0_outputs(3076));
    layer1_outputs(7394) <= not(layer0_outputs(6079));
    layer1_outputs(7395) <= '0';
    layer1_outputs(7396) <= layer0_outputs(6259);
    layer1_outputs(7397) <= not(layer0_outputs(733)) or (layer0_outputs(4245));
    layer1_outputs(7398) <= not((layer0_outputs(7141)) and (layer0_outputs(7241)));
    layer1_outputs(7399) <= not(layer0_outputs(2378));
    layer1_outputs(7400) <= layer0_outputs(893);
    layer1_outputs(7401) <= not(layer0_outputs(5311));
    layer1_outputs(7402) <= not(layer0_outputs(1344));
    layer1_outputs(7403) <= not((layer0_outputs(5335)) or (layer0_outputs(3480)));
    layer1_outputs(7404) <= not(layer0_outputs(4699));
    layer1_outputs(7405) <= layer0_outputs(5484);
    layer1_outputs(7406) <= layer0_outputs(5897);
    layer1_outputs(7407) <= (layer0_outputs(1866)) or (layer0_outputs(1835));
    layer1_outputs(7408) <= '0';
    layer1_outputs(7409) <= '1';
    layer1_outputs(7410) <= not(layer0_outputs(3857)) or (layer0_outputs(4408));
    layer1_outputs(7411) <= not(layer0_outputs(2649)) or (layer0_outputs(3033));
    layer1_outputs(7412) <= not((layer0_outputs(397)) and (layer0_outputs(7104)));
    layer1_outputs(7413) <= (layer0_outputs(4098)) and not (layer0_outputs(526));
    layer1_outputs(7414) <= not(layer0_outputs(7220));
    layer1_outputs(7415) <= (layer0_outputs(5672)) and (layer0_outputs(760));
    layer1_outputs(7416) <= not((layer0_outputs(4630)) or (layer0_outputs(5752)));
    layer1_outputs(7417) <= '1';
    layer1_outputs(7418) <= (layer0_outputs(2832)) and not (layer0_outputs(7179));
    layer1_outputs(7419) <= layer0_outputs(4725);
    layer1_outputs(7420) <= not(layer0_outputs(1209)) or (layer0_outputs(3765));
    layer1_outputs(7421) <= (layer0_outputs(53)) or (layer0_outputs(5291));
    layer1_outputs(7422) <= not(layer0_outputs(6547));
    layer1_outputs(7423) <= layer0_outputs(5155);
    layer1_outputs(7424) <= '1';
    layer1_outputs(7425) <= (layer0_outputs(5273)) or (layer0_outputs(5481));
    layer1_outputs(7426) <= not(layer0_outputs(5598));
    layer1_outputs(7427) <= not(layer0_outputs(7250));
    layer1_outputs(7428) <= not(layer0_outputs(5610));
    layer1_outputs(7429) <= not(layer0_outputs(7122)) or (layer0_outputs(4154));
    layer1_outputs(7430) <= not(layer0_outputs(4332)) or (layer0_outputs(3495));
    layer1_outputs(7431) <= (layer0_outputs(3390)) or (layer0_outputs(3445));
    layer1_outputs(7432) <= not((layer0_outputs(5356)) or (layer0_outputs(6088)));
    layer1_outputs(7433) <= '1';
    layer1_outputs(7434) <= not(layer0_outputs(6210));
    layer1_outputs(7435) <= layer0_outputs(2253);
    layer1_outputs(7436) <= not((layer0_outputs(4134)) and (layer0_outputs(3694)));
    layer1_outputs(7437) <= not(layer0_outputs(1655)) or (layer0_outputs(4334));
    layer1_outputs(7438) <= not(layer0_outputs(1400));
    layer1_outputs(7439) <= not(layer0_outputs(1180)) or (layer0_outputs(311));
    layer1_outputs(7440) <= layer0_outputs(1127);
    layer1_outputs(7441) <= (layer0_outputs(4504)) and (layer0_outputs(6344));
    layer1_outputs(7442) <= not(layer0_outputs(6508));
    layer1_outputs(7443) <= (layer0_outputs(4820)) and not (layer0_outputs(6813));
    layer1_outputs(7444) <= layer0_outputs(1660);
    layer1_outputs(7445) <= not(layer0_outputs(810));
    layer1_outputs(7446) <= '0';
    layer1_outputs(7447) <= (layer0_outputs(7428)) and not (layer0_outputs(7156));
    layer1_outputs(7448) <= (layer0_outputs(4009)) or (layer0_outputs(5752));
    layer1_outputs(7449) <= not(layer0_outputs(1579)) or (layer0_outputs(6381));
    layer1_outputs(7450) <= '1';
    layer1_outputs(7451) <= layer0_outputs(751);
    layer1_outputs(7452) <= '0';
    layer1_outputs(7453) <= not((layer0_outputs(4992)) and (layer0_outputs(1237)));
    layer1_outputs(7454) <= layer0_outputs(4160);
    layer1_outputs(7455) <= layer0_outputs(7028);
    layer1_outputs(7456) <= not((layer0_outputs(6724)) and (layer0_outputs(2256)));
    layer1_outputs(7457) <= not(layer0_outputs(3692)) or (layer0_outputs(4325));
    layer1_outputs(7458) <= not(layer0_outputs(222));
    layer1_outputs(7459) <= not(layer0_outputs(4434)) or (layer0_outputs(4462));
    layer1_outputs(7460) <= layer0_outputs(7666);
    layer1_outputs(7461) <= (layer0_outputs(4461)) and not (layer0_outputs(47));
    layer1_outputs(7462) <= not((layer0_outputs(1824)) and (layer0_outputs(5143)));
    layer1_outputs(7463) <= (layer0_outputs(1805)) and not (layer0_outputs(1444));
    layer1_outputs(7464) <= not(layer0_outputs(6974)) or (layer0_outputs(687));
    layer1_outputs(7465) <= '0';
    layer1_outputs(7466) <= (layer0_outputs(594)) and not (layer0_outputs(6332));
    layer1_outputs(7467) <= layer0_outputs(6672);
    layer1_outputs(7468) <= not(layer0_outputs(4278));
    layer1_outputs(7469) <= not(layer0_outputs(981)) or (layer0_outputs(2481));
    layer1_outputs(7470) <= not(layer0_outputs(524));
    layer1_outputs(7471) <= not((layer0_outputs(7126)) or (layer0_outputs(3456)));
    layer1_outputs(7472) <= not(layer0_outputs(3548));
    layer1_outputs(7473) <= not(layer0_outputs(3293));
    layer1_outputs(7474) <= layer0_outputs(834);
    layer1_outputs(7475) <= not((layer0_outputs(2724)) or (layer0_outputs(23)));
    layer1_outputs(7476) <= (layer0_outputs(2143)) and not (layer0_outputs(3121));
    layer1_outputs(7477) <= not((layer0_outputs(3439)) and (layer0_outputs(1165)));
    layer1_outputs(7478) <= (layer0_outputs(5247)) or (layer0_outputs(6453));
    layer1_outputs(7479) <= not((layer0_outputs(3910)) or (layer0_outputs(7358)));
    layer1_outputs(7480) <= not(layer0_outputs(7659)) or (layer0_outputs(6959));
    layer1_outputs(7481) <= not(layer0_outputs(3222)) or (layer0_outputs(1554));
    layer1_outputs(7482) <= (layer0_outputs(2266)) or (layer0_outputs(248));
    layer1_outputs(7483) <= not((layer0_outputs(670)) or (layer0_outputs(6844)));
    layer1_outputs(7484) <= '0';
    layer1_outputs(7485) <= not((layer0_outputs(1881)) or (layer0_outputs(5621)));
    layer1_outputs(7486) <= (layer0_outputs(6932)) and (layer0_outputs(6291));
    layer1_outputs(7487) <= not(layer0_outputs(5009));
    layer1_outputs(7488) <= layer0_outputs(4473);
    layer1_outputs(7489) <= not(layer0_outputs(6471));
    layer1_outputs(7490) <= not((layer0_outputs(7142)) and (layer0_outputs(7142)));
    layer1_outputs(7491) <= not(layer0_outputs(5855)) or (layer0_outputs(3624));
    layer1_outputs(7492) <= not(layer0_outputs(4080));
    layer1_outputs(7493) <= not((layer0_outputs(5098)) and (layer0_outputs(2124)));
    layer1_outputs(7494) <= layer0_outputs(2406);
    layer1_outputs(7495) <= not(layer0_outputs(4863));
    layer1_outputs(7496) <= not(layer0_outputs(2286));
    layer1_outputs(7497) <= (layer0_outputs(3230)) and not (layer0_outputs(3045));
    layer1_outputs(7498) <= layer0_outputs(5413);
    layer1_outputs(7499) <= not(layer0_outputs(3552)) or (layer0_outputs(1033));
    layer1_outputs(7500) <= (layer0_outputs(251)) or (layer0_outputs(2153));
    layer1_outputs(7501) <= not((layer0_outputs(5399)) and (layer0_outputs(6715)));
    layer1_outputs(7502) <= not(layer0_outputs(6227)) or (layer0_outputs(3732));
    layer1_outputs(7503) <= not(layer0_outputs(933)) or (layer0_outputs(1257));
    layer1_outputs(7504) <= not((layer0_outputs(672)) and (layer0_outputs(4210)));
    layer1_outputs(7505) <= not(layer0_outputs(7182)) or (layer0_outputs(1283));
    layer1_outputs(7506) <= '1';
    layer1_outputs(7507) <= (layer0_outputs(6358)) and not (layer0_outputs(1911));
    layer1_outputs(7508) <= not((layer0_outputs(969)) xor (layer0_outputs(2444)));
    layer1_outputs(7509) <= layer0_outputs(971);
    layer1_outputs(7510) <= not(layer0_outputs(2452));
    layer1_outputs(7511) <= not((layer0_outputs(6534)) xor (layer0_outputs(6161)));
    layer1_outputs(7512) <= not(layer0_outputs(5307)) or (layer0_outputs(5831));
    layer1_outputs(7513) <= (layer0_outputs(1652)) and (layer0_outputs(2905));
    layer1_outputs(7514) <= (layer0_outputs(548)) or (layer0_outputs(461));
    layer1_outputs(7515) <= not((layer0_outputs(5696)) and (layer0_outputs(5421)));
    layer1_outputs(7516) <= not((layer0_outputs(1326)) xor (layer0_outputs(7370)));
    layer1_outputs(7517) <= (layer0_outputs(4890)) and not (layer0_outputs(5713));
    layer1_outputs(7518) <= not((layer0_outputs(1209)) and (layer0_outputs(7341)));
    layer1_outputs(7519) <= (layer0_outputs(2399)) and (layer0_outputs(6549));
    layer1_outputs(7520) <= not((layer0_outputs(1167)) and (layer0_outputs(5772)));
    layer1_outputs(7521) <= not(layer0_outputs(6353)) or (layer0_outputs(1150));
    layer1_outputs(7522) <= not(layer0_outputs(2561));
    layer1_outputs(7523) <= (layer0_outputs(672)) xor (layer0_outputs(1809));
    layer1_outputs(7524) <= layer0_outputs(107);
    layer1_outputs(7525) <= not((layer0_outputs(831)) and (layer0_outputs(5242)));
    layer1_outputs(7526) <= (layer0_outputs(6620)) and (layer0_outputs(6629));
    layer1_outputs(7527) <= not(layer0_outputs(4316));
    layer1_outputs(7528) <= not(layer0_outputs(4941));
    layer1_outputs(7529) <= not(layer0_outputs(2173)) or (layer0_outputs(2266));
    layer1_outputs(7530) <= not(layer0_outputs(7215)) or (layer0_outputs(386));
    layer1_outputs(7531) <= not((layer0_outputs(570)) and (layer0_outputs(6897)));
    layer1_outputs(7532) <= not(layer0_outputs(6857));
    layer1_outputs(7533) <= (layer0_outputs(3161)) or (layer0_outputs(7670));
    layer1_outputs(7534) <= '0';
    layer1_outputs(7535) <= '1';
    layer1_outputs(7536) <= not((layer0_outputs(3193)) and (layer0_outputs(1907)));
    layer1_outputs(7537) <= (layer0_outputs(6128)) and (layer0_outputs(6179));
    layer1_outputs(7538) <= '0';
    layer1_outputs(7539) <= not((layer0_outputs(5186)) xor (layer0_outputs(4194)));
    layer1_outputs(7540) <= layer0_outputs(830);
    layer1_outputs(7541) <= (layer0_outputs(6875)) and not (layer0_outputs(2998));
    layer1_outputs(7542) <= layer0_outputs(921);
    layer1_outputs(7543) <= not((layer0_outputs(2466)) and (layer0_outputs(6416)));
    layer1_outputs(7544) <= (layer0_outputs(1953)) and not (layer0_outputs(1804));
    layer1_outputs(7545) <= (layer0_outputs(5606)) or (layer0_outputs(3436));
    layer1_outputs(7546) <= not(layer0_outputs(3933));
    layer1_outputs(7547) <= layer0_outputs(48);
    layer1_outputs(7548) <= (layer0_outputs(6300)) and not (layer0_outputs(1812));
    layer1_outputs(7549) <= not(layer0_outputs(5231));
    layer1_outputs(7550) <= not((layer0_outputs(5025)) or (layer0_outputs(2467)));
    layer1_outputs(7551) <= (layer0_outputs(5011)) or (layer0_outputs(5613));
    layer1_outputs(7552) <= layer0_outputs(3233);
    layer1_outputs(7553) <= (layer0_outputs(2726)) and (layer0_outputs(1612));
    layer1_outputs(7554) <= not(layer0_outputs(7103)) or (layer0_outputs(4295));
    layer1_outputs(7555) <= not((layer0_outputs(5864)) xor (layer0_outputs(6716)));
    layer1_outputs(7556) <= not(layer0_outputs(5386));
    layer1_outputs(7557) <= (layer0_outputs(4666)) and (layer0_outputs(1842));
    layer1_outputs(7558) <= (layer0_outputs(2517)) or (layer0_outputs(6927));
    layer1_outputs(7559) <= (layer0_outputs(1039)) and not (layer0_outputs(2018));
    layer1_outputs(7560) <= not((layer0_outputs(1832)) or (layer0_outputs(5151)));
    layer1_outputs(7561) <= layer0_outputs(1891);
    layer1_outputs(7562) <= not(layer0_outputs(3307));
    layer1_outputs(7563) <= not(layer0_outputs(1011)) or (layer0_outputs(2276));
    layer1_outputs(7564) <= (layer0_outputs(847)) and not (layer0_outputs(45));
    layer1_outputs(7565) <= not(layer0_outputs(4254));
    layer1_outputs(7566) <= '0';
    layer1_outputs(7567) <= not(layer0_outputs(5183));
    layer1_outputs(7568) <= (layer0_outputs(3399)) and (layer0_outputs(6786));
    layer1_outputs(7569) <= not(layer0_outputs(332)) or (layer0_outputs(4512));
    layer1_outputs(7570) <= not(layer0_outputs(6513));
    layer1_outputs(7571) <= layer0_outputs(2193);
    layer1_outputs(7572) <= (layer0_outputs(844)) and not (layer0_outputs(7469));
    layer1_outputs(7573) <= not((layer0_outputs(7516)) xor (layer0_outputs(7312)));
    layer1_outputs(7574) <= (layer0_outputs(4487)) and not (layer0_outputs(2423));
    layer1_outputs(7575) <= not(layer0_outputs(4578));
    layer1_outputs(7576) <= (layer0_outputs(5062)) and not (layer0_outputs(2244));
    layer1_outputs(7577) <= not(layer0_outputs(1301)) or (layer0_outputs(4591));
    layer1_outputs(7578) <= layer0_outputs(5459);
    layer1_outputs(7579) <= not(layer0_outputs(4078));
    layer1_outputs(7580) <= not(layer0_outputs(837)) or (layer0_outputs(5655));
    layer1_outputs(7581) <= (layer0_outputs(2911)) and not (layer0_outputs(2146));
    layer1_outputs(7582) <= (layer0_outputs(4801)) and (layer0_outputs(7039));
    layer1_outputs(7583) <= (layer0_outputs(5223)) and (layer0_outputs(6877));
    layer1_outputs(7584) <= not(layer0_outputs(1485));
    layer1_outputs(7585) <= (layer0_outputs(6480)) and (layer0_outputs(5630));
    layer1_outputs(7586) <= layer0_outputs(5508);
    layer1_outputs(7587) <= not(layer0_outputs(5485));
    layer1_outputs(7588) <= not(layer0_outputs(4888)) or (layer0_outputs(1825));
    layer1_outputs(7589) <= (layer0_outputs(7339)) and not (layer0_outputs(5359));
    layer1_outputs(7590) <= '0';
    layer1_outputs(7591) <= layer0_outputs(2831);
    layer1_outputs(7592) <= not((layer0_outputs(5288)) xor (layer0_outputs(217)));
    layer1_outputs(7593) <= not(layer0_outputs(5268));
    layer1_outputs(7594) <= '0';
    layer1_outputs(7595) <= (layer0_outputs(5233)) or (layer0_outputs(7408));
    layer1_outputs(7596) <= (layer0_outputs(7110)) and not (layer0_outputs(5914));
    layer1_outputs(7597) <= not((layer0_outputs(2663)) and (layer0_outputs(2599)));
    layer1_outputs(7598) <= not((layer0_outputs(4006)) and (layer0_outputs(3372)));
    layer1_outputs(7599) <= (layer0_outputs(2447)) and not (layer0_outputs(3545));
    layer1_outputs(7600) <= layer0_outputs(4649);
    layer1_outputs(7601) <= layer0_outputs(974);
    layer1_outputs(7602) <= not(layer0_outputs(5468)) or (layer0_outputs(117));
    layer1_outputs(7603) <= layer0_outputs(2850);
    layer1_outputs(7604) <= layer0_outputs(88);
    layer1_outputs(7605) <= not((layer0_outputs(6982)) or (layer0_outputs(7038)));
    layer1_outputs(7606) <= not(layer0_outputs(6235));
    layer1_outputs(7607) <= (layer0_outputs(4374)) or (layer0_outputs(2798));
    layer1_outputs(7608) <= layer0_outputs(4718);
    layer1_outputs(7609) <= layer0_outputs(6024);
    layer1_outputs(7610) <= not((layer0_outputs(3457)) or (layer0_outputs(4283)));
    layer1_outputs(7611) <= not(layer0_outputs(6666));
    layer1_outputs(7612) <= not(layer0_outputs(1235));
    layer1_outputs(7613) <= not(layer0_outputs(3513)) or (layer0_outputs(6985));
    layer1_outputs(7614) <= (layer0_outputs(6945)) and not (layer0_outputs(7501));
    layer1_outputs(7615) <= (layer0_outputs(3657)) and (layer0_outputs(5896));
    layer1_outputs(7616) <= layer0_outputs(492);
    layer1_outputs(7617) <= not((layer0_outputs(6634)) and (layer0_outputs(4259)));
    layer1_outputs(7618) <= not((layer0_outputs(6937)) or (layer0_outputs(5978)));
    layer1_outputs(7619) <= layer0_outputs(6898);
    layer1_outputs(7620) <= not(layer0_outputs(5984));
    layer1_outputs(7621) <= layer0_outputs(6824);
    layer1_outputs(7622) <= (layer0_outputs(4467)) xor (layer0_outputs(7262));
    layer1_outputs(7623) <= layer0_outputs(1956);
    layer1_outputs(7624) <= '0';
    layer1_outputs(7625) <= '0';
    layer1_outputs(7626) <= not(layer0_outputs(1188));
    layer1_outputs(7627) <= layer0_outputs(4124);
    layer1_outputs(7628) <= not(layer0_outputs(3735));
    layer1_outputs(7629) <= (layer0_outputs(6357)) xor (layer0_outputs(5924));
    layer1_outputs(7630) <= (layer0_outputs(3263)) and not (layer0_outputs(4869));
    layer1_outputs(7631) <= not(layer0_outputs(1717)) or (layer0_outputs(2631));
    layer1_outputs(7632) <= not((layer0_outputs(720)) xor (layer0_outputs(5320)));
    layer1_outputs(7633) <= (layer0_outputs(4304)) or (layer0_outputs(3721));
    layer1_outputs(7634) <= not((layer0_outputs(3378)) and (layer0_outputs(6921)));
    layer1_outputs(7635) <= (layer0_outputs(628)) and (layer0_outputs(4497));
    layer1_outputs(7636) <= not((layer0_outputs(1664)) and (layer0_outputs(975)));
    layer1_outputs(7637) <= not(layer0_outputs(4832));
    layer1_outputs(7638) <= not((layer0_outputs(3019)) or (layer0_outputs(6405)));
    layer1_outputs(7639) <= not(layer0_outputs(6816)) or (layer0_outputs(758));
    layer1_outputs(7640) <= not(layer0_outputs(2928)) or (layer0_outputs(3651));
    layer1_outputs(7641) <= layer0_outputs(865);
    layer1_outputs(7642) <= not((layer0_outputs(3698)) xor (layer0_outputs(3034)));
    layer1_outputs(7643) <= not(layer0_outputs(4142));
    layer1_outputs(7644) <= layer0_outputs(5274);
    layer1_outputs(7645) <= (layer0_outputs(2252)) and not (layer0_outputs(239));
    layer1_outputs(7646) <= layer0_outputs(1562);
    layer1_outputs(7647) <= layer0_outputs(4203);
    layer1_outputs(7648) <= '1';
    layer1_outputs(7649) <= not(layer0_outputs(4839)) or (layer0_outputs(454));
    layer1_outputs(7650) <= not(layer0_outputs(1667));
    layer1_outputs(7651) <= not(layer0_outputs(5222)) or (layer0_outputs(3770));
    layer1_outputs(7652) <= '0';
    layer1_outputs(7653) <= (layer0_outputs(5231)) or (layer0_outputs(7256));
    layer1_outputs(7654) <= (layer0_outputs(6659)) and not (layer0_outputs(4071));
    layer1_outputs(7655) <= layer0_outputs(7356);
    layer1_outputs(7656) <= not((layer0_outputs(5962)) and (layer0_outputs(4600)));
    layer1_outputs(7657) <= not(layer0_outputs(1204)) or (layer0_outputs(6325));
    layer1_outputs(7658) <= not((layer0_outputs(27)) and (layer0_outputs(6140)));
    layer1_outputs(7659) <= not(layer0_outputs(5452));
    layer1_outputs(7660) <= layer0_outputs(6246);
    layer1_outputs(7661) <= not((layer0_outputs(3101)) or (layer0_outputs(4665)));
    layer1_outputs(7662) <= not((layer0_outputs(4555)) and (layer0_outputs(1843)));
    layer1_outputs(7663) <= not(layer0_outputs(5531));
    layer1_outputs(7664) <= not(layer0_outputs(6292)) or (layer0_outputs(6139));
    layer1_outputs(7665) <= not(layer0_outputs(3963));
    layer1_outputs(7666) <= not(layer0_outputs(231)) or (layer0_outputs(4952));
    layer1_outputs(7667) <= (layer0_outputs(4601)) or (layer0_outputs(6034));
    layer1_outputs(7668) <= not((layer0_outputs(5398)) xor (layer0_outputs(3038)));
    layer1_outputs(7669) <= not(layer0_outputs(7004)) or (layer0_outputs(6521));
    layer1_outputs(7670) <= not(layer0_outputs(6676));
    layer1_outputs(7671) <= (layer0_outputs(3358)) or (layer0_outputs(379));
    layer1_outputs(7672) <= '0';
    layer1_outputs(7673) <= not((layer0_outputs(1718)) xor (layer0_outputs(2752)));
    layer1_outputs(7674) <= not((layer0_outputs(4307)) and (layer0_outputs(3131)));
    layer1_outputs(7675) <= not(layer0_outputs(3477));
    layer1_outputs(7676) <= layer0_outputs(2110);
    layer1_outputs(7677) <= layer0_outputs(1998);
    layer1_outputs(7678) <= '1';
    layer1_outputs(7679) <= not(layer0_outputs(2601)) or (layer0_outputs(1945));
    layer2_outputs(0) <= not(layer1_outputs(7516));
    layer2_outputs(1) <= not(layer1_outputs(5646)) or (layer1_outputs(418));
    layer2_outputs(2) <= not(layer1_outputs(3819));
    layer2_outputs(3) <= not(layer1_outputs(2882));
    layer2_outputs(4) <= '0';
    layer2_outputs(5) <= not(layer1_outputs(2800));
    layer2_outputs(6) <= (layer1_outputs(2772)) or (layer1_outputs(197));
    layer2_outputs(7) <= not(layer1_outputs(4676));
    layer2_outputs(8) <= not(layer1_outputs(7324));
    layer2_outputs(9) <= layer1_outputs(547);
    layer2_outputs(10) <= (layer1_outputs(1407)) xor (layer1_outputs(7616));
    layer2_outputs(11) <= (layer1_outputs(3619)) and not (layer1_outputs(7284));
    layer2_outputs(12) <= layer1_outputs(919);
    layer2_outputs(13) <= not(layer1_outputs(2585));
    layer2_outputs(14) <= (layer1_outputs(5889)) or (layer1_outputs(1617));
    layer2_outputs(15) <= (layer1_outputs(4313)) or (layer1_outputs(5066));
    layer2_outputs(16) <= not(layer1_outputs(5902)) or (layer1_outputs(2367));
    layer2_outputs(17) <= layer1_outputs(366);
    layer2_outputs(18) <= layer1_outputs(6038);
    layer2_outputs(19) <= layer1_outputs(5062);
    layer2_outputs(20) <= (layer1_outputs(3775)) or (layer1_outputs(1843));
    layer2_outputs(21) <= (layer1_outputs(6638)) or (layer1_outputs(5351));
    layer2_outputs(22) <= layer1_outputs(122);
    layer2_outputs(23) <= '0';
    layer2_outputs(24) <= layer1_outputs(5822);
    layer2_outputs(25) <= (layer1_outputs(4351)) and (layer1_outputs(6882));
    layer2_outputs(26) <= (layer1_outputs(3851)) and not (layer1_outputs(5305));
    layer2_outputs(27) <= (layer1_outputs(1584)) and not (layer1_outputs(4505));
    layer2_outputs(28) <= not(layer1_outputs(5277));
    layer2_outputs(29) <= (layer1_outputs(47)) and (layer1_outputs(1463));
    layer2_outputs(30) <= not(layer1_outputs(2035)) or (layer1_outputs(7436));
    layer2_outputs(31) <= layer1_outputs(5024);
    layer2_outputs(32) <= (layer1_outputs(1050)) and not (layer1_outputs(1786));
    layer2_outputs(33) <= (layer1_outputs(1341)) and (layer1_outputs(7165));
    layer2_outputs(34) <= not(layer1_outputs(2968));
    layer2_outputs(35) <= not(layer1_outputs(4127));
    layer2_outputs(36) <= not((layer1_outputs(6866)) or (layer1_outputs(2939)));
    layer2_outputs(37) <= layer1_outputs(4746);
    layer2_outputs(38) <= (layer1_outputs(1193)) and (layer1_outputs(739));
    layer2_outputs(39) <= (layer1_outputs(2190)) and (layer1_outputs(1679));
    layer2_outputs(40) <= layer1_outputs(4242);
    layer2_outputs(41) <= not(layer1_outputs(6386)) or (layer1_outputs(2847));
    layer2_outputs(42) <= not((layer1_outputs(4701)) or (layer1_outputs(1398)));
    layer2_outputs(43) <= '0';
    layer2_outputs(44) <= (layer1_outputs(4187)) and not (layer1_outputs(37));
    layer2_outputs(45) <= not((layer1_outputs(3824)) or (layer1_outputs(5123)));
    layer2_outputs(46) <= layer1_outputs(1673);
    layer2_outputs(47) <= layer1_outputs(5397);
    layer2_outputs(48) <= not(layer1_outputs(2710));
    layer2_outputs(49) <= layer1_outputs(30);
    layer2_outputs(50) <= (layer1_outputs(4999)) and (layer1_outputs(5722));
    layer2_outputs(51) <= (layer1_outputs(3353)) and not (layer1_outputs(2669));
    layer2_outputs(52) <= (layer1_outputs(2395)) and (layer1_outputs(2956));
    layer2_outputs(53) <= not(layer1_outputs(5758));
    layer2_outputs(54) <= not(layer1_outputs(7437));
    layer2_outputs(55) <= layer1_outputs(1892);
    layer2_outputs(56) <= not(layer1_outputs(129));
    layer2_outputs(57) <= not(layer1_outputs(1761));
    layer2_outputs(58) <= (layer1_outputs(2427)) and not (layer1_outputs(1125));
    layer2_outputs(59) <= not(layer1_outputs(556)) or (layer1_outputs(2420));
    layer2_outputs(60) <= not(layer1_outputs(3479));
    layer2_outputs(61) <= not(layer1_outputs(3079));
    layer2_outputs(62) <= not((layer1_outputs(5899)) and (layer1_outputs(2906)));
    layer2_outputs(63) <= not(layer1_outputs(2767)) or (layer1_outputs(7644));
    layer2_outputs(64) <= not(layer1_outputs(6234));
    layer2_outputs(65) <= (layer1_outputs(558)) and not (layer1_outputs(3065));
    layer2_outputs(66) <= layer1_outputs(4261);
    layer2_outputs(67) <= (layer1_outputs(4750)) xor (layer1_outputs(2364));
    layer2_outputs(68) <= not((layer1_outputs(5964)) and (layer1_outputs(5232)));
    layer2_outputs(69) <= not(layer1_outputs(689));
    layer2_outputs(70) <= '1';
    layer2_outputs(71) <= layer1_outputs(7521);
    layer2_outputs(72) <= not(layer1_outputs(6645)) or (layer1_outputs(1870));
    layer2_outputs(73) <= (layer1_outputs(5511)) and not (layer1_outputs(393));
    layer2_outputs(74) <= not(layer1_outputs(5827));
    layer2_outputs(75) <= not(layer1_outputs(3894));
    layer2_outputs(76) <= not(layer1_outputs(7390)) or (layer1_outputs(2955));
    layer2_outputs(77) <= not((layer1_outputs(4331)) and (layer1_outputs(1722)));
    layer2_outputs(78) <= layer1_outputs(5475);
    layer2_outputs(79) <= layer1_outputs(321);
    layer2_outputs(80) <= (layer1_outputs(2309)) and not (layer1_outputs(3153));
    layer2_outputs(81) <= not((layer1_outputs(5290)) xor (layer1_outputs(1845)));
    layer2_outputs(82) <= not((layer1_outputs(2767)) and (layer1_outputs(717)));
    layer2_outputs(83) <= '1';
    layer2_outputs(84) <= not(layer1_outputs(4109));
    layer2_outputs(85) <= (layer1_outputs(5464)) and not (layer1_outputs(3627));
    layer2_outputs(86) <= not(layer1_outputs(2999)) or (layer1_outputs(6540));
    layer2_outputs(87) <= (layer1_outputs(5622)) and not (layer1_outputs(364));
    layer2_outputs(88) <= (layer1_outputs(2150)) and (layer1_outputs(7581));
    layer2_outputs(89) <= layer1_outputs(4484);
    layer2_outputs(90) <= '1';
    layer2_outputs(91) <= not(layer1_outputs(174));
    layer2_outputs(92) <= not((layer1_outputs(7385)) and (layer1_outputs(3487)));
    layer2_outputs(93) <= not((layer1_outputs(4982)) and (layer1_outputs(1030)));
    layer2_outputs(94) <= not(layer1_outputs(5227));
    layer2_outputs(95) <= not(layer1_outputs(3641)) or (layer1_outputs(3256));
    layer2_outputs(96) <= layer1_outputs(1540);
    layer2_outputs(97) <= (layer1_outputs(4579)) and not (layer1_outputs(3840));
    layer2_outputs(98) <= (layer1_outputs(242)) and not (layer1_outputs(4597));
    layer2_outputs(99) <= not((layer1_outputs(3283)) or (layer1_outputs(7499)));
    layer2_outputs(100) <= (layer1_outputs(661)) and (layer1_outputs(5054));
    layer2_outputs(101) <= layer1_outputs(6513);
    layer2_outputs(102) <= layer1_outputs(6877);
    layer2_outputs(103) <= layer1_outputs(7364);
    layer2_outputs(104) <= not(layer1_outputs(3141)) or (layer1_outputs(3615));
    layer2_outputs(105) <= not(layer1_outputs(6564)) or (layer1_outputs(7053));
    layer2_outputs(106) <= not(layer1_outputs(2449));
    layer2_outputs(107) <= (layer1_outputs(7249)) and (layer1_outputs(6117));
    layer2_outputs(108) <= not((layer1_outputs(6044)) and (layer1_outputs(3455)));
    layer2_outputs(109) <= (layer1_outputs(947)) and not (layer1_outputs(6086));
    layer2_outputs(110) <= layer1_outputs(3623);
    layer2_outputs(111) <= (layer1_outputs(5457)) and not (layer1_outputs(1891));
    layer2_outputs(112) <= layer1_outputs(7585);
    layer2_outputs(113) <= (layer1_outputs(5478)) or (layer1_outputs(666));
    layer2_outputs(114) <= not(layer1_outputs(3684));
    layer2_outputs(115) <= not(layer1_outputs(5285));
    layer2_outputs(116) <= (layer1_outputs(7470)) or (layer1_outputs(950));
    layer2_outputs(117) <= layer1_outputs(1982);
    layer2_outputs(118) <= not(layer1_outputs(5635)) or (layer1_outputs(681));
    layer2_outputs(119) <= not(layer1_outputs(6703)) or (layer1_outputs(2250));
    layer2_outputs(120) <= '0';
    layer2_outputs(121) <= not(layer1_outputs(5695));
    layer2_outputs(122) <= (layer1_outputs(2306)) xor (layer1_outputs(3254));
    layer2_outputs(123) <= layer1_outputs(6320);
    layer2_outputs(124) <= not((layer1_outputs(5614)) and (layer1_outputs(7004)));
    layer2_outputs(125) <= layer1_outputs(5460);
    layer2_outputs(126) <= (layer1_outputs(5345)) and not (layer1_outputs(6598));
    layer2_outputs(127) <= layer1_outputs(6646);
    layer2_outputs(128) <= not((layer1_outputs(4797)) and (layer1_outputs(5784)));
    layer2_outputs(129) <= (layer1_outputs(7241)) or (layer1_outputs(1415));
    layer2_outputs(130) <= not(layer1_outputs(2135));
    layer2_outputs(131) <= layer1_outputs(6932);
    layer2_outputs(132) <= layer1_outputs(4986);
    layer2_outputs(133) <= (layer1_outputs(6475)) and not (layer1_outputs(3509));
    layer2_outputs(134) <= not(layer1_outputs(3135)) or (layer1_outputs(1690));
    layer2_outputs(135) <= not(layer1_outputs(2126));
    layer2_outputs(136) <= (layer1_outputs(5018)) and not (layer1_outputs(5770));
    layer2_outputs(137) <= layer1_outputs(6853);
    layer2_outputs(138) <= layer1_outputs(6863);
    layer2_outputs(139) <= (layer1_outputs(2201)) or (layer1_outputs(3158));
    layer2_outputs(140) <= not(layer1_outputs(6900));
    layer2_outputs(141) <= (layer1_outputs(852)) or (layer1_outputs(6412));
    layer2_outputs(142) <= '0';
    layer2_outputs(143) <= layer1_outputs(1157);
    layer2_outputs(144) <= (layer1_outputs(480)) and not (layer1_outputs(7026));
    layer2_outputs(145) <= layer1_outputs(764);
    layer2_outputs(146) <= not(layer1_outputs(4571));
    layer2_outputs(147) <= not(layer1_outputs(6772));
    layer2_outputs(148) <= not((layer1_outputs(1196)) and (layer1_outputs(1912)));
    layer2_outputs(149) <= not((layer1_outputs(2779)) and (layer1_outputs(7011)));
    layer2_outputs(150) <= layer1_outputs(5939);
    layer2_outputs(151) <= (layer1_outputs(574)) and (layer1_outputs(1417));
    layer2_outputs(152) <= (layer1_outputs(306)) and (layer1_outputs(661));
    layer2_outputs(153) <= not((layer1_outputs(3581)) and (layer1_outputs(3751)));
    layer2_outputs(154) <= layer1_outputs(288);
    layer2_outputs(155) <= not((layer1_outputs(3121)) or (layer1_outputs(6988)));
    layer2_outputs(156) <= layer1_outputs(2804);
    layer2_outputs(157) <= (layer1_outputs(993)) and (layer1_outputs(4805));
    layer2_outputs(158) <= not((layer1_outputs(960)) or (layer1_outputs(3339)));
    layer2_outputs(159) <= (layer1_outputs(6178)) and not (layer1_outputs(3763));
    layer2_outputs(160) <= not((layer1_outputs(185)) or (layer1_outputs(3795)));
    layer2_outputs(161) <= layer1_outputs(4803);
    layer2_outputs(162) <= (layer1_outputs(2457)) and not (layer1_outputs(4876));
    layer2_outputs(163) <= not(layer1_outputs(4019));
    layer2_outputs(164) <= layer1_outputs(7442);
    layer2_outputs(165) <= layer1_outputs(1664);
    layer2_outputs(166) <= (layer1_outputs(6970)) and not (layer1_outputs(130));
    layer2_outputs(167) <= not(layer1_outputs(381));
    layer2_outputs(168) <= (layer1_outputs(5670)) and (layer1_outputs(3640));
    layer2_outputs(169) <= not(layer1_outputs(1334)) or (layer1_outputs(3943));
    layer2_outputs(170) <= layer1_outputs(7009);
    layer2_outputs(171) <= not((layer1_outputs(4646)) and (layer1_outputs(4379)));
    layer2_outputs(172) <= (layer1_outputs(207)) and not (layer1_outputs(3774));
    layer2_outputs(173) <= layer1_outputs(6248);
    layer2_outputs(174) <= not((layer1_outputs(6162)) or (layer1_outputs(1507)));
    layer2_outputs(175) <= not(layer1_outputs(5289)) or (layer1_outputs(6963));
    layer2_outputs(176) <= '1';
    layer2_outputs(177) <= (layer1_outputs(3971)) xor (layer1_outputs(1082));
    layer2_outputs(178) <= '0';
    layer2_outputs(179) <= (layer1_outputs(1733)) and not (layer1_outputs(6658));
    layer2_outputs(180) <= not(layer1_outputs(7593));
    layer2_outputs(181) <= '1';
    layer2_outputs(182) <= (layer1_outputs(4298)) xor (layer1_outputs(7608));
    layer2_outputs(183) <= layer1_outputs(4441);
    layer2_outputs(184) <= layer1_outputs(2505);
    layer2_outputs(185) <= not(layer1_outputs(6686)) or (layer1_outputs(3123));
    layer2_outputs(186) <= not(layer1_outputs(2088)) or (layer1_outputs(2194));
    layer2_outputs(187) <= layer1_outputs(5706);
    layer2_outputs(188) <= not(layer1_outputs(7019));
    layer2_outputs(189) <= layer1_outputs(1758);
    layer2_outputs(190) <= (layer1_outputs(3808)) and not (layer1_outputs(1827));
    layer2_outputs(191) <= not(layer1_outputs(6864)) or (layer1_outputs(7343));
    layer2_outputs(192) <= '0';
    layer2_outputs(193) <= layer1_outputs(7440);
    layer2_outputs(194) <= not(layer1_outputs(5227));
    layer2_outputs(195) <= (layer1_outputs(305)) or (layer1_outputs(7079));
    layer2_outputs(196) <= not(layer1_outputs(2510));
    layer2_outputs(197) <= (layer1_outputs(7671)) or (layer1_outputs(3334));
    layer2_outputs(198) <= (layer1_outputs(2361)) and not (layer1_outputs(5181));
    layer2_outputs(199) <= layer1_outputs(5140);
    layer2_outputs(200) <= not(layer1_outputs(475));
    layer2_outputs(201) <= not(layer1_outputs(7236));
    layer2_outputs(202) <= layer1_outputs(7661);
    layer2_outputs(203) <= (layer1_outputs(7193)) and not (layer1_outputs(1472));
    layer2_outputs(204) <= not(layer1_outputs(3747)) or (layer1_outputs(1369));
    layer2_outputs(205) <= (layer1_outputs(5136)) and (layer1_outputs(7237));
    layer2_outputs(206) <= not(layer1_outputs(3895));
    layer2_outputs(207) <= (layer1_outputs(1031)) and not (layer1_outputs(5057));
    layer2_outputs(208) <= layer1_outputs(5048);
    layer2_outputs(209) <= (layer1_outputs(6529)) and not (layer1_outputs(7439));
    layer2_outputs(210) <= layer1_outputs(6587);
    layer2_outputs(211) <= not(layer1_outputs(210)) or (layer1_outputs(4303));
    layer2_outputs(212) <= not(layer1_outputs(5495)) or (layer1_outputs(834));
    layer2_outputs(213) <= not(layer1_outputs(6499));
    layer2_outputs(214) <= not((layer1_outputs(1342)) or (layer1_outputs(4113)));
    layer2_outputs(215) <= (layer1_outputs(4847)) and not (layer1_outputs(192));
    layer2_outputs(216) <= not(layer1_outputs(2740));
    layer2_outputs(217) <= (layer1_outputs(6949)) or (layer1_outputs(4384));
    layer2_outputs(218) <= '0';
    layer2_outputs(219) <= '0';
    layer2_outputs(220) <= (layer1_outputs(6594)) and not (layer1_outputs(4095));
    layer2_outputs(221) <= layer1_outputs(5153);
    layer2_outputs(222) <= not(layer1_outputs(3997));
    layer2_outputs(223) <= (layer1_outputs(1360)) or (layer1_outputs(5838));
    layer2_outputs(224) <= not(layer1_outputs(2188));
    layer2_outputs(225) <= not(layer1_outputs(3838)) or (layer1_outputs(7032));
    layer2_outputs(226) <= layer1_outputs(4231);
    layer2_outputs(227) <= not((layer1_outputs(3572)) or (layer1_outputs(2406)));
    layer2_outputs(228) <= not((layer1_outputs(6188)) or (layer1_outputs(420)));
    layer2_outputs(229) <= (layer1_outputs(1402)) or (layer1_outputs(7248));
    layer2_outputs(230) <= not(layer1_outputs(1895));
    layer2_outputs(231) <= (layer1_outputs(3810)) xor (layer1_outputs(754));
    layer2_outputs(232) <= (layer1_outputs(6261)) and not (layer1_outputs(3608));
    layer2_outputs(233) <= not(layer1_outputs(7180)) or (layer1_outputs(4263));
    layer2_outputs(234) <= '1';
    layer2_outputs(235) <= (layer1_outputs(1623)) and (layer1_outputs(5593));
    layer2_outputs(236) <= not(layer1_outputs(4575));
    layer2_outputs(237) <= layer1_outputs(1050);
    layer2_outputs(238) <= (layer1_outputs(2418)) or (layer1_outputs(5362));
    layer2_outputs(239) <= '0';
    layer2_outputs(240) <= layer1_outputs(7640);
    layer2_outputs(241) <= not(layer1_outputs(4840));
    layer2_outputs(242) <= not(layer1_outputs(527));
    layer2_outputs(243) <= layer1_outputs(2441);
    layer2_outputs(244) <= (layer1_outputs(7607)) and (layer1_outputs(3154));
    layer2_outputs(245) <= not(layer1_outputs(7675));
    layer2_outputs(246) <= (layer1_outputs(4867)) xor (layer1_outputs(4950));
    layer2_outputs(247) <= not(layer1_outputs(5344)) or (layer1_outputs(5542));
    layer2_outputs(248) <= '0';
    layer2_outputs(249) <= layer1_outputs(7597);
    layer2_outputs(250) <= not(layer1_outputs(6430)) or (layer1_outputs(2291));
    layer2_outputs(251) <= (layer1_outputs(2982)) and not (layer1_outputs(2258));
    layer2_outputs(252) <= not(layer1_outputs(5260)) or (layer1_outputs(4774));
    layer2_outputs(253) <= (layer1_outputs(1754)) and (layer1_outputs(6455));
    layer2_outputs(254) <= (layer1_outputs(4340)) or (layer1_outputs(4123));
    layer2_outputs(255) <= not(layer1_outputs(3747));
    layer2_outputs(256) <= '0';
    layer2_outputs(257) <= layer1_outputs(5059);
    layer2_outputs(258) <= layer1_outputs(6650);
    layer2_outputs(259) <= (layer1_outputs(5756)) and not (layer1_outputs(5028));
    layer2_outputs(260) <= not(layer1_outputs(3199)) or (layer1_outputs(2007));
    layer2_outputs(261) <= (layer1_outputs(3945)) and not (layer1_outputs(6539));
    layer2_outputs(262) <= not(layer1_outputs(1630));
    layer2_outputs(263) <= layer1_outputs(4839);
    layer2_outputs(264) <= not((layer1_outputs(2589)) and (layer1_outputs(2658)));
    layer2_outputs(265) <= not(layer1_outputs(2784)) or (layer1_outputs(2452));
    layer2_outputs(266) <= layer1_outputs(3057);
    layer2_outputs(267) <= not((layer1_outputs(6304)) and (layer1_outputs(658)));
    layer2_outputs(268) <= not(layer1_outputs(3913)) or (layer1_outputs(6152));
    layer2_outputs(269) <= layer1_outputs(5832);
    layer2_outputs(270) <= not((layer1_outputs(118)) or (layer1_outputs(5269)));
    layer2_outputs(271) <= not((layer1_outputs(6060)) or (layer1_outputs(6781)));
    layer2_outputs(272) <= layer1_outputs(5210);
    layer2_outputs(273) <= not(layer1_outputs(3430));
    layer2_outputs(274) <= not(layer1_outputs(3984)) or (layer1_outputs(6084));
    layer2_outputs(275) <= layer1_outputs(2543);
    layer2_outputs(276) <= not((layer1_outputs(589)) and (layer1_outputs(4247)));
    layer2_outputs(277) <= not(layer1_outputs(560)) or (layer1_outputs(216));
    layer2_outputs(278) <= not((layer1_outputs(1523)) and (layer1_outputs(2821)));
    layer2_outputs(279) <= not(layer1_outputs(4102)) or (layer1_outputs(811));
    layer2_outputs(280) <= (layer1_outputs(3125)) and not (layer1_outputs(3445));
    layer2_outputs(281) <= not(layer1_outputs(1370)) or (layer1_outputs(7509));
    layer2_outputs(282) <= not(layer1_outputs(3364));
    layer2_outputs(283) <= (layer1_outputs(1286)) and (layer1_outputs(272));
    layer2_outputs(284) <= layer1_outputs(1116);
    layer2_outputs(285) <= (layer1_outputs(5557)) and (layer1_outputs(3212));
    layer2_outputs(286) <= not(layer1_outputs(449)) or (layer1_outputs(2493));
    layer2_outputs(287) <= (layer1_outputs(3827)) or (layer1_outputs(574));
    layer2_outputs(288) <= not((layer1_outputs(3922)) and (layer1_outputs(6499)));
    layer2_outputs(289) <= layer1_outputs(1596);
    layer2_outputs(290) <= not(layer1_outputs(6456));
    layer2_outputs(291) <= not((layer1_outputs(1598)) and (layer1_outputs(5683)));
    layer2_outputs(292) <= not(layer1_outputs(5927));
    layer2_outputs(293) <= '1';
    layer2_outputs(294) <= not((layer1_outputs(3580)) or (layer1_outputs(3635)));
    layer2_outputs(295) <= not(layer1_outputs(5264));
    layer2_outputs(296) <= (layer1_outputs(6352)) and not (layer1_outputs(5523));
    layer2_outputs(297) <= not((layer1_outputs(4669)) xor (layer1_outputs(3759)));
    layer2_outputs(298) <= not(layer1_outputs(320));
    layer2_outputs(299) <= (layer1_outputs(1515)) xor (layer1_outputs(6151));
    layer2_outputs(300) <= not(layer1_outputs(7676));
    layer2_outputs(301) <= layer1_outputs(5995);
    layer2_outputs(302) <= layer1_outputs(5714);
    layer2_outputs(303) <= layer1_outputs(4097);
    layer2_outputs(304) <= not((layer1_outputs(2052)) and (layer1_outputs(867)));
    layer2_outputs(305) <= (layer1_outputs(3010)) and not (layer1_outputs(1559));
    layer2_outputs(306) <= (layer1_outputs(5457)) and not (layer1_outputs(962));
    layer2_outputs(307) <= (layer1_outputs(7071)) and (layer1_outputs(5737));
    layer2_outputs(308) <= not(layer1_outputs(4310));
    layer2_outputs(309) <= not((layer1_outputs(2829)) and (layer1_outputs(6465)));
    layer2_outputs(310) <= not(layer1_outputs(4311));
    layer2_outputs(311) <= not(layer1_outputs(1795)) or (layer1_outputs(6722));
    layer2_outputs(312) <= (layer1_outputs(3076)) or (layer1_outputs(7068));
    layer2_outputs(313) <= layer1_outputs(4837);
    layer2_outputs(314) <= not(layer1_outputs(2616));
    layer2_outputs(315) <= not(layer1_outputs(4688));
    layer2_outputs(316) <= (layer1_outputs(7369)) and not (layer1_outputs(3124));
    layer2_outputs(317) <= (layer1_outputs(1501)) and not (layer1_outputs(3341));
    layer2_outputs(318) <= '1';
    layer2_outputs(319) <= (layer1_outputs(1636)) or (layer1_outputs(5553));
    layer2_outputs(320) <= layer1_outputs(6621);
    layer2_outputs(321) <= layer1_outputs(4544);
    layer2_outputs(322) <= not(layer1_outputs(2155));
    layer2_outputs(323) <= not((layer1_outputs(2846)) and (layer1_outputs(7621)));
    layer2_outputs(324) <= (layer1_outputs(2733)) and (layer1_outputs(740));
    layer2_outputs(325) <= (layer1_outputs(2018)) and not (layer1_outputs(7016));
    layer2_outputs(326) <= layer1_outputs(6763);
    layer2_outputs(327) <= layer1_outputs(2388);
    layer2_outputs(328) <= (layer1_outputs(423)) and not (layer1_outputs(2835));
    layer2_outputs(329) <= layer1_outputs(428);
    layer2_outputs(330) <= not(layer1_outputs(6512));
    layer2_outputs(331) <= not(layer1_outputs(5906));
    layer2_outputs(332) <= layer1_outputs(684);
    layer2_outputs(333) <= '1';
    layer2_outputs(334) <= not(layer1_outputs(7460));
    layer2_outputs(335) <= not(layer1_outputs(4625));
    layer2_outputs(336) <= not(layer1_outputs(5813));
    layer2_outputs(337) <= (layer1_outputs(4944)) and not (layer1_outputs(1205));
    layer2_outputs(338) <= layer1_outputs(5360);
    layer2_outputs(339) <= not(layer1_outputs(3649)) or (layer1_outputs(559));
    layer2_outputs(340) <= (layer1_outputs(5966)) or (layer1_outputs(5388));
    layer2_outputs(341) <= '0';
    layer2_outputs(342) <= not(layer1_outputs(845)) or (layer1_outputs(524));
    layer2_outputs(343) <= layer1_outputs(1014);
    layer2_outputs(344) <= layer1_outputs(3530);
    layer2_outputs(345) <= layer1_outputs(7201);
    layer2_outputs(346) <= layer1_outputs(4991);
    layer2_outputs(347) <= not(layer1_outputs(1322)) or (layer1_outputs(1565));
    layer2_outputs(348) <= not((layer1_outputs(6526)) or (layer1_outputs(2329)));
    layer2_outputs(349) <= layer1_outputs(4201);
    layer2_outputs(350) <= not((layer1_outputs(5786)) or (layer1_outputs(1946)));
    layer2_outputs(351) <= (layer1_outputs(6623)) and not (layer1_outputs(7024));
    layer2_outputs(352) <= (layer1_outputs(2371)) and (layer1_outputs(7325));
    layer2_outputs(353) <= (layer1_outputs(2939)) xor (layer1_outputs(1702));
    layer2_outputs(354) <= (layer1_outputs(793)) or (layer1_outputs(5231));
    layer2_outputs(355) <= not((layer1_outputs(7376)) and (layer1_outputs(2465)));
    layer2_outputs(356) <= (layer1_outputs(7152)) xor (layer1_outputs(7090));
    layer2_outputs(357) <= not(layer1_outputs(743));
    layer2_outputs(358) <= layer1_outputs(521);
    layer2_outputs(359) <= not((layer1_outputs(5145)) and (layer1_outputs(3090)));
    layer2_outputs(360) <= '1';
    layer2_outputs(361) <= (layer1_outputs(4180)) and not (layer1_outputs(7296));
    layer2_outputs(362) <= not((layer1_outputs(5787)) or (layer1_outputs(2551)));
    layer2_outputs(363) <= not(layer1_outputs(5812));
    layer2_outputs(364) <= not((layer1_outputs(92)) or (layer1_outputs(2789)));
    layer2_outputs(365) <= not(layer1_outputs(1587)) or (layer1_outputs(6055));
    layer2_outputs(366) <= not(layer1_outputs(4952));
    layer2_outputs(367) <= not(layer1_outputs(3389));
    layer2_outputs(368) <= (layer1_outputs(869)) and not (layer1_outputs(1918));
    layer2_outputs(369) <= (layer1_outputs(6055)) and not (layer1_outputs(4977));
    layer2_outputs(370) <= not(layer1_outputs(2610)) or (layer1_outputs(7076));
    layer2_outputs(371) <= layer1_outputs(6689);
    layer2_outputs(372) <= (layer1_outputs(745)) and not (layer1_outputs(4998));
    layer2_outputs(373) <= '1';
    layer2_outputs(374) <= layer1_outputs(6991);
    layer2_outputs(375) <= '1';
    layer2_outputs(376) <= layer1_outputs(4060);
    layer2_outputs(377) <= (layer1_outputs(716)) and (layer1_outputs(1537));
    layer2_outputs(378) <= not(layer1_outputs(3626)) or (layer1_outputs(6382));
    layer2_outputs(379) <= '0';
    layer2_outputs(380) <= (layer1_outputs(3541)) and not (layer1_outputs(4872));
    layer2_outputs(381) <= (layer1_outputs(6086)) and not (layer1_outputs(2224));
    layer2_outputs(382) <= layer1_outputs(4740);
    layer2_outputs(383) <= layer1_outputs(3477);
    layer2_outputs(384) <= layer1_outputs(6030);
    layer2_outputs(385) <= not(layer1_outputs(4739)) or (layer1_outputs(4569));
    layer2_outputs(386) <= not(layer1_outputs(6196)) or (layer1_outputs(7254));
    layer2_outputs(387) <= (layer1_outputs(2104)) and not (layer1_outputs(6750));
    layer2_outputs(388) <= layer1_outputs(7152);
    layer2_outputs(389) <= layer1_outputs(1888);
    layer2_outputs(390) <= layer1_outputs(4775);
    layer2_outputs(391) <= not(layer1_outputs(5315)) or (layer1_outputs(1696));
    layer2_outputs(392) <= not(layer1_outputs(236));
    layer2_outputs(393) <= layer1_outputs(5911);
    layer2_outputs(394) <= (layer1_outputs(2489)) or (layer1_outputs(1339));
    layer2_outputs(395) <= (layer1_outputs(5968)) and (layer1_outputs(1804));
    layer2_outputs(396) <= not((layer1_outputs(5981)) or (layer1_outputs(1364)));
    layer2_outputs(397) <= (layer1_outputs(6679)) or (layer1_outputs(4831));
    layer2_outputs(398) <= layer1_outputs(3990);
    layer2_outputs(399) <= not((layer1_outputs(3037)) and (layer1_outputs(366)));
    layer2_outputs(400) <= not((layer1_outputs(3327)) and (layer1_outputs(4304)));
    layer2_outputs(401) <= not(layer1_outputs(518));
    layer2_outputs(402) <= '0';
    layer2_outputs(403) <= layer1_outputs(2340);
    layer2_outputs(404) <= layer1_outputs(1638);
    layer2_outputs(405) <= layer1_outputs(7199);
    layer2_outputs(406) <= not(layer1_outputs(641));
    layer2_outputs(407) <= not(layer1_outputs(1231));
    layer2_outputs(408) <= not((layer1_outputs(4261)) or (layer1_outputs(6652)));
    layer2_outputs(409) <= not((layer1_outputs(7500)) or (layer1_outputs(1240)));
    layer2_outputs(410) <= (layer1_outputs(4893)) or (layer1_outputs(239));
    layer2_outputs(411) <= (layer1_outputs(4813)) or (layer1_outputs(4371));
    layer2_outputs(412) <= (layer1_outputs(789)) and not (layer1_outputs(6026));
    layer2_outputs(413) <= '1';
    layer2_outputs(414) <= layer1_outputs(5256);
    layer2_outputs(415) <= not(layer1_outputs(2305)) or (layer1_outputs(4211));
    layer2_outputs(416) <= (layer1_outputs(6228)) and not (layer1_outputs(3312));
    layer2_outputs(417) <= not(layer1_outputs(3740));
    layer2_outputs(418) <= not(layer1_outputs(5829)) or (layer1_outputs(2932));
    layer2_outputs(419) <= layer1_outputs(2822);
    layer2_outputs(420) <= (layer1_outputs(3145)) and (layer1_outputs(6171));
    layer2_outputs(421) <= not(layer1_outputs(1190));
    layer2_outputs(422) <= not((layer1_outputs(971)) or (layer1_outputs(5081)));
    layer2_outputs(423) <= not(layer1_outputs(3035)) or (layer1_outputs(2441));
    layer2_outputs(424) <= not(layer1_outputs(3402));
    layer2_outputs(425) <= layer1_outputs(154);
    layer2_outputs(426) <= (layer1_outputs(6522)) and (layer1_outputs(3558));
    layer2_outputs(427) <= (layer1_outputs(2137)) and (layer1_outputs(2374));
    layer2_outputs(428) <= (layer1_outputs(6483)) or (layer1_outputs(7599));
    layer2_outputs(429) <= not(layer1_outputs(7178));
    layer2_outputs(430) <= layer1_outputs(5186);
    layer2_outputs(431) <= layer1_outputs(2610);
    layer2_outputs(432) <= not((layer1_outputs(444)) xor (layer1_outputs(2690)));
    layer2_outputs(433) <= (layer1_outputs(6685)) and not (layer1_outputs(5559));
    layer2_outputs(434) <= (layer1_outputs(6859)) and (layer1_outputs(888));
    layer2_outputs(435) <= (layer1_outputs(5650)) or (layer1_outputs(5721));
    layer2_outputs(436) <= (layer1_outputs(590)) and not (layer1_outputs(912));
    layer2_outputs(437) <= layer1_outputs(4918);
    layer2_outputs(438) <= not((layer1_outputs(1864)) and (layer1_outputs(6057)));
    layer2_outputs(439) <= not((layer1_outputs(7169)) or (layer1_outputs(2392)));
    layer2_outputs(440) <= not(layer1_outputs(6829)) or (layer1_outputs(1058));
    layer2_outputs(441) <= (layer1_outputs(2830)) and not (layer1_outputs(6186));
    layer2_outputs(442) <= layer1_outputs(2100);
    layer2_outputs(443) <= (layer1_outputs(503)) and not (layer1_outputs(1239));
    layer2_outputs(444) <= layer1_outputs(5811);
    layer2_outputs(445) <= not(layer1_outputs(4001));
    layer2_outputs(446) <= layer1_outputs(5771);
    layer2_outputs(447) <= layer1_outputs(6874);
    layer2_outputs(448) <= not(layer1_outputs(5165)) or (layer1_outputs(5432));
    layer2_outputs(449) <= not(layer1_outputs(5446)) or (layer1_outputs(5474));
    layer2_outputs(450) <= (layer1_outputs(3663)) and not (layer1_outputs(2496));
    layer2_outputs(451) <= not(layer1_outputs(2503));
    layer2_outputs(452) <= not(layer1_outputs(315));
    layer2_outputs(453) <= layer1_outputs(2635);
    layer2_outputs(454) <= layer1_outputs(6743);
    layer2_outputs(455) <= (layer1_outputs(5414)) and (layer1_outputs(6876));
    layer2_outputs(456) <= not(layer1_outputs(5087));
    layer2_outputs(457) <= not((layer1_outputs(7031)) and (layer1_outputs(7367)));
    layer2_outputs(458) <= not(layer1_outputs(4144));
    layer2_outputs(459) <= layer1_outputs(5255);
    layer2_outputs(460) <= layer1_outputs(3552);
    layer2_outputs(461) <= not(layer1_outputs(5234));
    layer2_outputs(462) <= not(layer1_outputs(4372));
    layer2_outputs(463) <= layer1_outputs(5116);
    layer2_outputs(464) <= layer1_outputs(5371);
    layer2_outputs(465) <= not(layer1_outputs(2801));
    layer2_outputs(466) <= not(layer1_outputs(409));
    layer2_outputs(467) <= not(layer1_outputs(6917));
    layer2_outputs(468) <= layer1_outputs(479);
    layer2_outputs(469) <= not(layer1_outputs(2715)) or (layer1_outputs(5991));
    layer2_outputs(470) <= (layer1_outputs(6984)) and not (layer1_outputs(910));
    layer2_outputs(471) <= not(layer1_outputs(3665));
    layer2_outputs(472) <= not(layer1_outputs(2485)) or (layer1_outputs(6005));
    layer2_outputs(473) <= not(layer1_outputs(5149));
    layer2_outputs(474) <= '1';
    layer2_outputs(475) <= (layer1_outputs(1059)) or (layer1_outputs(229));
    layer2_outputs(476) <= not(layer1_outputs(5110)) or (layer1_outputs(3138));
    layer2_outputs(477) <= not((layer1_outputs(6233)) and (layer1_outputs(3286)));
    layer2_outputs(478) <= not((layer1_outputs(6002)) and (layer1_outputs(6062)));
    layer2_outputs(479) <= not((layer1_outputs(1099)) or (layer1_outputs(5959)));
    layer2_outputs(480) <= (layer1_outputs(1718)) and not (layer1_outputs(7011));
    layer2_outputs(481) <= (layer1_outputs(2715)) and (layer1_outputs(2034));
    layer2_outputs(482) <= (layer1_outputs(693)) or (layer1_outputs(5278));
    layer2_outputs(483) <= (layer1_outputs(3252)) and not (layer1_outputs(4361));
    layer2_outputs(484) <= layer1_outputs(985);
    layer2_outputs(485) <= (layer1_outputs(1913)) and not (layer1_outputs(278));
    layer2_outputs(486) <= '0';
    layer2_outputs(487) <= not((layer1_outputs(6848)) and (layer1_outputs(3061)));
    layer2_outputs(488) <= (layer1_outputs(5031)) and not (layer1_outputs(4497));
    layer2_outputs(489) <= (layer1_outputs(410)) and not (layer1_outputs(951));
    layer2_outputs(490) <= (layer1_outputs(207)) and not (layer1_outputs(5501));
    layer2_outputs(491) <= '1';
    layer2_outputs(492) <= (layer1_outputs(6162)) or (layer1_outputs(6421));
    layer2_outputs(493) <= not(layer1_outputs(7551));
    layer2_outputs(494) <= not(layer1_outputs(1692));
    layer2_outputs(495) <= layer1_outputs(5629);
    layer2_outputs(496) <= not(layer1_outputs(6194)) or (layer1_outputs(4140));
    layer2_outputs(497) <= not(layer1_outputs(3311)) or (layer1_outputs(6519));
    layer2_outputs(498) <= not((layer1_outputs(1440)) and (layer1_outputs(1372)));
    layer2_outputs(499) <= not(layer1_outputs(1165));
    layer2_outputs(500) <= not((layer1_outputs(6106)) and (layer1_outputs(211)));
    layer2_outputs(501) <= layer1_outputs(5128);
    layer2_outputs(502) <= not(layer1_outputs(325));
    layer2_outputs(503) <= not((layer1_outputs(2470)) or (layer1_outputs(1770)));
    layer2_outputs(504) <= (layer1_outputs(1560)) and not (layer1_outputs(4654));
    layer2_outputs(505) <= not(layer1_outputs(4109)) or (layer1_outputs(1954));
    layer2_outputs(506) <= '0';
    layer2_outputs(507) <= layer1_outputs(554);
    layer2_outputs(508) <= layer1_outputs(7013);
    layer2_outputs(509) <= (layer1_outputs(696)) or (layer1_outputs(291));
    layer2_outputs(510) <= (layer1_outputs(2976)) and not (layer1_outputs(795));
    layer2_outputs(511) <= (layer1_outputs(3044)) xor (layer1_outputs(3470));
    layer2_outputs(512) <= not(layer1_outputs(6634));
    layer2_outputs(513) <= (layer1_outputs(7618)) and not (layer1_outputs(7449));
    layer2_outputs(514) <= (layer1_outputs(5808)) and (layer1_outputs(4866));
    layer2_outputs(515) <= '1';
    layer2_outputs(516) <= layer1_outputs(706);
    layer2_outputs(517) <= layer1_outputs(3323);
    layer2_outputs(518) <= (layer1_outputs(157)) or (layer1_outputs(22));
    layer2_outputs(519) <= (layer1_outputs(3003)) and (layer1_outputs(4633));
    layer2_outputs(520) <= (layer1_outputs(3677)) xor (layer1_outputs(1071));
    layer2_outputs(521) <= not(layer1_outputs(3621));
    layer2_outputs(522) <= '1';
    layer2_outputs(523) <= (layer1_outputs(4488)) and not (layer1_outputs(6673));
    layer2_outputs(524) <= not((layer1_outputs(7545)) or (layer1_outputs(1854)));
    layer2_outputs(525) <= (layer1_outputs(5860)) and not (layer1_outputs(1904));
    layer2_outputs(526) <= (layer1_outputs(3618)) xor (layer1_outputs(2091));
    layer2_outputs(527) <= not(layer1_outputs(4720)) or (layer1_outputs(2612));
    layer2_outputs(528) <= (layer1_outputs(2433)) and not (layer1_outputs(2878));
    layer2_outputs(529) <= layer1_outputs(1808);
    layer2_outputs(530) <= not(layer1_outputs(3468));
    layer2_outputs(531) <= not(layer1_outputs(5736));
    layer2_outputs(532) <= not((layer1_outputs(2792)) or (layer1_outputs(6679)));
    layer2_outputs(533) <= (layer1_outputs(2218)) and (layer1_outputs(5224));
    layer2_outputs(534) <= (layer1_outputs(2796)) or (layer1_outputs(6616));
    layer2_outputs(535) <= layer1_outputs(2513);
    layer2_outputs(536) <= not(layer1_outputs(3807));
    layer2_outputs(537) <= not(layer1_outputs(7639));
    layer2_outputs(538) <= not(layer1_outputs(7034)) or (layer1_outputs(3668));
    layer2_outputs(539) <= (layer1_outputs(897)) and not (layer1_outputs(749));
    layer2_outputs(540) <= (layer1_outputs(3385)) or (layer1_outputs(3685));
    layer2_outputs(541) <= '1';
    layer2_outputs(542) <= not(layer1_outputs(6576)) or (layer1_outputs(1920));
    layer2_outputs(543) <= (layer1_outputs(1917)) and not (layer1_outputs(6369));
    layer2_outputs(544) <= not(layer1_outputs(6042)) or (layer1_outputs(4921));
    layer2_outputs(545) <= not((layer1_outputs(3186)) xor (layer1_outputs(5958)));
    layer2_outputs(546) <= (layer1_outputs(119)) and (layer1_outputs(4823));
    layer2_outputs(547) <= not(layer1_outputs(5806)) or (layer1_outputs(1184));
    layer2_outputs(548) <= not(layer1_outputs(5392)) or (layer1_outputs(5550));
    layer2_outputs(549) <= (layer1_outputs(4173)) or (layer1_outputs(4074));
    layer2_outputs(550) <= not(layer1_outputs(623)) or (layer1_outputs(5677));
    layer2_outputs(551) <= (layer1_outputs(1622)) and not (layer1_outputs(4484));
    layer2_outputs(552) <= not(layer1_outputs(2557));
    layer2_outputs(553) <= not(layer1_outputs(264)) or (layer1_outputs(499));
    layer2_outputs(554) <= not((layer1_outputs(6290)) or (layer1_outputs(7311)));
    layer2_outputs(555) <= not(layer1_outputs(4839)) or (layer1_outputs(6937));
    layer2_outputs(556) <= not(layer1_outputs(2995));
    layer2_outputs(557) <= (layer1_outputs(6435)) or (layer1_outputs(3639));
    layer2_outputs(558) <= '1';
    layer2_outputs(559) <= (layer1_outputs(6682)) and (layer1_outputs(3302));
    layer2_outputs(560) <= (layer1_outputs(649)) or (layer1_outputs(3399));
    layer2_outputs(561) <= layer1_outputs(6173);
    layer2_outputs(562) <= layer1_outputs(6884);
    layer2_outputs(563) <= (layer1_outputs(6281)) and not (layer1_outputs(2279));
    layer2_outputs(564) <= not(layer1_outputs(4561));
    layer2_outputs(565) <= layer1_outputs(6182);
    layer2_outputs(566) <= layer1_outputs(3231);
    layer2_outputs(567) <= not((layer1_outputs(7497)) and (layer1_outputs(2582)));
    layer2_outputs(568) <= layer1_outputs(3520);
    layer2_outputs(569) <= not((layer1_outputs(4098)) or (layer1_outputs(95)));
    layer2_outputs(570) <= layer1_outputs(3526);
    layer2_outputs(571) <= layer1_outputs(124);
    layer2_outputs(572) <= not(layer1_outputs(1934));
    layer2_outputs(573) <= not(layer1_outputs(6487));
    layer2_outputs(574) <= (layer1_outputs(5167)) and not (layer1_outputs(2321));
    layer2_outputs(575) <= (layer1_outputs(6568)) and not (layer1_outputs(7634));
    layer2_outputs(576) <= '1';
    layer2_outputs(577) <= (layer1_outputs(2990)) or (layer1_outputs(2714));
    layer2_outputs(578) <= layer1_outputs(3597);
    layer2_outputs(579) <= not((layer1_outputs(4919)) and (layer1_outputs(5629)));
    layer2_outputs(580) <= not((layer1_outputs(713)) xor (layer1_outputs(4142)));
    layer2_outputs(581) <= not(layer1_outputs(435)) or (layer1_outputs(5337));
    layer2_outputs(582) <= not(layer1_outputs(4942));
    layer2_outputs(583) <= layer1_outputs(2698);
    layer2_outputs(584) <= not(layer1_outputs(7637));
    layer2_outputs(585) <= layer1_outputs(7236);
    layer2_outputs(586) <= (layer1_outputs(4519)) and (layer1_outputs(7082));
    layer2_outputs(587) <= not(layer1_outputs(4018));
    layer2_outputs(588) <= layer1_outputs(7127);
    layer2_outputs(589) <= layer1_outputs(2687);
    layer2_outputs(590) <= not(layer1_outputs(3826));
    layer2_outputs(591) <= (layer1_outputs(1387)) and not (layer1_outputs(5938));
    layer2_outputs(592) <= not((layer1_outputs(1649)) or (layer1_outputs(3538)));
    layer2_outputs(593) <= not(layer1_outputs(46));
    layer2_outputs(594) <= not((layer1_outputs(2982)) and (layer1_outputs(7530)));
    layer2_outputs(595) <= not(layer1_outputs(7483));
    layer2_outputs(596) <= not(layer1_outputs(2116));
    layer2_outputs(597) <= (layer1_outputs(3262)) and not (layer1_outputs(6326));
    layer2_outputs(598) <= not(layer1_outputs(1411));
    layer2_outputs(599) <= '1';
    layer2_outputs(600) <= (layer1_outputs(2695)) and (layer1_outputs(792));
    layer2_outputs(601) <= '0';
    layer2_outputs(602) <= layer1_outputs(3938);
    layer2_outputs(603) <= not((layer1_outputs(7544)) xor (layer1_outputs(4121)));
    layer2_outputs(604) <= layer1_outputs(6253);
    layer2_outputs(605) <= (layer1_outputs(5176)) and (layer1_outputs(4404));
    layer2_outputs(606) <= not(layer1_outputs(6993));
    layer2_outputs(607) <= not((layer1_outputs(5369)) or (layer1_outputs(1885)));
    layer2_outputs(608) <= (layer1_outputs(5547)) and not (layer1_outputs(6408));
    layer2_outputs(609) <= layer1_outputs(5376);
    layer2_outputs(610) <= not((layer1_outputs(4680)) or (layer1_outputs(1046)));
    layer2_outputs(611) <= not(layer1_outputs(772));
    layer2_outputs(612) <= not(layer1_outputs(4423)) or (layer1_outputs(2059));
    layer2_outputs(613) <= '1';
    layer2_outputs(614) <= (layer1_outputs(6803)) and not (layer1_outputs(905));
    layer2_outputs(615) <= '1';
    layer2_outputs(616) <= not(layer1_outputs(6837)) or (layer1_outputs(5600));
    layer2_outputs(617) <= not(layer1_outputs(4067)) or (layer1_outputs(4628));
    layer2_outputs(618) <= (layer1_outputs(1834)) and (layer1_outputs(7175));
    layer2_outputs(619) <= (layer1_outputs(2016)) and (layer1_outputs(25));
    layer2_outputs(620) <= layer1_outputs(7532);
    layer2_outputs(621) <= (layer1_outputs(3668)) and (layer1_outputs(3387));
    layer2_outputs(622) <= not(layer1_outputs(273));
    layer2_outputs(623) <= (layer1_outputs(602)) and not (layer1_outputs(1534));
    layer2_outputs(624) <= not((layer1_outputs(3366)) and (layer1_outputs(2085)));
    layer2_outputs(625) <= layer1_outputs(238);
    layer2_outputs(626) <= not((layer1_outputs(5181)) xor (layer1_outputs(2828)));
    layer2_outputs(627) <= layer1_outputs(7589);
    layer2_outputs(628) <= layer1_outputs(4390);
    layer2_outputs(629) <= (layer1_outputs(6342)) or (layer1_outputs(7098));
    layer2_outputs(630) <= not(layer1_outputs(1496));
    layer2_outputs(631) <= (layer1_outputs(5532)) and not (layer1_outputs(1234));
    layer2_outputs(632) <= layer1_outputs(5675);
    layer2_outputs(633) <= not((layer1_outputs(792)) or (layer1_outputs(2113)));
    layer2_outputs(634) <= not(layer1_outputs(6971));
    layer2_outputs(635) <= (layer1_outputs(6502)) and not (layer1_outputs(3080));
    layer2_outputs(636) <= '1';
    layer2_outputs(637) <= not(layer1_outputs(4876));
    layer2_outputs(638) <= (layer1_outputs(2914)) or (layer1_outputs(280));
    layer2_outputs(639) <= '0';
    layer2_outputs(640) <= not((layer1_outputs(569)) and (layer1_outputs(2175)));
    layer2_outputs(641) <= '1';
    layer2_outputs(642) <= not(layer1_outputs(3068));
    layer2_outputs(643) <= (layer1_outputs(1120)) and (layer1_outputs(6785));
    layer2_outputs(644) <= '0';
    layer2_outputs(645) <= layer1_outputs(2664);
    layer2_outputs(646) <= layer1_outputs(2172);
    layer2_outputs(647) <= '1';
    layer2_outputs(648) <= not(layer1_outputs(6074));
    layer2_outputs(649) <= (layer1_outputs(5684)) and not (layer1_outputs(2957));
    layer2_outputs(650) <= layer1_outputs(3689);
    layer2_outputs(651) <= (layer1_outputs(4027)) and (layer1_outputs(5090));
    layer2_outputs(652) <= not(layer1_outputs(2010));
    layer2_outputs(653) <= not((layer1_outputs(4661)) or (layer1_outputs(2744)));
    layer2_outputs(654) <= layer1_outputs(4687);
    layer2_outputs(655) <= (layer1_outputs(5915)) or (layer1_outputs(6274));
    layer2_outputs(656) <= (layer1_outputs(123)) and not (layer1_outputs(7199));
    layer2_outputs(657) <= layer1_outputs(2948);
    layer2_outputs(658) <= not(layer1_outputs(5642));
    layer2_outputs(659) <= layer1_outputs(1774);
    layer2_outputs(660) <= not((layer1_outputs(2290)) and (layer1_outputs(3416)));
    layer2_outputs(661) <= (layer1_outputs(3605)) and not (layer1_outputs(6893));
    layer2_outputs(662) <= layer1_outputs(530);
    layer2_outputs(663) <= (layer1_outputs(6400)) and (layer1_outputs(371));
    layer2_outputs(664) <= not(layer1_outputs(1232)) or (layer1_outputs(1028));
    layer2_outputs(665) <= not((layer1_outputs(1623)) and (layer1_outputs(5322)));
    layer2_outputs(666) <= not(layer1_outputs(2598));
    layer2_outputs(667) <= layer1_outputs(508);
    layer2_outputs(668) <= not(layer1_outputs(1143)) or (layer1_outputs(1671));
    layer2_outputs(669) <= '1';
    layer2_outputs(670) <= layer1_outputs(4940);
    layer2_outputs(671) <= '0';
    layer2_outputs(672) <= not(layer1_outputs(64)) or (layer1_outputs(1953));
    layer2_outputs(673) <= not(layer1_outputs(57));
    layer2_outputs(674) <= not((layer1_outputs(5586)) xor (layer1_outputs(6373)));
    layer2_outputs(675) <= (layer1_outputs(6073)) and not (layer1_outputs(6090));
    layer2_outputs(676) <= not((layer1_outputs(4040)) xor (layer1_outputs(5241)));
    layer2_outputs(677) <= not(layer1_outputs(3611)) or (layer1_outputs(6164));
    layer2_outputs(678) <= not(layer1_outputs(3899));
    layer2_outputs(679) <= not((layer1_outputs(146)) and (layer1_outputs(2021)));
    layer2_outputs(680) <= not(layer1_outputs(2078));
    layer2_outputs(681) <= (layer1_outputs(3398)) or (layer1_outputs(4451));
    layer2_outputs(682) <= layer1_outputs(3942);
    layer2_outputs(683) <= layer1_outputs(7403);
    layer2_outputs(684) <= layer1_outputs(2912);
    layer2_outputs(685) <= (layer1_outputs(5676)) and not (layer1_outputs(7216));
    layer2_outputs(686) <= not(layer1_outputs(1422)) or (layer1_outputs(549));
    layer2_outputs(687) <= not(layer1_outputs(7575));
    layer2_outputs(688) <= not(layer1_outputs(4656)) or (layer1_outputs(2607));
    layer2_outputs(689) <= not(layer1_outputs(899)) or (layer1_outputs(4821));
    layer2_outputs(690) <= (layer1_outputs(3700)) and (layer1_outputs(917));
    layer2_outputs(691) <= (layer1_outputs(2776)) and (layer1_outputs(5223));
    layer2_outputs(692) <= not(layer1_outputs(5778)) or (layer1_outputs(132));
    layer2_outputs(693) <= not(layer1_outputs(2025));
    layer2_outputs(694) <= (layer1_outputs(2216)) and not (layer1_outputs(3162));
    layer2_outputs(695) <= layer1_outputs(3875);
    layer2_outputs(696) <= not(layer1_outputs(7565)) or (layer1_outputs(2106));
    layer2_outputs(697) <= not((layer1_outputs(4833)) or (layer1_outputs(6953)));
    layer2_outputs(698) <= (layer1_outputs(2959)) or (layer1_outputs(3900));
    layer2_outputs(699) <= not(layer1_outputs(5898)) or (layer1_outputs(7007));
    layer2_outputs(700) <= layer1_outputs(7261);
    layer2_outputs(701) <= not(layer1_outputs(4787));
    layer2_outputs(702) <= not((layer1_outputs(5336)) and (layer1_outputs(940)));
    layer2_outputs(703) <= layer1_outputs(3650);
    layer2_outputs(704) <= not(layer1_outputs(3260));
    layer2_outputs(705) <= not((layer1_outputs(3272)) or (layer1_outputs(3840)));
    layer2_outputs(706) <= (layer1_outputs(59)) and (layer1_outputs(2031));
    layer2_outputs(707) <= not(layer1_outputs(3066));
    layer2_outputs(708) <= not(layer1_outputs(1771));
    layer2_outputs(709) <= not(layer1_outputs(1910));
    layer2_outputs(710) <= not(layer1_outputs(1456)) or (layer1_outputs(4320));
    layer2_outputs(711) <= not(layer1_outputs(5911));
    layer2_outputs(712) <= layer1_outputs(5142);
    layer2_outputs(713) <= layer1_outputs(685);
    layer2_outputs(714) <= (layer1_outputs(6867)) and not (layer1_outputs(4750));
    layer2_outputs(715) <= not(layer1_outputs(3317)) or (layer1_outputs(7084));
    layer2_outputs(716) <= not(layer1_outputs(1733));
    layer2_outputs(717) <= layer1_outputs(6717);
    layer2_outputs(718) <= not(layer1_outputs(6051)) or (layer1_outputs(3843));
    layer2_outputs(719) <= (layer1_outputs(7125)) and not (layer1_outputs(6330));
    layer2_outputs(720) <= (layer1_outputs(2253)) or (layer1_outputs(6544));
    layer2_outputs(721) <= (layer1_outputs(4600)) and not (layer1_outputs(2507));
    layer2_outputs(722) <= layer1_outputs(1016);
    layer2_outputs(723) <= not(layer1_outputs(3301)) or (layer1_outputs(3012));
    layer2_outputs(724) <= layer1_outputs(7101);
    layer2_outputs(725) <= not(layer1_outputs(4598)) or (layer1_outputs(3696));
    layer2_outputs(726) <= (layer1_outputs(4106)) and (layer1_outputs(4777));
    layer2_outputs(727) <= layer1_outputs(7401);
    layer2_outputs(728) <= '0';
    layer2_outputs(729) <= layer1_outputs(5044);
    layer2_outputs(730) <= not(layer1_outputs(2960)) or (layer1_outputs(1822));
    layer2_outputs(731) <= (layer1_outputs(5689)) and not (layer1_outputs(3564));
    layer2_outputs(732) <= (layer1_outputs(1277)) and (layer1_outputs(315));
    layer2_outputs(733) <= not((layer1_outputs(1759)) and (layer1_outputs(3764)));
    layer2_outputs(734) <= layer1_outputs(2494);
    layer2_outputs(735) <= (layer1_outputs(2434)) and (layer1_outputs(1329));
    layer2_outputs(736) <= (layer1_outputs(3463)) xor (layer1_outputs(2046));
    layer2_outputs(737) <= not((layer1_outputs(3610)) xor (layer1_outputs(676)));
    layer2_outputs(738) <= (layer1_outputs(5583)) and not (layer1_outputs(1999));
    layer2_outputs(739) <= layer1_outputs(7088);
    layer2_outputs(740) <= not(layer1_outputs(5698));
    layer2_outputs(741) <= not(layer1_outputs(4390)) or (layer1_outputs(5286));
    layer2_outputs(742) <= '0';
    layer2_outputs(743) <= not(layer1_outputs(3108));
    layer2_outputs(744) <= not((layer1_outputs(7304)) and (layer1_outputs(3539)));
    layer2_outputs(745) <= layer1_outputs(4428);
    layer2_outputs(746) <= layer1_outputs(738);
    layer2_outputs(747) <= layer1_outputs(818);
    layer2_outputs(748) <= '1';
    layer2_outputs(749) <= (layer1_outputs(7475)) and not (layer1_outputs(1991));
    layer2_outputs(750) <= layer1_outputs(5458);
    layer2_outputs(751) <= layer1_outputs(48);
    layer2_outputs(752) <= (layer1_outputs(5578)) and not (layer1_outputs(4061));
    layer2_outputs(753) <= not(layer1_outputs(2578));
    layer2_outputs(754) <= not(layer1_outputs(1753));
    layer2_outputs(755) <= (layer1_outputs(4888)) and (layer1_outputs(4491));
    layer2_outputs(756) <= not(layer1_outputs(6272));
    layer2_outputs(757) <= not(layer1_outputs(2457));
    layer2_outputs(758) <= not(layer1_outputs(5966)) or (layer1_outputs(1211));
    layer2_outputs(759) <= layer1_outputs(742);
    layer2_outputs(760) <= not(layer1_outputs(3201));
    layer2_outputs(761) <= '1';
    layer2_outputs(762) <= not(layer1_outputs(2533));
    layer2_outputs(763) <= layer1_outputs(3585);
    layer2_outputs(764) <= layer1_outputs(853);
    layer2_outputs(765) <= (layer1_outputs(1995)) and not (layer1_outputs(4005));
    layer2_outputs(766) <= layer1_outputs(2618);
    layer2_outputs(767) <= not((layer1_outputs(726)) or (layer1_outputs(4176)));
    layer2_outputs(768) <= layer1_outputs(2211);
    layer2_outputs(769) <= (layer1_outputs(7598)) and (layer1_outputs(490));
    layer2_outputs(770) <= (layer1_outputs(4898)) and (layer1_outputs(1657));
    layer2_outputs(771) <= not(layer1_outputs(5595)) or (layer1_outputs(5160));
    layer2_outputs(772) <= layer1_outputs(5566);
    layer2_outputs(773) <= (layer1_outputs(3832)) xor (layer1_outputs(7144));
    layer2_outputs(774) <= not(layer1_outputs(2516)) or (layer1_outputs(7663));
    layer2_outputs(775) <= (layer1_outputs(2793)) and (layer1_outputs(3590));
    layer2_outputs(776) <= (layer1_outputs(6510)) and not (layer1_outputs(3940));
    layer2_outputs(777) <= not(layer1_outputs(4512));
    layer2_outputs(778) <= not((layer1_outputs(4075)) or (layer1_outputs(7333)));
    layer2_outputs(779) <= (layer1_outputs(5980)) and (layer1_outputs(1635));
    layer2_outputs(780) <= '0';
    layer2_outputs(781) <= not(layer1_outputs(5198)) or (layer1_outputs(1131));
    layer2_outputs(782) <= not(layer1_outputs(1350));
    layer2_outputs(783) <= not(layer1_outputs(5797));
    layer2_outputs(784) <= not(layer1_outputs(1674));
    layer2_outputs(785) <= not(layer1_outputs(4243));
    layer2_outputs(786) <= not(layer1_outputs(476));
    layer2_outputs(787) <= layer1_outputs(7494);
    layer2_outputs(788) <= layer1_outputs(4063);
    layer2_outputs(789) <= '1';
    layer2_outputs(790) <= not((layer1_outputs(6285)) or (layer1_outputs(753)));
    layer2_outputs(791) <= (layer1_outputs(6619)) and not (layer1_outputs(5170));
    layer2_outputs(792) <= not((layer1_outputs(2370)) and (layer1_outputs(7074)));
    layer2_outputs(793) <= not(layer1_outputs(5051)) or (layer1_outputs(1838));
    layer2_outputs(794) <= layer1_outputs(1648);
    layer2_outputs(795) <= layer1_outputs(6641);
    layer2_outputs(796) <= not(layer1_outputs(7242)) or (layer1_outputs(5873));
    layer2_outputs(797) <= (layer1_outputs(7226)) or (layer1_outputs(3956));
    layer2_outputs(798) <= not(layer1_outputs(5172)) or (layer1_outputs(3547));
    layer2_outputs(799) <= not((layer1_outputs(2272)) xor (layer1_outputs(385)));
    layer2_outputs(800) <= (layer1_outputs(6182)) and not (layer1_outputs(7111));
    layer2_outputs(801) <= not((layer1_outputs(3935)) or (layer1_outputs(267)));
    layer2_outputs(802) <= not(layer1_outputs(1339));
    layer2_outputs(803) <= (layer1_outputs(5812)) or (layer1_outputs(414));
    layer2_outputs(804) <= not(layer1_outputs(118));
    layer2_outputs(805) <= (layer1_outputs(980)) and not (layer1_outputs(1239));
    layer2_outputs(806) <= not((layer1_outputs(460)) or (layer1_outputs(3803)));
    layer2_outputs(807) <= (layer1_outputs(4087)) and (layer1_outputs(4049));
    layer2_outputs(808) <= not(layer1_outputs(3122)) or (layer1_outputs(1522));
    layer2_outputs(809) <= layer1_outputs(7401);
    layer2_outputs(810) <= layer1_outputs(3741);
    layer2_outputs(811) <= not(layer1_outputs(5941)) or (layer1_outputs(3729));
    layer2_outputs(812) <= not((layer1_outputs(7547)) or (layer1_outputs(2762)));
    layer2_outputs(813) <= not((layer1_outputs(3191)) and (layer1_outputs(257)));
    layer2_outputs(814) <= not((layer1_outputs(3974)) or (layer1_outputs(5323)));
    layer2_outputs(815) <= not(layer1_outputs(734));
    layer2_outputs(816) <= not((layer1_outputs(639)) and (layer1_outputs(3128)));
    layer2_outputs(817) <= layer1_outputs(5410);
    layer2_outputs(818) <= not(layer1_outputs(1598)) or (layer1_outputs(2774));
    layer2_outputs(819) <= '0';
    layer2_outputs(820) <= layer1_outputs(7161);
    layer2_outputs(821) <= not((layer1_outputs(6192)) and (layer1_outputs(2089)));
    layer2_outputs(822) <= not(layer1_outputs(84)) or (layer1_outputs(2769));
    layer2_outputs(823) <= layer1_outputs(5959);
    layer2_outputs(824) <= (layer1_outputs(6671)) and (layer1_outputs(5099));
    layer2_outputs(825) <= not((layer1_outputs(4078)) or (layer1_outputs(7107)));
    layer2_outputs(826) <= not(layer1_outputs(141));
    layer2_outputs(827) <= not(layer1_outputs(2407)) or (layer1_outputs(1313));
    layer2_outputs(828) <= not((layer1_outputs(3451)) and (layer1_outputs(1923)));
    layer2_outputs(829) <= layer1_outputs(7140);
    layer2_outputs(830) <= layer1_outputs(4666);
    layer2_outputs(831) <= layer1_outputs(6549);
    layer2_outputs(832) <= not(layer1_outputs(565));
    layer2_outputs(833) <= '0';
    layer2_outputs(834) <= not((layer1_outputs(3280)) and (layer1_outputs(3438)));
    layer2_outputs(835) <= not((layer1_outputs(765)) or (layer1_outputs(2373)));
    layer2_outputs(836) <= not(layer1_outputs(3472));
    layer2_outputs(837) <= not(layer1_outputs(6440));
    layer2_outputs(838) <= not((layer1_outputs(543)) and (layer1_outputs(5855)));
    layer2_outputs(839) <= not(layer1_outputs(433));
    layer2_outputs(840) <= '0';
    layer2_outputs(841) <= '0';
    layer2_outputs(842) <= layer1_outputs(1289);
    layer2_outputs(843) <= layer1_outputs(7027);
    layer2_outputs(844) <= not(layer1_outputs(5819)) or (layer1_outputs(867));
    layer2_outputs(845) <= not(layer1_outputs(4111));
    layer2_outputs(846) <= (layer1_outputs(5104)) and not (layer1_outputs(6550));
    layer2_outputs(847) <= (layer1_outputs(2304)) xor (layer1_outputs(4889));
    layer2_outputs(848) <= not(layer1_outputs(4830));
    layer2_outputs(849) <= not(layer1_outputs(2906)) or (layer1_outputs(1322));
    layer2_outputs(850) <= '0';
    layer2_outputs(851) <= layer1_outputs(3981);
    layer2_outputs(852) <= layer1_outputs(2137);
    layer2_outputs(853) <= (layer1_outputs(4790)) or (layer1_outputs(2031));
    layer2_outputs(854) <= not(layer1_outputs(3823)) or (layer1_outputs(822));
    layer2_outputs(855) <= not(layer1_outputs(294)) or (layer1_outputs(3422));
    layer2_outputs(856) <= not(layer1_outputs(2654)) or (layer1_outputs(4238));
    layer2_outputs(857) <= (layer1_outputs(1626)) xor (layer1_outputs(4679));
    layer2_outputs(858) <= not(layer1_outputs(2060));
    layer2_outputs(859) <= layer1_outputs(2014);
    layer2_outputs(860) <= not((layer1_outputs(158)) and (layer1_outputs(3204)));
    layer2_outputs(861) <= layer1_outputs(6290);
    layer2_outputs(862) <= not(layer1_outputs(1659));
    layer2_outputs(863) <= layer1_outputs(2336);
    layer2_outputs(864) <= not((layer1_outputs(5803)) and (layer1_outputs(6391)));
    layer2_outputs(865) <= layer1_outputs(2541);
    layer2_outputs(866) <= (layer1_outputs(7158)) and not (layer1_outputs(2435));
    layer2_outputs(867) <= (layer1_outputs(2915)) or (layer1_outputs(4800));
    layer2_outputs(868) <= not(layer1_outputs(3070)) or (layer1_outputs(625));
    layer2_outputs(869) <= '1';
    layer2_outputs(870) <= not(layer1_outputs(1966));
    layer2_outputs(871) <= not(layer1_outputs(2593));
    layer2_outputs(872) <= not(layer1_outputs(4139));
    layer2_outputs(873) <= layer1_outputs(4379);
    layer2_outputs(874) <= not(layer1_outputs(5627)) or (layer1_outputs(1004));
    layer2_outputs(875) <= not(layer1_outputs(4821));
    layer2_outputs(876) <= not(layer1_outputs(646));
    layer2_outputs(877) <= (layer1_outputs(7658)) and not (layer1_outputs(5126));
    layer2_outputs(878) <= not(layer1_outputs(7499)) or (layer1_outputs(1262));
    layer2_outputs(879) <= not(layer1_outputs(407));
    layer2_outputs(880) <= not(layer1_outputs(4144)) or (layer1_outputs(7105));
    layer2_outputs(881) <= (layer1_outputs(5666)) and (layer1_outputs(5661));
    layer2_outputs(882) <= layer1_outputs(5114);
    layer2_outputs(883) <= not(layer1_outputs(7050));
    layer2_outputs(884) <= layer1_outputs(3781);
    layer2_outputs(885) <= not((layer1_outputs(6429)) and (layer1_outputs(2592)));
    layer2_outputs(886) <= (layer1_outputs(6947)) and not (layer1_outputs(763));
    layer2_outputs(887) <= (layer1_outputs(6840)) and (layer1_outputs(2587));
    layer2_outputs(888) <= layer1_outputs(6205);
    layer2_outputs(889) <= not(layer1_outputs(5674)) or (layer1_outputs(2299));
    layer2_outputs(890) <= (layer1_outputs(308)) and not (layer1_outputs(6263));
    layer2_outputs(891) <= not(layer1_outputs(1772));
    layer2_outputs(892) <= not((layer1_outputs(4902)) xor (layer1_outputs(6704)));
    layer2_outputs(893) <= (layer1_outputs(5088)) and not (layer1_outputs(3373));
    layer2_outputs(894) <= not(layer1_outputs(2063));
    layer2_outputs(895) <= (layer1_outputs(4779)) and not (layer1_outputs(287));
    layer2_outputs(896) <= layer1_outputs(7301);
    layer2_outputs(897) <= not(layer1_outputs(3658));
    layer2_outputs(898) <= (layer1_outputs(7489)) and (layer1_outputs(290));
    layer2_outputs(899) <= (layer1_outputs(6577)) and (layer1_outputs(7252));
    layer2_outputs(900) <= (layer1_outputs(1867)) and (layer1_outputs(2760));
    layer2_outputs(901) <= (layer1_outputs(5950)) or (layer1_outputs(6759));
    layer2_outputs(902) <= not(layer1_outputs(914));
    layer2_outputs(903) <= not(layer1_outputs(439));
    layer2_outputs(904) <= not(layer1_outputs(72));
    layer2_outputs(905) <= not(layer1_outputs(5077));
    layer2_outputs(906) <= layer1_outputs(353);
    layer2_outputs(907) <= not(layer1_outputs(6905));
    layer2_outputs(908) <= not(layer1_outputs(2161));
    layer2_outputs(909) <= (layer1_outputs(6839)) xor (layer1_outputs(1914));
    layer2_outputs(910) <= (layer1_outputs(3336)) and not (layer1_outputs(1979));
    layer2_outputs(911) <= layer1_outputs(932);
    layer2_outputs(912) <= layer1_outputs(817);
    layer2_outputs(913) <= not(layer1_outputs(5682)) or (layer1_outputs(2136));
    layer2_outputs(914) <= not(layer1_outputs(2555));
    layer2_outputs(915) <= not(layer1_outputs(3338)) or (layer1_outputs(5210));
    layer2_outputs(916) <= '1';
    layer2_outputs(917) <= not(layer1_outputs(6153));
    layer2_outputs(918) <= not(layer1_outputs(2326));
    layer2_outputs(919) <= (layer1_outputs(1669)) xor (layer1_outputs(3108));
    layer2_outputs(920) <= (layer1_outputs(2323)) and (layer1_outputs(2055));
    layer2_outputs(921) <= layer1_outputs(171);
    layer2_outputs(922) <= layer1_outputs(3244);
    layer2_outputs(923) <= '1';
    layer2_outputs(924) <= layer1_outputs(6067);
    layer2_outputs(925) <= layer1_outputs(6527);
    layer2_outputs(926) <= layer1_outputs(1779);
    layer2_outputs(927) <= (layer1_outputs(905)) and (layer1_outputs(1119));
    layer2_outputs(928) <= not((layer1_outputs(1022)) and (layer1_outputs(6910)));
    layer2_outputs(929) <= not((layer1_outputs(839)) and (layer1_outputs(4282)));
    layer2_outputs(930) <= layer1_outputs(1876);
    layer2_outputs(931) <= not((layer1_outputs(1465)) and (layer1_outputs(3033)));
    layer2_outputs(932) <= '1';
    layer2_outputs(933) <= not(layer1_outputs(2762));
    layer2_outputs(934) <= not((layer1_outputs(1926)) or (layer1_outputs(515)));
    layer2_outputs(935) <= layer1_outputs(2211);
    layer2_outputs(936) <= (layer1_outputs(1128)) xor (layer1_outputs(1516));
    layer2_outputs(937) <= not(layer1_outputs(7670));
    layer2_outputs(938) <= not(layer1_outputs(1072));
    layer2_outputs(939) <= not(layer1_outputs(3247)) or (layer1_outputs(6610));
    layer2_outputs(940) <= (layer1_outputs(71)) or (layer1_outputs(2664));
    layer2_outputs(941) <= (layer1_outputs(2951)) and not (layer1_outputs(6331));
    layer2_outputs(942) <= not((layer1_outputs(611)) or (layer1_outputs(1533)));
    layer2_outputs(943) <= not((layer1_outputs(6303)) xor (layer1_outputs(5018)));
    layer2_outputs(944) <= not(layer1_outputs(2185)) or (layer1_outputs(6626));
    layer2_outputs(945) <= (layer1_outputs(7570)) or (layer1_outputs(2070));
    layer2_outputs(946) <= layer1_outputs(6321);
    layer2_outputs(947) <= not(layer1_outputs(2452));
    layer2_outputs(948) <= not(layer1_outputs(2998));
    layer2_outputs(949) <= not(layer1_outputs(7662)) or (layer1_outputs(1074));
    layer2_outputs(950) <= not((layer1_outputs(4709)) or (layer1_outputs(3281)));
    layer2_outputs(951) <= not((layer1_outputs(6385)) xor (layer1_outputs(187)));
    layer2_outputs(952) <= layer1_outputs(5516);
    layer2_outputs(953) <= (layer1_outputs(3558)) and not (layer1_outputs(7587));
    layer2_outputs(954) <= (layer1_outputs(2859)) and not (layer1_outputs(1405));
    layer2_outputs(955) <= layer1_outputs(5773);
    layer2_outputs(956) <= not((layer1_outputs(1292)) or (layer1_outputs(5746)));
    layer2_outputs(957) <= '1';
    layer2_outputs(958) <= layer1_outputs(263);
    layer2_outputs(959) <= not((layer1_outputs(1318)) or (layer1_outputs(6882)));
    layer2_outputs(960) <= (layer1_outputs(4758)) and not (layer1_outputs(6799));
    layer2_outputs(961) <= not(layer1_outputs(3009));
    layer2_outputs(962) <= (layer1_outputs(5669)) and not (layer1_outputs(7650));
    layer2_outputs(963) <= (layer1_outputs(6242)) or (layer1_outputs(5126));
    layer2_outputs(964) <= not(layer1_outputs(4677));
    layer2_outputs(965) <= layer1_outputs(6523);
    layer2_outputs(966) <= not(layer1_outputs(6401)) or (layer1_outputs(4958));
    layer2_outputs(967) <= not(layer1_outputs(4122));
    layer2_outputs(968) <= not((layer1_outputs(6703)) and (layer1_outputs(2592)));
    layer2_outputs(969) <= (layer1_outputs(1382)) and not (layer1_outputs(4973));
    layer2_outputs(970) <= not((layer1_outputs(2097)) or (layer1_outputs(4907)));
    layer2_outputs(971) <= '0';
    layer2_outputs(972) <= '0';
    layer2_outputs(973) <= not((layer1_outputs(7634)) or (layer1_outputs(5157)));
    layer2_outputs(974) <= '0';
    layer2_outputs(975) <= not(layer1_outputs(4258));
    layer2_outputs(976) <= not((layer1_outputs(1983)) or (layer1_outputs(1972)));
    layer2_outputs(977) <= not(layer1_outputs(3670));
    layer2_outputs(978) <= not(layer1_outputs(4899));
    layer2_outputs(979) <= '0';
    layer2_outputs(980) <= layer1_outputs(4452);
    layer2_outputs(981) <= not(layer1_outputs(1126));
    layer2_outputs(982) <= not(layer1_outputs(45));
    layer2_outputs(983) <= not(layer1_outputs(1530)) or (layer1_outputs(7573));
    layer2_outputs(984) <= (layer1_outputs(456)) and not (layer1_outputs(7007));
    layer2_outputs(985) <= not((layer1_outputs(2474)) or (layer1_outputs(2368)));
    layer2_outputs(986) <= not(layer1_outputs(1414));
    layer2_outputs(987) <= (layer1_outputs(1226)) and not (layer1_outputs(1441));
    layer2_outputs(988) <= layer1_outputs(5763);
    layer2_outputs(989) <= not(layer1_outputs(2720)) or (layer1_outputs(4545));
    layer2_outputs(990) <= not((layer1_outputs(4847)) xor (layer1_outputs(4679)));
    layer2_outputs(991) <= layer1_outputs(6857);
    layer2_outputs(992) <= '1';
    layer2_outputs(993) <= not(layer1_outputs(572)) or (layer1_outputs(892));
    layer2_outputs(994) <= not(layer1_outputs(3174));
    layer2_outputs(995) <= (layer1_outputs(125)) and not (layer1_outputs(4113));
    layer2_outputs(996) <= '0';
    layer2_outputs(997) <= not(layer1_outputs(1873));
    layer2_outputs(998) <= not((layer1_outputs(2854)) or (layer1_outputs(3788)));
    layer2_outputs(999) <= (layer1_outputs(6159)) and not (layer1_outputs(1809));
    layer2_outputs(1000) <= (layer1_outputs(161)) or (layer1_outputs(6560));
    layer2_outputs(1001) <= not(layer1_outputs(1256)) or (layer1_outputs(1185));
    layer2_outputs(1002) <= (layer1_outputs(6079)) and (layer1_outputs(1819));
    layer2_outputs(1003) <= layer1_outputs(6843);
    layer2_outputs(1004) <= layer1_outputs(6104);
    layer2_outputs(1005) <= layer1_outputs(303);
    layer2_outputs(1006) <= layer1_outputs(1600);
    layer2_outputs(1007) <= layer1_outputs(200);
    layer2_outputs(1008) <= (layer1_outputs(6890)) and (layer1_outputs(539));
    layer2_outputs(1009) <= layer1_outputs(6710);
    layer2_outputs(1010) <= (layer1_outputs(4332)) and not (layer1_outputs(597));
    layer2_outputs(1011) <= (layer1_outputs(3915)) and not (layer1_outputs(7326));
    layer2_outputs(1012) <= (layer1_outputs(2620)) and not (layer1_outputs(3755));
    layer2_outputs(1013) <= (layer1_outputs(6018)) and not (layer1_outputs(2446));
    layer2_outputs(1014) <= '0';
    layer2_outputs(1015) <= layer1_outputs(3524);
    layer2_outputs(1016) <= layer1_outputs(4861);
    layer2_outputs(1017) <= '0';
    layer2_outputs(1018) <= not((layer1_outputs(3428)) and (layer1_outputs(4434)));
    layer2_outputs(1019) <= not((layer1_outputs(6025)) or (layer1_outputs(7444)));
    layer2_outputs(1020) <= not(layer1_outputs(6066));
    layer2_outputs(1021) <= not((layer1_outputs(7004)) and (layer1_outputs(2325)));
    layer2_outputs(1022) <= not(layer1_outputs(3612));
    layer2_outputs(1023) <= not(layer1_outputs(4487));
    layer2_outputs(1024) <= (layer1_outputs(2478)) or (layer1_outputs(1721));
    layer2_outputs(1025) <= '1';
    layer2_outputs(1026) <= not(layer1_outputs(6745)) or (layer1_outputs(6064));
    layer2_outputs(1027) <= '0';
    layer2_outputs(1028) <= not(layer1_outputs(581));
    layer2_outputs(1029) <= not((layer1_outputs(5839)) and (layer1_outputs(4640)));
    layer2_outputs(1030) <= layer1_outputs(3710);
    layer2_outputs(1031) <= layer1_outputs(7142);
    layer2_outputs(1032) <= not(layer1_outputs(3354)) or (layer1_outputs(2836));
    layer2_outputs(1033) <= not(layer1_outputs(7582));
    layer2_outputs(1034) <= (layer1_outputs(3410)) or (layer1_outputs(5158));
    layer2_outputs(1035) <= (layer1_outputs(7286)) and (layer1_outputs(3670));
    layer2_outputs(1036) <= not(layer1_outputs(3476));
    layer2_outputs(1037) <= '1';
    layer2_outputs(1038) <= not((layer1_outputs(446)) or (layer1_outputs(809)));
    layer2_outputs(1039) <= not(layer1_outputs(4696));
    layer2_outputs(1040) <= layer1_outputs(2064);
    layer2_outputs(1041) <= not(layer1_outputs(6726)) or (layer1_outputs(2045));
    layer2_outputs(1042) <= not(layer1_outputs(7575)) or (layer1_outputs(3875));
    layer2_outputs(1043) <= layer1_outputs(7438);
    layer2_outputs(1044) <= not(layer1_outputs(6881));
    layer2_outputs(1045) <= not(layer1_outputs(3320));
    layer2_outputs(1046) <= layer1_outputs(2705);
    layer2_outputs(1047) <= not(layer1_outputs(4013)) or (layer1_outputs(1374));
    layer2_outputs(1048) <= not(layer1_outputs(2781)) or (layer1_outputs(3563));
    layer2_outputs(1049) <= not(layer1_outputs(317)) or (layer1_outputs(2820));
    layer2_outputs(1050) <= (layer1_outputs(6838)) xor (layer1_outputs(705));
    layer2_outputs(1051) <= not(layer1_outputs(3572));
    layer2_outputs(1052) <= not(layer1_outputs(6078));
    layer2_outputs(1053) <= not((layer1_outputs(3337)) or (layer1_outputs(3028)));
    layer2_outputs(1054) <= '0';
    layer2_outputs(1055) <= not(layer1_outputs(4342)) or (layer1_outputs(3911));
    layer2_outputs(1056) <= not(layer1_outputs(7387)) or (layer1_outputs(421));
    layer2_outputs(1057) <= (layer1_outputs(6627)) and not (layer1_outputs(6810));
    layer2_outputs(1058) <= (layer1_outputs(5433)) xor (layer1_outputs(2570));
    layer2_outputs(1059) <= not(layer1_outputs(4624));
    layer2_outputs(1060) <= (layer1_outputs(1187)) or (layer1_outputs(2135));
    layer2_outputs(1061) <= not(layer1_outputs(2026));
    layer2_outputs(1062) <= not(layer1_outputs(6946));
    layer2_outputs(1063) <= layer1_outputs(5970);
    layer2_outputs(1064) <= (layer1_outputs(5729)) xor (layer1_outputs(2522));
    layer2_outputs(1065) <= not(layer1_outputs(3045)) or (layer1_outputs(4220));
    layer2_outputs(1066) <= not(layer1_outputs(44));
    layer2_outputs(1067) <= not(layer1_outputs(6437));
    layer2_outputs(1068) <= layer1_outputs(6640);
    layer2_outputs(1069) <= not((layer1_outputs(7141)) or (layer1_outputs(5768)));
    layer2_outputs(1070) <= not(layer1_outputs(429));
    layer2_outputs(1071) <= (layer1_outputs(1309)) and not (layer1_outputs(6855));
    layer2_outputs(1072) <= (layer1_outputs(965)) or (layer1_outputs(827));
    layer2_outputs(1073) <= not(layer1_outputs(7539)) or (layer1_outputs(2529));
    layer2_outputs(1074) <= not(layer1_outputs(4154)) or (layer1_outputs(4220));
    layer2_outputs(1075) <= not(layer1_outputs(4451));
    layer2_outputs(1076) <= not(layer1_outputs(7633)) or (layer1_outputs(2658));
    layer2_outputs(1077) <= not(layer1_outputs(7218));
    layer2_outputs(1078) <= not(layer1_outputs(4724));
    layer2_outputs(1079) <= layer1_outputs(77);
    layer2_outputs(1080) <= not(layer1_outputs(4389));
    layer2_outputs(1081) <= not(layer1_outputs(6460));
    layer2_outputs(1082) <= (layer1_outputs(4351)) xor (layer1_outputs(6588));
    layer2_outputs(1083) <= (layer1_outputs(5535)) and (layer1_outputs(4697));
    layer2_outputs(1084) <= not(layer1_outputs(6336));
    layer2_outputs(1085) <= not((layer1_outputs(626)) and (layer1_outputs(6166)));
    layer2_outputs(1086) <= '1';
    layer2_outputs(1087) <= not(layer1_outputs(3100));
    layer2_outputs(1088) <= (layer1_outputs(1431)) and (layer1_outputs(5259));
    layer2_outputs(1089) <= layer1_outputs(6780);
    layer2_outputs(1090) <= not(layer1_outputs(1561));
    layer2_outputs(1091) <= layer1_outputs(4919);
    layer2_outputs(1092) <= not(layer1_outputs(5723));
    layer2_outputs(1093) <= (layer1_outputs(3681)) and (layer1_outputs(4127));
    layer2_outputs(1094) <= not(layer1_outputs(7227)) or (layer1_outputs(1920));
    layer2_outputs(1095) <= not(layer1_outputs(6934)) or (layer1_outputs(7429));
    layer2_outputs(1096) <= layer1_outputs(1268);
    layer2_outputs(1097) <= not(layer1_outputs(7654)) or (layer1_outputs(3321));
    layer2_outputs(1098) <= layer1_outputs(2758);
    layer2_outputs(1099) <= not(layer1_outputs(5600)) or (layer1_outputs(3646));
    layer2_outputs(1100) <= not((layer1_outputs(4457)) or (layer1_outputs(7204)));
    layer2_outputs(1101) <= '0';
    layer2_outputs(1102) <= layer1_outputs(1996);
    layer2_outputs(1103) <= not((layer1_outputs(6411)) and (layer1_outputs(4190)));
    layer2_outputs(1104) <= layer1_outputs(762);
    layer2_outputs(1105) <= (layer1_outputs(6434)) or (layer1_outputs(1187));
    layer2_outputs(1106) <= (layer1_outputs(1638)) and (layer1_outputs(4265));
    layer2_outputs(1107) <= layer1_outputs(3086);
    layer2_outputs(1108) <= not(layer1_outputs(5211));
    layer2_outputs(1109) <= not((layer1_outputs(7264)) or (layer1_outputs(4342)));
    layer2_outputs(1110) <= not(layer1_outputs(80));
    layer2_outputs(1111) <= layer1_outputs(5272);
    layer2_outputs(1112) <= not(layer1_outputs(2816));
    layer2_outputs(1113) <= layer1_outputs(1025);
    layer2_outputs(1114) <= (layer1_outputs(2905)) or (layer1_outputs(5521));
    layer2_outputs(1115) <= (layer1_outputs(3001)) and (layer1_outputs(602));
    layer2_outputs(1116) <= not((layer1_outputs(3734)) or (layer1_outputs(6500)));
    layer2_outputs(1117) <= layer1_outputs(2600);
    layer2_outputs(1118) <= '1';
    layer2_outputs(1119) <= not((layer1_outputs(4782)) and (layer1_outputs(3219)));
    layer2_outputs(1120) <= (layer1_outputs(3835)) and (layer1_outputs(6341));
    layer2_outputs(1121) <= not((layer1_outputs(6467)) or (layer1_outputs(1203)));
    layer2_outputs(1122) <= not(layer1_outputs(6750));
    layer2_outputs(1123) <= not(layer1_outputs(4065));
    layer2_outputs(1124) <= not((layer1_outputs(4848)) and (layer1_outputs(335)));
    layer2_outputs(1125) <= not(layer1_outputs(5390));
    layer2_outputs(1126) <= layer1_outputs(5768);
    layer2_outputs(1127) <= not(layer1_outputs(2782));
    layer2_outputs(1128) <= (layer1_outputs(6804)) and (layer1_outputs(2235));
    layer2_outputs(1129) <= not(layer1_outputs(5361));
    layer2_outputs(1130) <= (layer1_outputs(6395)) and not (layer1_outputs(1531));
    layer2_outputs(1131) <= '0';
    layer2_outputs(1132) <= not(layer1_outputs(3931));
    layer2_outputs(1133) <= not(layer1_outputs(4078));
    layer2_outputs(1134) <= '1';
    layer2_outputs(1135) <= layer1_outputs(4307);
    layer2_outputs(1136) <= (layer1_outputs(2283)) and (layer1_outputs(4060));
    layer2_outputs(1137) <= layer1_outputs(3663);
    layer2_outputs(1138) <= not(layer1_outputs(7170)) or (layer1_outputs(6977));
    layer2_outputs(1139) <= (layer1_outputs(830)) xor (layer1_outputs(105));
    layer2_outputs(1140) <= not((layer1_outputs(5019)) and (layer1_outputs(2671)));
    layer2_outputs(1141) <= not(layer1_outputs(5286)) or (layer1_outputs(6357));
    layer2_outputs(1142) <= (layer1_outputs(6802)) and not (layer1_outputs(5079));
    layer2_outputs(1143) <= layer1_outputs(3231);
    layer2_outputs(1144) <= not(layer1_outputs(1369));
    layer2_outputs(1145) <= not((layer1_outputs(7048)) and (layer1_outputs(724)));
    layer2_outputs(1146) <= not(layer1_outputs(4398)) or (layer1_outputs(32));
    layer2_outputs(1147) <= not((layer1_outputs(4461)) and (layer1_outputs(2623)));
    layer2_outputs(1148) <= not(layer1_outputs(517)) or (layer1_outputs(7051));
    layer2_outputs(1149) <= (layer1_outputs(4000)) or (layer1_outputs(6563));
    layer2_outputs(1150) <= not(layer1_outputs(3304));
    layer2_outputs(1151) <= (layer1_outputs(6410)) and not (layer1_outputs(5512));
    layer2_outputs(1152) <= layer1_outputs(5355);
    layer2_outputs(1153) <= (layer1_outputs(6899)) and (layer1_outputs(49));
    layer2_outputs(1154) <= not(layer1_outputs(5309));
    layer2_outputs(1155) <= not(layer1_outputs(2600));
    layer2_outputs(1156) <= layer1_outputs(3517);
    layer2_outputs(1157) <= not(layer1_outputs(794)) or (layer1_outputs(5732));
    layer2_outputs(1158) <= (layer1_outputs(4715)) and not (layer1_outputs(5041));
    layer2_outputs(1159) <= (layer1_outputs(7548)) and not (layer1_outputs(4207));
    layer2_outputs(1160) <= not(layer1_outputs(5789));
    layer2_outputs(1161) <= layer1_outputs(2780);
    layer2_outputs(1162) <= '0';
    layer2_outputs(1163) <= layer1_outputs(267);
    layer2_outputs(1164) <= not(layer1_outputs(2269)) or (layer1_outputs(5713));
    layer2_outputs(1165) <= '0';
    layer2_outputs(1166) <= not((layer1_outputs(3676)) or (layer1_outputs(6561)));
    layer2_outputs(1167) <= (layer1_outputs(5739)) and not (layer1_outputs(4654));
    layer2_outputs(1168) <= '1';
    layer2_outputs(1169) <= layer1_outputs(2871);
    layer2_outputs(1170) <= layer1_outputs(1362);
    layer2_outputs(1171) <= (layer1_outputs(7461)) and not (layer1_outputs(58));
    layer2_outputs(1172) <= layer1_outputs(4393);
    layer2_outputs(1173) <= not(layer1_outputs(6101));
    layer2_outputs(1174) <= (layer1_outputs(1291)) or (layer1_outputs(3329));
    layer2_outputs(1175) <= not(layer1_outputs(154));
    layer2_outputs(1176) <= not(layer1_outputs(2689)) or (layer1_outputs(3968));
    layer2_outputs(1177) <= layer1_outputs(3112);
    layer2_outputs(1178) <= '1';
    layer2_outputs(1179) <= (layer1_outputs(7445)) and not (layer1_outputs(5039));
    layer2_outputs(1180) <= not(layer1_outputs(2568));
    layer2_outputs(1181) <= not((layer1_outputs(6439)) or (layer1_outputs(5499)));
    layer2_outputs(1182) <= not((layer1_outputs(4023)) and (layer1_outputs(2888)));
    layer2_outputs(1183) <= not(layer1_outputs(2289));
    layer2_outputs(1184) <= layer1_outputs(2424);
    layer2_outputs(1185) <= not(layer1_outputs(1217));
    layer2_outputs(1186) <= (layer1_outputs(459)) and not (layer1_outputs(4900));
    layer2_outputs(1187) <= not((layer1_outputs(6586)) and (layer1_outputs(1207)));
    layer2_outputs(1188) <= layer1_outputs(4543);
    layer2_outputs(1189) <= (layer1_outputs(4099)) xor (layer1_outputs(2974));
    layer2_outputs(1190) <= not(layer1_outputs(6069));
    layer2_outputs(1191) <= not(layer1_outputs(4823));
    layer2_outputs(1192) <= '1';
    layer2_outputs(1193) <= not((layer1_outputs(1379)) or (layer1_outputs(7292)));
    layer2_outputs(1194) <= layer1_outputs(3921);
    layer2_outputs(1195) <= not((layer1_outputs(6368)) and (layer1_outputs(4866)));
    layer2_outputs(1196) <= not(layer1_outputs(4309));
    layer2_outputs(1197) <= layer1_outputs(6559);
    layer2_outputs(1198) <= not(layer1_outputs(7145));
    layer2_outputs(1199) <= layer1_outputs(6553);
    layer2_outputs(1200) <= not((layer1_outputs(4321)) or (layer1_outputs(3426)));
    layer2_outputs(1201) <= (layer1_outputs(2353)) and not (layer1_outputs(4841));
    layer2_outputs(1202) <= (layer1_outputs(1778)) xor (layer1_outputs(3023));
    layer2_outputs(1203) <= '1';
    layer2_outputs(1204) <= layer1_outputs(3454);
    layer2_outputs(1205) <= layer1_outputs(1093);
    layer2_outputs(1206) <= layer1_outputs(6147);
    layer2_outputs(1207) <= '0';
    layer2_outputs(1208) <= not((layer1_outputs(2980)) or (layer1_outputs(1627)));
    layer2_outputs(1209) <= not(layer1_outputs(15)) or (layer1_outputs(5138));
    layer2_outputs(1210) <= layer1_outputs(3811);
    layer2_outputs(1211) <= (layer1_outputs(604)) xor (layer1_outputs(2303));
    layer2_outputs(1212) <= (layer1_outputs(4667)) and not (layer1_outputs(2858));
    layer2_outputs(1213) <= (layer1_outputs(6441)) and (layer1_outputs(6919));
    layer2_outputs(1214) <= (layer1_outputs(663)) and (layer1_outputs(1006));
    layer2_outputs(1215) <= not(layer1_outputs(5109)) or (layer1_outputs(6186));
    layer2_outputs(1216) <= not(layer1_outputs(6908));
    layer2_outputs(1217) <= layer1_outputs(7543);
    layer2_outputs(1218) <= layer1_outputs(1959);
    layer2_outputs(1219) <= not((layer1_outputs(4134)) xor (layer1_outputs(1458)));
    layer2_outputs(1220) <= layer1_outputs(2597);
    layer2_outputs(1221) <= not(layer1_outputs(6121));
    layer2_outputs(1222) <= layer1_outputs(7046);
    layer2_outputs(1223) <= not((layer1_outputs(6854)) or (layer1_outputs(7527)));
    layer2_outputs(1224) <= not((layer1_outputs(4500)) or (layer1_outputs(6397)));
    layer2_outputs(1225) <= layer1_outputs(2702);
    layer2_outputs(1226) <= '0';
    layer2_outputs(1227) <= (layer1_outputs(199)) or (layer1_outputs(5794));
    layer2_outputs(1228) <= (layer1_outputs(2170)) or (layer1_outputs(392));
    layer2_outputs(1229) <= layer1_outputs(6666);
    layer2_outputs(1230) <= not(layer1_outputs(3186)) or (layer1_outputs(1246));
    layer2_outputs(1231) <= '0';
    layer2_outputs(1232) <= layer1_outputs(1874);
    layer2_outputs(1233) <= not((layer1_outputs(3636)) or (layer1_outputs(7113)));
    layer2_outputs(1234) <= not((layer1_outputs(6859)) and (layer1_outputs(7508)));
    layer2_outputs(1235) <= '0';
    layer2_outputs(1236) <= layer1_outputs(4713);
    layer2_outputs(1237) <= not(layer1_outputs(6584));
    layer2_outputs(1238) <= not(layer1_outputs(2165));
    layer2_outputs(1239) <= not((layer1_outputs(3740)) and (layer1_outputs(3241)));
    layer2_outputs(1240) <= not((layer1_outputs(1714)) and (layer1_outputs(6771)));
    layer2_outputs(1241) <= layer1_outputs(1686);
    layer2_outputs(1242) <= not((layer1_outputs(47)) or (layer1_outputs(3953)));
    layer2_outputs(1243) <= (layer1_outputs(6960)) xor (layer1_outputs(136));
    layer2_outputs(1244) <= '0';
    layer2_outputs(1245) <= (layer1_outputs(5489)) or (layer1_outputs(4433));
    layer2_outputs(1246) <= layer1_outputs(589);
    layer2_outputs(1247) <= layer1_outputs(2362);
    layer2_outputs(1248) <= not(layer1_outputs(5378));
    layer2_outputs(1249) <= not((layer1_outputs(1041)) and (layer1_outputs(4913)));
    layer2_outputs(1250) <= (layer1_outputs(7060)) and not (layer1_outputs(4273));
    layer2_outputs(1251) <= not((layer1_outputs(6392)) or (layer1_outputs(4329)));
    layer2_outputs(1252) <= (layer1_outputs(3876)) and not (layer1_outputs(6758));
    layer2_outputs(1253) <= (layer1_outputs(3657)) and not (layer1_outputs(4522));
    layer2_outputs(1254) <= layer1_outputs(4770);
    layer2_outputs(1255) <= not(layer1_outputs(3492)) or (layer1_outputs(7623));
    layer2_outputs(1256) <= layer1_outputs(3806);
    layer2_outputs(1257) <= layer1_outputs(1213);
    layer2_outputs(1258) <= (layer1_outputs(5147)) and not (layer1_outputs(731));
    layer2_outputs(1259) <= not(layer1_outputs(362));
    layer2_outputs(1260) <= not(layer1_outputs(7229));
    layer2_outputs(1261) <= layer1_outputs(4969);
    layer2_outputs(1262) <= layer1_outputs(2988);
    layer2_outputs(1263) <= not(layer1_outputs(1057)) or (layer1_outputs(3804));
    layer2_outputs(1264) <= not(layer1_outputs(339)) or (layer1_outputs(7271));
    layer2_outputs(1265) <= not(layer1_outputs(798));
    layer2_outputs(1266) <= layer1_outputs(7340);
    layer2_outputs(1267) <= '1';
    layer2_outputs(1268) <= not(layer1_outputs(3661)) or (layer1_outputs(4643));
    layer2_outputs(1269) <= not(layer1_outputs(4549));
    layer2_outputs(1270) <= layer1_outputs(6325);
    layer2_outputs(1271) <= not(layer1_outputs(6169));
    layer2_outputs(1272) <= (layer1_outputs(7319)) and (layer1_outputs(1150));
    layer2_outputs(1273) <= layer1_outputs(3634);
    layer2_outputs(1274) <= (layer1_outputs(5249)) and not (layer1_outputs(1883));
    layer2_outputs(1275) <= layer1_outputs(1783);
    layer2_outputs(1276) <= '1';
    layer2_outputs(1277) <= not((layer1_outputs(40)) and (layer1_outputs(6100)));
    layer2_outputs(1278) <= layer1_outputs(7415);
    layer2_outputs(1279) <= not(layer1_outputs(7458));
    layer2_outputs(1280) <= not((layer1_outputs(1206)) or (layer1_outputs(2039)));
    layer2_outputs(1281) <= not(layer1_outputs(23));
    layer2_outputs(1282) <= not(layer1_outputs(3707)) or (layer1_outputs(4516));
    layer2_outputs(1283) <= '0';
    layer2_outputs(1284) <= not(layer1_outputs(6958)) or (layer1_outputs(4027));
    layer2_outputs(1285) <= not(layer1_outputs(5271));
    layer2_outputs(1286) <= layer1_outputs(2345);
    layer2_outputs(1287) <= (layer1_outputs(495)) and not (layer1_outputs(1286));
    layer2_outputs(1288) <= not(layer1_outputs(5242));
    layer2_outputs(1289) <= (layer1_outputs(4104)) or (layer1_outputs(1901));
    layer2_outputs(1290) <= layer1_outputs(1118);
    layer2_outputs(1291) <= (layer1_outputs(3857)) and (layer1_outputs(1677));
    layer2_outputs(1292) <= layer1_outputs(4781);
    layer2_outputs(1293) <= layer1_outputs(3127);
    layer2_outputs(1294) <= layer1_outputs(7462);
    layer2_outputs(1295) <= (layer1_outputs(6986)) and (layer1_outputs(6537));
    layer2_outputs(1296) <= not((layer1_outputs(113)) or (layer1_outputs(6927)));
    layer2_outputs(1297) <= layer1_outputs(6714);
    layer2_outputs(1298) <= '1';
    layer2_outputs(1299) <= (layer1_outputs(3887)) and (layer1_outputs(2745));
    layer2_outputs(1300) <= (layer1_outputs(3557)) xor (layer1_outputs(2506));
    layer2_outputs(1301) <= not((layer1_outputs(5613)) or (layer1_outputs(7407)));
    layer2_outputs(1302) <= layer1_outputs(850);
    layer2_outputs(1303) <= not((layer1_outputs(7389)) or (layer1_outputs(7596)));
    layer2_outputs(1304) <= (layer1_outputs(1854)) and not (layer1_outputs(3647));
    layer2_outputs(1305) <= '1';
    layer2_outputs(1306) <= layer1_outputs(5570);
    layer2_outputs(1307) <= (layer1_outputs(5086)) or (layer1_outputs(7164));
    layer2_outputs(1308) <= not((layer1_outputs(6779)) or (layer1_outputs(6207)));
    layer2_outputs(1309) <= layer1_outputs(108);
    layer2_outputs(1310) <= (layer1_outputs(6377)) and not (layer1_outputs(5709));
    layer2_outputs(1311) <= (layer1_outputs(33)) and not (layer1_outputs(3034));
    layer2_outputs(1312) <= not(layer1_outputs(945));
    layer2_outputs(1313) <= layer1_outputs(4986);
    layer2_outputs(1314) <= (layer1_outputs(1510)) and not (layer1_outputs(7143));
    layer2_outputs(1315) <= not(layer1_outputs(5067)) or (layer1_outputs(3188));
    layer2_outputs(1316) <= not(layer1_outputs(4458));
    layer2_outputs(1317) <= (layer1_outputs(3505)) xor (layer1_outputs(7491));
    layer2_outputs(1318) <= not(layer1_outputs(2000)) or (layer1_outputs(3141));
    layer2_outputs(1319) <= (layer1_outputs(6481)) and not (layer1_outputs(7099));
    layer2_outputs(1320) <= (layer1_outputs(4806)) xor (layer1_outputs(4058));
    layer2_outputs(1321) <= (layer1_outputs(2411)) and not (layer1_outputs(5040));
    layer2_outputs(1322) <= not(layer1_outputs(3203));
    layer2_outputs(1323) <= not((layer1_outputs(6572)) xor (layer1_outputs(3458)));
    layer2_outputs(1324) <= not(layer1_outputs(6288));
    layer2_outputs(1325) <= layer1_outputs(2605);
    layer2_outputs(1326) <= not(layer1_outputs(1118));
    layer2_outputs(1327) <= '0';
    layer2_outputs(1328) <= not((layer1_outputs(6049)) and (layer1_outputs(7157)));
    layer2_outputs(1329) <= (layer1_outputs(438)) and (layer1_outputs(546));
    layer2_outputs(1330) <= (layer1_outputs(3449)) and not (layer1_outputs(6378));
    layer2_outputs(1331) <= not(layer1_outputs(6)) or (layer1_outputs(5041));
    layer2_outputs(1332) <= not(layer1_outputs(3562));
    layer2_outputs(1333) <= (layer1_outputs(176)) and not (layer1_outputs(4536));
    layer2_outputs(1334) <= not(layer1_outputs(6525));
    layer2_outputs(1335) <= not(layer1_outputs(6979));
    layer2_outputs(1336) <= layer1_outputs(3025);
    layer2_outputs(1337) <= (layer1_outputs(781)) and not (layer1_outputs(986));
    layer2_outputs(1338) <= not(layer1_outputs(6999));
    layer2_outputs(1339) <= not(layer1_outputs(5970)) or (layer1_outputs(4259));
    layer2_outputs(1340) <= layer1_outputs(7602);
    layer2_outputs(1341) <= not((layer1_outputs(1377)) and (layer1_outputs(4819)));
    layer2_outputs(1342) <= not(layer1_outputs(5468));
    layer2_outputs(1343) <= layer1_outputs(3982);
    layer2_outputs(1344) <= not((layer1_outputs(6446)) or (layer1_outputs(2783)));
    layer2_outputs(1345) <= not((layer1_outputs(2319)) or (layer1_outputs(1714)));
    layer2_outputs(1346) <= layer1_outputs(4922);
    layer2_outputs(1347) <= layer1_outputs(5713);
    layer2_outputs(1348) <= not(layer1_outputs(1143)) or (layer1_outputs(3336));
    layer2_outputs(1349) <= layer1_outputs(1354);
    layer2_outputs(1350) <= not(layer1_outputs(608));
    layer2_outputs(1351) <= (layer1_outputs(2280)) and not (layer1_outputs(3407));
    layer2_outputs(1352) <= not(layer1_outputs(3110)) or (layer1_outputs(6044));
    layer2_outputs(1353) <= (layer1_outputs(4531)) and not (layer1_outputs(396));
    layer2_outputs(1354) <= (layer1_outputs(4857)) and not (layer1_outputs(567));
    layer2_outputs(1355) <= layer1_outputs(6027);
    layer2_outputs(1356) <= not(layer1_outputs(4518));
    layer2_outputs(1357) <= (layer1_outputs(4462)) or (layer1_outputs(975));
    layer2_outputs(1358) <= layer1_outputs(6217);
    layer2_outputs(1359) <= not((layer1_outputs(5539)) xor (layer1_outputs(674)));
    layer2_outputs(1360) <= layer1_outputs(4303);
    layer2_outputs(1361) <= layer1_outputs(7344);
    layer2_outputs(1362) <= not((layer1_outputs(5569)) or (layer1_outputs(5270)));
    layer2_outputs(1363) <= not(layer1_outputs(1401)) or (layer1_outputs(1351));
    layer2_outputs(1364) <= not(layer1_outputs(157)) or (layer1_outputs(1737));
    layer2_outputs(1365) <= '1';
    layer2_outputs(1366) <= not(layer1_outputs(5431));
    layer2_outputs(1367) <= not(layer1_outputs(7502));
    layer2_outputs(1368) <= not(layer1_outputs(1001)) or (layer1_outputs(5583));
    layer2_outputs(1369) <= not(layer1_outputs(7411)) or (layer1_outputs(942));
    layer2_outputs(1370) <= not(layer1_outputs(4503));
    layer2_outputs(1371) <= (layer1_outputs(7665)) xor (layer1_outputs(6171));
    layer2_outputs(1372) <= (layer1_outputs(1955)) and (layer1_outputs(7154));
    layer2_outputs(1373) <= not(layer1_outputs(4486));
    layer2_outputs(1374) <= (layer1_outputs(6994)) and not (layer1_outputs(6720));
    layer2_outputs(1375) <= (layer1_outputs(5296)) and not (layer1_outputs(5895));
    layer2_outputs(1376) <= not((layer1_outputs(4512)) or (layer1_outputs(1979)));
    layer2_outputs(1377) <= (layer1_outputs(3050)) and not (layer1_outputs(871));
    layer2_outputs(1378) <= (layer1_outputs(3673)) and not (layer1_outputs(6622));
    layer2_outputs(1379) <= not(layer1_outputs(7633));
    layer2_outputs(1380) <= not(layer1_outputs(1764));
    layer2_outputs(1381) <= layer1_outputs(6317);
    layer2_outputs(1382) <= layer1_outputs(4020);
    layer2_outputs(1383) <= (layer1_outputs(3579)) or (layer1_outputs(1317));
    layer2_outputs(1384) <= (layer1_outputs(2870)) and not (layer1_outputs(5573));
    layer2_outputs(1385) <= not((layer1_outputs(318)) or (layer1_outputs(7372)));
    layer2_outputs(1386) <= layer1_outputs(3294);
    layer2_outputs(1387) <= not((layer1_outputs(2139)) or (layer1_outputs(6757)));
    layer2_outputs(1388) <= not(layer1_outputs(4032)) or (layer1_outputs(3770));
    layer2_outputs(1389) <= not(layer1_outputs(6613));
    layer2_outputs(1390) <= (layer1_outputs(1194)) and not (layer1_outputs(519));
    layer2_outputs(1391) <= layer1_outputs(5575);
    layer2_outputs(1392) <= layer1_outputs(6972);
    layer2_outputs(1393) <= '1';
    layer2_outputs(1394) <= not((layer1_outputs(4199)) xor (layer1_outputs(882)));
    layer2_outputs(1395) <= not(layer1_outputs(6896)) or (layer1_outputs(3701));
    layer2_outputs(1396) <= layer1_outputs(5161);
    layer2_outputs(1397) <= (layer1_outputs(576)) xor (layer1_outputs(1117));
    layer2_outputs(1398) <= layer1_outputs(20);
    layer2_outputs(1399) <= '0';
    layer2_outputs(1400) <= (layer1_outputs(6483)) and not (layer1_outputs(2542));
    layer2_outputs(1401) <= '0';
    layer2_outputs(1402) <= layer1_outputs(4846);
    layer2_outputs(1403) <= not((layer1_outputs(4856)) or (layer1_outputs(5328)));
    layer2_outputs(1404) <= not(layer1_outputs(2357));
    layer2_outputs(1405) <= (layer1_outputs(5385)) and (layer1_outputs(7668));
    layer2_outputs(1406) <= not(layer1_outputs(3453)) or (layer1_outputs(996));
    layer2_outputs(1407) <= (layer1_outputs(1998)) and not (layer1_outputs(1768));
    layer2_outputs(1408) <= not(layer1_outputs(4213));
    layer2_outputs(1409) <= not(layer1_outputs(7263)) or (layer1_outputs(1739));
    layer2_outputs(1410) <= '1';
    layer2_outputs(1411) <= not((layer1_outputs(5200)) and (layer1_outputs(944)));
    layer2_outputs(1412) <= (layer1_outputs(1932)) and not (layer1_outputs(1769));
    layer2_outputs(1413) <= not(layer1_outputs(319));
    layer2_outputs(1414) <= '0';
    layer2_outputs(1415) <= (layer1_outputs(2717)) or (layer1_outputs(6133));
    layer2_outputs(1416) <= layer1_outputs(4296);
    layer2_outputs(1417) <= '0';
    layer2_outputs(1418) <= not(layer1_outputs(5258)) or (layer1_outputs(7606));
    layer2_outputs(1419) <= not(layer1_outputs(6586)) or (layer1_outputs(5485));
    layer2_outputs(1420) <= layer1_outputs(4925);
    layer2_outputs(1421) <= (layer1_outputs(3014)) or (layer1_outputs(2327));
    layer2_outputs(1422) <= not(layer1_outputs(1459));
    layer2_outputs(1423) <= (layer1_outputs(6449)) and not (layer1_outputs(1497));
    layer2_outputs(1424) <= (layer1_outputs(3425)) and not (layer1_outputs(627));
    layer2_outputs(1425) <= layer1_outputs(656);
    layer2_outputs(1426) <= (layer1_outputs(955)) or (layer1_outputs(375));
    layer2_outputs(1427) <= not(layer1_outputs(2976));
    layer2_outputs(1428) <= (layer1_outputs(2352)) or (layer1_outputs(7075));
    layer2_outputs(1429) <= '0';
    layer2_outputs(1430) <= not(layer1_outputs(7228));
    layer2_outputs(1431) <= not(layer1_outputs(2897)) or (layer1_outputs(5261));
    layer2_outputs(1432) <= layer1_outputs(6472);
    layer2_outputs(1433) <= (layer1_outputs(3385)) and (layer1_outputs(4553));
    layer2_outputs(1434) <= (layer1_outputs(4240)) xor (layer1_outputs(4670));
    layer2_outputs(1435) <= (layer1_outputs(6303)) or (layer1_outputs(740));
    layer2_outputs(1436) <= not(layer1_outputs(4051));
    layer2_outputs(1437) <= (layer1_outputs(3654)) and not (layer1_outputs(5068));
    layer2_outputs(1438) <= (layer1_outputs(5988)) and (layer1_outputs(4617));
    layer2_outputs(1439) <= not(layer1_outputs(5263));
    layer2_outputs(1440) <= layer1_outputs(4600);
    layer2_outputs(1441) <= not(layer1_outputs(3261)) or (layer1_outputs(904));
    layer2_outputs(1442) <= not(layer1_outputs(4480)) or (layer1_outputs(1609));
    layer2_outputs(1443) <= not((layer1_outputs(3567)) or (layer1_outputs(3213)));
    layer2_outputs(1444) <= (layer1_outputs(3793)) and (layer1_outputs(7351));
    layer2_outputs(1445) <= layer1_outputs(3706);
    layer2_outputs(1446) <= not((layer1_outputs(5660)) or (layer1_outputs(1612)));
    layer2_outputs(1447) <= not(layer1_outputs(535));
    layer2_outputs(1448) <= (layer1_outputs(1862)) xor (layer1_outputs(4734));
    layer2_outputs(1449) <= (layer1_outputs(3687)) and not (layer1_outputs(2055));
    layer2_outputs(1450) <= (layer1_outputs(5456)) and (layer1_outputs(4325));
    layer2_outputs(1451) <= layer1_outputs(4437);
    layer2_outputs(1452) <= not(layer1_outputs(2405)) or (layer1_outputs(4695));
    layer2_outputs(1453) <= not(layer1_outputs(2721)) or (layer1_outputs(3179));
    layer2_outputs(1454) <= layer1_outputs(2517);
    layer2_outputs(1455) <= not(layer1_outputs(3496)) or (layer1_outputs(5332));
    layer2_outputs(1456) <= not((layer1_outputs(1393)) and (layer1_outputs(6313)));
    layer2_outputs(1457) <= (layer1_outputs(457)) and (layer1_outputs(2044));
    layer2_outputs(1458) <= not(layer1_outputs(2678)) or (layer1_outputs(142));
    layer2_outputs(1459) <= (layer1_outputs(6496)) and (layer1_outputs(5617));
    layer2_outputs(1460) <= '0';
    layer2_outputs(1461) <= (layer1_outputs(6105)) xor (layer1_outputs(1878));
    layer2_outputs(1462) <= '0';
    layer2_outputs(1463) <= not(layer1_outputs(5046)) or (layer1_outputs(1994));
    layer2_outputs(1464) <= not(layer1_outputs(6854));
    layer2_outputs(1465) <= layer1_outputs(2708);
    layer2_outputs(1466) <= '0';
    layer2_outputs(1467) <= layer1_outputs(1557);
    layer2_outputs(1468) <= layer1_outputs(5166);
    layer2_outputs(1469) <= not(layer1_outputs(952)) or (layer1_outputs(7572));
    layer2_outputs(1470) <= not(layer1_outputs(4865));
    layer2_outputs(1471) <= layer1_outputs(2447);
    layer2_outputs(1472) <= (layer1_outputs(4210)) xor (layer1_outputs(430));
    layer2_outputs(1473) <= (layer1_outputs(5874)) and (layer1_outputs(4444));
    layer2_outputs(1474) <= not(layer1_outputs(4278)) or (layer1_outputs(427));
    layer2_outputs(1475) <= layer1_outputs(1846);
    layer2_outputs(1476) <= not(layer1_outputs(227)) or (layer1_outputs(4979));
    layer2_outputs(1477) <= (layer1_outputs(443)) and not (layer1_outputs(4369));
    layer2_outputs(1478) <= not(layer1_outputs(4274));
    layer2_outputs(1479) <= (layer1_outputs(2932)) and not (layer1_outputs(1607));
    layer2_outputs(1480) <= layer1_outputs(2659);
    layer2_outputs(1481) <= (layer1_outputs(3022)) and (layer1_outputs(248));
    layer2_outputs(1482) <= not(layer1_outputs(826));
    layer2_outputs(1483) <= layer1_outputs(6767);
    layer2_outputs(1484) <= (layer1_outputs(6202)) or (layer1_outputs(1226));
    layer2_outputs(1485) <= (layer1_outputs(2971)) and (layer1_outputs(1277));
    layer2_outputs(1486) <= layer1_outputs(1889);
    layer2_outputs(1487) <= not(layer1_outputs(7212));
    layer2_outputs(1488) <= (layer1_outputs(6125)) and not (layer1_outputs(7391));
    layer2_outputs(1489) <= not(layer1_outputs(784));
    layer2_outputs(1490) <= '1';
    layer2_outputs(1491) <= layer1_outputs(2268);
    layer2_outputs(1492) <= layer1_outputs(3632);
    layer2_outputs(1493) <= not(layer1_outputs(160)) or (layer1_outputs(2466));
    layer2_outputs(1494) <= layer1_outputs(1747);
    layer2_outputs(1495) <= '0';
    layer2_outputs(1496) <= not(layer1_outputs(4819)) or (layer1_outputs(1141));
    layer2_outputs(1497) <= (layer1_outputs(1547)) and not (layer1_outputs(4275));
    layer2_outputs(1498) <= layer1_outputs(7554);
    layer2_outputs(1499) <= (layer1_outputs(7441)) and not (layer1_outputs(7383));
    layer2_outputs(1500) <= not(layer1_outputs(7627)) or (layer1_outputs(3928));
    layer2_outputs(1501) <= layer1_outputs(1726);
    layer2_outputs(1502) <= not(layer1_outputs(7156)) or (layer1_outputs(6268));
    layer2_outputs(1503) <= (layer1_outputs(4855)) and not (layer1_outputs(6978));
    layer2_outputs(1504) <= layer1_outputs(6000);
    layer2_outputs(1505) <= layer1_outputs(4869);
    layer2_outputs(1506) <= layer1_outputs(2973);
    layer2_outputs(1507) <= layer1_outputs(4743);
    layer2_outputs(1508) <= not((layer1_outputs(358)) xor (layer1_outputs(6657)));
    layer2_outputs(1509) <= layer1_outputs(7217);
    layer2_outputs(1510) <= (layer1_outputs(3773)) and not (layer1_outputs(5275));
    layer2_outputs(1511) <= not((layer1_outputs(4652)) or (layer1_outputs(4735)));
    layer2_outputs(1512) <= layer1_outputs(5510);
    layer2_outputs(1513) <= (layer1_outputs(6736)) and not (layer1_outputs(1741));
    layer2_outputs(1514) <= layer1_outputs(622);
    layer2_outputs(1515) <= (layer1_outputs(584)) or (layer1_outputs(538));
    layer2_outputs(1516) <= layer1_outputs(6481);
    layer2_outputs(1517) <= '1';
    layer2_outputs(1518) <= not((layer1_outputs(4033)) or (layer1_outputs(1576)));
    layer2_outputs(1519) <= layer1_outputs(555);
    layer2_outputs(1520) <= not(layer1_outputs(833)) or (layer1_outputs(5074));
    layer2_outputs(1521) <= not(layer1_outputs(1543));
    layer2_outputs(1522) <= layer1_outputs(2274);
    layer2_outputs(1523) <= layer1_outputs(5239);
    layer2_outputs(1524) <= not(layer1_outputs(717)) or (layer1_outputs(5396));
    layer2_outputs(1525) <= not(layer1_outputs(3699));
    layer2_outputs(1526) <= not((layer1_outputs(471)) and (layer1_outputs(5836)));
    layer2_outputs(1527) <= '0';
    layer2_outputs(1528) <= not((layer1_outputs(3849)) or (layer1_outputs(842)));
    layer2_outputs(1529) <= (layer1_outputs(2166)) and not (layer1_outputs(5308));
    layer2_outputs(1530) <= not(layer1_outputs(1856));
    layer2_outputs(1531) <= not(layer1_outputs(2061)) or (layer1_outputs(4772));
    layer2_outputs(1532) <= layer1_outputs(4700);
    layer2_outputs(1533) <= layer1_outputs(1019);
    layer2_outputs(1534) <= not((layer1_outputs(4714)) or (layer1_outputs(6016)));
    layer2_outputs(1535) <= not(layer1_outputs(3347)) or (layer1_outputs(7546));
    layer2_outputs(1536) <= not(layer1_outputs(228));
    layer2_outputs(1537) <= not(layer1_outputs(60)) or (layer1_outputs(2036));
    layer2_outputs(1538) <= not((layer1_outputs(2391)) and (layer1_outputs(6881)));
    layer2_outputs(1539) <= layer1_outputs(3481);
    layer2_outputs(1540) <= layer1_outputs(4858);
    layer2_outputs(1541) <= layer1_outputs(3519);
    layer2_outputs(1542) <= not(layer1_outputs(116)) or (layer1_outputs(7607));
    layer2_outputs(1543) <= (layer1_outputs(5537)) and (layer1_outputs(4837));
    layer2_outputs(1544) <= not(layer1_outputs(3818));
    layer2_outputs(1545) <= not(layer1_outputs(7182));
    layer2_outputs(1546) <= (layer1_outputs(4981)) and not (layer1_outputs(2175));
    layer2_outputs(1547) <= not(layer1_outputs(3735));
    layer2_outputs(1548) <= '0';
    layer2_outputs(1549) <= not(layer1_outputs(3464));
    layer2_outputs(1550) <= not(layer1_outputs(7261)) or (layer1_outputs(1926));
    layer2_outputs(1551) <= not(layer1_outputs(4912));
    layer2_outputs(1552) <= layer1_outputs(4345);
    layer2_outputs(1553) <= layer1_outputs(6718);
    layer2_outputs(1554) <= (layer1_outputs(4766)) or (layer1_outputs(2832));
    layer2_outputs(1555) <= not(layer1_outputs(4842));
    layer2_outputs(1556) <= not(layer1_outputs(5158));
    layer2_outputs(1557) <= not(layer1_outputs(5300)) or (layer1_outputs(6375));
    layer2_outputs(1558) <= not(layer1_outputs(4994));
    layer2_outputs(1559) <= layer1_outputs(3695);
    layer2_outputs(1560) <= '0';
    layer2_outputs(1561) <= '0';
    layer2_outputs(1562) <= not(layer1_outputs(3718));
    layer2_outputs(1563) <= not((layer1_outputs(6422)) xor (layer1_outputs(2401)));
    layer2_outputs(1564) <= (layer1_outputs(5965)) or (layer1_outputs(4057));
    layer2_outputs(1565) <= not(layer1_outputs(855));
    layer2_outputs(1566) <= not(layer1_outputs(1777));
    layer2_outputs(1567) <= not(layer1_outputs(6551));
    layer2_outputs(1568) <= not(layer1_outputs(5859));
    layer2_outputs(1569) <= layer1_outputs(7302);
    layer2_outputs(1570) <= not((layer1_outputs(347)) or (layer1_outputs(4039)));
    layer2_outputs(1571) <= not(layer1_outputs(688));
    layer2_outputs(1572) <= layer1_outputs(3596);
    layer2_outputs(1573) <= not((layer1_outputs(5687)) and (layer1_outputs(6466)));
    layer2_outputs(1574) <= not(layer1_outputs(7153));
    layer2_outputs(1575) <= layer1_outputs(5659);
    layer2_outputs(1576) <= not(layer1_outputs(5347));
    layer2_outputs(1577) <= (layer1_outputs(2437)) and not (layer1_outputs(2978));
    layer2_outputs(1578) <= not(layer1_outputs(5782)) or (layer1_outputs(1732));
    layer2_outputs(1579) <= layer1_outputs(6385);
    layer2_outputs(1580) <= (layer1_outputs(5834)) or (layer1_outputs(7405));
    layer2_outputs(1581) <= layer1_outputs(404);
    layer2_outputs(1582) <= '1';
    layer2_outputs(1583) <= not(layer1_outputs(3418)) or (layer1_outputs(4190));
    layer2_outputs(1584) <= (layer1_outputs(5143)) and (layer1_outputs(599));
    layer2_outputs(1585) <= (layer1_outputs(3559)) or (layer1_outputs(832));
    layer2_outputs(1586) <= layer1_outputs(7559);
    layer2_outputs(1587) <= not(layer1_outputs(3733));
    layer2_outputs(1588) <= not((layer1_outputs(1477)) and (layer1_outputs(5727)));
    layer2_outputs(1589) <= '0';
    layer2_outputs(1590) <= (layer1_outputs(1703)) and not (layer1_outputs(7416));
    layer2_outputs(1591) <= (layer1_outputs(3223)) and not (layer1_outputs(2947));
    layer2_outputs(1592) <= not(layer1_outputs(34)) or (layer1_outputs(1620));
    layer2_outputs(1593) <= not(layer1_outputs(1571));
    layer2_outputs(1594) <= not(layer1_outputs(3625)) or (layer1_outputs(1303));
    layer2_outputs(1595) <= layer1_outputs(1261);
    layer2_outputs(1596) <= (layer1_outputs(736)) or (layer1_outputs(2042));
    layer2_outputs(1597) <= not(layer1_outputs(4042));
    layer2_outputs(1598) <= not(layer1_outputs(115)) or (layer1_outputs(6507));
    layer2_outputs(1599) <= layer1_outputs(2776);
    layer2_outputs(1600) <= not(layer1_outputs(2159)) or (layer1_outputs(3185));
    layer2_outputs(1601) <= not((layer1_outputs(2295)) and (layer1_outputs(2577)));
    layer2_outputs(1602) <= (layer1_outputs(4798)) or (layer1_outputs(3325));
    layer2_outputs(1603) <= not(layer1_outputs(7478));
    layer2_outputs(1604) <= layer1_outputs(755);
    layer2_outputs(1605) <= layer1_outputs(2924);
    layer2_outputs(1606) <= not(layer1_outputs(5318));
    layer2_outputs(1607) <= not(layer1_outputs(6871));
    layer2_outputs(1608) <= not(layer1_outputs(390));
    layer2_outputs(1609) <= '1';
    layer2_outputs(1610) <= not((layer1_outputs(3649)) or (layer1_outputs(3903)));
    layer2_outputs(1611) <= not(layer1_outputs(2974));
    layer2_outputs(1612) <= not((layer1_outputs(1723)) or (layer1_outputs(376)));
    layer2_outputs(1613) <= layer1_outputs(3441);
    layer2_outputs(1614) <= not(layer1_outputs(2476));
    layer2_outputs(1615) <= (layer1_outputs(3103)) and (layer1_outputs(647));
    layer2_outputs(1616) <= not((layer1_outputs(6601)) or (layer1_outputs(6639)));
    layer2_outputs(1617) <= (layer1_outputs(6052)) and (layer1_outputs(65));
    layer2_outputs(1618) <= not(layer1_outputs(7657));
    layer2_outputs(1619) <= not(layer1_outputs(4726));
    layer2_outputs(1620) <= not((layer1_outputs(3718)) or (layer1_outputs(771)));
    layer2_outputs(1621) <= not(layer1_outputs(885));
    layer2_outputs(1622) <= not(layer1_outputs(7054));
    layer2_outputs(1623) <= (layer1_outputs(1595)) and not (layer1_outputs(2426));
    layer2_outputs(1624) <= layer1_outputs(3076);
    layer2_outputs(1625) <= not(layer1_outputs(168));
    layer2_outputs(1626) <= not((layer1_outputs(298)) and (layer1_outputs(2040)));
    layer2_outputs(1627) <= not(layer1_outputs(4537)) or (layer1_outputs(2238));
    layer2_outputs(1628) <= not(layer1_outputs(4801));
    layer2_outputs(1629) <= layer1_outputs(3147);
    layer2_outputs(1630) <= (layer1_outputs(2657)) and not (layer1_outputs(6456));
    layer2_outputs(1631) <= not((layer1_outputs(4173)) or (layer1_outputs(7208)));
    layer2_outputs(1632) <= (layer1_outputs(4751)) and (layer1_outputs(6017));
    layer2_outputs(1633) <= (layer1_outputs(5413)) and not (layer1_outputs(1762));
    layer2_outputs(1634) <= not((layer1_outputs(2217)) or (layer1_outputs(5894)));
    layer2_outputs(1635) <= not((layer1_outputs(5199)) and (layer1_outputs(1554)));
    layer2_outputs(1636) <= not((layer1_outputs(1315)) or (layer1_outputs(3932)));
    layer2_outputs(1637) <= '1';
    layer2_outputs(1638) <= not(layer1_outputs(6741));
    layer2_outputs(1639) <= (layer1_outputs(1731)) and not (layer1_outputs(6022));
    layer2_outputs(1640) <= not((layer1_outputs(2713)) or (layer1_outputs(5334)));
    layer2_outputs(1641) <= not(layer1_outputs(2308)) or (layer1_outputs(5916));
    layer2_outputs(1642) <= (layer1_outputs(28)) and not (layer1_outputs(3376));
    layer2_outputs(1643) <= not(layer1_outputs(6300)) or (layer1_outputs(5271));
    layer2_outputs(1644) <= layer1_outputs(5319);
    layer2_outputs(1645) <= (layer1_outputs(4294)) xor (layer1_outputs(6063));
    layer2_outputs(1646) <= layer1_outputs(732);
    layer2_outputs(1647) <= layer1_outputs(3644);
    layer2_outputs(1648) <= (layer1_outputs(3163)) and not (layer1_outputs(3227));
    layer2_outputs(1649) <= layer1_outputs(388);
    layer2_outputs(1650) <= (layer1_outputs(4430)) xor (layer1_outputs(76));
    layer2_outputs(1651) <= layer1_outputs(4501);
    layer2_outputs(1652) <= not(layer1_outputs(6082)) or (layer1_outputs(3720));
    layer2_outputs(1653) <= not(layer1_outputs(4026));
    layer2_outputs(1654) <= not(layer1_outputs(4736));
    layer2_outputs(1655) <= not((layer1_outputs(2690)) or (layer1_outputs(851)));
    layer2_outputs(1656) <= not(layer1_outputs(1965));
    layer2_outputs(1657) <= not(layer1_outputs(4402));
    layer2_outputs(1658) <= '1';
    layer2_outputs(1659) <= (layer1_outputs(2672)) and not (layer1_outputs(3275));
    layer2_outputs(1660) <= '1';
    layer2_outputs(1661) <= layer1_outputs(2748);
    layer2_outputs(1662) <= layer1_outputs(6841);
    layer2_outputs(1663) <= not((layer1_outputs(3748)) and (layer1_outputs(7012)));
    layer2_outputs(1664) <= layer1_outputs(6624);
    layer2_outputs(1665) <= layer1_outputs(486);
    layer2_outputs(1666) <= layer1_outputs(7134);
    layer2_outputs(1667) <= layer1_outputs(5884);
    layer2_outputs(1668) <= not(layer1_outputs(3805));
    layer2_outputs(1669) <= layer1_outputs(2946);
    layer2_outputs(1670) <= layer1_outputs(2465);
    layer2_outputs(1671) <= (layer1_outputs(4191)) and (layer1_outputs(2521));
    layer2_outputs(1672) <= (layer1_outputs(1537)) and not (layer1_outputs(6380));
    layer2_outputs(1673) <= layer1_outputs(5329);
    layer2_outputs(1674) <= not(layer1_outputs(6734));
    layer2_outputs(1675) <= (layer1_outputs(2823)) and (layer1_outputs(2636));
    layer2_outputs(1676) <= '0';
    layer2_outputs(1677) <= (layer1_outputs(4867)) or (layer1_outputs(6762));
    layer2_outputs(1678) <= (layer1_outputs(6154)) or (layer1_outputs(3595));
    layer2_outputs(1679) <= not(layer1_outputs(3288)) or (layer1_outputs(5919));
    layer2_outputs(1680) <= not((layer1_outputs(4124)) or (layer1_outputs(5776)));
    layer2_outputs(1681) <= not((layer1_outputs(1635)) and (layer1_outputs(1907)));
    layer2_outputs(1682) <= layer1_outputs(5029);
    layer2_outputs(1683) <= not(layer1_outputs(3496));
    layer2_outputs(1684) <= '0';
    layer2_outputs(1685) <= not(layer1_outputs(7561)) or (layer1_outputs(143));
    layer2_outputs(1686) <= layer1_outputs(1619);
    layer2_outputs(1687) <= (layer1_outputs(4290)) and not (layer1_outputs(7090));
    layer2_outputs(1688) <= (layer1_outputs(5951)) and (layer1_outputs(626));
    layer2_outputs(1689) <= not(layer1_outputs(3585)) or (layer1_outputs(1345));
    layer2_outputs(1690) <= layer1_outputs(7228);
    layer2_outputs(1691) <= layer1_outputs(3594);
    layer2_outputs(1692) <= layer1_outputs(7438);
    layer2_outputs(1693) <= not((layer1_outputs(1265)) or (layer1_outputs(7577)));
    layer2_outputs(1694) <= not(layer1_outputs(3196)) or (layer1_outputs(6967));
    layer2_outputs(1695) <= not((layer1_outputs(6231)) and (layer1_outputs(858)));
    layer2_outputs(1696) <= not(layer1_outputs(3588)) or (layer1_outputs(359));
    layer2_outputs(1697) <= (layer1_outputs(4090)) or (layer1_outputs(5872));
    layer2_outputs(1698) <= (layer1_outputs(2103)) and not (layer1_outputs(7400));
    layer2_outputs(1699) <= (layer1_outputs(2561)) and not (layer1_outputs(7584));
    layer2_outputs(1700) <= layer1_outputs(5748);
    layer2_outputs(1701) <= not(layer1_outputs(7057)) or (layer1_outputs(6633));
    layer2_outputs(1702) <= layer1_outputs(4421);
    layer2_outputs(1703) <= not(layer1_outputs(2072));
    layer2_outputs(1704) <= layer1_outputs(224);
    layer2_outputs(1705) <= layer1_outputs(7321);
    layer2_outputs(1706) <= not(layer1_outputs(5985));
    layer2_outputs(1707) <= '1';
    layer2_outputs(1708) <= (layer1_outputs(7476)) and (layer1_outputs(1879));
    layer2_outputs(1709) <= layer1_outputs(4694);
    layer2_outputs(1710) <= not(layer1_outputs(896));
    layer2_outputs(1711) <= not((layer1_outputs(5594)) and (layer1_outputs(1903)));
    layer2_outputs(1712) <= layer1_outputs(196);
    layer2_outputs(1713) <= not(layer1_outputs(2732)) or (layer1_outputs(7000));
    layer2_outputs(1714) <= not((layer1_outputs(5618)) and (layer1_outputs(4648)));
    layer2_outputs(1715) <= layer1_outputs(3453);
    layer2_outputs(1716) <= layer1_outputs(4599);
    layer2_outputs(1717) <= not(layer1_outputs(2443)) or (layer1_outputs(4671));
    layer2_outputs(1718) <= not((layer1_outputs(6071)) and (layer1_outputs(5163)));
    layer2_outputs(1719) <= not(layer1_outputs(2165));
    layer2_outputs(1720) <= (layer1_outputs(3922)) xor (layer1_outputs(4384));
    layer2_outputs(1721) <= (layer1_outputs(7107)) and (layer1_outputs(1902));
    layer2_outputs(1722) <= (layer1_outputs(7166)) and not (layer1_outputs(3195));
    layer2_outputs(1723) <= layer1_outputs(2947);
    layer2_outputs(1724) <= layer1_outputs(2355);
    layer2_outputs(1725) <= not(layer1_outputs(1685)) or (layer1_outputs(3617));
    layer2_outputs(1726) <= '1';
    layer2_outputs(1727) <= (layer1_outputs(1752)) and (layer1_outputs(1823));
    layer2_outputs(1728) <= not(layer1_outputs(621));
    layer2_outputs(1729) <= not(layer1_outputs(6429));
    layer2_outputs(1730) <= (layer1_outputs(2287)) and (layer1_outputs(7305));
    layer2_outputs(1731) <= (layer1_outputs(5140)) and (layer1_outputs(248));
    layer2_outputs(1732) <= (layer1_outputs(1929)) and not (layer1_outputs(3856));
    layer2_outputs(1733) <= not(layer1_outputs(5412));
    layer2_outputs(1734) <= not(layer1_outputs(1698)) or (layer1_outputs(6339));
    layer2_outputs(1735) <= (layer1_outputs(6355)) or (layer1_outputs(243));
    layer2_outputs(1736) <= layer1_outputs(1034);
    layer2_outputs(1737) <= not((layer1_outputs(1122)) xor (layer1_outputs(109)));
    layer2_outputs(1738) <= layer1_outputs(2698);
    layer2_outputs(1739) <= (layer1_outputs(928)) or (layer1_outputs(5467));
    layer2_outputs(1740) <= (layer1_outputs(3460)) and (layer1_outputs(6015));
    layer2_outputs(1741) <= (layer1_outputs(4596)) and not (layer1_outputs(3620));
    layer2_outputs(1742) <= not((layer1_outputs(94)) and (layer1_outputs(1831)));
    layer2_outputs(1743) <= not(layer1_outputs(5156)) or (layer1_outputs(4350));
    layer2_outputs(1744) <= layer1_outputs(1403);
    layer2_outputs(1745) <= layer1_outputs(2899);
    layer2_outputs(1746) <= layer1_outputs(5245);
    layer2_outputs(1747) <= (layer1_outputs(1973)) and not (layer1_outputs(3513));
    layer2_outputs(1748) <= '1';
    layer2_outputs(1749) <= not(layer1_outputs(1219));
    layer2_outputs(1750) <= not((layer1_outputs(2839)) xor (layer1_outputs(812)));
    layer2_outputs(1751) <= layer1_outputs(5401);
    layer2_outputs(1752) <= layer1_outputs(1730);
    layer2_outputs(1753) <= (layer1_outputs(5730)) and not (layer1_outputs(2413));
    layer2_outputs(1754) <= not(layer1_outputs(2525));
    layer2_outputs(1755) <= layer1_outputs(6325);
    layer2_outputs(1756) <= '0';
    layer2_outputs(1757) <= layer1_outputs(4009);
    layer2_outputs(1758) <= (layer1_outputs(935)) and not (layer1_outputs(466));
    layer2_outputs(1759) <= not(layer1_outputs(1316)) or (layer1_outputs(5427));
    layer2_outputs(1760) <= layer1_outputs(3946);
    layer2_outputs(1761) <= '1';
    layer2_outputs(1762) <= layer1_outputs(3800);
    layer2_outputs(1763) <= not(layer1_outputs(1432));
    layer2_outputs(1764) <= layer1_outputs(6383);
    layer2_outputs(1765) <= (layer1_outputs(1036)) and (layer1_outputs(3602));
    layer2_outputs(1766) <= not(layer1_outputs(525));
    layer2_outputs(1767) <= (layer1_outputs(1454)) or (layer1_outputs(2288));
    layer2_outputs(1768) <= (layer1_outputs(591)) and not (layer1_outputs(1429));
    layer2_outputs(1769) <= (layer1_outputs(2022)) or (layer1_outputs(7207));
    layer2_outputs(1770) <= (layer1_outputs(3374)) and not (layer1_outputs(3972));
    layer2_outputs(1771) <= not(layer1_outputs(7614));
    layer2_outputs(1772) <= layer1_outputs(7510);
    layer2_outputs(1773) <= not(layer1_outputs(268)) or (layer1_outputs(3467));
    layer2_outputs(1774) <= '1';
    layer2_outputs(1775) <= not(layer1_outputs(3982)) or (layer1_outputs(5545));
    layer2_outputs(1776) <= '1';
    layer2_outputs(1777) <= not((layer1_outputs(1546)) or (layer1_outputs(1910)));
    layer2_outputs(1778) <= '0';
    layer2_outputs(1779) <= (layer1_outputs(4334)) and not (layer1_outputs(467));
    layer2_outputs(1780) <= not(layer1_outputs(1641)) or (layer1_outputs(6306));
    layer2_outputs(1781) <= not((layer1_outputs(5454)) and (layer1_outputs(2941)));
    layer2_outputs(1782) <= not(layer1_outputs(5975));
    layer2_outputs(1783) <= (layer1_outputs(4438)) xor (layer1_outputs(6796));
    layer2_outputs(1784) <= layer1_outputs(5633);
    layer2_outputs(1785) <= not(layer1_outputs(2573)) or (layer1_outputs(6495));
    layer2_outputs(1786) <= layer1_outputs(5034);
    layer2_outputs(1787) <= (layer1_outputs(604)) or (layer1_outputs(7153));
    layer2_outputs(1788) <= not(layer1_outputs(6681));
    layer2_outputs(1789) <= (layer1_outputs(5848)) and (layer1_outputs(7666));
    layer2_outputs(1790) <= (layer1_outputs(1746)) and not (layer1_outputs(6751));
    layer2_outputs(1791) <= layer1_outputs(336);
    layer2_outputs(1792) <= (layer1_outputs(1003)) and (layer1_outputs(304));
    layer2_outputs(1793) <= not(layer1_outputs(6110));
    layer2_outputs(1794) <= not(layer1_outputs(3738)) or (layer1_outputs(7173));
    layer2_outputs(1795) <= not(layer1_outputs(1959));
    layer2_outputs(1796) <= '1';
    layer2_outputs(1797) <= not((layer1_outputs(3346)) and (layer1_outputs(5275)));
    layer2_outputs(1798) <= (layer1_outputs(4035)) and (layer1_outputs(3960));
    layer2_outputs(1799) <= not((layer1_outputs(939)) and (layer1_outputs(6090)));
    layer2_outputs(1800) <= layer1_outputs(3246);
    layer2_outputs(1801) <= not((layer1_outputs(1653)) and (layer1_outputs(5408)));
    layer2_outputs(1802) <= not(layer1_outputs(813));
    layer2_outputs(1803) <= not(layer1_outputs(3927));
    layer2_outputs(1804) <= not(layer1_outputs(485));
    layer2_outputs(1805) <= (layer1_outputs(6900)) or (layer1_outputs(3662));
    layer2_outputs(1806) <= '1';
    layer2_outputs(1807) <= '1';
    layer2_outputs(1808) <= not(layer1_outputs(2048));
    layer2_outputs(1809) <= (layer1_outputs(1397)) xor (layer1_outputs(1503));
    layer2_outputs(1810) <= layer1_outputs(327);
    layer2_outputs(1811) <= not(layer1_outputs(6230));
    layer2_outputs(1812) <= (layer1_outputs(4744)) or (layer1_outputs(3877));
    layer2_outputs(1813) <= (layer1_outputs(3041)) and not (layer1_outputs(5805));
    layer2_outputs(1814) <= layer1_outputs(1524);
    layer2_outputs(1815) <= not(layer1_outputs(189)) or (layer1_outputs(2255));
    layer2_outputs(1816) <= layer1_outputs(6544);
    layer2_outputs(1817) <= not((layer1_outputs(482)) or (layer1_outputs(1462)));
    layer2_outputs(1818) <= layer1_outputs(5613);
    layer2_outputs(1819) <= not((layer1_outputs(4761)) xor (layer1_outputs(2837)));
    layer2_outputs(1820) <= layer1_outputs(5552);
    layer2_outputs(1821) <= not(layer1_outputs(2249));
    layer2_outputs(1822) <= (layer1_outputs(325)) and not (layer1_outputs(6825));
    layer2_outputs(1823) <= not(layer1_outputs(2132));
    layer2_outputs(1824) <= (layer1_outputs(5754)) or (layer1_outputs(1746));
    layer2_outputs(1825) <= not((layer1_outputs(7224)) and (layer1_outputs(603)));
    layer2_outputs(1826) <= layer1_outputs(3824);
    layer2_outputs(1827) <= not((layer1_outputs(7581)) or (layer1_outputs(5777)));
    layer2_outputs(1828) <= not((layer1_outputs(3067)) or (layer1_outputs(262)));
    layer2_outputs(1829) <= (layer1_outputs(5900)) xor (layer1_outputs(2347));
    layer2_outputs(1830) <= not(layer1_outputs(2311));
    layer2_outputs(1831) <= (layer1_outputs(586)) and (layer1_outputs(3930));
    layer2_outputs(1832) <= (layer1_outputs(632)) xor (layer1_outputs(5373));
    layer2_outputs(1833) <= layer1_outputs(4801);
    layer2_outputs(1834) <= layer1_outputs(4636);
    layer2_outputs(1835) <= layer1_outputs(3020);
    layer2_outputs(1836) <= not(layer1_outputs(2038));
    layer2_outputs(1837) <= layer1_outputs(640);
    layer2_outputs(1838) <= not(layer1_outputs(4003));
    layer2_outputs(1839) <= (layer1_outputs(4885)) and not (layer1_outputs(1490));
    layer2_outputs(1840) <= not((layer1_outputs(2472)) xor (layer1_outputs(7231)));
    layer2_outputs(1841) <= (layer1_outputs(3468)) and (layer1_outputs(4243));
    layer2_outputs(1842) <= layer1_outputs(1935);
    layer2_outputs(1843) <= not((layer1_outputs(1949)) or (layer1_outputs(2237)));
    layer2_outputs(1844) <= not(layer1_outputs(7528));
    layer2_outputs(1845) <= not((layer1_outputs(1078)) or (layer1_outputs(5980)));
    layer2_outputs(1846) <= layer1_outputs(889);
    layer2_outputs(1847) <= not((layer1_outputs(2069)) and (layer1_outputs(4603)));
    layer2_outputs(1848) <= not(layer1_outputs(4685));
    layer2_outputs(1849) <= layer1_outputs(6213);
    layer2_outputs(1850) <= layer1_outputs(4651);
    layer2_outputs(1851) <= not(layer1_outputs(6206)) or (layer1_outputs(3923));
    layer2_outputs(1852) <= (layer1_outputs(5303)) xor (layer1_outputs(6445));
    layer2_outputs(1853) <= not((layer1_outputs(2533)) xor (layer1_outputs(379)));
    layer2_outputs(1854) <= (layer1_outputs(4005)) and not (layer1_outputs(5677));
    layer2_outputs(1855) <= (layer1_outputs(1945)) and (layer1_outputs(5442));
    layer2_outputs(1856) <= not(layer1_outputs(4043));
    layer2_outputs(1857) <= (layer1_outputs(677)) xor (layer1_outputs(51));
    layer2_outputs(1858) <= not(layer1_outputs(2705));
    layer2_outputs(1859) <= '0';
    layer2_outputs(1860) <= layer1_outputs(286);
    layer2_outputs(1861) <= (layer1_outputs(3767)) and not (layer1_outputs(1668));
    layer2_outputs(1862) <= '1';
    layer2_outputs(1863) <= not(layer1_outputs(5508)) or (layer1_outputs(4044));
    layer2_outputs(1864) <= not(layer1_outputs(3777)) or (layer1_outputs(6309));
    layer2_outputs(1865) <= layer1_outputs(1194);
    layer2_outputs(1866) <= layer1_outputs(492);
    layer2_outputs(1867) <= not(layer1_outputs(3149)) or (layer1_outputs(6096));
    layer2_outputs(1868) <= layer1_outputs(1482);
    layer2_outputs(1869) <= not(layer1_outputs(3205));
    layer2_outputs(1870) <= (layer1_outputs(4408)) and not (layer1_outputs(6396));
    layer2_outputs(1871) <= not(layer1_outputs(5631));
    layer2_outputs(1872) <= (layer1_outputs(3230)) or (layer1_outputs(2752));
    layer2_outputs(1873) <= not(layer1_outputs(2538));
    layer2_outputs(1874) <= layer1_outputs(3909);
    layer2_outputs(1875) <= layer1_outputs(6759);
    layer2_outputs(1876) <= (layer1_outputs(654)) and (layer1_outputs(6801));
    layer2_outputs(1877) <= layer1_outputs(5550);
    layer2_outputs(1878) <= layer1_outputs(2397);
    layer2_outputs(1879) <= not(layer1_outputs(4010));
    layer2_outputs(1880) <= (layer1_outputs(6830)) or (layer1_outputs(4103));
    layer2_outputs(1881) <= (layer1_outputs(4580)) and not (layer1_outputs(388));
    layer2_outputs(1882) <= layer1_outputs(1521);
    layer2_outputs(1883) <= layer1_outputs(2222);
    layer2_outputs(1884) <= not(layer1_outputs(1940));
    layer2_outputs(1885) <= '1';
    layer2_outputs(1886) <= (layer1_outputs(2537)) and not (layer1_outputs(4125));
    layer2_outputs(1887) <= not(layer1_outputs(6599));
    layer2_outputs(1888) <= not(layer1_outputs(3488)) or (layer1_outputs(2584));
    layer2_outputs(1889) <= not(layer1_outputs(527));
    layer2_outputs(1890) <= '0';
    layer2_outputs(1891) <= not(layer1_outputs(4548));
    layer2_outputs(1892) <= '1';
    layer2_outputs(1893) <= layer1_outputs(3743);
    layer2_outputs(1894) <= (layer1_outputs(7353)) or (layer1_outputs(4301));
    layer2_outputs(1895) <= not(layer1_outputs(1964));
    layer2_outputs(1896) <= layer1_outputs(2155);
    layer2_outputs(1897) <= layer1_outputs(1375);
    layer2_outputs(1898) <= layer1_outputs(5319);
    layer2_outputs(1899) <= not(layer1_outputs(3021));
    layer2_outputs(1900) <= not((layer1_outputs(2739)) and (layer1_outputs(984)));
    layer2_outputs(1901) <= (layer1_outputs(6749)) or (layer1_outputs(3008));
    layer2_outputs(1902) <= not(layer1_outputs(455)) or (layer1_outputs(5542));
    layer2_outputs(1903) <= (layer1_outputs(6036)) and not (layer1_outputs(5863));
    layer2_outputs(1904) <= (layer1_outputs(1389)) xor (layer1_outputs(2182));
    layer2_outputs(1905) <= layer1_outputs(5224);
    layer2_outputs(1906) <= not((layer1_outputs(4925)) and (layer1_outputs(1149)));
    layer2_outputs(1907) <= (layer1_outputs(5990)) and (layer1_outputs(1839));
    layer2_outputs(1908) <= not(layer1_outputs(823));
    layer2_outputs(1909) <= not((layer1_outputs(2912)) and (layer1_outputs(117)));
    layer2_outputs(1910) <= not(layer1_outputs(2241));
    layer2_outputs(1911) <= layer1_outputs(854);
    layer2_outputs(1912) <= layer1_outputs(5779);
    layer2_outputs(1913) <= not((layer1_outputs(2962)) or (layer1_outputs(5549)));
    layer2_outputs(1914) <= layer1_outputs(824);
    layer2_outputs(1915) <= '0';
    layer2_outputs(1916) <= (layer1_outputs(2285)) and (layer1_outputs(67));
    layer2_outputs(1917) <= not(layer1_outputs(4771));
    layer2_outputs(1918) <= '1';
    layer2_outputs(1919) <= not(layer1_outputs(4297));
    layer2_outputs(1920) <= layer1_outputs(5701);
    layer2_outputs(1921) <= (layer1_outputs(830)) or (layer1_outputs(2742));
    layer2_outputs(1922) <= '1';
    layer2_outputs(1923) <= (layer1_outputs(1208)) and (layer1_outputs(1776));
    layer2_outputs(1924) <= (layer1_outputs(5849)) and (layer1_outputs(5746));
    layer2_outputs(1925) <= not(layer1_outputs(2120));
    layer2_outputs(1926) <= not(layer1_outputs(422));
    layer2_outputs(1927) <= (layer1_outputs(3994)) or (layer1_outputs(7069));
    layer2_outputs(1928) <= (layer1_outputs(3263)) and not (layer1_outputs(933));
    layer2_outputs(1929) <= (layer1_outputs(2334)) and not (layer1_outputs(5455));
    layer2_outputs(1930) <= not(layer1_outputs(2645));
    layer2_outputs(1931) <= not(layer1_outputs(5799)) or (layer1_outputs(1760));
    layer2_outputs(1932) <= (layer1_outputs(7493)) and (layer1_outputs(4927));
    layer2_outputs(1933) <= not(layer1_outputs(5314));
    layer2_outputs(1934) <= (layer1_outputs(609)) or (layer1_outputs(1056));
    layer2_outputs(1935) <= not(layer1_outputs(4526));
    layer2_outputs(1936) <= not((layer1_outputs(735)) xor (layer1_outputs(3314)));
    layer2_outputs(1937) <= not(layer1_outputs(3508)) or (layer1_outputs(5883));
    layer2_outputs(1938) <= (layer1_outputs(6068)) and not (layer1_outputs(5852));
    layer2_outputs(1939) <= not(layer1_outputs(3911)) or (layer1_outputs(3961));
    layer2_outputs(1940) <= (layer1_outputs(5280)) or (layer1_outputs(3030));
    layer2_outputs(1941) <= not(layer1_outputs(1744));
    layer2_outputs(1942) <= not(layer1_outputs(4620));
    layer2_outputs(1943) <= '1';
    layer2_outputs(1944) <= not(layer1_outputs(2359)) or (layer1_outputs(6299));
    layer2_outputs(1945) <= layer1_outputs(3706);
    layer2_outputs(1946) <= layer1_outputs(814);
    layer2_outputs(1947) <= not((layer1_outputs(270)) or (layer1_outputs(3170)));
    layer2_outputs(1948) <= (layer1_outputs(5390)) and (layer1_outputs(6826));
    layer2_outputs(1949) <= not(layer1_outputs(6363));
    layer2_outputs(1950) <= (layer1_outputs(4678)) and not (layer1_outputs(5799));
    layer2_outputs(1951) <= not(layer1_outputs(1138));
    layer2_outputs(1952) <= (layer1_outputs(4183)) or (layer1_outputs(5850));
    layer2_outputs(1953) <= (layer1_outputs(7538)) and (layer1_outputs(537));
    layer2_outputs(1954) <= not(layer1_outputs(685));
    layer2_outputs(1955) <= (layer1_outputs(4970)) and not (layer1_outputs(4628));
    layer2_outputs(1956) <= (layer1_outputs(4505)) and not (layer1_outputs(3893));
    layer2_outputs(1957) <= (layer1_outputs(1628)) and not (layer1_outputs(6521));
    layer2_outputs(1958) <= not(layer1_outputs(4590)) or (layer1_outputs(3113));
    layer2_outputs(1959) <= not(layer1_outputs(5698));
    layer2_outputs(1960) <= (layer1_outputs(920)) or (layer1_outputs(5483));
    layer2_outputs(1961) <= not((layer1_outputs(3574)) and (layer1_outputs(5480)));
    layer2_outputs(1962) <= layer1_outputs(4369);
    layer2_outputs(1963) <= not(layer1_outputs(5689)) or (layer1_outputs(7162));
    layer2_outputs(1964) <= layer1_outputs(1373);
    layer2_outputs(1965) <= layer1_outputs(1487);
    layer2_outputs(1966) <= (layer1_outputs(2214)) and (layer1_outputs(2255));
    layer2_outputs(1967) <= layer1_outputs(2400);
    layer2_outputs(1968) <= (layer1_outputs(3586)) and not (layer1_outputs(804));
    layer2_outputs(1969) <= layer1_outputs(2675);
    layer2_outputs(1970) <= not(layer1_outputs(7033)) or (layer1_outputs(5298));
    layer2_outputs(1971) <= not(layer1_outputs(6408));
    layer2_outputs(1972) <= not(layer1_outputs(3736));
    layer2_outputs(1973) <= layer1_outputs(266);
    layer2_outputs(1974) <= '1';
    layer2_outputs(1975) <= layer1_outputs(4778);
    layer2_outputs(1976) <= '0';
    layer2_outputs(1977) <= not((layer1_outputs(6467)) or (layer1_outputs(4708)));
    layer2_outputs(1978) <= not(layer1_outputs(7219)) or (layer1_outputs(1607));
    layer2_outputs(1979) <= (layer1_outputs(3638)) and not (layer1_outputs(4411));
    layer2_outputs(1980) <= not(layer1_outputs(5094));
    layer2_outputs(1981) <= layer1_outputs(3648);
    layer2_outputs(1982) <= layer1_outputs(1911);
    layer2_outputs(1983) <= not(layer1_outputs(3315));
    layer2_outputs(1984) <= not(layer1_outputs(2948));
    layer2_outputs(1985) <= (layer1_outputs(5910)) or (layer1_outputs(5714));
    layer2_outputs(1986) <= layer1_outputs(2012);
    layer2_outputs(1987) <= not(layer1_outputs(1698));
    layer2_outputs(1988) <= layer1_outputs(260);
    layer2_outputs(1989) <= not(layer1_outputs(7094)) or (layer1_outputs(2054));
    layer2_outputs(1990) <= layer1_outputs(1124);
    layer2_outputs(1991) <= (layer1_outputs(1331)) and not (layer1_outputs(1719));
    layer2_outputs(1992) <= layer1_outputs(3040);
    layer2_outputs(1993) <= '0';
    layer2_outputs(1994) <= not(layer1_outputs(5325));
    layer2_outputs(1995) <= not(layer1_outputs(6323));
    layer2_outputs(1996) <= (layer1_outputs(4124)) and not (layer1_outputs(4458));
    layer2_outputs(1997) <= layer1_outputs(4583);
    layer2_outputs(1998) <= layer1_outputs(3671);
    layer2_outputs(1999) <= not((layer1_outputs(6376)) and (layer1_outputs(1257)));
    layer2_outputs(2000) <= not(layer1_outputs(562)) or (layer1_outputs(1960));
    layer2_outputs(2001) <= '0';
    layer2_outputs(2002) <= layer1_outputs(3622);
    layer2_outputs(2003) <= (layer1_outputs(4937)) or (layer1_outputs(1912));
    layer2_outputs(2004) <= not(layer1_outputs(2963));
    layer2_outputs(2005) <= layer1_outputs(4498);
    layer2_outputs(2006) <= not(layer1_outputs(2316));
    layer2_outputs(2007) <= layer1_outputs(3160);
    layer2_outputs(2008) <= (layer1_outputs(5442)) and (layer1_outputs(1713));
    layer2_outputs(2009) <= not(layer1_outputs(7640)) or (layer1_outputs(6861));
    layer2_outputs(2010) <= (layer1_outputs(2240)) xor (layer1_outputs(6087));
    layer2_outputs(2011) <= not(layer1_outputs(3537)) or (layer1_outputs(1478));
    layer2_outputs(2012) <= layer1_outputs(6251);
    layer2_outputs(2013) <= (layer1_outputs(6936)) and not (layer1_outputs(5461));
    layer2_outputs(2014) <= not(layer1_outputs(4613)) or (layer1_outputs(5809));
    layer2_outputs(2015) <= layer1_outputs(442);
    layer2_outputs(2016) <= layer1_outputs(3425);
    layer2_outputs(2017) <= not((layer1_outputs(400)) and (layer1_outputs(6345)));
    layer2_outputs(2018) <= (layer1_outputs(2117)) or (layer1_outputs(7196));
    layer2_outputs(2019) <= layer1_outputs(4325);
    layer2_outputs(2020) <= not(layer1_outputs(72));
    layer2_outputs(2021) <= not(layer1_outputs(6270));
    layer2_outputs(2022) <= layer1_outputs(4029);
    layer2_outputs(2023) <= not((layer1_outputs(6266)) or (layer1_outputs(7271)));
    layer2_outputs(2024) <= layer1_outputs(4233);
    layer2_outputs(2025) <= layer1_outputs(2673);
    layer2_outputs(2026) <= not(layer1_outputs(6342));
    layer2_outputs(2027) <= '1';
    layer2_outputs(2028) <= '1';
    layer2_outputs(2029) <= (layer1_outputs(1573)) xor (layer1_outputs(5214));
    layer2_outputs(2030) <= layer1_outputs(4665);
    layer2_outputs(2031) <= not(layer1_outputs(2920));
    layer2_outputs(2032) <= '0';
    layer2_outputs(2033) <= not(layer1_outputs(1572));
    layer2_outputs(2034) <= '0';
    layer2_outputs(2035) <= '1';
    layer2_outputs(2036) <= '1';
    layer2_outputs(2037) <= layer1_outputs(7631);
    layer2_outputs(2038) <= not(layer1_outputs(2724));
    layer2_outputs(2039) <= (layer1_outputs(6694)) and (layer1_outputs(129));
    layer2_outputs(2040) <= (layer1_outputs(1128)) and not (layer1_outputs(6075));
    layer2_outputs(2041) <= layer1_outputs(5885);
    layer2_outputs(2042) <= (layer1_outputs(5128)) and not (layer1_outputs(5724));
    layer2_outputs(2043) <= (layer1_outputs(2790)) xor (layer1_outputs(6476));
    layer2_outputs(2044) <= layer1_outputs(565);
    layer2_outputs(2045) <= layer1_outputs(6295);
    layer2_outputs(2046) <= not((layer1_outputs(6242)) or (layer1_outputs(182)));
    layer2_outputs(2047) <= not((layer1_outputs(4884)) or (layer1_outputs(6827)));
    layer2_outputs(2048) <= not(layer1_outputs(3536));
    layer2_outputs(2049) <= not(layer1_outputs(3924));
    layer2_outputs(2050) <= not(layer1_outputs(239)) or (layer1_outputs(5234));
    layer2_outputs(2051) <= not(layer1_outputs(6699));
    layer2_outputs(2052) <= not((layer1_outputs(2453)) or (layer1_outputs(5776)));
    layer2_outputs(2053) <= not(layer1_outputs(2408)) or (layer1_outputs(2115));
    layer2_outputs(2054) <= not(layer1_outputs(819));
    layer2_outputs(2055) <= (layer1_outputs(1683)) xor (layer1_outputs(5328));
    layer2_outputs(2056) <= not((layer1_outputs(7256)) xor (layer1_outputs(163)));
    layer2_outputs(2057) <= (layer1_outputs(6582)) and (layer1_outputs(6444));
    layer2_outputs(2058) <= not(layer1_outputs(3345)) or (layer1_outputs(3765));
    layer2_outputs(2059) <= not((layer1_outputs(6364)) xor (layer1_outputs(2741)));
    layer2_outputs(2060) <= layer1_outputs(3379);
    layer2_outputs(2061) <= not(layer1_outputs(1643)) or (layer1_outputs(3919));
    layer2_outputs(2062) <= not((layer1_outputs(2415)) and (layer1_outputs(3367)));
    layer2_outputs(2063) <= (layer1_outputs(7423)) xor (layer1_outputs(5854));
    layer2_outputs(2064) <= not((layer1_outputs(349)) xor (layer1_outputs(417)));
    layer2_outputs(2065) <= layer1_outputs(4471);
    layer2_outputs(2066) <= layer1_outputs(6065);
    layer2_outputs(2067) <= (layer1_outputs(3442)) and not (layer1_outputs(4680));
    layer2_outputs(2068) <= (layer1_outputs(7454)) and (layer1_outputs(4119));
    layer2_outputs(2069) <= (layer1_outputs(6933)) and (layer1_outputs(4211));
    layer2_outputs(2070) <= (layer1_outputs(6477)) or (layer1_outputs(5518));
    layer2_outputs(2071) <= (layer1_outputs(2840)) xor (layer1_outputs(1682));
    layer2_outputs(2072) <= not(layer1_outputs(6625));
    layer2_outputs(2073) <= (layer1_outputs(4031)) or (layer1_outputs(1402));
    layer2_outputs(2074) <= not(layer1_outputs(4029));
    layer2_outputs(2075) <= not(layer1_outputs(7057));
    layer2_outputs(2076) <= (layer1_outputs(6579)) and not (layer1_outputs(4407));
    layer2_outputs(2077) <= not(layer1_outputs(5505));
    layer2_outputs(2078) <= not((layer1_outputs(2157)) and (layer1_outputs(2626)));
    layer2_outputs(2079) <= layer1_outputs(3970);
    layer2_outputs(2080) <= layer1_outputs(4720);
    layer2_outputs(2081) <= (layer1_outputs(6082)) and not (layer1_outputs(4433));
    layer2_outputs(2082) <= (layer1_outputs(2925)) xor (layer1_outputs(137));
    layer2_outputs(2083) <= (layer1_outputs(3084)) and not (layer1_outputs(5969));
    layer2_outputs(2084) <= '1';
    layer2_outputs(2085) <= not(layer1_outputs(6439));
    layer2_outputs(2086) <= '1';
    layer2_outputs(2087) <= not(layer1_outputs(1071)) or (layer1_outputs(4089));
    layer2_outputs(2088) <= not((layer1_outputs(1896)) or (layer1_outputs(6373)));
    layer2_outputs(2089) <= not(layer1_outputs(5630)) or (layer1_outputs(1853));
    layer2_outputs(2090) <= not((layer1_outputs(1412)) and (layer1_outputs(6222)));
    layer2_outputs(2091) <= (layer1_outputs(990)) and not (layer1_outputs(2668));
    layer2_outputs(2092) <= (layer1_outputs(7435)) or (layer1_outputs(3357));
    layer2_outputs(2093) <= not(layer1_outputs(911));
    layer2_outputs(2094) <= not(layer1_outputs(607)) or (layer1_outputs(1654));
    layer2_outputs(2095) <= not(layer1_outputs(4721)) or (layer1_outputs(6963));
    layer2_outputs(2096) <= layer1_outputs(557);
    layer2_outputs(2097) <= not((layer1_outputs(6454)) or (layer1_outputs(3776)));
    layer2_outputs(2098) <= (layer1_outputs(3839)) xor (layer1_outputs(5179));
    layer2_outputs(2099) <= layer1_outputs(6016);
    layer2_outputs(2100) <= not(layer1_outputs(6574));
    layer2_outputs(2101) <= not(layer1_outputs(308)) or (layer1_outputs(4374));
    layer2_outputs(2102) <= not((layer1_outputs(2047)) xor (layer1_outputs(4155)));
    layer2_outputs(2103) <= layer1_outputs(324);
    layer2_outputs(2104) <= not(layer1_outputs(6386));
    layer2_outputs(2105) <= layer1_outputs(7306);
    layer2_outputs(2106) <= not(layer1_outputs(1978));
    layer2_outputs(2107) <= (layer1_outputs(3855)) and not (layer1_outputs(4829));
    layer2_outputs(2108) <= (layer1_outputs(4148)) and not (layer1_outputs(919));
    layer2_outputs(2109) <= layer1_outputs(3293);
    layer2_outputs(2110) <= layer1_outputs(7015);
    layer2_outputs(2111) <= layer1_outputs(5556);
    layer2_outputs(2112) <= (layer1_outputs(6953)) and (layer1_outputs(902));
    layer2_outputs(2113) <= not((layer1_outputs(1886)) and (layer1_outputs(1811)));
    layer2_outputs(2114) <= layer1_outputs(5500);
    layer2_outputs(2115) <= (layer1_outputs(2949)) or (layer1_outputs(5248));
    layer2_outputs(2116) <= '0';
    layer2_outputs(2117) <= (layer1_outputs(927)) and (layer1_outputs(4418));
    layer2_outputs(2118) <= not(layer1_outputs(1435)) or (layer1_outputs(3412));
    layer2_outputs(2119) <= (layer1_outputs(5983)) and (layer1_outputs(3255));
    layer2_outputs(2120) <= not(layer1_outputs(7354)) or (layer1_outputs(7370));
    layer2_outputs(2121) <= (layer1_outputs(4039)) and (layer1_outputs(3514));
    layer2_outputs(2122) <= not(layer1_outputs(3845));
    layer2_outputs(2123) <= not(layer1_outputs(7170));
    layer2_outputs(2124) <= (layer1_outputs(3820)) and not (layer1_outputs(465));
    layer2_outputs(2125) <= layer1_outputs(2630);
    layer2_outputs(2126) <= not(layer1_outputs(4365)) or (layer1_outputs(1352));
    layer2_outputs(2127) <= (layer1_outputs(6406)) and not (layer1_outputs(3816));
    layer2_outputs(2128) <= not(layer1_outputs(489)) or (layer1_outputs(6393));
    layer2_outputs(2129) <= (layer1_outputs(429)) xor (layer1_outputs(5270));
    layer2_outputs(2130) <= layer1_outputs(5112);
    layer2_outputs(2131) <= (layer1_outputs(2196)) and (layer1_outputs(276));
    layer2_outputs(2132) <= not(layer1_outputs(947));
    layer2_outputs(2133) <= (layer1_outputs(5033)) and (layer1_outputs(98));
    layer2_outputs(2134) <= not(layer1_outputs(3573));
    layer2_outputs(2135) <= (layer1_outputs(5998)) or (layer1_outputs(3858));
    layer2_outputs(2136) <= layer1_outputs(2676);
    layer2_outputs(2137) <= '1';
    layer2_outputs(2138) <= (layer1_outputs(6202)) and (layer1_outputs(6976));
    layer2_outputs(2139) <= not(layer1_outputs(2683)) or (layer1_outputs(445));
    layer2_outputs(2140) <= (layer1_outputs(7540)) and (layer1_outputs(513));
    layer2_outputs(2141) <= '1';
    layer2_outputs(2142) <= layer1_outputs(4298);
    layer2_outputs(2143) <= layer1_outputs(3963);
    layer2_outputs(2144) <= (layer1_outputs(5974)) or (layer1_outputs(7600));
    layer2_outputs(2145) <= not((layer1_outputs(7373)) or (layer1_outputs(7358)));
    layer2_outputs(2146) <= not(layer1_outputs(2861));
    layer2_outputs(2147) <= (layer1_outputs(1144)) and (layer1_outputs(14));
    layer2_outputs(2148) <= '0';
    layer2_outputs(2149) <= not(layer1_outputs(1379));
    layer2_outputs(2150) <= (layer1_outputs(3490)) and (layer1_outputs(2389));
    layer2_outputs(2151) <= not((layer1_outputs(5463)) and (layer1_outputs(4881)));
    layer2_outputs(2152) <= (layer1_outputs(4535)) and (layer1_outputs(609));
    layer2_outputs(2153) <= not((layer1_outputs(365)) xor (layer1_outputs(2072)));
    layer2_outputs(2154) <= not(layer1_outputs(1335));
    layer2_outputs(2155) <= not(layer1_outputs(5655)) or (layer1_outputs(3817));
    layer2_outputs(2156) <= (layer1_outputs(5575)) and not (layer1_outputs(6175));
    layer2_outputs(2157) <= layer1_outputs(6243);
    layer2_outputs(2158) <= (layer1_outputs(5423)) and (layer1_outputs(3989));
    layer2_outputs(2159) <= not((layer1_outputs(882)) or (layer1_outputs(7407)));
    layer2_outputs(2160) <= not(layer1_outputs(6222));
    layer2_outputs(2161) <= not(layer1_outputs(2771));
    layer2_outputs(2162) <= '1';
    layer2_outputs(2163) <= not((layer1_outputs(7163)) xor (layer1_outputs(4158)));
    layer2_outputs(2164) <= (layer1_outputs(6292)) and (layer1_outputs(323));
    layer2_outputs(2165) <= layer1_outputs(6234);
    layer2_outputs(2166) <= (layer1_outputs(1299)) and not (layer1_outputs(571));
    layer2_outputs(2167) <= layer1_outputs(1697);
    layer2_outputs(2168) <= '0';
    layer2_outputs(2169) <= not(layer1_outputs(6676));
    layer2_outputs(2170) <= not(layer1_outputs(2777));
    layer2_outputs(2171) <= (layer1_outputs(2116)) and (layer1_outputs(573));
    layer2_outputs(2172) <= not((layer1_outputs(2335)) or (layer1_outputs(1897)));
    layer2_outputs(2173) <= not((layer1_outputs(329)) or (layer1_outputs(7518)));
    layer2_outputs(2174) <= not((layer1_outputs(7628)) or (layer1_outputs(4778)));
    layer2_outputs(2175) <= (layer1_outputs(1517)) or (layer1_outputs(7167));
    layer2_outputs(2176) <= (layer1_outputs(6987)) and not (layer1_outputs(7455));
    layer2_outputs(2177) <= not(layer1_outputs(4041));
    layer2_outputs(2178) <= layer1_outputs(4743);
    layer2_outputs(2179) <= not((layer1_outputs(6721)) and (layer1_outputs(7342)));
    layer2_outputs(2180) <= (layer1_outputs(4551)) or (layer1_outputs(2780));
    layer2_outputs(2181) <= layer1_outputs(3067);
    layer2_outputs(2182) <= (layer1_outputs(3351)) and (layer1_outputs(3604));
    layer2_outputs(2183) <= layer1_outputs(1749);
    layer2_outputs(2184) <= not((layer1_outputs(924)) and (layer1_outputs(5876)));
    layer2_outputs(2185) <= (layer1_outputs(5102)) and not (layer1_outputs(5935));
    layer2_outputs(2186) <= not(layer1_outputs(1474));
    layer2_outputs(2187) <= layer1_outputs(1769);
    layer2_outputs(2188) <= layer1_outputs(5046);
    layer2_outputs(2189) <= not((layer1_outputs(5196)) xor (layer1_outputs(3420)));
    layer2_outputs(2190) <= not((layer1_outputs(2608)) and (layer1_outputs(5419)));
    layer2_outputs(2191) <= layer1_outputs(2199);
    layer2_outputs(2192) <= (layer1_outputs(3598)) and (layer1_outputs(3414));
    layer2_outputs(2193) <= not(layer1_outputs(3214));
    layer2_outputs(2194) <= (layer1_outputs(2412)) or (layer1_outputs(6839));
    layer2_outputs(2195) <= not((layer1_outputs(4723)) xor (layer1_outputs(6989)));
    layer2_outputs(2196) <= not(layer1_outputs(1396)) or (layer1_outputs(3637));
    layer2_outputs(2197) <= (layer1_outputs(5024)) and not (layer1_outputs(2440));
    layer2_outputs(2198) <= (layer1_outputs(288)) and not (layer1_outputs(6706));
    layer2_outputs(2199) <= not(layer1_outputs(4244));
    layer2_outputs(2200) <= (layer1_outputs(572)) and not (layer1_outputs(944));
    layer2_outputs(2201) <= not(layer1_outputs(348));
    layer2_outputs(2202) <= not(layer1_outputs(3104));
    layer2_outputs(2203) <= not((layer1_outputs(3600)) xor (layer1_outputs(2858)));
    layer2_outputs(2204) <= (layer1_outputs(3947)) and not (layer1_outputs(4417));
    layer2_outputs(2205) <= layer1_outputs(3353);
    layer2_outputs(2206) <= not(layer1_outputs(5481)) or (layer1_outputs(7671));
    layer2_outputs(2207) <= not(layer1_outputs(6796));
    layer2_outputs(2208) <= not(layer1_outputs(321)) or (layer1_outputs(1993));
    layer2_outputs(2209) <= not(layer1_outputs(2723)) or (layer1_outputs(3269));
    layer2_outputs(2210) <= not(layer1_outputs(2158));
    layer2_outputs(2211) <= layer1_outputs(2404);
    layer2_outputs(2212) <= not(layer1_outputs(5145));
    layer2_outputs(2213) <= (layer1_outputs(4293)) and not (layer1_outputs(2396));
    layer2_outputs(2214) <= (layer1_outputs(6250)) xor (layer1_outputs(7525));
    layer2_outputs(2215) <= not(layer1_outputs(6692)) or (layer1_outputs(5831));
    layer2_outputs(2216) <= not((layer1_outputs(3499)) or (layer1_outputs(6337)));
    layer2_outputs(2217) <= layer1_outputs(4577);
    layer2_outputs(2218) <= (layer1_outputs(584)) and not (layer1_outputs(2106));
    layer2_outputs(2219) <= not(layer1_outputs(3888));
    layer2_outputs(2220) <= '1';
    layer2_outputs(2221) <= not(layer1_outputs(797)) or (layer1_outputs(1217));
    layer2_outputs(2222) <= (layer1_outputs(2042)) and not (layer1_outputs(541));
    layer2_outputs(2223) <= (layer1_outputs(6506)) xor (layer1_outputs(1168));
    layer2_outputs(2224) <= (layer1_outputs(6099)) and not (layer1_outputs(2755));
    layer2_outputs(2225) <= '1';
    layer2_outputs(2226) <= layer1_outputs(511);
    layer2_outputs(2227) <= not(layer1_outputs(5327)) or (layer1_outputs(3296));
    layer2_outputs(2228) <= not(layer1_outputs(487)) or (layer1_outputs(415));
    layer2_outputs(2229) <= not((layer1_outputs(26)) or (layer1_outputs(2243)));
    layer2_outputs(2230) <= not(layer1_outputs(322)) or (layer1_outputs(76));
    layer2_outputs(2231) <= not((layer1_outputs(5287)) xor (layer1_outputs(2848)));
    layer2_outputs(2232) <= (layer1_outputs(964)) and not (layer1_outputs(2349));
    layer2_outputs(2233) <= layer1_outputs(3477);
    layer2_outputs(2234) <= '1';
    layer2_outputs(2235) <= '0';
    layer2_outputs(2236) <= not((layer1_outputs(467)) and (layer1_outputs(3163)));
    layer2_outputs(2237) <= (layer1_outputs(4228)) and not (layer1_outputs(63));
    layer2_outputs(2238) <= '1';
    layer2_outputs(2239) <= (layer1_outputs(2179)) or (layer1_outputs(5193));
    layer2_outputs(2240) <= '1';
    layer2_outputs(2241) <= not((layer1_outputs(6029)) and (layer1_outputs(7624)));
    layer2_outputs(2242) <= not(layer1_outputs(6955));
    layer2_outputs(2243) <= layer1_outputs(1147);
    layer2_outputs(2244) <= '0';
    layer2_outputs(2245) <= layer1_outputs(7070);
    layer2_outputs(2246) <= not(layer1_outputs(5887));
    layer2_outputs(2247) <= not(layer1_outputs(7252));
    layer2_outputs(2248) <= not(layer1_outputs(1169));
    layer2_outputs(2249) <= not((layer1_outputs(731)) and (layer1_outputs(2667)));
    layer2_outputs(2250) <= not(layer1_outputs(6361));
    layer2_outputs(2251) <= (layer1_outputs(5582)) and (layer1_outputs(2436));
    layer2_outputs(2252) <= (layer1_outputs(2694)) and not (layer1_outputs(4893));
    layer2_outputs(2253) <= not(layer1_outputs(1275));
    layer2_outputs(2254) <= '1';
    layer2_outputs(2255) <= not(layer1_outputs(3193));
    layer2_outputs(2256) <= (layer1_outputs(5991)) and not (layer1_outputs(1399));
    layer2_outputs(2257) <= (layer1_outputs(3711)) and not (layer1_outputs(4768));
    layer2_outputs(2258) <= not(layer1_outputs(3934)) or (layer1_outputs(6518));
    layer2_outputs(2259) <= (layer1_outputs(4121)) and not (layer1_outputs(4151));
    layer2_outputs(2260) <= (layer1_outputs(3828)) and (layer1_outputs(2574));
    layer2_outputs(2261) <= not((layer1_outputs(3575)) and (layer1_outputs(906)));
    layer2_outputs(2262) <= layer1_outputs(5531);
    layer2_outputs(2263) <= not(layer1_outputs(1100));
    layer2_outputs(2264) <= not((layer1_outputs(4019)) and (layer1_outputs(5208)));
    layer2_outputs(2265) <= not(layer1_outputs(53));
    layer2_outputs(2266) <= (layer1_outputs(6143)) and (layer1_outputs(2143));
    layer2_outputs(2267) <= layer1_outputs(2861);
    layer2_outputs(2268) <= (layer1_outputs(6695)) and not (layer1_outputs(4507));
    layer2_outputs(2269) <= not(layer1_outputs(2539));
    layer2_outputs(2270) <= not(layer1_outputs(2862));
    layer2_outputs(2271) <= (layer1_outputs(757)) xor (layer1_outputs(3207));
    layer2_outputs(2272) <= '0';
    layer2_outputs(2273) <= not((layer1_outputs(7244)) or (layer1_outputs(3406)));
    layer2_outputs(2274) <= not(layer1_outputs(7558));
    layer2_outputs(2275) <= '0';
    layer2_outputs(2276) <= layer1_outputs(4470);
    layer2_outputs(2277) <= layer1_outputs(876);
    layer2_outputs(2278) <= '1';
    layer2_outputs(2279) <= (layer1_outputs(4730)) and not (layer1_outputs(2236));
    layer2_outputs(2280) <= not((layer1_outputs(4852)) or (layer1_outputs(7097)));
    layer2_outputs(2281) <= not(layer1_outputs(5766));
    layer2_outputs(2282) <= not((layer1_outputs(4179)) and (layer1_outputs(560)));
    layer2_outputs(2283) <= layer1_outputs(6296);
    layer2_outputs(2284) <= (layer1_outputs(6277)) and not (layer1_outputs(4301));
    layer2_outputs(2285) <= not(layer1_outputs(6596)) or (layer1_outputs(1616));
    layer2_outputs(2286) <= '1';
    layer2_outputs(2287) <= '1';
    layer2_outputs(2288) <= not((layer1_outputs(2885)) or (layer1_outputs(3313)));
    layer2_outputs(2289) <= not(layer1_outputs(3669));
    layer2_outputs(2290) <= (layer1_outputs(7497)) or (layer1_outputs(1254));
    layer2_outputs(2291) <= not((layer1_outputs(4244)) and (layer1_outputs(5857)));
    layer2_outputs(2292) <= (layer1_outputs(4718)) and not (layer1_outputs(2518));
    layer2_outputs(2293) <= layer1_outputs(2524);
    layer2_outputs(2294) <= (layer1_outputs(97)) and not (layer1_outputs(5473));
    layer2_outputs(2295) <= not((layer1_outputs(6012)) and (layer1_outputs(295)));
    layer2_outputs(2296) <= (layer1_outputs(7413)) and not (layer1_outputs(545));
    layer2_outputs(2297) <= not((layer1_outputs(4316)) or (layer1_outputs(6505)));
    layer2_outputs(2298) <= not(layer1_outputs(228));
    layer2_outputs(2299) <= not(layer1_outputs(4877)) or (layer1_outputs(3867));
    layer2_outputs(2300) <= (layer1_outputs(183)) and not (layer1_outputs(3012));
    layer2_outputs(2301) <= not((layer1_outputs(554)) and (layer1_outputs(7253)));
    layer2_outputs(2302) <= (layer1_outputs(2640)) or (layer1_outputs(3262));
    layer2_outputs(2303) <= layer1_outputs(4891);
    layer2_outputs(2304) <= not((layer1_outputs(5185)) or (layer1_outputs(1761)));
    layer2_outputs(2305) <= not(layer1_outputs(1812)) or (layer1_outputs(300));
    layer2_outputs(2306) <= (layer1_outputs(7471)) and not (layer1_outputs(262));
    layer2_outputs(2307) <= not((layer1_outputs(3044)) and (layer1_outputs(6235)));
    layer2_outputs(2308) <= (layer1_outputs(7545)) or (layer1_outputs(1872));
    layer2_outputs(2309) <= layer1_outputs(4426);
    layer2_outputs(2310) <= not((layer1_outputs(3976)) or (layer1_outputs(1102)));
    layer2_outputs(2311) <= not((layer1_outputs(7616)) or (layer1_outputs(6853)));
    layer2_outputs(2312) <= (layer1_outputs(1365)) and not (layer1_outputs(3973));
    layer2_outputs(2313) <= not(layer1_outputs(4047)) or (layer1_outputs(3199));
    layer2_outputs(2314) <= not(layer1_outputs(1982));
    layer2_outputs(2315) <= (layer1_outputs(6737)) and (layer1_outputs(3683));
    layer2_outputs(2316) <= not((layer1_outputs(4115)) or (layer1_outputs(203)));
    layer2_outputs(2317) <= not(layer1_outputs(6878));
    layer2_outputs(2318) <= (layer1_outputs(3637)) and (layer1_outputs(5301));
    layer2_outputs(2319) <= layer1_outputs(1782);
    layer2_outputs(2320) <= not(layer1_outputs(2640)) or (layer1_outputs(499));
    layer2_outputs(2321) <= layer1_outputs(214);
    layer2_outputs(2322) <= layer1_outputs(5226);
    layer2_outputs(2323) <= layer1_outputs(4482);
    layer2_outputs(2324) <= layer1_outputs(4904);
    layer2_outputs(2325) <= layer1_outputs(1613);
    layer2_outputs(2326) <= not((layer1_outputs(2517)) or (layer1_outputs(2114)));
    layer2_outputs(2327) <= layer1_outputs(7404);
    layer2_outputs(2328) <= not(layer1_outputs(3533));
    layer2_outputs(2329) <= '0';
    layer2_outputs(2330) <= not(layer1_outputs(772));
    layer2_outputs(2331) <= not(layer1_outputs(4742)) or (layer1_outputs(4258));
    layer2_outputs(2332) <= not(layer1_outputs(1161)) or (layer1_outputs(2358));
    layer2_outputs(2333) <= not(layer1_outputs(3541));
    layer2_outputs(2334) <= (layer1_outputs(4686)) and not (layer1_outputs(6391));
    layer2_outputs(2335) <= (layer1_outputs(316)) and (layer1_outputs(6251));
    layer2_outputs(2336) <= not((layer1_outputs(821)) and (layer1_outputs(7096)));
    layer2_outputs(2337) <= not(layer1_outputs(7292));
    layer2_outputs(2338) <= not(layer1_outputs(3337));
    layer2_outputs(2339) <= (layer1_outputs(890)) and not (layer1_outputs(6681));
    layer2_outputs(2340) <= not((layer1_outputs(3391)) and (layer1_outputs(6073)));
    layer2_outputs(2341) <= not(layer1_outputs(7490)) or (layer1_outputs(1479));
    layer2_outputs(2342) <= (layer1_outputs(687)) xor (layer1_outputs(5469));
    layer2_outputs(2343) <= (layer1_outputs(1853)) and not (layer1_outputs(3778));
    layer2_outputs(2344) <= (layer1_outputs(428)) and (layer1_outputs(7266));
    layer2_outputs(2345) <= not(layer1_outputs(5555));
    layer2_outputs(2346) <= (layer1_outputs(4590)) and not (layer1_outputs(1538));
    layer2_outputs(2347) <= (layer1_outputs(298)) xor (layer1_outputs(2657));
    layer2_outputs(2348) <= (layer1_outputs(4788)) or (layer1_outputs(5587));
    layer2_outputs(2349) <= (layer1_outputs(600)) and not (layer1_outputs(2530));
    layer2_outputs(2350) <= '1';
    layer2_outputs(2351) <= not(layer1_outputs(6564));
    layer2_outputs(2352) <= not(layer1_outputs(3293)) or (layer1_outputs(890));
    layer2_outputs(2353) <= not(layer1_outputs(1515));
    layer2_outputs(2354) <= not((layer1_outputs(6217)) or (layer1_outputs(5350)));
    layer2_outputs(2355) <= not(layer1_outputs(12));
    layer2_outputs(2356) <= not(layer1_outputs(5901)) or (layer1_outputs(5099));
    layer2_outputs(2357) <= not((layer1_outputs(453)) or (layer1_outputs(1171)));
    layer2_outputs(2358) <= (layer1_outputs(2930)) or (layer1_outputs(3860));
    layer2_outputs(2359) <= (layer1_outputs(4589)) and not (layer1_outputs(6620));
    layer2_outputs(2360) <= not((layer1_outputs(3443)) and (layer1_outputs(7060)));
    layer2_outputs(2361) <= not(layer1_outputs(5518));
    layer2_outputs(2362) <= (layer1_outputs(6038)) and (layer1_outputs(1230));
    layer2_outputs(2363) <= not((layer1_outputs(3331)) or (layer1_outputs(3368)));
    layer2_outputs(2364) <= not(layer1_outputs(2107));
    layer2_outputs(2365) <= not(layer1_outputs(4182));
    layer2_outputs(2366) <= not(layer1_outputs(1643));
    layer2_outputs(2367) <= (layer1_outputs(2022)) and (layer1_outputs(2714));
    layer2_outputs(2368) <= (layer1_outputs(5878)) and not (layer1_outputs(4340));
    layer2_outputs(2369) <= not(layer1_outputs(4143));
    layer2_outputs(2370) <= not(layer1_outputs(2739)) or (layer1_outputs(4910));
    layer2_outputs(2371) <= layer1_outputs(657);
    layer2_outputs(2372) <= layer1_outputs(5264);
    layer2_outputs(2373) <= (layer1_outputs(3580)) or (layer1_outputs(5779));
    layer2_outputs(2374) <= not(layer1_outputs(4289));
    layer2_outputs(2375) <= (layer1_outputs(4138)) and not (layer1_outputs(3916));
    layer2_outputs(2376) <= (layer1_outputs(828)) and not (layer1_outputs(1358));
    layer2_outputs(2377) <= layer1_outputs(4658);
    layer2_outputs(2378) <= (layer1_outputs(4188)) and not (layer1_outputs(480));
    layer2_outputs(2379) <= not(layer1_outputs(6012)) or (layer1_outputs(7285));
    layer2_outputs(2380) <= (layer1_outputs(4984)) and (layer1_outputs(5585));
    layer2_outputs(2381) <= not((layer1_outputs(5136)) or (layer1_outputs(2774)));
    layer2_outputs(2382) <= layer1_outputs(2105);
    layer2_outputs(2383) <= not((layer1_outputs(6413)) or (layer1_outputs(2363)));
    layer2_outputs(2384) <= not(layer1_outputs(53));
    layer2_outputs(2385) <= (layer1_outputs(3985)) or (layer1_outputs(3503));
    layer2_outputs(2386) <= (layer1_outputs(4951)) xor (layer1_outputs(56));
    layer2_outputs(2387) <= (layer1_outputs(3429)) xor (layer1_outputs(1563));
    layer2_outputs(2388) <= (layer1_outputs(6666)) and not (layer1_outputs(5251));
    layer2_outputs(2389) <= (layer1_outputs(6799)) and (layer1_outputs(5621));
    layer2_outputs(2390) <= not(layer1_outputs(4980));
    layer2_outputs(2391) <= (layer1_outputs(7667)) and not (layer1_outputs(3898));
    layer2_outputs(2392) <= not((layer1_outputs(6651)) xor (layer1_outputs(7318)));
    layer2_outputs(2393) <= (layer1_outputs(6168)) and not (layer1_outputs(7002));
    layer2_outputs(2394) <= layer1_outputs(3472);
    layer2_outputs(2395) <= '1';
    layer2_outputs(2396) <= layer1_outputs(204);
    layer2_outputs(2397) <= not(layer1_outputs(7115)) or (layer1_outputs(5701));
    layer2_outputs(2398) <= '1';
    layer2_outputs(2399) <= (layer1_outputs(3130)) and not (layer1_outputs(7042));
    layer2_outputs(2400) <= not(layer1_outputs(805));
    layer2_outputs(2401) <= layer1_outputs(7040);
    layer2_outputs(2402) <= (layer1_outputs(398)) and not (layer1_outputs(2500));
    layer2_outputs(2403) <= (layer1_outputs(1751)) and not (layer1_outputs(5443));
    layer2_outputs(2404) <= layer1_outputs(7420);
    layer2_outputs(2405) <= layer1_outputs(4009);
    layer2_outputs(2406) <= layer1_outputs(6938);
    layer2_outputs(2407) <= not((layer1_outputs(2013)) xor (layer1_outputs(7514)));
    layer2_outputs(2408) <= not(layer1_outputs(1895));
    layer2_outputs(2409) <= layer1_outputs(5161);
    layer2_outputs(2410) <= (layer1_outputs(4731)) and (layer1_outputs(462));
    layer2_outputs(2411) <= (layer1_outputs(7455)) or (layer1_outputs(328));
    layer2_outputs(2412) <= not(layer1_outputs(662));
    layer2_outputs(2413) <= not((layer1_outputs(6753)) and (layer1_outputs(1058)));
    layer2_outputs(2414) <= '0';
    layer2_outputs(2415) <= not((layer1_outputs(6110)) or (layer1_outputs(1097)));
    layer2_outputs(2416) <= (layer1_outputs(3892)) and not (layer1_outputs(3583));
    layer2_outputs(2417) <= (layer1_outputs(4629)) and not (layer1_outputs(4287));
    layer2_outputs(2418) <= (layer1_outputs(5169)) and (layer1_outputs(598));
    layer2_outputs(2419) <= not(layer1_outputs(3691));
    layer2_outputs(2420) <= layer1_outputs(4391);
    layer2_outputs(2421) <= (layer1_outputs(642)) and (layer1_outputs(3867));
    layer2_outputs(2422) <= layer1_outputs(5608);
    layer2_outputs(2423) <= '0';
    layer2_outputs(2424) <= not(layer1_outputs(1324));
    layer2_outputs(2425) <= not(layer1_outputs(3224));
    layer2_outputs(2426) <= layer1_outputs(1508);
    layer2_outputs(2427) <= (layer1_outputs(2807)) and not (layer1_outputs(1800));
    layer2_outputs(2428) <= '0';
    layer2_outputs(2429) <= not(layer1_outputs(1368)) or (layer1_outputs(3758));
    layer2_outputs(2430) <= layer1_outputs(1243);
    layer2_outputs(2431) <= not((layer1_outputs(2880)) and (layer1_outputs(6137)));
    layer2_outputs(2432) <= not(layer1_outputs(1739)) or (layer1_outputs(1025));
    layer2_outputs(2433) <= not(layer1_outputs(5510));
    layer2_outputs(2434) <= '1';
    layer2_outputs(2435) <= not(layer1_outputs(506));
    layer2_outputs(2436) <= not(layer1_outputs(5349));
    layer2_outputs(2437) <= layer1_outputs(1701);
    layer2_outputs(2438) <= layer1_outputs(1984);
    layer2_outputs(2439) <= layer1_outputs(5871);
    layer2_outputs(2440) <= not(layer1_outputs(234));
    layer2_outputs(2441) <= not(layer1_outputs(2162));
    layer2_outputs(2442) <= not((layer1_outputs(139)) and (layer1_outputs(5216)));
    layer2_outputs(2443) <= (layer1_outputs(6021)) or (layer1_outputs(7197));
    layer2_outputs(2444) <= layer1_outputs(6918);
    layer2_outputs(2445) <= (layer1_outputs(2750)) and not (layer1_outputs(6915));
    layer2_outputs(2446) <= not((layer1_outputs(2646)) or (layer1_outputs(5857)));
    layer2_outputs(2447) <= not(layer1_outputs(169));
    layer2_outputs(2448) <= not(layer1_outputs(6445)) or (layer1_outputs(7322));
    layer2_outputs(2449) <= not(layer1_outputs(470));
    layer2_outputs(2450) <= not((layer1_outputs(692)) or (layer1_outputs(6770)));
    layer2_outputs(2451) <= not((layer1_outputs(6026)) and (layer1_outputs(4740)));
    layer2_outputs(2452) <= not((layer1_outputs(5306)) or (layer1_outputs(5093)));
    layer2_outputs(2453) <= not((layer1_outputs(970)) or (layer1_outputs(1525)));
    layer2_outputs(2454) <= '0';
    layer2_outputs(2455) <= (layer1_outputs(5155)) and (layer1_outputs(3137));
    layer2_outputs(2456) <= (layer1_outputs(7494)) or (layer1_outputs(6209));
    layer2_outputs(2457) <= layer1_outputs(4825);
    layer2_outputs(2458) <= layer1_outputs(4607);
    layer2_outputs(2459) <= layer1_outputs(5215);
    layer2_outputs(2460) <= not((layer1_outputs(5807)) or (layer1_outputs(6300)));
    layer2_outputs(2461) <= (layer1_outputs(5670)) and not (layer1_outputs(4616));
    layer2_outputs(2462) <= not((layer1_outputs(4153)) and (layer1_outputs(5095)));
    layer2_outputs(2463) <= not(layer1_outputs(4382)) or (layer1_outputs(969));
    layer2_outputs(2464) <= not(layer1_outputs(6203));
    layer2_outputs(2465) <= not(layer1_outputs(754));
    layer2_outputs(2466) <= not(layer1_outputs(5954));
    layer2_outputs(2467) <= not(layer1_outputs(5047));
    layer2_outputs(2468) <= (layer1_outputs(4419)) and (layer1_outputs(6034));
    layer2_outputs(2469) <= layer1_outputs(6404);
    layer2_outputs(2470) <= not(layer1_outputs(1367)) or (layer1_outputs(1085));
    layer2_outputs(2471) <= not((layer1_outputs(2017)) or (layer1_outputs(5597)));
    layer2_outputs(2472) <= '1';
    layer2_outputs(2473) <= not((layer1_outputs(7542)) or (layer1_outputs(2204)));
    layer2_outputs(2474) <= not(layer1_outputs(979));
    layer2_outputs(2475) <= layer1_outputs(2257);
    layer2_outputs(2476) <= not(layer1_outputs(3276));
    layer2_outputs(2477) <= layer1_outputs(6219);
    layer2_outputs(2478) <= not((layer1_outputs(4477)) or (layer1_outputs(6094)));
    layer2_outputs(2479) <= (layer1_outputs(3941)) xor (layer1_outputs(2238));
    layer2_outputs(2480) <= not(layer1_outputs(7533));
    layer2_outputs(2481) <= layer1_outputs(5492);
    layer2_outputs(2482) <= '1';
    layer2_outputs(2483) <= layer1_outputs(3482);
    layer2_outputs(2484) <= not(layer1_outputs(5976)) or (layer1_outputs(1528));
    layer2_outputs(2485) <= layer1_outputs(4460);
    layer2_outputs(2486) <= layer1_outputs(2074);
    layer2_outputs(2487) <= not(layer1_outputs(144)) or (layer1_outputs(7535));
    layer2_outputs(2488) <= layer1_outputs(2020);
    layer2_outputs(2489) <= (layer1_outputs(3168)) or (layer1_outputs(4112));
    layer2_outputs(2490) <= not(layer1_outputs(4687));
    layer2_outputs(2491) <= layer1_outputs(735);
    layer2_outputs(2492) <= not(layer1_outputs(4727)) or (layer1_outputs(1590));
    layer2_outputs(2493) <= (layer1_outputs(4017)) or (layer1_outputs(4436));
    layer2_outputs(2494) <= not((layer1_outputs(5745)) and (layer1_outputs(3008)));
    layer2_outputs(2495) <= (layer1_outputs(1104)) and (layer1_outputs(2833));
    layer2_outputs(2496) <= (layer1_outputs(3319)) and not (layer1_outputs(5733));
    layer2_outputs(2497) <= not((layer1_outputs(4241)) or (layer1_outputs(615)));
    layer2_outputs(2498) <= layer1_outputs(6639);
    layer2_outputs(2499) <= not(layer1_outputs(1922)) or (layer1_outputs(5933));
    layer2_outputs(2500) <= not((layer1_outputs(1302)) and (layer1_outputs(3608)));
    layer2_outputs(2501) <= not((layer1_outputs(2394)) or (layer1_outputs(1741)));
    layer2_outputs(2502) <= not((layer1_outputs(4485)) or (layer1_outputs(165)));
    layer2_outputs(2503) <= not(layer1_outputs(6566));
    layer2_outputs(2504) <= layer1_outputs(4605);
    layer2_outputs(2505) <= not(layer1_outputs(55));
    layer2_outputs(2506) <= not(layer1_outputs(5908));
    layer2_outputs(2507) <= not(layer1_outputs(835));
    layer2_outputs(2508) <= not((layer1_outputs(6066)) xor (layer1_outputs(5089)));
    layer2_outputs(2509) <= not((layer1_outputs(1541)) xor (layer1_outputs(1947)));
    layer2_outputs(2510) <= not(layer1_outputs(7611));
    layer2_outputs(2511) <= layer1_outputs(5133);
    layer2_outputs(2512) <= not(layer1_outputs(3886));
    layer2_outputs(2513) <= not(layer1_outputs(1359)) or (layer1_outputs(3283));
    layer2_outputs(2514) <= layer1_outputs(2879);
    layer2_outputs(2515) <= not(layer1_outputs(5607));
    layer2_outputs(2516) <= layer1_outputs(1385);
    layer2_outputs(2517) <= not((layer1_outputs(1303)) and (layer1_outputs(4073)));
    layer2_outputs(2518) <= (layer1_outputs(3138)) and not (layer1_outputs(520));
    layer2_outputs(2519) <= layer1_outputs(727);
    layer2_outputs(2520) <= layer1_outputs(7041);
    layer2_outputs(2521) <= not(layer1_outputs(5374)) or (layer1_outputs(4067));
    layer2_outputs(2522) <= (layer1_outputs(2825)) and (layer1_outputs(4477));
    layer2_outputs(2523) <= not(layer1_outputs(2409)) or (layer1_outputs(2269));
    layer2_outputs(2524) <= not(layer1_outputs(4818)) or (layer1_outputs(3443));
    layer2_outputs(2525) <= not((layer1_outputs(1805)) or (layer1_outputs(7536)));
    layer2_outputs(2526) <= (layer1_outputs(4791)) and not (layer1_outputs(5762));
    layer2_outputs(2527) <= not(layer1_outputs(2057));
    layer2_outputs(2528) <= not((layer1_outputs(3802)) or (layer1_outputs(1838)));
    layer2_outputs(2529) <= not((layer1_outputs(2576)) or (layer1_outputs(4650)));
    layer2_outputs(2530) <= not((layer1_outputs(3799)) and (layer1_outputs(1708)));
    layer2_outputs(2531) <= not(layer1_outputs(6982));
    layer2_outputs(2532) <= not(layer1_outputs(7240));
    layer2_outputs(2533) <= not(layer1_outputs(4181));
    layer2_outputs(2534) <= layer1_outputs(6815);
    layer2_outputs(2535) <= layer1_outputs(5333);
    layer2_outputs(2536) <= layer1_outputs(4011);
    layer2_outputs(2537) <= layer1_outputs(16);
    layer2_outputs(2538) <= not(layer1_outputs(3324));
    layer2_outputs(2539) <= (layer1_outputs(4196)) and (layer1_outputs(4878));
    layer2_outputs(2540) <= not(layer1_outputs(391)) or (layer1_outputs(4076));
    layer2_outputs(2541) <= not(layer1_outputs(463));
    layer2_outputs(2542) <= '1';
    layer2_outputs(2543) <= not(layer1_outputs(3506));
    layer2_outputs(2544) <= not(layer1_outputs(233)) or (layer1_outputs(7375));
    layer2_outputs(2545) <= not(layer1_outputs(2673));
    layer2_outputs(2546) <= not(layer1_outputs(1220));
    layer2_outputs(2547) <= not(layer1_outputs(7259)) or (layer1_outputs(1361));
    layer2_outputs(2548) <= (layer1_outputs(1711)) and not (layer1_outputs(2635));
    layer2_outputs(2549) <= '1';
    layer2_outputs(2550) <= not(layer1_outputs(7046));
    layer2_outputs(2551) <= (layer1_outputs(3731)) and not (layer1_outputs(1011));
    layer2_outputs(2552) <= (layer1_outputs(7513)) and not (layer1_outputs(5526));
    layer2_outputs(2553) <= (layer1_outputs(2362)) and (layer1_outputs(3864));
    layer2_outputs(2554) <= (layer1_outputs(67)) and not (layer1_outputs(4097));
    layer2_outputs(2555) <= not(layer1_outputs(2163)) or (layer1_outputs(511));
    layer2_outputs(2556) <= layer1_outputs(7381);
    layer2_outputs(2557) <= not(layer1_outputs(7125));
    layer2_outputs(2558) <= layer1_outputs(3318);
    layer2_outputs(2559) <= not((layer1_outputs(6200)) or (layer1_outputs(1224)));
    layer2_outputs(2560) <= not((layer1_outputs(1689)) and (layer1_outputs(2033)));
    layer2_outputs(2561) <= layer1_outputs(1842);
    layer2_outputs(2562) <= (layer1_outputs(1137)) or (layer1_outputs(2989));
    layer2_outputs(2563) <= (layer1_outputs(4538)) and (layer1_outputs(1759));
    layer2_outputs(2564) <= not((layer1_outputs(5387)) or (layer1_outputs(4271)));
    layer2_outputs(2565) <= not(layer1_outputs(6778)) or (layer1_outputs(2950));
    layer2_outputs(2566) <= not((layer1_outputs(4498)) or (layer1_outputs(7298)));
    layer2_outputs(2567) <= '0';
    layer2_outputs(2568) <= not(layer1_outputs(3204)) or (layer1_outputs(6405));
    layer2_outputs(2569) <= layer1_outputs(2514);
    layer2_outputs(2570) <= not((layer1_outputs(1736)) or (layer1_outputs(2921)));
    layer2_outputs(2571) <= (layer1_outputs(6668)) xor (layer1_outputs(7512));
    layer2_outputs(2572) <= (layer1_outputs(2459)) or (layer1_outputs(2766));
    layer2_outputs(2573) <= not((layer1_outputs(3433)) and (layer1_outputs(2949)));
    layer2_outputs(2574) <= (layer1_outputs(2710)) and not (layer1_outputs(789));
    layer2_outputs(2575) <= (layer1_outputs(4394)) and (layer1_outputs(2156));
    layer2_outputs(2576) <= not(layer1_outputs(3053));
    layer2_outputs(2577) <= (layer1_outputs(1604)) and (layer1_outputs(4018));
    layer2_outputs(2578) <= not((layer1_outputs(583)) xor (layer1_outputs(3258)));
    layer2_outputs(2579) <= not(layer1_outputs(5396));
    layer2_outputs(2580) <= (layer1_outputs(1652)) and not (layer1_outputs(7246));
    layer2_outputs(2581) <= not((layer1_outputs(1861)) or (layer1_outputs(4764)));
    layer2_outputs(2582) <= layer1_outputs(2654);
    layer2_outputs(2583) <= not((layer1_outputs(3181)) and (layer1_outputs(6183)));
    layer2_outputs(2584) <= not(layer1_outputs(2960));
    layer2_outputs(2585) <= not((layer1_outputs(2602)) and (layer1_outputs(5056)));
    layer2_outputs(2586) <= layer1_outputs(24);
    layer2_outputs(2587) <= (layer1_outputs(651)) and not (layer1_outputs(5747));
    layer2_outputs(2588) <= layer1_outputs(3750);
    layer2_outputs(2589) <= layer1_outputs(3447);
    layer2_outputs(2590) <= '0';
    layer2_outputs(2591) <= (layer1_outputs(1459)) or (layer1_outputs(1793));
    layer2_outputs(2592) <= layer1_outputs(3945);
    layer2_outputs(2593) <= not((layer1_outputs(1189)) and (layer1_outputs(2979)));
    layer2_outputs(2594) <= layer1_outputs(1887);
    layer2_outputs(2595) <= not(layer1_outputs(6486));
    layer2_outputs(2596) <= layer1_outputs(6228);
    layer2_outputs(2597) <= layer1_outputs(6944);
    layer2_outputs(2598) <= layer1_outputs(2697);
    layer2_outputs(2599) <= not(layer1_outputs(6157));
    layer2_outputs(2600) <= layer1_outputs(240);
    layer2_outputs(2601) <= not(layer1_outputs(5353)) or (layer1_outputs(1923));
    layer2_outputs(2602) <= not(layer1_outputs(5653));
    layer2_outputs(2603) <= (layer1_outputs(1279)) xor (layer1_outputs(4224));
    layer2_outputs(2604) <= not(layer1_outputs(6955));
    layer2_outputs(2605) <= not((layer1_outputs(4974)) or (layer1_outputs(5395)));
    layer2_outputs(2606) <= (layer1_outputs(6112)) and not (layer1_outputs(3682));
    layer2_outputs(2607) <= not(layer1_outputs(4202)) or (layer1_outputs(7529));
    layer2_outputs(2608) <= not(layer1_outputs(3470)) or (layer1_outputs(4376));
    layer2_outputs(2609) <= layer1_outputs(1165);
    layer2_outputs(2610) <= (layer1_outputs(5506)) and not (layer1_outputs(3853));
    layer2_outputs(2611) <= not(layer1_outputs(6806)) or (layer1_outputs(13));
    layer2_outputs(2612) <= not((layer1_outputs(5221)) or (layer1_outputs(3189)));
    layer2_outputs(2613) <= '1';
    layer2_outputs(2614) <= not((layer1_outputs(4644)) and (layer1_outputs(2028)));
    layer2_outputs(2615) <= (layer1_outputs(3823)) and (layer1_outputs(563));
    layer2_outputs(2616) <= not(layer1_outputs(4114));
    layer2_outputs(2617) <= '1';
    layer2_outputs(2618) <= (layer1_outputs(3120)) and not (layer1_outputs(7285));
    layer2_outputs(2619) <= (layer1_outputs(7126)) and not (layer1_outputs(2754));
    layer2_outputs(2620) <= not(layer1_outputs(3957));
    layer2_outputs(2621) <= not(layer1_outputs(4992));
    layer2_outputs(2622) <= (layer1_outputs(5504)) and (layer1_outputs(6229));
    layer2_outputs(2623) <= layer1_outputs(162);
    layer2_outputs(2624) <= layer1_outputs(6824);
    layer2_outputs(2625) <= not(layer1_outputs(3077));
    layer2_outputs(2626) <= layer1_outputs(6372);
    layer2_outputs(2627) <= (layer1_outputs(5621)) and not (layer1_outputs(5384));
    layer2_outputs(2628) <= layer1_outputs(5905);
    layer2_outputs(2629) <= (layer1_outputs(1422)) or (layer1_outputs(6273));
    layer2_outputs(2630) <= layer1_outputs(5645);
    layer2_outputs(2631) <= '0';
    layer2_outputs(2632) <= (layer1_outputs(1646)) xor (layer1_outputs(3990));
    layer2_outputs(2633) <= not((layer1_outputs(659)) and (layer1_outputs(1363)));
    layer2_outputs(2634) <= layer1_outputs(5411);
    layer2_outputs(2635) <= layer1_outputs(5052);
    layer2_outputs(2636) <= layer1_outputs(4817);
    layer2_outputs(2637) <= not((layer1_outputs(4293)) or (layer1_outputs(1191)));
    layer2_outputs(2638) <= '1';
    layer2_outputs(2639) <= layer1_outputs(4168);
    layer2_outputs(2640) <= not(layer1_outputs(7287)) or (layer1_outputs(2803));
    layer2_outputs(2641) <= layer1_outputs(5606);
    layer2_outputs(2642) <= not(layer1_outputs(1034));
    layer2_outputs(2643) <= layer1_outputs(7005);
    layer2_outputs(2644) <= (layer1_outputs(1734)) and not (layer1_outputs(2950));
    layer2_outputs(2645) <= not(layer1_outputs(5305));
    layer2_outputs(2646) <= layer1_outputs(3307);
    layer2_outputs(2647) <= layer1_outputs(2805);
    layer2_outputs(2648) <= '0';
    layer2_outputs(2649) <= not((layer1_outputs(7498)) and (layer1_outputs(5602)));
    layer2_outputs(2650) <= layer1_outputs(7579);
    layer2_outputs(2651) <= layer1_outputs(1211);
    layer2_outputs(2652) <= not(layer1_outputs(2098));
    layer2_outputs(2653) <= (layer1_outputs(2004)) or (layer1_outputs(3140));
    layer2_outputs(2654) <= layer1_outputs(7307);
    layer2_outputs(2655) <= not(layer1_outputs(1072));
    layer2_outputs(2656) <= not(layer1_outputs(1881));
    layer2_outputs(2657) <= (layer1_outputs(2265)) and (layer1_outputs(3603));
    layer2_outputs(2658) <= (layer1_outputs(5828)) and not (layer1_outputs(6693));
    layer2_outputs(2659) <= not(layer1_outputs(722));
    layer2_outputs(2660) <= not(layer1_outputs(5907)) or (layer1_outputs(4358));
    layer2_outputs(2661) <= not(layer1_outputs(4333));
    layer2_outputs(2662) <= layer1_outputs(630);
    layer2_outputs(2663) <= layer1_outputs(585);
    layer2_outputs(2664) <= (layer1_outputs(5680)) or (layer1_outputs(806));
    layer2_outputs(2665) <= layer1_outputs(5866);
    layer2_outputs(2666) <= not(layer1_outputs(2347)) or (layer1_outputs(4872));
    layer2_outputs(2667) <= '0';
    layer2_outputs(2668) <= '0';
    layer2_outputs(2669) <= layer1_outputs(1237);
    layer2_outputs(2670) <= '1';
    layer2_outputs(2671) <= not(layer1_outputs(5889)) or (layer1_outputs(5453));
    layer2_outputs(2672) <= (layer1_outputs(1133)) and not (layer1_outputs(4965));
    layer2_outputs(2673) <= not(layer1_outputs(4603)) or (layer1_outputs(5700));
    layer2_outputs(2674) <= (layer1_outputs(6646)) and not (layer1_outputs(2056));
    layer2_outputs(2675) <= not(layer1_outputs(2778)) or (layer1_outputs(1527));
    layer2_outputs(2676) <= not((layer1_outputs(1944)) or (layer1_outputs(3441)));
    layer2_outputs(2677) <= layer1_outputs(7400);
    layer2_outputs(2678) <= (layer1_outputs(6126)) and not (layer1_outputs(7653));
    layer2_outputs(2679) <= '0';
    layer2_outputs(2680) <= (layer1_outputs(5225)) and not (layer1_outputs(368));
    layer2_outputs(2681) <= '0';
    layer2_outputs(2682) <= not(layer1_outputs(1427));
    layer2_outputs(2683) <= not(layer1_outputs(4946));
    layer2_outputs(2684) <= (layer1_outputs(3893)) and (layer1_outputs(689));
    layer2_outputs(2685) <= layer1_outputs(3381);
    layer2_outputs(2686) <= not((layer1_outputs(4796)) or (layer1_outputs(7384)));
    layer2_outputs(2687) <= layer1_outputs(7079);
    layer2_outputs(2688) <= not((layer1_outputs(1624)) or (layer1_outputs(7351)));
    layer2_outputs(2689) <= (layer1_outputs(7052)) and not (layer1_outputs(7611));
    layer2_outputs(2690) <= layer1_outputs(7339);
    layer2_outputs(2691) <= (layer1_outputs(74)) or (layer1_outputs(5316));
    layer2_outputs(2692) <= (layer1_outputs(4614)) or (layer1_outputs(313));
    layer2_outputs(2693) <= not(layer1_outputs(6384)) or (layer1_outputs(4383));
    layer2_outputs(2694) <= layer1_outputs(2464);
    layer2_outputs(2695) <= not(layer1_outputs(7213));
    layer2_outputs(2696) <= (layer1_outputs(3458)) or (layer1_outputs(4454));
    layer2_outputs(2697) <= not(layer1_outputs(3439)) or (layer1_outputs(6827));
    layer2_outputs(2698) <= layer1_outputs(5404);
    layer2_outputs(2699) <= (layer1_outputs(3721)) or (layer1_outputs(4755));
    layer2_outputs(2700) <= layer1_outputs(5393);
    layer2_outputs(2701) <= layer1_outputs(3201);
    layer2_outputs(2702) <= layer1_outputs(4672);
    layer2_outputs(2703) <= (layer1_outputs(6236)) and not (layer1_outputs(3392));
    layer2_outputs(2704) <= '1';
    layer2_outputs(2705) <= not(layer1_outputs(6332));
    layer2_outputs(2706) <= (layer1_outputs(2874)) and not (layer1_outputs(5023));
    layer2_outputs(2707) <= not(layer1_outputs(1259));
    layer2_outputs(2708) <= layer1_outputs(3023);
    layer2_outputs(2709) <= not((layer1_outputs(3932)) and (layer1_outputs(4794)));
    layer2_outputs(2710) <= not(layer1_outputs(2254));
    layer2_outputs(2711) <= not((layer1_outputs(3036)) xor (layer1_outputs(6837)));
    layer2_outputs(2712) <= (layer1_outputs(7564)) xor (layer1_outputs(355));
    layer2_outputs(2713) <= not((layer1_outputs(7191)) and (layer1_outputs(3170)));
    layer2_outputs(2714) <= not(layer1_outputs(4583));
    layer2_outputs(2715) <= not(layer1_outputs(509));
    layer2_outputs(2716) <= '0';
    layer2_outputs(2717) <= layer1_outputs(5229);
    layer2_outputs(2718) <= not((layer1_outputs(5480)) or (layer1_outputs(612)));
    layer2_outputs(2719) <= layer1_outputs(690);
    layer2_outputs(2720) <= (layer1_outputs(7443)) and (layer1_outputs(6797));
    layer2_outputs(2721) <= not((layer1_outputs(567)) and (layer1_outputs(70)));
    layer2_outputs(2722) <= not(layer1_outputs(3675)) or (layer1_outputs(6493));
    layer2_outputs(2723) <= layer1_outputs(6312);
    layer2_outputs(2724) <= (layer1_outputs(5157)) or (layer1_outputs(2144));
    layer2_outputs(2725) <= not(layer1_outputs(7119));
    layer2_outputs(2726) <= layer1_outputs(1435);
    layer2_outputs(2727) <= not(layer1_outputs(3400)) or (layer1_outputs(533));
    layer2_outputs(2728) <= (layer1_outputs(1467)) or (layer1_outputs(2129));
    layer2_outputs(2729) <= (layer1_outputs(1819)) or (layer1_outputs(4271));
    layer2_outputs(2730) <= layer1_outputs(3058);
    layer2_outputs(2731) <= not(layer1_outputs(4855)) or (layer1_outputs(2913));
    layer2_outputs(2732) <= not((layer1_outputs(7626)) and (layer1_outputs(5459)));
    layer2_outputs(2733) <= '0';
    layer2_outputs(2734) <= layer1_outputs(2082);
    layer2_outputs(2735) <= '0';
    layer2_outputs(2736) <= not(layer1_outputs(5)) or (layer1_outputs(2387));
    layer2_outputs(2737) <= not((layer1_outputs(532)) or (layer1_outputs(3694)));
    layer2_outputs(2738) <= (layer1_outputs(1886)) or (layer1_outputs(1301));
    layer2_outputs(2739) <= not(layer1_outputs(2560)) or (layer1_outputs(4334));
    layer2_outputs(2740) <= (layer1_outputs(1558)) and not (layer1_outputs(6254));
    layer2_outputs(2741) <= (layer1_outputs(3210)) or (layer1_outputs(5833));
    layer2_outputs(2742) <= (layer1_outputs(561)) and not (layer1_outputs(6431));
    layer2_outputs(2743) <= not(layer1_outputs(6088));
    layer2_outputs(2744) <= layer1_outputs(2675);
    layer2_outputs(2745) <= (layer1_outputs(6588)) or (layer1_outputs(3308));
    layer2_outputs(2746) <= '1';
    layer2_outputs(2747) <= (layer1_outputs(7154)) or (layer1_outputs(7450));
    layer2_outputs(2748) <= layer1_outputs(290);
    layer2_outputs(2749) <= (layer1_outputs(6144)) and not (layer1_outputs(2985));
    layer2_outputs(2750) <= not(layer1_outputs(255)) or (layer1_outputs(5107));
    layer2_outputs(2751) <= not(layer1_outputs(7329));
    layer2_outputs(2752) <= (layer1_outputs(6640)) or (layer1_outputs(5406));
    layer2_outputs(2753) <= not(layer1_outputs(468));
    layer2_outputs(2754) <= (layer1_outputs(4602)) and (layer1_outputs(4544));
    layer2_outputs(2755) <= (layer1_outputs(5740)) and not (layer1_outputs(2938));
    layer2_outputs(2756) <= (layer1_outputs(4887)) and not (layer1_outputs(4422));
    layer2_outputs(2757) <= (layer1_outputs(7636)) and not (layer1_outputs(2514));
    layer2_outputs(2758) <= not(layer1_outputs(5042));
    layer2_outputs(2759) <= not(layer1_outputs(6102));
    layer2_outputs(2760) <= (layer1_outputs(39)) and (layer1_outputs(5672));
    layer2_outputs(2761) <= (layer1_outputs(4530)) xor (layer1_outputs(6981));
    layer2_outputs(2762) <= (layer1_outputs(3730)) and not (layer1_outputs(7551));
    layer2_outputs(2763) <= layer1_outputs(5850);
    layer2_outputs(2764) <= not(layer1_outputs(2980));
    layer2_outputs(2765) <= layer1_outputs(6458);
    layer2_outputs(2766) <= not((layer1_outputs(6828)) or (layer1_outputs(1295)));
    layer2_outputs(2767) <= '1';
    layer2_outputs(2768) <= not(layer1_outputs(111)) or (layer1_outputs(7635));
    layer2_outputs(2769) <= not(layer1_outputs(5451));
    layer2_outputs(2770) <= layer1_outputs(4326);
    layer2_outputs(2771) <= (layer1_outputs(7445)) xor (layer1_outputs(568));
    layer2_outputs(2772) <= not(layer1_outputs(1863)) or (layer1_outputs(3723));
    layer2_outputs(2773) <= not(layer1_outputs(3522));
    layer2_outputs(2774) <= (layer1_outputs(4580)) and not (layer1_outputs(2665));
    layer2_outputs(2775) <= layer1_outputs(1214);
    layer2_outputs(2776) <= not(layer1_outputs(5652)) or (layer1_outputs(4432));
    layer2_outputs(2777) <= not(layer1_outputs(719));
    layer2_outputs(2778) <= not(layer1_outputs(1248));
    layer2_outputs(2779) <= layer1_outputs(4123);
    layer2_outputs(2780) <= not(layer1_outputs(128));
    layer2_outputs(2781) <= '1';
    layer2_outputs(2782) <= not((layer1_outputs(5278)) and (layer1_outputs(6680)));
    layer2_outputs(2783) <= layer1_outputs(1963);
    layer2_outputs(2784) <= not(layer1_outputs(1033)) or (layer1_outputs(4072));
    layer2_outputs(2785) <= not(layer1_outputs(1608)) or (layer1_outputs(3869));
    layer2_outputs(2786) <= (layer1_outputs(1654)) and not (layer1_outputs(4321));
    layer2_outputs(2787) <= (layer1_outputs(6733)) and (layer1_outputs(1178));
    layer2_outputs(2788) <= layer1_outputs(2637);
    layer2_outputs(2789) <= '0';
    layer2_outputs(2790) <= (layer1_outputs(2077)) and not (layer1_outputs(6747));
    layer2_outputs(2791) <= not(layer1_outputs(2721));
    layer2_outputs(2792) <= not((layer1_outputs(2951)) and (layer1_outputs(4619)));
    layer2_outputs(2793) <= (layer1_outputs(6961)) and not (layer1_outputs(1079));
    layer2_outputs(2794) <= (layer1_outputs(6773)) or (layer1_outputs(3377));
    layer2_outputs(2795) <= not(layer1_outputs(3554));
    layer2_outputs(2796) <= not((layer1_outputs(6687)) or (layer1_outputs(4989)));
    layer2_outputs(2797) <= layer1_outputs(5406);
    layer2_outputs(2798) <= '0';
    layer2_outputs(2799) <= not(layer1_outputs(1202)) or (layer1_outputs(3848));
    layer2_outputs(2800) <= not(layer1_outputs(6993)) or (layer1_outputs(5420));
    layer2_outputs(2801) <= (layer1_outputs(534)) xor (layer1_outputs(461));
    layer2_outputs(2802) <= not(layer1_outputs(1310)) or (layer1_outputs(4572));
    layer2_outputs(2803) <= not((layer1_outputs(4246)) and (layer1_outputs(7480)));
    layer2_outputs(2804) <= '1';
    layer2_outputs(2805) <= not((layer1_outputs(5711)) or (layer1_outputs(1154)));
    layer2_outputs(2806) <= layer1_outputs(5715);
    layer2_outputs(2807) <= (layer1_outputs(3349)) and not (layer1_outputs(4356));
    layer2_outputs(2808) <= '0';
    layer2_outputs(2809) <= layer1_outputs(1813);
    layer2_outputs(2810) <= layer1_outputs(6364);
    layer2_outputs(2811) <= (layer1_outputs(7149)) and not (layer1_outputs(5478));
    layer2_outputs(2812) <= (layer1_outputs(6113)) and (layer1_outputs(3511));
    layer2_outputs(2813) <= layer1_outputs(326);
    layer2_outputs(2814) <= layer1_outputs(2876);
    layer2_outputs(2815) <= not(layer1_outputs(2971)) or (layer1_outputs(7648));
    layer2_outputs(2816) <= not((layer1_outputs(6886)) or (layer1_outputs(7089)));
    layer2_outputs(2817) <= not((layer1_outputs(1851)) and (layer1_outputs(3722)));
    layer2_outputs(2818) <= not(layer1_outputs(6160));
    layer2_outputs(2819) <= layer1_outputs(4789);
    layer2_outputs(2820) <= not(layer1_outputs(1962));
    layer2_outputs(2821) <= not(layer1_outputs(1783)) or (layer1_outputs(4084));
    layer2_outputs(2822) <= not(layer1_outputs(3783)) or (layer1_outputs(5921));
    layer2_outputs(2823) <= not((layer1_outputs(225)) or (layer1_outputs(926)));
    layer2_outputs(2824) <= not((layer1_outputs(520)) or (layer1_outputs(3403)));
    layer2_outputs(2825) <= layer1_outputs(2806);
    layer2_outputs(2826) <= '1';
    layer2_outputs(2827) <= not(layer1_outputs(7627)) or (layer1_outputs(2383));
    layer2_outputs(2828) <= not(layer1_outputs(1969));
    layer2_outputs(2829) <= layer1_outputs(1943);
    layer2_outputs(2830) <= not(layer1_outputs(268));
    layer2_outputs(2831) <= not(layer1_outputs(3457));
    layer2_outputs(2832) <= not((layer1_outputs(5661)) and (layer1_outputs(3097)));
    layer2_outputs(2833) <= (layer1_outputs(7185)) and not (layer1_outputs(4933));
    layer2_outputs(2834) <= (layer1_outputs(975)) and (layer1_outputs(1464));
    layer2_outputs(2835) <= not(layer1_outputs(2310));
    layer2_outputs(2836) <= (layer1_outputs(4838)) and not (layer1_outputs(2318));
    layer2_outputs(2837) <= (layer1_outputs(54)) and not (layer1_outputs(2208));
    layer2_outputs(2838) <= not((layer1_outputs(870)) xor (layer1_outputs(3109)));
    layer2_outputs(2839) <= layer1_outputs(5408);
    layer2_outputs(2840) <= not(layer1_outputs(3827)) or (layer1_outputs(3165));
    layer2_outputs(2841) <= (layer1_outputs(566)) and (layer1_outputs(5004));
    layer2_outputs(2842) <= layer1_outputs(218);
    layer2_outputs(2843) <= (layer1_outputs(3907)) or (layer1_outputs(5764));
    layer2_outputs(2844) <= (layer1_outputs(3742)) and not (layer1_outputs(6442));
    layer2_outputs(2845) <= (layer1_outputs(3756)) or (layer1_outputs(3837));
    layer2_outputs(2846) <= not(layer1_outputs(6665)) or (layer1_outputs(3393));
    layer2_outputs(2847) <= layer1_outputs(4829);
    layer2_outputs(2848) <= (layer1_outputs(1796)) and not (layer1_outputs(1308));
    layer2_outputs(2849) <= (layer1_outputs(698)) xor (layer1_outputs(3758));
    layer2_outputs(2850) <= not((layer1_outputs(2412)) xor (layer1_outputs(191)));
    layer2_outputs(2851) <= not(layer1_outputs(2634));
    layer2_outputs(2852) <= not((layer1_outputs(7555)) and (layer1_outputs(1423)));
    layer2_outputs(2853) <= not(layer1_outputs(4323));
    layer2_outputs(2854) <= (layer1_outputs(7507)) or (layer1_outputs(5364));
    layer2_outputs(2855) <= not(layer1_outputs(6187));
    layer2_outputs(2856) <= '1';
    layer2_outputs(2857) <= not(layer1_outputs(1833)) or (layer1_outputs(5368));
    layer2_outputs(2858) <= (layer1_outputs(2066)) and not (layer1_outputs(983));
    layer2_outputs(2859) <= layer1_outputs(5705);
    layer2_outputs(2860) <= not((layer1_outputs(6204)) or (layer1_outputs(3413)));
    layer2_outputs(2861) <= (layer1_outputs(1345)) xor (layer1_outputs(768));
    layer2_outputs(2862) <= not(layer1_outputs(4054)) or (layer1_outputs(5669));
    layer2_outputs(2863) <= not(layer1_outputs(7332)) or (layer1_outputs(7320));
    layer2_outputs(2864) <= (layer1_outputs(91)) and not (layer1_outputs(1800));
    layer2_outputs(2865) <= not(layer1_outputs(19)) or (layer1_outputs(1418));
    layer2_outputs(2866) <= (layer1_outputs(6966)) xor (layer1_outputs(1419));
    layer2_outputs(2867) <= (layer1_outputs(7229)) and (layer1_outputs(2594));
    layer2_outputs(2868) <= layer1_outputs(4608);
    layer2_outputs(2869) <= layer1_outputs(3495);
    layer2_outputs(2870) <= not(layer1_outputs(2737)) or (layer1_outputs(1106));
    layer2_outputs(2871) <= not(layer1_outputs(1192));
    layer2_outputs(2872) <= layer1_outputs(1354);
    layer2_outputs(2873) <= not(layer1_outputs(7269));
    layer2_outputs(2874) <= layer1_outputs(5834);
    layer2_outputs(2875) <= '0';
    layer2_outputs(2876) <= not(layer1_outputs(6896)) or (layer1_outputs(7591));
    layer2_outputs(2877) <= layer1_outputs(4691);
    layer2_outputs(2878) <= not(layer1_outputs(6534)) or (layer1_outputs(3800));
    layer2_outputs(2879) <= (layer1_outputs(6059)) and (layer1_outputs(6422));
    layer2_outputs(2880) <= (layer1_outputs(4069)) and not (layer1_outputs(1253));
    layer2_outputs(2881) <= (layer1_outputs(1259)) and not (layer1_outputs(5975));
    layer2_outputs(2882) <= not((layer1_outputs(358)) and (layer1_outputs(4145)));
    layer2_outputs(2883) <= not(layer1_outputs(1708));
    layer2_outputs(2884) <= not(layer1_outputs(5903));
    layer2_outputs(2885) <= not((layer1_outputs(6940)) and (layer1_outputs(5156)));
    layer2_outputs(2886) <= (layer1_outputs(6844)) and (layer1_outputs(350));
    layer2_outputs(2887) <= not(layer1_outputs(1400)) or (layer1_outputs(1044));
    layer2_outputs(2888) <= '1';
    layer2_outputs(2889) <= layer1_outputs(1518);
    layer2_outputs(2890) <= (layer1_outputs(5904)) xor (layer1_outputs(2248));
    layer2_outputs(2891) <= layer1_outputs(4865);
    layer2_outputs(2892) <= (layer1_outputs(6937)) or (layer1_outputs(3032));
    layer2_outputs(2893) <= not((layer1_outputs(382)) and (layer1_outputs(4070)));
    layer2_outputs(2894) <= layer1_outputs(1866);
    layer2_outputs(2895) <= (layer1_outputs(7202)) or (layer1_outputs(5469));
    layer2_outputs(2896) <= (layer1_outputs(7504)) and not (layer1_outputs(3829));
    layer2_outputs(2897) <= '1';
    layer2_outputs(2898) <= layer1_outputs(4061);
    layer2_outputs(2899) <= layer1_outputs(641);
    layer2_outputs(2900) <= not(layer1_outputs(4764));
    layer2_outputs(2901) <= not(layer1_outputs(2844));
    layer2_outputs(2902) <= layer1_outputs(5956);
    layer2_outputs(2903) <= layer1_outputs(1344);
    layer2_outputs(2904) <= (layer1_outputs(1670)) or (layer1_outputs(5654));
    layer2_outputs(2905) <= not(layer1_outputs(6371));
    layer2_outputs(2906) <= not(layer1_outputs(397));
    layer2_outputs(2907) <= (layer1_outputs(3709)) and not (layer1_outputs(3217));
    layer2_outputs(2908) <= (layer1_outputs(5577)) and not (layer1_outputs(2252));
    layer2_outputs(2909) <= not(layer1_outputs(6682)) or (layer1_outputs(1632));
    layer2_outputs(2910) <= not(layer1_outputs(6764)) or (layer1_outputs(3297));
    layer2_outputs(2911) <= layer1_outputs(7522);
    layer2_outputs(2912) <= not(layer1_outputs(394));
    layer2_outputs(2913) <= not(layer1_outputs(2194)) or (layer1_outputs(3894));
    layer2_outputs(2914) <= not(layer1_outputs(2093));
    layer2_outputs(2915) <= layer1_outputs(1799);
    layer2_outputs(2916) <= not(layer1_outputs(2201));
    layer2_outputs(2917) <= layer1_outputs(492);
    layer2_outputs(2918) <= not((layer1_outputs(3275)) or (layer1_outputs(2163)));
    layer2_outputs(2919) <= layer1_outputs(3456);
    layer2_outputs(2920) <= layer1_outputs(5233);
    layer2_outputs(2921) <= (layer1_outputs(5466)) and not (layer1_outputs(5822));
    layer2_outputs(2922) <= (layer1_outputs(4081)) or (layer1_outputs(5248));
    layer2_outputs(2923) <= layer1_outputs(3073);
    layer2_outputs(2924) <= not(layer1_outputs(998)) or (layer1_outputs(6954));
    layer2_outputs(2925) <= not(layer1_outputs(6723));
    layer2_outputs(2926) <= (layer1_outputs(4403)) or (layer1_outputs(4401));
    layer2_outputs(2927) <= not(layer1_outputs(6370));
    layer2_outputs(2928) <= (layer1_outputs(4943)) or (layer1_outputs(6961));
    layer2_outputs(2929) <= not(layer1_outputs(704));
    layer2_outputs(2930) <= not((layer1_outputs(4856)) xor (layer1_outputs(6098)));
    layer2_outputs(2931) <= not(layer1_outputs(1037));
    layer2_outputs(2932) <= '0';
    layer2_outputs(2933) <= not(layer1_outputs(1333));
    layer2_outputs(2934) <= layer1_outputs(1273);
    layer2_outputs(2935) <= not(layer1_outputs(3268));
    layer2_outputs(2936) <= '1';
    layer2_outputs(2937) <= not(layer1_outputs(6845));
    layer2_outputs(2938) <= layer1_outputs(3297);
    layer2_outputs(2939) <= not(layer1_outputs(1987));
    layer2_outputs(2940) <= layer1_outputs(1391);
    layer2_outputs(2941) <= (layer1_outputs(6656)) and not (layer1_outputs(1294));
    layer2_outputs(2942) <= not(layer1_outputs(2062));
    layer2_outputs(2943) <= layer1_outputs(5209);
    layer2_outputs(2944) <= not((layer1_outputs(6476)) or (layer1_outputs(7336)));
    layer2_outputs(2945) <= layer1_outputs(3513);
    layer2_outputs(2946) <= (layer1_outputs(7138)) and not (layer1_outputs(5766));
    layer2_outputs(2947) <= layer1_outputs(1146);
    layer2_outputs(2948) <= not(layer1_outputs(3542)) or (layer1_outputs(6694));
    layer2_outputs(2949) <= not(layer1_outputs(7137)) or (layer1_outputs(7093));
    layer2_outputs(2950) <= layer1_outputs(5943);
    layer2_outputs(2951) <= (layer1_outputs(7350)) or (layer1_outputs(2063));
    layer2_outputs(2952) <= not(layer1_outputs(5584));
    layer2_outputs(2953) <= (layer1_outputs(544)) or (layer1_outputs(683));
    layer2_outputs(2954) <= layer1_outputs(6148);
    layer2_outputs(2955) <= (layer1_outputs(3298)) and not (layer1_outputs(6141));
    layer2_outputs(2956) <= layer1_outputs(725);
    layer2_outputs(2957) <= not(layer1_outputs(550));
    layer2_outputs(2958) <= not(layer1_outputs(5423)) or (layer1_outputs(7512));
    layer2_outputs(2959) <= (layer1_outputs(3420)) and not (layer1_outputs(1142));
    layer2_outputs(2960) <= not((layer1_outputs(2471)) and (layer1_outputs(4024)));
    layer2_outputs(2961) <= not(layer1_outputs(3921)) or (layer1_outputs(683));
    layer2_outputs(2962) <= not(layer1_outputs(2372)) or (layer1_outputs(7659));
    layer2_outputs(2963) <= layer1_outputs(7155);
    layer2_outputs(2964) <= layer1_outputs(6883);
    layer2_outputs(2965) <= (layer1_outputs(6720)) and (layer1_outputs(5823));
    layer2_outputs(2966) <= not((layer1_outputs(2611)) and (layer1_outputs(3484)));
    layer2_outputs(2967) <= not(layer1_outputs(5146)) or (layer1_outputs(2992));
    layer2_outputs(2968) <= (layer1_outputs(6956)) and (layer1_outputs(640));
    layer2_outputs(2969) <= (layer1_outputs(2679)) and not (layer1_outputs(7669));
    layer2_outputs(2970) <= (layer1_outputs(3889)) and not (layer1_outputs(6409));
    layer2_outputs(2971) <= not(layer1_outputs(4128)) or (layer1_outputs(5659));
    layer2_outputs(2972) <= (layer1_outputs(4036)) and not (layer1_outputs(2344));
    layer2_outputs(2973) <= layer1_outputs(2553);
    layer2_outputs(2974) <= not(layer1_outputs(5077)) or (layer1_outputs(2272));
    layer2_outputs(2975) <= (layer1_outputs(5708)) and (layer1_outputs(1218));
    layer2_outputs(2976) <= layer1_outputs(1978);
    layer2_outputs(2977) <= (layer1_outputs(48)) and not (layer1_outputs(3819));
    layer2_outputs(2978) <= not((layer1_outputs(1617)) or (layer1_outputs(3752)));
    layer2_outputs(2979) <= not((layer1_outputs(4057)) and (layer1_outputs(1363)));
    layer2_outputs(2980) <= '0';
    layer2_outputs(2981) <= (layer1_outputs(5253)) or (layer1_outputs(2150));
    layer2_outputs(2982) <= '1';
    layer2_outputs(2983) <= not((layer1_outputs(6635)) xor (layer1_outputs(335)));
    layer2_outputs(2984) <= layer1_outputs(5202);
    layer2_outputs(2985) <= not((layer1_outputs(1556)) xor (layer1_outputs(6155)));
    layer2_outputs(2986) <= not((layer1_outputs(1075)) and (layer1_outputs(4519)));
    layer2_outputs(2987) <= layer1_outputs(1163);
    layer2_outputs(2988) <= (layer1_outputs(4212)) or (layer1_outputs(2079));
    layer2_outputs(2989) <= (layer1_outputs(1434)) and not (layer1_outputs(2284));
    layer2_outputs(2990) <= not(layer1_outputs(2508)) or (layer1_outputs(6287));
    layer2_outputs(2991) <= '0';
    layer2_outputs(2992) <= not(layer1_outputs(201));
    layer2_outputs(2993) <= layer1_outputs(1556);
    layer2_outputs(2994) <= not((layer1_outputs(6498)) or (layer1_outputs(6607)));
    layer2_outputs(2995) <= '1';
    layer2_outputs(2996) <= (layer1_outputs(7447)) and not (layer1_outputs(4681));
    layer2_outputs(2997) <= (layer1_outputs(7074)) and not (layer1_outputs(2359));
    layer2_outputs(2998) <= not(layer1_outputs(5943)) or (layer1_outputs(5483));
    layer2_outputs(2999) <= (layer1_outputs(4)) xor (layer1_outputs(1544));
    layer2_outputs(3000) <= not(layer1_outputs(714));
    layer2_outputs(3001) <= '1';
    layer2_outputs(3002) <= not(layer1_outputs(861));
    layer2_outputs(3003) <= not((layer1_outputs(831)) and (layer1_outputs(7268)));
    layer2_outputs(3004) <= not(layer1_outputs(6939));
    layer2_outputs(3005) <= not((layer1_outputs(6978)) or (layer1_outputs(6573)));
    layer2_outputs(3006) <= not((layer1_outputs(461)) or (layer1_outputs(5837)));
    layer2_outputs(3007) <= not(layer1_outputs(2911));
    layer2_outputs(3008) <= not(layer1_outputs(1592));
    layer2_outputs(3009) <= not(layer1_outputs(3576));
    layer2_outputs(3010) <= layer1_outputs(3704);
    layer2_outputs(3011) <= '0';
    layer2_outputs(3012) <= (layer1_outputs(1992)) or (layer1_outputs(5819));
    layer2_outputs(3013) <= layer1_outputs(5840);
    layer2_outputs(3014) <= not(layer1_outputs(2757)) or (layer1_outputs(5516));
    layer2_outputs(3015) <= '0';
    layer2_outputs(3016) <= (layer1_outputs(841)) and (layer1_outputs(2439));
    layer2_outputs(3017) <= layer1_outputs(5964);
    layer2_outputs(3018) <= (layer1_outputs(4308)) and (layer1_outputs(4887));
    layer2_outputs(3019) <= not(layer1_outputs(7330));
    layer2_outputs(3020) <= (layer1_outputs(1673)) or (layer1_outputs(2469));
    layer2_outputs(3021) <= not(layer1_outputs(5115)) or (layer1_outputs(1873));
    layer2_outputs(3022) <= layer1_outputs(4759);
    layer2_outputs(3023) <= '1';
    layer2_outputs(3024) <= layer1_outputs(1634);
    layer2_outputs(3025) <= not((layer1_outputs(2390)) and (layer1_outputs(3708)));
    layer2_outputs(3026) <= layer1_outputs(3401);
    layer2_outputs(3027) <= not((layer1_outputs(3950)) or (layer1_outputs(61)));
    layer2_outputs(3028) <= not(layer1_outputs(1715));
    layer2_outputs(3029) <= not((layer1_outputs(1966)) and (layer1_outputs(5352)));
    layer2_outputs(3030) <= not(layer1_outputs(6366)) or (layer1_outputs(5482));
    layer2_outputs(3031) <= not(layer1_outputs(6752));
    layer2_outputs(3032) <= '1';
    layer2_outputs(3033) <= layer1_outputs(5426);
    layer2_outputs(3034) <= not(layer1_outputs(1555)) or (layer1_outputs(4279));
    layer2_outputs(3035) <= '0';
    layer2_outputs(3036) <= (layer1_outputs(4762)) xor (layer1_outputs(3229));
    layer2_outputs(3037) <= not(layer1_outputs(2130)) or (layer1_outputs(2655));
    layer2_outputs(3038) <= (layer1_outputs(7023)) and (layer1_outputs(4223));
    layer2_outputs(3039) <= layer1_outputs(948);
    layer2_outputs(3040) <= not(layer1_outputs(5726));
    layer2_outputs(3041) <= not((layer1_outputs(2178)) and (layer1_outputs(6064)));
    layer2_outputs(3042) <= (layer1_outputs(6276)) and not (layer1_outputs(4647));
    layer2_outputs(3043) <= layer1_outputs(587);
    layer2_outputs(3044) <= not(layer1_outputs(3522));
    layer2_outputs(3045) <= layer1_outputs(5164);
    layer2_outputs(3046) <= '1';
    layer2_outputs(3047) <= '1';
    layer2_outputs(3048) <= '1';
    layer2_outputs(3049) <= not((layer1_outputs(2577)) and (layer1_outputs(1007)));
    layer2_outputs(3050) <= not((layer1_outputs(6557)) and (layer1_outputs(1020)));
    layer2_outputs(3051) <= layer1_outputs(1744);
    layer2_outputs(3052) <= not((layer1_outputs(7112)) and (layer1_outputs(401)));
    layer2_outputs(3053) <= (layer1_outputs(4445)) and (layer1_outputs(2900));
    layer2_outputs(3054) <= (layer1_outputs(5688)) and not (layer1_outputs(5162));
    layer2_outputs(3055) <= (layer1_outputs(4725)) and not (layer1_outputs(2695));
    layer2_outputs(3056) <= not(layer1_outputs(898)) or (layer1_outputs(2220));
    layer2_outputs(3057) <= (layer1_outputs(418)) and not (layer1_outputs(7518));
    layer2_outputs(3058) <= (layer1_outputs(2834)) or (layer1_outputs(4166));
    layer2_outputs(3059) <= (layer1_outputs(2864)) and (layer1_outputs(4981));
    layer2_outputs(3060) <= not((layer1_outputs(1609)) or (layer1_outputs(6136)));
    layer2_outputs(3061) <= not(layer1_outputs(6546));
    layer2_outputs(3062) <= not((layer1_outputs(618)) xor (layer1_outputs(7289)));
    layer2_outputs(3063) <= layer1_outputs(5638);
    layer2_outputs(3064) <= (layer1_outputs(279)) and not (layer1_outputs(5297));
    layer2_outputs(3065) <= not((layer1_outputs(566)) xor (layer1_outputs(6672)));
    layer2_outputs(3066) <= not((layer1_outputs(2445)) or (layer1_outputs(4723)));
    layer2_outputs(3067) <= (layer1_outputs(5277)) and not (layer1_outputs(7118));
    layer2_outputs(3068) <= layer1_outputs(4033);
    layer2_outputs(3069) <= (layer1_outputs(4414)) and not (layer1_outputs(4915));
    layer2_outputs(3070) <= not(layer1_outputs(6764));
    layer2_outputs(3071) <= (layer1_outputs(2953)) and not (layer1_outputs(2857));
    layer2_outputs(3072) <= not(layer1_outputs(1014));
    layer2_outputs(3073) <= (layer1_outputs(6951)) or (layer1_outputs(6657));
    layer2_outputs(3074) <= not(layer1_outputs(3754)) or (layer1_outputs(5058));
    layer2_outputs(3075) <= not(layer1_outputs(4492)) or (layer1_outputs(1536));
    layer2_outputs(3076) <= not((layer1_outputs(3647)) or (layer1_outputs(7412)));
    layer2_outputs(3077) <= layer1_outputs(6440);
    layer2_outputs(3078) <= not(layer1_outputs(2120));
    layer2_outputs(3079) <= layer1_outputs(5242);
    layer2_outputs(3080) <= not((layer1_outputs(968)) or (layer1_outputs(4932)));
    layer2_outputs(3081) <= not(layer1_outputs(635));
    layer2_outputs(3082) <= (layer1_outputs(813)) and not (layer1_outputs(1235));
    layer2_outputs(3083) <= layer1_outputs(7593);
    layer2_outputs(3084) <= not(layer1_outputs(7320)) or (layer1_outputs(3808));
    layer2_outputs(3085) <= not((layer1_outputs(7431)) or (layer1_outputs(6875)));
    layer2_outputs(3086) <= not(layer1_outputs(3287));
    layer2_outputs(3087) <= layer1_outputs(2065);
    layer2_outputs(3088) <= layer1_outputs(4037);
    layer2_outputs(3089) <= not(layer1_outputs(5061)) or (layer1_outputs(4563));
    layer2_outputs(3090) <= '0';
    layer2_outputs(3091) <= not((layer1_outputs(1588)) and (layer1_outputs(4429)));
    layer2_outputs(3092) <= not(layer1_outputs(7589));
    layer2_outputs(3093) <= not(layer1_outputs(414));
    layer2_outputs(3094) <= not(layer1_outputs(6192));
    layer2_outputs(3095) <= (layer1_outputs(6284)) or (layer1_outputs(7386));
    layer2_outputs(3096) <= not(layer1_outputs(491));
    layer2_outputs(3097) <= (layer1_outputs(3255)) and not (layer1_outputs(3352));
    layer2_outputs(3098) <= (layer1_outputs(766)) or (layer1_outputs(1511));
    layer2_outputs(3099) <= (layer1_outputs(4122)) and not (layer1_outputs(3722));
    layer2_outputs(3100) <= not((layer1_outputs(2074)) or (layer1_outputs(4873)));
    layer2_outputs(3101) <= (layer1_outputs(6167)) or (layer1_outputs(4096));
    layer2_outputs(3102) <= (layer1_outputs(5976)) or (layer1_outputs(5488));
    layer2_outputs(3103) <= (layer1_outputs(4989)) and not (layer1_outputs(485));
    layer2_outputs(3104) <= not(layer1_outputs(1621));
    layer2_outputs(3105) <= layer1_outputs(197);
    layer2_outputs(3106) <= not((layer1_outputs(3914)) xor (layer1_outputs(6701)));
    layer2_outputs(3107) <= (layer1_outputs(2531)) and (layer1_outputs(2668));
    layer2_outputs(3108) <= '1';
    layer2_outputs(3109) <= not((layer1_outputs(3925)) xor (layer1_outputs(2786)));
    layer2_outputs(3110) <= (layer1_outputs(3190)) and not (layer1_outputs(5382));
    layer2_outputs(3111) <= (layer1_outputs(6793)) and (layer1_outputs(122));
    layer2_outputs(3112) <= not(layer1_outputs(2907));
    layer2_outputs(3113) <= not(layer1_outputs(3069)) or (layer1_outputs(6346));
    layer2_outputs(3114) <= not(layer1_outputs(4860)) or (layer1_outputs(4120));
    layer2_outputs(3115) <= layer1_outputs(2527);
    layer2_outputs(3116) <= not((layer1_outputs(4624)) and (layer1_outputs(7337)));
    layer2_outputs(3117) <= not(layer1_outputs(5863));
    layer2_outputs(3118) <= not(layer1_outputs(2913)) or (layer1_outputs(7565));
    layer2_outputs(3119) <= '1';
    layer2_outputs(3120) <= layer1_outputs(3645);
    layer2_outputs(3121) <= layer1_outputs(3628);
    layer2_outputs(3122) <= not(layer1_outputs(1777));
    layer2_outputs(3123) <= (layer1_outputs(7446)) xor (layer1_outputs(5735));
    layer2_outputs(3124) <= not(layer1_outputs(448)) or (layer1_outputs(387));
    layer2_outputs(3125) <= (layer1_outputs(1448)) and (layer1_outputs(1750));
    layer2_outputs(3126) <= layer1_outputs(7428);
    layer2_outputs(3127) <= not((layer1_outputs(2662)) xor (layer1_outputs(7111)));
    layer2_outputs(3128) <= (layer1_outputs(7265)) and not (layer1_outputs(3292));
    layer2_outputs(3129) <= not(layer1_outputs(5206));
    layer2_outputs(3130) <= not(layer1_outputs(2629)) or (layer1_outputs(7486));
    layer2_outputs(3131) <= not(layer1_outputs(7314)) or (layer1_outputs(4646));
    layer2_outputs(3132) <= not(layer1_outputs(7531)) or (layer1_outputs(1758));
    layer2_outputs(3133) <= (layer1_outputs(2501)) and not (layer1_outputs(5596));
    layer2_outputs(3134) <= not(layer1_outputs(2606)) or (layer1_outputs(6913));
    layer2_outputs(3135) <= (layer1_outputs(6378)) and not (layer1_outputs(503));
    layer2_outputs(3136) <= not((layer1_outputs(5194)) and (layer1_outputs(6593)));
    layer2_outputs(3137) <= not(layer1_outputs(4232));
    layer2_outputs(3138) <= (layer1_outputs(5843)) or (layer1_outputs(1002));
    layer2_outputs(3139) <= (layer1_outputs(4638)) and not (layer1_outputs(1815));
    layer2_outputs(3140) <= not((layer1_outputs(5649)) and (layer1_outputs(3495)));
    layer2_outputs(3141) <= (layer1_outputs(3218)) and not (layer1_outputs(3397));
    layer2_outputs(3142) <= not((layer1_outputs(3501)) or (layer1_outputs(2277)));
    layer2_outputs(3143) <= not((layer1_outputs(3421)) or (layer1_outputs(7361)));
    layer2_outputs(3144) <= (layer1_outputs(4777)) or (layer1_outputs(5178));
    layer2_outputs(3145) <= (layer1_outputs(4528)) and (layer1_outputs(2109));
    layer2_outputs(3146) <= not((layer1_outputs(7095)) or (layer1_outputs(3445)));
    layer2_outputs(3147) <= '1';
    layer2_outputs(3148) <= not((layer1_outputs(1906)) and (layer1_outputs(2067)));
    layer2_outputs(3149) <= not(layer1_outputs(6903));
    layer2_outputs(3150) <= layer1_outputs(2967);
    layer2_outputs(3151) <= not(layer1_outputs(6225));
    layer2_outputs(3152) <= layer1_outputs(7032);
    layer2_outputs(3153) <= (layer1_outputs(4546)) and (layer1_outputs(1229));
    layer2_outputs(3154) <= not(layer1_outputs(6058));
    layer2_outputs(3155) <= layer1_outputs(3955);
    layer2_outputs(3156) <= layer1_outputs(4101);
    layer2_outputs(3157) <= (layer1_outputs(376)) and not (layer1_outputs(4066));
    layer2_outputs(3158) <= not(layer1_outputs(967));
    layer2_outputs(3159) <= layer1_outputs(665);
    layer2_outputs(3160) <= (layer1_outputs(387)) or (layer1_outputs(585));
    layer2_outputs(3161) <= not(layer1_outputs(2245));
    layer2_outputs(3162) <= (layer1_outputs(5948)) or (layer1_outputs(7340));
    layer2_outputs(3163) <= not((layer1_outputs(5045)) or (layer1_outputs(7140)));
    layer2_outputs(3164) <= layer1_outputs(5823);
    layer2_outputs(3165) <= not(layer1_outputs(1110)) or (layer1_outputs(7642));
    layer2_outputs(3166) <= not(layer1_outputs(6665));
    layer2_outputs(3167) <= not((layer1_outputs(999)) and (layer1_outputs(6643)));
    layer2_outputs(3168) <= not(layer1_outputs(3403));
    layer2_outputs(3169) <= layer1_outputs(7070);
    layer2_outputs(3170) <= layer1_outputs(7219);
    layer2_outputs(3171) <= layer1_outputs(7022);
    layer2_outputs(3172) <= not(layer1_outputs(5765));
    layer2_outputs(3173) <= '1';
    layer2_outputs(3174) <= not(layer1_outputs(7557));
    layer2_outputs(3175) <= (layer1_outputs(949)) or (layer1_outputs(5415));
    layer2_outputs(3176) <= not((layer1_outputs(4566)) or (layer1_outputs(6260)));
    layer2_outputs(3177) <= (layer1_outputs(1734)) and not (layer1_outputs(3253));
    layer2_outputs(3178) <= (layer1_outputs(416)) and not (layer1_outputs(7539));
    layer2_outputs(3179) <= (layer1_outputs(5648)) and not (layer1_outputs(7549));
    layer2_outputs(3180) <= layer1_outputs(7121);
    layer2_outputs(3181) <= not(layer1_outputs(625));
    layer2_outputs(3182) <= layer1_outputs(1070);
    layer2_outputs(3183) <= not(layer1_outputs(6794));
    layer2_outputs(3184) <= (layer1_outputs(1749)) and (layer1_outputs(2494));
    layer2_outputs(3185) <= layer1_outputs(7546);
    layer2_outputs(3186) <= not((layer1_outputs(5372)) or (layer1_outputs(311)));
    layer2_outputs(3187) <= layer1_outputs(2047);
    layer2_outputs(3188) <= layer1_outputs(6363);
    layer2_outputs(3189) <= (layer1_outputs(2328)) and (layer1_outputs(6497));
    layer2_outputs(3190) <= (layer1_outputs(1818)) or (layer1_outputs(4609));
    layer2_outputs(3191) <= layer1_outputs(7481);
    layer2_outputs(3192) <= layer1_outputs(7305);
    layer2_outputs(3193) <= not(layer1_outputs(6153));
    layer2_outputs(3194) <= not((layer1_outputs(2204)) and (layer1_outputs(1115)));
    layer2_outputs(3195) <= not(layer1_outputs(5021)) or (layer1_outputs(6555));
    layer2_outputs(3196) <= (layer1_outputs(39)) and not (layer1_outputs(4115));
    layer2_outputs(3197) <= not(layer1_outputs(2535));
    layer2_outputs(3198) <= not((layer1_outputs(995)) and (layer1_outputs(6311)));
    layer2_outputs(3199) <= not(layer1_outputs(2491));
    layer2_outputs(3200) <= (layer1_outputs(6661)) and not (layer1_outputs(5403));
    layer2_outputs(3201) <= layer1_outputs(6870);
    layer2_outputs(3202) <= not(layer1_outputs(3062));
    layer2_outputs(3203) <= (layer1_outputs(5921)) or (layer1_outputs(6263));
    layer2_outputs(3204) <= not(layer1_outputs(4699)) or (layer1_outputs(5798));
    layer2_outputs(3205) <= '1';
    layer2_outputs(3206) <= not(layer1_outputs(1138));
    layer2_outputs(3207) <= (layer1_outputs(5013)) and (layer1_outputs(494));
    layer2_outputs(3208) <= not(layer1_outputs(5930)) or (layer1_outputs(924));
    layer2_outputs(3209) <= '1';
    layer2_outputs(3210) <= not(layer1_outputs(709));
    layer2_outputs(3211) <= layer1_outputs(2511);
    layer2_outputs(3212) <= (layer1_outputs(1610)) and not (layer1_outputs(800));
    layer2_outputs(3213) <= (layer1_outputs(3205)) xor (layer1_outputs(2641));
    layer2_outputs(3214) <= not(layer1_outputs(4160));
    layer2_outputs(3215) <= not(layer1_outputs(587));
    layer2_outputs(3216) <= not(layer1_outputs(5000)) or (layer1_outputs(2164));
    layer2_outputs(3217) <= (layer1_outputs(7274)) and (layer1_outputs(4264));
    layer2_outputs(3218) <= (layer1_outputs(1078)) or (layer1_outputs(3962));
    layer2_outputs(3219) <= not((layer1_outputs(7418)) or (layer1_outputs(6631)));
    layer2_outputs(3220) <= (layer1_outputs(5023)) and (layer1_outputs(2802));
    layer2_outputs(3221) <= (layer1_outputs(1850)) and (layer1_outputs(5641));
    layer2_outputs(3222) <= (layer1_outputs(1309)) and (layer1_outputs(1680));
    layer2_outputs(3223) <= (layer1_outputs(1306)) or (layer1_outputs(5856));
    layer2_outputs(3224) <= not(layer1_outputs(2599)) or (layer1_outputs(7039));
    layer2_outputs(3225) <= '1';
    layer2_outputs(3226) <= (layer1_outputs(6920)) and not (layer1_outputs(2330));
    layer2_outputs(3227) <= not(layer1_outputs(6897)) or (layer1_outputs(3370));
    layer2_outputs(3228) <= not(layer1_outputs(1216));
    layer2_outputs(3229) <= layer1_outputs(120);
    layer2_outputs(3230) <= '1';
    layer2_outputs(3231) <= '0';
    layer2_outputs(3232) <= (layer1_outputs(7001)) xor (layer1_outputs(5418));
    layer2_outputs(3233) <= (layer1_outputs(723)) or (layer1_outputs(3954));
    layer2_outputs(3234) <= layer1_outputs(3609);
    layer2_outputs(3235) <= (layer1_outputs(2430)) and not (layer1_outputs(344));
    layer2_outputs(3236) <= not(layer1_outputs(5026)) or (layer1_outputs(1090));
    layer2_outputs(3237) <= (layer1_outputs(680)) and not (layer1_outputs(6109));
    layer2_outputs(3238) <= not(layer1_outputs(6128));
    layer2_outputs(3239) <= not(layer1_outputs(1840)) or (layer1_outputs(4871));
    layer2_outputs(3240) <= layer1_outputs(954);
    layer2_outputs(3241) <= layer1_outputs(4815);
    layer2_outputs(3242) <= not((layer1_outputs(5403)) xor (layer1_outputs(4525)));
    layer2_outputs(3243) <= not((layer1_outputs(5790)) or (layer1_outputs(7391)));
    layer2_outputs(3244) <= layer1_outputs(5977);
    layer2_outputs(3245) <= not((layer1_outputs(2701)) xor (layer1_outputs(254)));
    layer2_outputs(3246) <= (layer1_outputs(2131)) or (layer1_outputs(2784));
    layer2_outputs(3247) <= (layer1_outputs(2472)) xor (layer1_outputs(5530));
    layer2_outputs(3248) <= layer1_outputs(5896);
    layer2_outputs(3249) <= not(layer1_outputs(2504)) or (layer1_outputs(7625));
    layer2_outputs(3250) <= not((layer1_outputs(6)) or (layer1_outputs(798)));
    layer2_outputs(3251) <= not(layer1_outputs(7290));
    layer2_outputs(3252) <= not(layer1_outputs(6635)) or (layer1_outputs(1008));
    layer2_outputs(3253) <= (layer1_outputs(3548)) and not (layer1_outputs(515));
    layer2_outputs(3254) <= (layer1_outputs(4391)) or (layer1_outputs(3));
    layer2_outputs(3255) <= (layer1_outputs(151)) and not (layer1_outputs(7500));
    layer2_outputs(3256) <= not(layer1_outputs(4291));
    layer2_outputs(3257) <= '0';
    layer2_outputs(3258) <= not(layer1_outputs(2688));
    layer2_outputs(3259) <= not((layer1_outputs(7286)) and (layer1_outputs(1990)));
    layer2_outputs(3260) <= not((layer1_outputs(5268)) or (layer1_outputs(4712)));
    layer2_outputs(3261) <= (layer1_outputs(4348)) or (layer1_outputs(3266));
    layer2_outputs(3262) <= not(layer1_outputs(320));
    layer2_outputs(3263) <= not(layer1_outputs(3311));
    layer2_outputs(3264) <= layer1_outputs(1067);
    layer2_outputs(3265) <= not(layer1_outputs(7661)) or (layer1_outputs(1218));
    layer2_outputs(3266) <= not(layer1_outputs(5417));
    layer2_outputs(3267) <= layer1_outputs(3810);
    layer2_outputs(3268) <= not(layer1_outputs(3330));
    layer2_outputs(3269) <= not(layer1_outputs(6817));
    layer2_outputs(3270) <= layer1_outputs(6794);
    layer2_outputs(3271) <= not(layer1_outputs(6520));
    layer2_outputs(3272) <= layer1_outputs(2409);
    layer2_outputs(3273) <= not((layer1_outputs(475)) or (layer1_outputs(3739)));
    layer2_outputs(3274) <= (layer1_outputs(6801)) or (layer1_outputs(3675));
    layer2_outputs(3275) <= not(layer1_outputs(2662));
    layer2_outputs(3276) <= not(layer1_outputs(4471));
    layer2_outputs(3277) <= not(layer1_outputs(2159));
    layer2_outputs(3278) <= layer1_outputs(875);
    layer2_outputs(3279) <= (layer1_outputs(4622)) and not (layer1_outputs(3356));
    layer2_outputs(3280) <= layer1_outputs(484);
    layer2_outputs(3281) <= not((layer1_outputs(1432)) and (layer1_outputs(5265)));
    layer2_outputs(3282) <= not(layer1_outputs(3151));
    layer2_outputs(3283) <= (layer1_outputs(7677)) and (layer1_outputs(3407));
    layer2_outputs(3284) <= not(layer1_outputs(6739)) or (layer1_outputs(4874));
    layer2_outputs(3285) <= layer1_outputs(4984);
    layer2_outputs(3286) <= not(layer1_outputs(6939));
    layer2_outputs(3287) <= not((layer1_outputs(4114)) or (layer1_outputs(7590)));
    layer2_outputs(3288) <= not((layer1_outputs(6618)) xor (layer1_outputs(4218)));
    layer2_outputs(3289) <= not((layer1_outputs(1439)) and (layer1_outputs(3267)));
    layer2_outputs(3290) <= (layer1_outputs(2723)) and not (layer1_outputs(5728));
    layer2_outputs(3291) <= not(layer1_outputs(200));
    layer2_outputs(3292) <= not(layer1_outputs(2368));
    layer2_outputs(3293) <= not(layer1_outputs(232)) or (layer1_outputs(6869));
    layer2_outputs(3294) <= not((layer1_outputs(7297)) or (layer1_outputs(1330)));
    layer2_outputs(3295) <= '1';
    layer2_outputs(3296) <= '1';
    layer2_outputs(3297) <= '0';
    layer2_outputs(3298) <= layer1_outputs(6804);
    layer2_outputs(3299) <= (layer1_outputs(4704)) and not (layer1_outputs(2141));
    layer2_outputs(3300) <= layer1_outputs(6952);
    layer2_outputs(3301) <= not(layer1_outputs(4564));
    layer2_outputs(3302) <= layer1_outputs(7051);
    layer2_outputs(3303) <= not((layer1_outputs(648)) xor (layer1_outputs(1630)));
    layer2_outputs(3304) <= layer1_outputs(1406);
    layer2_outputs(3305) <= layer1_outputs(732);
    layer2_outputs(3306) <= not(layer1_outputs(1083)) or (layer1_outputs(1586));
    layer2_outputs(3307) <= (layer1_outputs(7570)) and not (layer1_outputs(4645));
    layer2_outputs(3308) <= layer1_outputs(2154);
    layer2_outputs(3309) <= (layer1_outputs(1275)) xor (layer1_outputs(6508));
    layer2_outputs(3310) <= '1';
    layer2_outputs(3311) <= layer1_outputs(2382);
    layer2_outputs(3312) <= (layer1_outputs(710)) or (layer1_outputs(5502));
    layer2_outputs(3313) <= (layer1_outputs(7280)) and (layer1_outputs(4517));
    layer2_outputs(3314) <= not(layer1_outputs(3025));
    layer2_outputs(3315) <= not(layer1_outputs(6163));
    layer2_outputs(3316) <= (layer1_outputs(3947)) and not (layer1_outputs(783));
    layer2_outputs(3317) <= layer1_outputs(2158);
    layer2_outputs(3318) <= not(layer1_outputs(377));
    layer2_outputs(3319) <= '1';
    layer2_outputs(3320) <= (layer1_outputs(2649)) or (layer1_outputs(7475));
    layer2_outputs(3321) <= not((layer1_outputs(1390)) and (layer1_outputs(6992)));
    layer2_outputs(3322) <= not(layer1_outputs(2110)) or (layer1_outputs(1297));
    layer2_outputs(3323) <= layer1_outputs(1629);
    layer2_outputs(3324) <= layer1_outputs(71);
    layer2_outputs(3325) <= '1';
    layer2_outputs(3326) <= not(layer1_outputs(2899));
    layer2_outputs(3327) <= not((layer1_outputs(943)) or (layer1_outputs(737)));
    layer2_outputs(3328) <= (layer1_outputs(460)) and not (layer1_outputs(4941));
    layer2_outputs(3329) <= not(layer1_outputs(4034));
    layer2_outputs(3330) <= not(layer1_outputs(5568));
    layer2_outputs(3331) <= (layer1_outputs(1485)) or (layer1_outputs(7471));
    layer2_outputs(3332) <= not((layer1_outputs(3413)) and (layer1_outputs(3251)));
    layer2_outputs(3333) <= (layer1_outputs(903)) and not (layer1_outputs(5346));
    layer2_outputs(3334) <= not(layer1_outputs(4537));
    layer2_outputs(3335) <= not(layer1_outputs(4715));
    layer2_outputs(3336) <= layer1_outputs(5576);
    layer2_outputs(3337) <= not(layer1_outputs(3528));
    layer2_outputs(3338) <= not(layer1_outputs(7304));
    layer2_outputs(3339) <= not(layer1_outputs(981));
    layer2_outputs(3340) <= not(layer1_outputs(518));
    layer2_outputs(3341) <= (layer1_outputs(2718)) and (layer1_outputs(7453));
    layer2_outputs(3342) <= (layer1_outputs(5450)) and (layer1_outputs(4335));
    layer2_outputs(3343) <= layer1_outputs(7200);
    layer2_outputs(3344) <= not((layer1_outputs(2606)) or (layer1_outputs(4219)));
    layer2_outputs(3345) <= (layer1_outputs(6755)) or (layer1_outputs(3226));
    layer2_outputs(3346) <= layer1_outputs(4966);
    layer2_outputs(3347) <= not(layer1_outputs(330));
    layer2_outputs(3348) <= layer1_outputs(5841);
    layer2_outputs(3349) <= not((layer1_outputs(31)) or (layer1_outputs(4786)));
    layer2_outputs(3350) <= layer1_outputs(1248);
    layer2_outputs(3351) <= not(layer1_outputs(1849));
    layer2_outputs(3352) <= not(layer1_outputs(6479));
    layer2_outputs(3353) <= not(layer1_outputs(2787));
    layer2_outputs(3354) <= not(layer1_outputs(3967));
    layer2_outputs(3355) <= layer1_outputs(1068);
    layer2_outputs(3356) <= not((layer1_outputs(4550)) or (layer1_outputs(3161)));
    layer2_outputs(3357) <= not(layer1_outputs(4141));
    layer2_outputs(3358) <= not(layer1_outputs(5321)) or (layer1_outputs(303));
    layer2_outputs(3359) <= (layer1_outputs(4450)) and (layer1_outputs(7592));
    layer2_outputs(3360) <= (layer1_outputs(1791)) and not (layer1_outputs(2634));
    layer2_outputs(3361) <= '0';
    layer2_outputs(3362) <= not(layer1_outputs(3989));
    layer2_outputs(3363) <= (layer1_outputs(6286)) and not (layer1_outputs(6877));
    layer2_outputs(3364) <= not((layer1_outputs(4908)) and (layer1_outputs(4521)));
    layer2_outputs(3365) <= '1';
    layer2_outputs(3366) <= not(layer1_outputs(5565)) or (layer1_outputs(2030));
    layer2_outputs(3367) <= '0';
    layer2_outputs(3368) <= layer1_outputs(2438);
    layer2_outputs(3369) <= (layer1_outputs(1113)) and (layer1_outputs(1632));
    layer2_outputs(3370) <= not(layer1_outputs(6068));
    layer2_outputs(3371) <= not(layer1_outputs(3693));
    layer2_outputs(3372) <= not((layer1_outputs(6539)) or (layer1_outputs(3024)));
    layer2_outputs(3373) <= layer1_outputs(7563);
    layer2_outputs(3374) <= (layer1_outputs(6508)) and (layer1_outputs(7452));
    layer2_outputs(3375) <= not(layer1_outputs(405)) or (layer1_outputs(6745));
    layer2_outputs(3376) <= not((layer1_outputs(7560)) and (layer1_outputs(2699)));
    layer2_outputs(3377) <= not(layer1_outputs(7024)) or (layer1_outputs(1054));
    layer2_outputs(3378) <= '1';
    layer2_outputs(3379) <= (layer1_outputs(453)) or (layer1_outputs(5322));
    layer2_outputs(3380) <= (layer1_outputs(6145)) and not (layer1_outputs(7224));
    layer2_outputs(3381) <= not(layer1_outputs(4410));
    layer2_outputs(3382) <= layer1_outputs(3);
    layer2_outputs(3383) <= not(layer1_outputs(6218));
    layer2_outputs(3384) <= '0';
    layer2_outputs(3385) <= not(layer1_outputs(6170)) or (layer1_outputs(4795));
    layer2_outputs(3386) <= (layer1_outputs(4627)) or (layer1_outputs(6813));
    layer2_outputs(3387) <= not((layer1_outputs(3016)) or (layer1_outputs(5679)));
    layer2_outputs(3388) <= '0';
    layer2_outputs(3389) <= (layer1_outputs(2154)) and (layer1_outputs(5731));
    layer2_outputs(3390) <= (layer1_outputs(6847)) and (layer1_outputs(2839));
    layer2_outputs(3391) <= not((layer1_outputs(403)) and (layer1_outputs(2429)));
    layer2_outputs(3392) <= not(layer1_outputs(2552)) or (layer1_outputs(7211));
    layer2_outputs(3393) <= not((layer1_outputs(7655)) or (layer1_outputs(1601)));
    layer2_outputs(3394) <= not((layer1_outputs(4904)) xor (layer1_outputs(327)));
    layer2_outputs(3395) <= '1';
    layer2_outputs(3396) <= not(layer1_outputs(4987));
    layer2_outputs(3397) <= not(layer1_outputs(6960)) or (layer1_outputs(6871));
    layer2_outputs(3398) <= not(layer1_outputs(1367));
    layer2_outputs(3399) <= not((layer1_outputs(5645)) or (layer1_outputs(2700)));
    layer2_outputs(3400) <= not(layer1_outputs(274)) or (layer1_outputs(1204));
    layer2_outputs(3401) <= not(layer1_outputs(50));
    layer2_outputs(3402) <= (layer1_outputs(3968)) and not (layer1_outputs(6769));
    layer2_outputs(3403) <= layer1_outputs(131);
    layer2_outputs(3404) <= (layer1_outputs(2716)) or (layer1_outputs(6333));
    layer2_outputs(3405) <= (layer1_outputs(6008)) and not (layer1_outputs(6766));
    layer2_outputs(3406) <= (layer1_outputs(7310)) and not (layer1_outputs(5709));
    layer2_outputs(3407) <= not(layer1_outputs(286));
    layer2_outputs(3408) <= (layer1_outputs(3633)) or (layer1_outputs(7299));
    layer2_outputs(3409) <= layer1_outputs(7098);
    layer2_outputs(3410) <= not(layer1_outputs(5394));
    layer2_outputs(3411) <= not(layer1_outputs(5236)) or (layer1_outputs(1387));
    layer2_outputs(3412) <= not(layer1_outputs(5022));
    layer2_outputs(3413) <= not((layer1_outputs(2075)) and (layer1_outputs(204)));
    layer2_outputs(3414) <= not(layer1_outputs(2629)) or (layer1_outputs(3532));
    layer2_outputs(3415) <= not(layer1_outputs(3325)) or (layer1_outputs(1688));
    layer2_outputs(3416) <= (layer1_outputs(4353)) and not (layer1_outputs(3904));
    layer2_outputs(3417) <= (layer1_outputs(2144)) and (layer1_outputs(3832));
    layer2_outputs(3418) <= not(layer1_outputs(5894));
    layer2_outputs(3419) <= layer1_outputs(3749);
    layer2_outputs(3420) <= not(layer1_outputs(2863)) or (layer1_outputs(5479));
    layer2_outputs(3421) <= not(layer1_outputs(459)) or (layer1_outputs(920));
    layer2_outputs(3422) <= not((layer1_outputs(3290)) and (layer1_outputs(6532)));
    layer2_outputs(3423) <= not((layer1_outputs(2263)) xor (layer1_outputs(5841)));
    layer2_outputs(3424) <= not((layer1_outputs(5909)) and (layer1_outputs(4820)));
    layer2_outputs(3425) <= layer1_outputs(4224);
    layer2_outputs(3426) <= not(layer1_outputs(3655));
    layer2_outputs(3427) <= (layer1_outputs(7424)) or (layer1_outputs(6161));
    layer2_outputs(3428) <= (layer1_outputs(6277)) and not (layer1_outputs(6688));
    layer2_outputs(3429) <= not(layer1_outputs(281));
    layer2_outputs(3430) <= layer1_outputs(5734);
    layer2_outputs(3431) <= layer1_outputs(1682);
    layer2_outputs(3432) <= not(layer1_outputs(4532));
    layer2_outputs(3433) <= not(layer1_outputs(3791));
    layer2_outputs(3434) <= not((layer1_outputs(4527)) or (layer1_outputs(3222)));
    layer2_outputs(3435) <= layer1_outputs(3779);
    layer2_outputs(3436) <= not((layer1_outputs(3369)) and (layer1_outputs(2094)));
    layer2_outputs(3437) <= not(layer1_outputs(900));
    layer2_outputs(3438) <= layer1_outputs(2633);
    layer2_outputs(3439) <= not((layer1_outputs(715)) or (layer1_outputs(2310)));
    layer2_outputs(3440) <= not(layer1_outputs(5279));
    layer2_outputs(3441) <= (layer1_outputs(3156)) and not (layer1_outputs(3139));
    layer2_outputs(3442) <= '1';
    layer2_outputs(3443) <= layer1_outputs(5849);
    layer2_outputs(3444) <= not(layer1_outputs(1869));
    layer2_outputs(3445) <= not(layer1_outputs(2393));
    layer2_outputs(3446) <= not(layer1_outputs(1656));
    layer2_outputs(3447) <= not(layer1_outputs(420));
    layer2_outputs(3448) <= (layer1_outputs(5235)) and not (layer1_outputs(2421));
    layer2_outputs(3449) <= not(layer1_outputs(5266));
    layer2_outputs(3450) <= layer1_outputs(372);
    layer2_outputs(3451) <= not((layer1_outputs(3972)) or (layer1_outputs(3290)));
    layer2_outputs(3452) <= layer1_outputs(756);
    layer2_outputs(3453) <= layer1_outputs(356);
    layer2_outputs(3454) <= (layer1_outputs(488)) and not (layer1_outputs(7387));
    layer2_outputs(3455) <= not(layer1_outputs(2437)) or (layer1_outputs(1015));
    layer2_outputs(3456) <= not(layer1_outputs(7194));
    layer2_outputs(3457) <= (layer1_outputs(4961)) and not (layer1_outputs(5113));
    layer2_outputs(3458) <= (layer1_outputs(6732)) and not (layer1_outputs(7028));
    layer2_outputs(3459) <= layer1_outputs(7069);
    layer2_outputs(3460) <= (layer1_outputs(3599)) and not (layer1_outputs(2856));
    layer2_outputs(3461) <= (layer1_outputs(7601)) xor (layer1_outputs(5331));
    layer2_outputs(3462) <= not(layer1_outputs(86)) or (layer1_outputs(3410));
    layer2_outputs(3463) <= (layer1_outputs(5923)) xor (layer1_outputs(1639));
    layer2_outputs(3464) <= (layer1_outputs(3642)) and not (layer1_outputs(1641));
    layer2_outputs(3465) <= (layer1_outputs(1967)) and not (layer1_outputs(624));
    layer2_outputs(3466) <= not(layer1_outputs(1930)) or (layer1_outputs(4118));
    layer2_outputs(3467) <= not((layer1_outputs(6686)) and (layer1_outputs(5880)));
    layer2_outputs(3468) <= not(layer1_outputs(2364)) or (layer1_outputs(4217));
    layer2_outputs(3469) <= not(layer1_outputs(4704));
    layer2_outputs(3470) <= layer1_outputs(1538);
    layer2_outputs(3471) <= not(layer1_outputs(939)) or (layer1_outputs(282));
    layer2_outputs(3472) <= layer1_outputs(2704);
    layer2_outputs(3473) <= '0';
    layer2_outputs(3474) <= '0';
    layer2_outputs(3475) <= (layer1_outputs(5697)) or (layer1_outputs(4021));
    layer2_outputs(3476) <= layer1_outputs(399);
    layer2_outputs(3477) <= layer1_outputs(1866);
    layer2_outputs(3478) <= layer1_outputs(241);
    layer2_outputs(3479) <= not(layer1_outputs(3868));
    layer2_outputs(3480) <= not(layer1_outputs(2219)) or (layer1_outputs(1832));
    layer2_outputs(3481) <= layer1_outputs(1681);
    layer2_outputs(3482) <= (layer1_outputs(1255)) and (layer1_outputs(6221));
    layer2_outputs(3483) <= not(layer1_outputs(1811)) or (layer1_outputs(2994));
    layer2_outputs(3484) <= not((layer1_outputs(5383)) and (layer1_outputs(1574)));
    layer2_outputs(3485) <= layer1_outputs(5060);
    layer2_outputs(3486) <= not(layer1_outputs(5994)) or (layer1_outputs(279));
    layer2_outputs(3487) <= not(layer1_outputs(645));
    layer2_outputs(3488) <= '1';
    layer2_outputs(3489) <= (layer1_outputs(5330)) and not (layer1_outputs(2944));
    layer2_outputs(3490) <= layer1_outputs(2497);
    layer2_outputs(3491) <= not(layer1_outputs(5015));
    layer2_outputs(3492) <= not(layer1_outputs(7553)) or (layer1_outputs(4125));
    layer2_outputs(3493) <= layer1_outputs(1547);
    layer2_outputs(3494) <= not(layer1_outputs(1260)) or (layer1_outputs(4524));
    layer2_outputs(3495) <= layer1_outputs(758);
    layer2_outputs(3496) <= not(layer1_outputs(5189));
    layer2_outputs(3497) <= (layer1_outputs(3716)) and not (layer1_outputs(7222));
    layer2_outputs(3498) <= not((layer1_outputs(6173)) or (layer1_outputs(3784)));
    layer2_outputs(3499) <= (layer1_outputs(2136)) and not (layer1_outputs(6074));
    layer2_outputs(3500) <= '1';
    layer2_outputs(3501) <= not((layer1_outputs(5055)) and (layer1_outputs(5544)));
    layer2_outputs(3502) <= (layer1_outputs(3236)) and not (layer1_outputs(496));
    layer2_outputs(3503) <= layer1_outputs(4993);
    layer2_outputs(3504) <= not(layer1_outputs(1528));
    layer2_outputs(3505) <= not((layer1_outputs(1918)) and (layer1_outputs(4808)));
    layer2_outputs(3506) <= '0';
    layer2_outputs(3507) <= layer1_outputs(334);
    layer2_outputs(3508) <= (layer1_outputs(5576)) and not (layer1_outputs(916));
    layer2_outputs(3509) <= (layer1_outputs(1662)) and (layer1_outputs(1091));
    layer2_outputs(3510) <= not((layer1_outputs(2099)) and (layer1_outputs(4894)));
    layer2_outputs(3511) <= layer1_outputs(957);
    layer2_outputs(3512) <= '0';
    layer2_outputs(3513) <= layer1_outputs(948);
    layer2_outputs(3514) <= layer1_outputs(850);
    layer2_outputs(3515) <= not(layer1_outputs(7604));
    layer2_outputs(3516) <= not((layer1_outputs(719)) or (layer1_outputs(2146)));
    layer2_outputs(3517) <= layer1_outputs(198);
    layer2_outputs(3518) <= not(layer1_outputs(875));
    layer2_outputs(3519) <= layer1_outputs(283);
    layer2_outputs(3520) <= (layer1_outputs(5021)) or (layer1_outputs(5294));
    layer2_outputs(3521) <= (layer1_outputs(3483)) xor (layer1_outputs(4441));
    layer2_outputs(3522) <= not(layer1_outputs(2181)) or (layer1_outputs(7606));
    layer2_outputs(3523) <= layer1_outputs(1922);
    layer2_outputs(3524) <= layer1_outputs(2648);
    layer2_outputs(3525) <= not(layer1_outputs(5466));
    layer2_outputs(3526) <= (layer1_outputs(5357)) and not (layer1_outputs(7544));
    layer2_outputs(3527) <= (layer1_outputs(4462)) xor (layer1_outputs(5751));
    layer2_outputs(3528) <= layer1_outputs(3389);
    layer2_outputs(3529) <= (layer1_outputs(4064)) and (layer1_outputs(6015));
    layer2_outputs(3530) <= not(layer1_outputs(3355));
    layer2_outputs(3531) <= not(layer1_outputs(104));
    layer2_outputs(3532) <= not((layer1_outputs(5639)) or (layer1_outputs(3291)));
    layer2_outputs(3533) <= not(layer1_outputs(6821));
    layer2_outputs(3534) <= (layer1_outputs(2358)) or (layer1_outputs(7273));
    layer2_outputs(3535) <= not((layer1_outputs(3288)) or (layer1_outputs(3437)));
    layer2_outputs(3536) <= not((layer1_outputs(5280)) or (layer1_outputs(4157)));
    layer2_outputs(3537) <= (layer1_outputs(199)) xor (layer1_outputs(2824));
    layer2_outputs(3538) <= not((layer1_outputs(2706)) and (layer1_outputs(3652)));
    layer2_outputs(3539) <= not(layer1_outputs(113));
    layer2_outputs(3540) <= not((layer1_outputs(7612)) and (layer1_outputs(2028)));
    layer2_outputs(3541) <= not(layer1_outputs(6023));
    layer2_outputs(3542) <= (layer1_outputs(7138)) and (layer1_outputs(937));
    layer2_outputs(3543) <= (layer1_outputs(2230)) or (layer1_outputs(4953));
    layer2_outputs(3544) <= '1';
    layer2_outputs(3545) <= not((layer1_outputs(729)) xor (layer1_outputs(1942)));
    layer2_outputs(3546) <= (layer1_outputs(1313)) or (layer1_outputs(6822));
    layer2_outputs(3547) <= layer1_outputs(1092);
    layer2_outputs(3548) <= not(layer1_outputs(2560));
    layer2_outputs(3549) <= not((layer1_outputs(6925)) and (layer1_outputs(2529)));
    layer2_outputs(3550) <= not(layer1_outputs(3238));
    layer2_outputs(3551) <= (layer1_outputs(1835)) or (layer1_outputs(6433));
    layer2_outputs(3552) <= '1';
    layer2_outputs(3553) <= (layer1_outputs(5177)) or (layer1_outputs(6414));
    layer2_outputs(3554) <= (layer1_outputs(5338)) and (layer1_outputs(2428));
    layer2_outputs(3555) <= not(layer1_outputs(4412));
    layer2_outputs(3556) <= (layer1_outputs(1266)) or (layer1_outputs(2156));
    layer2_outputs(3557) <= layer1_outputs(4393);
    layer2_outputs(3558) <= not(layer1_outputs(4711));
    layer2_outputs(3559) <= layer1_outputs(1845);
    layer2_outputs(3560) <= layer1_outputs(6880);
    layer2_outputs(3561) <= layer1_outputs(2527);
    layer2_outputs(3562) <= not((layer1_outputs(4153)) or (layer1_outputs(6156)));
    layer2_outputs(3563) <= not((layer1_outputs(5485)) or (layer1_outputs(4511)));
    layer2_outputs(3564) <= layer1_outputs(2450);
    layer2_outputs(3565) <= not(layer1_outputs(3678));
    layer2_outputs(3566) <= not(layer1_outputs(4024)) or (layer1_outputs(929));
    layer2_outputs(3567) <= not((layer1_outputs(4811)) or (layer1_outputs(1220)));
    layer2_outputs(3568) <= not(layer1_outputs(5627)) or (layer1_outputs(3059));
    layer2_outputs(3569) <= (layer1_outputs(3225)) or (layer1_outputs(887));
    layer2_outputs(3570) <= (layer1_outputs(1227)) or (layer1_outputs(4234));
    layer2_outputs(3571) <= layer1_outputs(4615);
    layer2_outputs(3572) <= (layer1_outputs(4151)) and not (layer1_outputs(4972));
    layer2_outputs(3573) <= not((layer1_outputs(3301)) and (layer1_outputs(4517)));
    layer2_outputs(3574) <= not(layer1_outputs(3620)) or (layer1_outputs(2522));
    layer2_outputs(3575) <= layer1_outputs(6338);
    layer2_outputs(3576) <= '0';
    layer2_outputs(3577) <= not(layer1_outputs(6131));
    layer2_outputs(3578) <= not(layer1_outputs(5946));
    layer2_outputs(3579) <= not((layer1_outputs(7629)) xor (layer1_outputs(1965)));
    layer2_outputs(3580) <= (layer1_outputs(6091)) and not (layer1_outputs(1472));
    layer2_outputs(3581) <= (layer1_outputs(7189)) xor (layer1_outputs(2198));
    layer2_outputs(3582) <= (layer1_outputs(3329)) or (layer1_outputs(4703));
    layer2_outputs(3583) <= not((layer1_outputs(915)) or (layer1_outputs(3976)));
    layer2_outputs(3584) <= '0';
    layer2_outputs(3585) <= (layer1_outputs(5293)) and (layer1_outputs(3846));
    layer2_outputs(3586) <= not(layer1_outputs(2747)) or (layer1_outputs(3658));
    layer2_outputs(3587) <= not(layer1_outputs(3152)) or (layer1_outputs(3869));
    layer2_outputs(3588) <= not(layer1_outputs(6879)) or (layer1_outputs(432));
    layer2_outputs(3589) <= (layer1_outputs(7036)) and (layer1_outputs(5332));
    layer2_outputs(3590) <= layer1_outputs(3136);
    layer2_outputs(3591) <= '0';
    layer2_outputs(3592) <= not((layer1_outputs(2160)) and (layer1_outputs(5932)));
    layer2_outputs(3593) <= not(layer1_outputs(1989));
    layer2_outputs(3594) <= (layer1_outputs(2423)) and not (layer1_outputs(4987));
    layer2_outputs(3595) <= (layer1_outputs(184)) and not (layer1_outputs(488));
    layer2_outputs(3596) <= (layer1_outputs(6172)) and not (layer1_outputs(6301));
    layer2_outputs(3597) <= layer1_outputs(6345);
    layer2_outputs(3598) <= not((layer1_outputs(1147)) and (layer1_outputs(5108)));
    layer2_outputs(3599) <= not((layer1_outputs(6983)) and (layer1_outputs(675)));
    layer2_outputs(3600) <= layer1_outputs(3764);
    layer2_outputs(3601) <= layer1_outputs(2805);
    layer2_outputs(3602) <= layer1_outputs(6348);
    layer2_outputs(3603) <= (layer1_outputs(2892)) and not (layer1_outputs(2346));
    layer2_outputs(3604) <= layer1_outputs(7363);
    layer2_outputs(3605) <= (layer1_outputs(1625)) and not (layer1_outputs(859));
    layer2_outputs(3606) <= not(layer1_outputs(309)) or (layer1_outputs(4692));
    layer2_outputs(3607) <= not(layer1_outputs(7421));
    layer2_outputs(3608) <= not(layer1_outputs(3791)) or (layer1_outputs(4494));
    layer2_outputs(3609) <= layer1_outputs(4272);
    layer2_outputs(3610) <= not(layer1_outputs(5963));
    layer2_outputs(3611) <= (layer1_outputs(3002)) and not (layer1_outputs(2793));
    layer2_outputs(3612) <= (layer1_outputs(2726)) or (layer1_outputs(1645));
    layer2_outputs(3613) <= '0';
    layer2_outputs(3614) <= not(layer1_outputs(5654));
    layer2_outputs(3615) <= layer1_outputs(1027);
    layer2_outputs(3616) <= '0';
    layer2_outputs(3617) <= (layer1_outputs(7328)) and not (layer1_outputs(3880));
    layer2_outputs(3618) <= not((layer1_outputs(6709)) and (layer1_outputs(2324)));
    layer2_outputs(3619) <= (layer1_outputs(6615)) and not (layer1_outputs(3958));
    layer2_outputs(3620) <= not(layer1_outputs(791)) or (layer1_outputs(434));
    layer2_outputs(3621) <= '1';
    layer2_outputs(3622) <= layer1_outputs(1457);
    layer2_outputs(3623) <= layer1_outputs(713);
    layer2_outputs(3624) <= not(layer1_outputs(336));
    layer2_outputs(3625) <= layer1_outputs(3103);
    layer2_outputs(3626) <= layer1_outputs(3798);
    layer2_outputs(3627) <= not(layer1_outputs(848)) or (layer1_outputs(5673));
    layer2_outputs(3628) <= layer1_outputs(5073);
    layer2_outputs(3629) <= layer1_outputs(1876);
    layer2_outputs(3630) <= layer1_outputs(6744);
    layer2_outputs(3631) <= not((layer1_outputs(5814)) xor (layer1_outputs(6240)));
    layer2_outputs(3632) <= not(layer1_outputs(3175));
    layer2_outputs(3633) <= (layer1_outputs(3866)) and (layer1_outputs(4259));
    layer2_outputs(3634) <= not((layer1_outputs(3439)) and (layer1_outputs(2351)));
    layer2_outputs(3635) <= not(layer1_outputs(6060)) or (layer1_outputs(4022));
    layer2_outputs(3636) <= not(layer1_outputs(4719));
    layer2_outputs(3637) <= layer1_outputs(6797);
    layer2_outputs(3638) <= not((layer1_outputs(1027)) and (layer1_outputs(752)));
    layer2_outputs(3639) <= not((layer1_outputs(494)) and (layer1_outputs(4035)));
    layer2_outputs(3640) <= layer1_outputs(4570);
    layer2_outputs(3641) <= (layer1_outputs(2843)) and (layer1_outputs(5083));
    layer2_outputs(3642) <= layer1_outputs(6398);
    layer2_outputs(3643) <= not(layer1_outputs(2073));
    layer2_outputs(3644) <= layer1_outputs(6324);
    layer2_outputs(3645) <= not((layer1_outputs(1015)) and (layer1_outputs(6390)));
    layer2_outputs(3646) <= (layer1_outputs(3235)) and not (layer1_outputs(4130));
    layer2_outputs(3647) <= (layer1_outputs(4762)) or (layer1_outputs(1409));
    layer2_outputs(3648) <= layer1_outputs(3405);
    layer2_outputs(3649) <= (layer1_outputs(7101)) and not (layer1_outputs(7503));
    layer2_outputs(3650) <= not((layer1_outputs(6104)) or (layer1_outputs(2934)));
    layer2_outputs(3651) <= not(layer1_outputs(5682));
    layer2_outputs(3652) <= layer1_outputs(3793);
    layer2_outputs(3653) <= '1';
    layer2_outputs(3654) <= layer1_outputs(271);
    layer2_outputs(3655) <= not(layer1_outputs(5993)) or (layer1_outputs(1975));
    layer2_outputs(3656) <= not(layer1_outputs(2413));
    layer2_outputs(3657) <= not((layer1_outputs(6149)) and (layer1_outputs(2094)));
    layer2_outputs(3658) <= not((layer1_outputs(4349)) or (layer1_outputs(1263)));
    layer2_outputs(3659) <= not(layer1_outputs(1660)) or (layer1_outputs(3988));
    layer2_outputs(3660) <= not((layer1_outputs(3019)) or (layer1_outputs(3877)));
    layer2_outputs(3661) <= not((layer1_outputs(2743)) xor (layer1_outputs(2242)));
    layer2_outputs(3662) <= not(layer1_outputs(6766)) or (layer1_outputs(2896));
    layer2_outputs(3663) <= not((layer1_outputs(7431)) and (layer1_outputs(5604)));
    layer2_outputs(3664) <= not(layer1_outputs(7562));
    layer2_outputs(3665) <= not(layer1_outputs(5767));
    layer2_outputs(3666) <= not(layer1_outputs(902)) or (layer1_outputs(7049));
    layer2_outputs(3667) <= layer1_outputs(2997);
    layer2_outputs(3668) <= layer1_outputs(3465);
    layer2_outputs(3669) <= layer1_outputs(3602);
    layer2_outputs(3670) <= (layer1_outputs(2320)) and (layer1_outputs(5365));
    layer2_outputs(3671) <= not(layer1_outputs(2054));
    layer2_outputs(3672) <= (layer1_outputs(7176)) or (layer1_outputs(4639));
    layer2_outputs(3673) <= (layer1_outputs(1395)) or (layer1_outputs(721));
    layer2_outputs(3674) <= not((layer1_outputs(2528)) and (layer1_outputs(4967)));
    layer2_outputs(3675) <= '0';
    layer2_outputs(3676) <= not((layer1_outputs(860)) or (layer1_outputs(2016)));
    layer2_outputs(3677) <= not(layer1_outputs(6180));
    layer2_outputs(3678) <= layer1_outputs(3874);
    layer2_outputs(3679) <= not(layer1_outputs(4790));
    layer2_outputs(3680) <= not(layer1_outputs(1175));
    layer2_outputs(3681) <= (layer1_outputs(4356)) xor (layer1_outputs(193));
    layer2_outputs(3682) <= not((layer1_outputs(6127)) and (layer1_outputs(2708)));
    layer2_outputs(3683) <= not((layer1_outputs(6574)) or (layer1_outputs(5333)));
    layer2_outputs(3684) <= '1';
    layer2_outputs(3685) <= layer1_outputs(2250);
    layer2_outputs(3686) <= (layer1_outputs(6714)) and (layer1_outputs(1328));
    layer2_outputs(3687) <= not(layer1_outputs(4760));
    layer2_outputs(3688) <= not((layer1_outputs(6019)) or (layer1_outputs(1225)));
    layer2_outputs(3689) <= (layer1_outputs(1948)) and (layer1_outputs(2735));
    layer2_outputs(3690) <= not(layer1_outputs(4612));
    layer2_outputs(3691) <= not(layer1_outputs(4760));
    layer2_outputs(3692) <= not(layer1_outputs(1051)) or (layer1_outputs(5150));
    layer2_outputs(3693) <= layer1_outputs(69);
    layer2_outputs(3694) <= not(layer1_outputs(1583));
    layer2_outputs(3695) <= layer1_outputs(694);
    layer2_outputs(3696) <= not(layer1_outputs(4890));
    layer2_outputs(3697) <= not(layer1_outputs(6604)) or (layer1_outputs(6139));
    layer2_outputs(3698) <= (layer1_outputs(3338)) and not (layer1_outputs(601));
    layer2_outputs(3699) <= not((layer1_outputs(4396)) xor (layer1_outputs(5998)));
    layer2_outputs(3700) <= '0';
    layer2_outputs(3701) <= (layer1_outputs(7410)) and not (layer1_outputs(1481));
    layer2_outputs(3702) <= not((layer1_outputs(4916)) xor (layer1_outputs(5062)));
    layer2_outputs(3703) <= (layer1_outputs(425)) and not (layer1_outputs(6846));
    layer2_outputs(3704) <= (layer1_outputs(7367)) and not (layer1_outputs(837));
    layer2_outputs(3705) <= layer1_outputs(6970);
    layer2_outputs(3706) <= (layer1_outputs(6029)) or (layer1_outputs(3657));
    layer2_outputs(3707) <= (layer1_outputs(1884)) and not (layer1_outputs(6647));
    layer2_outputs(3708) <= layer1_outputs(5509);
    layer2_outputs(3709) <= not(layer1_outputs(360)) or (layer1_outputs(2958));
    layer2_outputs(3710) <= (layer1_outputs(1488)) and (layer1_outputs(1323));
    layer2_outputs(3711) <= not((layer1_outputs(4753)) and (layer1_outputs(7580)));
    layer2_outputs(3712) <= (layer1_outputs(3803)) and not (layer1_outputs(4944));
    layer2_outputs(3713) <= not(layer1_outputs(2107)) or (layer1_outputs(2869));
    layer2_outputs(3714) <= '1';
    layer2_outputs(3715) <= layer1_outputs(1766);
    layer2_outputs(3716) <= not((layer1_outputs(2740)) or (layer1_outputs(7501)));
    layer2_outputs(3717) <= (layer1_outputs(3925)) or (layer1_outputs(2625));
    layer2_outputs(3718) <= not((layer1_outputs(5996)) and (layer1_outputs(7469)));
    layer2_outputs(3719) <= not(layer1_outputs(1743)) or (layer1_outputs(2205));
    layer2_outputs(3720) <= (layer1_outputs(5791)) and not (layer1_outputs(4473));
    layer2_outputs(3721) <= not(layer1_outputs(3366));
    layer2_outputs(3722) <= (layer1_outputs(5639)) and not (layer1_outputs(4506));
    layer2_outputs(3723) <= (layer1_outputs(6428)) or (layer1_outputs(4710));
    layer2_outputs(3724) <= not(layer1_outputs(2293)) or (layer1_outputs(3854));
    layer2_outputs(3725) <= not(layer1_outputs(7663));
    layer2_outputs(3726) <= not(layer1_outputs(5879)) or (layer1_outputs(7591));
    layer2_outputs(3727) <= layer1_outputs(3444);
    layer2_outputs(3728) <= not(layer1_outputs(6577)) or (layer1_outputs(6195));
    layer2_outputs(3729) <= '0';
    layer2_outputs(3730) <= not(layer1_outputs(5064)) or (layer1_outputs(5781));
    layer2_outputs(3731) <= not(layer1_outputs(5350)) or (layer1_outputs(7080));
    layer2_outputs(3732) <= not(layer1_outputs(7382));
    layer2_outputs(3733) <= not(layer1_outputs(7408));
    layer2_outputs(3734) <= not(layer1_outputs(3047)) or (layer1_outputs(1244));
    layer2_outputs(3735) <= (layer1_outputs(3371)) xor (layer1_outputs(7323));
    layer2_outputs(3736) <= not(layer1_outputs(1175));
    layer2_outputs(3737) <= layer1_outputs(4227);
    layer2_outputs(3738) <= not(layer1_outputs(2320)) or (layer1_outputs(81));
    layer2_outputs(3739) <= not(layer1_outputs(4730));
    layer2_outputs(3740) <= (layer1_outputs(4863)) and not (layer1_outputs(3043));
    layer2_outputs(3741) <= not((layer1_outputs(3870)) and (layer1_outputs(6556)));
    layer2_outputs(3742) <= (layer1_outputs(7174)) and not (layer1_outputs(3489));
    layer2_outputs(3743) <= not(layer1_outputs(6663));
    layer2_outputs(3744) <= (layer1_outputs(4327)) and not (layer1_outputs(1921));
    layer2_outputs(3745) <= '1';
    layer2_outputs(3746) <= not(layer1_outputs(294));
    layer2_outputs(3747) <= '0';
    layer2_outputs(3748) <= not(layer1_outputs(6699));
    layer2_outputs(3749) <= (layer1_outputs(156)) and (layer1_outputs(3071));
    layer2_outputs(3750) <= (layer1_outputs(6561)) and not (layer1_outputs(6572));
    layer2_outputs(3751) <= (layer1_outputs(6244)) and not (layer1_outputs(6257));
    layer2_outputs(3752) <= not((layer1_outputs(3172)) xor (layer1_outputs(6712)));
    layer2_outputs(3753) <= layer1_outputs(2918);
    layer2_outputs(3754) <= not(layer1_outputs(6585));
    layer2_outputs(3755) <= not(layer1_outputs(477)) or (layer1_outputs(500));
    layer2_outputs(3756) <= not((layer1_outputs(2167)) and (layer1_outputs(2993)));
    layer2_outputs(3757) <= (layer1_outputs(1805)) and (layer1_outputs(7354));
    layer2_outputs(3758) <= (layer1_outputs(7526)) and (layer1_outputs(1665));
    layer2_outputs(3759) <= (layer1_outputs(2495)) and not (layer1_outputs(2261));
    layer2_outputs(3760) <= not(layer1_outputs(6968));
    layer2_outputs(3761) <= not((layer1_outputs(4990)) and (layer1_outputs(5174)));
    layer2_outputs(3762) <= (layer1_outputs(2341)) and (layer1_outputs(5190));
    layer2_outputs(3763) <= '1';
    layer2_outputs(3764) <= (layer1_outputs(1481)) or (layer1_outputs(2315));
    layer2_outputs(3765) <= not(layer1_outputs(4130));
    layer2_outputs(3766) <= layer1_outputs(7130);
    layer2_outputs(3767) <= not(layer1_outputs(7109));
    layer2_outputs(3768) <= not(layer1_outputs(4053));
    layer2_outputs(3769) <= (layer1_outputs(715)) and not (layer1_outputs(3561));
    layer2_outputs(3770) <= layer1_outputs(466);
    layer2_outputs(3771) <= not(layer1_outputs(5490)) or (layer1_outputs(4620));
    layer2_outputs(3772) <= layer1_outputs(4249);
    layer2_outputs(3773) <= not(layer1_outputs(7132));
    layer2_outputs(3774) <= not(layer1_outputs(6831));
    layer2_outputs(3775) <= not(layer1_outputs(3750));
    layer2_outputs(3776) <= layer1_outputs(1705);
    layer2_outputs(3777) <= not(layer1_outputs(7045));
    layer2_outputs(3778) <= not(layer1_outputs(269));
    layer2_outputs(3779) <= (layer1_outputs(3055)) and not (layer1_outputs(508));
    layer2_outputs(3780) <= (layer1_outputs(7432)) and (layer1_outputs(6916));
    layer2_outputs(3781) <= (layer1_outputs(3615)) and not (layer1_outputs(672));
    layer2_outputs(3782) <= layer1_outputs(6003);
    layer2_outputs(3783) <= layer1_outputs(1306);
    layer2_outputs(3784) <= layer1_outputs(59);
    layer2_outputs(3785) <= not(layer1_outputs(4645)) or (layer1_outputs(2877));
    layer2_outputs(3786) <= layer1_outputs(1006);
    layer2_outputs(3787) <= (layer1_outputs(6835)) or (layer1_outputs(1045));
    layer2_outputs(3788) <= layer1_outputs(246);
    layer2_outputs(3789) <= (layer1_outputs(3788)) and (layer1_outputs(4945));
    layer2_outputs(3790) <= not((layer1_outputs(3987)) or (layer1_outputs(2261)));
    layer2_outputs(3791) <= '0';
    layer2_outputs(3792) <= not(layer1_outputs(4737));
    layer2_outputs(3793) <= (layer1_outputs(5180)) or (layer1_outputs(7204));
    layer2_outputs(3794) <= (layer1_outputs(6746)) or (layer1_outputs(1631));
    layer2_outputs(3795) <= layer1_outputs(5171);
    layer2_outputs(3796) <= layer1_outputs(5115);
    layer2_outputs(3797) <= (layer1_outputs(1073)) and not (layer1_outputs(7353));
    layer2_outputs(3798) <= '0';
    layer2_outputs(3799) <= layer1_outputs(4971);
    layer2_outputs(3800) <= layer1_outputs(3376);
    layer2_outputs(3801) <= not(layer1_outputs(5132));
    layer2_outputs(3802) <= '0';
    layer2_outputs(3803) <= layer1_outputs(1394);
    layer2_outputs(3804) <= (layer1_outputs(3461)) and (layer1_outputs(2105));
    layer2_outputs(3805) <= not(layer1_outputs(1035)) or (layer1_outputs(2623));
    layer2_outputs(3806) <= layer1_outputs(2168);
    layer2_outputs(3807) <= (layer1_outputs(399)) xor (layer1_outputs(6341));
    layer2_outputs(3808) <= not(layer1_outputs(2354));
    layer2_outputs(3809) <= (layer1_outputs(1160)) and not (layer1_outputs(296));
    layer2_outputs(3810) <= layer1_outputs(5815);
    layer2_outputs(3811) <= not(layer1_outputs(6307));
    layer2_outputs(3812) <= layer1_outputs(2617);
    layer2_outputs(3813) <= not(layer1_outputs(6198));
    layer2_outputs(3814) <= not(layer1_outputs(4118));
    layer2_outputs(3815) <= not(layer1_outputs(4662)) or (layer1_outputs(7449));
    layer2_outputs(3816) <= (layer1_outputs(7406)) or (layer1_outputs(2979));
    layer2_outputs(3817) <= (layer1_outputs(1689)) and (layer1_outputs(1973));
    layer2_outputs(3818) <= not((layer1_outputs(7366)) or (layer1_outputs(4442)));
    layer2_outputs(3819) <= layer1_outputs(4264);
    layer2_outputs(3820) <= not(layer1_outputs(3100));
    layer2_outputs(3821) <= not(layer1_outputs(6004));
    layer2_outputs(3822) <= (layer1_outputs(1581)) and not (layer1_outputs(194));
    layer2_outputs(3823) <= (layer1_outputs(4164)) or (layer1_outputs(56));
    layer2_outputs(3824) <= (layer1_outputs(5484)) and not (layer1_outputs(691));
    layer2_outputs(3825) <= layer1_outputs(6811);
    layer2_outputs(3826) <= layer1_outputs(6581);
    layer2_outputs(3827) <= not(layer1_outputs(2720)) or (layer1_outputs(1256));
    layer2_outputs(3828) <= layer1_outputs(1197);
    layer2_outputs(3829) <= (layer1_outputs(3282)) and (layer1_outputs(2917));
    layer2_outputs(3830) <= (layer1_outputs(2538)) and not (layer1_outputs(3316));
    layer2_outputs(3831) <= not(layer1_outputs(5759));
    layer2_outputs(3832) <= not(layer1_outputs(3437));
    layer2_outputs(3833) <= not(layer1_outputs(1495));
    layer2_outputs(3834) <= (layer1_outputs(3331)) and not (layer1_outputs(2724));
    layer2_outputs(3835) <= (layer1_outputs(4187)) or (layer1_outputs(4233));
    layer2_outputs(3836) <= not((layer1_outputs(2004)) and (layer1_outputs(2689)));
    layer2_outputs(3837) <= (layer1_outputs(5065)) and (layer1_outputs(2247));
    layer2_outputs(3838) <= (layer1_outputs(1121)) and (layer1_outputs(1830));
    layer2_outputs(3839) <= (layer1_outputs(3862)) and not (layer1_outputs(2536));
    layer2_outputs(3840) <= layer1_outputs(5218);
    layer2_outputs(3841) <= '0';
    layer2_outputs(3842) <= not(layer1_outputs(3577));
    layer2_outputs(3843) <= not(layer1_outputs(1489));
    layer2_outputs(3844) <= (layer1_outputs(6723)) or (layer1_outputs(6045));
    layer2_outputs(3845) <= (layer1_outputs(6512)) or (layer1_outputs(4469));
    layer2_outputs(3846) <= not((layer1_outputs(3399)) or (layer1_outputs(5418)));
    layer2_outputs(3847) <= layer1_outputs(52);
    layer2_outputs(3848) <= (layer1_outputs(6914)) and (layer1_outputs(5050));
    layer2_outputs(3849) <= not(layer1_outputs(2551));
    layer2_outputs(3850) <= not(layer1_outputs(1667)) or (layer1_outputs(4920));
    layer2_outputs(3851) <= not(layer1_outputs(4509));
    layer2_outputs(3852) <= not((layer1_outputs(1957)) and (layer1_outputs(4602)));
    layer2_outputs(3853) <= not((layer1_outputs(4236)) or (layer1_outputs(3191)));
    layer2_outputs(3854) <= not(layer1_outputs(1421)) or (layer1_outputs(771));
    layer2_outputs(3855) <= not(layer1_outputs(7670));
    layer2_outputs(3856) <= not(layer1_outputs(1603)) or (layer1_outputs(3802));
    layer2_outputs(3857) <= not(layer1_outputs(1662));
    layer2_outputs(3858) <= (layer1_outputs(4610)) and not (layer1_outputs(3794));
    layer2_outputs(3859) <= (layer1_outputs(4747)) and not (layer1_outputs(3268));
    layer2_outputs(3860) <= (layer1_outputs(367)) and not (layer1_outputs(2019));
    layer2_outputs(3861) <= not(layer1_outputs(4879)) or (layer1_outputs(2924));
    layer2_outputs(3862) <= not(layer1_outputs(7238));
    layer2_outputs(3863) <= not((layer1_outputs(863)) or (layer1_outputs(1646)));
    layer2_outputs(3864) <= not((layer1_outputs(5620)) or (layer1_outputs(4601)));
    layer2_outputs(3865) <= (layer1_outputs(6506)) and not (layer1_outputs(1621));
    layer2_outputs(3866) <= not(layer1_outputs(4621));
    layer2_outputs(3867) <= not((layer1_outputs(322)) xor (layer1_outputs(997)));
    layer2_outputs(3868) <= (layer1_outputs(680)) or (layer1_outputs(801));
    layer2_outputs(3869) <= (layer1_outputs(2225)) and (layer1_outputs(3131));
    layer2_outputs(3870) <= not((layer1_outputs(164)) or (layer1_outputs(6011)));
    layer2_outputs(3871) <= not(layer1_outputs(6210)) or (layer1_outputs(3026));
    layer2_outputs(3872) <= not(layer1_outputs(3547)) or (layer1_outputs(4138));
    layer2_outputs(3873) <= not(layer1_outputs(3730));
    layer2_outputs(3874) <= (layer1_outputs(2872)) and (layer1_outputs(784));
    layer2_outputs(3875) <= (layer1_outputs(1064)) and not (layer1_outputs(582));
    layer2_outputs(3876) <= (layer1_outputs(6236)) and (layer1_outputs(1588));
    layer2_outputs(3877) <= not(layer1_outputs(5988));
    layer2_outputs(3878) <= not(layer1_outputs(4528));
    layer2_outputs(3879) <= layer1_outputs(5127);
    layer2_outputs(3880) <= '0';
    layer2_outputs(3881) <= layer1_outputs(103);
    layer2_outputs(3882) <= layer1_outputs(7533);
    layer2_outputs(3883) <= (layer1_outputs(941)) or (layer1_outputs(4909));
    layer2_outputs(3884) <= '0';
    layer2_outputs(3885) <= not(layer1_outputs(4960));
    layer2_outputs(3886) <= not(layer1_outputs(4267));
    layer2_outputs(3887) <= not(layer1_outputs(1312));
    layer2_outputs(3888) <= not(layer1_outputs(6324)) or (layer1_outputs(2071));
    layer2_outputs(3889) <= (layer1_outputs(3999)) and (layer1_outputs(5503));
    layer2_outputs(3890) <= not((layer1_outputs(2468)) or (layer1_outputs(5391)));
    layer2_outputs(3891) <= (layer1_outputs(2301)) and not (layer1_outputs(5527));
    layer2_outputs(3892) <= not(layer1_outputs(3908));
    layer2_outputs(3893) <= (layer1_outputs(1633)) and (layer1_outputs(2919));
    layer2_outputs(3894) <= not((layer1_outputs(219)) and (layer1_outputs(5900)));
    layer2_outputs(3895) <= not((layer1_outputs(7480)) xor (layer1_outputs(1776)));
    layer2_outputs(3896) <= not((layer1_outputs(6379)) or (layer1_outputs(5006)));
    layer2_outputs(3897) <= (layer1_outputs(2458)) or (layer1_outputs(7653));
    layer2_outputs(3898) <= not((layer1_outputs(345)) and (layer1_outputs(4465)));
    layer2_outputs(3899) <= (layer1_outputs(551)) and not (layer1_outputs(7515));
    layer2_outputs(3900) <= not((layer1_outputs(7133)) or (layer1_outputs(119)));
    layer2_outputs(3901) <= not(layer1_outputs(3057));
    layer2_outputs(3902) <= not(layer1_outputs(958));
    layer2_outputs(3903) <= (layer1_outputs(756)) or (layer1_outputs(6922));
    layer2_outputs(3904) <= '1';
    layer2_outputs(3905) <= (layer1_outputs(1377)) and (layer1_outputs(7302));
    layer2_outputs(3906) <= layer1_outputs(4677);
    layer2_outputs(3907) <= not((layer1_outputs(4547)) or (layer1_outputs(4957)));
    layer2_outputs(3908) <= layer1_outputs(1767);
    layer2_outputs(3909) <= (layer1_outputs(36)) or (layer1_outputs(2336));
    layer2_outputs(3910) <= not(layer1_outputs(2790)) or (layer1_outputs(7368));
    layer2_outputs(3911) <= (layer1_outputs(1134)) xor (layer1_outputs(4107));
    layer2_outputs(3912) <= not(layer1_outputs(2995)) or (layer1_outputs(3021));
    layer2_outputs(3913) <= not(layer1_outputs(1452)) or (layer1_outputs(4268));
    layer2_outputs(3914) <= '0';
    layer2_outputs(3915) <= not(layer1_outputs(1527));
    layer2_outputs(3916) <= layer1_outputs(5728);
    layer2_outputs(3917) <= layer1_outputs(6820);
    layer2_outputs(3918) <= layer1_outputs(6258);
    layer2_outputs(3919) <= (layer1_outputs(1518)) and (layer1_outputs(655));
    layer2_outputs(3920) <= not(layer1_outputs(1640)) or (layer1_outputs(879));
    layer2_outputs(3921) <= not(layer1_outputs(6715));
    layer2_outputs(3922) <= not((layer1_outputs(6636)) xor (layer1_outputs(2807)));
    layer2_outputs(3923) <= (layer1_outputs(4976)) and not (layer1_outputs(6629));
    layer2_outputs(3924) <= not(layer1_outputs(1683)) or (layer1_outputs(7479));
    layer2_outputs(3925) <= '1';
    layer2_outputs(3926) <= (layer1_outputs(3700)) or (layer1_outputs(5831));
    layer2_outputs(3927) <= (layer1_outputs(1792)) and not (layer1_outputs(2114));
    layer2_outputs(3928) <= not(layer1_outputs(3966)) or (layer1_outputs(2648));
    layer2_outputs(3929) <= '0';
    layer2_outputs(3930) <= (layer1_outputs(208)) xor (layer1_outputs(6604));
    layer2_outputs(3931) <= '0';
    layer2_outputs(3932) <= (layer1_outputs(3561)) and not (layer1_outputs(1232));
    layer2_outputs(3933) <= (layer1_outputs(3446)) and not (layer1_outputs(3122));
    layer2_outputs(3934) <= (layer1_outputs(6734)) and not (layer1_outputs(3215));
    layer2_outputs(3935) <= not(layer1_outputs(4359));
    layer2_outputs(3936) <= not(layer1_outputs(3951));
    layer2_outputs(3937) <= not((layer1_outputs(6578)) or (layer1_outputs(5507)));
    layer2_outputs(3938) <= '0';
    layer2_outputs(3939) <= not(layer1_outputs(2811));
    layer2_outputs(3940) <= not((layer1_outputs(3340)) and (layer1_outputs(2656)));
    layer2_outputs(3941) <= not((layer1_outputs(1498)) and (layer1_outputs(3863)));
    layer2_outputs(3942) <= (layer1_outputs(6840)) and not (layer1_outputs(1475));
    layer2_outputs(3943) <= not((layer1_outputs(6028)) xor (layer1_outputs(6757)));
    layer2_outputs(3944) <= not(layer1_outputs(1562)) or (layer1_outputs(7277));
    layer2_outputs(3945) <= '1';
    layer2_outputs(3946) <= not(layer1_outputs(2224)) or (layer1_outputs(4248));
    layer2_outputs(3947) <= (layer1_outputs(3220)) and not (layer1_outputs(313));
    layer2_outputs(3948) <= layer1_outputs(7122);
    layer2_outputs(3949) <= (layer1_outputs(4933)) and (layer1_outputs(4171));
    layer2_outputs(3950) <= not(layer1_outputs(4792)) or (layer1_outputs(1857));
    layer2_outputs(3951) <= layer1_outputs(5534);
    layer2_outputs(3952) <= layer1_outputs(3206);
    layer2_outputs(3953) <= layer1_outputs(2145);
    layer2_outputs(3954) <= not(layer1_outputs(4722)) or (layer1_outputs(7307));
    layer2_outputs(3955) <= (layer1_outputs(4068)) and (layer1_outputs(6230));
    layer2_outputs(3956) <= not(layer1_outputs(3863)) or (layer1_outputs(616));
    layer2_outputs(3957) <= (layer1_outputs(6645)) and not (layer1_outputs(4427));
    layer2_outputs(3958) <= (layer1_outputs(6443)) and (layer1_outputs(5760));
    layer2_outputs(3959) <= (layer1_outputs(5116)) and not (layer1_outputs(3136));
    layer2_outputs(3960) <= layer1_outputs(6006);
    layer2_outputs(3961) <= (layer1_outputs(6427)) and not (layer1_outputs(464));
    layer2_outputs(3962) <= (layer1_outputs(6240)) and not (layer1_outputs(1520));
    layer2_outputs(3963) <= layer1_outputs(1357);
    layer2_outputs(3964) <= (layer1_outputs(4425)) or (layer1_outputs(4835));
    layer2_outputs(3965) <= (layer1_outputs(4761)) or (layer1_outputs(4751));
    layer2_outputs(3966) <= not(layer1_outputs(1042));
    layer2_outputs(3967) <= not((layer1_outputs(2369)) and (layer1_outputs(7355)));
    layer2_outputs(3968) <= '0';
    layer2_outputs(3969) <= not((layer1_outputs(6913)) or (layer1_outputs(78)));
    layer2_outputs(3970) <= not(layer1_outputs(6314));
    layer2_outputs(3971) <= '0';
    layer2_outputs(3972) <= layer1_outputs(6495);
    layer2_outputs(3973) <= (layer1_outputs(504)) and not (layer1_outputs(1672));
    layer2_outputs(3974) <= (layer1_outputs(7345)) xor (layer1_outputs(3809));
    layer2_outputs(3975) <= (layer1_outputs(1693)) and not (layer1_outputs(3552));
    layer2_outputs(3976) <= not((layer1_outputs(5620)) and (layer1_outputs(2331)));
    layer2_outputs(3977) <= (layer1_outputs(1675)) and not (layer1_outputs(7162));
    layer2_outputs(3978) <= not(layer1_outputs(4681)) or (layer1_outputs(3284));
    layer2_outputs(3979) <= not(layer1_outputs(5726)) or (layer1_outputs(3134));
    layer2_outputs(3980) <= not(layer1_outputs(7623));
    layer2_outputs(3981) <= (layer1_outputs(4809)) and not (layer1_outputs(2822));
    layer2_outputs(3982) <= (layer1_outputs(6692)) or (layer1_outputs(4864));
    layer2_outputs(3983) <= (layer1_outputs(5861)) and not (layer1_outputs(5549));
    layer2_outputs(3984) <= not(layer1_outputs(5859)) or (layer1_outputs(5993));
    layer2_outputs(3985) <= (layer1_outputs(445)) and (layer1_outputs(1466));
    layer2_outputs(3986) <= not((layer1_outputs(7326)) or (layer1_outputs(3743)));
    layer2_outputs(3987) <= (layer1_outputs(1130)) and (layer1_outputs(773));
    layer2_outputs(3988) <= (layer1_outputs(7058)) or (layer1_outputs(2066));
    layer2_outputs(3989) <= not(layer1_outputs(3017)) or (layer1_outputs(3853));
    layer2_outputs(3990) <= not(layer1_outputs(215));
    layer2_outputs(3991) <= not((layer1_outputs(4318)) and (layer1_outputs(1952)));
    layer2_outputs(3992) <= layer1_outputs(5008);
    layer2_outputs(3993) <= '1';
    layer2_outputs(3994) <= (layer1_outputs(1276)) and (layer1_outputs(3180));
    layer2_outputs(3995) <= not(layer1_outputs(2011)) or (layer1_outputs(4795));
    layer2_outputs(3996) <= not((layer1_outputs(2306)) or (layer1_outputs(3779)));
    layer2_outputs(3997) <= not((layer1_outputs(2671)) or (layer1_outputs(3498)));
    layer2_outputs(3998) <= layer1_outputs(894);
    layer2_outputs(3999) <= '0';
    layer2_outputs(4000) <= not(layer1_outputs(2170));
    layer2_outputs(4001) <= layer1_outputs(1424);
    layer2_outputs(4002) <= (layer1_outputs(2548)) and not (layer1_outputs(5610));
    layer2_outputs(4003) <= layer1_outputs(1111);
    layer2_outputs(4004) <= (layer1_outputs(1154)) or (layer1_outputs(2189));
    layer2_outputs(4005) <= layer1_outputs(6817);
    layer2_outputs(4006) <= (layer1_outputs(6252)) or (layer1_outputs(4));
    layer2_outputs(4007) <= layer1_outputs(775);
    layer2_outputs(4008) <= not((layer1_outputs(5624)) xor (layer1_outputs(2424)));
    layer2_outputs(4009) <= not((layer1_outputs(3031)) or (layer1_outputs(4635)));
    layer2_outputs(4010) <= not((layer1_outputs(5741)) and (layer1_outputs(7210)));
    layer2_outputs(4011) <= '1';
    layer2_outputs(4012) <= layer1_outputs(4838);
    layer2_outputs(4013) <= not(layer1_outputs(6952));
    layer2_outputs(4014) <= (layer1_outputs(7382)) or (layer1_outputs(523));
    layer2_outputs(4015) <= not(layer1_outputs(796)) or (layer1_outputs(5896));
    layer2_outputs(4016) <= (layer1_outputs(4869)) and not (layer1_outputs(4599));
    layer2_outputs(4017) <= not(layer1_outputs(4707));
    layer2_outputs(4018) <= not((layer1_outputs(7066)) and (layer1_outputs(2850)));
    layer2_outputs(4019) <= layer1_outputs(2067);
    layer2_outputs(4020) <= not(layer1_outputs(1650)) or (layer1_outputs(5775));
    layer2_outputs(4021) <= '1';
    layer2_outputs(4022) <= '0';
    layer2_outputs(4023) <= not((layer1_outputs(3857)) and (layer1_outputs(1029)));
    layer2_outputs(4024) <= layer1_outputs(4276);
    layer2_outputs(4025) <= layer1_outputs(3977);
    layer2_outputs(4026) <= '1';
    layer2_outputs(4027) <= not(layer1_outputs(5283));
    layer2_outputs(4028) <= not(layer1_outputs(864));
    layer2_outputs(4029) <= layer1_outputs(3998);
    layer2_outputs(4030) <= '0';
    layer2_outputs(4031) <= layer1_outputs(4731);
    layer2_outputs(4032) <= not(layer1_outputs(6814));
    layer2_outputs(4033) <= (layer1_outputs(970)) and not (layer1_outputs(5907));
    layer2_outputs(4034) <= not((layer1_outputs(1099)) and (layer1_outputs(915)));
    layer2_outputs(4035) <= layer1_outputs(2381);
    layer2_outputs(4036) <= layer1_outputs(6381);
    layer2_outputs(4037) <= not(layer1_outputs(6384)) or (layer1_outputs(5869));
    layer2_outputs(4038) <= layer1_outputs(7531);
    layer2_outputs(4039) <= '0';
    layer2_outputs(4040) <= not(layer1_outputs(6612)) or (layer1_outputs(6852));
    layer2_outputs(4041) <= (layer1_outputs(2423)) and not (layer1_outputs(4179));
    layer2_outputs(4042) <= not((layer1_outputs(1765)) and (layer1_outputs(4434)));
    layer2_outputs(4043) <= not(layer1_outputs(696)) or (layer1_outputs(7414));
    layer2_outputs(4044) <= not(layer1_outputs(3521));
    layer2_outputs(4045) <= not(layer1_outputs(1927));
    layer2_outputs(4046) <= not(layer1_outputs(3052));
    layer2_outputs(4047) <= layer1_outputs(4362);
    layer2_outputs(4048) <= not(layer1_outputs(2381));
    layer2_outputs(4049) <= (layer1_outputs(620)) or (layer1_outputs(950));
    layer2_outputs(4050) <= '1';
    layer2_outputs(4051) <= not((layer1_outputs(2617)) or (layer1_outputs(2751)));
    layer2_outputs(4052) <= not((layer1_outputs(3352)) and (layer1_outputs(5915)));
    layer2_outputs(4053) <= (layer1_outputs(5130)) and not (layer1_outputs(5856));
    layer2_outputs(4054) <= (layer1_outputs(1687)) and not (layer1_outputs(5890));
    layer2_outputs(4055) <= (layer1_outputs(3004)) or (layer1_outputs(4894));
    layer2_outputs(4056) <= not(layer1_outputs(5068)) or (layer1_outputs(2274));
    layer2_outputs(4057) <= (layer1_outputs(3478)) or (layer1_outputs(5377));
    layer2_outputs(4058) <= layer1_outputs(4059);
    layer2_outputs(4059) <= not((layer1_outputs(4442)) and (layer1_outputs(595)));
    layer2_outputs(4060) <= (layer1_outputs(2679)) and not (layer1_outputs(299));
    layer2_outputs(4061) <= not(layer1_outputs(7130));
    layer2_outputs(4062) <= not(layer1_outputs(4880));
    layer2_outputs(4063) <= (layer1_outputs(1599)) and not (layer1_outputs(5061));
    layer2_outputs(4064) <= (layer1_outputs(1157)) or (layer1_outputs(6297));
    layer2_outputs(4065) <= not(layer1_outputs(474)) or (layer1_outputs(3818));
    layer2_outputs(4066) <= (layer1_outputs(5944)) and not (layer1_outputs(2019));
    layer2_outputs(4067) <= layer1_outputs(1553);
    layer2_outputs(4068) <= layer1_outputs(2879);
    layer2_outputs(4069) <= (layer1_outputs(6356)) and (layer1_outputs(7272));
    layer2_outputs(4070) <= layer1_outputs(3235);
    layer2_outputs(4071) <= not(layer1_outputs(7526)) or (layer1_outputs(7406));
    layer2_outputs(4072) <= not((layer1_outputs(7388)) or (layer1_outputs(2542)));
    layer2_outputs(4073) <= layer1_outputs(7468);
    layer2_outputs(4074) <= not(layer1_outputs(7509));
    layer2_outputs(4075) <= (layer1_outputs(4262)) or (layer1_outputs(2366));
    layer2_outputs(4076) <= (layer1_outputs(333)) and not (layer1_outputs(3214));
    layer2_outputs(4077) <= '1';
    layer2_outputs(4078) <= not((layer1_outputs(3273)) or (layer1_outputs(4921)));
    layer2_outputs(4079) <= not(layer1_outputs(4997));
    layer2_outputs(4080) <= not(layer1_outputs(2991)) or (layer1_outputs(6713));
    layer2_outputs(4081) <= not(layer1_outputs(3466));
    layer2_outputs(4082) <= layer1_outputs(192);
    layer2_outputs(4083) <= (layer1_outputs(6322)) and (layer1_outputs(3272));
    layer2_outputs(4084) <= (layer1_outputs(5443)) and not (layer1_outputs(1606));
    layer2_outputs(4085) <= (layer1_outputs(6040)) and not (layer1_outputs(1951));
    layer2_outputs(4086) <= layer1_outputs(6488);
    layer2_outputs(4087) <= layer1_outputs(7082);
    layer2_outputs(4088) <= layer1_outputs(3938);
    layer2_outputs(4089) <= (layer1_outputs(2510)) or (layer1_outputs(3417));
    layer2_outputs(4090) <= not((layer1_outputs(1125)) xor (layer1_outputs(1198)));
    layer2_outputs(4091) <= layer1_outputs(3302);
    layer2_outputs(4092) <= not((layer1_outputs(6077)) xor (layer1_outputs(6615)));
    layer2_outputs(4093) <= not(layer1_outputs(743)) or (layer1_outputs(6969));
    layer2_outputs(4094) <= not(layer1_outputs(3878));
    layer2_outputs(4095) <= not(layer1_outputs(3375)) or (layer1_outputs(5783));
    layer2_outputs(4096) <= not(layer1_outputs(3937));
    layer2_outputs(4097) <= layer1_outputs(2087);
    layer2_outputs(4098) <= (layer1_outputs(7128)) and (layer1_outputs(778));
    layer2_outputs(4099) <= '0';
    layer2_outputs(4100) <= not((layer1_outputs(5830)) and (layer1_outputs(523)));
    layer2_outputs(4101) <= (layer1_outputs(3139)) or (layer1_outputs(4225));
    layer2_outputs(4102) <= not(layer1_outputs(3660)) or (layer1_outputs(1203));
    layer2_outputs(4103) <= layer1_outputs(1950);
    layer2_outputs(4104) <= not(layer1_outputs(5339));
    layer2_outputs(4105) <= not(layer1_outputs(3890));
    layer2_outputs(4106) <= layer1_outputs(6409);
    layer2_outputs(4107) <= (layer1_outputs(6562)) and (layer1_outputs(2176));
    layer2_outputs(4108) <= layer1_outputs(345);
    layer2_outputs(4109) <= '0';
    layer2_outputs(4110) <= layer1_outputs(634);
    layer2_outputs(4111) <= not(layer1_outputs(2127)) or (layer1_outputs(2661));
    layer2_outputs(4112) <= not(layer1_outputs(1591)) or (layer1_outputs(3335));
    layer2_outputs(4113) <= (layer1_outputs(2984)) or (layer1_outputs(1802));
    layer2_outputs(4114) <= (layer1_outputs(5664)) or (layer1_outputs(1464));
    layer2_outputs(4115) <= not(layer1_outputs(1180));
    layer2_outputs(4116) <= not(layer1_outputs(4135)) or (layer1_outputs(7559));
    layer2_outputs(4117) <= '0';
    layer2_outputs(4118) <= not(layer1_outputs(3834));
    layer2_outputs(4119) <= not(layer1_outputs(2706));
    layer2_outputs(4120) <= layer1_outputs(2087);
    layer2_outputs(4121) <= layer1_outputs(3179);
    layer2_outputs(4122) <= not(layer1_outputs(4275));
    layer2_outputs(4123) <= not((layer1_outputs(3544)) and (layer1_outputs(3081)));
    layer2_outputs(4124) <= not((layer1_outputs(2282)) xor (layer1_outputs(7615)));
    layer2_outputs(4125) <= not((layer1_outputs(3726)) and (layer1_outputs(7251)));
    layer2_outputs(4126) <= (layer1_outputs(5137)) and not (layer1_outputs(3134));
    layer2_outputs(4127) <= (layer1_outputs(5739)) or (layer1_outputs(3792));
    layer2_outputs(4128) <= not(layer1_outputs(3333));
    layer2_outputs(4129) <= not(layer1_outputs(2513));
    layer2_outputs(4130) <= (layer1_outputs(6603)) and (layer1_outputs(3380));
    layer2_outputs(4131) <= not((layer1_outputs(106)) xor (layer1_outputs(4682)));
    layer2_outputs(4132) <= not(layer1_outputs(6072));
    layer2_outputs(4133) <= not(layer1_outputs(2580));
    layer2_outputs(4134) <= (layer1_outputs(4554)) or (layer1_outputs(2318));
    layer2_outputs(4135) <= (layer1_outputs(3277)) and not (layer1_outputs(5763));
    layer2_outputs(4136) <= not(layer1_outputs(133));
    layer2_outputs(4137) <= not(layer1_outputs(2032));
    layer2_outputs(4138) <= not(layer1_outputs(569));
    layer2_outputs(4139) <= not((layer1_outputs(5617)) xor (layer1_outputs(3280)));
    layer2_outputs(4140) <= '1';
    layer2_outputs(4141) <= not((layer1_outputs(5705)) and (layer1_outputs(6291)));
    layer2_outputs(4142) <= (layer1_outputs(1500)) and not (layer1_outputs(1411));
    layer2_outputs(4143) <= layer1_outputs(5892);
    layer2_outputs(4144) <= '1';
    layer2_outputs(4145) <= (layer1_outputs(5699)) or (layer1_outputs(4785));
    layer2_outputs(4146) <= not((layer1_outputs(4706)) or (layer1_outputs(582)));
    layer2_outputs(4147) <= (layer1_outputs(4406)) and not (layer1_outputs(2480));
    layer2_outputs(4148) <= '1';
    layer2_outputs(4149) <= '0';
    layer2_outputs(4150) <= not(layer1_outputs(4358));
    layer2_outputs(4151) <= (layer1_outputs(5960)) and not (layer1_outputs(1114));
    layer2_outputs(4152) <= not(layer1_outputs(232)) or (layer1_outputs(3089));
    layer2_outputs(4153) <= layer1_outputs(5927);
    layer2_outputs(4154) <= (layer1_outputs(4825)) and not (layer1_outputs(159));
    layer2_outputs(4155) <= not(layer1_outputs(5543));
    layer2_outputs(4156) <= not(layer1_outputs(4495));
    layer2_outputs(4157) <= (layer1_outputs(1114)) and not (layer1_outputs(3117));
    layer2_outputs(4158) <= not(layer1_outputs(3813));
    layer2_outputs(4159) <= not(layer1_outputs(4176)) or (layer1_outputs(4782));
    layer2_outputs(4160) <= not(layer1_outputs(2166));
    layer2_outputs(4161) <= layer1_outputs(6224);
    layer2_outputs(4162) <= (layer1_outputs(4763)) or (layer1_outputs(3245));
    layer2_outputs(4163) <= layer1_outputs(5292);
    layer2_outputs(4164) <= '1';
    layer2_outputs(4165) <= not((layer1_outputs(5306)) or (layer1_outputs(1471)));
    layer2_outputs(4166) <= (layer1_outputs(250)) and not (layer1_outputs(4143));
    layer2_outputs(4167) <= not((layer1_outputs(2078)) xor (layer1_outputs(6295)));
    layer2_outputs(4168) <= '1';
    layer2_outputs(4169) <= layer1_outputs(2005);
    layer2_outputs(4170) <= (layer1_outputs(5107)) and (layer1_outputs(5348));
    layer2_outputs(4171) <= (layer1_outputs(5809)) and (layer1_outputs(4105));
    layer2_outputs(4172) <= not(layer1_outputs(4625));
    layer2_outputs(4173) <= not(layer1_outputs(5288));
    layer2_outputs(4174) <= (layer1_outputs(2330)) or (layer1_outputs(2666));
    layer2_outputs(4175) <= not((layer1_outputs(5792)) and (layer1_outputs(2371)));
    layer2_outputs(4176) <= (layer1_outputs(1404)) or (layer1_outputs(132));
    layer2_outputs(4177) <= not(layer1_outputs(4702)) or (layer1_outputs(4552));
    layer2_outputs(4178) <= (layer1_outputs(6798)) or (layer1_outputs(7071));
    layer2_outputs(4179) <= '0';
    layer2_outputs(4180) <= not((layer1_outputs(1871)) and (layer1_outputs(6490)));
    layer2_outputs(4181) <= layer1_outputs(6724);
    layer2_outputs(4182) <= not(layer1_outputs(4611));
    layer2_outputs(4183) <= layer1_outputs(7201);
    layer2_outputs(4184) <= layer1_outputs(1932);
    layer2_outputs(4185) <= '0';
    layer2_outputs(4186) <= not(layer1_outputs(3559));
    layer2_outputs(4187) <= not(layer1_outputs(7226));
    layer2_outputs(4188) <= not(layer1_outputs(760));
    layer2_outputs(4189) <= not(layer1_outputs(2225));
    layer2_outputs(4190) <= layer1_outputs(4363);
    layer2_outputs(4191) <= not(layer1_outputs(4920));
    layer2_outputs(4192) <= (layer1_outputs(5968)) and (layer1_outputs(7352));
    layer2_outputs(4193) <= not((layer1_outputs(857)) or (layer1_outputs(6984)));
    layer2_outputs(4194) <= not(layer1_outputs(1065));
    layer2_outputs(4195) <= not((layer1_outputs(6181)) and (layer1_outputs(7550)));
    layer2_outputs(4196) <= (layer1_outputs(3129)) and not (layer1_outputs(4805));
    layer2_outputs(4197) <= layer1_outputs(3691);
    layer2_outputs(4198) <= '0';
    layer2_outputs(4199) <= layer1_outputs(2332);
    layer2_outputs(4200) <= (layer1_outputs(5774)) and not (layer1_outputs(6708));
    layer2_outputs(4201) <= not(layer1_outputs(3384));
    layer2_outputs(4202) <= (layer1_outputs(1358)) and (layer1_outputs(3264));
    layer2_outputs(4203) <= layer1_outputs(362);
    layer2_outputs(4204) <= not(layer1_outputs(2348)) or (layer1_outputs(7167));
    layer2_outputs(4205) <= not(layer1_outputs(4576)) or (layer1_outputs(3442));
    layer2_outputs(4206) <= not(layer1_outputs(7073));
    layer2_outputs(4207) <= not(layer1_outputs(4798)) or (layer1_outputs(1871));
    layer2_outputs(4208) <= layer1_outputs(1346);
    layer2_outputs(4209) <= layer1_outputs(4562);
    layer2_outputs(4210) <= layer1_outputs(2614);
    layer2_outputs(4211) <= (layer1_outputs(6808)) and not (layer1_outputs(3806));
    layer2_outputs(4212) <= not(layer1_outputs(43)) or (layer1_outputs(6013));
    layer2_outputs(4213) <= layer1_outputs(1695);
    layer2_outputs(4214) <= '0';
    layer2_outputs(4215) <= (layer1_outputs(7669)) or (layer1_outputs(6350));
    layer2_outputs(4216) <= not((layer1_outputs(4899)) and (layer1_outputs(580)));
    layer2_outputs(4217) <= layer1_outputs(868);
    layer2_outputs(4218) <= not(layer1_outputs(7184)) or (layer1_outputs(2842));
    layer2_outputs(4219) <= not(layer1_outputs(1702)) or (layer1_outputs(4931));
    layer2_outputs(4220) <= layer1_outputs(2179);
    layer2_outputs(4221) <= layer1_outputs(1670);
    layer2_outputs(4222) <= layer1_outputs(5124);
    layer2_outputs(4223) <= layer1_outputs(6959);
    layer2_outputs(4224) <= layer1_outputs(3979);
    layer2_outputs(4225) <= '1';
    layer2_outputs(4226) <= not(layer1_outputs(3022));
    layer2_outputs(4227) <= not(layer1_outputs(2278));
    layer2_outputs(4228) <= layer1_outputs(1526);
    layer2_outputs(4229) <= layer1_outputs(4665);
    layer2_outputs(4230) <= layer1_outputs(3219);
    layer2_outputs(4231) <= not((layer1_outputs(1974)) or (layer1_outputs(3109)));
    layer2_outputs(4232) <= not(layer1_outputs(6232));
    layer2_outputs(4233) <= not(layer1_outputs(4660));
    layer2_outputs(4234) <= (layer1_outputs(653)) and (layer1_outputs(4376));
    layer2_outputs(4235) <= (layer1_outputs(6624)) or (layer1_outputs(507));
    layer2_outputs(4236) <= (layer1_outputs(4496)) or (layer1_outputs(2549));
    layer2_outputs(4237) <= layer1_outputs(2043);
    layer2_outputs(4238) <= not(layer1_outputs(3237)) or (layer1_outputs(530));
    layer2_outputs(4239) <= not((layer1_outputs(1738)) xor (layer1_outputs(3148)));
    layer2_outputs(4240) <= layer1_outputs(2302);
    layer2_outputs(4241) <= not((layer1_outputs(2590)) or (layer1_outputs(2534)));
    layer2_outputs(4242) <= not(layer1_outputs(7414)) or (layer1_outputs(7524));
    layer2_outputs(4243) <= (layer1_outputs(6477)) and (layer1_outputs(7266));
    layer2_outputs(4244) <= (layer1_outputs(2039)) or (layer1_outputs(4928));
    layer2_outputs(4245) <= not((layer1_outputs(3772)) or (layer1_outputs(1192)));
    layer2_outputs(4246) <= (layer1_outputs(6678)) and not (layer1_outputs(5043));
    layer2_outputs(4247) <= not(layer1_outputs(3252));
    layer2_outputs(4248) <= not(layer1_outputs(5537));
    layer2_outputs(4249) <= (layer1_outputs(7442)) and not (layer1_outputs(3695));
    layer2_outputs(4250) <= '0';
    layer2_outputs(4251) <= (layer1_outputs(2153)) and not (layer1_outputs(839));
    layer2_outputs(4252) <= (layer1_outputs(5592)) or (layer1_outputs(1998));
    layer2_outputs(4253) <= not((layer1_outputs(3133)) and (layer1_outputs(965)));
    layer2_outputs(4254) <= not(layer1_outputs(1927));
    layer2_outputs(4255) <= not(layer1_outputs(342));
    layer2_outputs(4256) <= layer1_outputs(2121);
    layer2_outputs(4257) <= layer1_outputs(4685);
    layer2_outputs(4258) <= (layer1_outputs(840)) and not (layer1_outputs(4794));
    layer2_outputs(4259) <= (layer1_outputs(5179)) or (layer1_outputs(1162));
    layer2_outputs(4260) <= (layer1_outputs(3345)) and not (layer1_outputs(2259));
    layer2_outputs(4261) <= not(layer1_outputs(7330));
    layer2_outputs(4262) <= layer1_outputs(7279);
    layer2_outputs(4263) <= layer1_outputs(5177);
    layer2_outputs(4264) <= not(layer1_outputs(5489));
    layer2_outputs(4265) <= (layer1_outputs(7087)) xor (layer1_outputs(7434));
    layer2_outputs(4266) <= '0';
    layer2_outputs(4267) <= not(layer1_outputs(5105)) or (layer1_outputs(5574));
    layer2_outputs(4268) <= not((layer1_outputs(5169)) and (layer1_outputs(6596)));
    layer2_outputs(4269) <= (layer1_outputs(4431)) and not (layer1_outputs(4330));
    layer2_outputs(4270) <= '1';
    layer2_outputs(4271) <= layer1_outputs(3528);
    layer2_outputs(4272) <= (layer1_outputs(4178)) and not (layer1_outputs(5494));
    layer2_outputs(4273) <= not(layer1_outputs(5785));
    layer2_outputs(4274) <= not(layer1_outputs(2942)) or (layer1_outputs(3940));
    layer2_outputs(4275) <= layer1_outputs(749);
    layer2_outputs(4276) <= layer1_outputs(11);
    layer2_outputs(4277) <= not(layer1_outputs(2537));
    layer2_outputs(4278) <= not(layer1_outputs(3510));
    layer2_outputs(4279) <= not(layer1_outputs(1510));
    layer2_outputs(4280) <= layer1_outputs(832);
    layer2_outputs(4281) <= (layer1_outputs(218)) and not (layer1_outputs(3836));
    layer2_outputs(4282) <= layer1_outputs(5955);
    layer2_outputs(4283) <= layer1_outputs(4479);
    layer2_outputs(4284) <= not((layer1_outputs(3963)) and (layer1_outputs(2439)));
    layer2_outputs(4285) <= layer1_outputs(4964);
    layer2_outputs(4286) <= layer1_outputs(6061);
    layer2_outputs(4287) <= not(layer1_outputs(1989));
    layer2_outputs(4288) <= (layer1_outputs(2886)) or (layer1_outputs(4952));
    layer2_outputs(4289) <= layer1_outputs(5520);
    layer2_outputs(4290) <= not(layer1_outputs(3184)) or (layer1_outputs(7490));
    layer2_outputs(4291) <= not(layer1_outputs(3284));
    layer2_outputs(4292) <= not((layer1_outputs(6298)) xor (layer1_outputs(3120)));
    layer2_outputs(4293) <= layer1_outputs(7223);
    layer2_outputs(4294) <= not((layer1_outputs(6292)) and (layer1_outputs(5400)));
    layer2_outputs(4295) <= not(layer1_outputs(3797));
    layer2_outputs(4296) <= layer1_outputs(694);
    layer2_outputs(4297) <= (layer1_outputs(7265)) and (layer1_outputs(5193));
    layer2_outputs(4298) <= not((layer1_outputs(5276)) xor (layer1_outputs(1656)));
    layer2_outputs(4299) <= not(layer1_outputs(3391));
    layer2_outputs(4300) <= not((layer1_outputs(6127)) and (layer1_outputs(6677)));
    layer2_outputs(4301) <= layer1_outputs(1278);
    layer2_outputs(4302) <= (layer1_outputs(3427)) and (layer1_outputs(7641));
    layer2_outputs(4303) <= not((layer1_outputs(5686)) or (layer1_outputs(606)));
    layer2_outputs(4304) <= layer1_outputs(2414);
    layer2_outputs(4305) <= not(layer1_outputs(2596)) or (layer1_outputs(6161));
    layer2_outputs(4306) <= layer1_outputs(6203);
    layer2_outputs(4307) <= '0';
    layer2_outputs(4308) <= not(layer1_outputs(7135));
    layer2_outputs(4309) <= not((layer1_outputs(3492)) and (layer1_outputs(6014)));
    layer2_outputs(4310) <= not(layer1_outputs(5944)) or (layer1_outputs(4279));
    layer2_outputs(4311) <= not((layer1_outputs(247)) or (layer1_outputs(1446)));
    layer2_outputs(4312) <= not(layer1_outputs(1672));
    layer2_outputs(4313) <= layer1_outputs(1875);
    layer2_outputs(4314) <= layer1_outputs(1249);
    layer2_outputs(4315) <= not(layer1_outputs(457));
    layer2_outputs(4316) <= (layer1_outputs(1410)) and not (layer1_outputs(6605));
    layer2_outputs(4317) <= layer1_outputs(6768);
    layer2_outputs(4318) <= '0';
    layer2_outputs(4319) <= not((layer1_outputs(5737)) or (layer1_outputs(1299)));
    layer2_outputs(4320) <= layer1_outputs(6143);
    layer2_outputs(4321) <= (layer1_outputs(4016)) or (layer1_outputs(5113));
    layer2_outputs(4322) <= '0';
    layer2_outputs(4323) <= not((layer1_outputs(3883)) or (layer1_outputs(3285)));
    layer2_outputs(4324) <= not((layer1_outputs(6146)) xor (layer1_outputs(2506)));
    layer2_outputs(4325) <= (layer1_outputs(1347)) and not (layer1_outputs(1767));
    layer2_outputs(4326) <= not((layer1_outputs(6614)) or (layer1_outputs(2177)));
    layer2_outputs(4327) <= not(layer1_outputs(4395)) or (layer1_outputs(6301));
    layer2_outputs(4328) <= (layer1_outputs(1351)) and not (layer1_outputs(2200));
    layer2_outputs(4329) <= (layer1_outputs(1583)) and not (layer1_outputs(6189));
    layer2_outputs(4330) <= (layer1_outputs(5744)) xor (layer1_outputs(2384));
    layer2_outputs(4331) <= layer1_outputs(1568);
    layer2_outputs(4332) <= '1';
    layer2_outputs(4333) <= (layer1_outputs(167)) and not (layer1_outputs(2125));
    layer2_outputs(4334) <= not(layer1_outputs(6271));
    layer2_outputs(4335) <= not(layer1_outputs(1386));
    layer2_outputs(4336) <= '0';
    layer2_outputs(4337) <= '0';
    layer2_outputs(4338) <= not(layer1_outputs(7159)) or (layer1_outputs(3597));
    layer2_outputs(4339) <= '0';
    layer2_outputs(4340) <= not(layer1_outputs(3777)) or (layer1_outputs(2508));
    layer2_outputs(4341) <= not(layer1_outputs(2812));
    layer2_outputs(4342) <= not(layer1_outputs(6771));
    layer2_outputs(4343) <= (layer1_outputs(5147)) or (layer1_outputs(2108));
    layer2_outputs(4344) <= not(layer1_outputs(1680)) or (layer1_outputs(710));
    layer2_outputs(4345) <= not(layer1_outputs(2046)) or (layer1_outputs(6855));
    layer2_outputs(4346) <= (layer1_outputs(989)) and not (layer1_outputs(2628));
    layer2_outputs(4347) <= '0';
    layer2_outputs(4348) <= layer1_outputs(1119);
    layer2_outputs(4349) <= not((layer1_outputs(6351)) xor (layer1_outputs(6347)));
    layer2_outputs(4350) <= layer1_outputs(3939);
    layer2_outputs(4351) <= (layer1_outputs(1691)) and (layer1_outputs(1131));
    layer2_outputs(4352) <= layer1_outputs(6305);
    layer2_outputs(4353) <= not(layer1_outputs(4389));
    layer2_outputs(4354) <= not(layer1_outputs(6838));
    layer2_outputs(4355) <= not((layer1_outputs(512)) and (layer1_outputs(6911)));
    layer2_outputs(4356) <= layer1_outputs(18);
    layer2_outputs(4357) <= not((layer1_outputs(2952)) and (layer1_outputs(5110)));
    layer2_outputs(4358) <= not(layer1_outputs(4332));
    layer2_outputs(4359) <= layer1_outputs(4013);
    layer2_outputs(4360) <= not(layer1_outputs(1605)) or (layer1_outputs(2052));
    layer2_outputs(4361) <= layer1_outputs(6382);
    layer2_outputs(4362) <= (layer1_outputs(7588)) and not (layer1_outputs(42));
    layer2_outputs(4363) <= not(layer1_outputs(4142));
    layer2_outputs(4364) <= not((layer1_outputs(6609)) or (layer1_outputs(4699)));
    layer2_outputs(4365) <= '0';
    layer2_outputs(4366) <= (layer1_outputs(7177)) and not (layer1_outputs(6590));
    layer2_outputs(4367) <= (layer1_outputs(6504)) and (layer1_outputs(711));
    layer2_outputs(4368) <= layer1_outputs(4559);
    layer2_outputs(4369) <= layer1_outputs(5962);
    layer2_outputs(4370) <= (layer1_outputs(4056)) and not (layer1_outputs(6035));
    layer2_outputs(4371) <= layer1_outputs(3629);
    layer2_outputs(4372) <= not((layer1_outputs(330)) or (layer1_outputs(5212)));
    layer2_outputs(4373) <= (layer1_outputs(5060)) and not (layer1_outputs(1517));
    layer2_outputs(4374) <= not(layer1_outputs(4845));
    layer2_outputs(4375) <= '1';
    layer2_outputs(4376) <= layer1_outputs(5183);
    layer2_outputs(4377) <= not((layer1_outputs(6438)) or (layer1_outputs(1667)));
    layer2_outputs(4378) <= (layer1_outputs(594)) and not (layer1_outputs(6630));
    layer2_outputs(4379) <= not(layer1_outputs(5258));
    layer2_outputs(4380) <= not((layer1_outputs(2488)) and (layer1_outputs(3725)));
    layer2_outputs(4381) <= layer1_outputs(5030);
    layer2_outputs(4382) <= '1';
    layer2_outputs(4383) <= not(layer1_outputs(7635));
    layer2_outputs(4384) <= not(layer1_outputs(1990)) or (layer1_outputs(6259));
    layer2_outputs(4385) <= layer1_outputs(2852);
    layer2_outputs(4386) <= not((layer1_outputs(4467)) or (layer1_outputs(934)));
    layer2_outputs(4387) <= not(layer1_outputs(5539));
    layer2_outputs(4388) <= (layer1_outputs(5636)) or (layer1_outputs(5842));
    layer2_outputs(4389) <= not(layer1_outputs(932)) or (layer1_outputs(900));
    layer2_outputs(4390) <= not((layer1_outputs(3132)) and (layer1_outputs(714)));
    layer2_outputs(4391) <= (layer1_outputs(6261)) or (layer1_outputs(3505));
    layer2_outputs(4392) <= '1';
    layer2_outputs(4393) <= layer1_outputs(2397);
    layer2_outputs(4394) <= not(layer1_outputs(6144));
    layer2_outputs(4395) <= (layer1_outputs(7241)) and (layer1_outputs(6315));
    layer2_outputs(4396) <= (layer1_outputs(1928)) and not (layer1_outputs(513));
    layer2_outputs(4397) <= not(layer1_outputs(4375));
    layer2_outputs(4398) <= not(layer1_outputs(3846));
    layer2_outputs(4399) <= not(layer1_outputs(1018)) or (layer1_outputs(5754));
    layer2_outputs(4400) <= layer1_outputs(5838);
    layer2_outputs(4401) <= not(layer1_outputs(3594));
    layer2_outputs(4402) <= layer1_outputs(2889);
    layer2_outputs(4403) <= layer1_outputs(2276);
    layer2_outputs(4404) <= not(layer1_outputs(1885));
    layer2_outputs(4405) <= layer1_outputs(805);
    layer2_outputs(4406) <= '0';
    layer2_outputs(4407) <= not(layer1_outputs(4656));
    layer2_outputs(4408) <= layer1_outputs(2903);
    layer2_outputs(4409) <= not((layer1_outputs(670)) xor (layer1_outputs(5032)));
    layer2_outputs(4410) <= '1';
    layer2_outputs(4411) <= not(layer1_outputs(4571)) or (layer1_outputs(668));
    layer2_outputs(4412) <= not(layer1_outputs(4435));
    layer2_outputs(4413) <= not(layer1_outputs(3378)) or (layer1_outputs(2601));
    layer2_outputs(4414) <= not(layer1_outputs(6749));
    layer2_outputs(4415) <= not(layer1_outputs(2422));
    layer2_outputs(4416) <= layer1_outputs(7076);
    layer2_outputs(4417) <= layer1_outputs(6527);
    layer2_outputs(4418) <= not(layer1_outputs(3847)) or (layer1_outputs(1444));
    layer2_outputs(4419) <= not((layer1_outputs(5312)) or (layer1_outputs(2015)));
    layer2_outputs(4420) <= not((layer1_outputs(4126)) xor (layer1_outputs(2519)));
    layer2_outputs(4421) <= not(layer1_outputs(7675));
    layer2_outputs(4422) <= not(layer1_outputs(2962)) or (layer1_outputs(2953));
    layer2_outputs(4423) <= not(layer1_outputs(6966));
    layer2_outputs(4424) <= (layer1_outputs(6597)) or (layer1_outputs(3762));
    layer2_outputs(4425) <= (layer1_outputs(2579)) and not (layer1_outputs(4797));
    layer2_outputs(4426) <= '1';
    layer2_outputs(4427) <= layer1_outputs(3540);
    layer2_outputs(4428) <= not(layer1_outputs(231));
    layer2_outputs(4429) <= not((layer1_outputs(4658)) and (layer1_outputs(4524)));
    layer2_outputs(4430) <= not(layer1_outputs(1207));
    layer2_outputs(4431) <= (layer1_outputs(4148)) and not (layer1_outputs(353));
    layer2_outputs(4432) <= not(layer1_outputs(5801));
    layer2_outputs(4433) <= not(layer1_outputs(5228));
    layer2_outputs(4434) <= not(layer1_outputs(4831));
    layer2_outputs(4435) <= layer1_outputs(2262);
    layer2_outputs(4436) <= not(layer1_outputs(6155)) or (layer1_outputs(5696));
    layer2_outputs(4437) <= '1';
    layer2_outputs(4438) <= not((layer1_outputs(165)) and (layer1_outputs(722)));
    layer2_outputs(4439) <= (layer1_outputs(2922)) and not (layer1_outputs(5430));
    layer2_outputs(4440) <= not(layer1_outputs(2799)) or (layer1_outputs(5355));
    layer2_outputs(4441) <= (layer1_outputs(2768)) and not (layer1_outputs(3236));
    layer2_outputs(4442) <= (layer1_outputs(3200)) xor (layer1_outputs(5005));
    layer2_outputs(4443) <= not(layer1_outputs(2525));
    layer2_outputs(4444) <= layer1_outputs(6111);
    layer2_outputs(4445) <= not((layer1_outputs(4295)) and (layer1_outputs(1237)));
    layer2_outputs(4446) <= not(layer1_outputs(5710));
    layer2_outputs(4447) <= not(layer1_outputs(4948));
    layer2_outputs(4448) <= layer1_outputs(3626);
    layer2_outputs(4449) <= not(layer1_outputs(1136)) or (layer1_outputs(4140));
    layer2_outputs(4450) <= not(layer1_outputs(614));
    layer2_outputs(4451) <= not((layer1_outputs(2251)) xor (layer1_outputs(7216)));
    layer2_outputs(4452) <= not(layer1_outputs(6902));
    layer2_outputs(4453) <= layer1_outputs(4366);
    layer2_outputs(4454) <= layer1_outputs(1055);
    layer2_outputs(4455) <= not(layer1_outputs(6337)) or (layer1_outputs(6200));
    layer2_outputs(4456) <= not((layer1_outputs(3092)) or (layer1_outputs(3884)));
    layer2_outputs(4457) <= layer1_outputs(1637);
    layer2_outputs(4458) <= (layer1_outputs(2470)) or (layer1_outputs(3881));
    layer2_outputs(4459) <= not(layer1_outputs(7003));
    layer2_outputs(4460) <= not(layer1_outputs(1210)) or (layer1_outputs(4766));
    layer2_outputs(4461) <= layer1_outputs(5486);
    layer2_outputs(4462) <= not(layer1_outputs(3697));
    layer2_outputs(4463) <= not((layer1_outputs(1506)) xor (layer1_outputs(1430)));
    layer2_outputs(4464) <= (layer1_outputs(3322)) and not (layer1_outputs(1970));
    layer2_outputs(4465) <= (layer1_outputs(3556)) and not (layer1_outputs(4202));
    layer2_outputs(4466) <= not(layer1_outputs(5772)) or (layer1_outputs(3046));
    layer2_outputs(4467) <= not((layer1_outputs(4662)) or (layer1_outputs(7541)));
    layer2_outputs(4468) <= (layer1_outputs(679)) and (layer1_outputs(7132));
    layer2_outputs(4469) <= '1';
    layer2_outputs(4470) <= not((layer1_outputs(7383)) or (layer1_outputs(2061)));
    layer2_outputs(4471) <= layer1_outputs(3746);
    layer2_outputs(4472) <= '0';
    layer2_outputs(4473) <= layer1_outputs(1404);
    layer2_outputs(4474) <= not(layer1_outputs(6244));
    layer2_outputs(4475) <= not(layer1_outputs(130));
    layer2_outputs(4476) <= '1';
    layer2_outputs(4477) <= not(layer1_outputs(3359)) or (layer1_outputs(1173));
    layer2_outputs(4478) <= (layer1_outputs(1716)) or (layer1_outputs(6052));
    layer2_outputs(4479) <= (layer1_outputs(425)) and (layer1_outputs(3380));
    layer2_outputs(4480) <= (layer1_outputs(3858)) and not (layer1_outputs(6462));
    layer2_outputs(4481) <= not((layer1_outputs(5676)) xor (layer1_outputs(3674)));
    layer2_outputs(4482) <= not(layer1_outputs(1916));
    layer2_outputs(4483) <= '0';
    layer2_outputs(4484) <= (layer1_outputs(233)) and not (layer1_outputs(3083));
    layer2_outputs(4485) <= not(layer1_outputs(4851)) or (layer1_outputs(6861));
    layer2_outputs(4486) <= layer1_outputs(2197);
    layer2_outputs(4487) <= not(layer1_outputs(2921));
    layer2_outputs(4488) <= layer1_outputs(6157);
    layer2_outputs(4489) <= (layer1_outputs(2603)) and not (layer1_outputs(5596));
    layer2_outputs(4490) <= not((layer1_outputs(6327)) and (layer1_outputs(1228)));
    layer2_outputs(4491) <= '1';
    layer2_outputs(4492) <= not(layer1_outputs(5901));
    layer2_outputs(4493) <= not((layer1_outputs(6792)) or (layer1_outputs(2563)));
    layer2_outputs(4494) <= not((layer1_outputs(1451)) xor (layer1_outputs(4971)));
    layer2_outputs(4495) <= layer1_outputs(5579);
    layer2_outputs(4496) <= '1';
    layer2_outputs(4497) <= layer1_outputs(3423);
    layer2_outputs(4498) <= not((layer1_outputs(1305)) and (layer1_outputs(6233)));
    layer2_outputs(4499) <= not((layer1_outputs(5956)) and (layer1_outputs(2314)));
    layer2_outputs(4500) <= not((layer1_outputs(4943)) or (layer1_outputs(5125)));
    layer2_outputs(4501) <= (layer1_outputs(1542)) or (layer1_outputs(7398));
    layer2_outputs(4502) <= (layer1_outputs(5341)) and not (layer1_outputs(5826));
    layer2_outputs(4503) <= (layer1_outputs(1570)) and not (layer1_outputs(4678));
    layer2_outputs(4504) <= not((layer1_outputs(7083)) and (layer1_outputs(3322)));
    layer2_outputs(4505) <= (layer1_outputs(2444)) and (layer1_outputs(1516));
    layer2_outputs(4506) <= not((layer1_outputs(4979)) and (layer1_outputs(4377)));
    layer2_outputs(4507) <= not(layer1_outputs(2716));
    layer2_outputs(4508) <= (layer1_outputs(6355)) or (layer1_outputs(4937));
    layer2_outputs(4509) <= layer1_outputs(6387);
    layer2_outputs(4510) <= layer1_outputs(5441);
    layer2_outputs(4511) <= (layer1_outputs(4674)) and (layer1_outputs(1829));
    layer2_outputs(4512) <= (layer1_outputs(2685)) and not (layer1_outputs(7230));
    layer2_outputs(4513) <= layer1_outputs(6034);
    layer2_outputs(4514) <= '1';
    layer2_outputs(4515) <= layer1_outputs(2523);
    layer2_outputs(4516) <= (layer1_outputs(1872)) and not (layer1_outputs(1967));
    layer2_outputs(4517) <= not(layer1_outputs(149));
    layer2_outputs(4518) <= layer1_outputs(3491);
    layer2_outputs(4519) <= (layer1_outputs(2547)) and not (layer1_outputs(2312));
    layer2_outputs(4520) <= layer1_outputs(6614);
    layer2_outputs(4521) <= (layer1_outputs(7617)) or (layer1_outputs(7592));
    layer2_outputs(4522) <= (layer1_outputs(6923)) and (layer1_outputs(645));
    layer2_outputs(4523) <= not(layer1_outputs(4661));
    layer2_outputs(4524) <= not(layer1_outputs(817));
    layer2_outputs(4525) <= not(layer1_outputs(1311));
    layer2_outputs(4526) <= (layer1_outputs(4492)) and not (layer1_outputs(6622));
    layer2_outputs(4527) <= not(layer1_outputs(6580)) or (layer1_outputs(4523));
    layer2_outputs(4528) <= (layer1_outputs(7641)) xor (layer1_outputs(289));
    layer2_outputs(4529) <= '0';
    layer2_outputs(4530) <= (layer1_outputs(2145)) or (layer1_outputs(3997));
    layer2_outputs(4531) <= not(layer1_outputs(620));
    layer2_outputs(4532) <= (layer1_outputs(1824)) and not (layer1_outputs(2545));
    layer2_outputs(4533) <= not((layer1_outputs(6545)) xor (layer1_outputs(226)));
    layer2_outputs(4534) <= (layer1_outputs(6492)) and not (layer1_outputs(2119));
    layer2_outputs(4535) <= layer1_outputs(2637);
    layer2_outputs(4536) <= not(layer1_outputs(5541)) or (layer1_outputs(2365));
    layer2_outputs(4537) <= not(layer1_outputs(6805));
    layer2_outputs(4538) <= not((layer1_outputs(5498)) and (layer1_outputs(7099)));
    layer2_outputs(4539) <= not((layer1_outputs(1726)) and (layer1_outputs(821)));
    layer2_outputs(4540) <= not(layer1_outputs(1221));
    layer2_outputs(4541) <= not((layer1_outputs(4555)) xor (layer1_outputs(7149)));
    layer2_outputs(4542) <= not(layer1_outputs(7430));
    layer2_outputs(4543) <= layer1_outputs(3636);
    layer2_outputs(4544) <= not(layer1_outputs(7466)) or (layer1_outputs(1835));
    layer2_outputs(4545) <= not(layer1_outputs(7451)) or (layer1_outputs(6995));
    layer2_outputs(4546) <= not((layer1_outputs(2515)) and (layer1_outputs(7303)));
    layer2_outputs(4547) <= not((layer1_outputs(4649)) or (layer1_outputs(1371)));
    layer2_outputs(4548) <= not(layer1_outputs(259)) or (layer1_outputs(5917));
    layer2_outputs(4549) <= not(layer1_outputs(7339));
    layer2_outputs(4550) <= not(layer1_outputs(1195));
    layer2_outputs(4551) <= not(layer1_outputs(5848));
    layer2_outputs(4552) <= not((layer1_outputs(403)) or (layer1_outputs(1798)));
    layer2_outputs(4553) <= layer1_outputs(2746);
    layer2_outputs(4554) <= layer1_outputs(2206);
    layer2_outputs(4555) <= not(layer1_outputs(3679));
    layer2_outputs(4556) <= (layer1_outputs(2670)) and not (layer1_outputs(1285));
    layer2_outputs(4557) <= (layer1_outputs(4209)) and not (layer1_outputs(747));
    layer2_outputs(4558) <= (layer1_outputs(4991)) and not (layer1_outputs(6111));
    layer2_outputs(4559) <= layer1_outputs(231);
    layer2_outputs(4560) <= not(layer1_outputs(2219));
    layer2_outputs(4561) <= not((layer1_outputs(1591)) or (layer1_outputs(5787)));
    layer2_outputs(4562) <= not(layer1_outputs(100));
    layer2_outputs(4563) <= '1';
    layer2_outputs(4564) <= (layer1_outputs(6388)) and (layer1_outputs(2216));
    layer2_outputs(4565) <= layer1_outputs(2377);
    layer2_outputs(4566) <= (layer1_outputs(2619)) and (layer1_outputs(6005));
    layer2_outputs(4567) <= '0';
    layer2_outputs(4568) <= not((layer1_outputs(4100)) or (layer1_outputs(1356)));
    layer2_outputs(4569) <= layer1_outputs(876);
    layer2_outputs(4570) <= not(layer1_outputs(3711));
    layer2_outputs(4571) <= not(layer1_outputs(987)) or (layer1_outputs(6091));
    layer2_outputs(4572) <= (layer1_outputs(1101)) and not (layer1_outputs(2387));
    layer2_outputs(4573) <= not(layer1_outputs(5002)) or (layer1_outputs(6888));
    layer2_outputs(4574) <= not(layer1_outputs(4807)) or (layer1_outputs(441));
    layer2_outputs(4575) <= (layer1_outputs(6602)) and (layer1_outputs(6374));
    layer2_outputs(4576) <= layer1_outputs(4482);
    layer2_outputs(4577) <= layer1_outputs(1005);
    layer2_outputs(4578) <= layer1_outputs(110);
    layer2_outputs(4579) <= not(layer1_outputs(992)) or (layer1_outputs(801));
    layer2_outputs(4580) <= (layer1_outputs(992)) or (layer1_outputs(7552));
    layer2_outputs(4581) <= not(layer1_outputs(3479));
    layer2_outputs(4582) <= not((layer1_outputs(6177)) or (layer1_outputs(7303)));
    layer2_outputs(4583) <= (layer1_outputs(2895)) xor (layer1_outputs(145));
    layer2_outputs(4584) <= not(layer1_outputs(5492)) or (layer1_outputs(42));
    layer2_outputs(4585) <= layer1_outputs(6751);
    layer2_outputs(4586) <= '0';
    layer2_outputs(4587) <= not(layer1_outputs(1867));
    layer2_outputs(4588) <= not(layer1_outputs(126)) or (layer1_outputs(292));
    layer2_outputs(4589) <= (layer1_outputs(7335)) xor (layer1_outputs(1703));
    layer2_outputs(4590) <= not(layer1_outputs(1826)) or (layer1_outputs(7166));
    layer2_outputs(4591) <= layer1_outputs(5923);
    layer2_outputs(4592) <= not(layer1_outputs(4449));
    layer2_outputs(4593) <= (layer1_outputs(5644)) or (layer1_outputs(3712));
    layer2_outputs(4594) <= not(layer1_outputs(2832));
    layer2_outputs(4595) <= (layer1_outputs(2239)) and (layer1_outputs(1706));
    layer2_outputs(4596) <= layer1_outputs(3693);
    layer2_outputs(4597) <= (layer1_outputs(361)) and (layer1_outputs(1602));
    layer2_outputs(4598) <= not(layer1_outputs(3106));
    layer2_outputs(4599) <= not((layer1_outputs(3521)) and (layer1_outputs(2376)));
    layer2_outputs(4600) <= (layer1_outputs(2226)) or (layer1_outputs(6451));
    layer2_outputs(4601) <= '1';
    layer2_outputs(4602) <= not((layer1_outputs(4015)) and (layer1_outputs(3450)));
    layer2_outputs(4603) <= not((layer1_outputs(4812)) xor (layer1_outputs(6599)));
    layer2_outputs(4604) <= (layer1_outputs(2304)) or (layer1_outputs(5003));
    layer2_outputs(4605) <= not((layer1_outputs(3967)) and (layer1_outputs(1076)));
    layer2_outputs(4606) <= (layer1_outputs(7242)) and not (layer1_outputs(6892));
    layer2_outputs(4607) <= '1';
    layer2_outputs(4608) <= not(layer1_outputs(3848)) or (layer1_outputs(33));
    layer2_outputs(4609) <= (layer1_outputs(3993)) and (layer1_outputs(434));
    layer2_outputs(4610) <= not(layer1_outputs(5449));
    layer2_outputs(4611) <= (layer1_outputs(450)) or (layer1_outputs(3489));
    layer2_outputs(4612) <= (layer1_outputs(4094)) and not (layer1_outputs(3118));
    layer2_outputs(4613) <= layer1_outputs(5951);
    layer2_outputs(4614) <= layer1_outputs(4059);
    layer2_outputs(4615) <= (layer1_outputs(6070)) and (layer1_outputs(6742));
    layer2_outputs(4616) <= (layer1_outputs(794)) and not (layer1_outputs(2475));
    layer2_outputs(4617) <= not(layer1_outputs(3809));
    layer2_outputs(4618) <= '1';
    layer2_outputs(4619) <= not((layer1_outputs(5476)) or (layer1_outputs(4612)));
    layer2_outputs(4620) <= not(layer1_outputs(4673)) or (layer1_outputs(2009));
    layer2_outputs(4621) <= not(layer1_outputs(7157)) or (layer1_outputs(973));
    layer2_outputs(4622) <= not(layer1_outputs(6452));
    layer2_outputs(4623) <= (layer1_outputs(5982)) or (layer1_outputs(5820));
    layer2_outputs(4624) <= layer1_outputs(2247);
    layer2_outputs(4625) <= layer1_outputs(2554);
    layer2_outputs(4626) <= not(layer1_outputs(380));
    layer2_outputs(4627) <= '0';
    layer2_outputs(4628) <= not(layer1_outputs(2388)) or (layer1_outputs(891));
    layer2_outputs(4629) <= not((layer1_outputs(5824)) or (layer1_outputs(5103)));
    layer2_outputs(4630) <= not((layer1_outputs(4022)) and (layer1_outputs(6448)));
    layer2_outputs(4631) <= not(layer1_outputs(5154));
    layer2_outputs(4632) <= (layer1_outputs(4641)) and (layer1_outputs(4182));
    layer2_outputs(4633) <= layer1_outputs(2638);
    layer2_outputs(4634) <= (layer1_outputs(7429)) and not (layer1_outputs(7306));
    layer2_outputs(4635) <= (layer1_outputs(7572)) and not (layer1_outputs(5986));
    layer2_outputs(4636) <= layer1_outputs(3350);
    layer2_outputs(4637) <= (layer1_outputs(5750)) xor (layer1_outputs(6076));
    layer2_outputs(4638) <= (layer1_outputs(2382)) and (layer1_outputs(2386));
    layer2_outputs(4639) <= (layer1_outputs(1433)) or (layer1_outputs(6141));
    layer2_outputs(4640) <= (layer1_outputs(1742)) and not (layer1_outputs(7299));
    layer2_outputs(4641) <= not(layer1_outputs(1980));
    layer2_outputs(4642) <= not(layer1_outputs(5690)) or (layer1_outputs(1180));
    layer2_outputs(4643) <= layer1_outputs(6975);
    layer2_outputs(4644) <= '1';
    layer2_outputs(4645) <= (layer1_outputs(1460)) and not (layer1_outputs(4833));
    layer2_outputs(4646) <= (layer1_outputs(215)) and not (layer1_outputs(4895));
    layer2_outputs(4647) <= layer1_outputs(6776);
    layer2_outputs(4648) <= not(layer1_outputs(4892)) or (layer1_outputs(5154));
    layer2_outputs(4649) <= not(layer1_outputs(2146)) or (layer1_outputs(5416));
    layer2_outputs(4650) <= '0';
    layer2_outputs(4651) <= layer1_outputs(1504);
    layer2_outputs(4652) <= not(layer1_outputs(241)) or (layer1_outputs(1476));
    layer2_outputs(4653) <= not((layer1_outputs(3063)) or (layer1_outputs(7275)));
    layer2_outputs(4654) <= layer1_outputs(4268);
    layer2_outputs(4655) <= not(layer1_outputs(1039));
    layer2_outputs(4656) <= '0';
    layer2_outputs(4657) <= (layer1_outputs(7171)) and (layer1_outputs(2796));
    layer2_outputs(4658) <= not(layer1_outputs(7001));
    layer2_outputs(4659) <= (layer1_outputs(3428)) xor (layer1_outputs(404));
    layer2_outputs(4660) <= layer1_outputs(2917);
    layer2_outputs(4661) <= not(layer1_outputs(6450));
    layer2_outputs(4662) <= not(layer1_outputs(5265)) or (layer1_outputs(6923));
    layer2_outputs(4663) <= not((layer1_outputs(1785)) or (layer1_outputs(5428)));
    layer2_outputs(4664) <= (layer1_outputs(3266)) or (layer1_outputs(2217));
    layer2_outputs(4665) <= layer1_outputs(5871);
    layer2_outputs(4666) <= layer1_outputs(4198);
    layer2_outputs(4667) <= not((layer1_outputs(4676)) and (layer1_outputs(5544)));
    layer2_outputs(4668) <= not(layer1_outputs(4435));
    layer2_outputs(4669) <= layer1_outputs(1293);
    layer2_outputs(4670) <= (layer1_outputs(1144)) and (layer1_outputs(7179));
    layer2_outputs(4671) <= (layer1_outputs(4824)) and not (layer1_outputs(7106));
    layer2_outputs(4672) <= (layer1_outputs(3011)) and (layer1_outputs(2485));
    layer2_outputs(4673) <= (layer1_outputs(5855)) and (layer1_outputs(6163));
    layer2_outputs(4674) <= layer1_outputs(2428);
    layer2_outputs(4675) <= not((layer1_outputs(844)) or (layer1_outputs(5680)));
    layer2_outputs(4676) <= layer1_outputs(1061);
    layer2_outputs(4677) <= (layer1_outputs(538)) and not (layer1_outputs(2868));
    layer2_outputs(4678) <= not((layer1_outputs(5802)) or (layer1_outputs(4834)));
    layer2_outputs(4679) <= (layer1_outputs(85)) and (layer1_outputs(3641));
    layer2_outputs(4680) <= '0';
    layer2_outputs(4681) <= (layer1_outputs(3475)) and not (layer1_outputs(6637));
    layer2_outputs(4682) <= layer1_outputs(2588);
    layer2_outputs(4683) <= not(layer1_outputs(2799)) or (layer1_outputs(4154));
    layer2_outputs(4684) <= not(layer1_outputs(5096)) or (layer1_outputs(7086));
    layer2_outputs(4685) <= layer1_outputs(946);
    layer2_outputs(4686) <= not(layer1_outputs(5255));
    layer2_outputs(4687) <= layer1_outputs(6769);
    layer2_outputs(4688) <= not(layer1_outputs(3126));
    layer2_outputs(4689) <= (layer1_outputs(2909)) and not (layer1_outputs(4316));
    layer2_outputs(4690) <= layer1_outputs(6009);
    layer2_outputs(4691) <= (layer1_outputs(1659)) or (layer1_outputs(5237));
    layer2_outputs(4692) <= layer1_outputs(4506);
    layer2_outputs(4693) <= layer1_outputs(2992);
    layer2_outputs(4694) <= (layer1_outputs(1368)) and (layer1_outputs(2851));
    layer2_outputs(4695) <= layer1_outputs(5358);
    layer2_outputs(4696) <= not(layer1_outputs(7378)) or (layer1_outputs(6387));
    layer2_outputs(4697) <= not((layer1_outputs(4550)) or (layer1_outputs(3188)));
    layer2_outputs(4698) <= layer1_outputs(7027);
    layer2_outputs(4699) <= layer1_outputs(5038);
    layer2_outputs(4700) <= not(layer1_outputs(4361)) or (layer1_outputs(1182));
    layer2_outputs(4701) <= '1';
    layer2_outputs(4702) <= layer1_outputs(1053);
    layer2_outputs(4703) <= layer1_outputs(3081);
    layer2_outputs(4704) <= not((layer1_outputs(4266)) or (layer1_outputs(5087)));
    layer2_outputs(4705) <= not(layer1_outputs(1330));
    layer2_outputs(4706) <= not(layer1_outputs(857));
    layer2_outputs(4707) <= not((layer1_outputs(3347)) or (layer1_outputs(1593)));
    layer2_outputs(4708) <= (layer1_outputs(3694)) and not (layer1_outputs(3013));
    layer2_outputs(4709) <= layer1_outputs(3386);
    layer2_outputs(4710) <= not(layer1_outputs(6701));
    layer2_outputs(4711) <= layer1_outputs(4371);
    layer2_outputs(4712) <= '0';
    layer2_outputs(4713) <= layer1_outputs(2480);
    layer2_outputs(4714) <= not((layer1_outputs(1658)) xor (layer1_outputs(6788)));
    layer2_outputs(4715) <= not(layer1_outputs(6239));
    layer2_outputs(4716) <= layer1_outputs(5712);
    layer2_outputs(4717) <= layer1_outputs(141);
    layer2_outputs(4718) <= not((layer1_outputs(2555)) and (layer1_outputs(1169)));
    layer2_outputs(4719) <= (layer1_outputs(2649)) and not (layer1_outputs(6218));
    layer2_outputs(4720) <= layer1_outputs(7362);
    layer2_outputs(4721) <= not(layer1_outputs(342));
    layer2_outputs(4722) <= (layer1_outputs(3873)) and (layer1_outputs(4648));
    layer2_outputs(4723) <= not((layer1_outputs(5167)) and (layer1_outputs(13)));
    layer2_outputs(4724) <= not(layer1_outputs(6533));
    layer2_outputs(4725) <= (layer1_outputs(495)) and not (layer1_outputs(5918));
    layer2_outputs(4726) <= not(layer1_outputs(840)) or (layer1_outputs(855));
    layer2_outputs(4727) <= layer1_outputs(4549);
    layer2_outputs(4728) <= layer1_outputs(7038);
    layer2_outputs(4729) <= (layer1_outputs(4283)) or (layer1_outputs(737));
    layer2_outputs(4730) <= not((layer1_outputs(5175)) xor (layer1_outputs(5057)));
    layer2_outputs(4731) <= (layer1_outputs(2859)) and not (layer1_outputs(1444));
    layer2_outputs(4732) <= not(layer1_outputs(3358)) or (layer1_outputs(6484));
    layer2_outputs(4733) <= layer1_outputs(1199);
    layer2_outputs(4734) <= not(layer1_outputs(4632));
    layer2_outputs(4735) <= (layer1_outputs(3346)) or (layer1_outputs(531));
    layer2_outputs(4736) <= layer1_outputs(7062);
    layer2_outputs(4737) <= '1';
    layer2_outputs(4738) <= not(layer1_outputs(5890));
    layer2_outputs(4739) <= (layer1_outputs(2681)) and (layer1_outputs(2773));
    layer2_outputs(4740) <= not(layer1_outputs(1400));
    layer2_outputs(4741) <= not(layer1_outputs(7067));
    layer2_outputs(4742) <= (layer1_outputs(7393)) or (layer1_outputs(4635));
    layer2_outputs(4743) <= (layer1_outputs(4940)) and not (layer1_outputs(3473));
    layer2_outputs(4744) <= (layer1_outputs(1522)) or (layer1_outputs(3720));
    layer2_outputs(4745) <= layer1_outputs(4793);
    layer2_outputs(4746) <= not(layer1_outputs(6925)) or (layer1_outputs(3087));
    layer2_outputs(4747) <= layer1_outputs(5571);
    layer2_outputs(4748) <= not(layer1_outputs(3119));
    layer2_outputs(4749) <= (layer1_outputs(6992)) and (layer1_outputs(1636));
    layer2_outputs(4750) <= not(layer1_outputs(820));
    layer2_outputs(4751) <= not((layer1_outputs(6425)) and (layer1_outputs(3017)));
    layer2_outputs(4752) <= not(layer1_outputs(6260)) or (layer1_outputs(5201));
    layer2_outputs(4753) <= layer1_outputs(7537);
    layer2_outputs(4754) <= (layer1_outputs(251)) and not (layer1_outputs(5141));
    layer2_outputs(4755) <= layer1_outputs(6843);
    layer2_outputs(4756) <= layer1_outputs(5440);
    layer2_outputs(4757) <= (layer1_outputs(27)) and not (layer1_outputs(4004));
    layer2_outputs(4758) <= (layer1_outputs(4147)) and not (layer1_outputs(6238));
    layer2_outputs(4759) <= not((layer1_outputs(5212)) and (layer1_outputs(6188)));
    layer2_outputs(4760) <= not((layer1_outputs(6998)) or (layer1_outputs(7156)));
    layer2_outputs(4761) <= layer1_outputs(1344);
    layer2_outputs(4762) <= (layer1_outputs(275)) and (layer1_outputs(502));
    layer2_outputs(4763) <= not(layer1_outputs(6990));
    layer2_outputs(4764) <= layer1_outputs(289);
    layer2_outputs(4765) <= not((layer1_outputs(3635)) and (layer1_outputs(4741)));
    layer2_outputs(4766) <= not((layer1_outputs(7586)) or (layer1_outputs(1712)));
    layer2_outputs(4767) <= layer1_outputs(1828);
    layer2_outputs(4768) <= layer1_outputs(2294);
    layer2_outputs(4769) <= not(layer1_outputs(2389));
    layer2_outputs(4770) <= (layer1_outputs(2373)) or (layer1_outputs(6247));
    layer2_outputs(4771) <= (layer1_outputs(1711)) and not (layer1_outputs(7566));
    layer2_outputs(4772) <= not(layer1_outputs(2872));
    layer2_outputs(4773) <= layer1_outputs(2956);
    layer2_outputs(4774) <= layer1_outputs(7346);
    layer2_outputs(4775) <= '1';
    layer2_outputs(4776) <= not(layer1_outputs(7278)) or (layer1_outputs(5678));
    layer2_outputs(4777) <= not((layer1_outputs(6249)) and (layer1_outputs(5851)));
    layer2_outputs(4778) <= not((layer1_outputs(5693)) and (layer1_outputs(2674)));
    layer2_outputs(4779) <= not(layer1_outputs(3350)) or (layer1_outputs(7373));
    layer2_outputs(4780) <= layer1_outputs(4748);
    layer2_outputs(4781) <= not(layer1_outputs(6914)) or (layer1_outputs(5862));
    layer2_outputs(4782) <= not((layer1_outputs(1242)) or (layer1_outputs(3075)));
    layer2_outputs(4783) <= not(layer1_outputs(2001));
    layer2_outputs(4784) <= (layer1_outputs(5010)) and not (layer1_outputs(4728));
    layer2_outputs(4785) <= (layer1_outputs(3370)) or (layer1_outputs(3961));
    layer2_outputs(4786) <= not(layer1_outputs(6818)) or (layer1_outputs(708));
    layer2_outputs(4787) <= not(layer1_outputs(5904)) or (layer1_outputs(6013));
    layer2_outputs(4788) <= (layer1_outputs(6406)) and (layer1_outputs(5972));
    layer2_outputs(4789) <= not(layer1_outputs(1937));
    layer2_outputs(4790) <= '1';
    layer2_outputs(4791) <= (layer1_outputs(5692)) and (layer1_outputs(6021));
    layer2_outputs(4792) <= '1';
    layer2_outputs(4793) <= (layer1_outputs(7315)) and (layer1_outputs(243));
    layer2_outputs(4794) <= (layer1_outputs(3169)) and (layer1_outputs(1710));
    layer2_outputs(4795) <= not(layer1_outputs(6775));
    layer2_outputs(4796) <= '0';
    layer2_outputs(4797) <= layer1_outputs(7232);
    layer2_outputs(4798) <= not((layer1_outputs(4748)) xor (layer1_outputs(4560)));
    layer2_outputs(4799) <= not(layer1_outputs(2746));
    layer2_outputs(4800) <= not(layer1_outputs(3923));
    layer2_outputs(4801) <= not(layer1_outputs(3761));
    layer2_outputs(4802) <= '0';
    layer2_outputs(4803) <= (layer1_outputs(3289)) or (layer1_outputs(1686));
    layer2_outputs(4804) <= (layer1_outputs(6102)) and not (layer1_outputs(4578));
    layer2_outputs(4805) <= not(layer1_outputs(3299));
    layer2_outputs(4806) <= not(layer1_outputs(7482));
    layer2_outputs(4807) <= (layer1_outputs(6517)) and not (layer1_outputs(4897));
    layer2_outputs(4808) <= (layer1_outputs(7194)) and not (layer1_outputs(6212));
    layer2_outputs(4809) <= layer1_outputs(3193);
    layer2_outputs(4810) <= (layer1_outputs(4669)) or (layer1_outputs(277));
    layer2_outputs(4811) <= not(layer1_outputs(861));
    layer2_outputs(4812) <= not(layer1_outputs(371));
    layer2_outputs(4813) <= layer1_outputs(3912);
    layer2_outputs(4814) <= not((layer1_outputs(5717)) and (layer1_outputs(5249)));
    layer2_outputs(4815) <= layer1_outputs(1113);
    layer2_outputs(4816) <= not((layer1_outputs(605)) or (layer1_outputs(4799)));
    layer2_outputs(4817) <= '1';
    layer2_outputs(4818) <= not((layer1_outputs(4236)) and (layer1_outputs(1647)));
    layer2_outputs(4819) <= not(layer1_outputs(4210));
    layer2_outputs(4820) <= not((layer1_outputs(3291)) xor (layer1_outputs(2813)));
    layer2_outputs(4821) <= (layer1_outputs(1827)) and not (layer1_outputs(4314));
    layer2_outputs(4822) <= (layer1_outputs(7235)) and not (layer1_outputs(1314));
    layer2_outputs(4823) <= '0';
    layer2_outputs(4824) <= not(layer1_outputs(6617)) or (layer1_outputs(7468));
    layer2_outputs(4825) <= (layer1_outputs(5807)) and not (layer1_outputs(2264));
    layer2_outputs(4826) <= not(layer1_outputs(577));
    layer2_outputs(4827) <= not((layer1_outputs(4653)) xor (layer1_outputs(6553)));
    layer2_outputs(4828) <= layer1_outputs(4988);
    layer2_outputs(4829) <= layer1_outputs(4558);
    layer2_outputs(4830) <= (layer1_outputs(1140)) and (layer1_outputs(5788));
    layer2_outputs(4831) <= layer1_outputs(746);
    layer2_outputs(4832) <= layer1_outputs(6862);
    layer2_outputs(4833) <= not(layer1_outputs(2367));
    layer2_outputs(4834) <= not((layer1_outputs(2040)) and (layer1_outputs(1810)));
    layer2_outputs(4835) <= not((layer1_outputs(4058)) xor (layer1_outputs(5195)));
    layer2_outputs(4836) <= '0';
    layer2_outputs(4837) <= not((layer1_outputs(3102)) or (layer1_outputs(2873)));
    layer2_outputs(4838) <= (layer1_outputs(537)) and (layer1_outputs(4631));
    layer2_outputs(4839) <= layer1_outputs(4902);
    layer2_outputs(4840) <= not(layer1_outputs(1213));
    layer2_outputs(4841) <= layer1_outputs(1319);
    layer2_outputs(4842) <= not(layer1_outputs(3332)) or (layer1_outputs(7131));
    layer2_outputs(4843) <= (layer1_outputs(4083)) and not (layer1_outputs(6567));
    layer2_outputs(4844) <= not(layer1_outputs(1720));
    layer2_outputs(4845) <= not(layer1_outputs(2043));
    layer2_outputs(4846) <= layer1_outputs(5637);
    layer2_outputs(4847) <= (layer1_outputs(1461)) and not (layer1_outputs(1350));
    layer2_outputs(4848) <= not(layer1_outputs(4336));
    layer2_outputs(4849) <= not(layer1_outputs(7267));
    layer2_outputs(4850) <= (layer1_outputs(2111)) and (layer1_outputs(1442));
    layer2_outputs(4851) <= not(layer1_outputs(1740));
    layer2_outputs(4852) <= (layer1_outputs(5070)) or (layer1_outputs(981));
    layer2_outputs(4853) <= '1';
    layer2_outputs(4854) <= (layer1_outputs(4260)) and (layer1_outputs(135));
    layer2_outputs(4855) <= (layer1_outputs(3732)) or (layer1_outputs(4752));
    layer2_outputs(4856) <= not((layer1_outputs(2138)) or (layer1_outputs(4055)));
    layer2_outputs(4857) <= not(layer1_outputs(586));
    layer2_outputs(4858) <= not(layer1_outputs(5935));
    layer2_outputs(4859) <= layer1_outputs(4888);
    layer2_outputs(4860) <= (layer1_outputs(3114)) xor (layer1_outputs(2791));
    layer2_outputs(4861) <= (layer1_outputs(5977)) and not (layer1_outputs(2526));
    layer2_outputs(4862) <= '0';
    layer2_outputs(4863) <= '1';
    layer2_outputs(4864) <= (layer1_outputs(4946)) or (layer1_outputs(7037));
    layer2_outputs(4865) <= not(layer1_outputs(6735));
    layer2_outputs(4866) <= not(layer1_outputs(3124));
    layer2_outputs(4867) <= layer1_outputs(236);
    layer2_outputs(4868) <= '0';
    layer2_outputs(4869) <= (layer1_outputs(4042)) and (layer1_outputs(4373));
    layer2_outputs(4870) <= not(layer1_outputs(9));
    layer2_outputs(4871) <= not(layer1_outputs(6037));
    layer2_outputs(4872) <= not(layer1_outputs(6302));
    layer2_outputs(4873) <= (layer1_outputs(3177)) and (layer1_outputs(7514));
    layer2_outputs(4874) <= not(layer1_outputs(6583)) or (layer1_outputs(7474));
    layer2_outputs(4875) <= layer1_outputs(5574);
    layer2_outputs(4876) <= layer1_outputs(6421);
    layer2_outputs(4877) <= (layer1_outputs(2286)) or (layer1_outputs(3098));
    layer2_outputs(4878) <= not((layer1_outputs(7276)) or (layer1_outputs(3415)));
    layer2_outputs(4879) <= (layer1_outputs(2999)) and (layer1_outputs(1650));
    layer2_outputs(4880) <= (layer1_outputs(6981)) and (layer1_outputs(1156));
    layer2_outputs(4881) <= '0';
    layer2_outputs(4882) <= not(layer1_outputs(2571));
    layer2_outputs(4883) <= layer1_outputs(123);
    layer2_outputs(4884) <= layer1_outputs(2559);
    layer2_outputs(4885) <= not(layer1_outputs(4896));
    layer2_outputs(4886) <= '0';
    layer2_outputs(4887) <= (layer1_outputs(534)) and not (layer1_outputs(5214));
    layer2_outputs(4888) <= not((layer1_outputs(6035)) and (layer1_outputs(6175)));
    layer2_outputs(4889) <= not((layer1_outputs(4618)) and (layer1_outputs(1942)));
    layer2_outputs(4890) <= layer1_outputs(2015);
    layer2_outputs(4891) <= layer1_outputs(6380);
    layer2_outputs(4892) <= (layer1_outputs(3390)) and not (layer1_outputs(4568));
    layer2_outputs(4893) <= (layer1_outputs(6535)) and not (layer1_outputs(4073));
    layer2_outputs(4894) <= layer1_outputs(5338);
    layer2_outputs(4895) <= (layer1_outputs(4584)) and not (layer1_outputs(3927));
    layer2_outputs(4896) <= (layer1_outputs(6866)) and not (layer1_outputs(525));
    layer2_outputs(4897) <= layer1_outputs(2131);
    layer2_outputs(4898) <= not(layer1_outputs(6231));
    layer2_outputs(4899) <= not(layer1_outputs(5607));
    layer2_outputs(4900) <= (layer1_outputs(5528)) and (layer1_outputs(779));
    layer2_outputs(4901) <= layer1_outputs(2878);
    layer2_outputs(4902) <= (layer1_outputs(2826)) and (layer1_outputs(2142));
    layer2_outputs(4903) <= not((layer1_outputs(7257)) or (layer1_outputs(238)));
    layer2_outputs(4904) <= not(layer1_outputs(3926));
    layer2_outputs(4905) <= not(layer1_outputs(1181));
    layer2_outputs(4906) <= not((layer1_outputs(886)) or (layer1_outputs(2297)));
    layer2_outputs(4907) <= not(layer1_outputs(2650));
    layer2_outputs(4908) <= layer1_outputs(5025);
    layer2_outputs(4909) <= not(layer1_outputs(5238)) or (layer1_outputs(2996));
    layer2_outputs(4910) <= layer1_outputs(2215);
    layer2_outputs(4911) <= layer1_outputs(3616);
    layer2_outputs(4912) <= not(layer1_outputs(6466));
    layer2_outputs(4913) <= (layer1_outputs(3667)) or (layer1_outputs(3029));
    layer2_outputs(4914) <= layer1_outputs(7630);
    layer2_outputs(4915) <= layer1_outputs(864);
    layer2_outputs(4916) <= not(layer1_outputs(6557)) or (layer1_outputs(6328));
    layer2_outputs(4917) <= not(layer1_outputs(2071)) or (layer1_outputs(1133));
    layer2_outputs(4918) <= not((layer1_outputs(3396)) and (layer1_outputs(6625)));
    layer2_outputs(4919) <= not(layer1_outputs(3471));
    layer2_outputs(4920) <= not(layer1_outputs(6929));
    layer2_outputs(4921) <= layer1_outputs(5312);
    layer2_outputs(4922) <= not(layer1_outputs(3746)) or (layer1_outputs(3042));
    layer2_outputs(4923) <= not(layer1_outputs(7558)) or (layer1_outputs(4473));
    layer2_outputs(4924) <= layer1_outputs(5070);
    layer2_outputs(4925) <= not(layer1_outputs(4167));
    layer2_outputs(4926) <= (layer1_outputs(811)) and not (layer1_outputs(1023));
    layer2_outputs(4927) <= not((layer1_outputs(4050)) and (layer1_outputs(1353)));
    layer2_outputs(4928) <= not(layer1_outputs(1887));
    layer2_outputs(4929) <= layer1_outputs(1825);
    layer2_outputs(4930) <= layer1_outputs(1359);
    layer2_outputs(4931) <= layer1_outputs(1722);
    layer2_outputs(4932) <= '1';
    layer2_outputs(4933) <= not(layer1_outputs(7615)) or (layer1_outputs(5667));
    layer2_outputs(4934) <= not(layer1_outputs(2624)) or (layer1_outputs(657));
    layer2_outputs(4935) <= layer1_outputs(6740);
    layer2_outputs(4936) <= not(layer1_outputs(7467)) or (layer1_outputs(3431));
    layer2_outputs(4937) <= not((layer1_outputs(4079)) and (layer1_outputs(7279)));
    layer2_outputs(4938) <= not((layer1_outputs(2609)) and (layer1_outputs(2977)));
    layer2_outputs(4939) <= not((layer1_outputs(925)) or (layer1_outputs(5085)));
    layer2_outputs(4940) <= not(layer1_outputs(5175));
    layer2_outputs(4941) <= not(layer1_outputs(5222)) or (layer1_outputs(6834));
    layer2_outputs(4942) <= not(layer1_outputs(3042));
    layer2_outputs(4943) <= not(layer1_outputs(4306)) or (layer1_outputs(724));
    layer2_outputs(4944) <= layer1_outputs(4086);
    layer2_outputs(4945) <= not(layer1_outputs(4159));
    layer2_outputs(4946) <= not(layer1_outputs(6001));
    layer2_outputs(4947) <= layer1_outputs(5405);
    layer2_outputs(4948) <= layer1_outputs(3259);
    layer2_outputs(4949) <= (layer1_outputs(4229)) and not (layer1_outputs(2518));
    layer2_outputs(4950) <= not(layer1_outputs(6565)) or (layer1_outputs(4080));
    layer2_outputs(4951) <= (layer1_outputs(3467)) and not (layer1_outputs(1205));
    layer2_outputs(4952) <= not(layer1_outputs(6812)) or (layer1_outputs(926));
    layer2_outputs(4953) <= '1';
    layer2_outputs(4954) <= '0';
    layer2_outputs(4955) <= not(layer1_outputs(7597));
    layer2_outputs(4956) <= not(layer1_outputs(3928));
    layer2_outputs(4957) <= layer1_outputs(617);
    layer2_outputs(4958) <= layer1_outputs(3686);
    layer2_outputs(4959) <= layer1_outputs(1964);
    layer2_outputs(4960) <= (layer1_outputs(6778)) and not (layer1_outputs(5456));
    layer2_outputs(4961) <= not(layer1_outputs(3364)) or (layer1_outputs(7061));
    layer2_outputs(4962) <= (layer1_outputs(2298)) or (layer1_outputs(6538));
    layer2_outputs(4963) <= not(layer1_outputs(3768)) or (layer1_outputs(4420));
    layer2_outputs(4964) <= not(layer1_outputs(7485));
    layer2_outputs(4965) <= not(layer1_outputs(3587)) or (layer1_outputs(6264));
    layer2_outputs(4966) <= not(layer1_outputs(1890));
    layer2_outputs(4967) <= not((layer1_outputs(3825)) and (layer1_outputs(102)));
    layer2_outputs(4968) <= not(layer1_outputs(6056));
    layer2_outputs(4969) <= not(layer1_outputs(5668));
    layer2_outputs(4970) <= (layer1_outputs(6149)) or (layer1_outputs(6199));
    layer2_outputs(4971) <= '0';
    layer2_outputs(4972) <= not(layer1_outputs(4606));
    layer2_outputs(4973) <= layer1_outputs(312);
    layer2_outputs(4974) <= not((layer1_outputs(5304)) xor (layer1_outputs(6176)));
    layer2_outputs(4975) <= not(layer1_outputs(349));
    layer2_outputs(4976) <= not(layer1_outputs(1919));
    layer2_outputs(4977) <= not(layer1_outputs(4565)) or (layer1_outputs(7495));
    layer2_outputs(4978) <= (layer1_outputs(1957)) and (layer1_outputs(2436));
    layer2_outputs(4979) <= not((layer1_outputs(5345)) xor (layer1_outputs(7525)));
    layer2_outputs(4980) <= '0';
    layer2_outputs(4981) <= not(layer1_outputs(6317));
    layer2_outputs(4982) <= not((layer1_outputs(860)) xor (layer1_outputs(4896)));
    layer2_outputs(4983) <= not((layer1_outputs(3596)) or (layer1_outputs(3053)));
    layer2_outputs(4984) <= not(layer1_outputs(4643));
    layer2_outputs(4985) <= (layer1_outputs(4100)) and not (layer1_outputs(2575));
    layer2_outputs(4986) <= not(layer1_outputs(5146)) or (layer1_outputs(2451));
    layer2_outputs(4987) <= not((layer1_outputs(1407)) or (layer1_outputs(415)));
    layer2_outputs(4988) <= (layer1_outputs(3018)) and not (layer1_outputs(820));
    layer2_outputs(4989) <= (layer1_outputs(595)) and (layer1_outputs(4914));
    layer2_outputs(4990) <= not((layer1_outputs(2983)) and (layer1_outputs(2938)));
    layer2_outputs(4991) <= not(layer1_outputs(4367));
    layer2_outputs(4992) <= layer1_outputs(5926);
    layer2_outputs(4993) <= (layer1_outputs(5206)) or (layer1_outputs(4345));
    layer2_outputs(4994) <= (layer1_outputs(4513)) and (layer1_outputs(6358));
    layer2_outputs(4995) <= not(layer1_outputs(7586));
    layer2_outputs(4996) <= not(layer1_outputs(5118));
    layer2_outputs(4997) <= layer1_outputs(3178);
    layer2_outputs(4998) <= (layer1_outputs(6591)) and (layer1_outputs(5665));
    layer2_outputs(4999) <= not((layer1_outputs(235)) or (layer1_outputs(787)));
    layer2_outputs(5000) <= not(layer1_outputs(478)) or (layer1_outputs(5755));
    layer2_outputs(5001) <= not((layer1_outputs(4763)) and (layer1_outputs(5522)));
    layer2_outputs(5002) <= (layer1_outputs(3300)) and not (layer1_outputs(2357));
    layer2_outputs(5003) <= not((layer1_outputs(869)) and (layer1_outputs(3460)));
    layer2_outputs(5004) <= not(layer1_outputs(3034));
    layer2_outputs(5005) <= not((layer1_outputs(1882)) xor (layer1_outputs(1061)));
    layer2_outputs(5006) <= (layer1_outputs(1660)) xor (layer1_outputs(1896));
    layer2_outputs(5007) <= '0';
    layer2_outputs(5008) <= not(layer1_outputs(7150));
    layer2_outputs(5009) <= layer1_outputs(3504);
    layer2_outputs(5010) <= not(layer1_outputs(2666)) or (layer1_outputs(5470));
    layer2_outputs(5011) <= not((layer1_outputs(2526)) and (layer1_outputs(3709)));
    layer2_outputs(5012) <= not((layer1_outputs(2946)) and (layer1_outputs(5250)));
    layer2_outputs(5013) <= (layer1_outputs(4575)) and (layer1_outputs(1019));
    layer2_outputs(5014) <= (layer1_outputs(6221)) and (layer1_outputs(4252));
    layer2_outputs(5015) <= (layer1_outputs(6430)) and (layer1_outputs(3101));
    layer2_outputs(5016) <= layer1_outputs(4292);
    layer2_outputs(5017) <= not((layer1_outputs(295)) or (layer1_outputs(5623)));
    layer2_outputs(5018) <= not((layer1_outputs(2133)) or (layer1_outputs(6095)));
    layer2_outputs(5019) <= layer1_outputs(3130);
    layer2_outputs(5020) <= (layer1_outputs(2910)) and not (layer1_outputs(4255));
    layer2_outputs(5021) <= layer1_outputs(2036);
    layer2_outputs(5022) <= not((layer1_outputs(7347)) and (layer1_outputs(5845)));
    layer2_outputs(5023) <= not(layer1_outputs(2942));
    layer2_outputs(5024) <= layer1_outputs(3634);
    layer2_outputs(5025) <= (layer1_outputs(5604)) xor (layer1_outputs(6352));
    layer2_outputs(5026) <= (layer1_outputs(4717)) and not (layer1_outputs(6677));
    layer2_outputs(5027) <= not(layer1_outputs(1035)) or (layer1_outputs(5473));
    layer2_outputs(5028) <= not((layer1_outputs(3305)) and (layer1_outputs(6662)));
    layer2_outputs(5029) <= not((layer1_outputs(3662)) and (layer1_outputs(6708)));
    layer2_outputs(5030) <= (layer1_outputs(5336)) and not (layer1_outputs(4012));
    layer2_outputs(5031) <= not(layer1_outputs(1159));
    layer2_outputs(5032) <= not(layer1_outputs(3046));
    layer2_outputs(5033) <= layer1_outputs(578);
    layer2_outputs(5034) <= '1';
    layer2_outputs(5035) <= (layer1_outputs(3488)) or (layer1_outputs(7574));
    layer2_outputs(5036) <= not(layer1_outputs(2049)) or (layer1_outputs(4093));
    layer2_outputs(5037) <= layer1_outputs(4974);
    layer2_outputs(5038) <= not(layer1_outputs(5660));
    layer2_outputs(5039) <= layer1_outputs(5272);
    layer2_outputs(5040) <= not(layer1_outputs(6715)) or (layer1_outputs(5790));
    layer2_outputs(5041) <= (layer1_outputs(6547)) or (layer1_outputs(472));
    layer2_outputs(5042) <= not(layer1_outputs(644)) or (layer1_outputs(6897));
    layer2_outputs(5043) <= not((layer1_outputs(7422)) and (layer1_outputs(4717)));
    layer2_outputs(5044) <= layer1_outputs(1486);
    layer2_outputs(5045) <= layer1_outputs(7432);
    layer2_outputs(5046) <= not((layer1_outputs(2659)) or (layer1_outputs(3395)));
    layer2_outputs(5047) <= layer1_outputs(733);
    layer2_outputs(5048) <= layer1_outputs(1817);
    layer2_outputs(5049) <= (layer1_outputs(302)) and not (layer1_outputs(4197));
    layer2_outputs(5050) <= (layer1_outputs(6379)) and (layer1_outputs(6548));
    layer2_outputs(5051) <= not(layer1_outputs(2931));
    layer2_outputs(5052) <= (layer1_outputs(880)) and not (layer1_outputs(4773));
    layer2_outputs(5053) <= layer1_outputs(5371);
    layer2_outputs(5054) <= (layer1_outputs(3598)) xor (layer1_outputs(6819));
    layer2_outputs(5055) <= not(layer1_outputs(4036));
    layer2_outputs(5056) <= not(layer1_outputs(5170));
    layer2_outputs(5057) <= not((layer1_outputs(6193)) xor (layer1_outputs(5883)));
    layer2_outputs(5058) <= layer1_outputs(7415);
    layer2_outputs(5059) <= (layer1_outputs(2222)) and (layer1_outputs(412));
    layer2_outputs(5060) <= '0';
    layer2_outputs(5061) <= layer1_outputs(7136);
    layer2_outputs(5062) <= not((layer1_outputs(2379)) and (layer1_outputs(5027)));
    layer2_outputs(5063) <= layer1_outputs(1409);
    layer2_outputs(5064) <= not(layer1_outputs(1426));
    layer2_outputs(5065) <= '1';
    layer2_outputs(5066) <= layer1_outputs(5683);
    layer2_outputs(5067) <= not(layer1_outputs(4994));
    layer2_outputs(5068) <= not(layer1_outputs(3409));
    layer2_outputs(5069) <= layer1_outputs(2356);
    layer2_outputs(5070) <= (layer1_outputs(143)) or (layer1_outputs(4728));
    layer2_outputs(5071) <= (layer1_outputs(1639)) or (layer1_outputs(1801));
    layer2_outputs(5072) <= layer1_outputs(3785);
    layer2_outputs(5073) <= layer1_outputs(1221);
    layer2_outputs(5074) <= (layer1_outputs(712)) or (layer1_outputs(2752));
    layer2_outputs(5075) <= '1';
    layer2_outputs(5076) <= layer1_outputs(3616);
    layer2_outputs(5077) <= layer1_outputs(378);
    layer2_outputs(5078) <= layer1_outputs(1877);
    layer2_outputs(5079) <= (layer1_outputs(3421)) and not (layer1_outputs(2983));
    layer2_outputs(5080) <= not(layer1_outputs(1178));
    layer2_outputs(5081) <= not((layer1_outputs(4596)) and (layer1_outputs(2230)));
    layer2_outputs(5082) <= not(layer1_outputs(2687));
    layer2_outputs(5083) <= not(layer1_outputs(6372));
    layer2_outputs(5084) <= (layer1_outputs(4826)) and not (layer1_outputs(5536));
    layer2_outputs(5085) <= '0';
    layer2_outputs(5086) <= layer1_outputs(7460);
    layer2_outputs(5087) <= (layer1_outputs(1493)) xor (layer1_outputs(699));
    layer2_outputs(5088) <= not((layer1_outputs(6537)) and (layer1_outputs(2770)));
    layer2_outputs(5089) <= layer1_outputs(3837);
    layer2_outputs(5090) <= (layer1_outputs(3484)) and not (layer1_outputs(2922));
    layer2_outputs(5091) <= not((layer1_outputs(5854)) and (layer1_outputs(7005)));
    layer2_outputs(5092) <= '1';
    layer2_outputs(5093) <= layer1_outputs(1958);
    layer2_outputs(5094) <= layer1_outputs(941);
    layer2_outputs(5095) <= not(layer1_outputs(630));
    layer2_outputs(5096) <= layer1_outputs(2843);
    layer2_outputs(5097) <= (layer1_outputs(5865)) or (layer1_outputs(140));
    layer2_outputs(5098) <= not(layer1_outputs(5906)) or (layer1_outputs(596));
    layer2_outputs(5099) <= (layer1_outputs(5503)) and not (layer1_outputs(4663));
    layer2_outputs(5100) <= not(layer1_outputs(3070));
    layer2_outputs(5101) <= not(layer1_outputs(1852));
    layer2_outputs(5102) <= not(layer1_outputs(746));
    layer2_outputs(5103) <= not((layer1_outputs(5228)) or (layer1_outputs(6264)));
    layer2_outputs(5104) <= not(layer1_outputs(1924)) or (layer1_outputs(2442));
    layer2_outputs(5105) <= (layer1_outputs(2303)) and not (layer1_outputs(4657));
    layer2_outputs(5106) <= '1';
    layer2_outputs(5107) <= not(layer1_outputs(2128)) or (layer1_outputs(2756));
    layer2_outputs(5108) <= not(layer1_outputs(931));
    layer2_outputs(5109) <= layer1_outputs(2003);
    layer2_outputs(5110) <= not(layer1_outputs(6458)) or (layer1_outputs(3434));
    layer2_outputs(5111) <= (layer1_outputs(3888)) and (layer1_outputs(6047));
    layer2_outputs(5112) <= not((layer1_outputs(2049)) and (layer1_outputs(4784)));
    layer2_outputs(5113) <= (layer1_outputs(7448)) and not (layer1_outputs(198));
    layer2_outputs(5114) <= not(layer1_outputs(1506));
    layer2_outputs(5115) <= layer1_outputs(1357);
    layer2_outputs(5116) <= layer1_outputs(1929);
    layer2_outputs(5117) <= not(layer1_outputs(3696));
    layer2_outputs(5118) <= layer1_outputs(5873);
    layer2_outputs(5119) <= '1';
    layer2_outputs(5120) <= not(layer1_outputs(3890)) or (layer1_outputs(69));
    layer2_outputs(5121) <= layer1_outputs(7077);
    layer2_outputs(5122) <= not((layer1_outputs(2419)) and (layer1_outputs(5877)));
    layer2_outputs(5123) <= not((layer1_outputs(1940)) and (layer1_outputs(5616)));
    layer2_outputs(5124) <= (layer1_outputs(3805)) and not (layer1_outputs(7253));
    layer2_outputs(5125) <= layer1_outputs(4312);
    layer2_outputs(5126) <= (layer1_outputs(114)) or (layer1_outputs(5112));
    layer2_outputs(5127) <= layer1_outputs(3591);
    layer2_outputs(5128) <= layer1_outputs(5513);
    layer2_outputs(5129) <= layer1_outputs(1215);
    layer2_outputs(5130) <= not(layer1_outputs(6108)) or (layer1_outputs(4131));
    layer2_outputs(5131) <= layer1_outputs(6946);
    layer2_outputs(5132) <= '0';
    layer2_outputs(5133) <= layer1_outputs(6469);
    layer2_outputs(5134) <= not(layer1_outputs(2312)) or (layer1_outputs(5804));
    layer2_outputs(5135) <= not(layer1_outputs(2639));
    layer2_outputs(5136) <= not(layer1_outputs(5886));
    layer2_outputs(5137) <= '0';
    layer2_outputs(5138) <= (layer1_outputs(1710)) or (layer1_outputs(1824));
    layer2_outputs(5139) <= layer1_outputs(5897);
    layer2_outputs(5140) <= not(layer1_outputs(2519));
    layer2_outputs(5141) <= (layer1_outputs(2928)) xor (layer1_outputs(5307));
    layer2_outputs(5142) <= not(layer1_outputs(150));
    layer2_outputs(5143) <= (layer1_outputs(5033)) and (layer1_outputs(7334));
    layer2_outputs(5144) <= not(layer1_outputs(5448));
    layer2_outputs(5145) <= not((layer1_outputs(1155)) and (layer1_outputs(1302)));
    layer2_outputs(5146) <= layer1_outputs(6834);
    layer2_outputs(5147) <= not(layer1_outputs(7178));
    layer2_outputs(5148) <= not(layer1_outputs(2376));
    layer2_outputs(5149) <= not(layer1_outputs(7198)) or (layer1_outputs(6419));
    layer2_outputs(5150) <= (layer1_outputs(5137)) and not (layer1_outputs(1952));
    layer2_outputs(5151) <= (layer1_outputs(7366)) and not (layer1_outputs(7168));
    layer2_outputs(5152) <= layer1_outputs(1318);
    layer2_outputs(5153) <= (layer1_outputs(3579)) xor (layer1_outputs(2765));
    layer2_outputs(5154) <= not(layer1_outputs(3181));
    layer2_outputs(5155) <= not(layer1_outputs(4388));
    layer2_outputs(5156) <= not(layer1_outputs(1479));
    layer2_outputs(5157) <= layer1_outputs(3512);
    layer2_outputs(5158) <= not((layer1_outputs(4404)) xor (layer1_outputs(5340)));
    layer2_outputs(5159) <= not(layer1_outputs(2030));
    layer2_outputs(5160) <= (layer1_outputs(4387)) xor (layer1_outputs(1064));
    layer2_outputs(5161) <= layer1_outputs(5317);
    layer2_outputs(5162) <= not(layer1_outputs(1797)) or (layer1_outputs(1619));
    layer2_outputs(5163) <= layer1_outputs(742);
    layer2_outputs(5164) <= layer1_outputs(4272);
    layer2_outputs(5165) <= layer1_outputs(1599);
    layer2_outputs(5166) <= (layer1_outputs(621)) and not (layer1_outputs(1361));
    layer2_outputs(5167) <= (layer1_outputs(5300)) and not (layer1_outputs(2392));
    layer2_outputs(5168) <= not(layer1_outputs(3207)) or (layer1_outputs(6014));
    layer2_outputs(5169) <= layer1_outputs(3891);
    layer2_outputs(5170) <= '1';
    layer2_outputs(5171) <= layer1_outputs(4862);
    layer2_outputs(5172) <= not(layer1_outputs(3348)) or (layer1_outputs(3273));
    layer2_outputs(5173) <= not(layer1_outputs(409)) or (layer1_outputs(2901));
    layer2_outputs(5174) <= (layer1_outputs(2220)) and not (layer1_outputs(1748));
    layer2_outputs(5175) <= layer1_outputs(607);
    layer2_outputs(5176) <= not((layer1_outputs(7609)) and (layer1_outputs(6893)));
    layer2_outputs(5177) <= not(layer1_outputs(6929));
    layer2_outputs(5178) <= (layer1_outputs(99)) and (layer1_outputs(1341));
    layer2_outputs(5179) <= (layer1_outputs(4189)) and not (layer1_outputs(2540));
    layer2_outputs(5180) <= not(layer1_outputs(3702));
    layer2_outputs(5181) <= (layer1_outputs(4397)) or (layer1_outputs(5538));
    layer2_outputs(5182) <= not(layer1_outputs(6289)) or (layer1_outputs(4930));
    layer2_outputs(5183) <= (layer1_outputs(7629)) xor (layer1_outputs(5329));
    layer2_outputs(5184) <= not(layer1_outputs(4152)) or (layer1_outputs(662));
    layer2_outputs(5185) <= not(layer1_outputs(7083));
    layer2_outputs(5186) <= not(layer1_outputs(7655));
    layer2_outputs(5187) <= not(layer1_outputs(6969));
    layer2_outputs(5188) <= not(layer1_outputs(2608));
    layer2_outputs(5189) <= not(layer1_outputs(4660));
    layer2_outputs(5190) <= not(layer1_outputs(2883));
    layer2_outputs(5191) <= (layer1_outputs(6042)) and (layer1_outputs(3178));
    layer2_outputs(5192) <= (layer1_outputs(2722)) xor (layer1_outputs(6208));
    layer2_outputs(5193) <= not(layer1_outputs(6833));
    layer2_outputs(5194) <= not(layer1_outputs(5044)) or (layer1_outputs(5022));
    layer2_outputs(5195) <= (layer1_outputs(392)) and (layer1_outputs(6307));
    layer2_outputs(5196) <= (layer1_outputs(4295)) and (layer1_outputs(7203));
    layer2_outputs(5197) <= not((layer1_outputs(148)) xor (layer1_outputs(5205)));
    layer2_outputs(5198) <= not(layer1_outputs(5375)) or (layer1_outputs(7668));
    layer2_outputs(5199) <= not(layer1_outputs(3357)) or (layer1_outputs(1666));
    layer2_outputs(5200) <= (layer1_outputs(3073)) and not (layer1_outputs(6119));
    layer2_outputs(5201) <= not(layer1_outputs(1784)) or (layer1_outputs(7434));
    layer2_outputs(5202) <= not(layer1_outputs(7462));
    layer2_outputs(5203) <= not(layer1_outputs(5842));
    layer2_outputs(5204) <= layer1_outputs(5638);
    layer2_outputs(5205) <= '0';
    layer2_outputs(5206) <= not(layer1_outputs(1955));
    layer2_outputs(5207) <= not(layer1_outputs(2232));
    layer2_outputs(5208) <= not((layer1_outputs(3995)) and (layer1_outputs(2812)));
    layer2_outputs(5209) <= (layer1_outputs(3504)) xor (layer1_outputs(7093));
    layer2_outputs(5210) <= not(layer1_outputs(4609));
    layer2_outputs(5211) <= not((layer1_outputs(1649)) or (layer1_outputs(6043)));
    layer2_outputs(5212) <= not(layer1_outputs(2288)) or (layer1_outputs(6050));
    layer2_outputs(5213) <= layer1_outputs(1250);
    layer2_outputs(5214) <= (layer1_outputs(942)) xor (layer1_outputs(5365));
    layer2_outputs(5215) <= not(layer1_outputs(4593)) or (layer1_outputs(6493));
    layer2_outputs(5216) <= not((layer1_outputs(1011)) or (layer1_outputs(1451)));
    layer2_outputs(5217) <= not((layer1_outputs(7394)) and (layer1_outputs(2050)));
    layer2_outputs(5218) <= layer1_outputs(7270);
    layer2_outputs(5219) <= not(layer1_outputs(1425)) or (layer1_outputs(1842));
    layer2_outputs(5220) <= not(layer1_outputs(254));
    layer2_outputs(5221) <= (layer1_outputs(3133)) and not (layer1_outputs(1721));
    layer2_outputs(5222) <= not(layer1_outputs(1555));
    layer2_outputs(5223) <= layer1_outputs(5385);
    layer2_outputs(5224) <= '1';
    layer2_outputs(5225) <= (layer1_outputs(6541)) and not (layer1_outputs(77));
    layer2_outputs(5226) <= layer1_outputs(5006);
    layer2_outputs(5227) <= not(layer1_outputs(1977));
    layer2_outputs(5228) <= '1';
    layer2_outputs(5229) <= (layer1_outputs(5794)) and (layer1_outputs(5732));
    layer2_outputs(5230) <= (layer1_outputs(5630)) or (layer1_outputs(751));
    layer2_outputs(5231) <= layer1_outputs(301);
    layer2_outputs(5232) <= layer1_outputs(4226);
    layer2_outputs(5233) <= '0';
    layer2_outputs(5234) <= (layer1_outputs(3507)) and not (layer1_outputs(3360));
    layer2_outputs(5235) <= not((layer1_outputs(3048)) or (layer1_outputs(6763)));
    layer2_outputs(5236) <= not((layer1_outputs(5898)) or (layer1_outputs(7523)));
    layer2_outputs(5237) <= not(layer1_outputs(966)) or (layer1_outputs(2210));
    layer2_outputs(5238) <= not(layer1_outputs(1485));
    layer2_outputs(5239) <= (layer1_outputs(3464)) and not (layer1_outputs(2213));
    layer2_outputs(5240) <= not(layer1_outputs(2448));
    layer2_outputs(5241) <= not((layer1_outputs(5462)) or (layer1_outputs(3424)));
    layer2_outputs(5242) <= (layer1_outputs(4461)) and not (layer1_outputs(1774));
    layer2_outputs(5243) <= not(layer1_outputs(2591));
    layer2_outputs(5244) <= '1';
    layer2_outputs(5245) <= not(layer1_outputs(1030)) or (layer1_outputs(3618));
    layer2_outputs(5246) <= not(layer1_outputs(4830)) or (layer1_outputs(4377));
    layer2_outputs(5247) <= not(layer1_outputs(1976));
    layer2_outputs(5248) <= layer1_outputs(4604);
    layer2_outputs(5249) <= not(layer1_outputs(6730)) or (layer1_outputs(4501));
    layer2_outputs(5250) <= (layer1_outputs(5651)) xor (layer1_outputs(5411));
    layer2_outputs(5251) <= (layer1_outputs(4098)) and (layer1_outputs(1323));
    layer2_outputs(5252) <= not((layer1_outputs(5050)) xor (layer1_outputs(831)));
    layer2_outputs(5253) <= layer1_outputs(3011);
    layer2_outputs(5254) <= not(layer1_outputs(5409));
    layer2_outputs(5255) <= not(layer1_outputs(1168)) or (layer1_outputs(7371));
    layer2_outputs(5256) <= '0';
    layer2_outputs(5257) <= not(layer1_outputs(3752));
    layer2_outputs(5258) <= (layer1_outputs(3816)) and (layer1_outputs(1241));
    layer2_outputs(5259) <= layer1_outputs(2963);
    layer2_outputs(5260) <= layer1_outputs(2800);
    layer2_outputs(5261) <= layer1_outputs(5180);
    layer2_outputs(5262) <= (layer1_outputs(6279)) and not (layer1_outputs(652));
    layer2_outputs(5263) <= layer1_outputs(7638);
    layer2_outputs(5264) <= layer1_outputs(4573);
    layer2_outputs(5265) <= not(layer1_outputs(4754)) or (layer1_outputs(3648));
    layer2_outputs(5266) <= not(layer1_outputs(7158)) or (layer1_outputs(4941));
    layer2_outputs(5267) <= (layer1_outputs(1160)) and (layer1_outputs(7426));
    layer2_outputs(5268) <= not((layer1_outputs(4936)) or (layer1_outputs(3688)));
    layer2_outputs(5269) <= not(layer1_outputs(1418));
    layer2_outputs(5270) <= layer1_outputs(3047);
    layer2_outputs(5271) <= not(layer1_outputs(3708)) or (layer1_outputs(2184));
    layer2_outputs(5272) <= not((layer1_outputs(7423)) or (layer1_outputs(4542)));
    layer2_outputs(5273) <= not(layer1_outputs(3776));
    layer2_outputs(5274) <= (layer1_outputs(6612)) and (layer1_outputs(3560));
    layer2_outputs(5275) <= not(layer1_outputs(6420));
    layer2_outputs(5276) <= not(layer1_outputs(4705));
    layer2_outputs(5277) <= (layer1_outputs(4253)) and not (layer1_outputs(6459));
    layer2_outputs(5278) <= (layer1_outputs(2609)) xor (layer1_outputs(7419));
    layer2_outputs(5279) <= (layer1_outputs(563)) and not (layer1_outputs(2857));
    layer2_outputs(5280) <= not((layer1_outputs(5957)) or (layer1_outputs(4201)));
    layer2_outputs(5281) <= layer1_outputs(5846);
    layer2_outputs(5282) <= (layer1_outputs(3651)) and not (layer1_outputs(4134));
    layer2_outputs(5283) <= not(layer1_outputs(887));
    layer2_outputs(5284) <= layer1_outputs(1360);
    layer2_outputs(5285) <= layer1_outputs(6519);
    layer2_outputs(5286) <= (layer1_outputs(5893)) or (layer1_outputs(2734));
    layer2_outputs(5287) <= (layer1_outputs(961)) and (layer1_outputs(4842));
    layer2_outputs(5288) <= not(layer1_outputs(2403));
    layer2_outputs(5289) <= layer1_outputs(1785);
    layer2_outputs(5290) <= not(layer1_outputs(2809));
    layer2_outputs(5291) <= not((layer1_outputs(2108)) and (layer1_outputs(3493)));
    layer2_outputs(5292) <= not(layer1_outputs(5399));
    layer2_outputs(5293) <= not(layer1_outputs(1453));
    layer2_outputs(5294) <= (layer1_outputs(2152)) and not (layer1_outputs(436));
    layer2_outputs(5295) <= (layer1_outputs(1109)) and not (layer1_outputs(49));
    layer2_outputs(5296) <= (layer1_outputs(5407)) and (layer1_outputs(4884));
    layer2_outputs(5297) <= layer1_outputs(5150);
    layer2_outputs(5298) <= not(layer1_outputs(7290));
    layer2_outputs(5299) <= (layer1_outputs(5591)) or (layer1_outputs(6332));
    layer2_outputs(5300) <= layer1_outputs(3904);
    layer2_outputs(5301) <= not(layer1_outputs(1206));
    layer2_outputs(5302) <= not((layer1_outputs(4631)) or (layer1_outputs(4490)));
    layer2_outputs(5303) <= not((layer1_outputs(4322)) or (layer1_outputs(6045)));
    layer2_outputs(5304) <= not((layer1_outputs(5437)) xor (layer1_outputs(190)));
    layer2_outputs(5305) <= not(layer1_outputs(5521)) or (layer1_outputs(5525));
    layer2_outputs(5306) <= layer1_outputs(4690);
    layer2_outputs(5307) <= (layer1_outputs(1661)) and not (layer1_outputs(4529));
    layer2_outputs(5308) <= (layer1_outputs(1622)) and not (layer1_outputs(6181));
    layer2_outputs(5309) <= layer1_outputs(4197);
    layer2_outputs(5310) <= layer1_outputs(5360);
    layer2_outputs(5311) <= not(layer1_outputs(5285));
    layer2_outputs(5312) <= not(layer1_outputs(3466));
    layer2_outputs(5313) <= not((layer1_outputs(3452)) or (layer1_outputs(4045)));
    layer2_outputs(5314) <= not(layer1_outputs(5984));
    layer2_outputs(5315) <= '0';
    layer2_outputs(5316) <= not(layer1_outputs(1391));
    layer2_outputs(5317) <= layer1_outputs(374);
    layer2_outputs(5318) <= layer1_outputs(1898);
    layer2_outputs(5319) <= layer1_outputs(3245);
    layer2_outputs(5320) <= not(layer1_outputs(4732)) or (layer1_outputs(1669));
    layer2_outputs(5321) <= not(layer1_outputs(1166));
    layer2_outputs(5322) <= not(layer1_outputs(4567)) or (layer1_outputs(4653));
    layer2_outputs(5323) <= not(layer1_outputs(7487));
    layer2_outputs(5324) <= (layer1_outputs(2203)) and (layer1_outputs(7473));
    layer2_outputs(5325) <= not((layer1_outputs(3880)) or (layer1_outputs(7316)));
    layer2_outputs(5326) <= layer1_outputs(1468);
    layer2_outputs(5327) <= (layer1_outputs(4421)) and (layer1_outputs(2920));
    layer2_outputs(5328) <= not((layer1_outputs(3052)) or (layer1_outputs(1719)));
    layer2_outputs(5329) <= not(layer1_outputs(1613)) or (layer1_outputs(5063));
    layer2_outputs(5330) <= not(layer1_outputs(1394)) or (layer1_outputs(125));
    layer2_outputs(5331) <= (layer1_outputs(6438)) or (layer1_outputs(3043));
    layer2_outputs(5332) <= (layer1_outputs(2713)) and (layer1_outputs(3897));
    layer2_outputs(5333) <= '1';
    layer2_outputs(5334) <= not(layer1_outputs(3016));
    layer2_outputs(5335) <= '1';
    layer2_outputs(5336) <= not((layer1_outputs(2645)) or (layer1_outputs(4729)));
    layer2_outputs(5337) <= not(layer1_outputs(2463)) or (layer1_outputs(6457));
    layer2_outputs(5338) <= not(layer1_outputs(670));
    layer2_outputs(5339) <= not((layer1_outputs(3060)) or (layer1_outputs(5308)));
    layer2_outputs(5340) <= layer1_outputs(7604);
    layer2_outputs(5341) <= '1';
    layer2_outputs(5342) <= (layer1_outputs(6712)) and not (layer1_outputs(7342));
    layer2_outputs(5343) <= not(layer1_outputs(1378));
    layer2_outputs(5344) <= layer1_outputs(4367);
    layer2_outputs(5345) <= not((layer1_outputs(4290)) xor (layer1_outputs(2761)));
    layer2_outputs(5346) <= (layer1_outputs(3631)) and (layer1_outputs(1324));
    layer2_outputs(5347) <= not((layer1_outputs(181)) or (layer1_outputs(3654)));
    layer2_outputs(5348) <= not((layer1_outputs(7519)) and (layer1_outputs(6500)));
    layer2_outputs(5349) <= not((layer1_outputs(961)) and (layer1_outputs(6807)));
    layer2_outputs(5350) <= (layer1_outputs(5120)) or (layer1_outputs(1044));
    layer2_outputs(5351) <= not(layer1_outputs(6641));
    layer2_outputs(5352) <= not(layer1_outputs(5119));
    layer2_outputs(5353) <= not(layer1_outputs(7612));
    layer2_outputs(5354) <= (layer1_outputs(5082)) or (layer1_outputs(184));
    layer2_outputs(5355) <= not(layer1_outputs(4812));
    layer2_outputs(5356) <= layer1_outputs(529);
    layer2_outputs(5357) <= not((layer1_outputs(3228)) or (layer1_outputs(6020)));
    layer2_outputs(5358) <= layer1_outputs(4843);
    layer2_outputs(5359) <= '0';
    layer2_outputs(5360) <= not((layer1_outputs(3014)) and (layer1_outputs(4383)));
    layer2_outputs(5361) <= not(layer1_outputs(2618));
    layer2_outputs(5362) <= not((layer1_outputs(916)) and (layer1_outputs(2149)));
    layer2_outputs(5363) <= (layer1_outputs(2037)) and (layer1_outputs(3482));
    layer2_outputs(5364) <= layer1_outputs(3512);
    layer2_outputs(5365) <= not((layer1_outputs(6522)) xor (layer1_outputs(6597)));
    layer2_outputs(5366) <= (layer1_outputs(1374)) and not (layer1_outputs(1807));
    layer2_outputs(5367) <= layer1_outputs(3277);
    layer2_outputs(5368) <= (layer1_outputs(1985)) and not (layer1_outputs(633));
    layer2_outputs(5369) <= '1';
    layer2_outputs(5370) <= (layer1_outputs(5354)) xor (layer1_outputs(253));
    layer2_outputs(5371) <= not(layer1_outputs(3190));
    layer2_outputs(5372) <= not(layer1_outputs(2425)) or (layer1_outputs(2563));
    layer2_outputs(5373) <= (layer1_outputs(5666)) and not (layer1_outputs(1655));
    layer2_outputs(5374) <= (layer1_outputs(6936)) and not (layer1_outputs(6194));
    layer2_outputs(5375) <= not((layer1_outputs(3054)) or (layer1_outputs(2123)));
    layer2_outputs(5376) <= not(layer1_outputs(78));
    layer2_outputs(5377) <= '1';
    layer2_outputs(5378) <= '1';
    layer2_outputs(5379) <= '1';
    layer2_outputs(5380) <= layer1_outputs(865);
    layer2_outputs(5381) <= layer1_outputs(1893);
    layer2_outputs(5382) <= (layer1_outputs(2987)) and not (layer1_outputs(7557));
    layer2_outputs(5383) <= not(layer1_outputs(7033)) or (layer1_outputs(4102));
    layer2_outputs(5384) <= (layer1_outputs(7516)) or (layer1_outputs(7456));
    layer2_outputs(5385) <= not((layer1_outputs(5697)) and (layer1_outputs(319)));
    layer2_outputs(5386) <= (layer1_outputs(1725)) or (layer1_outputs(5108));
    layer2_outputs(5387) <= not((layer1_outputs(1024)) and (layer1_outputs(7331)));
    layer2_outputs(5388) <= not((layer1_outputs(2965)) or (layer1_outputs(7679)));
    layer2_outputs(5389) <= not((layer1_outputs(5731)) and (layer1_outputs(1191)));
    layer2_outputs(5390) <= not(layer1_outputs(5513));
    layer2_outputs(5391) <= layer1_outputs(5593);
    layer2_outputs(5392) <= not(layer1_outputs(300));
    layer2_outputs(5393) <= '1';
    layer2_outputs(5394) <= not(layer1_outputs(2794));
    layer2_outputs(5395) <= not(layer1_outputs(564)) or (layer1_outputs(1806));
    layer2_outputs(5396) <= not((layer1_outputs(117)) or (layer1_outputs(4489)));
    layer2_outputs(5397) <= (layer1_outputs(4453)) and not (layer1_outputs(3206));
    layer2_outputs(5398) <= not(layer1_outputs(5736));
    layer2_outputs(5399) <= not(layer1_outputs(3996));
    layer2_outputs(5400) <= not((layer1_outputs(5801)) or (layer1_outputs(6128)));
    layer2_outputs(5401) <= (layer1_outputs(7498)) and not (layer1_outputs(426));
    layer2_outputs(5402) <= not(layer1_outputs(2142)) or (layer1_outputs(6548));
    layer2_outputs(5403) <= layer1_outputs(259);
    layer2_outputs(5404) <= (layer1_outputs(6610)) and not (layer1_outputs(2191));
    layer2_outputs(5405) <= (layer1_outputs(478)) and not (layer1_outputs(2589));
    layer2_outputs(5406) <= (layer1_outputs(7275)) and (layer1_outputs(968));
    layer2_outputs(5407) <= not(layer1_outputs(3704));
    layer2_outputs(5408) <= not(layer1_outputs(3332)) or (layer1_outputs(6407));
    layer2_outputs(5409) <= (layer1_outputs(4774)) and not (layer1_outputs(5240));
    layer2_outputs(5410) <= layer1_outputs(2981);
    layer2_outputs(5411) <= not(layer1_outputs(4768));
    layer2_outputs(5412) <= layer1_outputs(1692);
    layer2_outputs(5413) <= not(layer1_outputs(1295));
    layer2_outputs(5414) <= not(layer1_outputs(4675));
    layer2_outputs(5415) <= (layer1_outputs(4104)) and not (layer1_outputs(454));
    layer2_outputs(5416) <= layer1_outputs(1559);
    layer2_outputs(5417) <= '0';
    layer2_outputs(5418) <= not(layer1_outputs(660));
    layer2_outputs(5419) <= layer1_outputs(5570);
    layer2_outputs(5420) <= (layer1_outputs(7458)) and not (layer1_outputs(2395));
    layer2_outputs(5421) <= (layer1_outputs(6000)) and not (layer1_outputs(6878));
    layer2_outputs(5422) <= '1';
    layer2_outputs(5423) <= (layer1_outputs(3308)) or (layer1_outputs(4747));
    layer2_outputs(5424) <= not(layer1_outputs(2402)) or (layer1_outputs(2711));
    layer2_outputs(5425) <= layer1_outputs(6129);
    layer2_outputs(5426) <= (layer1_outputs(3960)) and not (layer1_outputs(4604));
    layer2_outputs(5427) <= not(layer1_outputs(2520));
    layer2_outputs(5428) <= not(layer1_outputs(128));
    layer2_outputs(5429) <= (layer1_outputs(6542)) and not (layer1_outputs(4470));
    layer2_outputs(5430) <= not(layer1_outputs(874)) or (layer1_outputs(3726));
    layer2_outputs(5431) <= layer1_outputs(2965);
    layer2_outputs(5432) <= (layer1_outputs(598)) and not (layer1_outputs(557));
    layer2_outputs(5433) <= not((layer1_outputs(1987)) and (layer1_outputs(2489)));
    layer2_outputs(5434) <= not((layer1_outputs(5612)) and (layer1_outputs(1161)));
    layer2_outputs(5435) <= (layer1_outputs(3948)) and not (layer1_outputs(1141));
    layer2_outputs(5436) <= not((layer1_outputs(470)) and (layer1_outputs(5100)));
    layer2_outputs(5437) <= (layer1_outputs(3679)) and not (layer1_outputs(4329));
    layer2_outputs(5438) <= (layer1_outputs(5928)) and not (layer1_outputs(7171));
    layer2_outputs(5439) <= layer1_outputs(3304);
    layer2_outputs(5440) <= not(layer1_outputs(6524));
    layer2_outputs(5441) <= not(layer1_outputs(5772)) or (layer1_outputs(6272));
    layer2_outputs(5442) <= (layer1_outputs(5611)) or (layer1_outputs(4954));
    layer2_outputs(5443) <= (layer1_outputs(6931)) and (layer1_outputs(1336));
    layer2_outputs(5444) <= not(layer1_outputs(2408));
    layer2_outputs(5445) <= '0';
    layer2_outputs(5446) <= (layer1_outputs(1816)) and not (layer1_outputs(1557));
    layer2_outputs(5447) <= not(layer1_outputs(1728));
    layer2_outputs(5448) <= not((layer1_outputs(6283)) and (layer1_outputs(1566)));
    layer2_outputs(5449) <= not(layer1_outputs(1139));
    layer2_outputs(5450) <= (layer1_outputs(3039)) or (layer1_outputs(2933));
    layer2_outputs(5451) <= layer1_outputs(255);
    layer2_outputs(5452) <= layer1_outputs(5196);
    layer2_outputs(5453) <= not(layer1_outputs(5501)) or (layer1_outputs(4416));
    layer2_outputs(5454) <= (layer1_outputs(4300)) xor (layer1_outputs(1618));
    layer2_outputs(5455) <= not((layer1_outputs(7116)) and (layer1_outputs(5934)));
    layer2_outputs(5456) <= layer1_outputs(3253);
    layer2_outputs(5457) <= (layer1_outputs(7529)) and not (layer1_outputs(6271));
    layer2_outputs(5458) <= '0';
    layer2_outputs(5459) <= layer1_outputs(6308);
    layer2_outputs(5460) <= layer1_outputs(7321);
    layer2_outputs(5461) <= not((layer1_outputs(2446)) and (layer1_outputs(4474)));
    layer2_outputs(5462) <= '0';
    layer2_outputs(5463) <= not(layer1_outputs(2898)) or (layer1_outputs(4663));
    layer2_outputs(5464) <= not((layer1_outputs(318)) or (layer1_outputs(2033)));
    layer2_outputs(5465) <= layer1_outputs(4617);
    layer2_outputs(5466) <= not(layer1_outputs(2056));
    layer2_outputs(5467) <= (layer1_outputs(7422)) xor (layer1_outputs(1988));
    layer2_outputs(5468) <= not(layer1_outputs(3629));
    layer2_outputs(5469) <= not(layer1_outputs(3089)) or (layer1_outputs(2855));
    layer2_outputs(5470) <= '0';
    layer2_outputs(5471) <= not((layer1_outputs(5765)) or (layer1_outputs(4257)));
    layer2_outputs(5472) <= (layer1_outputs(107)) or (layer1_outputs(5263));
    layer2_outputs(5473) <= not(layer1_outputs(7233));
    layer2_outputs(5474) <= (layer1_outputs(4824)) and (layer1_outputs(2558));
    layer2_outputs(5475) <= (layer1_outputs(2820)) and not (layer1_outputs(6436));
    layer2_outputs(5476) <= not(layer1_outputs(6562));
    layer2_outputs(5477) <= '0';
    layer2_outputs(5478) <= layer1_outputs(4028);
    layer2_outputs(5479) <= not(layer1_outputs(5567)) or (layer1_outputs(4185));
    layer2_outputs(5480) <= not(layer1_outputs(2725));
    layer2_outputs(5481) <= not(layer1_outputs(3786));
    layer2_outputs(5482) <= not((layer1_outputs(1261)) or (layer1_outputs(3112)));
    layer2_outputs(5483) <= '0';
    layer2_outputs(5484) <= (layer1_outputs(5832)) and (layer1_outputs(6423));
    layer2_outputs(5485) <= not((layer1_outputs(7129)) or (layer1_outputs(4614)));
    layer2_outputs(5486) <= layer1_outputs(1438);
    layer2_outputs(5487) <= not(layer1_outputs(7245)) or (layer1_outputs(1604));
    layer2_outputs(5488) <= not(layer1_outputs(4163));
    layer2_outputs(5489) <= (layer1_outputs(4205)) or (layer1_outputs(3755));
    layer2_outputs(5490) <= layer1_outputs(4889);
    layer2_outputs(5491) <= '1';
    layer2_outputs(5492) <= layer1_outputs(62);
    layer2_outputs(5493) <= not(layer1_outputs(2445));
    layer2_outputs(5494) <= not(layer1_outputs(7026));
    layer2_outputs(5495) <= (layer1_outputs(3617)) and not (layer1_outputs(721));
    layer2_outputs(5496) <= (layer1_outputs(3543)) and not (layer1_outputs(4149));
    layer2_outputs(5497) <= not((layer1_outputs(4370)) or (layer1_outputs(2313)));
    layer2_outputs(5498) <= layer1_outputs(505);
    layer2_outputs(5499) <= (layer1_outputs(4221)) or (layer1_outputs(2837));
    layer2_outputs(5500) <= (layer1_outputs(2595)) and (layer1_outputs(4926));
    layer2_outputs(5501) <= (layer1_outputs(7327)) and not (layer1_outputs(2267));
    layer2_outputs(5502) <= (layer1_outputs(6658)) and (layer1_outputs(5562));
    layer2_outputs(5503) <= not((layer1_outputs(7209)) and (layer1_outputs(369)));
    layer2_outputs(5504) <= not(layer1_outputs(5273));
    layer2_outputs(5505) <= (layer1_outputs(30)) and not (layer1_outputs(4954));
    layer2_outputs(5506) <= (layer1_outputs(3019)) and not (layer1_outputs(5589));
    layer2_outputs(5507) <= not(layer1_outputs(3980));
    layer2_outputs(5508) <= '1';
    layer2_outputs(5509) <= (layer1_outputs(4927)) and (layer1_outputs(173));
    layer2_outputs(5510) <= (layer1_outputs(2195)) and not (layer1_outputs(6973));
    layer2_outputs(5511) <= not((layer1_outputs(2006)) and (layer1_outputs(5967)));
    layer2_outputs(5512) <= (layer1_outputs(701)) xor (layer1_outputs(2233));
    layer2_outputs(5513) <= not(layer1_outputs(4038));
    layer2_outputs(5514) <= layer1_outputs(4592);
    layer2_outputs(5515) <= (layer1_outputs(1439)) and (layer1_outputs(6349));
    layer2_outputs(5516) <= not(layer1_outputs(5475)) or (layer1_outputs(373));
    layer2_outputs(5517) <= (layer1_outputs(115)) and not (layer1_outputs(6449));
    layer2_outputs(5518) <= not(layer1_outputs(3211));
    layer2_outputs(5519) <= not(layer1_outputs(1491));
    layer2_outputs(5520) <= not(layer1_outputs(386)) or (layer1_outputs(5932));
    layer2_outputs(5521) <= not(layer1_outputs(7225));
    layer2_outputs(5522) <= not((layer1_outputs(4903)) xor (layer1_outputs(5708)));
    layer2_outputs(5523) <= not((layer1_outputs(3931)) and (layer1_outputs(6756)));
    layer2_outputs(5524) <= (layer1_outputs(6321)) and (layer1_outputs(6394));
    layer2_outputs(5525) <= not(layer1_outputs(4344)) or (layer1_outputs(5450));
    layer2_outputs(5526) <= '0';
    layer2_outputs(5527) <= '0';
    layer2_outputs(5528) <= layer1_outputs(5533);
    layer2_outputs(5529) <= not(layer1_outputs(4533));
    layer2_outputs(5530) <= (layer1_outputs(7358)) and not (layer1_outputs(6362));
    layer2_outputs(5531) <= layer1_outputs(5064);
    layer2_outputs(5532) <= not((layer1_outputs(4803)) and (layer1_outputs(5317)));
    layer2_outputs(5533) <= '1';
    layer2_outputs(5534) <= not((layer1_outputs(1585)) or (layer1_outputs(3748)));
    layer2_outputs(5535) <= not(layer1_outputs(496));
    layer2_outputs(5536) <= not(layer1_outputs(3171));
    layer2_outputs(5537) <= (layer1_outputs(3929)) and (layer1_outputs(6942));
    layer2_outputs(5538) <= (layer1_outputs(5)) and (layer1_outputs(4091));
    layer2_outputs(5539) <= (layer1_outputs(2954)) and not (layer1_outputs(3820));
    layer2_outputs(5540) <= not((layer1_outputs(3469)) or (layer1_outputs(3924)));
    layer2_outputs(5541) <= not(layer1_outputs(3050));
    layer2_outputs(5542) <= not(layer1_outputs(4368));
    layer2_outputs(5543) <= (layer1_outputs(3416)) and not (layer1_outputs(654));
    layer2_outputs(5544) <= not(layer1_outputs(6713));
    layer2_outputs(5545) <= layer1_outputs(1347);
    layer2_outputs(5546) <= (layer1_outputs(6541)) or (layer1_outputs(3525));
    layer2_outputs(5547) <= '1';
    layer2_outputs(5548) <= layer1_outputs(2148);
    layer2_outputs(5549) <= (layer1_outputs(4365)) and not (layer1_outputs(5003));
    layer2_outputs(5550) <= layer1_outputs(7372);
    layer2_outputs(5551) <= not(layer1_outputs(5918)) or (layer1_outputs(3831));
    layer2_outputs(5552) <= layer1_outputs(859);
    layer2_outputs(5553) <= not(layer1_outputs(382)) or (layer1_outputs(1009));
    layer2_outputs(5554) <= (layer1_outputs(5704)) xor (layer1_outputs(866));
    layer2_outputs(5555) <= not(layer1_outputs(173));
    layer2_outputs(5556) <= (layer1_outputs(138)) and not (layer1_outputs(3902));
    layer2_outputs(5557) <= '1';
    layer2_outputs(5558) <= layer1_outputs(5436);
    layer2_outputs(5559) <= layer1_outputs(6865);
    layer2_outputs(5560) <= not(layer1_outputs(2231));
    layer2_outputs(5561) <= (layer1_outputs(479)) and not (layer1_outputs(542));
    layer2_outputs(5562) <= layer1_outputs(4975);
    layer2_outputs(5563) <= (layer1_outputs(7002)) or (layer1_outputs(6113));
    layer2_outputs(5564) <= layer1_outputs(2667);
    layer2_outputs(5565) <= not((layer1_outputs(7574)) or (layer1_outputs(6507)));
    layer2_outputs(5566) <= not(layer1_outputs(2556));
    layer2_outputs(5567) <= layer1_outputs(6353);
    layer2_outputs(5568) <= not((layer1_outputs(1569)) and (layer1_outputs(3078)));
    layer2_outputs(5569) <= not(layer1_outputs(1862));
    layer2_outputs(5570) <= layer1_outputs(3038);
    layer2_outputs(5571) <= not(layer1_outputs(1502)) or (layer1_outputs(3027));
    layer2_outputs(5572) <= not(layer1_outputs(3902));
    layer2_outputs(5573) <= not(layer1_outputs(7025)) or (layer1_outputs(2684));
    layer2_outputs(5574) <= (layer1_outputs(4062)) and not (layer1_outputs(1606));
    layer2_outputs(5575) <= (layer1_outputs(5611)) xor (layer1_outputs(6170));
    layer2_outputs(5576) <= not(layer1_outputs(3182)) or (layer1_outputs(6515));
    layer2_outputs(5577) <= not(layer1_outputs(3871));
    layer2_outputs(5578) <= '1';
    layer2_outputs(5579) <= not(layer1_outputs(3613));
    layer2_outputs(5580) <= not(layer1_outputs(6790));
    layer2_outputs(5581) <= not(layer1_outputs(4818)) or (layer1_outputs(5092));
    layer2_outputs(5582) <= not(layer1_outputs(3760));
    layer2_outputs(5583) <= layer1_outputs(3986);
    layer2_outputs(5584) <= (layer1_outputs(9)) and not (layer1_outputs(2692));
    layer2_outputs(5585) <= not(layer1_outputs(4895));
    layer2_outputs(5586) <= not(layer1_outputs(1993));
    layer2_outputs(5587) <= not((layer1_outputs(1525)) and (layer1_outputs(397)));
    layer2_outputs(5588) <= '1';
    layer2_outputs(5589) <= (layer1_outputs(7348)) or (layer1_outputs(4010));
    layer2_outputs(5590) <= (layer1_outputs(894)) and not (layer1_outputs(7548));
    layer2_outputs(5591) <= not(layer1_outputs(2622));
    layer2_outputs(5592) <= not(layer1_outputs(5633)) or (layer1_outputs(5874));
    layer2_outputs(5593) <= (layer1_outputs(5284)) or (layer1_outputs(1566));
    layer2_outputs(5594) <= layer1_outputs(583);
    layer2_outputs(5595) <= not(layer1_outputs(7249)) or (layer1_outputs(6124));
    layer2_outputs(5596) <= not(layer1_outputs(5103));
    layer2_outputs(5597) <= (layer1_outputs(1284)) and (layer1_outputs(2566));
    layer2_outputs(5598) <= (layer1_outputs(6777)) and (layer1_outputs(1584));
    layer2_outputs(5599) <= not(layer1_outputs(1049)) or (layer1_outputs(2095));
    layer2_outputs(5600) <= '0';
    layer2_outputs(5601) <= not(layer1_outputs(6672));
    layer2_outputs(5602) <= (layer1_outputs(4326)) or (layer1_outputs(6513));
    layer2_outputs(5603) <= layer1_outputs(151);
    layer2_outputs(5604) <= layer1_outputs(1603);
    layer2_outputs(5605) <= not(layer1_outputs(1855));
    layer2_outputs(5606) <= layer1_outputs(152);
    layer2_outputs(5607) <= layer1_outputs(6246);
    layer2_outputs(5608) <= not(layer1_outputs(1228)) or (layer1_outputs(2100));
    layer2_outputs(5609) <= '0';
    layer2_outputs(5610) <= not(layer1_outputs(6116));
    layer2_outputs(5611) <= not((layer1_outputs(3152)) or (layer1_outputs(6494)));
    layer2_outputs(5612) <= not(layer1_outputs(4180));
    layer2_outputs(5613) <= not(layer1_outputs(3101));
    layer2_outputs(5614) <= not(layer1_outputs(5950));
    layer2_outputs(5615) <= not(layer1_outputs(2221)) or (layer1_outputs(6847));
    layer2_outputs(5616) <= '1';
    layer2_outputs(5617) <= not((layer1_outputs(3221)) or (layer1_outputs(5386)));
    layer2_outputs(5618) <= not((layer1_outputs(544)) and (layer1_outputs(412)));
    layer2_outputs(5619) <= not((layer1_outputs(6705)) or (layer1_outputs(908)));
    layer2_outputs(5620) <= not(layer1_outputs(136));
    layer2_outputs(5621) <= not(layer1_outputs(6462));
    layer2_outputs(5622) <= not((layer1_outputs(360)) or (layer1_outputs(5738)));
    layer2_outputs(5623) <= not(layer1_outputs(5337));
    layer2_outputs(5624) <= (layer1_outputs(155)) and (layer1_outputs(5012));
    layer2_outputs(5625) <= layer1_outputs(4161);
    layer2_outputs(5626) <= not(layer1_outputs(649));
    layer2_outputs(5627) <= not((layer1_outputs(7477)) and (layer1_outputs(4735)));
    layer2_outputs(5628) <= not(layer1_outputs(3847));
    layer2_outputs(5629) <= not((layer1_outputs(348)) or (layer1_outputs(1508)));
    layer2_outputs(5630) <= (layer1_outputs(6039)) and (layer1_outputs(2719));
    layer2_outputs(5631) <= layer1_outputs(3368);
    layer2_outputs(5632) <= not((layer1_outputs(3094)) xor (layer1_outputs(7245)));
    layer2_outputs(5633) <= layer1_outputs(4566);
    layer2_outputs(5634) <= not(layer1_outputs(5274));
    layer2_outputs(5635) <= not(layer1_outputs(5461));
    layer2_outputs(5636) <= layer1_outputs(3644);
    layer2_outputs(5637) <= not(layer1_outputs(16)) or (layer1_outputs(5315));
    layer2_outputs(5638) <= layer1_outputs(4429);
    layer2_outputs(5639) <= layer1_outputs(6526);
    layer2_outputs(5640) <= (layer1_outputs(469)) and (layer1_outputs(1655));
    layer2_outputs(5641) <= layer1_outputs(1098);
    layer2_outputs(5642) <= not(layer1_outputs(760));
    layer2_outputs(5643) <= (layer1_outputs(2643)) and (layer1_outputs(5722));
    layer2_outputs(5644) <= not((layer1_outputs(3546)) or (layer1_outputs(648)));
    layer2_outputs(5645) <= layer1_outputs(5144);
    layer2_outputs(5646) <= not((layer1_outputs(2581)) or (layer1_outputs(3189)));
    layer2_outputs(5647) <= not(layer1_outputs(4729)) or (layer1_outputs(6047));
    layer2_outputs(5648) <= layer1_outputs(3555);
    layer2_outputs(5649) <= not((layer1_outputs(2122)) or (layer1_outputs(7519)));
    layer2_outputs(5650) <= '0';
    layer2_outputs(5651) <= not((layer1_outputs(1223)) or (layer1_outputs(1675)));
    layer2_outputs(5652) <= not(layer1_outputs(998));
    layer2_outputs(5653) <= layer1_outputs(6468);
    layer2_outputs(5654) <= (layer1_outputs(3828)) and not (layer1_outputs(2865));
    layer2_outputs(5655) <= not(layer1_outputs(6214));
    layer2_outputs(5656) <= not(layer1_outputs(6920)) or (layer1_outputs(3560));
    layer2_outputs(5657) <= not(layer1_outputs(4776));
    layer2_outputs(5658) <= not(layer1_outputs(1449));
    layer2_outputs(5659) <= not(layer1_outputs(7010));
    layer2_outputs(5660) <= not(layer1_outputs(3506));
    layer2_outputs(5661) <= not((layer1_outputs(6156)) or (layer1_outputs(5720)));
    layer2_outputs(5662) <= not(layer1_outputs(6944));
    layer2_outputs(5663) <= '0';
    layer2_outputs(5664) <= (layer1_outputs(4542)) and (layer1_outputs(6530));
    layer2_outputs(5665) <= not(layer1_outputs(6485)) or (layer1_outputs(3970));
    layer2_outputs(5666) <= (layer1_outputs(1437)) and (layer1_outputs(2567));
    layer2_outputs(5667) <= '1';
    layer2_outputs(5668) <= '1';
    layer2_outputs(5669) <= not((layer1_outputs(2758)) or (layer1_outputs(1340)));
    layer2_outputs(5670) <= not(layer1_outputs(2241));
    layer2_outputs(5671) <= not(layer1_outputs(2069));
    layer2_outputs(5672) <= not((layer1_outputs(1792)) and (layer1_outputs(5869)));
    layer2_outputs(5673) <= (layer1_outputs(7489)) xor (layer1_outputs(6267));
    layer2_outputs(5674) <= (layer1_outputs(1861)) or (layer1_outputs(3258));
    layer2_outputs(5675) <= not(layer1_outputs(6849));
    layer2_outputs(5676) <= not((layer1_outputs(3242)) or (layer1_outputs(3382)));
    layer2_outputs(5677) <= '1';
    layer2_outputs(5678) <= not(layer1_outputs(5796)) or (layer1_outputs(7435));
    layer2_outputs(5679) <= (layer1_outputs(5184)) and not (layer1_outputs(4288));
    layer2_outputs(5680) <= not((layer1_outputs(110)) and (layer1_outputs(6762)));
    layer2_outputs(5681) <= '1';
    layer2_outputs(5682) <= not(layer1_outputs(6719));
    layer2_outputs(5683) <= layer1_outputs(815);
    layer2_outputs(5684) <= (layer1_outputs(6864)) and not (layer1_outputs(3119));
    layer2_outputs(5685) <= not((layer1_outputs(3516)) or (layer1_outputs(5082)));
    layer2_outputs(5686) <= (layer1_outputs(3418)) and (layer1_outputs(814));
    layer2_outputs(5687) <= (layer1_outputs(6890)) and not (layer1_outputs(1265));
    layer2_outputs(5688) <= layer1_outputs(257);
    layer2_outputs(5689) <= not(layer1_outputs(7136)) or (layer1_outputs(3909));
    layer2_outputs(5690) <= not(layer1_outputs(2945)) or (layer1_outputs(5114));
    layer2_outputs(5691) <= (layer1_outputs(4216)) and (layer1_outputs(815));
    layer2_outputs(5692) <= (layer1_outputs(5370)) and (layer1_outputs(2884));
    layer2_outputs(5693) <= not((layer1_outputs(5913)) or (layer1_outputs(2370)));
    layer2_outputs(5694) <= not((layer1_outputs(6446)) xor (layer1_outputs(6443)));
    layer2_outputs(5695) <= not(layer1_outputs(891)) or (layer1_outputs(5267));
    layer2_outputs(5696) <= layer1_outputs(748);
    layer2_outputs(5697) <= not(layer1_outputs(1663));
    layer2_outputs(5698) <= (layer1_outputs(4922)) and not (layer1_outputs(3054));
    layer2_outputs(5699) <= not(layer1_outputs(7205));
    layer2_outputs(5700) <= not(layer1_outputs(627)) or (layer1_outputs(2619));
    layer2_outputs(5701) <= not(layer1_outputs(535));
    layer2_outputs(5702) <= layer1_outputs(4741);
    layer2_outputs(5703) <= (layer1_outputs(7017)) and (layer1_outputs(1179));
    layer2_outputs(5704) <= not(layer1_outputs(1343)) or (layer1_outputs(4437));
    layer2_outputs(5705) <= not(layer1_outputs(2124));
    layer2_outputs(5706) <= layer1_outputs(6403);
    layer2_outputs(5707) <= not(layer1_outputs(1605));
    layer2_outputs(5708) <= not(layer1_outputs(5674));
    layer2_outputs(5709) <= (layer1_outputs(7058)) and (layer1_outputs(5007));
    layer2_outputs(5710) <= layer1_outputs(1326);
    layer2_outputs(5711) <= not((layer1_outputs(822)) xor (layer1_outputs(5514)));
    layer2_outputs(5712) <= not(layer1_outputs(4714));
    layer2_outputs(5713) <= not(layer1_outputs(1059));
    layer2_outputs(5714) <= (layer1_outputs(484)) and (layer1_outputs(6250));
    layer2_outputs(5715) <= not(layer1_outputs(1281));
    layer2_outputs(5716) <= not(layer1_outputs(723));
    layer2_outputs(5717) <= layer1_outputs(521);
    layer2_outputs(5718) <= not(layer1_outputs(863));
    layer2_outputs(5719) <= not(layer1_outputs(7276));
    layer2_outputs(5720) <= layer1_outputs(1039);
    layer2_outputs(5721) <= layer1_outputs(6434);
    layer2_outputs(5722) <= layer1_outputs(3051);
    layer2_outputs(5723) <= (layer1_outputs(2627)) and (layer1_outputs(5973));
    layer2_outputs(5724) <= layer1_outputs(4783);
    layer2_outputs(5725) <= (layer1_outputs(1498)) xor (layer1_outputs(2680));
    layer2_outputs(5726) <= (layer1_outputs(433)) or (layer1_outputs(5864));
    layer2_outputs(5727) <= not(layer1_outputs(6670));
    layer2_outputs(5728) <= not((layer1_outputs(6906)) and (layer1_outputs(7010)));
    layer2_outputs(5729) <= not(layer1_outputs(1283));
    layer2_outputs(5730) <= not(layer1_outputs(4756)) or (layer1_outputs(5016));
    layer2_outputs(5731) <= layer1_outputs(2060);
    layer2_outputs(5732) <= not(layer1_outputs(5717));
    layer2_outputs(5733) <= not((layer1_outputs(164)) and (layer1_outputs(3821)));
    layer2_outputs(5734) <= '1';
    layer2_outputs(5735) <= not((layer1_outputs(951)) or (layer1_outputs(4716)));
    layer2_outputs(5736) <= (layer1_outputs(7496)) and (layer1_outputs(741));
    layer2_outputs(5737) <= (layer1_outputs(895)) and not (layer1_outputs(6811));
    layer2_outputs(5738) <= layer1_outputs(43);
    layer2_outputs(5739) <= not(layer1_outputs(3090));
    layer2_outputs(5740) <= not((layer1_outputs(971)) or (layer1_outputs(6748)));
    layer2_outputs(5741) <= not(layer1_outputs(6511)) or (layer1_outputs(1729));
    layer2_outputs(5742) <= (layer1_outputs(1552)) and (layer1_outputs(4968));
    layer2_outputs(5743) <= (layer1_outputs(4252)) and (layer1_outputs(2011));
    layer2_outputs(5744) <= (layer1_outputs(7453)) and (layer1_outputs(6416));
    layer2_outputs(5745) <= layer1_outputs(430);
    layer2_outputs(5746) <= '1';
    layer2_outputs(5747) <= layer1_outputs(4495);
    layer2_outputs(5748) <= not(layer1_outputs(4518));
    layer2_outputs(5749) <= not(layer1_outputs(7362));
    layer2_outputs(5750) <= layer1_outputs(3680);
    layer2_outputs(5751) <= (layer1_outputs(3814)) and (layer1_outputs(6850));
    layer2_outputs(5752) <= layer1_outputs(3121);
    layer2_outputs(5753) <= (layer1_outputs(2048)) and not (layer1_outputs(7517));
    layer2_outputs(5754) <= not(layer1_outputs(4093));
    layer2_outputs(5755) <= (layer1_outputs(1216)) and not (layer1_outputs(2032));
    layer2_outputs(5756) <= '1';
    layer2_outputs(5757) <= not(layer1_outputs(2753)) or (layer1_outputs(5949));
    layer2_outputs(5758) <= not(layer1_outputs(1013));
    layer2_outputs(5759) <= layer1_outputs(673);
    layer2_outputs(5760) <= not(layer1_outputs(7568));
    layer2_outputs(5761) <= not(layer1_outputs(3295));
    layer2_outputs(5762) <= not(layer1_outputs(2929));
    layer2_outputs(5763) <= layer1_outputs(1210);
    layer2_outputs(5764) <= not(layer1_outputs(5891));
    layer2_outputs(5765) <= '0';
    layer2_outputs(5766) <= (layer1_outputs(4172)) or (layer1_outputs(1696));
    layer2_outputs(5767) <= layer1_outputs(6968);
    layer2_outputs(5768) <= (layer1_outputs(7428)) xor (layer1_outputs(3077));
    layer2_outputs(5769) <= not(layer1_outputs(1389));
    layer2_outputs(5770) <= (layer1_outputs(7179)) or (layer1_outputs(3936));
    layer2_outputs(5771) <= not(layer1_outputs(4948));
    layer2_outputs(5772) <= (layer1_outputs(2844)) and not (layer1_outputs(2101));
    layer2_outputs(5773) <= (layer1_outputs(2275)) or (layer1_outputs(5151));
    layer2_outputs(5774) <= not(layer1_outputs(4048)) or (layer1_outputs(4240));
    layer2_outputs(5775) <= '0';
    layer2_outputs(5776) <= not(layer1_outputs(4966));
    layer2_outputs(5777) <= (layer1_outputs(757)) and not (layer1_outputs(7013));
    layer2_outputs(5778) <= layer1_outputs(1934);
    layer2_outputs(5779) <= not(layer1_outputs(3564));
    layer2_outputs(5780) <= layer1_outputs(5511);
    layer2_outputs(5781) <= not(layer1_outputs(2901)) or (layer1_outputs(4467));
    layer2_outputs(5782) <= not(layer1_outputs(1801));
    layer2_outputs(5783) <= (layer1_outputs(5716)) and not (layer1_outputs(458));
    layer2_outputs(5784) <= layer1_outputs(6453);
    layer2_outputs(5785) <= not(layer1_outputs(6050)) or (layer1_outputs(765));
    layer2_outputs(5786) <= not(layer1_outputs(4087));
    layer2_outputs(5787) <= (layer1_outputs(5074)) and (layer1_outputs(7486));
    layer2_outputs(5788) <= not(layer1_outputs(2343));
    layer2_outputs(5789) <= layer1_outputs(1307);
    layer2_outputs(5790) <= not((layer1_outputs(4938)) xor (layer1_outputs(3086)));
    layer2_outputs(5791) <= not((layer1_outputs(4616)) or (layer1_outputs(5037)));
    layer2_outputs(5792) <= layer1_outputs(2086);
    layer2_outputs(5793) <= layer1_outputs(3933);
    layer2_outputs(5794) <= (layer1_outputs(4401)) xor (layer1_outputs(2969));
    layer2_outputs(5795) <= not(layer1_outputs(3633));
    layer2_outputs(5796) <= (layer1_outputs(6285)) and not (layer1_outputs(5071));
    layer2_outputs(5797) <= (layer1_outputs(1768)) or (layer1_outputs(720));
    layer2_outputs(5798) <= (layer1_outputs(2910)) and not (layer1_outputs(2075));
    layer2_outputs(5799) <= layer1_outputs(7003);
    layer2_outputs(5800) <= (layer1_outputs(4879)) and not (layer1_outputs(1490));
    layer2_outputs(5801) <= layer1_outputs(6010);
    layer2_outputs(5802) <= layer1_outputs(5484);
    layer2_outputs(5803) <= layer1_outputs(5519);
    layer2_outputs(5804) <= not((layer1_outputs(6407)) or (layer1_outputs(1620)));
    layer2_outputs(5805) <= (layer1_outputs(2491)) and not (layer1_outputs(6494));
    layer2_outputs(5806) <= not(layer1_outputs(6119)) or (layer1_outputs(4460));
    layer2_outputs(5807) <= not(layer1_outputs(5536)) or (layer1_outputs(3128));
    layer2_outputs(5808) <= layer1_outputs(3265);
    layer2_outputs(5809) <= '1';
    layer2_outputs(5810) <= layer1_outputs(7549);
    layer2_outputs(5811) <= not((layer1_outputs(1279)) and (layer1_outputs(8)));
    layer2_outputs(5812) <= layer1_outputs(4914);
    layer2_outputs(5813) <= not((layer1_outputs(6256)) and (layer1_outputs(2918)));
    layer2_outputs(5814) <= not(layer1_outputs(803));
    layer2_outputs(5815) <= (layer1_outputs(5075)) and not (layer1_outputs(1087));
    layer2_outputs(5816) <= (layer1_outputs(2369)) and (layer1_outputs(3474));
    layer2_outputs(5817) <= layer1_outputs(2257);
    layer2_outputs(5818) <= not(layer1_outputs(1086));
    layer2_outputs(5819) <= (layer1_outputs(6121)) and not (layer1_outputs(7348));
    layer2_outputs(5820) <= '0';
    layer2_outputs(5821) <= (layer1_outputs(593)) or (layer1_outputs(5302));
    layer2_outputs(5822) <= (layer1_outputs(2266)) or (layer1_outputs(3565));
    layer2_outputs(5823) <= '0';
    layer2_outputs(5824) <= not(layer1_outputs(528)) or (layer1_outputs(3689));
    layer2_outputs(5825) <= not(layer1_outputs(989)) or (layer1_outputs(7564));
    layer2_outputs(5826) <= not(layer1_outputs(4456)) or (layer1_outputs(7556));
    layer2_outputs(5827) <= (layer1_outputs(27)) and (layer1_outputs(5250));
    layer2_outputs(5828) <= layer1_outputs(2307);
    layer2_outputs(5829) <= '0';
    layer2_outputs(5830) <= '1';
    layer2_outputs(5831) <= not((layer1_outputs(7394)) xor (layer1_outputs(2574)));
    layer2_outputs(5832) <= not((layer1_outputs(3697)) or (layer1_outputs(6816)));
    layer2_outputs(5833) <= not((layer1_outputs(2492)) or (layer1_outputs(5828)));
    layer2_outputs(5834) <= not(layer1_outputs(1026)) or (layer1_outputs(2406));
    layer2_outputs(5835) <= '0';
    layer2_outputs(5836) <= not(layer1_outputs(2524)) or (layer1_outputs(3485));
    layer2_outputs(5837) <= (layer1_outputs(3582)) and (layer1_outputs(5476));
    layer2_outputs(5838) <= not((layer1_outputs(5756)) or (layer1_outputs(389)));
    layer2_outputs(5839) <= layer1_outputs(2929);
    layer2_outputs(5840) <= not(layer1_outputs(98));
    layer2_outputs(5841) <= layer1_outputs(7294);
    layer2_outputs(5842) <= '0';
    layer2_outputs(5843) <= '0';
    layer2_outputs(5844) <= layer1_outputs(3176);
    layer2_outputs(5845) <= not((layer1_outputs(6432)) xor (layer1_outputs(984)));
    layer2_outputs(5846) <= not((layer1_outputs(4146)) and (layer1_outputs(7537)));
    layer2_outputs(5847) <= '0';
    layer2_outputs(5848) <= (layer1_outputs(2245)) and not (layer1_outputs(825));
    layer2_outputs(5849) <= not(layer1_outputs(2134)) or (layer1_outputs(5577));
    layer2_outputs(5850) <= layer1_outputs(927);
    layer2_outputs(5851) <= layer1_outputs(2903);
    layer2_outputs(5852) <= layer1_outputs(7513);
    layer2_outputs(5853) <= not((layer1_outputs(2342)) or (layer1_outputs(4508)));
    layer2_outputs(5854) <= '1';
    layer2_outputs(5855) <= not((layer1_outputs(5134)) or (layer1_outputs(3759)));
    layer2_outputs(5856) <= not((layer1_outputs(4282)) or (layer1_outputs(5186)));
    layer2_outputs(5857) <= not(layer1_outputs(3166)) or (layer1_outputs(79));
    layer2_outputs(5858) <= not(layer1_outputs(7075));
    layer2_outputs(5859) <= not(layer1_outputs(5858));
    layer2_outputs(5860) <= layer1_outputs(4767);
    layer2_outputs(5861) <= not(layer1_outputs(2562));
    layer2_outputs(5862) <= (layer1_outputs(6399)) and (layer1_outputs(7139));
    layer2_outputs(5863) <= (layer1_outputs(4198)) and not (layer1_outputs(6417));
    layer2_outputs(5864) <= not(layer1_outputs(6555)) or (layer1_outputs(87));
    layer2_outputs(5865) <= layer1_outputs(5209);
    layer2_outputs(5866) <= layer1_outputs(2299);
    layer2_outputs(5867) <= (layer1_outputs(1167)) or (layer1_outputs(676));
    layer2_outputs(5868) <= layer1_outputs(7248);
    layer2_outputs(5869) <= (layer1_outputs(7012)) and (layer1_outputs(1782));
    layer2_outputs(5870) <= not(layer1_outputs(2205));
    layer2_outputs(5871) <= not((layer1_outputs(6402)) or (layer1_outputs(5159)));
    layer2_outputs(5872) <= not(layer1_outputs(3208));
    layer2_outputs(5873) <= not((layer1_outputs(4440)) and (layer1_outputs(3956)));
    layer2_outputs(5874) <= (layer1_outputs(6705)) and not (layer1_outputs(3269));
    layer2_outputs(5875) <= layer1_outputs(2271);
    layer2_outputs(5876) <= not(layer1_outputs(2886)) or (layer1_outputs(5590));
    layer2_outputs(5877) <= not(layer1_outputs(7077));
    layer2_outputs(5878) <= (layer1_outputs(6654)) or (layer1_outputs(4588));
    layer2_outputs(5879) <= layer1_outputs(5844);
    layer2_outputs(5880) <= (layer1_outputs(187)) and (layer1_outputs(2151));
    layer2_outputs(5881) <= not(layer1_outputs(6806));
    layer2_outputs(5882) <= not((layer1_outputs(7008)) and (layer1_outputs(3563)));
    layer2_outputs(5883) <= not(layer1_outputs(341));
    layer2_outputs(5884) <= (layer1_outputs(5949)) and not (layer1_outputs(83));
    layer2_outputs(5885) <= (layer1_outputs(84)) or (layer1_outputs(4353));
    layer2_outputs(5886) <= not(layer1_outputs(3763));
    layer2_outputs(5887) <= layer1_outputs(5743);
    layer2_outputs(5888) <= layer1_outputs(36);
    layer2_outputs(5889) <= not((layer1_outputs(6957)) xor (layer1_outputs(7045)));
    layer2_outputs(5890) <= not(layer1_outputs(1548));
    layer2_outputs(5891) <= (layer1_outputs(7067)) and (layer1_outputs(914));
    layer2_outputs(5892) <= not(layer1_outputs(5606));
    layer2_outputs(5893) <= (layer1_outputs(3849)) and not (layer1_outputs(5750));
    layer2_outputs(5894) <= not(layer1_outputs(4721));
    layer2_outputs(5895) <= (layer1_outputs(5681)) and (layer1_outputs(5500));
    layer2_outputs(5896) <= not(layer1_outputs(458));
    layer2_outputs(5897) <= (layer1_outputs(2193)) or (layer1_outputs(1484));
    layer2_outputs(5898) <= not((layer1_outputs(6051)) or (layer1_outputs(4407)));
    layer2_outputs(5899) <= not((layer1_outputs(767)) and (layer1_outputs(7243)));
    layer2_outputs(5900) <= layer1_outputs(5438);
    layer2_outputs(5901) <= not(layer1_outputs(2586)) or (layer1_outputs(3751));
    layer2_outputs(5902) <= (layer1_outputs(6653)) or (layer1_outputs(6781));
    layer2_outputs(5903) <= layer1_outputs(3240);
    layer2_outputs(5904) <= (layer1_outputs(775)) and not (layer1_outputs(1894));
    layer2_outputs(5905) <= not(layer1_outputs(6370)) or (layer1_outputs(178));
    layer2_outputs(5906) <= not(layer1_outputs(4001));
    layer2_outputs(5907) <= not(layer1_outputs(4032)) or (layer1_outputs(922));
    layer2_outputs(5908) <= not(layer1_outputs(172)) or (layer1_outputs(7622));
    layer2_outputs(5909) <= not(layer1_outputs(4117));
    layer2_outputs(5910) <= (layer1_outputs(133)) or (layer1_outputs(6746));
    layer2_outputs(5911) <= layer1_outputs(4330);
    layer2_outputs(5912) <= (layer1_outputs(1781)) or (layer1_outputs(3457));
    layer2_outputs(5913) <= not(layer1_outputs(6030));
    layer2_outputs(5914) <= not(layer1_outputs(1812));
    layer2_outputs(5915) <= not(layer1_outputs(395));
    layer2_outputs(5916) <= layer1_outputs(6489);
    layer2_outputs(5917) <= not(layer1_outputs(2199)) or (layer1_outputs(385));
    layer2_outputs(5918) <= not(layer1_outputs(7043));
    layer2_outputs(5919) <= not((layer1_outputs(346)) or (layer1_outputs(5434)));
    layer2_outputs(5920) <= (layer1_outputs(487)) and not (layer1_outputs(1894));
    layer2_outputs(5921) <= not((layer1_outputs(4520)) and (layer1_outputs(2596)));
    layer2_outputs(5922) <= not(layer1_outputs(6273)) or (layer1_outputs(3714));
    layer2_outputs(5923) <= not((layer1_outputs(1986)) and (layer1_outputs(2481)));
    layer2_outputs(5924) <= (layer1_outputs(1262)) and (layer1_outputs(3398));
    layer2_outputs(5925) <= (layer1_outputs(4674)) and not (layer1_outputs(7645));
    layer2_outputs(5926) <= not((layer1_outputs(3994)) or (layer1_outputs(1564)));
    layer2_outputs(5927) <= not((layer1_outputs(7678)) and (layer1_outputs(5745)));
    layer2_outputs(5928) <= (layer1_outputs(3140)) and (layer1_outputs(6146));
    layer2_outputs(5929) <= not(layer1_outputs(6549)) or (layer1_outputs(6740));
    layer2_outputs(5930) <= layer1_outputs(7021);
    layer2_outputs(5931) <= layer1_outputs(2875);
    layer2_outputs(5932) <= (layer1_outputs(3480)) and not (layer1_outputs(6511));
    layer2_outputs(5933) <= '0';
    layer2_outputs(5934) <= (layer1_outputs(3080)) and not (layer1_outputs(6965));
    layer2_outputs(5935) <= not(layer1_outputs(4023));
    layer2_outputs(5936) <= not(layer1_outputs(3548));
    layer2_outputs(5937) <= not((layer1_outputs(5225)) xor (layer1_outputs(6463)));
    layer2_outputs(5938) <= layer1_outputs(6214);
    layer2_outputs(5939) <= layer1_outputs(5367);
    layer2_outputs(5940) <= layer1_outputs(3032);
    layer2_outputs(5941) <= not(layer1_outputs(873)) or (layer1_outputs(1301));
    layer2_outputs(5942) <= '0';
    layer2_outputs(5943) <= not(layer1_outputs(2171));
    layer2_outputs(5944) <= layer1_outputs(6621);
    layer2_outputs(5945) <= not(layer1_outputs(4392)) or (layer1_outputs(7283));
    layer2_outputs(5946) <= (layer1_outputs(7379)) and (layer1_outputs(3173));
    layer2_outputs(5947) <= not(layer1_outputs(2086));
    layer2_outputs(5948) <= layer1_outputs(3549);
    layer2_outputs(5949) <= not(layer1_outputs(1177));
    layer2_outputs(5950) <= layer1_outputs(3762);
    layer2_outputs(5951) <= not(layer1_outputs(5309));
    layer2_outputs(5952) <= not(layer1_outputs(6617));
    layer2_outputs(5953) <= layer1_outputs(2602);
    layer2_outputs(5954) <= not(layer1_outputs(1911));
    layer2_outputs(5955) <= layer1_outputs(1348);
    layer2_outputs(5956) <= not(layer1_outputs(3197));
    layer2_outputs(5957) <= (layer1_outputs(6918)) and (layer1_outputs(3988));
    layer2_outputs(5958) <= not(layer1_outputs(193));
    layer2_outputs(5959) <= not((layer1_outputs(2928)) or (layer1_outputs(2501)));
    layer2_outputs(5960) <= not(layer1_outputs(638)) or (layer1_outputs(7135));
    layer2_outputs(5961) <= (layer1_outputs(1023)) and not (layer1_outputs(3446));
    layer2_outputs(5962) <= '0';
    layer2_outputs(5963) <= layer1_outputs(3671);
    layer2_outputs(5964) <= not((layer1_outputs(5016)) and (layer1_outputs(2394)));
    layer2_outputs(5965) <= not(layer1_outputs(5075)) or (layer1_outputs(3732));
    layer2_outputs(5966) <= layer1_outputs(5888);
    layer2_outputs(5967) <= not(layer1_outputs(7063));
    layer2_outputs(5968) <= not((layer1_outputs(1381)) or (layer1_outputs(2911)));
    layer2_outputs(5969) <= not(layer1_outputs(5962)) or (layer1_outputs(413));
    layer2_outputs(5970) <= not(layer1_outputs(3292));
    layer2_outputs(5971) <= not(layer1_outputs(1614));
    layer2_outputs(5972) <= (layer1_outputs(5870)) and (layer1_outputs(4976));
    layer2_outputs(5973) <= layer1_outputs(5402);
    layer2_outputs(5974) <= not(layer1_outputs(3474)) or (layer1_outputs(7197));
    layer2_outputs(5975) <= not(layer1_outputs(2203));
    layer2_outputs(5976) <= not(layer1_outputs(3154));
    layer2_outputs(5977) <= (layer1_outputs(363)) and (layer1_outputs(1107));
    layer2_outputs(5978) <= not(layer1_outputs(3249)) or (layer1_outputs(904));
    layer2_outputs(5979) <= layer1_outputs(4193);
    layer2_outputs(5980) <= not(layer1_outputs(4424)) or (layer1_outputs(6215));
    layer2_outputs(5981) <= not(layer1_outputs(4071));
    layer2_outputs(5982) <= not(layer1_outputs(5464));
    layer2_outputs(5983) <= not((layer1_outputs(201)) or (layer1_outputs(3194)));
    layer2_outputs(5984) <= (layer1_outputs(6756)) and not (layer1_outputs(6603));
    layer2_outputs(5985) <= (layer1_outputs(6490)) xor (layer1_outputs(4343));
    layer2_outputs(5986) <= layer1_outputs(6097);
    layer2_outputs(5987) <= layer1_outputs(6880);
    layer2_outputs(5988) <= not((layer1_outputs(1704)) or (layer1_outputs(384)));
    layer2_outputs(5989) <= (layer1_outputs(3951)) or (layer1_outputs(7035));
    layer2_outputs(5990) <= layer1_outputs(91);
    layer2_outputs(5991) <= not(layer1_outputs(1158)) or (layer1_outputs(7603));
    layer2_outputs(5992) <= not(layer1_outputs(6919)) or (layer1_outputs(6164));
    layer2_outputs(5993) <= not(layer1_outputs(2273));
    layer2_outputs(5994) <= not(layer1_outputs(3852));
    layer2_outputs(5995) <= (layer1_outputs(3202)) and not (layer1_outputs(5867));
    layer2_outputs(5996) <= '1';
    layer2_outputs(5997) <= not(layer1_outputs(5497));
    layer2_outputs(5998) <= layer1_outputs(5526);
    layer2_outputs(5999) <= not(layer1_outputs(4759)) or (layer1_outputs(6491));
    layer2_outputs(6000) <= (layer1_outputs(3642)) or (layer1_outputs(3661));
    layer2_outputs(6001) <= layer1_outputs(690);
    layer2_outputs(6002) <= not(layer1_outputs(3404));
    layer2_outputs(6003) <= layer1_outputs(3653);
    layer2_outputs(6004) <= not(layer1_outputs(3481)) or (layer1_outputs(6748));
    layer2_outputs(6005) <= not((layer1_outputs(1121)) and (layer1_outputs(1786)));
    layer2_outputs(6006) <= not(layer1_outputs(6738)) or (layer1_outputs(1038));
    layer2_outputs(6007) <= not(layer1_outputs(575)) or (layer1_outputs(4194));
    layer2_outputs(6008) <= (layer1_outputs(2467)) or (layer1_outputs(3451));
    layer2_outputs(6009) <= not(layer1_outputs(1384));
    layer2_outputs(6010) <= (layer1_outputs(2819)) and not (layer1_outputs(1787));
    layer2_outputs(6011) <= layer1_outputs(6693);
    layer2_outputs(6012) <= not(layer1_outputs(6912));
    layer2_outputs(6013) <= layer1_outputs(531);
    layer2_outputs(6014) <= (layer1_outputs(4309)) and not (layer1_outputs(3829));
    layer2_outputs(6015) <= not(layer1_outputs(3182));
    layer2_outputs(6016) <= (layer1_outputs(4923)) or (layer1_outputs(1029));
    layer2_outputs(6017) <= layer1_outputs(6040);
    layer2_outputs(6018) <= not(layer1_outputs(885)) or (layer1_outputs(1956));
    layer2_outputs(6019) <= layer1_outputs(1833);
    layer2_outputs(6020) <= not(layer1_outputs(1096)) or (layer1_outputs(206));
    layer2_outputs(6021) <= not(layer1_outputs(1399)) or (layer1_outputs(3781));
    layer2_outputs(6022) <= not(layer1_outputs(3971));
    layer2_outputs(6023) <= not((layer1_outputs(4726)) xor (layer1_outputs(6743)));
    layer2_outputs(6024) <= layer1_outputs(1856);
    layer2_outputs(6025) <= not(layer1_outputs(4091));
    layer2_outputs(6026) <= (layer1_outputs(6926)) and not (layer1_outputs(528));
    layer2_outputs(6027) <= (layer1_outputs(686)) and not (layer1_outputs(539));
    layer2_outputs(6028) <= not((layer1_outputs(2460)) or (layer1_outputs(5865)));
    layer2_outputs(6029) <= not(layer1_outputs(2625));
    layer2_outputs(6030) <= not(layer1_outputs(6041));
    layer2_outputs(6031) <= not((layer1_outputs(903)) xor (layer1_outputs(705)));
    layer2_outputs(6032) <= layer1_outputs(2831);
    layer2_outputs(6033) <= not(layer1_outputs(5835));
    layer2_outputs(6034) <= layer1_outputs(3935);
    layer2_outputs(6035) <= not(layer1_outputs(1715));
    layer2_outputs(6036) <= (layer1_outputs(1775)) and not (layer1_outputs(112));
    layer2_outputs(6037) <= '0';
    layer2_outputs(6038) <= not(layer1_outputs(858));
    layer2_outputs(6039) <= not(layer1_outputs(6795));
    layer2_outputs(6040) <= not((layer1_outputs(5487)) xor (layer1_outputs(2772)));
    layer2_outputs(6041) <= layer1_outputs(2333);
    layer2_outputs(6042) <= not(layer1_outputs(1891));
    layer2_outputs(6043) <= (layer1_outputs(37)) and not (layer1_outputs(999));
    layer2_outputs(6044) <= not(layer1_outputs(2757)) or (layer1_outputs(5486));
    layer2_outputs(6045) <= layer1_outputs(6319);
    layer2_outputs(6046) <= layer1_outputs(3664);
    layer2_outputs(6047) <= layer1_outputs(6587);
    layer2_outputs(6048) <= (layer1_outputs(3607)) and not (layer1_outputs(3864));
    layer2_outputs(6049) <= not(layer1_outputs(6320));
    layer2_outputs(6050) <= '1';
    layer2_outputs(6051) <= (layer1_outputs(5343)) or (layer1_outputs(2343));
    layer2_outputs(6052) <= not(layer1_outputs(2081));
    layer2_outputs(6053) <= not(layer1_outputs(6515));
    layer2_outputs(6054) <= layer1_outputs(96);
    layer2_outputs(6055) <= not(layer1_outputs(7293));
    layer2_outputs(6056) <= not(layer1_outputs(4629));
    layer2_outputs(6057) <= layer1_outputs(50);
    layer2_outputs(6058) <= not((layer1_outputs(4655)) xor (layer1_outputs(4781)));
    layer2_outputs(6059) <= layer1_outputs(5945);
    layer2_outputs(6060) <= (layer1_outputs(202)) and not (layer1_outputs(5829));
    layer2_outputs(6061) <= (layer1_outputs(5748)) and not (layer1_outputs(1483));
    layer2_outputs(6062) <= not(layer1_outputs(4312)) or (layer1_outputs(5725));
    layer2_outputs(6063) <= '1';
    layer2_outputs(6064) <= not(layer1_outputs(3539)) or (layer1_outputs(7122));
    layer2_outputs(6065) <= not((layer1_outputs(5592)) xor (layer1_outputs(2234)));
    layer2_outputs(6066) <= (layer1_outputs(896)) and (layer1_outputs(1699));
    layer2_outputs(6067) <= not((layer1_outputs(2191)) and (layer1_outputs(5868)));
    layer2_outputs(6068) <= not(layer1_outputs(7235));
    layer2_outputs(6069) <= (layer1_outputs(4246)) and not (layer1_outputs(5120));
    layer2_outputs(6070) <= (layer1_outputs(3713)) or (layer1_outputs(4267));
    layer2_outputs(6071) <= (layer1_outputs(1437)) and not (layer1_outputs(1267));
    layer2_outputs(6072) <= not(layer1_outputs(730));
    layer2_outputs(6073) <= not(layer1_outputs(966)) or (layer1_outputs(3306));
    layer2_outputs(6074) <= (layer1_outputs(3583)) and not (layer1_outputs(194));
    layer2_outputs(6075) <= layer1_outputs(3203);
    layer2_outputs(6076) <= not((layer1_outputs(7100)) or (layer1_outputs(5019)));
    layer2_outputs(6077) <= not(layer1_outputs(2174));
    layer2_outputs(6078) <= not(layer1_outputs(6788)) or (layer1_outputs(3724));
    layer2_outputs(6079) <= not(layer1_outputs(2676));
    layer2_outputs(6080) <= '0';
    layer2_outputs(6081) <= (layer1_outputs(3640)) and not (layer1_outputs(6911));
    layer2_outputs(6082) <= not((layer1_outputs(851)) xor (layer1_outputs(3142)));
    layer2_outputs(6083) <= layer1_outputs(1272);
    layer2_outputs(6084) <= (layer1_outputs(917)) and (layer1_outputs(1021));
    layer2_outputs(6085) <= not(layer1_outputs(7450));
    layer2_outputs(6086) <= not(layer1_outputs(1968)) or (layer1_outputs(4769));
    layer2_outputs(6087) <= layer1_outputs(522);
    layer2_outputs(6088) <= (layer1_outputs(2268)) and not (layer1_outputs(293));
    layer2_outputs(6089) <= '1';
    layer2_outputs(6090) <= (layer1_outputs(2185)) and not (layer1_outputs(6461));
    layer2_outputs(6091) <= (layer1_outputs(2711)) or (layer1_outputs(6774));
    layer2_outputs(6092) <= not(layer1_outputs(7065));
    layer2_outputs(6093) <= (layer1_outputs(5916)) xor (layer1_outputs(5404));
    layer2_outputs(6094) <= layer1_outputs(3250);
    layer2_outputs(6095) <= (layer1_outputs(7100)) and not (layer1_outputs(4160));
    layer2_outputs(6096) <= not(layer1_outputs(3966));
    layer2_outputs(6097) <= not(layer1_outputs(7405));
    layer2_outputs(6098) <= not(layer1_outputs(7073));
    layer2_outputs(6099) <= not(layer1_outputs(907));
    layer2_outputs(6100) <= layer1_outputs(7492);
    layer2_outputs(6101) <= (layer1_outputs(5880)) and not (layer1_outputs(1329));
    layer2_outputs(6102) <= not(layer1_outputs(4270));
    layer2_outputs(6103) <= layer1_outputs(698);
    layer2_outputs(6104) <= layer1_outputs(2123);
    layer2_outputs(6105) <= not(layer1_outputs(40)) or (layer1_outputs(3884));
    layer2_outputs(6106) <= (layer1_outputs(5440)) or (layer1_outputs(4070));
    layer2_outputs(6107) <= layer1_outputs(3064);
    layer2_outputs(6108) <= not(layer1_outputs(7501));
    layer2_outputs(6109) <= layer1_outputs(6536);
    layer2_outputs(6110) <= not(layer1_outputs(5835)) or (layer1_outputs(3343));
    layer2_outputs(6111) <= layer1_outputs(101);
    layer2_outputs(6112) <= (layer1_outputs(4249)) and not (layer1_outputs(389));
    layer2_outputs(6113) <= '0';
    layer2_outputs(6114) <= '1';
    layer2_outputs(6115) <= layer1_outputs(7463);
    layer2_outputs(6116) <= not(layer1_outputs(943)) or (layer1_outputs(2417));
    layer2_outputs(6117) <= not(layer1_outputs(5090));
    layer2_outputs(6118) <= layer1_outputs(5432);
    layer2_outputs(6119) <= not((layer1_outputs(2764)) and (layer1_outputs(7110)));
    layer2_outputs(6120) <= '1';
    layer2_outputs(6121) <= (layer1_outputs(5742)) and (layer1_outputs(2957));
    layer2_outputs(6122) <= (layer1_outputs(111)) and (layer1_outputs(2607));
    layer2_outputs(6123) <= not(layer1_outputs(1294));
    layer2_outputs(6124) <= '0';
    layer2_outputs(6125) <= '0';
    layer2_outputs(6126) <= not(layer1_outputs(6252));
    layer2_outputs(6127) <= (layer1_outputs(3447)) and (layer1_outputs(7146));
    layer2_outputs(6128) <= not((layer1_outputs(5276)) xor (layer1_outputs(6935)));
    layer2_outputs(6129) <= (layer1_outputs(370)) and (layer1_outputs(5979));
    layer2_outputs(6130) <= not(layer1_outputs(1321));
    layer2_outputs(6131) <= not((layer1_outputs(1062)) or (layer1_outputs(5813)));
    layer2_outputs(6132) <= not(layer1_outputs(6637)) or (layer1_outputs(3782));
    layer2_outputs(6133) <= layer1_outputs(4161);
    layer2_outputs(6134) <= not(layer1_outputs(5755));
    layer2_outputs(6135) <= not(layer1_outputs(637)) or (layer1_outputs(2260));
    layer2_outputs(6136) <= '0';
    layer2_outputs(6137) <= layer1_outputs(5165);
    layer2_outputs(6138) <= layer1_outputs(3588);
    layer2_outputs(6139) <= not(layer1_outputs(4428));
    layer2_outputs(6140) <= not(layer1_outputs(6103)) or (layer1_outputs(4490));
    layer2_outputs(6141) <= not(layer1_outputs(4205));
    layer2_outputs(6142) <= not(layer1_outputs(5398)) or (layer1_outputs(4924));
    layer2_outputs(6143) <= not((layer1_outputs(1020)) xor (layer1_outputs(1906)));
    layer2_outputs(6144) <= '0';
    layer2_outputs(6145) <= layer1_outputs(4416);
    layer2_outputs(6146) <= not(layer1_outputs(4044));
    layer2_outputs(6147) <= not(layer1_outputs(2440));
    layer2_outputs(6148) <= layer1_outputs(1271);
    layer2_outputs(6149) <= not(layer1_outputs(395));
    layer2_outputs(6150) <= not(layer1_outputs(7174));
    layer2_outputs(6151) <= (layer1_outputs(4667)) or (layer1_outputs(6326));
    layer2_outputs(6152) <= (layer1_outputs(1348)) and not (layer1_outputs(6130));
    layer2_outputs(6153) <= not(layer1_outputs(3886));
    layer2_outputs(6154) <= layer1_outputs(2233);
    layer2_outputs(6155) <= layer1_outputs(679);
    layer2_outputs(6156) <= (layer1_outputs(3553)) and (layer1_outputs(1009));
    layer2_outputs(6157) <= (layer1_outputs(4319)) or (layer1_outputs(7568));
    layer2_outputs(6158) <= not((layer1_outputs(4336)) or (layer1_outputs(2101)));
    layer2_outputs(6159) <= (layer1_outputs(6985)) xor (layer1_outputs(2246));
    layer2_outputs(6160) <= layer1_outputs(6534);
    layer2_outputs(6161) <= not((layer1_outputs(6529)) or (layer1_outputs(6727)));
    layer2_outputs(6162) <= not((layer1_outputs(2853)) or (layer1_outputs(1040)));
    layer2_outputs(6163) <= (layer1_outputs(2502)) or (layer1_outputs(4229));
    layer2_outputs(6164) <= not((layer1_outputs(5893)) or (layer1_outputs(4840)));
    layer2_outputs(6165) <= not(layer1_outputs(2644)) or (layer1_outputs(1326));
    layer2_outputs(6166) <= (layer1_outputs(7257)) and not (layer1_outputs(441));
    layer2_outputs(6167) <= (layer1_outputs(1757)) and (layer1_outputs(6437));
    layer2_outputs(6168) <= (layer1_outputs(8)) or (layer1_outputs(6451));
    layer2_outputs(6169) <= layer1_outputs(407);
    layer2_outputs(6170) <= layer1_outputs(4591);
    layer2_outputs(6171) <= (layer1_outputs(558)) or (layer1_outputs(6503));
    layer2_outputs(6172) <= not(layer1_outputs(1821)) or (layer1_outputs(895));
    layer2_outputs(6173) <= layer1_outputs(4820);
    layer2_outputs(6174) <= (layer1_outputs(3949)) and not (layer1_outputs(4425));
    layer2_outputs(6175) <= (layer1_outputs(1467)) and (layer1_outputs(848));
    layer2_outputs(6176) <= not(layer1_outputs(3913)) or (layer1_outputs(4338));
    layer2_outputs(6177) <= '0';
    layer2_outputs(6178) <= not((layer1_outputs(4410)) or (layer1_outputs(4385)));
    layer2_outputs(6179) <= not(layer1_outputs(1980));
    layer2_outputs(6180) <= layer1_outputs(2385);
    layer2_outputs(6181) <= (layer1_outputs(3500)) or (layer1_outputs(1355));
    layer2_outputs(6182) <= layer1_outputs(868);
    layer2_outputs(6183) <= not((layer1_outputs(3285)) or (layer1_outputs(833)));
    layer2_outputs(6184) <= (layer1_outputs(4756)) and not (layer1_outputs(1450));
    layer2_outputs(6185) <= not(layer1_outputs(3411));
    layer2_outputs(6186) <= not((layer1_outputs(3341)) or (layer1_outputs(5419)));
    layer2_outputs(6187) <= layer1_outputs(3436);
    layer2_outputs(6188) <= not((layer1_outputs(4186)) and (layer1_outputs(4701)));
    layer2_outputs(6189) <= '1';
    layer2_outputs(6190) <= (layer1_outputs(365)) and not (layer1_outputs(1671));
    layer2_outputs(6191) <= layer1_outputs(3036);
    layer2_outputs(6192) <= layer1_outputs(5072);
    layer2_outputs(6193) <= (layer1_outputs(1614)) or (layer1_outputs(828));
    layer2_outputs(6194) <= layer1_outputs(1390);
    layer2_outputs(6195) <= not(layer1_outputs(3075));
    layer2_outputs(6196) <= (layer1_outputs(3856)) and not (layer1_outputs(6977));
    layer2_outputs(6197) <= (layer1_outputs(3015)) and not (layer1_outputs(6514));
    layer2_outputs(6198) <= layer1_outputs(1296);
    layer2_outputs(6199) <= layer1_outputs(5005);
    layer2_outputs(6200) <= (layer1_outputs(3432)) and (layer1_outputs(2024));
    layer2_outputs(6201) <= not(layer1_outputs(5339));
    layer2_outputs(6202) <= (layer1_outputs(844)) or (layer1_outputs(1789));
    layer2_outputs(6203) <= not((layer1_outputs(1235)) and (layer1_outputs(3354)));
    layer2_outputs(6204) <= (layer1_outputs(1484)) and not (layer1_outputs(4862));
    layer2_outputs(6205) <= not((layer1_outputs(7464)) or (layer1_outputs(4157)));
    layer2_outputs(6206) <= (layer1_outputs(5563)) and not (layer1_outputs(2198));
    layer2_outputs(6207) <= '1';
    layer2_outputs(6208) <= layer1_outputs(2530);
    layer2_outputs(6209) <= (layer1_outputs(5833)) or (layer1_outputs(2743));
    layer2_outputs(6210) <= not(layer1_outputs(5373));
    layer2_outputs(6211) <= not(layer1_outputs(2916)) or (layer1_outputs(4870));
    layer2_outputs(6212) <= not((layer1_outputs(7309)) or (layer1_outputs(3745)));
    layer2_outputs(6213) <= (layer1_outputs(5171)) xor (layer1_outputs(3215));
    layer2_outputs(6214) <= '0';
    layer2_outputs(6215) <= layer1_outputs(5034);
    layer2_outputs(6216) <= (layer1_outputs(1988)) and (layer1_outputs(2169));
    layer2_outputs(6217) <= not(layer1_outputs(3015));
    layer2_outputs(6218) <= (layer1_outputs(6744)) xor (layer1_outputs(4972));
    layer2_outputs(6219) <= '1';
    layer2_outputs(6220) <= (layer1_outputs(1333)) and (layer1_outputs(5725));
    layer2_outputs(6221) <= not((layer1_outputs(2940)) or (layer1_outputs(5168)));
    layer2_outputs(6222) <= (layer1_outputs(2404)) or (layer1_outputs(4689));
    layer2_outputs(6223) <= not(layer1_outputs(728)) or (layer1_outputs(5798));
    layer2_outputs(6224) <= (layer1_outputs(1241)) and not (layer1_outputs(6268));
    layer2_outputs(6225) <= not(layer1_outputs(2365));
    layer2_outputs(6226) <= layer1_outputs(2296);
    layer2_outputs(6227) <= (layer1_outputs(1088)) and not (layer1_outputs(2422));
    layer2_outputs(6228) <= layer1_outputs(3438);
    layer2_outputs(6229) <= (layer1_outputs(7584)) and (layer1_outputs(1130));
    layer2_outputs(6230) <= not((layer1_outputs(7030)) and (layer1_outputs(4627)));
    layer2_outputs(6231) <= not((layer1_outputs(6123)) and (layer1_outputs(1661)));
    layer2_outputs(6232) <= layer1_outputs(7106);
    layer2_outputs(6233) <= '0';
    layer2_outputs(6234) <= not((layer1_outputs(3187)) and (layer1_outputs(1378)));
    layer2_outputs(6235) <= not(layer1_outputs(4950));
    layer2_outputs(6236) <= not((layer1_outputs(3497)) or (layer1_outputs(2697)));
    layer2_outputs(6237) <= (layer1_outputs(4775)) and not (layer1_outputs(4438));
    layer2_outputs(6238) <= (layer1_outputs(2414)) and (layer1_outputs(6752));
    layer2_outputs(6239) <= not(layer1_outputs(6659)) or (layer1_outputs(4020));
    layer2_outputs(6240) <= not(layer1_outputs(1545)) or (layer1_outputs(3148));
    layer2_outputs(6241) <= '1';
    layer2_outputs(6242) <= '1';
    layer2_outputs(6243) <= '0';
    layer2_outputs(6244) <= not(layer1_outputs(341));
    layer2_outputs(6245) <= '0';
    layer2_outputs(6246) <= not(layer1_outputs(4374));
    layer2_outputs(6247) <= (layer1_outputs(4745)) and (layer1_outputs(3126));
    layer2_outputs(6248) <= (layer1_outputs(2458)) and not (layer1_outputs(2897));
    layer2_outputs(6249) <= layer1_outputs(6774);
    layer2_outputs(6250) <= (layer1_outputs(709)) or (layer1_outputs(2024));
    layer2_outputs(6251) <= '0';
    layer2_outputs(6252) <= '0';
    layer2_outputs(6253) <= layer1_outputs(7193);
    layer2_outputs(6254) <= not(layer1_outputs(7436));
    layer2_outputs(6255) <= not((layer1_outputs(938)) or (layer1_outputs(2744)));
    layer2_outputs(6256) <= not(layer1_outputs(2892));
    layer2_outputs(6257) <= not(layer1_outputs(4924));
    layer2_outputs(6258) <= not(layer1_outputs(7505)) or (layer1_outputs(4003));
    layer2_outputs(6259) <= not(layer1_outputs(4853)) or (layer1_outputs(768));
    layer2_outputs(6260) <= layer1_outputs(5349);
    layer2_outputs(6261) <= layer1_outputs(5984);
    layer2_outputs(6262) <= not(layer1_outputs(2936));
    layer2_outputs(6263) <= not(layer1_outputs(4375));
    layer2_outputs(6264) <= '1';
    layer2_outputs(6265) <= (layer1_outputs(54)) and not (layer1_outputs(3508));
    layer2_outputs(6266) <= layer1_outputs(4012);
    layer2_outputs(6267) <= not(layer1_outputs(4426));
    layer2_outputs(6268) <= layer1_outputs(7676);
    layer2_outputs(6269) <= not(layer1_outputs(1884)) or (layer1_outputs(3766));
    layer2_outputs(6270) <= not(layer1_outputs(82));
    layer2_outputs(6271) <= not(layer1_outputs(1787)) or (layer1_outputs(6447));
    layer2_outputs(6272) <= (layer1_outputs(5704)) and not (layer1_outputs(2709));
    layer2_outputs(6273) <= not(layer1_outputs(6578)) or (layer1_outputs(5185));
    layer2_outputs(6274) <= layer1_outputs(4178);
    layer2_outputs(6275) <= layer1_outputs(1865);
    layer2_outputs(6276) <= layer1_outputs(2027);
    layer2_outputs(6277) <= not(layer1_outputs(5293));
    layer2_outputs(6278) <= not(layer1_outputs(57)) or (layer1_outputs(5808));
    layer2_outputs(6279) <= not(layer1_outputs(6220));
    layer2_outputs(6280) <= not((layer1_outputs(6010)) or (layer1_outputs(4063)));
    layer2_outputs(6281) <= not(layer1_outputs(6845));
    layer2_outputs(6282) <= '1';
    layer2_outputs(6283) <= not(layer1_outputs(1021));
    layer2_outputs(6284) <= not(layer1_outputs(3975)) or (layer1_outputs(5724));
    layer2_outputs(6285) <= layer1_outputs(5381);
    layer2_outputs(6286) <= '1';
    layer2_outputs(6287) <= layer1_outputs(2090);
    layer2_outputs(6288) <= (layer1_outputs(892)) xor (layer1_outputs(816));
    layer2_outputs(6289) <= '1';
    layer2_outputs(6290) <= not(layer1_outputs(2167));
    layer2_outputs(6291) <= '0';
    layer2_outputs(6292) <= layer1_outputs(3682);
    layer2_outputs(6293) <= layer1_outputs(5069);
    layer2_outputs(6294) <= (layer1_outputs(5729)) or (layer1_outputs(7175));
    layer2_outputs(6295) <= layer1_outputs(7595);
    layer2_outputs(6296) <= not(layer1_outputs(6067));
    layer2_outputs(6297) <= not((layer1_outputs(4584)) xor (layer1_outputs(4719)));
    layer2_outputs(6298) <= layer1_outputs(3996);
    layer2_outputs(6299) <= (layer1_outputs(3577)) and not (layer1_outputs(1529));
    layer2_outputs(6300) <= layer1_outputs(5119);
    layer2_outputs(6301) <= not(layer1_outputs(5706));
    layer2_outputs(6302) <= '0';
    layer2_outputs(6303) <= layer1_outputs(7487);
    layer2_outputs(6304) <= not(layer1_outputs(7210));
    layer2_outputs(6305) <= (layer1_outputs(3836)) or (layer1_outputs(4386));
    layer2_outputs(6306) <= layer1_outputs(777);
    layer2_outputs(6307) <= layer1_outputs(7103);
    layer2_outputs(6308) <= not(layer1_outputs(7547)) or (layer1_outputs(2828));
    layer2_outputs(6309) <= not((layer1_outputs(4368)) or (layer1_outputs(1945)));
    layer2_outputs(6310) <= not(layer1_outputs(2363));
    layer2_outputs(6311) <= (layer1_outputs(4320)) and not (layer1_outputs(6491));
    layer2_outputs(6312) <= not(layer1_outputs(3234));
    layer2_outputs(6313) <= not(layer1_outputs(643)) or (layer1_outputs(5002));
    layer2_outputs(6314) <= '0';
    layer2_outputs(6315) <= not(layer1_outputs(6868)) or (layer1_outputs(4659));
    layer2_outputs(6316) <= not(layer1_outputs(7311));
    layer2_outputs(6317) <= '1';
    layer2_outputs(6318) <= '1';
    layer2_outputs(6319) <= not(layer1_outputs(3226));
    layer2_outputs(6320) <= layer1_outputs(493);
    layer2_outputs(6321) <= not((layer1_outputs(4378)) or (layer1_outputs(6595)));
    layer2_outputs(6322) <= '0';
    layer2_outputs(6323) <= layer1_outputs(4089);
    layer2_outputs(6324) <= not((layer1_outputs(3192)) or (layer1_outputs(3876)));
    layer2_outputs(6325) <= layer1_outputs(1421);
    layer2_outputs(6326) <= not(layer1_outputs(6664));
    layer2_outputs(6327) <= not((layer1_outputs(5254)) or (layer1_outputs(5764)));
    layer2_outputs(6328) <= not(layer1_outputs(2958));
    layer2_outputs(6329) <= not(layer1_outputs(3062));
    layer2_outputs(6330) <= not((layer1_outputs(803)) or (layer1_outputs(3745)));
    layer2_outputs(6331) <= not(layer1_outputs(1046));
    layer2_outputs(6332) <= not(layer1_outputs(1162)) or (layer1_outputs(4204));
    layer2_outputs(6333) <= layer1_outputs(5226);
    layer2_outputs(6334) <= not(layer1_outputs(11));
    layer2_outputs(6335) <= '1';
    layer2_outputs(6336) <= layer1_outputs(5032);
    layer2_outputs(6337) <= not(layer1_outputs(5928)) or (layer1_outputs(7218));
    layer2_outputs(6338) <= not(layer1_outputs(2174));
    layer2_outputs(6339) <= not((layer1_outputs(5065)) or (layer1_outputs(5902)));
    layer2_outputs(6340) <= layer1_outputs(6696);
    layer2_outputs(6341) <= not((layer1_outputs(28)) and (layer1_outputs(6081)));
    layer2_outputs(6342) <= not(layer1_outputs(6901));
    layer2_outputs(6343) <= not(layer1_outputs(5605));
    layer2_outputs(6344) <= (layer1_outputs(3462)) and (layer1_outputs(5364));
    layer2_outputs(6345) <= (layer1_outputs(1325)) xor (layer1_outputs(3056));
    layer2_outputs(6346) <= not(layer1_outputs(3287)) or (layer1_outputs(4387));
    layer2_outputs(6347) <= layer1_outputs(4046);
    layer2_outputs(6348) <= layer1_outputs(6964);
    layer2_outputs(6349) <= (layer1_outputs(4694)) and not (layer1_outputs(7118));
    layer2_outputs(6350) <= not((layer1_outputs(5562)) and (layer1_outputs(2755)));
    layer2_outputs(6351) <= not((layer1_outputs(1839)) or (layer1_outputs(6760)));
    layer2_outputs(6352) <= not((layer1_outputs(7374)) and (layer1_outputs(144)));
    layer2_outputs(6353) <= not(layer1_outputs(7231)) or (layer1_outputs(5380));
    layer2_outputs(6354) <= not((layer1_outputs(4913)) or (layer1_outputs(5324)));
    layer2_outputs(6355) <= not(layer1_outputs(7644)) or (layer1_outputs(1941));
    layer2_outputs(6356) <= not(layer1_outputs(1705));
    layer2_outputs(6357) <= '1';
    layer2_outputs(6358) <= not(layer1_outputs(4513));
    layer2_outputs(6359) <= (layer1_outputs(1089)) and not (layer1_outputs(410));
    layer2_outputs(6360) <= layer1_outputs(1577);
    layer2_outputs(6361) <= (layer1_outputs(5983)) and not (layer1_outputs(4150));
    layer2_outputs(6362) <= not(layer1_outputs(2338)) or (layer1_outputs(2463));
    layer2_outputs(6363) <= not((layer1_outputs(473)) or (layer1_outputs(2753)));
    layer2_outputs(6364) <= layer1_outputs(6684);
    layer2_outputs(6365) <= layer1_outputs(6319);
    layer2_outputs(6366) <= (layer1_outputs(5987)) and not (layer1_outputs(5012));
    layer2_outputs(6367) <= not(layer1_outputs(2578));
    layer2_outputs(6368) <= (layer1_outputs(1264)) and not (layer1_outputs(6356));
    layer2_outputs(6369) <= layer1_outputs(2);
    layer2_outputs(6370) <= not(layer1_outputs(5796));
    layer2_outputs(6371) <= (layer1_outputs(2630)) and not (layer1_outputs(4724));
    layer2_outputs(6372) <= (layer1_outputs(5069)) and (layer1_outputs(7283));
    layer2_outputs(6373) <= not(layer1_outputs(2029)) or (layer1_outputs(3197));
    layer2_outputs(6374) <= not(layer1_outputs(3071));
    layer2_outputs(6375) <= layer1_outputs(1067);
    layer2_outputs(6376) <= '1';
    layer2_outputs(6377) <= (layer1_outputs(1080)) or (layer1_outputs(1051));
    layer2_outputs(6378) <= (layer1_outputs(6809)) or (layer1_outputs(7105));
    layer2_outputs(6379) <= not(layer1_outputs(3429));
    layer2_outputs(6380) <= layer1_outputs(3038);
    layer2_outputs(6381) <= (layer1_outputs(377)) and (layer1_outputs(5648));
    layer2_outputs(6382) <= layer1_outputs(4568);
    layer2_outputs(6383) <= (layer1_outputs(224)) and (layer1_outputs(3240));
    layer2_outputs(6384) <= not(layer1_outputs(6772)) or (layer1_outputs(1956));
    layer2_outputs(6385) <= (layer1_outputs(6975)) or (layer1_outputs(393));
    layer2_outputs(6386) <= not(layer1_outputs(1921)) or (layer1_outputs(4788));
    layer2_outputs(6387) <= layer1_outputs(390);
    layer2_outputs(6388) <= not(layer1_outputs(6304));
    layer2_outputs(6389) <= '0';
    layer2_outputs(6390) <= not(layer1_outputs(3143)) or (layer1_outputs(6415));
    layer2_outputs(6391) <= not(layer1_outputs(2138)) or (layer1_outputs(7660));
    layer2_outputs(6392) <= layer1_outputs(6634);
    layer2_outputs(6393) <= not(layer1_outputs(5853)) or (layer1_outputs(4534));
    layer2_outputs(6394) <= (layer1_outputs(5515)) and (layer1_outputs(2638));
    layer2_outputs(6395) <= '0';
    layer2_outputs(6396) <= '1';
    layer2_outputs(6397) <= not(layer1_outputs(4199));
    layer2_outputs(6398) <= layer1_outputs(5101);
    layer2_outputs(6399) <= layer1_outputs(2027);
    layer2_outputs(6400) <= '1';
    layer2_outputs(6401) <= not(layer1_outputs(7630)) or (layer1_outputs(1236));
    layer2_outputs(6402) <= (layer1_outputs(1536)) and (layer1_outputs(2322));
    layer2_outputs(6403) <= (layer1_outputs(7443)) and not (layer1_outputs(1055));
    layer2_outputs(6404) <= (layer1_outputs(4170)) and (layer1_outputs(2686));
    layer2_outputs(6405) <= layer1_outputs(5735);
    layer2_outputs(6406) <= not(layer1_outputs(6917));
    layer2_outputs(6407) <= not(layer1_outputs(3760));
    layer2_outputs(6408) <= not(layer1_outputs(3480));
    layer2_outputs(6409) <= (layer1_outputs(2693)) and not (layer1_outputs(3757));
    layer2_outputs(6410) <= not(layer1_outputs(6716));
    layer2_outputs(6411) <= not(layer1_outputs(6048));
    layer2_outputs(6412) <= (layer1_outputs(1251)) and (layer1_outputs(955));
    layer2_outputs(6413) <= (layer1_outputs(5367)) and (layer1_outputs(7022));
    layer2_outputs(6414) <= not(layer1_outputs(7331));
    layer2_outputs(6415) <= (layer1_outputs(3769)) and (layer1_outputs(6124));
    layer2_outputs(6416) <= layer1_outputs(5439);
    layer2_outputs(6417) <= layer1_outputs(578);
    layer2_outputs(6418) <= not((layer1_outputs(5410)) or (layer1_outputs(3584)));
    layer2_outputs(6419) <= layer1_outputs(3835);
    layer2_outputs(6420) <= not(layer1_outputs(3607)) or (layer1_outputs(1997));
    layer2_outputs(6421) <= (layer1_outputs(4671)) and not (layer1_outputs(5742));
    layer2_outputs(6422) <= not(layer1_outputs(5565));
    layer2_outputs(6423) <= (layer1_outputs(497)) or (layer1_outputs(1278));
    layer2_outputs(6424) <= layer1_outputs(2639);
    layer2_outputs(6425) <= (layer1_outputs(7246)) and not (layer1_outputs(5252));
    layer2_outputs(6426) <= (layer1_outputs(659)) and (layer1_outputs(1971));
    layer2_outputs(6427) <= layer1_outputs(1658);
    layer2_outputs(6428) <= layer1_outputs(7041);
    layer2_outputs(6429) <= (layer1_outputs(3575)) and not (layer1_outputs(5055));
    layer2_outputs(6430) <= '0';
    layer2_outputs(6431) <= layer1_outputs(2246);
    layer2_outputs(6432) <= not(layer1_outputs(6702));
    layer2_outputs(6433) <= (layer1_outputs(7047)) and not (layer1_outputs(5656));
    layer2_outputs(6434) <= '0';
    layer2_outputs(6435) <= layer1_outputs(81);
    layer2_outputs(6436) <= layer1_outputs(6631);
    layer2_outputs(6437) <= (layer1_outputs(1628)) and not (layer1_outputs(6683));
    layer2_outputs(6438) <= not(layer1_outputs(4235)) or (layer1_outputs(1215));
    layer2_outputs(6439) <= '0';
    layer2_outputs(6440) <= not((layer1_outputs(6789)) xor (layer1_outputs(265)));
    layer2_outputs(6441) <= not(layer1_outputs(159)) or (layer1_outputs(1202));
    layer2_outputs(6442) <= (layer1_outputs(2284)) and not (layer1_outputs(5240));
    layer2_outputs(6443) <= not(layer1_outputs(6786));
    layer2_outputs(6444) <= not(layer1_outputs(5121));
    layer2_outputs(6445) <= layer1_outputs(4297);
    layer2_outputs(6446) <= not(layer1_outputs(3514));
    layer2_outputs(6447) <= not(layer1_outputs(3132)) or (layer1_outputs(5509));
    layer2_outputs(6448) <= not(layer1_outputs(4092));
    layer2_outputs(6449) <= not(layer1_outputs(2926));
    layer2_outputs(6450) <= (layer1_outputs(6452)) and (layer1_outputs(6858));
    layer2_outputs(6451) <= (layer1_outputs(4515)) and (layer1_outputs(7160));
    layer2_outputs(6452) <= not(layer1_outputs(1804));
    layer2_outputs(6453) <= '0';
    layer2_outputs(6454) <= layer1_outputs(3686);
    layer2_outputs(6455) <= not(layer1_outputs(6424)) or (layer1_outputs(6949));
    layer2_outputs(6456) <= (layer1_outputs(3949)) and not (layer1_outputs(3167));
    layer2_outputs(6457) <= not(layer1_outputs(4137)) or (layer1_outputs(3959));
    layer2_outputs(6458) <= (layer1_outputs(3843)) and (layer1_outputs(1092));
    layer2_outputs(6459) <= not(layer1_outputs(6140)) or (layer1_outputs(6755));
    layer2_outputs(6460) <= not((layer1_outputs(2944)) and (layer1_outputs(1116)));
    layer2_outputs(6461) <= (layer1_outputs(1254)) and not (layer1_outputs(2162));
    layer2_outputs(6462) <= not(layer1_outputs(3404));
    layer2_outputs(6463) <= '0';
    layer2_outputs(6464) <= not((layer1_outputs(5017)) or (layer1_outputs(1541)));
    layer2_outputs(6465) <= layer1_outputs(4213);
    layer2_outputs(6466) <= not(layer1_outputs(706)) or (layer1_outputs(6818));
    layer2_outputs(6467) <= not(layer1_outputs(7659)) or (layer1_outputs(5733));
    layer2_outputs(6468) <= (layer1_outputs(1514)) and (layer1_outputs(5274));
    layer2_outputs(6469) <= not(layer1_outputs(7064));
    layer2_outputs(6470) <= not(layer1_outputs(10)) or (layer1_outputs(4214));
    layer2_outputs(6471) <= layer1_outputs(1937);
    layer2_outputs(6472) <= '1';
    layer2_outputs(6473) <= not(layer1_outputs(5445));
    layer2_outputs(6474) <= not(layer1_outputs(1438));
    layer2_outputs(6475) <= layer1_outputs(29);
    layer2_outputs(6476) <= not(layer1_outputs(3765));
    layer2_outputs(6477) <= not(layer1_outputs(505)) or (layer1_outputs(5887));
    layer2_outputs(6478) <= not(layer1_outputs(3098)) or (layer1_outputs(7164));
    layer2_outputs(6479) <= not((layer1_outputs(5299)) or (layer1_outputs(4352)));
    layer2_outputs(6480) <= not((layer1_outputs(1274)) and (layer1_outputs(5417)));
    layer2_outputs(6481) <= not(layer1_outputs(3716));
    layer2_outputs(6482) <= layer1_outputs(5091);
    layer2_outputs(6483) <= not(layer1_outputs(2684));
    layer2_outputs(6484) <= (layer1_outputs(2297)) and not (layer1_outputs(3051));
    layer2_outputs(6485) <= not((layer1_outputs(2824)) or (layer1_outputs(7127)));
    layer2_outputs(6486) <= (layer1_outputs(6022)) xor (layer1_outputs(3855));
    layer2_outputs(6487) <= layer1_outputs(6344);
    layer2_outputs(6488) <= (layer1_outputs(411)) and (layer1_outputs(2728));
    layer2_outputs(6489) <= not(layer1_outputs(923));
    layer2_outputs(6490) <= not(layer1_outputs(4395)) or (layer1_outputs(1098));
    layer2_outputs(6491) <= not(layer1_outputs(1424));
    layer2_outputs(6492) <= layer1_outputs(3906);
    layer2_outputs(6493) <= not((layer1_outputs(3717)) and (layer1_outputs(1944)));
    layer2_outputs(6494) <= not((layer1_outputs(4081)) or (layer1_outputs(7523)));
    layer2_outputs(6495) <= (layer1_outputs(3986)) and not (layer1_outputs(2435));
    layer2_outputs(6496) <= not(layer1_outputs(297));
    layer2_outputs(6497) <= (layer1_outputs(4810)) xor (layer1_outputs(1898));
    layer2_outputs(6498) <= not(layer1_outputs(2469));
    layer2_outputs(6499) <= (layer1_outputs(1963)) and not (layer1_outputs(5424));
    layer2_outputs(6500) <= layer1_outputs(4802);
    layer2_outputs(6501) <= not((layer1_outputs(4481)) or (layer1_outputs(3737)));
    layer2_outputs(6502) <= not(layer1_outputs(331)) or (layer1_outputs(2484));
    layer2_outputs(6503) <= not((layer1_outputs(3944)) or (layer1_outputs(638)));
    layer2_outputs(6504) <= not(layer1_outputs(2867));
    layer2_outputs(6505) <= (layer1_outputs(4324)) or (layer1_outputs(842));
    layer2_outputs(6506) <= not((layer1_outputs(7332)) or (layer1_outputs(2273)));
    layer2_outputs(6507) <= not(layer1_outputs(5133));
    layer2_outputs(6508) <= not(layer1_outputs(5217)) or (layer1_outputs(1589));
    layer2_outputs(6509) <= layer1_outputs(5244);
    layer2_outputs(6510) <= not(layer1_outputs(2095)) or (layer1_outputs(3099));
    layer2_outputs(6511) <= layer1_outputs(4034);
    layer2_outputs(6512) <= (layer1_outputs(5291)) or (layer1_outputs(4514));
    layer2_outputs(6513) <= (layer1_outputs(6243)) and not (layer1_outputs(5097));
    layer2_outputs(6514) <= (layer1_outputs(6605)) and not (layer1_outputs(2741));
    layer2_outputs(6515) <= not(layer1_outputs(6628));
    layer2_outputs(6516) <= (layer1_outputs(6328)) and not (layer1_outputs(3567));
    layer2_outputs(6517) <= not(layer1_outputs(3659)) or (layer1_outputs(4522));
    layer2_outputs(6518) <= not(layer1_outputs(3278)) or (layer1_outputs(3060));
    layer2_outputs(6519) <= not(layer1_outputs(1753)) or (layer1_outputs(2845));
    layer2_outputs(6520) <= not(layer1_outputs(631));
    layer2_outputs(6521) <= layer1_outputs(1080);
    layer2_outputs(6522) <= layer1_outputs(4324);
    layer2_outputs(6523) <= (layer1_outputs(7397)) and (layer1_outputs(5589));
    layer2_outputs(6524) <= layer1_outputs(2586);
    layer2_outputs(6525) <= layer1_outputs(3570);
    layer2_outputs(6526) <= not((layer1_outputs(1865)) or (layer1_outputs(4785)));
    layer2_outputs(6527) <= not(layer1_outputs(691));
    layer2_outputs(6528) <= layer1_outputs(2588);
    layer2_outputs(6529) <= not(layer1_outputs(936));
    layer2_outputs(6530) <= '0';
    layer2_outputs(6531) <= layer1_outputs(3830);
    layer2_outputs(6532) <= not(layer1_outputs(5202));
    layer2_outputs(6533) <= not(layer1_outputs(4132));
    layer2_outputs(6534) <= not(layer1_outputs(5073)) or (layer1_outputs(222));
    layer2_outputs(6535) <= layer1_outputs(3419);
    layer2_outputs(6536) <= not((layer1_outputs(6002)) xor (layer1_outputs(2111)));
    layer2_outputs(6537) <= layer1_outputs(3683);
    layer2_outputs(6538) <= (layer1_outputs(1070)) or (layer1_outputs(1883));
    layer2_outputs(6539) <= layer1_outputs(6191);
    layer2_outputs(6540) <= '1';
    layer2_outputs(6541) <= not(layer1_outputs(1961));
    layer2_outputs(6542) <= not(layer1_outputs(3174));
    layer2_outputs(6543) <= layer1_outputs(1681);
    layer2_outputs(6544) <= (layer1_outputs(1691)) and (layer1_outputs(4822));
    layer2_outputs(6545) <= not(layer1_outputs(1017));
    layer2_outputs(6546) <= not(layer1_outputs(6810));
    layer2_outputs(6547) <= not(layer1_outputs(5223));
    layer2_outputs(6548) <= not((layer1_outputs(7186)) or (layer1_outputs(7017)));
    layer2_outputs(6549) <= not(layer1_outputs(4873));
    layer2_outputs(6550) <= not(layer1_outputs(1069));
    layer2_outputs(6551) <= not(layer1_outputs(994));
    layer2_outputs(6552) <= not(layer1_outputs(2407));
    layer2_outputs(6553) <= (layer1_outputs(5301)) and (layer1_outputs(2876));
    layer2_outputs(6554) <= layer1_outputs(1897);
    layer2_outputs(6555) <= (layer1_outputs(6340)) and not (layer1_outputs(253));
    layer2_outputs(6556) <= (layer1_outputs(5468)) and not (layer1_outputs(1799));
    layer2_outputs(6557) <= not((layer1_outputs(4007)) or (layer1_outputs(3362)));
    layer2_outputs(6558) <= (layer1_outputs(1308)) or (layer1_outputs(4712));
    layer2_outputs(6559) <= not(layer1_outputs(6906));
    layer2_outputs(6560) <= layer1_outputs(4619);
    layer2_outputs(6561) <= not((layer1_outputs(2890)) xor (layer1_outputs(4885)));
    layer2_outputs(6562) <= (layer1_outputs(4241)) xor (layer1_outputs(3435));
    layer2_outputs(6563) <= not((layer1_outputs(1850)) xor (layer1_outputs(5310)));
    layer2_outputs(6564) <= (layer1_outputs(7674)) or (layer1_outputs(2102));
    layer2_outputs(6565) <= not(layer1_outputs(3950));
    layer2_outputs(6566) <= not((layer1_outputs(3333)) and (layer1_outputs(5078)));
    layer2_outputs(6567) <= not(layer1_outputs(55));
    layer2_outputs(6568) <= (layer1_outputs(6518)) or (layer1_outputs(4082));
    layer2_outputs(6569) <= layer1_outputs(2403);
    layer2_outputs(6570) <= layer1_outputs(6158);
    layer2_outputs(6571) <= (layer1_outputs(2838)) and not (layer1_outputs(938));
    layer2_outputs(6572) <= layer1_outputs(880);
    layer2_outputs(6573) <= not(layer1_outputs(1847));
    layer2_outputs(6574) <= (layer1_outputs(175)) xor (layer1_outputs(4072));
    layer2_outputs(6575) <= not((layer1_outputs(1577)) or (layer1_outputs(2133)));
    layer2_outputs(6576) <= layer1_outputs(5375);
    layer2_outputs(6577) <= layer1_outputs(4806);
    layer2_outputs(6578) <= layer1_outputs(6150);
    layer2_outputs(6579) <= (layer1_outputs(2779)) and not (layer1_outputs(1875));
    layer2_outputs(6580) <= (layer1_outputs(4905)) and not (layer1_outputs(97));
    layer2_outputs(6581) <= layer1_outputs(314);
    layer2_outputs(6582) <= (layer1_outputs(6076)) and (layer1_outputs(6671));
    layer2_outputs(6583) <= (layer1_outputs(6698)) and not (layer1_outputs(6528));
    layer2_outputs(6584) <= not((layer1_outputs(2294)) and (layer1_outputs(642)));
    layer2_outputs(6585) <= not(layer1_outputs(2795)) or (layer1_outputs(6199));
    layer2_outputs(6586) <= not(layer1_outputs(5646));
    layer2_outputs(6587) <= (layer1_outputs(2966)) and not (layer1_outputs(6947));
    layer2_outputs(6588) <= layer1_outputs(383);
    layer2_outputs(6589) <= not((layer1_outputs(2509)) and (layer1_outputs(7390)));
    layer2_outputs(6590) <= (layer1_outputs(3516)) and not (layer1_outputs(1196));
    layer2_outputs(6591) <= layer1_outputs(6874);
    layer2_outputs(6592) <= layer1_outputs(6626);
    layer2_outputs(6593) <= (layer1_outputs(7015)) and not (layer1_outputs(3362));
    layer2_outputs(6594) <= layer1_outputs(127);
    layer2_outputs(6595) <= not((layer1_outputs(2497)) or (layer1_outputs(712)));
    layer2_outputs(6596) <= (layer1_outputs(1905)) and not (layer1_outputs(2498));
    layer2_outputs(6597) <= (layer1_outputs(2461)) and (layer1_outputs(5994));
    layer2_outputs(6598) <= (layer1_outputs(2747)) or (layer1_outputs(4420));
    layer2_outputs(6599) <= not(layer1_outputs(6136)) or (layer1_outputs(1081));
    layer2_outputs(6600) <= (layer1_outputs(6118)) or (layer1_outputs(3621));
    layer2_outputs(6601) <= (layer1_outputs(1820)) and not (layer1_outputs(788));
    layer2_outputs(6602) <= not(layer1_outputs(7123)) or (layer1_outputs(1159));
    layer2_outputs(6603) <= layer1_outputs(2849);
    layer2_outputs(6604) <= not(layer1_outputs(3454)) or (layer1_outputs(6283));
    layer2_outputs(6605) <= not((layer1_outputs(1199)) and (layer1_outputs(1073)));
    layer2_outputs(6606) <= not(layer1_outputs(3270)) or (layer1_outputs(4898));
    layer2_outputs(6607) <= (layer1_outputs(2149)) and not (layer1_outputs(6357));
    layer2_outputs(6608) <= not(layer1_outputs(6367)) or (layer1_outputs(5836));
    layer2_outputs(6609) <= layer1_outputs(4659);
    layer2_outputs(6610) <= not(layer1_outputs(1406));
    layer2_outputs(6611) <= not((layer1_outputs(5231)) and (layer1_outputs(4002)));
    layer2_outputs(6612) <= not(layer1_outputs(7409));
    layer2_outputs(6613) <= not(layer1_outputs(1773));
    layer2_outputs(6614) <= not(layer1_outputs(1057));
    layer2_outputs(6615) <= not(layer1_outputs(4453)) or (layer1_outputs(73));
    layer2_outputs(6616) <= not((layer1_outputs(6084)) and (layer1_outputs(1969)));
    layer2_outputs(6617) <= (layer1_outputs(2334)) or (layer1_outputs(1000));
    layer2_outputs(6618) <= '1';
    layer2_outputs(6619) <= (layer1_outputs(4792)) and (layer1_outputs(6294));
    layer2_outputs(6620) <= not(layer1_outputs(356));
    layer2_outputs(6621) <= not(layer1_outputs(543)) or (layer1_outputs(3274));
    layer2_outputs(6622) <= (layer1_outputs(4082)) and not (layer1_outputs(1108));
    layer2_outputs(6623) <= not(layer1_outputs(573));
    layer2_outputs(6624) <= layer1_outputs(1666);
    layer2_outputs(6625) <= not(layer1_outputs(1864));
    layer2_outputs(6626) <= layer1_outputs(3929);
    layer2_outputs(6627) <= layer1_outputs(4459);
    layer2_outputs(6628) <= '0';
    layer2_outputs(6629) <= layer1_outputs(7298);
    layer2_outputs(6630) <= not(layer1_outputs(3554));
    layer2_outputs(6631) <= (layer1_outputs(21)) and not (layer1_outputs(2709));
    layer2_outputs(6632) <= layer1_outputs(4978);
    layer2_outputs(6633) <= not(layer1_outputs(979));
    layer2_outputs(6634) <= (layer1_outputs(6566)) or (layer1_outputs(4215));
    layer2_outputs(6635) <= layer1_outputs(3624);
    layer2_outputs(6636) <= not(layer1_outputs(778)) or (layer1_outputs(4637));
    layer2_outputs(6637) <= (layer1_outputs(7309)) and not (layer1_outputs(4936));
    layer2_outputs(6638) <= not((layer1_outputs(444)) and (layer1_outputs(846)));
    layer2_outputs(6639) <= not((layer1_outputs(2789)) or (layer1_outputs(1554)));
    layer2_outputs(6640) <= not((layer1_outputs(4749)) or (layer1_outputs(7602)));
    layer2_outputs(6641) <= not((layer1_outputs(4165)) or (layer1_outputs(471)));
    layer2_outputs(6642) <= not((layer1_outputs(4399)) or (layer1_outputs(4076)));
    layer2_outputs(6643) <= (layer1_outputs(497)) and (layer1_outputs(6620));
    layer2_outputs(6644) <= (layer1_outputs(5761)) and not (layer1_outputs(6909));
    layer2_outputs(6645) <= (layer1_outputs(4652)) and (layer1_outputs(3383));
    layer2_outputs(6646) <= (layer1_outputs(5937)) xor (layer1_outputs(7563));
    layer2_outputs(6647) <= layer1_outputs(4567);
    layer2_outputs(6648) <= layer1_outputs(5431);
    layer2_outputs(6649) <= not((layer1_outputs(2058)) or (layer1_outputs(532)));
    layer2_outputs(6650) <= (layer1_outputs(1117)) xor (layer1_outputs(6471));
    layer2_outputs(6651) <= not(layer1_outputs(5821)) or (layer1_outputs(5094));
    layer2_outputs(6652) <= layer1_outputs(1340);
    layer2_outputs(6653) <= not((layer1_outputs(3524)) or (layer1_outputs(1066)));
    layer2_outputs(6654) <= layer1_outputs(700);
    layer2_outputs(6655) <= not(layer1_outputs(3388)) or (layer1_outputs(612));
    layer2_outputs(6656) <= not((layer1_outputs(6684)) and (layer1_outputs(5899)));
    layer2_outputs(6657) <= (layer1_outputs(7150)) and not (layer1_outputs(5780));
    layer2_outputs(6658) <= not((layer1_outputs(93)) and (layer1_outputs(4800)));
    layer2_outputs(6659) <= layer1_outputs(6616);
    layer2_outputs(6660) <= not((layer1_outputs(3155)) xor (layer1_outputs(4998)));
    layer2_outputs(6661) <= not(layer1_outputs(2621));
    layer2_outputs(6662) <= layer1_outputs(301);
    layer2_outputs(6663) <= (layer1_outputs(437)) and not (layer1_outputs(613));
    layer2_outputs(6664) <= layer1_outputs(1298);
    layer2_outputs(6665) <= (layer1_outputs(982)) and (layer1_outputs(4071));
    layer2_outputs(6666) <= not(layer1_outputs(4708));
    layer2_outputs(6667) <= (layer1_outputs(6780)) and not (layer1_outputs(1105));
    layer2_outputs(6668) <= (layer1_outputs(5963)) and (layer1_outputs(3300));
    layer2_outputs(6669) <= layer1_outputs(1562);
    layer2_outputs(6670) <= layer1_outputs(1543);
    layer2_outputs(6671) <= (layer1_outputs(7481)) and not (layer1_outputs(3365));
    layer2_outputs(6672) <= layer1_outputs(6680);
    layer2_outputs(6673) <= layer1_outputs(6416);
    layer2_outputs(6674) <= not(layer1_outputs(6725));
    layer2_outputs(6675) <= not(layer1_outputs(5773)) or (layer1_outputs(35));
    layer2_outputs(6676) <= not(layer1_outputs(6432)) or (layer1_outputs(4615));
    layer2_outputs(6677) <= not(layer1_outputs(3159));
    layer2_outputs(6678) <= not(layer1_outputs(3850));
    layer2_outputs(6679) <= not(layer1_outputs(3790)) or (layer1_outputs(4493));
    layer2_outputs(6680) <= not(layer1_outputs(4262)) or (layer1_outputs(6504));
    layer2_outputs(6681) <= layer1_outputs(7200);
    layer2_outputs(6682) <= not(layer1_outputs(2765));
    layer2_outputs(6683) <= not(layer1_outputs(1597)) or (layer1_outputs(1283));
    layer2_outputs(6684) <= not(layer1_outputs(6227)) or (layer1_outputs(3209));
    layer2_outputs(6685) <= layer1_outputs(25);
    layer2_outputs(6686) <= (layer1_outputs(2694)) and not (layer1_outputs(1738));
    layer2_outputs(6687) <= (layer1_outputs(7665)) and (layer1_outputs(1445));
    layer2_outputs(6688) <= layer1_outputs(972);
    layer2_outputs(6689) <= not(layer1_outputs(302));
    layer2_outputs(6690) <= layer1_outputs(3247);
    layer2_outputs(6691) <= not(layer1_outputs(4858)) or (layer1_outputs(5320));
    layer2_outputs(6692) <= layer1_outputs(1108);
    layer2_outputs(6693) <= layer1_outputs(5989);
    layer2_outputs(6694) <= (layer1_outputs(5886)) or (layer1_outputs(6350));
    layer2_outputs(6695) <= not(layer1_outputs(2936)) or (layer1_outputs(4454));
    layer2_outputs(6696) <= (layer1_outputs(3672)) and not (layer1_outputs(6659));
    layer2_outputs(6697) <= not(layer1_outputs(2548));
    layer2_outputs(6698) <= layer1_outputs(1386);
    layer2_outputs(6699) <= (layer1_outputs(3605)) and not (layer1_outputs(4539));
    layer2_outputs(6700) <= not(layer1_outputs(2539));
    layer2_outputs(6701) <= layer1_outputs(6099);
    layer2_outputs(6702) <= layer1_outputs(89);
    layer2_outputs(6703) <= '1';
    layer2_outputs(6704) <= layer1_outputs(3811);
    layer2_outputs(6705) <= not((layer1_outputs(2547)) xor (layer1_outputs(3860)));
    layer2_outputs(6706) <= not((layer1_outputs(5009)) and (layer1_outputs(2425)));
    layer2_outputs(6707) <= (layer1_outputs(3244)) or (layer1_outputs(166));
    layer2_outputs(6708) <= (layer1_outputs(624)) and (layer1_outputs(5413));
    layer2_outputs(6709) <= not((layer1_outputs(6284)) and (layer1_outputs(2873)));
    layer2_outputs(6710) <= not(layer1_outputs(7610));
    layer2_outputs(6711) <= layer1_outputs(5354);
    layer2_outputs(6712) <= layer1_outputs(5453);
    layer2_outputs(6713) <= layer1_outputs(2631);
    layer2_outputs(6714) <= (layer1_outputs(4901)) and not (layer1_outputs(4319));
    layer2_outputs(6715) <= not((layer1_outputs(5525)) xor (layer1_outputs(6255)));
    layer2_outputs(6716) <= not(layer1_outputs(1829)) or (layer1_outputs(3527));
    layer2_outputs(6717) <= not(layer1_outputs(957));
    layer2_outputs(6718) <= (layer1_outputs(2044)) and (layer1_outputs(4692));
    layer2_outputs(6719) <= not(layer1_outputs(5885)) or (layer1_outputs(2532));
    layer2_outputs(6720) <= (layer1_outputs(4811)) and (layer1_outputs(6823));
    layer2_outputs(6721) <= not(layer1_outputs(4802));
    layer2_outputs(6722) <= not(layer1_outputs(884));
    layer2_outputs(6723) <= layer1_outputs(548);
    layer2_outputs(6724) <= not(layer1_outputs(1779)) or (layer1_outputs(3424));
    layer2_outputs(6725) <= (layer1_outputs(6258)) and not (layer1_outputs(3543));
    layer2_outputs(6726) <= not(layer1_outputs(2977)) or (layer1_outputs(7421));
    layer2_outputs(6727) <= (layer1_outputs(2139)) or (layer1_outputs(1112));
    layer2_outputs(6728) <= not((layer1_outputs(1847)) or (layer1_outputs(1962)));
    layer2_outputs(6729) <= (layer1_outputs(619)) and not (layer1_outputs(2651));
    layer2_outputs(6730) <= (layer1_outputs(1900)) and not (layer1_outputs(4499));
    layer2_outputs(6731) <= not(layer1_outputs(3363)) or (layer1_outputs(1441));
    layer2_outputs(6732) <= not(layer1_outputs(5771));
    layer2_outputs(6733) <= '0';
    layer2_outputs(6734) <= not(layer1_outputs(2935));
    layer2_outputs(6735) <= '0';
    layer2_outputs(6736) <= layer1_outputs(4472);
    layer2_outputs(6737) <= layer1_outputs(6829);
    layer2_outputs(6738) <= (layer1_outputs(4192)) and (layer1_outputs(1593));
    layer2_outputs(6739) <= (layer1_outputs(6783)) and not (layer1_outputs(1085));
    layer2_outputs(6740) <= (layer1_outputs(5936)) and not (layer1_outputs(270));
    layer2_outputs(6741) <= layer1_outputs(6697);
    layer2_outputs(6742) <= not(layer1_outputs(2169)) or (layer1_outputs(2157));
    layer2_outputs(6743) <= not(layer1_outputs(6700));
    layer2_outputs(6744) <= not(layer1_outputs(7620)) or (layer1_outputs(2141));
    layer2_outputs(6745) <= not(layer1_outputs(7488));
    layer2_outputs(6746) <= (layer1_outputs(3303)) or (layer1_outputs(6314));
    layer2_outputs(6747) <= not((layer1_outputs(6335)) xor (layer1_outputs(3260)));
    layer2_outputs(6748) <= (layer1_outputs(5204)) and not (layer1_outputs(6779));
    layer2_outputs(6749) <= not(layer1_outputs(3009));
    layer2_outputs(6750) <= not((layer1_outputs(7347)) and (layer1_outputs(4218)));
    layer2_outputs(6751) <= not(layer1_outputs(6479));
    layer2_outputs(6752) <= not(layer1_outputs(3728)) or (layer1_outputs(5830));
    layer2_outputs(6753) <= not(layer1_outputs(6642)) or (layer1_outputs(2012));
    layer2_outputs(6754) <= layer1_outputs(4581);
    layer2_outputs(6755) <= not(layer1_outputs(4791));
    layer2_outputs(6756) <= layer1_outputs(2875);
    layer2_outputs(6757) <= '0';
    layer2_outputs(6758) <= not(layer1_outputs(3211));
    layer2_outputs(6759) <= not(layer1_outputs(2781)) or (layer1_outputs(6411));
    layer2_outputs(6760) <= not(layer1_outputs(73));
    layer2_outputs(6761) <= '0';
    layer2_outputs(6762) <= not((layer1_outputs(1487)) xor (layer1_outputs(5941)));
    layer2_outputs(6763) <= layer1_outputs(7205);
    layer2_outputs(6764) <= (layer1_outputs(1179)) and not (layer1_outputs(834));
    layer2_outputs(6765) <= (layer1_outputs(1065)) and not (layer1_outputs(3494));
    layer2_outputs(6766) <= layer1_outputs(3841);
    layer2_outputs(6767) <= not(layer1_outputs(7095));
    layer2_outputs(6768) <= (layer1_outputs(6786)) and not (layer1_outputs(6126));
    layer2_outputs(6769) <= (layer1_outputs(501)) and not (layer1_outputs(3097));
    layer2_outputs(6770) <= not((layer1_outputs(4949)) or (layer1_outputs(6849)));
    layer2_outputs(6771) <= not((layer1_outputs(2401)) or (layer1_outputs(6930)));
    layer2_outputs(6772) <= not((layer1_outputs(6109)) or (layer1_outputs(5663)));
    layer2_outputs(6773) <= '1';
    layer2_outputs(6774) <= not((layer1_outputs(684)) or (layer1_outputs(2712)));
    layer2_outputs(6775) <= not(layer1_outputs(7258));
    layer2_outputs(6776) <= (layer1_outputs(1440)) xor (layer1_outputs(5295));
    layer2_outputs(6777) <= (layer1_outputs(6142)) and not (layer1_outputs(7369));
    layer2_outputs(6778) <= not(layer1_outputs(3908));
    layer2_outputs(6779) <= layer1_outputs(6747);
    layer2_outputs(6780) <= (layer1_outputs(3164)) and (layer1_outputs(1397));
    layer2_outputs(6781) <= not(layer1_outputs(3789)) or (layer1_outputs(7054));
    layer2_outputs(6782) <= (layer1_outputs(1602)) or (layer1_outputs(1008));
    layer2_outputs(6783) <= layer1_outputs(592);
    layer2_outputs(6784) <= (layer1_outputs(4400)) or (layer1_outputs(3494));
    layer2_outputs(6785) <= layer1_outputs(5554);
    layer2_outputs(6786) <= not(layer1_outputs(1858));
    layer2_outputs(6787) <= not(layer1_outputs(7019)) or (layer1_outputs(1252));
    layer2_outputs(6788) <= '1';
    layer2_outputs(6789) <= not(layer1_outputs(5144));
    layer2_outputs(6790) <= (layer1_outputs(3079)) and not (layer1_outputs(41));
    layer2_outputs(6791) <= layer1_outputs(7018);
    layer2_outputs(6792) <= not(layer1_outputs(6802));
    layer2_outputs(6793) <= (layer1_outputs(6973)) and not (layer1_outputs(6956));
    layer2_outputs(6794) <= not(layer1_outputs(7267));
    layer2_outputs(6795) <= not(layer1_outputs(5978)) or (layer1_outputs(4507));
    layer2_outputs(6796) <= '0';
    layer2_outputs(6797) <= (layer1_outputs(2553)) or (layer1_outputs(7578));
    layer2_outputs(6798) <= (layer1_outputs(1858)) and not (layer1_outputs(3172));
    layer2_outputs(6799) <= not(layer1_outputs(2730));
    layer2_outputs(6800) <= '1';
    layer2_outputs(6801) <= (layer1_outputs(4500)) and (layer1_outputs(4299));
    layer2_outputs(6802) <= (layer1_outputs(7521)) and (layer1_outputs(3910));
    layer2_outputs(6803) <= not(layer1_outputs(3286));
    layer2_outputs(6804) <= not(layer1_outputs(2641)) or (layer1_outputs(58));
    layer2_outputs(6805) <= layer1_outputs(4587);
    layer2_outputs(6806) <= not((layer1_outputs(843)) and (layer1_outputs(4563)));
    layer2_outputs(6807) <= not(layer1_outputs(1890));
    layer2_outputs(6808) <= layer1_outputs(3573);
    layer2_outputs(6809) <= not(layer1_outputs(3992));
    layer2_outputs(6810) <= not(layer1_outputs(2737));
    layer2_outputs(6811) <= (layer1_outputs(5362)) and (layer1_outputs(6107));
    layer2_outputs(6812) <= (layer1_outputs(3874)) or (layer1_outputs(1653));
    layer2_outputs(6813) <= layer1_outputs(6739);
    layer2_outputs(6814) <= (layer1_outputs(2455)) or (layer1_outputs(4875));
    layer2_outputs(6815) <= layer1_outputs(2891);
    layer2_outputs(6816) <= '0';
    layer2_outputs(6817) <= '0';
    layer2_outputs(6818) <= not(layer1_outputs(4906));
    layer2_outputs(6819) <= not(layer1_outputs(6475));
    layer2_outputs(6820) <= (layer1_outputs(581)) and not (layer1_outputs(2730));
    layer2_outputs(6821) <= layer1_outputs(2581);
    layer2_outputs(6822) <= not(layer1_outputs(1919)) or (layer1_outputs(4359));
    layer2_outputs(6823) <= (layer1_outputs(1855)) or (layer1_outputs(1869));
    layer2_outputs(6824) <= not((layer1_outputs(1907)) and (layer1_outputs(7469)));
    layer2_outputs(6825) <= (layer1_outputs(3703)) and (layer1_outputs(6820));
    layer2_outputs(6826) <= '0';
    layer2_outputs(6827) <= layer1_outputs(7510);
    layer2_outputs(6828) <= (layer1_outputs(7651)) or (layer1_outputs(2580));
    layer2_outputs(6829) <= layer1_outputs(1723);
    layer2_outputs(6830) <= not(layer1_outputs(4906));
    layer2_outputs(6831) <= layer1_outputs(1848);
    layer2_outputs(6832) <= (layer1_outputs(5805)) and (layer1_outputs(109));
    layer2_outputs(6833) <= (layer1_outputs(4815)) and not (layer1_outputs(1728));
    layer2_outputs(6834) <= not((layer1_outputs(451)) or (layer1_outputs(718)));
    layer2_outputs(6835) <= not(layer1_outputs(2644)) or (layer1_outputs(5482));
    layer2_outputs(6836) <= not(layer1_outputs(6551));
    layer2_outputs(6837) <= layer1_outputs(2051);
    layer2_outputs(6838) <= layer1_outputs(2798);
    layer2_outputs(6839) <= (layer1_outputs(4520)) and not (layer1_outputs(3954));
    layer2_outputs(6840) <= (layer1_outputs(1880)) or (layer1_outputs(4068));
    layer2_outputs(6841) <= (layer1_outputs(4588)) and not (layer1_outputs(7072));
    layer2_outputs(6842) <= (layer1_outputs(5220)) and (layer1_outputs(2785));
    layer2_outputs(6843) <= (layer1_outputs(1062)) and not (layer1_outputs(836));
    layer2_outputs(6844) <= layer1_outputs(6980);
    layer2_outputs(6845) <= layer1_outputs(6265);
    layer2_outputs(6846) <= not(layer1_outputs(4638));
    layer2_outputs(6847) <= not(layer1_outputs(6333));
    layer2_outputs(6848) <= not(layer1_outputs(6310));
    layer2_outputs(6849) <= not(layer1_outputs(1296));
    layer2_outputs(6850) <= (layer1_outputs(223)) and not (layer1_outputs(1493));
    layer2_outputs(6851) <= not(layer1_outputs(4559));
    layer2_outputs(6852) <= (layer1_outputs(1115)) and not (layer1_outputs(2583));
    layer2_outputs(6853) <= (layer1_outputs(5124)) and (layer1_outputs(2383));
    layer2_outputs(6854) <= not(layer1_outputs(1104));
    layer2_outputs(6855) <= (layer1_outputs(1247)) or (layer1_outputs(6979));
    layer2_outputs(6856) <= (layer1_outputs(4016)) xor (layer1_outputs(205));
    layer2_outputs(6857) <= layer1_outputs(5538);
    layer2_outputs(6858) <= not(layer1_outputs(2940)) or (layer1_outputs(4208));
    layer2_outputs(6859) <= layer1_outputs(5571);
    layer2_outputs(6860) <= layer1_outputs(908);
    layer2_outputs(6861) <= layer1_outputs(350);
    layer2_outputs(6862) <= layer1_outputs(2025);
    layer2_outputs(6863) <= not(layer1_outputs(3780)) or (layer1_outputs(5615));
    layer2_outputs(6864) <= (layer1_outputs(4854)) xor (layer1_outputs(2309));
    layer2_outputs(6865) <= not(layer1_outputs(3157));
    layer2_outputs(6866) <= not(layer1_outputs(3306));
    layer2_outputs(6867) <= not(layer1_outputs(5840));
    layer2_outputs(6868) <= not((layer1_outputs(2565)) or (layer1_outputs(7217)));
    layer2_outputs(6869) <= (layer1_outputs(3537)) and not (layer1_outputs(3578));
    layer2_outputs(6870) <= (layer1_outputs(5740)) and not (layer1_outputs(827));
    layer2_outputs(6871) <= (layer1_outputs(2835)) and (layer1_outputs(2496));
    layer2_outputs(6872) <= layer1_outputs(1063);
    layer2_outputs(6873) <= not(layer1_outputs(5291)) or (layer1_outputs(2504));
    layer2_outputs(6874) <= layer1_outputs(1079);
    layer2_outputs(6875) <= layer1_outputs(1346);
    layer2_outputs(6876) <= not(layer1_outputs(5978));
    layer2_outputs(6877) <= not((layer1_outputs(849)) and (layer1_outputs(3861)));
    layer2_outputs(6878) <= layer1_outputs(1371);
    layer2_outputs(6879) <= (layer1_outputs(5586)) or (layer1_outputs(550));
    layer2_outputs(6880) <= layer1_outputs(6848);
    layer2_outputs(6881) <= not(layer1_outputs(561));
    layer2_outputs(6882) <= not(layer1_outputs(4483)) or (layer1_outputs(4457));
    layer2_outputs(6883) <= (layer1_outputs(5383)) xor (layer1_outputs(3549));
    layer2_outputs(6884) <= layer1_outputs(1826);
    layer2_outputs(6885) <= layer1_outputs(6909);
    layer2_outputs(6886) <= (layer1_outputs(4386)) and not (layer1_outputs(1201));
    layer2_outputs(6887) <= not((layer1_outputs(4107)) xor (layer1_outputs(5982)));
    layer2_outputs(6888) <= (layer1_outputs(3239)) or (layer1_outputs(2328));
    layer2_outputs(6889) <= '0';
    layer2_outputs(6890) <= not(layer1_outputs(7129));
    layer2_outputs(6891) <= layer1_outputs(3500);
    layer2_outputs(6892) <= (layer1_outputs(5215)) and not (layer1_outputs(6957));
    layer2_outputs(6893) <= (layer1_outputs(7277)) and not (layer1_outputs(2665));
    layer2_outputs(6894) <= not(layer1_outputs(2536));
    layer2_outputs(6895) <= (layer1_outputs(4136)) or (layer1_outputs(7147));
    layer2_outputs(6896) <= not(layer1_outputs(1219));
    layer2_outputs(6897) <= not(layer1_outputs(5356)) or (layer1_outputs(3406));
    layer2_outputs(6898) <= '0';
    layer2_outputs(6899) <= not(layer1_outputs(75));
    layer2_outputs(6900) <= not((layer1_outputs(2616)) and (layer1_outputs(6392)));
    layer2_outputs(6901) <= not(layer1_outputs(6863));
    layer2_outputs(6902) <= layer1_outputs(7357);
    layer2_outputs(6903) <= not(layer1_outputs(2572)) or (layer1_outputs(6768));
    layer2_outputs(6904) <= not(layer1_outputs(1285));
    layer2_outputs(6905) <= layer1_outputs(692);
    layer2_outputs(6906) <= not(layer1_outputs(4439));
    layer2_outputs(6907) <= '0';
    layer2_outputs(6908) <= not((layer1_outputs(682)) xor (layer1_outputs(1730)));
    layer2_outputs(6909) <= layer1_outputs(4357);
    layer2_outputs(6910) <= not((layer1_outputs(7259)) or (layer1_outputs(1597)));
    layer2_outputs(6911) <= not((layer1_outputs(2104)) and (layer1_outputs(1917)));
    layer2_outputs(6912) <= not(layer1_outputs(4727)) or (layer1_outputs(4250));
    layer2_outputs(6913) <= layer1_outputs(7578);
    layer2_outputs(6914) <= not((layer1_outputs(5548)) or (layer1_outputs(5454)));
    layer2_outputs(6915) <= not((layer1_outputs(7188)) or (layer1_outputs(1170)));
    layer2_outputs(6916) <= not(layer1_outputs(5535)) or (layer1_outputs(4670));
    layer2_outputs(6917) <= (layer1_outputs(633)) or (layer1_outputs(5598));
    layer2_outputs(6918) <= not(layer1_outputs(1960)) or (layer1_outputs(5875));
    layer2_outputs(6919) <= (layer1_outputs(6600)) and (layer1_outputs(6627));
    layer2_outputs(6920) <= not(layer1_outputs(380)) or (layer1_outputs(3469));
    layer2_outputs(6921) <= layer1_outputs(3111);
    layer2_outputs(6922) <= layer1_outputs(2386);
    layer2_outputs(6923) <= (layer1_outputs(6291)) and not (layer1_outputs(2182));
    layer2_outputs(6924) <= not((layer1_outputs(1762)) or (layer1_outputs(1266)));
    layer2_outputs(6925) <= layer1_outputs(2543);
    layer2_outputs(6926) <= (layer1_outputs(5307)) and (layer1_outputs(1618));
    layer2_outputs(6927) <= not((layer1_outputs(5753)) or (layer1_outputs(5318)));
    layer2_outputs(6928) <= (layer1_outputs(6134)) and not (layer1_outputs(1122));
    layer2_outputs(6929) <= (layer1_outputs(189)) and not (layer1_outputs(6785));
    layer2_outputs(6930) <= (layer1_outputs(1452)) or (layer1_outputs(1766));
    layer2_outputs(6931) <= not(layer1_outputs(1475));
    layer2_outputs(6932) <= (layer1_outputs(1038)) and (layer1_outputs(5343));
    layer2_outputs(6933) <= (layer1_outputs(5504)) and not (layer1_outputs(4235));
    layer2_outputs(6934) <= layer1_outputs(6077);
    layer2_outputs(6935) <= layer1_outputs(7365);
    layer2_outputs(6936) <= not(layer1_outputs(1807));
    layer2_outputs(6937) <= '1';
    layer2_outputs(6938) <= (layer1_outputs(3055)) and not (layer1_outputs(2969));
    layer2_outputs(6939) <= not((layer1_outputs(7091)) and (layer1_outputs(4702)));
    layer2_outputs(6940) <= layer1_outputs(3317);
    layer2_outputs(6941) <= not(layer1_outputs(7511));
    layer2_outputs(6942) <= not(layer1_outputs(3655));
    layer2_outputs(6943) <= not((layer1_outputs(2112)) or (layer1_outputs(3735)));
    layer2_outputs(6944) <= not(layer1_outputs(2110));
    layer2_outputs(6945) <= not(layer1_outputs(7583)) or (layer1_outputs(5851));
    layer2_outputs(6946) <= not(layer1_outputs(3388));
    layer2_outputs(6947) <= not(layer1_outputs(2346)) or (layer1_outputs(263));
    layer2_outputs(6948) <= layer1_outputs(3498);
    layer2_outputs(6949) <= not(layer1_outputs(1900));
    layer2_outputs(6950) <= (layer1_outputs(1365)) xor (layer1_outputs(3256));
    layer2_outputs(6951) <= (layer1_outputs(6700)) and (layer1_outputs(2113));
    layer2_outputs(6952) <= '1';
    layer2_outputs(6953) <= (layer1_outputs(2188)) and not (layer1_outputs(4175));
    layer2_outputs(6954) <= not(layer1_outputs(5939));
    layer2_outputs(6955) <= not((layer1_outputs(3813)) xor (layer1_outputs(7247)));
    layer2_outputs(6956) <= (layer1_outputs(6092)) and (layer1_outputs(6721));
    layer2_outputs(6957) <= '1';
    layer2_outputs(6958) <= not((layer1_outputs(4666)) and (layer1_outputs(4995)));
    layer2_outputs(6959) <= (layer1_outputs(6883)) and (layer1_outputs(62));
    layer2_outputs(6960) <= (layer1_outputs(6758)) and (layer1_outputs(6353));
    layer2_outputs(6961) <= not(layer1_outputs(5054));
    layer2_outputs(6962) <= (layer1_outputs(5929)) or (layer1_outputs(6223));
    layer2_outputs(6963) <= not(layer1_outputs(3200));
    layer2_outputs(6964) <= (layer1_outputs(3409)) and (layer1_outputs(4557));
    layer2_outputs(6965) <= layer1_outputs(3687);
    layer2_outputs(6966) <= not(layer1_outputs(6717));
    layer2_outputs(6967) <= '1';
    layer2_outputs(6968) <= not((layer1_outputs(4167)) and (layer1_outputs(3519)));
    layer2_outputs(6969) <= (layer1_outputs(6985)) and (layer1_outputs(1288));
    layer2_outputs(6970) <= layer1_outputs(7237);
    layer2_outputs(6971) <= not(layer1_outputs(2584)) or (layer1_outputs(5955));
    layer2_outputs(6972) <= not(layer1_outputs(1129));
    layer2_outputs(6973) <= not(layer1_outputs(672));
    layer2_outputs(6974) <= not(layer1_outputs(5148));
    layer2_outputs(6975) <= layer1_outputs(3731);
    layer2_outputs(6976) <= not((layer1_outputs(1003)) and (layer1_outputs(5699)));
    layer2_outputs(6977) <= not((layer1_outputs(101)) xor (layer1_outputs(3551)));
    layer2_outputs(6978) <= (layer1_outputs(2896)) and not (layer1_outputs(2253));
    layer2_outputs(6979) <= (layer1_outputs(38)) and not (layer1_outputs(3833));
    layer2_outputs(6980) <= (layer1_outputs(4725)) and (layer1_outputs(2130));
    layer2_outputs(6981) <= (layer1_outputs(5129)) xor (layer1_outputs(4278));
    layer2_outputs(6982) <= '0';
    layer2_outputs(6983) <= (layer1_outputs(3862)) or (layer1_outputs(3973));
    layer2_outputs(6984) <= layer1_outputs(7553);
    layer2_outputs(6985) <= layer1_outputs(74);
    layer2_outputs(6986) <= layer1_outputs(5702);
    layer2_outputs(6987) <= layer1_outputs(3459);
    layer2_outputs(6988) <= layer1_outputs(6885);
    layer2_outputs(6989) <= layer1_outputs(2338);
    layer2_outputs(6990) <= (layer1_outputs(2621)) or (layer1_outputs(3387));
    layer2_outputs(6991) <= layer1_outputs(7181);
    layer2_outputs(6992) <= not(layer1_outputs(1342)) or (layer1_outputs(5862));
    layer2_outputs(6993) <= layer1_outputs(3355);
    layer2_outputs(6994) <= (layer1_outputs(5348)) and (layer1_outputs(2291));
    layer2_outputs(6995) <= not((layer1_outputs(6505)) and (layer1_outputs(2008)));
    layer2_outputs(6996) <= not(layer1_outputs(5778)) or (layer1_outputs(2998));
    layer2_outputs(6997) <= not(layer1_outputs(4346));
    layer2_outputs(6998) <= (layer1_outputs(3939)) or (layer1_outputs(5517));
    layer2_outputs(6999) <= not(layer1_outputs(7341));
    layer2_outputs(7000) <= '1';
    layer2_outputs(7001) <= not(layer1_outputs(6241));
    layer2_outputs(7002) <= not(layer1_outputs(3361));
    layer2_outputs(7003) <= (layer1_outputs(1707)) and (layer1_outputs(3360));
    layer2_outputs(7004) <= '0';
    layer2_outputs(7005) <= not(layer1_outputs(5316));
    layer2_outputs(7006) <= not(layer1_outputs(650));
    layer2_outputs(7007) <= not((layer1_outputs(7440)) and (layer1_outputs(7296)));
    layer2_outputs(7008) <= layer1_outputs(631);
    layer2_outputs(7009) <= layer1_outputs(3228);
    layer2_outputs(7010) <= not(layer1_outputs(2990));
    layer2_outputs(7011) <= layer1_outputs(4424);
    layer2_outputs(7012) <= (layer1_outputs(7660)) xor (layer1_outputs(3264));
    layer2_outputs(7013) <= not(layer1_outputs(3184)) or (layer1_outputs(2090));
    layer2_outputs(7014) <= layer1_outputs(752);
    layer2_outputs(7015) <= '1';
    layer2_outputs(7016) <= layer1_outputs(7316);
    layer2_outputs(7017) <= layer1_outputs(1031);
    layer2_outputs(7018) <= not(layer1_outputs(4877)) or (layer1_outputs(3948));
    layer2_outputs(7019) <= (layer1_outputs(6465)) and not (layer1_outputs(5560));
    layer2_outputs(7020) <= (layer1_outputs(2650)) and not (layer1_outputs(7399));
    layer2_outputs(7021) <= not((layer1_outputs(7588)) or (layer1_outputs(7472)));
    layer2_outputs(7022) <= layer1_outputs(3978);
    layer2_outputs(7023) <= (layer1_outputs(7020)) and not (layer1_outputs(3093));
    layer2_outputs(7024) <= layer1_outputs(2093);
    layer2_outputs(7025) <= not(layer1_outputs(2286));
    layer2_outputs(7026) <= not(layer1_outputs(6775));
    layer2_outputs(7027) <= not(layer1_outputs(1601)) or (layer1_outputs(3576));
    layer2_outputs(7028) <= not(layer1_outputs(2298)) or (layer1_outputs(334));
    layer2_outputs(7029) <= not((layer1_outputs(3872)) or (layer1_outputs(1222)));
    layer2_outputs(7030) <= not(layer1_outputs(6450));
    layer2_outputs(7031) <= not(layer1_outputs(1249));
    layer2_outputs(7032) <= (layer1_outputs(5122)) and (layer1_outputs(6343));
    layer2_outputs(7033) <= '0';
    layer2_outputs(7034) <= layer1_outputs(1142);
    layer2_outputs(7035) <= (layer1_outputs(854)) and (layer1_outputs(160));
    layer2_outputs(7036) <= not(layer1_outputs(977));
    layer2_outputs(7037) <= not(layer1_outputs(1544));
    layer2_outputs(7038) <= layer1_outputs(4982);
    layer2_outputs(7039) <= not((layer1_outputs(5039)) or (layer1_outputs(5979)));
    layer2_outputs(7040) <= not(layer1_outputs(5837));
    layer2_outputs(7041) <= not((layer1_outputs(2360)) and (layer1_outputs(1200)));
    layer2_outputs(7042) <= (layer1_outputs(1188)) and not (layer1_outputs(258));
    layer2_outputs(7043) <= layer1_outputs(190);
    layer2_outputs(7044) <= (layer1_outputs(3807)) and not (layer1_outputs(5428));
    layer2_outputs(7045) <= '1';
    layer2_outputs(7046) <= layer1_outputs(7569);
    layer2_outputs(7047) <= not(layer1_outputs(2455));
    layer2_outputs(7048) <= not(layer1_outputs(6842)) or (layer1_outputs(1123));
    layer2_outputs(7049) <= not(layer1_outputs(1338)) or (layer1_outputs(1208));
    layer2_outputs(7050) <= layer1_outputs(7646);
    layer2_outputs(7051) <= layer1_outputs(5421);
    layer2_outputs(7052) <= not(layer1_outputs(2171));
    layer2_outputs(7053) <= not(layer1_outputs(5341));
    layer2_outputs(7054) <= not(layer1_outputs(375));
    layer2_outputs(7055) <= layer1_outputs(3085);
    layer2_outputs(7056) <= not((layer1_outputs(2931)) or (layer1_outputs(3381)));
    layer2_outputs(7057) <= not(layer1_outputs(1504));
    layer2_outputs(7058) <= layer1_outputs(4447);
    layer2_outputs(7059) <= layer1_outputs(2952);
    layer2_outputs(7060) <= not(layer1_outputs(338));
    layer2_outputs(7061) <= (layer1_outputs(3529)) and (layer1_outputs(6589));
    layer2_outputs(7062) <= layer1_outputs(4930);
    layer2_outputs(7063) <= not(layer1_outputs(4363));
    layer2_outputs(7064) <= (layer1_outputs(7262)) and not (layer1_outputs(7195));
    layer2_outputs(7065) <= layer1_outputs(669);
    layer2_outputs(7066) <= layer1_outputs(5233);
    layer2_outputs(7067) <= not((layer1_outputs(367)) or (layer1_outputs(4413)));
    layer2_outputs(7068) <= not(layer1_outputs(5040));
    layer2_outputs(7069) <= layer1_outputs(4475);
    layer2_outputs(7070) <= not((layer1_outputs(1028)) or (layer1_outputs(5585)));
    layer2_outputs(7071) <= not(layer1_outputs(2825));
    layer2_outputs(7072) <= (layer1_outputs(2663)) and (layer1_outputs(6934));
    layer2_outputs(7073) <= not((layer1_outputs(593)) and (layer1_outputs(4006)));
    layer2_outputs(7074) <= (layer1_outputs(449)) and (layer1_outputs(266));
    layer2_outputs(7075) <= (layer1_outputs(343)) and (layer1_outputs(7636));
    layer2_outputs(7076) <= layer1_outputs(1385);
    layer2_outputs(7077) <= not((layer1_outputs(3900)) and (layer1_outputs(2808)));
    layer2_outputs(7078) <= (layer1_outputs(4607)) and not (layer1_outputs(4598));
    layer2_outputs(7079) <= (layer1_outputs(340)) and not (layer1_outputs(3780));
    layer2_outputs(7080) <= not(layer1_outputs(3787));
    layer2_outputs(7081) <= not(layer1_outputs(7133));
    layer2_outputs(7082) <= not(layer1_outputs(2732));
    layer2_outputs(7083) <= layer1_outputs(7515);
    layer2_outputs(7084) <= (layer1_outputs(6282)) xor (layer1_outputs(3144));
    layer2_outputs(7085) <= layer1_outputs(592);
    layer2_outputs(7086) <= not(layer1_outputs(4509));
    layer2_outputs(7087) <= not(layer1_outputs(6873)) or (layer1_outputs(3873));
    layer2_outputs(7088) <= (layer1_outputs(1676)) and not (layer1_outputs(3450));
    layer2_outputs(7089) <= not(layer1_outputs(3698));
    layer2_outputs(7090) <= not(layer1_outputs(2775));
    layer2_outputs(7091) <= (layer1_outputs(4169)) and not (layer1_outputs(2339));
    layer2_outputs(7092) <= not((layer1_outputs(4909)) or (layer1_outputs(6997)));
    layer2_outputs(7093) <= (layer1_outputs(6433)) and not (layer1_outputs(7268));
    layer2_outputs(7094) <= not((layer1_outputs(2964)) xor (layer1_outputs(3701)));
    layer2_outputs(7095) <= not((layer1_outputs(675)) and (layer1_outputs(3327)));
    layer2_outputs(7096) <= not((layer1_outputs(1915)) or (layer1_outputs(2565)));
    layer2_outputs(7097) <= (layer1_outputs(3952)) xor (layer1_outputs(3834));
    layer2_outputs(7098) <= not(layer1_outputs(249));
    layer2_outputs(7099) <= '1';
    layer2_outputs(7100) <= not((layer1_outputs(5303)) or (layer1_outputs(223)));
    layer2_outputs(7101) <= (layer1_outputs(2492)) or (layer1_outputs(1231));
    layer2_outputs(7102) <= layer1_outputs(5188);
    layer2_outputs(7103) <= not((layer1_outputs(2300)) or (layer1_outputs(6653)));
    layer2_outputs(7104) <= layer1_outputs(7244);
    layer2_outputs(7105) <= '1';
    layer2_outputs(7106) <= not(layer1_outputs(1984)) or (layer1_outputs(6075));
    layer2_outputs(7107) <= not(layer1_outputs(379));
    layer2_outputs(7108) <= not(layer1_outputs(3005));
    layer2_outputs(7109) <= not(layer1_outputs(1480)) or (layer1_outputs(490));
    layer2_outputs(7110) <= not((layer1_outputs(2622)) or (layer1_outputs(491)));
    layer2_outputs(7111) <= not(layer1_outputs(2696));
    layer2_outputs(7112) <= not(layer1_outputs(324));
    layer2_outputs(7113) <= not(layer1_outputs(4586)) or (layer1_outputs(1109));
    layer2_outputs(7114) <= (layer1_outputs(3979)) and (layer1_outputs(5030));
    layer2_outputs(7115) <= layer1_outputs(5173);
    layer2_outputs(7116) <= not(layer1_outputs(155));
    layer2_outputs(7117) <= not(layer1_outputs(4466)) or (layer1_outputs(3569));
    layer2_outputs(7118) <= (layer1_outputs(4883)) and not (layer1_outputs(483));
    layer2_outputs(7119) <= not(layer1_outputs(1615));
    layer2_outputs(7120) <= (layer1_outputs(4711)) and not (layer1_outputs(1553));
    layer2_outputs(7121) <= not(layer1_outputs(4539));
    layer2_outputs(7122) <= (layer1_outputs(1633)) or (layer1_outputs(559));
    layer2_outputs(7123) <= layer1_outputs(3091);
    layer2_outputs(7124) <= layer1_outputs(46);
    layer2_outputs(7125) <= not(layer1_outputs(6735)) or (layer1_outputs(5953));
    layer2_outputs(7126) <= not(layer1_outputs(6245));
    layer2_outputs(7127) <= not(layer1_outputs(6427));
    layer2_outputs(7128) <= not(layer1_outputs(5152)) or (layer1_outputs(4951));
    layer2_outputs(7129) <= '0';
    layer2_outputs(7130) <= not(layer1_outputs(4911)) or (layer1_outputs(1909));
    layer2_outputs(7131) <= not(layer1_outputs(6915));
    layer2_outputs(7132) <= (layer1_outputs(5459)) and not (layer1_outputs(5580));
    layer2_outputs(7133) <= not(layer1_outputs(3896));
    layer2_outputs(7134) <= (layer1_outputs(677)) or (layer1_outputs(7043));
    layer2_outputs(7135) <= not(layer1_outputs(7131));
    layer2_outputs(7136) <= not(layer1_outputs(1149)) or (layer1_outputs(4338));
    layer2_outputs(7137) <= not((layer1_outputs(7281)) xor (layer1_outputs(911)));
    layer2_outputs(7138) <= (layer1_outputs(2314)) and (layer1_outputs(6305));
    layer2_outputs(7139) <= layer1_outputs(4439);
    layer2_outputs(7140) <= layer1_outputs(6393);
    layer2_outputs(7141) <= not(layer1_outputs(142)) or (layer1_outputs(6569));
    layer2_outputs(7142) <= not(layer1_outputs(1273)) or (layer1_outputs(285));
    layer2_outputs(7143) <= (layer1_outputs(2296)) and (layer1_outputs(4969));
    layer2_outputs(7144) <= layer1_outputs(2483);
    layer2_outputs(7145) <= not(layer1_outputs(5818));
    layer2_outputs(7146) <= not(layer1_outputs(4673));
    layer2_outputs(7147) <= (layer1_outputs(2803)) and not (layer1_outputs(5121));
    layer2_outputs(7148) <= layer1_outputs(5254);
    layer2_outputs(7149) <= layer1_outputs(1315);
    layer2_outputs(7150) <= not(layer1_outputs(7255)) or (layer1_outputs(3882));
    layer2_outputs(7151) <= (layer1_outputs(4004)) and not (layer1_outputs(1182));
    layer2_outputs(7152) <= not(layer1_outputs(211)) or (layer1_outputs(5262));
    layer2_outputs(7153) <= not(layer1_outputs(2569));
    layer2_outputs(7154) <= (layer1_outputs(7301)) or (layer1_outputs(3804));
    layer2_outputs(7155) <= '1';
    layer2_outputs(7156) <= not(layer1_outputs(299)) or (layer1_outputs(3242));
    layer2_outputs(7157) <= layer1_outputs(1304);
    layer2_outputs(7158) <= not(layer1_outputs(6185));
    layer2_outputs(7159) <= layer1_outputs(29);
    layer2_outputs(7160) <= layer1_outputs(4171);
    layer2_outputs(7161) <= not((layer1_outputs(4065)) or (layer1_outputs(406)));
    layer2_outputs(7162) <= layer1_outputs(7520);
    layer2_outputs(7163) <= not(layer1_outputs(2930)) or (layer1_outputs(2308));
    layer2_outputs(7164) <= '1';
    layer2_outputs(7165) <= not((layer1_outputs(2570)) or (layer1_outputs(2295)));
    layer2_outputs(7166) <= not((layer1_outputs(5662)) and (layer1_outputs(4315)));
    layer2_outputs(7167) <= (layer1_outputs(1288)) or (layer1_outputs(4698));
    layer2_outputs(7168) <= layer1_outputs(1151);
    layer2_outputs(7169) <= layer1_outputs(3230);
    layer2_outputs(7170) <= not(layer1_outputs(3623));
    layer2_outputs(7171) <= (layer1_outputs(6702)) xor (layer1_outputs(1236));
    layer2_outputs(7172) <= not(layer1_outputs(4536)) or (layer1_outputs(7380));
    layer2_outputs(7173) <= '1';
    layer2_outputs(7174) <= not((layer1_outputs(3198)) xor (layer1_outputs(1383)));
    layer2_outputs(7175) <= not(layer1_outputs(6950));
    layer2_outputs(7176) <= (layer1_outputs(2569)) and (layer1_outputs(5702));
    layer2_outputs(7177) <= '0';
    layer2_outputs(7178) <= (layer1_outputs(1470)) and (layer1_outputs(5624));
    layer2_outputs(7179) <= (layer1_outputs(1795)) and (layer1_outputs(5201));
    layer2_outputs(7180) <= (layer1_outputs(674)) and not (layer1_outputs(2631));
    layer2_outputs(7181) <= not(layer1_outputs(2259)) or (layer1_outputs(2416));
    layer2_outputs(7182) <= not(layer1_outputs(6088)) or (layer1_outputs(1626));
    layer2_outputs(7183) <= '1';
    layer2_outputs(7184) <= not(layer1_outputs(5066));
    layer2_outputs(7185) <= (layer1_outputs(2615)) and not (layer1_outputs(4684));
    layer2_outputs(7186) <= '1';
    layer2_outputs(7187) <= layer1_outputs(121);
    layer2_outputs(7188) <= (layer1_outputs(4299)) and not (layer1_outputs(5718));
    layer2_outputs(7189) <= '0';
    layer2_outputs(7190) <= layer1_outputs(6678);
    layer2_outputs(7191) <= '1';
    layer2_outputs(7192) <= layer1_outputs(4688);
    layer2_outputs(7193) <= '0';
    layer2_outputs(7194) <= (layer1_outputs(3507)) and (layer1_outputs(762));
    layer2_outputs(7195) <= not(layer1_outputs(5230));
    layer2_outputs(7196) <= not(layer1_outputs(4445)) or (layer1_outputs(580));
    layer2_outputs(7197) <= (layer1_outputs(1724)) or (layer1_outputs(6112));
    layer2_outputs(7198) <= (layer1_outputs(4572)) and not (layer1_outputs(4188));
    layer2_outputs(7199) <= (layer1_outputs(4478)) and not (layer1_outputs(3545));
    layer2_outputs(7200) <= layer1_outputs(1127);
    layer2_outputs(7201) <= not(layer1_outputs(7576)) or (layer1_outputs(4935));
    layer2_outputs(7202) <= layer1_outputs(4366);
    layer2_outputs(7203) <= (layer1_outputs(2411)) and (layer1_outputs(736));
    layer2_outputs(7204) <= not(layer1_outputs(5868));
    layer2_outputs(7205) <= (layer1_outputs(4215)) and not (layer1_outputs(3392));
    layer2_outputs(7206) <= not(layer1_outputs(7055));
    layer2_outputs(7207) <= not((layer1_outputs(1135)) or (layer1_outputs(2893)));
    layer2_outputs(7208) <= '1';
    layer2_outputs(7209) <= not(layer1_outputs(5761)) or (layer1_outputs(4206));
    layer2_outputs(7210) <= '1';
    layer2_outputs(7211) <= not(layer1_outputs(2399));
    layer2_outputs(7212) <= not((layer1_outputs(186)) or (layer1_outputs(7078)));
    layer2_outputs(7213) <= not(layer1_outputs(758));
    layer2_outputs(7214) <= (layer1_outputs(7190)) and (layer1_outputs(3650));
    layer2_outputs(7215) <= (layer1_outputs(7341)) or (layer1_outputs(1287));
    layer2_outputs(7216) <= (layer1_outputs(3386)) or (layer1_outputs(7322));
    layer2_outputs(7217) <= layer1_outputs(6183);
    layer2_outputs(7218) <= (layer1_outputs(2909)) and not (layer1_outputs(7639));
    layer2_outputs(7219) <= not(layer1_outputs(1408)) or (layer1_outputs(6546));
    layer2_outputs(7220) <= (layer1_outputs(82)) or (layer1_outputs(7185));
    layer2_outputs(7221) <= layer1_outputs(4302);
    layer2_outputs(7222) <= layer1_outputs(226);
    layer2_outputs(7223) <= not(layer1_outputs(6024));
    layer2_outputs(7224) <= (layer1_outputs(3991)) or (layer1_outputs(2554));
    layer2_outputs(7225) <= not(layer1_outputs(7085));
    layer2_outputs(7226) <= not(layer1_outputs(6983));
    layer2_outputs(7227) <= not(layer1_outputs(6184));
    layer2_outputs(7228) <= not(layer1_outputs(2702));
    layer2_outputs(7229) <= not((layer1_outputs(2750)) xor (layer1_outputs(936)));
    layer2_outputs(7230) <= layer1_outputs(6580);
    layer2_outputs(7231) <= not(layer1_outputs(2500)) or (layer1_outputs(287));
    layer2_outputs(7232) <= layer1_outputs(2787);
    layer2_outputs(7233) <= (layer1_outputs(744)) and (layer1_outputs(220));
    layer2_outputs(7234) <= not(layer1_outputs(4328));
    layer2_outputs(7235) <= layer1_outputs(473);
    layer2_outputs(7236) <= not(layer1_outputs(608));
    layer2_outputs(7237) <= (layer1_outputs(7619)) and not (layer1_outputs(2178));
    layer2_outputs(7238) <= (layer1_outputs(4686)) or (layer1_outputs(6275));
    layer2_outputs(7239) <= not(layer1_outputs(6554));
    layer2_outputs(7240) <= not(layer1_outputs(2967));
    layer2_outputs(7241) <= layer1_outputs(6425);
    layer2_outputs(7242) <= not(layer1_outputs(3749));
    layer2_outputs(7243) <= (layer1_outputs(1426)) and not (layer1_outputs(618));
    layer2_outputs(7244) <= layer1_outputs(629);
    layer2_outputs(7245) <= not(layer1_outputs(221));
    layer2_outputs(7246) <= not(layer1_outputs(5029));
    layer2_outputs(7247) <= not(layer1_outputs(3613));
    layer2_outputs(7248) <= (layer1_outputs(7573)) and (layer1_outputs(2759));
    layer2_outputs(7249) <= (layer1_outputs(3742)) and not (layer1_outputs(5644));
    layer2_outputs(7250) <= not(layer1_outputs(1868)) or (layer1_outputs(1287));
    layer2_outputs(7251) <= (layer1_outputs(6216)) and not (layer1_outputs(3162));
    layer2_outputs(7252) <= not(layer1_outputs(121)) or (layer1_outputs(339));
    layer2_outputs(7253) <= layer1_outputs(4096);
    layer2_outputs(7254) <= (layer1_outputs(1533)) and (layer1_outputs(6517));
    layer2_outputs(7255) <= not(layer1_outputs(6089)) or (layer1_outputs(5767));
    layer2_outputs(7256) <= not((layer1_outputs(777)) or (layer1_outputs(426)));
    layer2_outputs(7257) <= not(layer1_outputs(2528));
    layer2_outputs(7258) <= not(layer1_outputs(5168));
    layer2_outputs(7259) <= layer1_outputs(3195);
    layer2_outputs(7260) <= '0';
    layer2_outputs(7261) <= '1';
    layer2_outputs(7262) <= '0';
    layer2_outputs(7263) <= not(layer1_outputs(2794)) or (layer1_outputs(6197));
    layer2_outputs(7264) <= layer1_outputs(6459);
    layer2_outputs(7265) <= layer1_outputs(1596);
    layer2_outputs(7266) <= not((layer1_outputs(4008)) or (layer1_outputs(1725)));
    layer2_outputs(7267) <= layer1_outputs(4281);
    layer2_outputs(7268) <= '1';
    layer2_outputs(7269) <= not(layer1_outputs(5914)) or (layer1_outputs(2285));
    layer2_outputs(7270) <= '0';
    layer2_outputs(7271) <= (layer1_outputs(6502)) and not (layer1_outputs(5000));
    layer2_outputs(7272) <= (layer1_outputs(7081)) or (layer1_outputs(6298));
    layer2_outputs(7273) <= layer1_outputs(3002);
    layer2_outputs(7274) <= (layer1_outputs(5426)) and (layer1_outputs(5687));
    layer2_outputs(7275) <= not((layer1_outputs(273)) and (layer1_outputs(5025)));
    layer2_outputs(7276) <= layer1_outputs(945);
    layer2_outputs(7277) <= not((layer1_outputs(6523)) and (layer1_outputs(3412)));
    layer2_outputs(7278) <= not((layer1_outputs(292)) xor (layer1_outputs(6509)));
    layer2_outputs(7279) <= not(layer1_outputs(5173)) or (layer1_outputs(1012));
    layer2_outputs(7280) <= layer1_outputs(4014);
    layer2_outputs(7281) <= not(layer1_outputs(1821));
    layer2_outputs(7282) <= not(layer1_outputs(2806));
    layer2_outputs(7283) <= '0';
    layer2_outputs(7284) <= (layer1_outputs(6368)) and not (layer1_outputs(3485));
    layer2_outputs(7285) <= not((layer1_outputs(2109)) or (layer1_outputs(1948)));
    layer2_outputs(7286) <= not(layer1_outputs(7567));
    layer2_outputs(7287) <= (layer1_outputs(748)) or (layer1_outputs(7273));
    layer2_outputs(7288) <= not(layer1_outputs(2612));
    layer2_outputs(7289) <= not(layer1_outputs(5192));
    layer2_outputs(7290) <= not(layer1_outputs(3826)) or (layer1_outputs(4630));
    layer2_outputs(7291) <= (layer1_outputs(1507)) and not (layer1_outputs(3222));
    layer2_outputs(7292) <= layer1_outputs(312);
    layer2_outputs(7293) <= (layer1_outputs(2582)) and (layer1_outputs(1512));
    layer2_outputs(7294) <= layer1_outputs(7120);
    layer2_outputs(7295) <= '1';
    layer2_outputs(7296) <= (layer1_outputs(5655)) and not (layer1_outputs(597));
    layer2_outputs(7297) <= not(layer1_outputs(829));
    layer2_outputs(7298) <= not(layer1_outputs(1794));
    layer2_outputs(7299) <= not(layer1_outputs(5817));
    layer2_outputs(7300) <= not(layer1_outputs(878));
    layer2_outputs(7301) <= not((layer1_outputs(3270)) xor (layer1_outputs(2842)));
    layer2_outputs(7302) <= (layer1_outputs(988)) and not (layer1_outputs(7392));
    layer2_outputs(7303) <= not((layer1_outputs(590)) and (layer1_outputs(4452)));
    layer2_outputs(7304) <= (layer1_outputs(3550)) and not (layer1_outputs(4289));
    layer2_outputs(7305) <= layer1_outputs(7561);
    layer2_outputs(7306) <= (layer1_outputs(4647)) and not (layer1_outputs(7014));
    layer2_outputs(7307) <= not(layer1_outputs(4350));
    layer2_outputs(7308) <= not((layer1_outputs(6753)) or (layer1_outputs(3314)));
    layer2_outputs(7309) <= not(layer1_outputs(3556)) or (layer1_outputs(6809));
    layer2_outputs(7310) <= not(layer1_outputs(7222));
    layer2_outputs(7311) <= layer1_outputs(2287);
    layer2_outputs(7312) <= (layer1_outputs(2766)) and (layer1_outputs(5452));
    layer2_outputs(7313) <= (layer1_outputs(6872)) and (layer1_outputs(3672));
    layer2_outputs(7314) <= (layer1_outputs(5649)) and (layer1_outputs(186));
    layer2_outputs(7315) <= not(layer1_outputs(6262));
    layer2_outputs(7316) <= layer1_outputs(5981);
    layer2_outputs(7317) <= not((layer1_outputs(7554)) or (layer1_outputs(2745)));
    layer2_outputs(7318) <= (layer1_outputs(209)) or (layer1_outputs(3169));
    layer2_outputs(7319) <= not(layer1_outputs(3667)) or (layer1_outputs(1486));
    layer2_outputs(7320) <= (layer1_outputs(5971)) or (layer1_outputs(6185));
    layer2_outputs(7321) <= '1';
    layer2_outputs(7322) <= not(layer1_outputs(4485));
    layer2_outputs(7323) <= not((layer1_outputs(1430)) or (layer1_outputs(5987)));
    layer2_outputs(7324) <= not(layer1_outputs(5422));
    layer2_outputs(7325) <= not((layer1_outputs(1832)) and (layer1_outputs(6867)));
    layer2_outputs(7326) <= layer1_outputs(5952);
    layer2_outputs(7327) <= not(layer1_outputs(87));
    layer2_outputs(7328) <= not(layer1_outputs(2023));
    layer2_outputs(7329) <= not(layer1_outputs(4511));
    layer2_outputs(7330) <= (layer1_outputs(3786)) xor (layer1_outputs(3534));
    layer2_outputs(7331) <= (layer1_outputs(3638)) and not (layer1_outputs(2451));
    layer2_outputs(7332) <= not((layer1_outputs(5135)) and (layer1_outputs(2079)));
    layer2_outputs(7333) <= (layer1_outputs(3744)) and not (layer1_outputs(6669));
    layer2_outputs(7334) <= not(layer1_outputs(5289));
    layer2_outputs(7335) <= not(layer1_outputs(3208));
    layer2_outputs(7336) <= not(layer1_outputs(5652));
    layer2_outputs(7337) <= not(layer1_outputs(3343)) or (layer1_outputs(3946));
    layer2_outputs(7338) <= (layer1_outputs(7233)) or (layer1_outputs(3766));
    layer2_outputs(7339) <= not(layer1_outputs(7361)) or (layer1_outputs(1110));
    layer2_outputs(7340) <= '1';
    layer2_outputs(7341) <= (layer1_outputs(1477)) or (layer1_outputs(5908));
    layer2_outputs(7342) <= (layer1_outputs(3061)) and (layer1_outputs(1931));
    layer2_outputs(7343) <= (layer1_outputs(5470)) and not (layer1_outputs(2302));
    layer2_outputs(7344) <= not(layer1_outputs(5967));
    layer2_outputs(7345) <= not((layer1_outputs(2281)) and (layer1_outputs(3719)));
    layer2_outputs(7346) <= not(layer1_outputs(493));
    layer2_outputs(7347) <= layer1_outputs(311);
    layer2_outputs(7348) <= not(layer1_outputs(2894)) or (layer1_outputs(2674));
    layer2_outputs(7349) <= not((layer1_outputs(2410)) or (layer1_outputs(5420)));
    layer2_outputs(7350) <= (layer1_outputs(2838)) and (layer1_outputs(383));
    layer2_outputs(7351) <= (layer1_outputs(6293)) or (layer1_outputs(1724));
    layer2_outputs(7352) <= not((layer1_outputs(2244)) or (layer1_outputs(4626)));
    layer2_outputs(7353) <= (layer1_outputs(7148)) or (layer1_outputs(1068));
    layer2_outputs(7354) <= layer1_outputs(5757);
    layer2_outputs(7355) <= (layer1_outputs(7209)) and not (layer1_outputs(5810));
    layer2_outputs(7356) <= (layer1_outputs(4597)) and not (layer1_outputs(2994));
    layer2_outputs(7357) <= not(layer1_outputs(4970)) or (layer1_outputs(230));
    layer2_outputs(7358) <= not(layer1_outputs(6365)) or (layer1_outputs(524));
    layer2_outputs(7359) <= '0';
    layer2_outputs(7360) <= '0';
    layer2_outputs(7361) <= not((layer1_outputs(5230)) xor (layer1_outputs(2736)));
    layer2_outputs(7362) <= (layer1_outputs(2815)) and not (layer1_outputs(2703));
    layer2_outputs(7363) <= (layer1_outputs(2181)) and not (layer1_outputs(6736));
    layer2_outputs(7364) <= layer1_outputs(5816);
    layer2_outputs(7365) <= '1';
    layer2_outputs(7366) <= not(layer1_outputs(6792));
    layer2_outputs(7367) <= not(layer1_outputs(6455));
    layer2_outputs(7368) <= (layer1_outputs(4200)) and (layer1_outputs(881));
    layer2_outputs(7369) <= (layer1_outputs(2498)) and not (layer1_outputs(5512));
    layer2_outputs(7370) <= not(layer1_outputs(1137));
    layer2_outputs(7371) <= layer1_outputs(373);
    layer2_outputs(7372) <= layer1_outputs(4713);
    layer2_outputs(7373) <= not((layer1_outputs(162)) and (layer1_outputs(6826)));
    layer2_outputs(7374) <= not((layer1_outputs(3493)) xor (layer1_outputs(3478)));
    layer2_outputs(7375) <= not((layer1_outputs(4446)) or (layer1_outputs(1902)));
    layer2_outputs(7376) <= layer1_outputs(4672);
    layer2_outputs(7377) <= not((layer1_outputs(5505)) and (layer1_outputs(3515)));
    layer2_outputs(7378) <= not(layer1_outputs(3361));
    layer2_outputs(7379) <= (layer1_outputs(4957)) and (layer1_outputs(394));
    layer2_outputs(7380) <= (layer1_outputs(7674)) and not (layer1_outputs(6789));
    layer2_outputs(7381) <= not(layer1_outputs(2187)) or (layer1_outputs(5281));
    layer2_outputs(7382) <= (layer1_outputs(6793)) or (layer1_outputs(3041));
    layer2_outputs(7383) <= not((layer1_outputs(2112)) and (layer1_outputs(5934)));
    layer2_outputs(7384) <= not((layer1_outputs(509)) xor (layer1_outputs(6559)));
    layer2_outputs(7385) <= (layer1_outputs(6901)) and not (layer1_outputs(7643));
    layer2_outputs(7386) <= not((layer1_outputs(3005)) and (layer1_outputs(2833)));
    layer2_outputs(7387) <= (layer1_outputs(1687)) and (layer1_outputs(2815));
    layer2_outputs(7388) <= '1';
    layer2_outputs(7389) <= not(layer1_outputs(3531));
    layer2_outputs(7390) <= not(layer1_outputs(5471));
    layer2_outputs(7391) <= layer1_outputs(1156);
    layer2_outputs(7392) <= (layer1_outputs(4165)) and (layer1_outputs(7198));
    layer2_outputs(7393) <= not(layer1_outputs(3194)) or (layer1_outputs(4521));
    layer2_outputs(7394) <= not((layer1_outputs(1581)) and (layer1_outputs(3868)));
    layer2_outputs(7395) <= '0';
    layer2_outputs(7396) <= not(layer1_outputs(2490));
    layer2_outputs(7397) <= layer1_outputs(4038);
    layer2_outputs(7398) <= (layer1_outputs(6423)) xor (layer1_outputs(884));
    layer2_outputs(7399) <= not(layer1_outputs(504));
    layer2_outputs(7400) <= not(layer1_outputs(6256));
    layer2_outputs(7401) <= not(layer1_outputs(1834));
    layer2_outputs(7402) <= layer1_outputs(4956);
    layer2_outputs(7403) <= (layer1_outputs(628)) and not (layer1_outputs(4402));
    layer2_outputs(7404) <= layer1_outputs(472);
    layer2_outputs(7405) <= not(layer1_outputs(3591));
    layer2_outputs(7406) <= (layer1_outputs(1549)) and (layer1_outputs(4822));
    layer2_outputs(7407) <= not(layer1_outputs(146));
    layer2_outputs(7408) <= '0';
    layer2_outputs(7409) <= not(layer1_outputs(5681));
    layer2_outputs(7410) <= not(layer1_outputs(3323));
    layer2_outputs(7411) <= '0';
    layer2_outputs(7412) <= not(layer1_outputs(4561));
    layer2_outputs(7413) <= layer1_outputs(5393);
    layer2_outputs(7414) <= not(layer1_outputs(6179));
    layer2_outputs(7415) <= not((layer1_outputs(4859)) or (layer1_outputs(3741)));
    layer2_outputs(7416) <= not(layer1_outputs(5719)) or (layer1_outputs(5743));
    layer2_outputs(7417) <= not(layer1_outputs(2183));
    layer2_outputs(7418) <= not(layer1_outputs(1684));
    layer2_outputs(7419) <= (layer1_outputs(1720)) or (layer1_outputs(1732));
    layer2_outputs(7420) <= not(layer1_outputs(3879));
    layer2_outputs(7421) <= (layer1_outputs(4481)) and not (layer1_outputs(7357));
    layer2_outputs(7422) <= (layer1_outputs(6444)) and not (layer1_outputs(92));
    layer2_outputs(7423) <= not(layer1_outputs(3402));
    layer2_outputs(7424) <= '0';
    layer2_outputs(7425) <= layer1_outputs(148);
    layer2_outputs(7426) <= '1';
    layer2_outputs(7427) <= not((layer1_outputs(3562)) xor (layer1_outputs(4119)));
    layer2_outputs(7428) <= layer1_outputs(1551);
    layer2_outputs(7429) <= not(layer1_outputs(3243));
    layer2_outputs(7430) <= layer1_outputs(837);
    layer2_outputs(7431) <= not(layer1_outputs(6025));
    layer2_outputs(7432) <= (layer1_outputs(222)) or (layer1_outputs(3448));
    layer2_outputs(7433) <= (layer1_outputs(1270)) or (layer1_outputs(10));
    layer2_outputs(7434) <= not(layer1_outputs(219)) or (layer1_outputs(2738));
    layer2_outputs(7435) <= not(layer1_outputs(1212));
    layer2_outputs(7436) <= (layer1_outputs(2278)) and (layer1_outputs(5387));
    layer2_outputs(7437) <= layer1_outputs(2290);
    layer2_outputs(7438) <= not((layer1_outputs(4541)) or (layer1_outputs(5052)));
    layer2_outputs(7439) <= not((layer1_outputs(790)) or (layer1_outputs(3006)));
    layer2_outputs(7440) <= not((layer1_outputs(5647)) and (layer1_outputs(2493)));
    layer2_outputs(7441) <= not((layer1_outputs(5465)) or (layer1_outputs(5612)));
    layer2_outputs(7442) <= not(layer1_outputs(3934)) or (layer1_outputs(4443));
    layer2_outputs(7443) <= layer1_outputs(1033);
    layer2_outputs(7444) <= layer1_outputs(3612);
    layer2_outputs(7445) <= not(layer1_outputs(6033));
    layer2_outputs(7446) <= '0';
    layer2_outputs(7447) <= (layer1_outputs(4050)) and (layer1_outputs(6398));
    layer2_outputs(7448) <= not((layer1_outputs(7050)) and (layer1_outputs(400)));
    layer2_outputs(7449) <= not(layer1_outputs(7029)) or (layer1_outputs(5244));
    layer2_outputs(7450) <= layer1_outputs(6412);
    layer2_outputs(7451) <= (layer1_outputs(2468)) or (layer1_outputs(5623));
    layer2_outputs(7452) <= not(layer1_outputs(4159));
    layer2_outputs(7453) <= (layer1_outputs(6728)) and not (layer1_outputs(3955));
    layer2_outputs(7454) <= (layer1_outputs(4655)) and not (layer1_outputs(4690));
    layer2_outputs(7455) <= not(layer1_outputs(7631));
    layer2_outputs(7456) <= not((layer1_outputs(7410)) xor (layer1_outputs(1567)));
    layer2_outputs(7457) <= layer1_outputs(6554);
    layer2_outputs(7458) <= (layer1_outputs(6190)) and (layer1_outputs(134));
    layer2_outputs(7459) <= not((layer1_outputs(5780)) and (layer1_outputs(3324)));
    layer2_outputs(7460) <= not(layer1_outputs(1284));
    layer2_outputs(7461) <= not(layer1_outputs(7571));
    layer2_outputs(7462) <= layer1_outputs(4228);
    layer2_outputs(7463) <= not(layer1_outputs(7091));
    layer2_outputs(7464) <= not(layer1_outputs(7021)) or (layer1_outputs(4337));
    layer2_outputs(7465) <= layer1_outputs(5775);
    layer2_outputs(7466) <= not(layer1_outputs(3490));
    layer2_outputs(7467) <= not(layer1_outputs(6286));
    layer2_outputs(7468) <= layer1_outputs(5049);
    layer2_outputs(7469) <= (layer1_outputs(2535)) and not (layer1_outputs(4947));
    layer2_outputs(7470) <= not((layer1_outputs(482)) and (layer1_outputs(4307)));
    layer2_outputs(7471) <= not((layer1_outputs(369)) or (layer1_outputs(5795)));
    layer2_outputs(7472) <= (layer1_outputs(2092)) and not (layer1_outputs(5540));
    layer2_outputs(7473) <= not(layer1_outputs(6471));
    layer2_outputs(7474) <= (layer1_outputs(1892)) and not (layer1_outputs(5187));
    layer2_outputs(7475) <= layer1_outputs(1928);
    layer2_outputs(7476) <= not(layer1_outputs(3502));
    layer2_outputs(7477) <= layer1_outputs(372);
    layer2_outputs(7478) <= not((layer1_outputs(4851)) and (layer1_outputs(6278)));
    layer2_outputs(7479) <= (layer1_outputs(1)) and (layer1_outputs(5691));
    layer2_outputs(7480) <= layer1_outputs(1427);
    layer2_outputs(7481) <= layer1_outputs(7473);
    layer2_outputs(7482) <= not(layer1_outputs(5009));
    layer2_outputs(7483) <= layer1_outputs(7103);
    layer2_outputs(7484) <= (layer1_outputs(2344)) and not (layer1_outputs(5945));
    layer2_outputs(7485) <= (layer1_outputs(7146)) or (layer1_outputs(3408));
    layer2_outputs(7486) <= not(layer1_outputs(3627));
    layer2_outputs(7487) <= not(layer1_outputs(3313)) or (layer1_outputs(3969));
    layer2_outputs(7488) <= layer1_outputs(103);
    layer2_outputs(7489) <= (layer1_outputs(2377)) or (layer1_outputs(2243));
    layer2_outputs(7490) <= (layer1_outputs(6783)) and (layer1_outputs(7215));
    layer2_outputs(7491) <= layer1_outputs(4245);
    layer2_outputs(7492) <= layer1_outputs(2307);
    layer2_outputs(7493) <= '0';
    layer2_outputs(7494) <= (layer1_outputs(5759)) and (layer1_outputs(3656));
    layer2_outputs(7495) <= (layer1_outputs(7637)) and not (layer1_outputs(3535));
    layer2_outputs(7496) <= layer1_outputs(1032);
    layer2_outputs(7497) <= not((layer1_outputs(4636)) and (layer1_outputs(3048)));
    layer2_outputs(7498) <= (layer1_outputs(6516)) xor (layer1_outputs(7349));
    layer2_outputs(7499) <= not((layer1_outputs(5386)) and (layer1_outputs(5474)));
    layer2_outputs(7500) <= '0';
    layer2_outputs(7501) <= not((layer1_outputs(1105)) and (layer1_outputs(7206)));
    layer2_outputs(7502) <= not(layer1_outputs(6647)) or (layer1_outputs(6053));
    layer2_outputs(7503) <= layer1_outputs(958);
    layer2_outputs(7504) <= not(layer1_outputs(3013));
    layer2_outputs(7505) <= not(layer1_outputs(355)) or (layer1_outputs(7569));
    layer2_outputs(7506) <= '1';
    layer2_outputs(7507) <= not(layer1_outputs(536));
    layer2_outputs(7508) <= (layer1_outputs(3164)) and not (layer1_outputs(2329));
    layer2_outputs(7509) <= (layer1_outputs(2380)) xor (layer1_outputs(6358));
    layer2_outputs(7510) <= '1';
    layer2_outputs(7511) <= not(layer1_outputs(5288));
    layer2_outputs(7512) <= (layer1_outputs(5035)) or (layer1_outputs(2160));
    layer2_outputs(7513) <= not(layer1_outputs(7282));
    layer2_outputs(7514) <= (layer1_outputs(2961)) and not (layer1_outputs(728));
    layer2_outputs(7515) <= layer1_outputs(3690);
    layer2_outputs(7516) <= not(layer1_outputs(4302));
    layer2_outputs(7517) <= not((layer1_outputs(284)) or (layer1_outputs(5700)));
    layer2_outputs(7518) <= not(layer1_outputs(1431));
    layer2_outputs(7519) <= layer1_outputs(6288);
    layer2_outputs(7520) <= (layer1_outputs(5014)) and not (layer1_outputs(7308));
    layer2_outputs(7521) <= (layer1_outputs(3738)) and not (layer1_outputs(6138));
    layer2_outputs(7522) <= not(layer1_outputs(7649)) or (layer1_outputs(7613));
    layer2_outputs(7523) <= layer1_outputs(3515);
    layer2_outputs(7524) <= layer1_outputs(2385);
    layer2_outputs(7525) <= not(layer1_outputs(6765));
    layer2_outputs(7526) <= (layer1_outputs(2841)) and not (layer1_outputs(6106));
    layer2_outputs(7527) <= not(layer1_outputs(3094));
    layer2_outputs(7528) <= layer1_outputs(1043);
    layer2_outputs(7529) <= not(layer1_outputs(6441)) or (layer1_outputs(1542));
    layer2_outputs(7530) <= (layer1_outputs(4589)) and not (layer1_outputs(6239));
    layer2_outputs(7531) <= (layer1_outputs(5758)) and not (layer1_outputs(3814));
    layer2_outputs(7532) <= (layer1_outputs(38)) or (layer1_outputs(4962));
    layer2_outputs(7533) <= not((layer1_outputs(1574)) or (layer1_outputs(4578)));
    layer2_outputs(7534) <= not((layer1_outputs(3160)) xor (layer1_outputs(3680)));
    layer2_outputs(7535) <= layer1_outputs(5803);
    layer2_outputs(7536) <= not(layer1_outputs(6176));
    layer2_outputs(7537) <= not(layer1_outputs(7225));
    layer2_outputs(7538) <= '1';
    layer2_outputs(7539) <= (layer1_outputs(6907)) xor (layer1_outputs(4496));
    layer2_outputs(7540) <= not(layer1_outputs(7413)) or (layer1_outputs(1453));
    layer2_outputs(7541) <= not(layer1_outputs(5793));
    layer2_outputs(7542) <= not(layer1_outputs(3072));
    layer2_outputs(7543) <= (layer1_outputs(3117)) xor (layer1_outputs(6935));
    layer2_outputs(7544) <= (layer1_outputs(7284)) and not (layer1_outputs(3571));
    layer2_outputs(7545) <= (layer1_outputs(3936)) and not (layer1_outputs(3225));
    layer2_outputs(7546) <= (layer1_outputs(261)) and (layer1_outputs(3265));
    layer2_outputs(7547) <= '0';
    layer2_outputs(7548) <= (layer1_outputs(3734)) or (layer1_outputs(5327));
    layer2_outputs(7549) <= not(layer1_outputs(5243));
    layer2_outputs(7550) <= not(layer1_outputs(5352));
    layer2_outputs(7551) <= layer1_outputs(7393);
    layer2_outputs(7552) <= not((layer1_outputs(3010)) or (layer1_outputs(1947)));
    layer2_outputs(7553) <= layer1_outputs(6905);
    layer2_outputs(7554) <= not((layer1_outputs(929)) and (layer1_outputs(6533)));
    layer2_outputs(7555) <= layer1_outputs(1523);
    layer2_outputs(7556) <= not(layer1_outputs(5182));
    layer2_outputs(7557) <= not((layer1_outputs(1624)) xor (layer1_outputs(3865)));
    layer2_outputs(7558) <= (layer1_outputs(838)) and not (layer1_outputs(635));
    layer2_outputs(7559) <= not(layer1_outputs(6083));
    layer2_outputs(7560) <= not(layer1_outputs(1594));
    layer2_outputs(7561) <= (layer1_outputs(4915)) or (layer1_outputs(4640));
    layer2_outputs(7562) <= '1';
    layer2_outputs(7563) <= layer1_outputs(2768);
    layer2_outputs(7564) <= layer1_outputs(6293);
    layer2_outputs(7565) <= (layer1_outputs(274)) and not (layer1_outputs(779));
    layer2_outputs(7566) <= (layer1_outputs(3007)) and (layer1_outputs(4256));
    layer2_outputs(7567) <= not(layer1_outputs(6990)) or (layer1_outputs(1840));
    layer2_outputs(7568) <= not(layer1_outputs(4878)) or (layer1_outputs(4052));
    layer2_outputs(7569) <= layer1_outputs(6825);
    layer2_outputs(7570) <= layer1_outputs(7472);
    layer2_outputs(7571) <= (layer1_outputs(2647)) and (layer1_outputs(829));
    layer2_outputs(7572) <= not(layer1_outputs(5080)) or (layer1_outputs(2080));
    layer2_outputs(7573) <= (layer1_outputs(522)) and not (layer1_outputs(7110));
    layer2_outputs(7574) <= '0';
    layer2_outputs(7575) <= not(layer1_outputs(2633)) or (layer1_outputs(7620));
    layer2_outputs(7576) <= (layer1_outputs(2717)) and not (layer1_outputs(1678));
    layer2_outputs(7577) <= not((layer1_outputs(2700)) and (layer1_outputs(2642)));
    layer2_outputs(7578) <= (layer1_outputs(3024)) and not (layer1_outputs(907));
    layer2_outputs(7579) <= (layer1_outputs(6767)) and not (layer1_outputs(1300));
    layer2_outputs(7580) <= not((layer1_outputs(4466)) or (layer1_outputs(2770)));
    layer2_outputs(7581) <= layer1_outputs(6056);
    layer2_outputs(7582) <= '1';
    layer2_outputs(7583) <= not(layer1_outputs(3229));
    layer2_outputs(7584) <= not(layer1_outputs(1936));
    layer2_outputs(7585) <= not(layer1_outputs(1997));
    layer2_outputs(7586) <= not(layer1_outputs(7020)) or (layer1_outputs(283));
    layer2_outputs(7587) <= not(layer1_outputs(6558));
    layer2_outputs(7588) <= layer1_outputs(976);
    layer2_outputs(7589) <= '1';
    layer2_outputs(7590) <= layer1_outputs(4308);
    layer2_outputs(7591) <= (layer1_outputs(1679)) and (layer1_outputs(2691));
    layer2_outputs(7592) <= (layer1_outputs(3082)) and not (layer1_outputs(1145));
    layer2_outputs(7593) <= (layer1_outputs(4162)) or (layer1_outputs(5707));
    layer2_outputs(7594) <= '0';
    layer2_outputs(7595) <= (layer1_outputs(4277)) and (layer1_outputs(1970));
    layer2_outputs(7596) <= not(layer1_outputs(260));
    layer2_outputs(7597) <= layer1_outputs(2870);
    layer2_outputs(7598) <= (layer1_outputs(2361)) or (layer1_outputs(6329));
    layer2_outputs(7599) <= layer1_outputs(4364);
    layer2_outputs(7600) <= not(layer1_outputs(5491));
    layer2_outputs(7601) <= not((layer1_outputs(297)) or (layer1_outputs(2002)));
    layer2_outputs(7602) <= layer1_outputs(6982);
    layer2_outputs(7603) <= not((layer1_outputs(6041)) and (layer1_outputs(3593)));
    layer2_outputs(7604) <= layer1_outputs(6470);
    layer2_outputs(7605) <= (layer1_outputs(3985)) xor (layer1_outputs(1000));
    layer2_outputs(7606) <= layer1_outputs(2212);
    layer2_outputs(7607) <= not((layer1_outputs(3632)) or (layer1_outputs(6207)));
    layer2_outputs(7608) <= layer1_outputs(3155);
    layer2_outputs(7609) <= (layer1_outputs(6716)) and (layer1_outputs(5366));
    layer2_outputs(7610) <= (layer1_outputs(7359)) or (layer1_outputs(3307));
    layer2_outputs(7611) <= (layer1_outputs(4850)) or (layer1_outputs(1497));
    layer2_outputs(7612) <= not(layer1_outputs(4709));
    layer2_outputs(7613) <= layer1_outputs(615);
    layer2_outputs(7614) <= '0';
    layer2_outputs(7615) <= layer1_outputs(780);
    layer2_outputs(7616) <= not(layer1_outputs(5122)) or (layer1_outputs(7599));
    layer2_outputs(7617) <= not(layer1_outputs(4184));
    layer2_outputs(7618) <= '1';
    layer2_outputs(7619) <= not((layer1_outputs(2447)) or (layer1_outputs(1094)));
    layer2_outputs(7620) <= layer1_outputs(4030);
    layer2_outputs(7621) <= not(layer1_outputs(2481)) or (layer1_outputs(2991));
    layer2_outputs(7622) <= layer1_outputs(4753);
    layer2_outputs(7623) <= not(layer1_outputs(4414));
    layer2_outputs(7624) <= (layer1_outputs(5533)) and not (layer1_outputs(2068));
    layer2_outputs(7625) <= (layer1_outputs(7527)) and not (layer1_outputs(6576));
    layer2_outputs(7626) <= layer1_outputs(1040);
    layer2_outputs(7627) <= (layer1_outputs(759)) and (layer1_outputs(3375));
    layer2_outputs(7628) <= (layer1_outputs(4315)) and not (layer1_outputs(4313));
    layer2_outputs(7629) <= layer1_outputs(5081);
    layer2_outputs(7630) <= layer1_outputs(5125);
    layer2_outputs(7631) <= not((layer1_outputs(741)) or (layer1_outputs(1271)));
    layer2_outputs(7632) <= not((layer1_outputs(3105)) or (layer1_outputs(647)));
    layer2_outputs(7633) <= '1';
    layer2_outputs(7634) <= (layer1_outputs(1524)) and (layer1_outputs(6309));
    layer2_outputs(7635) <= (layer1_outputs(2283)) and not (layer1_outputs(925));
    layer2_outputs(7636) <= not((layer1_outputs(5363)) xor (layer1_outputs(1788)));
    layer2_outputs(7637) <= (layer1_outputs(1878)) or (layer1_outputs(5738));
    layer2_outputs(7638) <= not(layer1_outputs(6650));
    layer2_outputs(7639) <= (layer1_outputs(4546)) xor (layer1_outputs(4116));
    layer2_outputs(7640) <= (layer1_outputs(5036)) and not (layer1_outputs(440));
    layer2_outputs(7641) <= (layer1_outputs(6072)) and not (layer1_outputs(2380));
    layer2_outputs(7642) <= '0';
    layer2_outputs(7643) <= not((layer1_outputs(4399)) or (layer1_outputs(3113)));
    layer2_outputs(7644) <= (layer1_outputs(2575)) and not (layer1_outputs(3991));
    layer2_outputs(7645) <= (layer1_outputs(3095)) and not (layer1_outputs(1412));
    layer2_outputs(7646) <= (layer1_outputs(1991)) and not (layer1_outputs(6418));
    layer2_outputs(7647) <= '1';
    layer2_outputs(7648) <= not(layer1_outputs(3212));
    layer2_outputs(7649) <= '0';
    layer2_outputs(7650) <= not(layer1_outputs(1754));
    layer2_outputs(7651) <= not(layer1_outputs(2316));
    layer2_outputs(7652) <= layer1_outputs(4816);
    layer2_outputs(7653) <= (layer1_outputs(6986)) xor (layer1_outputs(978));
    layer2_outputs(7654) <= (layer1_outputs(1727)) and (layer1_outputs(5031));
    layer2_outputs(7655) <= layer1_outputs(431);
    layer2_outputs(7656) <= not(layer1_outputs(3944));
    layer2_outputs(7657) <= layer1_outputs(6461);
    layer2_outputs(7658) <= not(layer1_outputs(4025)) or (layer1_outputs(1290));
    layer2_outputs(7659) <= (layer1_outputs(2430)) xor (layer1_outputs(3838));
    layer2_outputs(7660) <= layer1_outputs(1364);
    layer2_outputs(7661) <= not((layer1_outputs(6226)) or (layer1_outputs(6833)));
    layer2_outputs(7662) <= (layer1_outputs(4983)) or (layer1_outputs(6081));
    layer2_outputs(7663) <= not((layer1_outputs(2450)) or (layer1_outputs(988)));
    layer2_outputs(7664) <= not(layer1_outputs(4443));
    layer2_outputs(7665) <= not(layer1_outputs(5088));
    layer2_outputs(7666) <= not((layer1_outputs(3400)) and (layer1_outputs(5335)));
    layer2_outputs(7667) <= (layer1_outputs(847)) and not (layer1_outputs(1977));
    layer2_outputs(7668) <= not(layer1_outputs(6910)) or (layer1_outputs(1234));
    layer2_outputs(7669) <= not((layer1_outputs(6069)) or (layer1_outputs(802)));
    layer2_outputs(7670) <= (layer1_outputs(4564)) or (layer1_outputs(5777));
    layer2_outputs(7671) <= (layer1_outputs(2189)) and not (layer1_outputs(6987));
    layer2_outputs(7672) <= (layer1_outputs(4558)) xor (layer1_outputs(4967));
    layer2_outputs(7673) <= (layer1_outputs(1132)) and (layer1_outputs(6280));
    layer2_outputs(7674) <= layer1_outputs(7230);
    layer2_outputs(7675) <= '1';
    layer2_outputs(7676) <= layer1_outputs(1173);
    layer2_outputs(7677) <= (layer1_outputs(6375)) and (layer1_outputs(5973));
    layer2_outputs(7678) <= not(layer1_outputs(5261));
    layer2_outputs(7679) <= layer1_outputs(1380);
    layer3_outputs(0) <= not((layer2_outputs(4240)) and (layer2_outputs(6061)));
    layer3_outputs(1) <= not(layer2_outputs(4510)) or (layer2_outputs(635));
    layer3_outputs(2) <= not(layer2_outputs(7152));
    layer3_outputs(3) <= layer2_outputs(4234);
    layer3_outputs(4) <= (layer2_outputs(7598)) and not (layer2_outputs(3636));
    layer3_outputs(5) <= (layer2_outputs(6281)) and (layer2_outputs(3029));
    layer3_outputs(6) <= layer2_outputs(2570);
    layer3_outputs(7) <= (layer2_outputs(3623)) and not (layer2_outputs(1183));
    layer3_outputs(8) <= not(layer2_outputs(6445));
    layer3_outputs(9) <= not(layer2_outputs(4831));
    layer3_outputs(10) <= not((layer2_outputs(776)) and (layer2_outputs(2870)));
    layer3_outputs(11) <= (layer2_outputs(1826)) and not (layer2_outputs(7275));
    layer3_outputs(12) <= (layer2_outputs(7496)) and not (layer2_outputs(3775));
    layer3_outputs(13) <= '1';
    layer3_outputs(14) <= layer2_outputs(680);
    layer3_outputs(15) <= not(layer2_outputs(6025));
    layer3_outputs(16) <= '0';
    layer3_outputs(17) <= layer2_outputs(908);
    layer3_outputs(18) <= not(layer2_outputs(382));
    layer3_outputs(19) <= not(layer2_outputs(7425));
    layer3_outputs(20) <= (layer2_outputs(3263)) and not (layer2_outputs(6749));
    layer3_outputs(21) <= layer2_outputs(2751);
    layer3_outputs(22) <= layer2_outputs(841);
    layer3_outputs(23) <= not((layer2_outputs(3394)) or (layer2_outputs(233)));
    layer3_outputs(24) <= layer2_outputs(323);
    layer3_outputs(25) <= not(layer2_outputs(28)) or (layer2_outputs(6680));
    layer3_outputs(26) <= not((layer2_outputs(1104)) or (layer2_outputs(7193)));
    layer3_outputs(27) <= not(layer2_outputs(1204));
    layer3_outputs(28) <= layer2_outputs(4264);
    layer3_outputs(29) <= layer2_outputs(6648);
    layer3_outputs(30) <= not(layer2_outputs(5620)) or (layer2_outputs(6950));
    layer3_outputs(31) <= not(layer2_outputs(769));
    layer3_outputs(32) <= not(layer2_outputs(1559));
    layer3_outputs(33) <= layer2_outputs(5378);
    layer3_outputs(34) <= (layer2_outputs(2427)) xor (layer2_outputs(3702));
    layer3_outputs(35) <= not(layer2_outputs(2849));
    layer3_outputs(36) <= not(layer2_outputs(3958));
    layer3_outputs(37) <= layer2_outputs(920);
    layer3_outputs(38) <= (layer2_outputs(7088)) or (layer2_outputs(1847));
    layer3_outputs(39) <= (layer2_outputs(1934)) and not (layer2_outputs(7190));
    layer3_outputs(40) <= not(layer2_outputs(7092));
    layer3_outputs(41) <= not(layer2_outputs(778));
    layer3_outputs(42) <= not(layer2_outputs(3606));
    layer3_outputs(43) <= '1';
    layer3_outputs(44) <= not((layer2_outputs(5280)) or (layer2_outputs(391)));
    layer3_outputs(45) <= layer2_outputs(1567);
    layer3_outputs(46) <= layer2_outputs(7639);
    layer3_outputs(47) <= not(layer2_outputs(5971));
    layer3_outputs(48) <= (layer2_outputs(6438)) and not (layer2_outputs(6746));
    layer3_outputs(49) <= layer2_outputs(3889);
    layer3_outputs(50) <= layer2_outputs(3268);
    layer3_outputs(51) <= not((layer2_outputs(5834)) and (layer2_outputs(3423)));
    layer3_outputs(52) <= layer2_outputs(6575);
    layer3_outputs(53) <= (layer2_outputs(7482)) and (layer2_outputs(2698));
    layer3_outputs(54) <= layer2_outputs(5714);
    layer3_outputs(55) <= not((layer2_outputs(2762)) xor (layer2_outputs(6724)));
    layer3_outputs(56) <= (layer2_outputs(5467)) or (layer2_outputs(5429));
    layer3_outputs(57) <= layer2_outputs(1734);
    layer3_outputs(58) <= not((layer2_outputs(4037)) xor (layer2_outputs(1213)));
    layer3_outputs(59) <= not(layer2_outputs(6055));
    layer3_outputs(60) <= (layer2_outputs(2107)) or (layer2_outputs(453));
    layer3_outputs(61) <= (layer2_outputs(1079)) and not (layer2_outputs(4579));
    layer3_outputs(62) <= layer2_outputs(3244);
    layer3_outputs(63) <= (layer2_outputs(3898)) and (layer2_outputs(549));
    layer3_outputs(64) <= not(layer2_outputs(2818));
    layer3_outputs(65) <= not(layer2_outputs(1825)) or (layer2_outputs(7242));
    layer3_outputs(66) <= not((layer2_outputs(6631)) xor (layer2_outputs(3665)));
    layer3_outputs(67) <= not(layer2_outputs(5107));
    layer3_outputs(68) <= not(layer2_outputs(1557));
    layer3_outputs(69) <= (layer2_outputs(4225)) xor (layer2_outputs(4286));
    layer3_outputs(70) <= not(layer2_outputs(2292));
    layer3_outputs(71) <= (layer2_outputs(561)) and not (layer2_outputs(6980));
    layer3_outputs(72) <= '1';
    layer3_outputs(73) <= (layer2_outputs(799)) and not (layer2_outputs(6841));
    layer3_outputs(74) <= (layer2_outputs(5991)) and (layer2_outputs(3405));
    layer3_outputs(75) <= layer2_outputs(6737);
    layer3_outputs(76) <= layer2_outputs(6051);
    layer3_outputs(77) <= not(layer2_outputs(2948)) or (layer2_outputs(7645));
    layer3_outputs(78) <= (layer2_outputs(7440)) or (layer2_outputs(1470));
    layer3_outputs(79) <= not(layer2_outputs(6340));
    layer3_outputs(80) <= (layer2_outputs(1851)) xor (layer2_outputs(1337));
    layer3_outputs(81) <= not(layer2_outputs(3847)) or (layer2_outputs(2871));
    layer3_outputs(82) <= layer2_outputs(5014);
    layer3_outputs(83) <= not(layer2_outputs(665));
    layer3_outputs(84) <= not(layer2_outputs(5552)) or (layer2_outputs(3278));
    layer3_outputs(85) <= '1';
    layer3_outputs(86) <= not((layer2_outputs(3833)) or (layer2_outputs(5454)));
    layer3_outputs(87) <= not(layer2_outputs(2868));
    layer3_outputs(88) <= not((layer2_outputs(255)) and (layer2_outputs(2277)));
    layer3_outputs(89) <= layer2_outputs(7139);
    layer3_outputs(90) <= '0';
    layer3_outputs(91) <= not(layer2_outputs(5318)) or (layer2_outputs(5276));
    layer3_outputs(92) <= not(layer2_outputs(1013)) or (layer2_outputs(943));
    layer3_outputs(93) <= layer2_outputs(58);
    layer3_outputs(94) <= layer2_outputs(6705);
    layer3_outputs(95) <= (layer2_outputs(5742)) or (layer2_outputs(6509));
    layer3_outputs(96) <= (layer2_outputs(815)) or (layer2_outputs(9));
    layer3_outputs(97) <= not(layer2_outputs(2809));
    layer3_outputs(98) <= not((layer2_outputs(2437)) and (layer2_outputs(6563)));
    layer3_outputs(99) <= (layer2_outputs(5557)) and (layer2_outputs(3750));
    layer3_outputs(100) <= not(layer2_outputs(5309));
    layer3_outputs(101) <= layer2_outputs(2435);
    layer3_outputs(102) <= layer2_outputs(3288);
    layer3_outputs(103) <= (layer2_outputs(991)) and not (layer2_outputs(5174));
    layer3_outputs(104) <= layer2_outputs(6032);
    layer3_outputs(105) <= (layer2_outputs(6853)) and not (layer2_outputs(5413));
    layer3_outputs(106) <= not(layer2_outputs(2362));
    layer3_outputs(107) <= not(layer2_outputs(1382)) or (layer2_outputs(1533));
    layer3_outputs(108) <= layer2_outputs(7341);
    layer3_outputs(109) <= layer2_outputs(5763);
    layer3_outputs(110) <= '1';
    layer3_outputs(111) <= not((layer2_outputs(777)) or (layer2_outputs(2970)));
    layer3_outputs(112) <= (layer2_outputs(1217)) xor (layer2_outputs(3544));
    layer3_outputs(113) <= layer2_outputs(1208);
    layer3_outputs(114) <= not(layer2_outputs(4458));
    layer3_outputs(115) <= layer2_outputs(5624);
    layer3_outputs(116) <= not(layer2_outputs(5362));
    layer3_outputs(117) <= not(layer2_outputs(734));
    layer3_outputs(118) <= (layer2_outputs(6284)) and not (layer2_outputs(5566));
    layer3_outputs(119) <= not(layer2_outputs(2506)) or (layer2_outputs(7672));
    layer3_outputs(120) <= not(layer2_outputs(1828)) or (layer2_outputs(4610));
    layer3_outputs(121) <= layer2_outputs(6710);
    layer3_outputs(122) <= layer2_outputs(4925);
    layer3_outputs(123) <= layer2_outputs(1396);
    layer3_outputs(124) <= layer2_outputs(4403);
    layer3_outputs(125) <= layer2_outputs(6666);
    layer3_outputs(126) <= (layer2_outputs(6821)) and not (layer2_outputs(1992));
    layer3_outputs(127) <= (layer2_outputs(2258)) xor (layer2_outputs(3474));
    layer3_outputs(128) <= not(layer2_outputs(333)) or (layer2_outputs(2889));
    layer3_outputs(129) <= not(layer2_outputs(2344)) or (layer2_outputs(4336));
    layer3_outputs(130) <= (layer2_outputs(425)) and not (layer2_outputs(4018));
    layer3_outputs(131) <= not(layer2_outputs(2408));
    layer3_outputs(132) <= (layer2_outputs(3759)) and not (layer2_outputs(4030));
    layer3_outputs(133) <= layer2_outputs(4521);
    layer3_outputs(134) <= not(layer2_outputs(1988)) or (layer2_outputs(5484));
    layer3_outputs(135) <= not(layer2_outputs(2588));
    layer3_outputs(136) <= layer2_outputs(6661);
    layer3_outputs(137) <= not(layer2_outputs(7357)) or (layer2_outputs(2247));
    layer3_outputs(138) <= layer2_outputs(6048);
    layer3_outputs(139) <= layer2_outputs(3708);
    layer3_outputs(140) <= not((layer2_outputs(638)) or (layer2_outputs(3356)));
    layer3_outputs(141) <= not(layer2_outputs(3337)) or (layer2_outputs(6597));
    layer3_outputs(142) <= not(layer2_outputs(3871)) or (layer2_outputs(7624));
    layer3_outputs(143) <= not((layer2_outputs(1743)) and (layer2_outputs(5159)));
    layer3_outputs(144) <= not((layer2_outputs(7051)) or (layer2_outputs(7665)));
    layer3_outputs(145) <= layer2_outputs(5058);
    layer3_outputs(146) <= not(layer2_outputs(4199));
    layer3_outputs(147) <= not(layer2_outputs(4015)) or (layer2_outputs(693));
    layer3_outputs(148) <= layer2_outputs(3403);
    layer3_outputs(149) <= '1';
    layer3_outputs(150) <= (layer2_outputs(7609)) xor (layer2_outputs(7418));
    layer3_outputs(151) <= not(layer2_outputs(1901));
    layer3_outputs(152) <= (layer2_outputs(5302)) and not (layer2_outputs(769));
    layer3_outputs(153) <= layer2_outputs(5172);
    layer3_outputs(154) <= (layer2_outputs(3760)) and not (layer2_outputs(3605));
    layer3_outputs(155) <= layer2_outputs(2231);
    layer3_outputs(156) <= not(layer2_outputs(3293)) or (layer2_outputs(5412));
    layer3_outputs(157) <= (layer2_outputs(5451)) and (layer2_outputs(813));
    layer3_outputs(158) <= layer2_outputs(4784);
    layer3_outputs(159) <= not((layer2_outputs(5101)) or (layer2_outputs(2738)));
    layer3_outputs(160) <= (layer2_outputs(5727)) or (layer2_outputs(5142));
    layer3_outputs(161) <= not(layer2_outputs(4673));
    layer3_outputs(162) <= not((layer2_outputs(4032)) or (layer2_outputs(7658)));
    layer3_outputs(163) <= not((layer2_outputs(7053)) xor (layer2_outputs(546)));
    layer3_outputs(164) <= (layer2_outputs(6934)) or (layer2_outputs(4920));
    layer3_outputs(165) <= not((layer2_outputs(220)) xor (layer2_outputs(55)));
    layer3_outputs(166) <= (layer2_outputs(123)) and not (layer2_outputs(1548));
    layer3_outputs(167) <= '1';
    layer3_outputs(168) <= not(layer2_outputs(2756)) or (layer2_outputs(5226));
    layer3_outputs(169) <= (layer2_outputs(4172)) and (layer2_outputs(5282));
    layer3_outputs(170) <= layer2_outputs(2008);
    layer3_outputs(171) <= not(layer2_outputs(308));
    layer3_outputs(172) <= not(layer2_outputs(6095)) or (layer2_outputs(6487));
    layer3_outputs(173) <= layer2_outputs(5769);
    layer3_outputs(174) <= not(layer2_outputs(3476));
    layer3_outputs(175) <= layer2_outputs(5577);
    layer3_outputs(176) <= not((layer2_outputs(5833)) and (layer2_outputs(2371)));
    layer3_outputs(177) <= not(layer2_outputs(1024));
    layer3_outputs(178) <= not(layer2_outputs(7567)) or (layer2_outputs(5676));
    layer3_outputs(179) <= not(layer2_outputs(7361));
    layer3_outputs(180) <= not(layer2_outputs(3642));
    layer3_outputs(181) <= (layer2_outputs(3237)) and not (layer2_outputs(6287));
    layer3_outputs(182) <= not((layer2_outputs(5151)) and (layer2_outputs(5914)));
    layer3_outputs(183) <= layer2_outputs(648);
    layer3_outputs(184) <= (layer2_outputs(3895)) and (layer2_outputs(3373));
    layer3_outputs(185) <= layer2_outputs(3169);
    layer3_outputs(186) <= (layer2_outputs(2299)) or (layer2_outputs(6419));
    layer3_outputs(187) <= not((layer2_outputs(4754)) or (layer2_outputs(5476)));
    layer3_outputs(188) <= layer2_outputs(1547);
    layer3_outputs(189) <= (layer2_outputs(34)) and (layer2_outputs(5662));
    layer3_outputs(190) <= not(layer2_outputs(1148));
    layer3_outputs(191) <= not(layer2_outputs(4492));
    layer3_outputs(192) <= layer2_outputs(6560);
    layer3_outputs(193) <= not(layer2_outputs(5977));
    layer3_outputs(194) <= layer2_outputs(3924);
    layer3_outputs(195) <= '0';
    layer3_outputs(196) <= not(layer2_outputs(3805));
    layer3_outputs(197) <= (layer2_outputs(3680)) xor (layer2_outputs(2263));
    layer3_outputs(198) <= layer2_outputs(6017);
    layer3_outputs(199) <= (layer2_outputs(1618)) xor (layer2_outputs(872));
    layer3_outputs(200) <= not(layer2_outputs(7119));
    layer3_outputs(201) <= layer2_outputs(512);
    layer3_outputs(202) <= not(layer2_outputs(3565));
    layer3_outputs(203) <= (layer2_outputs(7152)) or (layer2_outputs(1870));
    layer3_outputs(204) <= not(layer2_outputs(4757)) or (layer2_outputs(7230));
    layer3_outputs(205) <= (layer2_outputs(4814)) or (layer2_outputs(1599));
    layer3_outputs(206) <= not(layer2_outputs(3027));
    layer3_outputs(207) <= layer2_outputs(7571);
    layer3_outputs(208) <= not((layer2_outputs(6779)) xor (layer2_outputs(1949)));
    layer3_outputs(209) <= not((layer2_outputs(4891)) and (layer2_outputs(1957)));
    layer3_outputs(210) <= layer2_outputs(1606);
    layer3_outputs(211) <= (layer2_outputs(4944)) or (layer2_outputs(322));
    layer3_outputs(212) <= layer2_outputs(2397);
    layer3_outputs(213) <= not((layer2_outputs(421)) and (layer2_outputs(3482)));
    layer3_outputs(214) <= not(layer2_outputs(3340));
    layer3_outputs(215) <= not(layer2_outputs(1690));
    layer3_outputs(216) <= not(layer2_outputs(6716)) or (layer2_outputs(2958));
    layer3_outputs(217) <= layer2_outputs(3889);
    layer3_outputs(218) <= layer2_outputs(2753);
    layer3_outputs(219) <= not(layer2_outputs(3673));
    layer3_outputs(220) <= layer2_outputs(1070);
    layer3_outputs(221) <= layer2_outputs(346);
    layer3_outputs(222) <= layer2_outputs(7412);
    layer3_outputs(223) <= not(layer2_outputs(5131));
    layer3_outputs(224) <= (layer2_outputs(6205)) xor (layer2_outputs(3977));
    layer3_outputs(225) <= not(layer2_outputs(5183));
    layer3_outputs(226) <= not(layer2_outputs(4380));
    layer3_outputs(227) <= not(layer2_outputs(588)) or (layer2_outputs(4059));
    layer3_outputs(228) <= not(layer2_outputs(3242)) or (layer2_outputs(330));
    layer3_outputs(229) <= (layer2_outputs(5181)) and (layer2_outputs(353));
    layer3_outputs(230) <= layer2_outputs(4995);
    layer3_outputs(231) <= '1';
    layer3_outputs(232) <= not(layer2_outputs(7453));
    layer3_outputs(233) <= not((layer2_outputs(6809)) and (layer2_outputs(3190)));
    layer3_outputs(234) <= not((layer2_outputs(558)) xor (layer2_outputs(2700)));
    layer3_outputs(235) <= not(layer2_outputs(7462));
    layer3_outputs(236) <= (layer2_outputs(4425)) xor (layer2_outputs(4961));
    layer3_outputs(237) <= (layer2_outputs(5686)) and not (layer2_outputs(7562));
    layer3_outputs(238) <= layer2_outputs(6522);
    layer3_outputs(239) <= not(layer2_outputs(7651));
    layer3_outputs(240) <= (layer2_outputs(3806)) xor (layer2_outputs(4409));
    layer3_outputs(241) <= not((layer2_outputs(5914)) or (layer2_outputs(2959)));
    layer3_outputs(242) <= not(layer2_outputs(4235));
    layer3_outputs(243) <= not(layer2_outputs(3939));
    layer3_outputs(244) <= not((layer2_outputs(1882)) or (layer2_outputs(6820)));
    layer3_outputs(245) <= '0';
    layer3_outputs(246) <= not(layer2_outputs(4583));
    layer3_outputs(247) <= (layer2_outputs(6263)) xor (layer2_outputs(1029));
    layer3_outputs(248) <= not((layer2_outputs(1504)) and (layer2_outputs(2161)));
    layer3_outputs(249) <= '1';
    layer3_outputs(250) <= (layer2_outputs(1181)) and not (layer2_outputs(5431));
    layer3_outputs(251) <= layer2_outputs(5553);
    layer3_outputs(252) <= not(layer2_outputs(433)) or (layer2_outputs(5145));
    layer3_outputs(253) <= '1';
    layer3_outputs(254) <= layer2_outputs(5024);
    layer3_outputs(255) <= not((layer2_outputs(4635)) and (layer2_outputs(7354)));
    layer3_outputs(256) <= not(layer2_outputs(6991));
    layer3_outputs(257) <= not(layer2_outputs(3547));
    layer3_outputs(258) <= (layer2_outputs(3701)) or (layer2_outputs(5414));
    layer3_outputs(259) <= (layer2_outputs(2372)) and not (layer2_outputs(5777));
    layer3_outputs(260) <= layer2_outputs(2422);
    layer3_outputs(261) <= not(layer2_outputs(4848));
    layer3_outputs(262) <= (layer2_outputs(1491)) and not (layer2_outputs(7354));
    layer3_outputs(263) <= not(layer2_outputs(2654)) or (layer2_outputs(5849));
    layer3_outputs(264) <= layer2_outputs(2652);
    layer3_outputs(265) <= layer2_outputs(5012);
    layer3_outputs(266) <= not(layer2_outputs(3531));
    layer3_outputs(267) <= not(layer2_outputs(521));
    layer3_outputs(268) <= not((layer2_outputs(1888)) or (layer2_outputs(3477)));
    layer3_outputs(269) <= (layer2_outputs(4144)) or (layer2_outputs(4107));
    layer3_outputs(270) <= not((layer2_outputs(5785)) or (layer2_outputs(3769)));
    layer3_outputs(271) <= (layer2_outputs(176)) xor (layer2_outputs(5123));
    layer3_outputs(272) <= layer2_outputs(1011);
    layer3_outputs(273) <= not(layer2_outputs(4775)) or (layer2_outputs(3911));
    layer3_outputs(274) <= (layer2_outputs(3375)) and (layer2_outputs(5243));
    layer3_outputs(275) <= not(layer2_outputs(3511));
    layer3_outputs(276) <= not(layer2_outputs(4967));
    layer3_outputs(277) <= not(layer2_outputs(19));
    layer3_outputs(278) <= (layer2_outputs(1821)) and (layer2_outputs(5389));
    layer3_outputs(279) <= (layer2_outputs(2159)) or (layer2_outputs(7484));
    layer3_outputs(280) <= layer2_outputs(862);
    layer3_outputs(281) <= layer2_outputs(1908);
    layer3_outputs(282) <= not((layer2_outputs(1654)) or (layer2_outputs(2719)));
    layer3_outputs(283) <= not(layer2_outputs(3812));
    layer3_outputs(284) <= not((layer2_outputs(7235)) or (layer2_outputs(3508)));
    layer3_outputs(285) <= not(layer2_outputs(5449));
    layer3_outputs(286) <= layer2_outputs(7185);
    layer3_outputs(287) <= not(layer2_outputs(3318));
    layer3_outputs(288) <= (layer2_outputs(210)) and (layer2_outputs(1449));
    layer3_outputs(289) <= '0';
    layer3_outputs(290) <= (layer2_outputs(4394)) and not (layer2_outputs(7127));
    layer3_outputs(291) <= not(layer2_outputs(5720));
    layer3_outputs(292) <= layer2_outputs(6797);
    layer3_outputs(293) <= not((layer2_outputs(7468)) and (layer2_outputs(1570)));
    layer3_outputs(294) <= layer2_outputs(3332);
    layer3_outputs(295) <= (layer2_outputs(7273)) and not (layer2_outputs(3486));
    layer3_outputs(296) <= not(layer2_outputs(7080)) or (layer2_outputs(1632));
    layer3_outputs(297) <= not(layer2_outputs(3664));
    layer3_outputs(298) <= layer2_outputs(4719);
    layer3_outputs(299) <= (layer2_outputs(947)) and not (layer2_outputs(3221));
    layer3_outputs(300) <= layer2_outputs(1913);
    layer3_outputs(301) <= not(layer2_outputs(4848));
    layer3_outputs(302) <= not(layer2_outputs(2601)) or (layer2_outputs(335));
    layer3_outputs(303) <= not((layer2_outputs(2425)) xor (layer2_outputs(4166)));
    layer3_outputs(304) <= not(layer2_outputs(6952));
    layer3_outputs(305) <= layer2_outputs(271);
    layer3_outputs(306) <= (layer2_outputs(4021)) or (layer2_outputs(241));
    layer3_outputs(307) <= not((layer2_outputs(486)) or (layer2_outputs(7166)));
    layer3_outputs(308) <= not(layer2_outputs(6834));
    layer3_outputs(309) <= (layer2_outputs(2079)) xor (layer2_outputs(2677));
    layer3_outputs(310) <= not(layer2_outputs(298));
    layer3_outputs(311) <= layer2_outputs(6319);
    layer3_outputs(312) <= not(layer2_outputs(2671)) or (layer2_outputs(6540));
    layer3_outputs(313) <= not((layer2_outputs(5299)) or (layer2_outputs(2727)));
    layer3_outputs(314) <= (layer2_outputs(4460)) and not (layer2_outputs(7128));
    layer3_outputs(315) <= layer2_outputs(1958);
    layer3_outputs(316) <= not(layer2_outputs(2071));
    layer3_outputs(317) <= (layer2_outputs(5612)) and not (layer2_outputs(3821));
    layer3_outputs(318) <= not(layer2_outputs(2972));
    layer3_outputs(319) <= layer2_outputs(30);
    layer3_outputs(320) <= layer2_outputs(6778);
    layer3_outputs(321) <= not(layer2_outputs(766));
    layer3_outputs(322) <= not(layer2_outputs(2327)) or (layer2_outputs(1919));
    layer3_outputs(323) <= '1';
    layer3_outputs(324) <= layer2_outputs(2587);
    layer3_outputs(325) <= not(layer2_outputs(3355));
    layer3_outputs(326) <= (layer2_outputs(4254)) and (layer2_outputs(374));
    layer3_outputs(327) <= not(layer2_outputs(6001));
    layer3_outputs(328) <= layer2_outputs(5422);
    layer3_outputs(329) <= (layer2_outputs(1858)) or (layer2_outputs(762));
    layer3_outputs(330) <= not((layer2_outputs(1772)) and (layer2_outputs(6174)));
    layer3_outputs(331) <= '0';
    layer3_outputs(332) <= not((layer2_outputs(2034)) or (layer2_outputs(3839)));
    layer3_outputs(333) <= not(layer2_outputs(7353));
    layer3_outputs(334) <= '0';
    layer3_outputs(335) <= not(layer2_outputs(1366));
    layer3_outputs(336) <= layer2_outputs(6260);
    layer3_outputs(337) <= (layer2_outputs(2802)) and not (layer2_outputs(2846));
    layer3_outputs(338) <= not(layer2_outputs(2573));
    layer3_outputs(339) <= layer2_outputs(1121);
    layer3_outputs(340) <= layer2_outputs(4630);
    layer3_outputs(341) <= layer2_outputs(445);
    layer3_outputs(342) <= layer2_outputs(1076);
    layer3_outputs(343) <= not(layer2_outputs(571));
    layer3_outputs(344) <= not(layer2_outputs(3857)) or (layer2_outputs(582));
    layer3_outputs(345) <= not(layer2_outputs(4704));
    layer3_outputs(346) <= not(layer2_outputs(7544));
    layer3_outputs(347) <= '1';
    layer3_outputs(348) <= not(layer2_outputs(3121));
    layer3_outputs(349) <= layer2_outputs(358);
    layer3_outputs(350) <= (layer2_outputs(3678)) xor (layer2_outputs(6338));
    layer3_outputs(351) <= layer2_outputs(1935);
    layer3_outputs(352) <= not(layer2_outputs(4945));
    layer3_outputs(353) <= (layer2_outputs(6377)) and not (layer2_outputs(6852));
    layer3_outputs(354) <= not((layer2_outputs(1550)) and (layer2_outputs(4450)));
    layer3_outputs(355) <= (layer2_outputs(4326)) and not (layer2_outputs(6542));
    layer3_outputs(356) <= '0';
    layer3_outputs(357) <= not((layer2_outputs(5325)) and (layer2_outputs(2379)));
    layer3_outputs(358) <= not(layer2_outputs(7337)) or (layer2_outputs(6458));
    layer3_outputs(359) <= not((layer2_outputs(3601)) or (layer2_outputs(6777)));
    layer3_outputs(360) <= layer2_outputs(2375);
    layer3_outputs(361) <= '0';
    layer3_outputs(362) <= not(layer2_outputs(5898));
    layer3_outputs(363) <= not((layer2_outputs(5861)) xor (layer2_outputs(3729)));
    layer3_outputs(364) <= '0';
    layer3_outputs(365) <= (layer2_outputs(1703)) or (layer2_outputs(3792));
    layer3_outputs(366) <= not(layer2_outputs(5864));
    layer3_outputs(367) <= not(layer2_outputs(1639));
    layer3_outputs(368) <= not((layer2_outputs(4665)) and (layer2_outputs(1211)));
    layer3_outputs(369) <= (layer2_outputs(1797)) and (layer2_outputs(455));
    layer3_outputs(370) <= not((layer2_outputs(7130)) and (layer2_outputs(314)));
    layer3_outputs(371) <= not((layer2_outputs(2415)) or (layer2_outputs(1649)));
    layer3_outputs(372) <= not(layer2_outputs(4282));
    layer3_outputs(373) <= not((layer2_outputs(5266)) xor (layer2_outputs(7055)));
    layer3_outputs(374) <= not(layer2_outputs(807)) or (layer2_outputs(6569));
    layer3_outputs(375) <= not(layer2_outputs(2978)) or (layer2_outputs(4692));
    layer3_outputs(376) <= layer2_outputs(1780);
    layer3_outputs(377) <= not(layer2_outputs(1180)) or (layer2_outputs(1232));
    layer3_outputs(378) <= not((layer2_outputs(5285)) and (layer2_outputs(4053)));
    layer3_outputs(379) <= not(layer2_outputs(2215));
    layer3_outputs(380) <= layer2_outputs(3364);
    layer3_outputs(381) <= not((layer2_outputs(6885)) or (layer2_outputs(1439)));
    layer3_outputs(382) <= not(layer2_outputs(5016));
    layer3_outputs(383) <= not(layer2_outputs(4475)) or (layer2_outputs(5849));
    layer3_outputs(384) <= (layer2_outputs(3203)) xor (layer2_outputs(763));
    layer3_outputs(385) <= not(layer2_outputs(2594));
    layer3_outputs(386) <= layer2_outputs(6331);
    layer3_outputs(387) <= not(layer2_outputs(3519));
    layer3_outputs(388) <= not((layer2_outputs(7128)) xor (layer2_outputs(5225)));
    layer3_outputs(389) <= not(layer2_outputs(1008)) or (layer2_outputs(5647));
    layer3_outputs(390) <= not((layer2_outputs(796)) xor (layer2_outputs(20)));
    layer3_outputs(391) <= layer2_outputs(3716);
    layer3_outputs(392) <= (layer2_outputs(1196)) or (layer2_outputs(5181));
    layer3_outputs(393) <= not(layer2_outputs(3525));
    layer3_outputs(394) <= (layer2_outputs(5124)) and not (layer2_outputs(2100));
    layer3_outputs(395) <= (layer2_outputs(6441)) and not (layer2_outputs(3249));
    layer3_outputs(396) <= not((layer2_outputs(6269)) or (layer2_outputs(4681)));
    layer3_outputs(397) <= layer2_outputs(4833);
    layer3_outputs(398) <= '1';
    layer3_outputs(399) <= not(layer2_outputs(6974));
    layer3_outputs(400) <= not(layer2_outputs(5340));
    layer3_outputs(401) <= layer2_outputs(655);
    layer3_outputs(402) <= layer2_outputs(4228);
    layer3_outputs(403) <= layer2_outputs(2140);
    layer3_outputs(404) <= (layer2_outputs(6818)) and not (layer2_outputs(5231));
    layer3_outputs(405) <= not(layer2_outputs(1670));
    layer3_outputs(406) <= (layer2_outputs(6316)) and not (layer2_outputs(5221));
    layer3_outputs(407) <= not((layer2_outputs(7389)) xor (layer2_outputs(2211)));
    layer3_outputs(408) <= not((layer2_outputs(1140)) xor (layer2_outputs(2767)));
    layer3_outputs(409) <= layer2_outputs(1761);
    layer3_outputs(410) <= not((layer2_outputs(206)) and (layer2_outputs(3507)));
    layer3_outputs(411) <= not(layer2_outputs(7355));
    layer3_outputs(412) <= not(layer2_outputs(4277));
    layer3_outputs(413) <= not(layer2_outputs(3551)) or (layer2_outputs(1705));
    layer3_outputs(414) <= '1';
    layer3_outputs(415) <= layer2_outputs(2426);
    layer3_outputs(416) <= not(layer2_outputs(5239)) or (layer2_outputs(1143));
    layer3_outputs(417) <= not((layer2_outputs(3825)) and (layer2_outputs(613)));
    layer3_outputs(418) <= not((layer2_outputs(3794)) or (layer2_outputs(3391)));
    layer3_outputs(419) <= layer2_outputs(5215);
    layer3_outputs(420) <= not(layer2_outputs(2156));
    layer3_outputs(421) <= (layer2_outputs(1342)) and not (layer2_outputs(4984));
    layer3_outputs(422) <= layer2_outputs(5135);
    layer3_outputs(423) <= not((layer2_outputs(1549)) or (layer2_outputs(343)));
    layer3_outputs(424) <= (layer2_outputs(6448)) and not (layer2_outputs(107));
    layer3_outputs(425) <= layer2_outputs(2692);
    layer3_outputs(426) <= (layer2_outputs(2989)) and not (layer2_outputs(6135));
    layer3_outputs(427) <= not(layer2_outputs(564));
    layer3_outputs(428) <= not(layer2_outputs(4444));
    layer3_outputs(429) <= not(layer2_outputs(1894)) or (layer2_outputs(4446));
    layer3_outputs(430) <= (layer2_outputs(2737)) and not (layer2_outputs(6687));
    layer3_outputs(431) <= not((layer2_outputs(5978)) or (layer2_outputs(5093)));
    layer3_outputs(432) <= not(layer2_outputs(4102));
    layer3_outputs(433) <= not(layer2_outputs(7018));
    layer3_outputs(434) <= not(layer2_outputs(3577));
    layer3_outputs(435) <= layer2_outputs(2328);
    layer3_outputs(436) <= not(layer2_outputs(5312)) or (layer2_outputs(7289));
    layer3_outputs(437) <= not((layer2_outputs(502)) or (layer2_outputs(423)));
    layer3_outputs(438) <= not((layer2_outputs(2771)) xor (layer2_outputs(3258)));
    layer3_outputs(439) <= not(layer2_outputs(6772)) or (layer2_outputs(2142));
    layer3_outputs(440) <= layer2_outputs(6693);
    layer3_outputs(441) <= '1';
    layer3_outputs(442) <= (layer2_outputs(6751)) and not (layer2_outputs(6403));
    layer3_outputs(443) <= not(layer2_outputs(4806)) or (layer2_outputs(4563));
    layer3_outputs(444) <= not(layer2_outputs(4738));
    layer3_outputs(445) <= layer2_outputs(115);
    layer3_outputs(446) <= not(layer2_outputs(1358));
    layer3_outputs(447) <= (layer2_outputs(6993)) and (layer2_outputs(4625));
    layer3_outputs(448) <= '1';
    layer3_outputs(449) <= (layer2_outputs(2183)) and (layer2_outputs(329));
    layer3_outputs(450) <= not(layer2_outputs(5708));
    layer3_outputs(451) <= not((layer2_outputs(3864)) or (layer2_outputs(4432)));
    layer3_outputs(452) <= not(layer2_outputs(2969)) or (layer2_outputs(1009));
    layer3_outputs(453) <= not((layer2_outputs(2411)) or (layer2_outputs(5581)));
    layer3_outputs(454) <= layer2_outputs(897);
    layer3_outputs(455) <= not(layer2_outputs(4017));
    layer3_outputs(456) <= not(layer2_outputs(4904));
    layer3_outputs(457) <= (layer2_outputs(7400)) and (layer2_outputs(1119));
    layer3_outputs(458) <= '1';
    layer3_outputs(459) <= (layer2_outputs(7256)) and not (layer2_outputs(6483));
    layer3_outputs(460) <= (layer2_outputs(3012)) and not (layer2_outputs(118));
    layer3_outputs(461) <= (layer2_outputs(7376)) and not (layer2_outputs(6152));
    layer3_outputs(462) <= not(layer2_outputs(3978));
    layer3_outputs(463) <= not(layer2_outputs(7267));
    layer3_outputs(464) <= not(layer2_outputs(2578)) or (layer2_outputs(2304));
    layer3_outputs(465) <= layer2_outputs(4113);
    layer3_outputs(466) <= not(layer2_outputs(1963)) or (layer2_outputs(5430));
    layer3_outputs(467) <= (layer2_outputs(1469)) and not (layer2_outputs(3778));
    layer3_outputs(468) <= not((layer2_outputs(7099)) or (layer2_outputs(2351)));
    layer3_outputs(469) <= not(layer2_outputs(6944));
    layer3_outputs(470) <= layer2_outputs(6762);
    layer3_outputs(471) <= not(layer2_outputs(4674));
    layer3_outputs(472) <= not((layer2_outputs(3061)) or (layer2_outputs(4732)));
    layer3_outputs(473) <= layer2_outputs(7247);
    layer3_outputs(474) <= not(layer2_outputs(4970));
    layer3_outputs(475) <= layer2_outputs(3751);
    layer3_outputs(476) <= not((layer2_outputs(6267)) or (layer2_outputs(782)));
    layer3_outputs(477) <= not((layer2_outputs(3341)) or (layer2_outputs(6852)));
    layer3_outputs(478) <= not(layer2_outputs(7568)) or (layer2_outputs(5300));
    layer3_outputs(479) <= layer2_outputs(4810);
    layer3_outputs(480) <= '0';
    layer3_outputs(481) <= '0';
    layer3_outputs(482) <= (layer2_outputs(4069)) or (layer2_outputs(2242));
    layer3_outputs(483) <= layer2_outputs(7221);
    layer3_outputs(484) <= not(layer2_outputs(401));
    layer3_outputs(485) <= (layer2_outputs(4296)) and not (layer2_outputs(6758));
    layer3_outputs(486) <= not(layer2_outputs(4471)) or (layer2_outputs(6959));
    layer3_outputs(487) <= layer2_outputs(1078);
    layer3_outputs(488) <= not((layer2_outputs(5327)) or (layer2_outputs(6320)));
    layer3_outputs(489) <= not((layer2_outputs(453)) and (layer2_outputs(7615)));
    layer3_outputs(490) <= not(layer2_outputs(5787)) or (layer2_outputs(2500));
    layer3_outputs(491) <= (layer2_outputs(334)) and not (layer2_outputs(2951));
    layer3_outputs(492) <= not((layer2_outputs(3414)) or (layer2_outputs(5418)));
    layer3_outputs(493) <= not(layer2_outputs(3638));
    layer3_outputs(494) <= not(layer2_outputs(5741));
    layer3_outputs(495) <= '0';
    layer3_outputs(496) <= '1';
    layer3_outputs(497) <= not(layer2_outputs(3157));
    layer3_outputs(498) <= layer2_outputs(5874);
    layer3_outputs(499) <= not((layer2_outputs(6204)) or (layer2_outputs(3370)));
    layer3_outputs(500) <= not(layer2_outputs(4477));
    layer3_outputs(501) <= not(layer2_outputs(936));
    layer3_outputs(502) <= layer2_outputs(4213);
    layer3_outputs(503) <= not(layer2_outputs(6244)) or (layer2_outputs(6192));
    layer3_outputs(504) <= layer2_outputs(3784);
    layer3_outputs(505) <= not((layer2_outputs(5330)) or (layer2_outputs(7091)));
    layer3_outputs(506) <= (layer2_outputs(5450)) xor (layer2_outputs(3667));
    layer3_outputs(507) <= (layer2_outputs(3786)) and not (layer2_outputs(4007));
    layer3_outputs(508) <= layer2_outputs(3072);
    layer3_outputs(509) <= (layer2_outputs(2806)) and (layer2_outputs(4399));
    layer3_outputs(510) <= not(layer2_outputs(4926)) or (layer2_outputs(1787));
    layer3_outputs(511) <= layer2_outputs(3510);
    layer3_outputs(512) <= (layer2_outputs(79)) and (layer2_outputs(3510));
    layer3_outputs(513) <= not(layer2_outputs(3324)) or (layer2_outputs(232));
    layer3_outputs(514) <= layer2_outputs(1951);
    layer3_outputs(515) <= (layer2_outputs(6342)) and not (layer2_outputs(1210));
    layer3_outputs(516) <= (layer2_outputs(4405)) or (layer2_outputs(619));
    layer3_outputs(517) <= layer2_outputs(2138);
    layer3_outputs(518) <= layer2_outputs(59);
    layer3_outputs(519) <= not((layer2_outputs(3267)) and (layer2_outputs(1020)));
    layer3_outputs(520) <= layer2_outputs(2581);
    layer3_outputs(521) <= (layer2_outputs(3515)) or (layer2_outputs(1551));
    layer3_outputs(522) <= not(layer2_outputs(7003));
    layer3_outputs(523) <= (layer2_outputs(3694)) and not (layer2_outputs(3735));
    layer3_outputs(524) <= not(layer2_outputs(895));
    layer3_outputs(525) <= (layer2_outputs(1323)) and (layer2_outputs(2393));
    layer3_outputs(526) <= '0';
    layer3_outputs(527) <= (layer2_outputs(2893)) and not (layer2_outputs(5486));
    layer3_outputs(528) <= (layer2_outputs(1428)) and not (layer2_outputs(4637));
    layer3_outputs(529) <= not(layer2_outputs(3070)) or (layer2_outputs(2905));
    layer3_outputs(530) <= layer2_outputs(7637);
    layer3_outputs(531) <= (layer2_outputs(2652)) xor (layer2_outputs(7332));
    layer3_outputs(532) <= not(layer2_outputs(2006));
    layer3_outputs(533) <= (layer2_outputs(3684)) and not (layer2_outputs(1189));
    layer3_outputs(534) <= not((layer2_outputs(1491)) or (layer2_outputs(5396)));
    layer3_outputs(535) <= not(layer2_outputs(5013)) or (layer2_outputs(6837));
    layer3_outputs(536) <= '0';
    layer3_outputs(537) <= (layer2_outputs(7457)) and (layer2_outputs(6034));
    layer3_outputs(538) <= (layer2_outputs(1210)) xor (layer2_outputs(2145));
    layer3_outputs(539) <= (layer2_outputs(7157)) and (layer2_outputs(1769));
    layer3_outputs(540) <= not(layer2_outputs(3077));
    layer3_outputs(541) <= not(layer2_outputs(1021));
    layer3_outputs(542) <= not((layer2_outputs(3970)) and (layer2_outputs(2914)));
    layer3_outputs(543) <= (layer2_outputs(2906)) and not (layer2_outputs(625));
    layer3_outputs(544) <= not(layer2_outputs(1198));
    layer3_outputs(545) <= layer2_outputs(1052);
    layer3_outputs(546) <= not((layer2_outputs(4308)) and (layer2_outputs(5153)));
    layer3_outputs(547) <= (layer2_outputs(5806)) or (layer2_outputs(6160));
    layer3_outputs(548) <= layer2_outputs(7331);
    layer3_outputs(549) <= not(layer2_outputs(2724)) or (layer2_outputs(5978));
    layer3_outputs(550) <= not((layer2_outputs(1572)) or (layer2_outputs(5522)));
    layer3_outputs(551) <= not(layer2_outputs(281));
    layer3_outputs(552) <= not((layer2_outputs(3907)) or (layer2_outputs(5807)));
    layer3_outputs(553) <= (layer2_outputs(4881)) and not (layer2_outputs(5224));
    layer3_outputs(554) <= layer2_outputs(3697);
    layer3_outputs(555) <= not(layer2_outputs(4543)) or (layer2_outputs(6468));
    layer3_outputs(556) <= (layer2_outputs(1182)) and not (layer2_outputs(185));
    layer3_outputs(557) <= (layer2_outputs(6368)) and (layer2_outputs(4312));
    layer3_outputs(558) <= layer2_outputs(847);
    layer3_outputs(559) <= layer2_outputs(188);
    layer3_outputs(560) <= (layer2_outputs(5681)) or (layer2_outputs(3844));
    layer3_outputs(561) <= (layer2_outputs(1179)) and not (layer2_outputs(7210));
    layer3_outputs(562) <= (layer2_outputs(4780)) and not (layer2_outputs(705));
    layer3_outputs(563) <= layer2_outputs(7282);
    layer3_outputs(564) <= not(layer2_outputs(6743)) or (layer2_outputs(3151));
    layer3_outputs(565) <= layer2_outputs(4998);
    layer3_outputs(566) <= (layer2_outputs(3024)) and not (layer2_outputs(1306));
    layer3_outputs(567) <= not(layer2_outputs(6067)) or (layer2_outputs(6846));
    layer3_outputs(568) <= (layer2_outputs(5819)) xor (layer2_outputs(1748));
    layer3_outputs(569) <= (layer2_outputs(6756)) xor (layer2_outputs(4365));
    layer3_outputs(570) <= layer2_outputs(4832);
    layer3_outputs(571) <= layer2_outputs(4162);
    layer3_outputs(572) <= (layer2_outputs(3161)) and not (layer2_outputs(5967));
    layer3_outputs(573) <= not((layer2_outputs(3381)) xor (layer2_outputs(6540)));
    layer3_outputs(574) <= layer2_outputs(6991);
    layer3_outputs(575) <= (layer2_outputs(3548)) and not (layer2_outputs(4585));
    layer3_outputs(576) <= '0';
    layer3_outputs(577) <= (layer2_outputs(884)) or (layer2_outputs(1348));
    layer3_outputs(578) <= '1';
    layer3_outputs(579) <= layer2_outputs(456);
    layer3_outputs(580) <= (layer2_outputs(2166)) and not (layer2_outputs(5860));
    layer3_outputs(581) <= not((layer2_outputs(5595)) or (layer2_outputs(3385)));
    layer3_outputs(582) <= (layer2_outputs(5095)) and (layer2_outputs(1051));
    layer3_outputs(583) <= (layer2_outputs(2960)) and (layer2_outputs(5885));
    layer3_outputs(584) <= not(layer2_outputs(6765));
    layer3_outputs(585) <= layer2_outputs(757);
    layer3_outputs(586) <= (layer2_outputs(7677)) or (layer2_outputs(4880));
    layer3_outputs(587) <= layer2_outputs(4981);
    layer3_outputs(588) <= not(layer2_outputs(1247));
    layer3_outputs(589) <= not(layer2_outputs(659));
    layer3_outputs(590) <= layer2_outputs(5438);
    layer3_outputs(591) <= not((layer2_outputs(6824)) or (layer2_outputs(3087)));
    layer3_outputs(592) <= layer2_outputs(7046);
    layer3_outputs(593) <= (layer2_outputs(3486)) and (layer2_outputs(3950));
    layer3_outputs(594) <= not(layer2_outputs(4488));
    layer3_outputs(595) <= layer2_outputs(230);
    layer3_outputs(596) <= not(layer2_outputs(4841)) or (layer2_outputs(423));
    layer3_outputs(597) <= (layer2_outputs(808)) or (layer2_outputs(6832));
    layer3_outputs(598) <= (layer2_outputs(5419)) and not (layer2_outputs(5859));
    layer3_outputs(599) <= '0';
    layer3_outputs(600) <= not(layer2_outputs(7530)) or (layer2_outputs(5852));
    layer3_outputs(601) <= (layer2_outputs(1629)) and (layer2_outputs(7255));
    layer3_outputs(602) <= (layer2_outputs(3287)) and not (layer2_outputs(1839));
    layer3_outputs(603) <= (layer2_outputs(2364)) and not (layer2_outputs(1675));
    layer3_outputs(604) <= layer2_outputs(3697);
    layer3_outputs(605) <= not((layer2_outputs(110)) or (layer2_outputs(1528)));
    layer3_outputs(606) <= layer2_outputs(7165);
    layer3_outputs(607) <= layer2_outputs(2384);
    layer3_outputs(608) <= not(layer2_outputs(6951));
    layer3_outputs(609) <= not(layer2_outputs(1525));
    layer3_outputs(610) <= layer2_outputs(1921);
    layer3_outputs(611) <= not(layer2_outputs(1702));
    layer3_outputs(612) <= (layer2_outputs(5805)) and not (layer2_outputs(5468));
    layer3_outputs(613) <= not(layer2_outputs(5175));
    layer3_outputs(614) <= '0';
    layer3_outputs(615) <= (layer2_outputs(504)) and not (layer2_outputs(7656));
    layer3_outputs(616) <= not(layer2_outputs(7670));
    layer3_outputs(617) <= (layer2_outputs(2577)) and not (layer2_outputs(7619));
    layer3_outputs(618) <= not(layer2_outputs(6685));
    layer3_outputs(619) <= (layer2_outputs(5270)) and not (layer2_outputs(5172));
    layer3_outputs(620) <= (layer2_outputs(285)) and (layer2_outputs(5542));
    layer3_outputs(621) <= not(layer2_outputs(2913));
    layer3_outputs(622) <= not(layer2_outputs(1097));
    layer3_outputs(623) <= not(layer2_outputs(5056));
    layer3_outputs(624) <= not(layer2_outputs(5380));
    layer3_outputs(625) <= not(layer2_outputs(6840));
    layer3_outputs(626) <= layer2_outputs(3668);
    layer3_outputs(627) <= not((layer2_outputs(5166)) or (layer2_outputs(3995)));
    layer3_outputs(628) <= not(layer2_outputs(5236));
    layer3_outputs(629) <= (layer2_outputs(6755)) and (layer2_outputs(586));
    layer3_outputs(630) <= not((layer2_outputs(6360)) xor (layer2_outputs(3080)));
    layer3_outputs(631) <= (layer2_outputs(5451)) and not (layer2_outputs(3620));
    layer3_outputs(632) <= '0';
    layer3_outputs(633) <= layer2_outputs(6910);
    layer3_outputs(634) <= not((layer2_outputs(6426)) or (layer2_outputs(2579)));
    layer3_outputs(635) <= layer2_outputs(2814);
    layer3_outputs(636) <= (layer2_outputs(5364)) and not (layer2_outputs(3212));
    layer3_outputs(637) <= not(layer2_outputs(7528));
    layer3_outputs(638) <= not((layer2_outputs(290)) and (layer2_outputs(3073)));
    layer3_outputs(639) <= (layer2_outputs(3526)) xor (layer2_outputs(5516));
    layer3_outputs(640) <= not(layer2_outputs(6791));
    layer3_outputs(641) <= not((layer2_outputs(7352)) and (layer2_outputs(3626)));
    layer3_outputs(642) <= not(layer2_outputs(213));
    layer3_outputs(643) <= not(layer2_outputs(2561));
    layer3_outputs(644) <= not(layer2_outputs(1352));
    layer3_outputs(645) <= (layer2_outputs(312)) and not (layer2_outputs(5496));
    layer3_outputs(646) <= (layer2_outputs(3667)) and not (layer2_outputs(4333));
    layer3_outputs(647) <= not(layer2_outputs(3708)) or (layer2_outputs(4248));
    layer3_outputs(648) <= not(layer2_outputs(4042));
    layer3_outputs(649) <= not(layer2_outputs(5887));
    layer3_outputs(650) <= not((layer2_outputs(6085)) and (layer2_outputs(738)));
    layer3_outputs(651) <= (layer2_outputs(5402)) and not (layer2_outputs(3360));
    layer3_outputs(652) <= not(layer2_outputs(242));
    layer3_outputs(653) <= not((layer2_outputs(1006)) or (layer2_outputs(7638)));
    layer3_outputs(654) <= layer2_outputs(1294);
    layer3_outputs(655) <= (layer2_outputs(4468)) and (layer2_outputs(6787));
    layer3_outputs(656) <= layer2_outputs(3188);
    layer3_outputs(657) <= (layer2_outputs(5578)) and not (layer2_outputs(3437));
    layer3_outputs(658) <= (layer2_outputs(5829)) and not (layer2_outputs(1637));
    layer3_outputs(659) <= layer2_outputs(7516);
    layer3_outputs(660) <= not(layer2_outputs(6697));
    layer3_outputs(661) <= not(layer2_outputs(5534));
    layer3_outputs(662) <= layer2_outputs(4255);
    layer3_outputs(663) <= not(layer2_outputs(1914));
    layer3_outputs(664) <= (layer2_outputs(5128)) and not (layer2_outputs(5780));
    layer3_outputs(665) <= not(layer2_outputs(4451)) or (layer2_outputs(6905));
    layer3_outputs(666) <= not((layer2_outputs(5248)) xor (layer2_outputs(1412)));
    layer3_outputs(667) <= not(layer2_outputs(6268));
    layer3_outputs(668) <= not((layer2_outputs(1845)) and (layer2_outputs(2612)));
    layer3_outputs(669) <= (layer2_outputs(2993)) and not (layer2_outputs(1220));
    layer3_outputs(670) <= not((layer2_outputs(2207)) xor (layer2_outputs(5121)));
    layer3_outputs(671) <= (layer2_outputs(7399)) and not (layer2_outputs(1842));
    layer3_outputs(672) <= (layer2_outputs(2419)) and not (layer2_outputs(676));
    layer3_outputs(673) <= not(layer2_outputs(3445));
    layer3_outputs(674) <= not(layer2_outputs(6769));
    layer3_outputs(675) <= not((layer2_outputs(5107)) xor (layer2_outputs(393)));
    layer3_outputs(676) <= not(layer2_outputs(911)) or (layer2_outputs(2242));
    layer3_outputs(677) <= not(layer2_outputs(6454));
    layer3_outputs(678) <= not(layer2_outputs(1830)) or (layer2_outputs(3523));
    layer3_outputs(679) <= (layer2_outputs(5999)) or (layer2_outputs(5043));
    layer3_outputs(680) <= (layer2_outputs(3518)) or (layer2_outputs(5185));
    layer3_outputs(681) <= layer2_outputs(2167);
    layer3_outputs(682) <= not(layer2_outputs(1806));
    layer3_outputs(683) <= not(layer2_outputs(56));
    layer3_outputs(684) <= not(layer2_outputs(6579));
    layer3_outputs(685) <= layer2_outputs(2575);
    layer3_outputs(686) <= '1';
    layer3_outputs(687) <= (layer2_outputs(2942)) and not (layer2_outputs(4209));
    layer3_outputs(688) <= not(layer2_outputs(4073));
    layer3_outputs(689) <= (layer2_outputs(2216)) or (layer2_outputs(6915));
    layer3_outputs(690) <= (layer2_outputs(5856)) and (layer2_outputs(653));
    layer3_outputs(691) <= '0';
    layer3_outputs(692) <= not(layer2_outputs(3845));
    layer3_outputs(693) <= not(layer2_outputs(5363)) or (layer2_outputs(7370));
    layer3_outputs(694) <= not((layer2_outputs(6195)) or (layer2_outputs(3718)));
    layer3_outputs(695) <= layer2_outputs(1451);
    layer3_outputs(696) <= layer2_outputs(127);
    layer3_outputs(697) <= (layer2_outputs(4695)) and not (layer2_outputs(1054));
    layer3_outputs(698) <= not((layer2_outputs(1065)) or (layer2_outputs(2314)));
    layer3_outputs(699) <= not(layer2_outputs(1133));
    layer3_outputs(700) <= (layer2_outputs(1782)) and (layer2_outputs(4633));
    layer3_outputs(701) <= not(layer2_outputs(2897));
    layer3_outputs(702) <= layer2_outputs(7291);
    layer3_outputs(703) <= (layer2_outputs(4816)) or (layer2_outputs(5033));
    layer3_outputs(704) <= (layer2_outputs(2369)) xor (layer2_outputs(2794));
    layer3_outputs(705) <= not(layer2_outputs(2787)) or (layer2_outputs(2390));
    layer3_outputs(706) <= not(layer2_outputs(5009));
    layer3_outputs(707) <= (layer2_outputs(1007)) and not (layer2_outputs(7601));
    layer3_outputs(708) <= layer2_outputs(3501);
    layer3_outputs(709) <= not(layer2_outputs(1611)) or (layer2_outputs(7468));
    layer3_outputs(710) <= not(layer2_outputs(4931)) or (layer2_outputs(7675));
    layer3_outputs(711) <= '0';
    layer3_outputs(712) <= (layer2_outputs(6532)) xor (layer2_outputs(4432));
    layer3_outputs(713) <= '0';
    layer3_outputs(714) <= not(layer2_outputs(4159));
    layer3_outputs(715) <= not(layer2_outputs(4302)) or (layer2_outputs(6010));
    layer3_outputs(716) <= not(layer2_outputs(3868)) or (layer2_outputs(3946));
    layer3_outputs(717) <= not((layer2_outputs(5374)) xor (layer2_outputs(3174)));
    layer3_outputs(718) <= (layer2_outputs(4064)) xor (layer2_outputs(2841));
    layer3_outputs(719) <= not(layer2_outputs(5424));
    layer3_outputs(720) <= not(layer2_outputs(6651));
    layer3_outputs(721) <= layer2_outputs(3799);
    layer3_outputs(722) <= not(layer2_outputs(415)) or (layer2_outputs(958));
    layer3_outputs(723) <= not(layer2_outputs(6599));
    layer3_outputs(724) <= not(layer2_outputs(4707));
    layer3_outputs(725) <= '0';
    layer3_outputs(726) <= layer2_outputs(665);
    layer3_outputs(727) <= layer2_outputs(3477);
    layer3_outputs(728) <= not(layer2_outputs(3937));
    layer3_outputs(729) <= not((layer2_outputs(6444)) and (layer2_outputs(7260)));
    layer3_outputs(730) <= (layer2_outputs(6070)) and not (layer2_outputs(4051));
    layer3_outputs(731) <= (layer2_outputs(7557)) or (layer2_outputs(1345));
    layer3_outputs(732) <= not(layer2_outputs(7531));
    layer3_outputs(733) <= not(layer2_outputs(3859)) or (layer2_outputs(1325));
    layer3_outputs(734) <= not((layer2_outputs(3630)) and (layer2_outputs(6428)));
    layer3_outputs(735) <= (layer2_outputs(1934)) and not (layer2_outputs(3611));
    layer3_outputs(736) <= layer2_outputs(7534);
    layer3_outputs(737) <= (layer2_outputs(2003)) and not (layer2_outputs(2996));
    layer3_outputs(738) <= layer2_outputs(2230);
    layer3_outputs(739) <= layer2_outputs(2775);
    layer3_outputs(740) <= not(layer2_outputs(7587));
    layer3_outputs(741) <= not(layer2_outputs(103));
    layer3_outputs(742) <= (layer2_outputs(464)) or (layer2_outputs(4141));
    layer3_outputs(743) <= layer2_outputs(4210);
    layer3_outputs(744) <= not(layer2_outputs(6440));
    layer3_outputs(745) <= not((layer2_outputs(1046)) and (layer2_outputs(3613)));
    layer3_outputs(746) <= layer2_outputs(2691);
    layer3_outputs(747) <= layer2_outputs(6348);
    layer3_outputs(748) <= layer2_outputs(2045);
    layer3_outputs(749) <= not(layer2_outputs(7523)) or (layer2_outputs(6634));
    layer3_outputs(750) <= not((layer2_outputs(5355)) and (layer2_outputs(4068)));
    layer3_outputs(751) <= not(layer2_outputs(3690)) or (layer2_outputs(7067));
    layer3_outputs(752) <= (layer2_outputs(1262)) and not (layer2_outputs(7600));
    layer3_outputs(753) <= not(layer2_outputs(1891));
    layer3_outputs(754) <= (layer2_outputs(5596)) and (layer2_outputs(1907));
    layer3_outputs(755) <= layer2_outputs(3113);
    layer3_outputs(756) <= not(layer2_outputs(4826));
    layer3_outputs(757) <= not(layer2_outputs(6716));
    layer3_outputs(758) <= (layer2_outputs(6222)) and not (layer2_outputs(889));
    layer3_outputs(759) <= layer2_outputs(832);
    layer3_outputs(760) <= not((layer2_outputs(2296)) or (layer2_outputs(3879)));
    layer3_outputs(761) <= not(layer2_outputs(6499)) or (layer2_outputs(5113));
    layer3_outputs(762) <= (layer2_outputs(82)) and (layer2_outputs(7512));
    layer3_outputs(763) <= not(layer2_outputs(227));
    layer3_outputs(764) <= not(layer2_outputs(6790));
    layer3_outputs(765) <= not((layer2_outputs(5665)) and (layer2_outputs(6292)));
    layer3_outputs(766) <= (layer2_outputs(6302)) and (layer2_outputs(4883));
    layer3_outputs(767) <= not(layer2_outputs(7205)) or (layer2_outputs(2060));
    layer3_outputs(768) <= (layer2_outputs(3586)) and (layer2_outputs(7020));
    layer3_outputs(769) <= layer2_outputs(7148);
    layer3_outputs(770) <= (layer2_outputs(5436)) and not (layer2_outputs(7511));
    layer3_outputs(771) <= not(layer2_outputs(1968));
    layer3_outputs(772) <= not(layer2_outputs(4979)) or (layer2_outputs(4996));
    layer3_outputs(773) <= layer2_outputs(2563);
    layer3_outputs(774) <= not((layer2_outputs(4395)) and (layer2_outputs(1279)));
    layer3_outputs(775) <= layer2_outputs(1804);
    layer3_outputs(776) <= layer2_outputs(3241);
    layer3_outputs(777) <= not(layer2_outputs(5723));
    layer3_outputs(778) <= layer2_outputs(5446);
    layer3_outputs(779) <= not((layer2_outputs(5803)) or (layer2_outputs(4056)));
    layer3_outputs(780) <= not((layer2_outputs(6070)) or (layer2_outputs(298)));
    layer3_outputs(781) <= (layer2_outputs(1572)) and (layer2_outputs(2659));
    layer3_outputs(782) <= not(layer2_outputs(4422));
    layer3_outputs(783) <= not(layer2_outputs(3369));
    layer3_outputs(784) <= layer2_outputs(3905);
    layer3_outputs(785) <= not(layer2_outputs(5607));
    layer3_outputs(786) <= '0';
    layer3_outputs(787) <= layer2_outputs(5528);
    layer3_outputs(788) <= not(layer2_outputs(5093));
    layer3_outputs(789) <= not(layer2_outputs(1788)) or (layer2_outputs(6008));
    layer3_outputs(790) <= '0';
    layer3_outputs(791) <= not(layer2_outputs(7156)) or (layer2_outputs(3816));
    layer3_outputs(792) <= (layer2_outputs(6049)) and (layer2_outputs(2112));
    layer3_outputs(793) <= not(layer2_outputs(1819));
    layer3_outputs(794) <= (layer2_outputs(6670)) and not (layer2_outputs(691));
    layer3_outputs(795) <= layer2_outputs(5353);
    layer3_outputs(796) <= (layer2_outputs(3788)) or (layer2_outputs(6477));
    layer3_outputs(797) <= not(layer2_outputs(1686));
    layer3_outputs(798) <= not(layer2_outputs(6388)) or (layer2_outputs(5066));
    layer3_outputs(799) <= (layer2_outputs(6875)) and (layer2_outputs(4902));
    layer3_outputs(800) <= not(layer2_outputs(5428)) or (layer2_outputs(7278));
    layer3_outputs(801) <= not(layer2_outputs(485)) or (layer2_outputs(2815));
    layer3_outputs(802) <= layer2_outputs(2431);
    layer3_outputs(803) <= layer2_outputs(5399);
    layer3_outputs(804) <= not((layer2_outputs(821)) or (layer2_outputs(3315)));
    layer3_outputs(805) <= (layer2_outputs(3233)) and (layer2_outputs(7179));
    layer3_outputs(806) <= (layer2_outputs(3587)) and not (layer2_outputs(7658));
    layer3_outputs(807) <= layer2_outputs(1066);
    layer3_outputs(808) <= not(layer2_outputs(4208));
    layer3_outputs(809) <= not(layer2_outputs(5352)) or (layer2_outputs(64));
    layer3_outputs(810) <= not(layer2_outputs(744));
    layer3_outputs(811) <= (layer2_outputs(7643)) and (layer2_outputs(921));
    layer3_outputs(812) <= layer2_outputs(6543);
    layer3_outputs(813) <= (layer2_outputs(1089)) or (layer2_outputs(4667));
    layer3_outputs(814) <= not(layer2_outputs(245)) or (layer2_outputs(3141));
    layer3_outputs(815) <= (layer2_outputs(7201)) and not (layer2_outputs(5675));
    layer3_outputs(816) <= (layer2_outputs(921)) and (layer2_outputs(6873));
    layer3_outputs(817) <= (layer2_outputs(1155)) and not (layer2_outputs(3003));
    layer3_outputs(818) <= not(layer2_outputs(5387)) or (layer2_outputs(3411));
    layer3_outputs(819) <= not((layer2_outputs(481)) and (layer2_outputs(1822)));
    layer3_outputs(820) <= not(layer2_outputs(4366)) or (layer2_outputs(5982));
    layer3_outputs(821) <= layer2_outputs(6832);
    layer3_outputs(822) <= layer2_outputs(1878);
    layer3_outputs(823) <= not(layer2_outputs(7636));
    layer3_outputs(824) <= layer2_outputs(6525);
    layer3_outputs(825) <= layer2_outputs(7327);
    layer3_outputs(826) <= (layer2_outputs(4873)) and not (layer2_outputs(6614));
    layer3_outputs(827) <= not(layer2_outputs(5887));
    layer3_outputs(828) <= (layer2_outputs(835)) and (layer2_outputs(6164));
    layer3_outputs(829) <= not(layer2_outputs(427));
    layer3_outputs(830) <= (layer2_outputs(16)) or (layer2_outputs(3224));
    layer3_outputs(831) <= '0';
    layer3_outputs(832) <= (layer2_outputs(6899)) xor (layer2_outputs(493));
    layer3_outputs(833) <= (layer2_outputs(6644)) and not (layer2_outputs(6386));
    layer3_outputs(834) <= not(layer2_outputs(130));
    layer3_outputs(835) <= (layer2_outputs(5390)) and not (layer2_outputs(292));
    layer3_outputs(836) <= (layer2_outputs(1824)) and not (layer2_outputs(147));
    layer3_outputs(837) <= (layer2_outputs(5127)) and not (layer2_outputs(1402));
    layer3_outputs(838) <= '0';
    layer3_outputs(839) <= not(layer2_outputs(2823));
    layer3_outputs(840) <= (layer2_outputs(4502)) and not (layer2_outputs(4470));
    layer3_outputs(841) <= '1';
    layer3_outputs(842) <= not((layer2_outputs(6610)) or (layer2_outputs(2607)));
    layer3_outputs(843) <= not(layer2_outputs(5143));
    layer3_outputs(844) <= (layer2_outputs(385)) and (layer2_outputs(3494));
    layer3_outputs(845) <= layer2_outputs(1813);
    layer3_outputs(846) <= (layer2_outputs(1284)) and not (layer2_outputs(3233));
    layer3_outputs(847) <= (layer2_outputs(3122)) and (layer2_outputs(1596));
    layer3_outputs(848) <= not(layer2_outputs(1872)) or (layer2_outputs(5316));
    layer3_outputs(849) <= not((layer2_outputs(1432)) or (layer2_outputs(1375)));
    layer3_outputs(850) <= (layer2_outputs(2801)) xor (layer2_outputs(2469));
    layer3_outputs(851) <= not(layer2_outputs(6147));
    layer3_outputs(852) <= not(layer2_outputs(711));
    layer3_outputs(853) <= not((layer2_outputs(4449)) and (layer2_outputs(7352)));
    layer3_outputs(854) <= not(layer2_outputs(149));
    layer3_outputs(855) <= layer2_outputs(3494);
    layer3_outputs(856) <= not(layer2_outputs(4616)) or (layer2_outputs(5989));
    layer3_outputs(857) <= not(layer2_outputs(6533)) or (layer2_outputs(4746));
    layer3_outputs(858) <= not(layer2_outputs(5591));
    layer3_outputs(859) <= not(layer2_outputs(7423));
    layer3_outputs(860) <= (layer2_outputs(1728)) and not (layer2_outputs(3172));
    layer3_outputs(861) <= (layer2_outputs(4715)) xor (layer2_outputs(6162));
    layer3_outputs(862) <= not((layer2_outputs(2786)) xor (layer2_outputs(4875)));
    layer3_outputs(863) <= (layer2_outputs(2840)) and (layer2_outputs(5593));
    layer3_outputs(864) <= not(layer2_outputs(5124));
    layer3_outputs(865) <= (layer2_outputs(4094)) xor (layer2_outputs(5374));
    layer3_outputs(866) <= not(layer2_outputs(918));
    layer3_outputs(867) <= layer2_outputs(3172);
    layer3_outputs(868) <= (layer2_outputs(109)) or (layer2_outputs(138));
    layer3_outputs(869) <= not(layer2_outputs(1320)) or (layer2_outputs(2107));
    layer3_outputs(870) <= not(layer2_outputs(5339));
    layer3_outputs(871) <= (layer2_outputs(3623)) and (layer2_outputs(5563));
    layer3_outputs(872) <= not(layer2_outputs(4773));
    layer3_outputs(873) <= not(layer2_outputs(2609));
    layer3_outputs(874) <= layer2_outputs(1013);
    layer3_outputs(875) <= '1';
    layer3_outputs(876) <= not(layer2_outputs(3979)) or (layer2_outputs(6287));
    layer3_outputs(877) <= not(layer2_outputs(6525));
    layer3_outputs(878) <= not(layer2_outputs(7383));
    layer3_outputs(879) <= not(layer2_outputs(2039));
    layer3_outputs(880) <= not(layer2_outputs(6856)) or (layer2_outputs(816));
    layer3_outputs(881) <= layer2_outputs(2650);
    layer3_outputs(882) <= not(layer2_outputs(1554)) or (layer2_outputs(6168));
    layer3_outputs(883) <= (layer2_outputs(4425)) and not (layer2_outputs(1771));
    layer3_outputs(884) <= not(layer2_outputs(4372));
    layer3_outputs(885) <= (layer2_outputs(2853)) or (layer2_outputs(6369));
    layer3_outputs(886) <= '1';
    layer3_outputs(887) <= '1';
    layer3_outputs(888) <= (layer2_outputs(4224)) or (layer2_outputs(5440));
    layer3_outputs(889) <= layer2_outputs(4487);
    layer3_outputs(890) <= not(layer2_outputs(5857)) or (layer2_outputs(6175));
    layer3_outputs(891) <= (layer2_outputs(5559)) and not (layer2_outputs(6759));
    layer3_outputs(892) <= not((layer2_outputs(3529)) or (layer2_outputs(2246)));
    layer3_outputs(893) <= layer2_outputs(4603);
    layer3_outputs(894) <= layer2_outputs(5748);
    layer3_outputs(895) <= not(layer2_outputs(3565));
    layer3_outputs(896) <= not((layer2_outputs(5984)) and (layer2_outputs(7261)));
    layer3_outputs(897) <= not((layer2_outputs(6914)) and (layer2_outputs(833)));
    layer3_outputs(898) <= (layer2_outputs(6683)) and not (layer2_outputs(734));
    layer3_outputs(899) <= (layer2_outputs(3460)) and (layer2_outputs(2707));
    layer3_outputs(900) <= layer2_outputs(4779);
    layer3_outputs(901) <= not(layer2_outputs(7216)) or (layer2_outputs(5643));
    layer3_outputs(902) <= (layer2_outputs(4287)) and not (layer2_outputs(2547));
    layer3_outputs(903) <= (layer2_outputs(5841)) xor (layer2_outputs(524));
    layer3_outputs(904) <= layer2_outputs(1374);
    layer3_outputs(905) <= not(layer2_outputs(5052));
    layer3_outputs(906) <= not(layer2_outputs(108));
    layer3_outputs(907) <= layer2_outputs(2976);
    layer3_outputs(908) <= not((layer2_outputs(1984)) or (layer2_outputs(4816)));
    layer3_outputs(909) <= (layer2_outputs(7666)) and not (layer2_outputs(1571));
    layer3_outputs(910) <= not(layer2_outputs(4604)) or (layer2_outputs(4942));
    layer3_outputs(911) <= not((layer2_outputs(7604)) xor (layer2_outputs(6100)));
    layer3_outputs(912) <= not((layer2_outputs(2823)) and (layer2_outputs(339)));
    layer3_outputs(913) <= (layer2_outputs(6365)) and not (layer2_outputs(2289));
    layer3_outputs(914) <= (layer2_outputs(7064)) and (layer2_outputs(6799));
    layer3_outputs(915) <= layer2_outputs(1764);
    layer3_outputs(916) <= not(layer2_outputs(3521));
    layer3_outputs(917) <= not((layer2_outputs(2024)) and (layer2_outputs(1243)));
    layer3_outputs(918) <= not(layer2_outputs(4467));
    layer3_outputs(919) <= layer2_outputs(4683);
    layer3_outputs(920) <= not((layer2_outputs(429)) and (layer2_outputs(1757)));
    layer3_outputs(921) <= not(layer2_outputs(4156)) or (layer2_outputs(2340));
    layer3_outputs(922) <= not(layer2_outputs(5592)) or (layer2_outputs(7477));
    layer3_outputs(923) <= (layer2_outputs(6361)) and not (layer2_outputs(1268));
    layer3_outputs(924) <= not((layer2_outputs(331)) and (layer2_outputs(6647)));
    layer3_outputs(925) <= not((layer2_outputs(5531)) or (layer2_outputs(230)));
    layer3_outputs(926) <= not(layer2_outputs(213));
    layer3_outputs(927) <= not((layer2_outputs(4668)) xor (layer2_outputs(4730)));
    layer3_outputs(928) <= (layer2_outputs(4792)) and (layer2_outputs(6797));
    layer3_outputs(929) <= not(layer2_outputs(1801)) or (layer2_outputs(2094));
    layer3_outputs(930) <= not((layer2_outputs(50)) or (layer2_outputs(3582)));
    layer3_outputs(931) <= not(layer2_outputs(3161));
    layer3_outputs(932) <= not(layer2_outputs(3779)) or (layer2_outputs(1555));
    layer3_outputs(933) <= (layer2_outputs(5836)) xor (layer2_outputs(351));
    layer3_outputs(934) <= (layer2_outputs(6599)) and not (layer2_outputs(7063));
    layer3_outputs(935) <= (layer2_outputs(5829)) and not (layer2_outputs(5472));
    layer3_outputs(936) <= layer2_outputs(1995);
    layer3_outputs(937) <= (layer2_outputs(3537)) and not (layer2_outputs(4220));
    layer3_outputs(938) <= layer2_outputs(5285);
    layer3_outputs(939) <= not((layer2_outputs(5154)) and (layer2_outputs(5098)));
    layer3_outputs(940) <= not((layer2_outputs(1731)) and (layer2_outputs(1965)));
    layer3_outputs(941) <= layer2_outputs(1047);
    layer3_outputs(942) <= not((layer2_outputs(6398)) and (layer2_outputs(7123)));
    layer3_outputs(943) <= not(layer2_outputs(4504)) or (layer2_outputs(4648));
    layer3_outputs(944) <= (layer2_outputs(7342)) or (layer2_outputs(2029));
    layer3_outputs(945) <= (layer2_outputs(3785)) or (layer2_outputs(4678));
    layer3_outputs(946) <= (layer2_outputs(7676)) xor (layer2_outputs(4739));
    layer3_outputs(947) <= '0';
    layer3_outputs(948) <= layer2_outputs(1820);
    layer3_outputs(949) <= (layer2_outputs(3937)) and not (layer2_outputs(1877));
    layer3_outputs(950) <= not(layer2_outputs(6844));
    layer3_outputs(951) <= not(layer2_outputs(3160)) or (layer2_outputs(6572));
    layer3_outputs(952) <= (layer2_outputs(6489)) or (layer2_outputs(1947));
    layer3_outputs(953) <= (layer2_outputs(5982)) xor (layer2_outputs(3379));
    layer3_outputs(954) <= layer2_outputs(345);
    layer3_outputs(955) <= layer2_outputs(474);
    layer3_outputs(956) <= layer2_outputs(6778);
    layer3_outputs(957) <= '0';
    layer3_outputs(958) <= layer2_outputs(3436);
    layer3_outputs(959) <= not((layer2_outputs(5447)) and (layer2_outputs(1307)));
    layer3_outputs(960) <= not(layer2_outputs(7607)) or (layer2_outputs(5678));
    layer3_outputs(961) <= not(layer2_outputs(36));
    layer3_outputs(962) <= layer2_outputs(6605);
    layer3_outputs(963) <= not(layer2_outputs(2441));
    layer3_outputs(964) <= layer2_outputs(3377);
    layer3_outputs(965) <= not((layer2_outputs(4196)) or (layer2_outputs(2488)));
    layer3_outputs(966) <= layer2_outputs(1034);
    layer3_outputs(967) <= not(layer2_outputs(1642));
    layer3_outputs(968) <= not(layer2_outputs(1596));
    layer3_outputs(969) <= layer2_outputs(2057);
    layer3_outputs(970) <= not(layer2_outputs(823));
    layer3_outputs(971) <= not(layer2_outputs(5684));
    layer3_outputs(972) <= not(layer2_outputs(3285));
    layer3_outputs(973) <= '1';
    layer3_outputs(974) <= not(layer2_outputs(6635));
    layer3_outputs(975) <= (layer2_outputs(135)) or (layer2_outputs(584));
    layer3_outputs(976) <= '1';
    layer3_outputs(977) <= not(layer2_outputs(3917));
    layer3_outputs(978) <= not(layer2_outputs(7174)) or (layer2_outputs(3532));
    layer3_outputs(979) <= (layer2_outputs(1651)) or (layer2_outputs(951));
    layer3_outputs(980) <= not((layer2_outputs(6795)) or (layer2_outputs(2091)));
    layer3_outputs(981) <= layer2_outputs(7616);
    layer3_outputs(982) <= not(layer2_outputs(3673));
    layer3_outputs(983) <= not((layer2_outputs(3179)) or (layer2_outputs(2173)));
    layer3_outputs(984) <= (layer2_outputs(5108)) and not (layer2_outputs(5098));
    layer3_outputs(985) <= (layer2_outputs(4368)) and not (layer2_outputs(1470));
    layer3_outputs(986) <= not(layer2_outputs(4352)) or (layer2_outputs(3389));
    layer3_outputs(987) <= not(layer2_outputs(6882));
    layer3_outputs(988) <= layer2_outputs(2507);
    layer3_outputs(989) <= not(layer2_outputs(3164));
    layer3_outputs(990) <= (layer2_outputs(5574)) or (layer2_outputs(54));
    layer3_outputs(991) <= not(layer2_outputs(2769));
    layer3_outputs(992) <= layer2_outputs(745);
    layer3_outputs(993) <= (layer2_outputs(2480)) and not (layer2_outputs(989));
    layer3_outputs(994) <= (layer2_outputs(2502)) and not (layer2_outputs(1184));
    layer3_outputs(995) <= not(layer2_outputs(6411));
    layer3_outputs(996) <= not((layer2_outputs(4511)) and (layer2_outputs(5272)));
    layer3_outputs(997) <= (layer2_outputs(5657)) and (layer2_outputs(2639));
    layer3_outputs(998) <= layer2_outputs(896);
    layer3_outputs(999) <= layer2_outputs(800);
    layer3_outputs(1000) <= (layer2_outputs(7056)) and not (layer2_outputs(5289));
    layer3_outputs(1001) <= not(layer2_outputs(4501));
    layer3_outputs(1002) <= not((layer2_outputs(709)) xor (layer2_outputs(2305)));
    layer3_outputs(1003) <= not((layer2_outputs(2372)) or (layer2_outputs(4279)));
    layer3_outputs(1004) <= (layer2_outputs(828)) and not (layer2_outputs(311));
    layer3_outputs(1005) <= not(layer2_outputs(3028));
    layer3_outputs(1006) <= not((layer2_outputs(2283)) and (layer2_outputs(1607)));
    layer3_outputs(1007) <= layer2_outputs(112);
    layer3_outputs(1008) <= '0';
    layer3_outputs(1009) <= not(layer2_outputs(4135));
    layer3_outputs(1010) <= layer2_outputs(5442);
    layer3_outputs(1011) <= not(layer2_outputs(853)) or (layer2_outputs(7476));
    layer3_outputs(1012) <= (layer2_outputs(1657)) and not (layer2_outputs(7291));
    layer3_outputs(1013) <= not(layer2_outputs(5861)) or (layer2_outputs(2026));
    layer3_outputs(1014) <= not(layer2_outputs(3863)) or (layer2_outputs(5008));
    layer3_outputs(1015) <= not(layer2_outputs(1975));
    layer3_outputs(1016) <= layer2_outputs(229);
    layer3_outputs(1017) <= (layer2_outputs(6202)) and not (layer2_outputs(7122));
    layer3_outputs(1018) <= (layer2_outputs(5509)) or (layer2_outputs(3737));
    layer3_outputs(1019) <= not(layer2_outputs(3660));
    layer3_outputs(1020) <= not(layer2_outputs(6283));
    layer3_outputs(1021) <= (layer2_outputs(7240)) or (layer2_outputs(5277));
    layer3_outputs(1022) <= layer2_outputs(2395);
    layer3_outputs(1023) <= not(layer2_outputs(1373));
    layer3_outputs(1024) <= '1';
    layer3_outputs(1025) <= not(layer2_outputs(5674));
    layer3_outputs(1026) <= not(layer2_outputs(2469)) or (layer2_outputs(4000));
    layer3_outputs(1027) <= (layer2_outputs(2783)) and not (layer2_outputs(3594));
    layer3_outputs(1028) <= layer2_outputs(532);
    layer3_outputs(1029) <= not(layer2_outputs(7341));
    layer3_outputs(1030) <= (layer2_outputs(4540)) and not (layer2_outputs(6017));
    layer3_outputs(1031) <= layer2_outputs(1544);
    layer3_outputs(1032) <= not(layer2_outputs(3855));
    layer3_outputs(1033) <= not(layer2_outputs(1467));
    layer3_outputs(1034) <= layer2_outputs(2632);
    layer3_outputs(1035) <= not(layer2_outputs(6961));
    layer3_outputs(1036) <= layer2_outputs(1536);
    layer3_outputs(1037) <= layer2_outputs(539);
    layer3_outputs(1038) <= '0';
    layer3_outputs(1039) <= not((layer2_outputs(4612)) or (layer2_outputs(1462)));
    layer3_outputs(1040) <= not((layer2_outputs(6456)) and (layer2_outputs(3530)));
    layer3_outputs(1041) <= (layer2_outputs(5840)) and not (layer2_outputs(3983));
    layer3_outputs(1042) <= not(layer2_outputs(5646));
    layer3_outputs(1043) <= not((layer2_outputs(2592)) or (layer2_outputs(5104)));
    layer3_outputs(1044) <= not(layer2_outputs(7548)) or (layer2_outputs(7031));
    layer3_outputs(1045) <= not((layer2_outputs(5390)) and (layer2_outputs(7655)));
    layer3_outputs(1046) <= not(layer2_outputs(4097));
    layer3_outputs(1047) <= not(layer2_outputs(7650));
    layer3_outputs(1048) <= not(layer2_outputs(1145));
    layer3_outputs(1049) <= not(layer2_outputs(187));
    layer3_outputs(1050) <= layer2_outputs(69);
    layer3_outputs(1051) <= not(layer2_outputs(4707));
    layer3_outputs(1052) <= (layer2_outputs(2756)) or (layer2_outputs(7302));
    layer3_outputs(1053) <= (layer2_outputs(730)) and not (layer2_outputs(1453));
    layer3_outputs(1054) <= (layer2_outputs(2376)) and not (layer2_outputs(7358));
    layer3_outputs(1055) <= not((layer2_outputs(2127)) xor (layer2_outputs(1678)));
    layer3_outputs(1056) <= not((layer2_outputs(838)) or (layer2_outputs(7617)));
    layer3_outputs(1057) <= layer2_outputs(3897);
    layer3_outputs(1058) <= not(layer2_outputs(6996)) or (layer2_outputs(1724));
    layer3_outputs(1059) <= not(layer2_outputs(67));
    layer3_outputs(1060) <= (layer2_outputs(7074)) xor (layer2_outputs(6986));
    layer3_outputs(1061) <= not(layer2_outputs(1389));
    layer3_outputs(1062) <= not(layer2_outputs(4525)) or (layer2_outputs(2682));
    layer3_outputs(1063) <= not(layer2_outputs(2277)) or (layer2_outputs(805));
    layer3_outputs(1064) <= not(layer2_outputs(4052)) or (layer2_outputs(7480));
    layer3_outputs(1065) <= layer2_outputs(5278);
    layer3_outputs(1066) <= not((layer2_outputs(792)) and (layer2_outputs(5680)));
    layer3_outputs(1067) <= (layer2_outputs(3945)) and (layer2_outputs(4240));
    layer3_outputs(1068) <= not(layer2_outputs(4441));
    layer3_outputs(1069) <= (layer2_outputs(545)) and not (layer2_outputs(384));
    layer3_outputs(1070) <= (layer2_outputs(48)) or (layer2_outputs(770));
    layer3_outputs(1071) <= (layer2_outputs(4393)) xor (layer2_outputs(5503));
    layer3_outputs(1072) <= not((layer2_outputs(2243)) and (layer2_outputs(4994)));
    layer3_outputs(1073) <= not(layer2_outputs(2378));
    layer3_outputs(1074) <= layer2_outputs(1680);
    layer3_outputs(1075) <= not(layer2_outputs(3743));
    layer3_outputs(1076) <= (layer2_outputs(1885)) or (layer2_outputs(5508));
    layer3_outputs(1077) <= not((layer2_outputs(6536)) or (layer2_outputs(1046)));
    layer3_outputs(1078) <= not(layer2_outputs(3126));
    layer3_outputs(1079) <= not((layer2_outputs(1912)) and (layer2_outputs(892)));
    layer3_outputs(1080) <= layer2_outputs(1009);
    layer3_outputs(1081) <= layer2_outputs(2786);
    layer3_outputs(1082) <= not(layer2_outputs(2743)) or (layer2_outputs(924));
    layer3_outputs(1083) <= (layer2_outputs(737)) and (layer2_outputs(7505));
    layer3_outputs(1084) <= not(layer2_outputs(3554));
    layer3_outputs(1085) <= (layer2_outputs(6473)) and not (layer2_outputs(4870));
    layer3_outputs(1086) <= not(layer2_outputs(3140));
    layer3_outputs(1087) <= not((layer2_outputs(4788)) xor (layer2_outputs(2627)));
    layer3_outputs(1088) <= not(layer2_outputs(3802));
    layer3_outputs(1089) <= (layer2_outputs(7435)) and not (layer2_outputs(1533));
    layer3_outputs(1090) <= not(layer2_outputs(3466)) or (layer2_outputs(2515));
    layer3_outputs(1091) <= (layer2_outputs(3493)) and (layer2_outputs(2937));
    layer3_outputs(1092) <= not(layer2_outputs(1549));
    layer3_outputs(1093) <= not(layer2_outputs(6965)) or (layer2_outputs(3259));
    layer3_outputs(1094) <= not(layer2_outputs(5192));
    layer3_outputs(1095) <= not(layer2_outputs(276));
    layer3_outputs(1096) <= layer2_outputs(4842);
    layer3_outputs(1097) <= layer2_outputs(4045);
    layer3_outputs(1098) <= (layer2_outputs(7037)) and (layer2_outputs(1913));
    layer3_outputs(1099) <= not(layer2_outputs(4676));
    layer3_outputs(1100) <= (layer2_outputs(4359)) and not (layer2_outputs(317));
    layer3_outputs(1101) <= layer2_outputs(1645);
    layer3_outputs(1102) <= not(layer2_outputs(3460));
    layer3_outputs(1103) <= layer2_outputs(2696);
    layer3_outputs(1104) <= (layer2_outputs(5678)) and not (layer2_outputs(6011));
    layer3_outputs(1105) <= layer2_outputs(3457);
    layer3_outputs(1106) <= layer2_outputs(2894);
    layer3_outputs(1107) <= (layer2_outputs(7022)) and not (layer2_outputs(4244));
    layer3_outputs(1108) <= (layer2_outputs(2881)) and (layer2_outputs(5595));
    layer3_outputs(1109) <= layer2_outputs(7551);
    layer3_outputs(1110) <= (layer2_outputs(3297)) and not (layer2_outputs(2784));
    layer3_outputs(1111) <= layer2_outputs(1433);
    layer3_outputs(1112) <= '0';
    layer3_outputs(1113) <= layer2_outputs(2974);
    layer3_outputs(1114) <= not(layer2_outputs(4235)) or (layer2_outputs(1568));
    layer3_outputs(1115) <= (layer2_outputs(1623)) or (layer2_outputs(2726));
    layer3_outputs(1116) <= '0';
    layer3_outputs(1117) <= not(layer2_outputs(2477)) or (layer2_outputs(6595));
    layer3_outputs(1118) <= layer2_outputs(4778);
    layer3_outputs(1119) <= '1';
    layer3_outputs(1120) <= not(layer2_outputs(2957));
    layer3_outputs(1121) <= not(layer2_outputs(1517));
    layer3_outputs(1122) <= not(layer2_outputs(2222)) or (layer2_outputs(6062));
    layer3_outputs(1123) <= not(layer2_outputs(2778));
    layer3_outputs(1124) <= not((layer2_outputs(2859)) xor (layer2_outputs(5656)));
    layer3_outputs(1125) <= layer2_outputs(3524);
    layer3_outputs(1126) <= not(layer2_outputs(4507));
    layer3_outputs(1127) <= not(layer2_outputs(6903));
    layer3_outputs(1128) <= (layer2_outputs(4106)) and (layer2_outputs(5492));
    layer3_outputs(1129) <= not(layer2_outputs(4764));
    layer3_outputs(1130) <= not(layer2_outputs(6209));
    layer3_outputs(1131) <= layer2_outputs(6750);
    layer3_outputs(1132) <= not((layer2_outputs(6305)) xor (layer2_outputs(4856)));
    layer3_outputs(1133) <= not(layer2_outputs(4358)) or (layer2_outputs(1621));
    layer3_outputs(1134) <= layer2_outputs(572);
    layer3_outputs(1135) <= not((layer2_outputs(2180)) or (layer2_outputs(2557)));
    layer3_outputs(1136) <= '0';
    layer3_outputs(1137) <= not(layer2_outputs(6307));
    layer3_outputs(1138) <= (layer2_outputs(5720)) and not (layer2_outputs(2285));
    layer3_outputs(1139) <= layer2_outputs(5688);
    layer3_outputs(1140) <= not((layer2_outputs(7074)) and (layer2_outputs(5784)));
    layer3_outputs(1141) <= not(layer2_outputs(4666));
    layer3_outputs(1142) <= layer2_outputs(875);
    layer3_outputs(1143) <= layer2_outputs(4530);
    layer3_outputs(1144) <= '0';
    layer3_outputs(1145) <= (layer2_outputs(3427)) xor (layer2_outputs(4989));
    layer3_outputs(1146) <= (layer2_outputs(7441)) and not (layer2_outputs(3920));
    layer3_outputs(1147) <= not(layer2_outputs(6326)) or (layer2_outputs(7209));
    layer3_outputs(1148) <= not((layer2_outputs(3543)) and (layer2_outputs(6418)));
    layer3_outputs(1149) <= layer2_outputs(6416);
    layer3_outputs(1150) <= not(layer2_outputs(1791)) or (layer2_outputs(1018));
    layer3_outputs(1151) <= not(layer2_outputs(2010));
    layer3_outputs(1152) <= (layer2_outputs(4345)) or (layer2_outputs(1293));
    layer3_outputs(1153) <= not((layer2_outputs(1)) or (layer2_outputs(6095)));
    layer3_outputs(1154) <= not(layer2_outputs(7211));
    layer3_outputs(1155) <= layer2_outputs(7136);
    layer3_outputs(1156) <= not(layer2_outputs(6941)) or (layer2_outputs(4335));
    layer3_outputs(1157) <= not(layer2_outputs(7648));
    layer3_outputs(1158) <= (layer2_outputs(2251)) and not (layer2_outputs(6335));
    layer3_outputs(1159) <= not(layer2_outputs(5722));
    layer3_outputs(1160) <= not(layer2_outputs(4653)) or (layer2_outputs(7385));
    layer3_outputs(1161) <= not((layer2_outputs(1498)) and (layer2_outputs(340)));
    layer3_outputs(1162) <= (layer2_outputs(7655)) and not (layer2_outputs(4995));
    layer3_outputs(1163) <= not(layer2_outputs(3352)) or (layer2_outputs(3185));
    layer3_outputs(1164) <= not(layer2_outputs(4795));
    layer3_outputs(1165) <= not(layer2_outputs(4452));
    layer3_outputs(1166) <= not(layer2_outputs(2818)) or (layer2_outputs(4772));
    layer3_outputs(1167) <= (layer2_outputs(5413)) xor (layer2_outputs(4170));
    layer3_outputs(1168) <= layer2_outputs(1031);
    layer3_outputs(1169) <= (layer2_outputs(2400)) or (layer2_outputs(5147));
    layer3_outputs(1170) <= not(layer2_outputs(687));
    layer3_outputs(1171) <= layer2_outputs(1);
    layer3_outputs(1172) <= '0';
    layer3_outputs(1173) <= not(layer2_outputs(396));
    layer3_outputs(1174) <= not((layer2_outputs(2785)) and (layer2_outputs(7080)));
    layer3_outputs(1175) <= not((layer2_outputs(4709)) or (layer2_outputs(5701)));
    layer3_outputs(1176) <= layer2_outputs(2117);
    layer3_outputs(1177) <= (layer2_outputs(4800)) or (layer2_outputs(3493));
    layer3_outputs(1178) <= (layer2_outputs(5890)) and (layer2_outputs(3840));
    layer3_outputs(1179) <= not(layer2_outputs(5400));
    layer3_outputs(1180) <= not(layer2_outputs(4062)) or (layer2_outputs(4790));
    layer3_outputs(1181) <= '1';
    layer3_outputs(1182) <= layer2_outputs(150);
    layer3_outputs(1183) <= not((layer2_outputs(4978)) and (layer2_outputs(2290)));
    layer3_outputs(1184) <= (layer2_outputs(2721)) and (layer2_outputs(3234));
    layer3_outputs(1185) <= not(layer2_outputs(4711));
    layer3_outputs(1186) <= not(layer2_outputs(6159)) or (layer2_outputs(3868));
    layer3_outputs(1187) <= not(layer2_outputs(6004));
    layer3_outputs(1188) <= layer2_outputs(7641);
    layer3_outputs(1189) <= layer2_outputs(4728);
    layer3_outputs(1190) <= not(layer2_outputs(2847));
    layer3_outputs(1191) <= not((layer2_outputs(7154)) and (layer2_outputs(1737)));
    layer3_outputs(1192) <= (layer2_outputs(2824)) and not (layer2_outputs(1283));
    layer3_outputs(1193) <= layer2_outputs(3627);
    layer3_outputs(1194) <= not(layer2_outputs(6379)) or (layer2_outputs(1849));
    layer3_outputs(1195) <= not(layer2_outputs(2959));
    layer3_outputs(1196) <= '1';
    layer3_outputs(1197) <= (layer2_outputs(4716)) and not (layer2_outputs(2697));
    layer3_outputs(1198) <= layer2_outputs(6698);
    layer3_outputs(1199) <= not(layer2_outputs(3596)) or (layer2_outputs(7294));
    layer3_outputs(1200) <= not((layer2_outputs(3662)) xor (layer2_outputs(679)));
    layer3_outputs(1201) <= not(layer2_outputs(5312)) or (layer2_outputs(5238));
    layer3_outputs(1202) <= not(layer2_outputs(5179));
    layer3_outputs(1203) <= (layer2_outputs(6707)) or (layer2_outputs(7138));
    layer3_outputs(1204) <= not((layer2_outputs(6709)) and (layer2_outputs(6)));
    layer3_outputs(1205) <= not(layer2_outputs(2685));
    layer3_outputs(1206) <= not(layer2_outputs(6101));
    layer3_outputs(1207) <= not((layer2_outputs(5806)) xor (layer2_outputs(1147)));
    layer3_outputs(1208) <= layer2_outputs(6324);
    layer3_outputs(1209) <= (layer2_outputs(5494)) and (layer2_outputs(835));
    layer3_outputs(1210) <= not(layer2_outputs(5036));
    layer3_outputs(1211) <= not(layer2_outputs(3515));
    layer3_outputs(1212) <= not(layer2_outputs(1158));
    layer3_outputs(1213) <= layer2_outputs(7251);
    layer3_outputs(1214) <= layer2_outputs(5906);
    layer3_outputs(1215) <= not(layer2_outputs(4095));
    layer3_outputs(1216) <= not((layer2_outputs(6434)) xor (layer2_outputs(4261)));
    layer3_outputs(1217) <= not(layer2_outputs(2047));
    layer3_outputs(1218) <= layer2_outputs(3034);
    layer3_outputs(1219) <= not((layer2_outputs(2895)) or (layer2_outputs(587)));
    layer3_outputs(1220) <= not(layer2_outputs(392));
    layer3_outputs(1221) <= layer2_outputs(49);
    layer3_outputs(1222) <= not(layer2_outputs(7541));
    layer3_outputs(1223) <= '1';
    layer3_outputs(1224) <= (layer2_outputs(6080)) and not (layer2_outputs(7191));
    layer3_outputs(1225) <= not((layer2_outputs(1061)) and (layer2_outputs(1507)));
    layer3_outputs(1226) <= (layer2_outputs(4684)) and not (layer2_outputs(39));
    layer3_outputs(1227) <= (layer2_outputs(4245)) and not (layer2_outputs(2815));
    layer3_outputs(1228) <= (layer2_outputs(1034)) xor (layer2_outputs(6729));
    layer3_outputs(1229) <= (layer2_outputs(1486)) or (layer2_outputs(1548));
    layer3_outputs(1230) <= '0';
    layer3_outputs(1231) <= not(layer2_outputs(2572));
    layer3_outputs(1232) <= layer2_outputs(4637);
    layer3_outputs(1233) <= (layer2_outputs(5081)) and (layer2_outputs(3220));
    layer3_outputs(1234) <= not((layer2_outputs(1861)) and (layer2_outputs(2059)));
    layer3_outputs(1235) <= not(layer2_outputs(632));
    layer3_outputs(1236) <= '0';
    layer3_outputs(1237) <= not(layer2_outputs(4835));
    layer3_outputs(1238) <= not((layer2_outputs(428)) and (layer2_outputs(1831)));
    layer3_outputs(1239) <= (layer2_outputs(4012)) and (layer2_outputs(6868));
    layer3_outputs(1240) <= layer2_outputs(5683);
    layer3_outputs(1241) <= not(layer2_outputs(2149));
    layer3_outputs(1242) <= not(layer2_outputs(1463));
    layer3_outputs(1243) <= not(layer2_outputs(344));
    layer3_outputs(1244) <= not(layer2_outputs(1767));
    layer3_outputs(1245) <= (layer2_outputs(1240)) or (layer2_outputs(7296));
    layer3_outputs(1246) <= (layer2_outputs(5571)) and not (layer2_outputs(7100));
    layer3_outputs(1247) <= (layer2_outputs(1055)) and not (layer2_outputs(3303));
    layer3_outputs(1248) <= layer2_outputs(3208);
    layer3_outputs(1249) <= (layer2_outputs(6142)) and (layer2_outputs(6877));
    layer3_outputs(1250) <= (layer2_outputs(3616)) and not (layer2_outputs(2988));
    layer3_outputs(1251) <= not(layer2_outputs(2099));
    layer3_outputs(1252) <= (layer2_outputs(1085)) and not (layer2_outputs(127));
    layer3_outputs(1253) <= not((layer2_outputs(2315)) xor (layer2_outputs(3932)));
    layer3_outputs(1254) <= (layer2_outputs(1774)) and not (layer2_outputs(6704));
    layer3_outputs(1255) <= layer2_outputs(2409);
    layer3_outputs(1256) <= layer2_outputs(1762);
    layer3_outputs(1257) <= (layer2_outputs(1822)) xor (layer2_outputs(2314));
    layer3_outputs(1258) <= (layer2_outputs(7616)) xor (layer2_outputs(4029));
    layer3_outputs(1259) <= not(layer2_outputs(1716));
    layer3_outputs(1260) <= not(layer2_outputs(3245));
    layer3_outputs(1261) <= not((layer2_outputs(2523)) xor (layer2_outputs(3252)));
    layer3_outputs(1262) <= not(layer2_outputs(3583)) or (layer2_outputs(5843));
    layer3_outputs(1263) <= not(layer2_outputs(4686));
    layer3_outputs(1264) <= not(layer2_outputs(5773)) or (layer2_outputs(808));
    layer3_outputs(1265) <= layer2_outputs(4372);
    layer3_outputs(1266) <= not(layer2_outputs(2553));
    layer3_outputs(1267) <= layer2_outputs(4283);
    layer3_outputs(1268) <= not(layer2_outputs(4962));
    layer3_outputs(1269) <= layer2_outputs(3081);
    layer3_outputs(1270) <= not(layer2_outputs(3378)) or (layer2_outputs(3907));
    layer3_outputs(1271) <= not((layer2_outputs(6929)) or (layer2_outputs(7200)));
    layer3_outputs(1272) <= (layer2_outputs(2116)) xor (layer2_outputs(4525));
    layer3_outputs(1273) <= not(layer2_outputs(1132));
    layer3_outputs(1274) <= layer2_outputs(2227);
    layer3_outputs(1275) <= layer2_outputs(4798);
    layer3_outputs(1276) <= (layer2_outputs(4435)) xor (layer2_outputs(6474));
    layer3_outputs(1277) <= (layer2_outputs(4102)) and (layer2_outputs(3105));
    layer3_outputs(1278) <= (layer2_outputs(162)) and not (layer2_outputs(2438));
    layer3_outputs(1279) <= not(layer2_outputs(1134)) or (layer2_outputs(6151));
    layer3_outputs(1280) <= not(layer2_outputs(4531)) or (layer2_outputs(1565));
    layer3_outputs(1281) <= not((layer2_outputs(4440)) and (layer2_outputs(4320)));
    layer3_outputs(1282) <= not(layer2_outputs(7283)) or (layer2_outputs(4376));
    layer3_outputs(1283) <= not(layer2_outputs(4559));
    layer3_outputs(1284) <= not(layer2_outputs(3878)) or (layer2_outputs(2204));
    layer3_outputs(1285) <= (layer2_outputs(3253)) or (layer2_outputs(2948));
    layer3_outputs(1286) <= (layer2_outputs(6282)) xor (layer2_outputs(2248));
    layer3_outputs(1287) <= not((layer2_outputs(5113)) and (layer2_outputs(4627)));
    layer3_outputs(1288) <= not(layer2_outputs(1664));
    layer3_outputs(1289) <= layer2_outputs(5268);
    layer3_outputs(1290) <= not(layer2_outputs(408)) or (layer2_outputs(597));
    layer3_outputs(1291) <= (layer2_outputs(4750)) and (layer2_outputs(4036));
    layer3_outputs(1292) <= not((layer2_outputs(2073)) or (layer2_outputs(7429)));
    layer3_outputs(1293) <= layer2_outputs(5896);
    layer3_outputs(1294) <= '0';
    layer3_outputs(1295) <= layer2_outputs(2882);
    layer3_outputs(1296) <= '0';
    layer3_outputs(1297) <= layer2_outputs(4041);
    layer3_outputs(1298) <= not(layer2_outputs(6015)) or (layer2_outputs(5436));
    layer3_outputs(1299) <= layer2_outputs(6413);
    layer3_outputs(1300) <= not(layer2_outputs(4443));
    layer3_outputs(1301) <= not(layer2_outputs(3376)) or (layer2_outputs(3831));
    layer3_outputs(1302) <= layer2_outputs(4925);
    layer3_outputs(1303) <= not((layer2_outputs(4212)) and (layer2_outputs(5759)));
    layer3_outputs(1304) <= '1';
    layer3_outputs(1305) <= (layer2_outputs(4791)) and not (layer2_outputs(440));
    layer3_outputs(1306) <= not(layer2_outputs(6406));
    layer3_outputs(1307) <= (layer2_outputs(7172)) and not (layer2_outputs(2433));
    layer3_outputs(1308) <= not((layer2_outputs(5059)) xor (layer2_outputs(6767)));
    layer3_outputs(1309) <= not((layer2_outputs(3424)) and (layer2_outputs(3318)));
    layer3_outputs(1310) <= not(layer2_outputs(6186)) or (layer2_outputs(5743));
    layer3_outputs(1311) <= (layer2_outputs(553)) and not (layer2_outputs(2763));
    layer3_outputs(1312) <= not(layer2_outputs(1165));
    layer3_outputs(1313) <= not(layer2_outputs(592));
    layer3_outputs(1314) <= not(layer2_outputs(4932));
    layer3_outputs(1315) <= not(layer2_outputs(5735));
    layer3_outputs(1316) <= '0';
    layer3_outputs(1317) <= not(layer2_outputs(2044));
    layer3_outputs(1318) <= not(layer2_outputs(6613));
    layer3_outputs(1319) <= (layer2_outputs(1422)) or (layer2_outputs(7507));
    layer3_outputs(1320) <= '1';
    layer3_outputs(1321) <= layer2_outputs(3444);
    layer3_outputs(1322) <= '1';
    layer3_outputs(1323) <= not(layer2_outputs(1194)) or (layer2_outputs(4699));
    layer3_outputs(1324) <= layer2_outputs(688);
    layer3_outputs(1325) <= not(layer2_outputs(5653)) or (layer2_outputs(4259));
    layer3_outputs(1326) <= not(layer2_outputs(4031));
    layer3_outputs(1327) <= not(layer2_outputs(6069));
    layer3_outputs(1328) <= not(layer2_outputs(6198));
    layer3_outputs(1329) <= (layer2_outputs(4777)) or (layer2_outputs(251));
    layer3_outputs(1330) <= (layer2_outputs(3346)) and not (layer2_outputs(3479));
    layer3_outputs(1331) <= not(layer2_outputs(3363));
    layer3_outputs(1332) <= (layer2_outputs(6888)) and not (layer2_outputs(2521));
    layer3_outputs(1333) <= (layer2_outputs(1311)) and not (layer2_outputs(6455));
    layer3_outputs(1334) <= not(layer2_outputs(1012));
    layer3_outputs(1335) <= layer2_outputs(6836);
    layer3_outputs(1336) <= layer2_outputs(4702);
    layer3_outputs(1337) <= not(layer2_outputs(7676));
    layer3_outputs(1338) <= (layer2_outputs(1026)) xor (layer2_outputs(4469));
    layer3_outputs(1339) <= not(layer2_outputs(3330));
    layer3_outputs(1340) <= not(layer2_outputs(238));
    layer3_outputs(1341) <= not((layer2_outputs(4201)) and (layer2_outputs(3850)));
    layer3_outputs(1342) <= (layer2_outputs(4203)) xor (layer2_outputs(3329));
    layer3_outputs(1343) <= not(layer2_outputs(6146));
    layer3_outputs(1344) <= not(layer2_outputs(4438)) or (layer2_outputs(3985));
    layer3_outputs(1345) <= (layer2_outputs(7277)) xor (layer2_outputs(4143));
    layer3_outputs(1346) <= (layer2_outputs(6271)) and (layer2_outputs(5271));
    layer3_outputs(1347) <= not((layer2_outputs(5204)) xor (layer2_outputs(5001)));
    layer3_outputs(1348) <= (layer2_outputs(2542)) or (layer2_outputs(5532));
    layer3_outputs(1349) <= not((layer2_outputs(2891)) or (layer2_outputs(2237)));
    layer3_outputs(1350) <= (layer2_outputs(5850)) and not (layer2_outputs(5895));
    layer3_outputs(1351) <= not(layer2_outputs(1381)) or (layer2_outputs(4363));
    layer3_outputs(1352) <= (layer2_outputs(5742)) or (layer2_outputs(2256));
    layer3_outputs(1353) <= layer2_outputs(4733);
    layer3_outputs(1354) <= layer2_outputs(2687);
    layer3_outputs(1355) <= not(layer2_outputs(1987));
    layer3_outputs(1356) <= not(layer2_outputs(2340)) or (layer2_outputs(89));
    layer3_outputs(1357) <= not(layer2_outputs(5437));
    layer3_outputs(1358) <= not((layer2_outputs(4555)) or (layer2_outputs(6007)));
    layer3_outputs(1359) <= not(layer2_outputs(200)) or (layer2_outputs(6405));
    layer3_outputs(1360) <= (layer2_outputs(4765)) and (layer2_outputs(7300));
    layer3_outputs(1361) <= not(layer2_outputs(4738));
    layer3_outputs(1362) <= (layer2_outputs(5214)) and not (layer2_outputs(7284));
    layer3_outputs(1363) <= not(layer2_outputs(320)) or (layer2_outputs(3528));
    layer3_outputs(1364) <= layer2_outputs(6699);
    layer3_outputs(1365) <= not(layer2_outputs(6308));
    layer3_outputs(1366) <= not((layer2_outputs(3138)) xor (layer2_outputs(1840)));
    layer3_outputs(1367) <= not(layer2_outputs(1372));
    layer3_outputs(1368) <= '0';
    layer3_outputs(1369) <= layer2_outputs(5368);
    layer3_outputs(1370) <= layer2_outputs(5011);
    layer3_outputs(1371) <= layer2_outputs(7532);
    layer3_outputs(1372) <= not(layer2_outputs(4165)) or (layer2_outputs(638));
    layer3_outputs(1373) <= '0';
    layer3_outputs(1374) <= (layer2_outputs(3242)) and not (layer2_outputs(2049));
    layer3_outputs(1375) <= not((layer2_outputs(285)) or (layer2_outputs(7555)));
    layer3_outputs(1376) <= layer2_outputs(350);
    layer3_outputs(1377) <= not(layer2_outputs(7246));
    layer3_outputs(1378) <= layer2_outputs(6662);
    layer3_outputs(1379) <= '0';
    layer3_outputs(1380) <= not(layer2_outputs(2326));
    layer3_outputs(1381) <= not(layer2_outputs(1202));
    layer3_outputs(1382) <= not(layer2_outputs(3343));
    layer3_outputs(1383) <= not(layer2_outputs(1115)) or (layer2_outputs(4171));
    layer3_outputs(1384) <= not((layer2_outputs(5610)) or (layer2_outputs(5013)));
    layer3_outputs(1385) <= layer2_outputs(2820);
    layer3_outputs(1386) <= layer2_outputs(4485);
    layer3_outputs(1387) <= not(layer2_outputs(1800));
    layer3_outputs(1388) <= (layer2_outputs(4974)) and not (layer2_outputs(5041));
    layer3_outputs(1389) <= (layer2_outputs(7041)) and (layer2_outputs(6562));
    layer3_outputs(1390) <= not((layer2_outputs(6462)) and (layer2_outputs(5948)));
    layer3_outputs(1391) <= layer2_outputs(6026);
    layer3_outputs(1392) <= '0';
    layer3_outputs(1393) <= not(layer2_outputs(4610)) or (layer2_outputs(6125));
    layer3_outputs(1394) <= (layer2_outputs(7301)) and not (layer2_outputs(5660));
    layer3_outputs(1395) <= not(layer2_outputs(754));
    layer3_outputs(1396) <= not((layer2_outputs(5918)) xor (layer2_outputs(1444)));
    layer3_outputs(1397) <= not(layer2_outputs(2545)) or (layer2_outputs(6333));
    layer3_outputs(1398) <= not(layer2_outputs(7292));
    layer3_outputs(1399) <= not((layer2_outputs(258)) and (layer2_outputs(5240)));
    layer3_outputs(1400) <= layer2_outputs(2535);
    layer3_outputs(1401) <= (layer2_outputs(4283)) and not (layer2_outputs(914));
    layer3_outputs(1402) <= not((layer2_outputs(6292)) xor (layer2_outputs(2519)));
    layer3_outputs(1403) <= not(layer2_outputs(6667));
    layer3_outputs(1404) <= (layer2_outputs(4616)) or (layer2_outputs(7133));
    layer3_outputs(1405) <= not((layer2_outputs(3095)) or (layer2_outputs(1315)));
    layer3_outputs(1406) <= (layer2_outputs(2642)) or (layer2_outputs(3109));
    layer3_outputs(1407) <= not(layer2_outputs(555));
    layer3_outputs(1408) <= (layer2_outputs(3634)) and (layer2_outputs(7042));
    layer3_outputs(1409) <= '1';
    layer3_outputs(1410) <= layer2_outputs(5408);
    layer3_outputs(1411) <= not(layer2_outputs(1334));
    layer3_outputs(1412) <= layer2_outputs(5502);
    layer3_outputs(1413) <= not(layer2_outputs(5498));
    layer3_outputs(1414) <= '1';
    layer3_outputs(1415) <= not(layer2_outputs(2588));
    layer3_outputs(1416) <= not(layer2_outputs(6674));
    layer3_outputs(1417) <= not(layer2_outputs(3689)) or (layer2_outputs(7049));
    layer3_outputs(1418) <= layer2_outputs(5572);
    layer3_outputs(1419) <= (layer2_outputs(4735)) and (layer2_outputs(3056));
    layer3_outputs(1420) <= (layer2_outputs(6519)) and not (layer2_outputs(54));
    layer3_outputs(1421) <= (layer2_outputs(2674)) and not (layer2_outputs(5792));
    layer3_outputs(1422) <= layer2_outputs(892);
    layer3_outputs(1423) <= not((layer2_outputs(1947)) and (layer2_outputs(5287)));
    layer3_outputs(1424) <= not(layer2_outputs(187));
    layer3_outputs(1425) <= layer2_outputs(3446);
    layer3_outputs(1426) <= (layer2_outputs(189)) and not (layer2_outputs(3463));
    layer3_outputs(1427) <= layer2_outputs(224);
    layer3_outputs(1428) <= (layer2_outputs(5737)) and not (layer2_outputs(1093));
    layer3_outputs(1429) <= layer2_outputs(7101);
    layer3_outputs(1430) <= '0';
    layer3_outputs(1431) <= layer2_outputs(3307);
    layer3_outputs(1432) <= not((layer2_outputs(5381)) or (layer2_outputs(4505)));
    layer3_outputs(1433) <= not(layer2_outputs(173));
    layer3_outputs(1434) <= (layer2_outputs(5765)) or (layer2_outputs(2353));
    layer3_outputs(1435) <= not(layer2_outputs(4437));
    layer3_outputs(1436) <= not((layer2_outputs(2455)) or (layer2_outputs(7503)));
    layer3_outputs(1437) <= not(layer2_outputs(4736));
    layer3_outputs(1438) <= not(layer2_outputs(1970));
    layer3_outputs(1439) <= layer2_outputs(5340);
    layer3_outputs(1440) <= (layer2_outputs(2480)) and (layer2_outputs(7324));
    layer3_outputs(1441) <= layer2_outputs(4658);
    layer3_outputs(1442) <= not(layer2_outputs(5599));
    layer3_outputs(1443) <= not((layer2_outputs(2568)) xor (layer2_outputs(3404)));
    layer3_outputs(1444) <= not((layer2_outputs(5028)) and (layer2_outputs(6132)));
    layer3_outputs(1445) <= layer2_outputs(148);
    layer3_outputs(1446) <= not(layer2_outputs(3163)) or (layer2_outputs(4958));
    layer3_outputs(1447) <= (layer2_outputs(3671)) xor (layer2_outputs(2728));
    layer3_outputs(1448) <= not((layer2_outputs(3292)) xor (layer2_outputs(6066)));
    layer3_outputs(1449) <= (layer2_outputs(5622)) and (layer2_outputs(5971));
    layer3_outputs(1450) <= (layer2_outputs(3913)) or (layer2_outputs(5633));
    layer3_outputs(1451) <= (layer2_outputs(985)) and not (layer2_outputs(4199));
    layer3_outputs(1452) <= not((layer2_outputs(4434)) or (layer2_outputs(5633)));
    layer3_outputs(1453) <= not((layer2_outputs(4998)) and (layer2_outputs(623)));
    layer3_outputs(1454) <= (layer2_outputs(1277)) and not (layer2_outputs(5658));
    layer3_outputs(1455) <= layer2_outputs(6199);
    layer3_outputs(1456) <= not((layer2_outputs(1408)) or (layer2_outputs(1161)));
    layer3_outputs(1457) <= (layer2_outputs(6382)) xor (layer2_outputs(5185));
    layer3_outputs(1458) <= (layer2_outputs(7010)) and not (layer2_outputs(299));
    layer3_outputs(1459) <= not(layer2_outputs(3614));
    layer3_outputs(1460) <= layer2_outputs(6825);
    layer3_outputs(1461) <= layer2_outputs(5621);
    layer3_outputs(1462) <= (layer2_outputs(7529)) and not (layer2_outputs(641));
    layer3_outputs(1463) <= not(layer2_outputs(1234)) or (layer2_outputs(5290));
    layer3_outputs(1464) <= '1';
    layer3_outputs(1465) <= layer2_outputs(5704);
    layer3_outputs(1466) <= not((layer2_outputs(1080)) and (layer2_outputs(6137)));
    layer3_outputs(1467) <= (layer2_outputs(5348)) and not (layer2_outputs(1501));
    layer3_outputs(1468) <= (layer2_outputs(5659)) and not (layer2_outputs(5825));
    layer3_outputs(1469) <= layer2_outputs(7203);
    layer3_outputs(1470) <= '1';
    layer3_outputs(1471) <= not(layer2_outputs(1536));
    layer3_outputs(1472) <= not((layer2_outputs(2740)) or (layer2_outputs(1545)));
    layer3_outputs(1473) <= (layer2_outputs(1430)) and not (layer2_outputs(151));
    layer3_outputs(1474) <= layer2_outputs(2432);
    layer3_outputs(1475) <= (layer2_outputs(6677)) and not (layer2_outputs(4846));
    layer3_outputs(1476) <= not(layer2_outputs(7064));
    layer3_outputs(1477) <= not(layer2_outputs(6539));
    layer3_outputs(1478) <= not(layer2_outputs(7670));
    layer3_outputs(1479) <= layer2_outputs(390);
    layer3_outputs(1480) <= not(layer2_outputs(2857)) or (layer2_outputs(4747));
    layer3_outputs(1481) <= (layer2_outputs(7454)) xor (layer2_outputs(1278));
    layer3_outputs(1482) <= not(layer2_outputs(5083));
    layer3_outputs(1483) <= not((layer2_outputs(1883)) or (layer2_outputs(468)));
    layer3_outputs(1484) <= '0';
    layer3_outputs(1485) <= (layer2_outputs(1222)) or (layer2_outputs(3276));
    layer3_outputs(1486) <= '1';
    layer3_outputs(1487) <= (layer2_outputs(7148)) or (layer2_outputs(7312));
    layer3_outputs(1488) <= not(layer2_outputs(7103)) or (layer2_outputs(2956));
    layer3_outputs(1489) <= (layer2_outputs(265)) and not (layer2_outputs(7210));
    layer3_outputs(1490) <= not(layer2_outputs(5653));
    layer3_outputs(1491) <= layer2_outputs(1108);
    layer3_outputs(1492) <= not(layer2_outputs(4991));
    layer3_outputs(1493) <= (layer2_outputs(7306)) xor (layer2_outputs(6491));
    layer3_outputs(1494) <= (layer2_outputs(5584)) and (layer2_outputs(3465));
    layer3_outputs(1495) <= (layer2_outputs(4014)) and (layer2_outputs(6182));
    layer3_outputs(1496) <= not(layer2_outputs(660));
    layer3_outputs(1497) <= (layer2_outputs(6801)) and not (layer2_outputs(1865));
    layer3_outputs(1498) <= layer2_outputs(4316);
    layer3_outputs(1499) <= not((layer2_outputs(7047)) xor (layer2_outputs(7)));
    layer3_outputs(1500) <= not(layer2_outputs(5421));
    layer3_outputs(1501) <= layer2_outputs(5685);
    layer3_outputs(1502) <= layer2_outputs(269);
    layer3_outputs(1503) <= layer2_outputs(4581);
    layer3_outputs(1504) <= not(layer2_outputs(7224)) or (layer2_outputs(6627));
    layer3_outputs(1505) <= layer2_outputs(5721);
    layer3_outputs(1506) <= not(layer2_outputs(579));
    layer3_outputs(1507) <= layer2_outputs(3826);
    layer3_outputs(1508) <= layer2_outputs(1990);
    layer3_outputs(1509) <= layer2_outputs(3589);
    layer3_outputs(1510) <= layer2_outputs(2503);
    layer3_outputs(1511) <= not((layer2_outputs(6255)) or (layer2_outputs(4584)));
    layer3_outputs(1512) <= not(layer2_outputs(5690));
    layer3_outputs(1513) <= not(layer2_outputs(4715));
    layer3_outputs(1514) <= (layer2_outputs(2921)) or (layer2_outputs(6515));
    layer3_outputs(1515) <= layer2_outputs(4948);
    layer3_outputs(1516) <= layer2_outputs(5381);
    layer3_outputs(1517) <= layer2_outputs(1502);
    layer3_outputs(1518) <= layer2_outputs(637);
    layer3_outputs(1519) <= not((layer2_outputs(6035)) xor (layer2_outputs(1659)));
    layer3_outputs(1520) <= not(layer2_outputs(7518)) or (layer2_outputs(7440));
    layer3_outputs(1521) <= not(layer2_outputs(5949)) or (layer2_outputs(3545));
    layer3_outputs(1522) <= not((layer2_outputs(2223)) and (layer2_outputs(6476)));
    layer3_outputs(1523) <= not(layer2_outputs(6854));
    layer3_outputs(1524) <= (layer2_outputs(2486)) and not (layer2_outputs(1690));
    layer3_outputs(1525) <= not(layer2_outputs(2276));
    layer3_outputs(1526) <= not(layer2_outputs(6237));
    layer3_outputs(1527) <= not((layer2_outputs(6083)) or (layer2_outputs(4914)));
    layer3_outputs(1528) <= (layer2_outputs(2534)) and not (layer2_outputs(3905));
    layer3_outputs(1529) <= not((layer2_outputs(7040)) and (layer2_outputs(7488)));
    layer3_outputs(1530) <= (layer2_outputs(4887)) and not (layer2_outputs(2704));
    layer3_outputs(1531) <= layer2_outputs(3210);
    layer3_outputs(1532) <= (layer2_outputs(6188)) and (layer2_outputs(6652));
    layer3_outputs(1533) <= not((layer2_outputs(4434)) or (layer2_outputs(1575)));
    layer3_outputs(1534) <= not((layer2_outputs(4885)) or (layer2_outputs(4138)));
    layer3_outputs(1535) <= layer2_outputs(1302);
    layer3_outputs(1536) <= not(layer2_outputs(7124));
    layer3_outputs(1537) <= not((layer2_outputs(6598)) and (layer2_outputs(6678)));
    layer3_outputs(1538) <= layer2_outputs(7056);
    layer3_outputs(1539) <= (layer2_outputs(654)) and not (layer2_outputs(1942));
    layer3_outputs(1540) <= layer2_outputs(377);
    layer3_outputs(1541) <= not(layer2_outputs(6532));
    layer3_outputs(1542) <= not((layer2_outputs(6547)) or (layer2_outputs(2484)));
    layer3_outputs(1543) <= not(layer2_outputs(5234)) or (layer2_outputs(7157));
    layer3_outputs(1544) <= '1';
    layer3_outputs(1545) <= not(layer2_outputs(6138));
    layer3_outputs(1546) <= not(layer2_outputs(5112));
    layer3_outputs(1547) <= not(layer2_outputs(843));
    layer3_outputs(1548) <= not(layer2_outputs(5208));
    layer3_outputs(1549) <= not(layer2_outputs(2087));
    layer3_outputs(1550) <= not(layer2_outputs(5421));
    layer3_outputs(1551) <= (layer2_outputs(2131)) and (layer2_outputs(1559));
    layer3_outputs(1552) <= layer2_outputs(4237);
    layer3_outputs(1553) <= not(layer2_outputs(338));
    layer3_outputs(1554) <= (layer2_outputs(4710)) and not (layer2_outputs(6464));
    layer3_outputs(1555) <= '1';
    layer3_outputs(1556) <= layer2_outputs(4931);
    layer3_outputs(1557) <= (layer2_outputs(215)) and not (layer2_outputs(6668));
    layer3_outputs(1558) <= layer2_outputs(4137);
    layer3_outputs(1559) <= '1';
    layer3_outputs(1560) <= not(layer2_outputs(6072));
    layer3_outputs(1561) <= not(layer2_outputs(2132)) or (layer2_outputs(7159));
    layer3_outputs(1562) <= (layer2_outputs(2571)) and not (layer2_outputs(5320));
    layer3_outputs(1563) <= layer2_outputs(2909);
    layer3_outputs(1564) <= not(layer2_outputs(2857)) or (layer2_outputs(3557));
    layer3_outputs(1565) <= layer2_outputs(1045);
    layer3_outputs(1566) <= layer2_outputs(5143);
    layer3_outputs(1567) <= (layer2_outputs(1280)) and (layer2_outputs(970));
    layer3_outputs(1568) <= not(layer2_outputs(452)) or (layer2_outputs(7135));
    layer3_outputs(1569) <= (layer2_outputs(6367)) and not (layer2_outputs(1950));
    layer3_outputs(1570) <= (layer2_outputs(7030)) and not (layer2_outputs(7084));
    layer3_outputs(1571) <= (layer2_outputs(6567)) or (layer2_outputs(7009));
    layer3_outputs(1572) <= not(layer2_outputs(6097)) or (layer2_outputs(3461));
    layer3_outputs(1573) <= not(layer2_outputs(5760));
    layer3_outputs(1574) <= '0';
    layer3_outputs(1575) <= not((layer2_outputs(7630)) and (layer2_outputs(1800)));
    layer3_outputs(1576) <= layer2_outputs(7326);
    layer3_outputs(1577) <= (layer2_outputs(7573)) and not (layer2_outputs(7077));
    layer3_outputs(1578) <= not(layer2_outputs(7439));
    layer3_outputs(1579) <= layer2_outputs(6442);
    layer3_outputs(1580) <= (layer2_outputs(2038)) and not (layer2_outputs(5424));
    layer3_outputs(1581) <= not(layer2_outputs(1170));
    layer3_outputs(1582) <= (layer2_outputs(420)) and not (layer2_outputs(5474));
    layer3_outputs(1583) <= (layer2_outputs(3712)) and not (layer2_outputs(1558));
    layer3_outputs(1584) <= not(layer2_outputs(2777)) or (layer2_outputs(2359));
    layer3_outputs(1585) <= layer2_outputs(3648);
    layer3_outputs(1586) <= not(layer2_outputs(6186));
    layer3_outputs(1587) <= not(layer2_outputs(4490));
    layer3_outputs(1588) <= (layer2_outputs(1841)) xor (layer2_outputs(1199));
    layer3_outputs(1589) <= (layer2_outputs(1355)) or (layer2_outputs(4060));
    layer3_outputs(1590) <= not(layer2_outputs(5269));
    layer3_outputs(1591) <= not(layer2_outputs(1537));
    layer3_outputs(1592) <= not(layer2_outputs(4232));
    layer3_outputs(1593) <= not(layer2_outputs(4761));
    layer3_outputs(1594) <= not((layer2_outputs(2587)) and (layer2_outputs(7223)));
    layer3_outputs(1595) <= not(layer2_outputs(5848));
    layer3_outputs(1596) <= not(layer2_outputs(6043)) or (layer2_outputs(1853));
    layer3_outputs(1597) <= not(layer2_outputs(3079));
    layer3_outputs(1598) <= (layer2_outputs(1101)) or (layer2_outputs(6447));
    layer3_outputs(1599) <= layer2_outputs(5478);
    layer3_outputs(1600) <= not(layer2_outputs(7046));
    layer3_outputs(1601) <= not(layer2_outputs(4076));
    layer3_outputs(1602) <= '1';
    layer3_outputs(1603) <= not(layer2_outputs(3286)) or (layer2_outputs(5153));
    layer3_outputs(1604) <= not(layer2_outputs(3326)) or (layer2_outputs(4081));
    layer3_outputs(1605) <= (layer2_outputs(5450)) and (layer2_outputs(2585));
    layer3_outputs(1606) <= (layer2_outputs(6156)) xor (layer2_outputs(4811));
    layer3_outputs(1607) <= (layer2_outputs(3988)) or (layer2_outputs(2118));
    layer3_outputs(1608) <= not(layer2_outputs(7513));
    layer3_outputs(1609) <= (layer2_outputs(937)) and not (layer2_outputs(4964));
    layer3_outputs(1610) <= layer2_outputs(1627);
    layer3_outputs(1611) <= not(layer2_outputs(5715));
    layer3_outputs(1612) <= layer2_outputs(1763);
    layer3_outputs(1613) <= not(layer2_outputs(4161));
    layer3_outputs(1614) <= not(layer2_outputs(946)) or (layer2_outputs(1704));
    layer3_outputs(1615) <= not((layer2_outputs(3835)) and (layer2_outputs(5649)));
    layer3_outputs(1616) <= not(layer2_outputs(6514)) or (layer2_outputs(7320));
    layer3_outputs(1617) <= (layer2_outputs(6752)) and (layer2_outputs(544));
    layer3_outputs(1618) <= (layer2_outputs(5198)) and not (layer2_outputs(1453));
    layer3_outputs(1619) <= not((layer2_outputs(388)) and (layer2_outputs(3549)));
    layer3_outputs(1620) <= not(layer2_outputs(4058));
    layer3_outputs(1621) <= (layer2_outputs(6729)) and not (layer2_outputs(2350));
    layer3_outputs(1622) <= '0';
    layer3_outputs(1623) <= not(layer2_outputs(585));
    layer3_outputs(1624) <= (layer2_outputs(6892)) and not (layer2_outputs(2265));
    layer3_outputs(1625) <= layer2_outputs(2416);
    layer3_outputs(1626) <= not((layer2_outputs(6636)) or (layer2_outputs(4119)));
    layer3_outputs(1627) <= not(layer2_outputs(4780));
    layer3_outputs(1628) <= not(layer2_outputs(7669));
    layer3_outputs(1629) <= layer2_outputs(3189);
    layer3_outputs(1630) <= (layer2_outputs(2599)) and (layer2_outputs(6128));
    layer3_outputs(1631) <= not(layer2_outputs(2776));
    layer3_outputs(1632) <= '0';
    layer3_outputs(1633) <= not(layer2_outputs(943));
    layer3_outputs(1634) <= (layer2_outputs(2111)) and (layer2_outputs(2693));
    layer3_outputs(1635) <= layer2_outputs(5518);
    layer3_outputs(1636) <= '1';
    layer3_outputs(1637) <= (layer2_outputs(3940)) and not (layer2_outputs(1553));
    layer3_outputs(1638) <= not(layer2_outputs(7213));
    layer3_outputs(1639) <= (layer2_outputs(7431)) and not (layer2_outputs(4860));
    layer3_outputs(1640) <= not(layer2_outputs(1110));
    layer3_outputs(1641) <= (layer2_outputs(208)) or (layer2_outputs(4787));
    layer3_outputs(1642) <= (layer2_outputs(5893)) or (layer2_outputs(2306));
    layer3_outputs(1643) <= layer2_outputs(836);
    layer3_outputs(1644) <= layer2_outputs(24);
    layer3_outputs(1645) <= (layer2_outputs(5094)) and not (layer2_outputs(445));
    layer3_outputs(1646) <= layer2_outputs(4864);
    layer3_outputs(1647) <= layer2_outputs(2080);
    layer3_outputs(1648) <= layer2_outputs(6573);
    layer3_outputs(1649) <= layer2_outputs(5053);
    layer3_outputs(1650) <= not(layer2_outputs(4120)) or (layer2_outputs(2629));
    layer3_outputs(1651) <= (layer2_outputs(3178)) or (layer2_outputs(5750));
    layer3_outputs(1652) <= not(layer2_outputs(6351));
    layer3_outputs(1653) <= not(layer2_outputs(5179));
    layer3_outputs(1654) <= not((layer2_outputs(7241)) and (layer2_outputs(2165)));
    layer3_outputs(1655) <= not(layer2_outputs(2503));
    layer3_outputs(1656) <= layer2_outputs(6452);
    layer3_outputs(1657) <= layer2_outputs(1540);
    layer3_outputs(1658) <= not((layer2_outputs(2339)) and (layer2_outputs(2512)));
    layer3_outputs(1659) <= not(layer2_outputs(6957));
    layer3_outputs(1660) <= layer2_outputs(5936);
    layer3_outputs(1661) <= not(layer2_outputs(6931)) or (layer2_outputs(392));
    layer3_outputs(1662) <= not(layer2_outputs(2303)) or (layer2_outputs(4427));
    layer3_outputs(1663) <= not(layer2_outputs(4408)) or (layer2_outputs(7397));
    layer3_outputs(1664) <= layer2_outputs(5244);
    layer3_outputs(1665) <= not((layer2_outputs(6943)) or (layer2_outputs(5626)));
    layer3_outputs(1666) <= not(layer2_outputs(1351));
    layer3_outputs(1667) <= layer2_outputs(6901);
    layer3_outputs(1668) <= (layer2_outputs(5620)) and not (layer2_outputs(4275));
    layer3_outputs(1669) <= layer2_outputs(1285);
    layer3_outputs(1670) <= '0';
    layer3_outputs(1671) <= not(layer2_outputs(4720));
    layer3_outputs(1672) <= not(layer2_outputs(7522)) or (layer2_outputs(81));
    layer3_outputs(1673) <= '0';
    layer3_outputs(1674) <= not(layer2_outputs(7055));
    layer3_outputs(1675) <= layer2_outputs(2520);
    layer3_outputs(1676) <= not((layer2_outputs(7475)) or (layer2_outputs(4441)));
    layer3_outputs(1677) <= not(layer2_outputs(99)) or (layer2_outputs(6602));
    layer3_outputs(1678) <= not(layer2_outputs(4420));
    layer3_outputs(1679) <= not(layer2_outputs(877));
    layer3_outputs(1680) <= layer2_outputs(283);
    layer3_outputs(1681) <= not(layer2_outputs(7345)) or (layer2_outputs(2493));
    layer3_outputs(1682) <= not((layer2_outputs(3027)) xor (layer2_outputs(6120)));
    layer3_outputs(1683) <= layer2_outputs(2813);
    layer3_outputs(1684) <= not((layer2_outputs(4341)) or (layer2_outputs(6996)));
    layer3_outputs(1685) <= (layer2_outputs(4768)) or (layer2_outputs(3883));
    layer3_outputs(1686) <= not(layer2_outputs(6014));
    layer3_outputs(1687) <= (layer2_outputs(727)) and not (layer2_outputs(912));
    layer3_outputs(1688) <= not(layer2_outputs(1735)) or (layer2_outputs(5207));
    layer3_outputs(1689) <= not(layer2_outputs(5198));
    layer3_outputs(1690) <= layer2_outputs(6987);
    layer3_outputs(1691) <= not(layer2_outputs(7384)) or (layer2_outputs(7520));
    layer3_outputs(1692) <= not(layer2_outputs(5383));
    layer3_outputs(1693) <= layer2_outputs(1059);
    layer3_outputs(1694) <= (layer2_outputs(740)) or (layer2_outputs(169));
    layer3_outputs(1695) <= not((layer2_outputs(3802)) xor (layer2_outputs(1482)));
    layer3_outputs(1696) <= not((layer2_outputs(6191)) or (layer2_outputs(5193)));
    layer3_outputs(1697) <= '1';
    layer3_outputs(1698) <= layer2_outputs(6023);
    layer3_outputs(1699) <= not(layer2_outputs(2455));
    layer3_outputs(1700) <= layer2_outputs(4138);
    layer3_outputs(1701) <= (layer2_outputs(5625)) and (layer2_outputs(7361));
    layer3_outputs(1702) <= not(layer2_outputs(859)) or (layer2_outputs(2349));
    layer3_outputs(1703) <= (layer2_outputs(640)) and (layer2_outputs(3153));
    layer3_outputs(1704) <= not(layer2_outputs(451));
    layer3_outputs(1705) <= layer2_outputs(7188);
    layer3_outputs(1706) <= not((layer2_outputs(2496)) and (layer2_outputs(1088)));
    layer3_outputs(1707) <= layer2_outputs(3272);
    layer3_outputs(1708) <= '1';
    layer3_outputs(1709) <= not((layer2_outputs(2465)) xor (layer2_outputs(7033)));
    layer3_outputs(1710) <= (layer2_outputs(7529)) and not (layer2_outputs(3900));
    layer3_outputs(1711) <= not((layer2_outputs(1917)) xor (layer2_outputs(6959)));
    layer3_outputs(1712) <= (layer2_outputs(6518)) and not (layer2_outputs(4778));
    layer3_outputs(1713) <= layer2_outputs(2205);
    layer3_outputs(1714) <= not((layer2_outputs(4645)) and (layer2_outputs(4861)));
    layer3_outputs(1715) <= not(layer2_outputs(2294));
    layer3_outputs(1716) <= not(layer2_outputs(7227));
    layer3_outputs(1717) <= not((layer2_outputs(416)) xor (layer2_outputs(4876)));
    layer3_outputs(1718) <= layer2_outputs(779);
    layer3_outputs(1719) <= (layer2_outputs(4834)) and not (layer2_outputs(4827));
    layer3_outputs(1720) <= (layer2_outputs(2281)) and not (layer2_outputs(2741));
    layer3_outputs(1721) <= not((layer2_outputs(6947)) xor (layer2_outputs(3331)));
    layer3_outputs(1722) <= not(layer2_outputs(1884));
    layer3_outputs(1723) <= layer2_outputs(2004);
    layer3_outputs(1724) <= not(layer2_outputs(3132)) or (layer2_outputs(1272));
    layer3_outputs(1725) <= not(layer2_outputs(3302));
    layer3_outputs(1726) <= not((layer2_outputs(6829)) or (layer2_outputs(1619)));
    layer3_outputs(1727) <= not(layer2_outputs(3998)) or (layer2_outputs(3473));
    layer3_outputs(1728) <= '0';
    layer3_outputs(1729) <= not(layer2_outputs(1440)) or (layer2_outputs(2799));
    layer3_outputs(1730) <= not((layer2_outputs(6413)) xor (layer2_outputs(4428)));
    layer3_outputs(1731) <= not(layer2_outputs(3610));
    layer3_outputs(1732) <= not(layer2_outputs(6618));
    layer3_outputs(1733) <= layer2_outputs(3096);
    layer3_outputs(1734) <= not(layer2_outputs(5880));
    layer3_outputs(1735) <= (layer2_outputs(5784)) and (layer2_outputs(1130));
    layer3_outputs(1736) <= (layer2_outputs(4877)) xor (layer2_outputs(6137));
    layer3_outputs(1737) <= layer2_outputs(2929);
    layer3_outputs(1738) <= (layer2_outputs(4459)) and not (layer2_outputs(6155));
    layer3_outputs(1739) <= not(layer2_outputs(3719));
    layer3_outputs(1740) <= not(layer2_outputs(281));
    layer3_outputs(1741) <= layer2_outputs(6652);
    layer3_outputs(1742) <= layer2_outputs(6992);
    layer3_outputs(1743) <= (layer2_outputs(1738)) and (layer2_outputs(5380));
    layer3_outputs(1744) <= (layer2_outputs(2220)) and not (layer2_outputs(5042));
    layer3_outputs(1745) <= not(layer2_outputs(6626));
    layer3_outputs(1746) <= not(layer2_outputs(2445));
    layer3_outputs(1747) <= (layer2_outputs(4976)) and not (layer2_outputs(899));
    layer3_outputs(1748) <= layer2_outputs(5254);
    layer3_outputs(1749) <= (layer2_outputs(6916)) and not (layer2_outputs(2642));
    layer3_outputs(1750) <= layer2_outputs(809);
    layer3_outputs(1751) <= (layer2_outputs(1077)) and (layer2_outputs(7025));
    layer3_outputs(1752) <= (layer2_outputs(6252)) and not (layer2_outputs(3190));
    layer3_outputs(1753) <= not(layer2_outputs(3016));
    layer3_outputs(1754) <= not((layer2_outputs(3273)) or (layer2_outputs(4986)));
    layer3_outputs(1755) <= layer2_outputs(4313);
    layer3_outputs(1756) <= (layer2_outputs(1056)) or (layer2_outputs(1220));
    layer3_outputs(1757) <= not(layer2_outputs(3883));
    layer3_outputs(1758) <= '0';
    layer3_outputs(1759) <= not(layer2_outputs(3649)) or (layer2_outputs(7561));
    layer3_outputs(1760) <= (layer2_outputs(5599)) and (layer2_outputs(2949));
    layer3_outputs(1761) <= not(layer2_outputs(3302));
    layer3_outputs(1762) <= (layer2_outputs(5365)) and not (layer2_outputs(6375));
    layer3_outputs(1763) <= not(layer2_outputs(4991));
    layer3_outputs(1764) <= '0';
    layer3_outputs(1765) <= '0';
    layer3_outputs(1766) <= not(layer2_outputs(1926));
    layer3_outputs(1767) <= (layer2_outputs(1698)) and not (layer2_outputs(22));
    layer3_outputs(1768) <= not(layer2_outputs(1816));
    layer3_outputs(1769) <= not((layer2_outputs(312)) xor (layer2_outputs(2352)));
    layer3_outputs(1770) <= not(layer2_outputs(7569));
    layer3_outputs(1771) <= (layer2_outputs(3265)) and (layer2_outputs(7168));
    layer3_outputs(1772) <= (layer2_outputs(4583)) and not (layer2_outputs(4574));
    layer3_outputs(1773) <= (layer2_outputs(5425)) and not (layer2_outputs(826));
    layer3_outputs(1774) <= not(layer2_outputs(7406)) or (layer2_outputs(1793));
    layer3_outputs(1775) <= not(layer2_outputs(4863)) or (layer2_outputs(5354));
    layer3_outputs(1776) <= not(layer2_outputs(359));
    layer3_outputs(1777) <= (layer2_outputs(1916)) and not (layer2_outputs(3223));
    layer3_outputs(1778) <= layer2_outputs(2614);
    layer3_outputs(1779) <= not(layer2_outputs(2772));
    layer3_outputs(1780) <= layer2_outputs(6421);
    layer3_outputs(1781) <= layer2_outputs(3299);
    layer3_outputs(1782) <= not((layer2_outputs(2515)) or (layer2_outputs(1740)));
    layer3_outputs(1783) <= layer2_outputs(7076);
    layer3_outputs(1784) <= not((layer2_outputs(4274)) xor (layer2_outputs(6518)));
    layer3_outputs(1785) <= (layer2_outputs(3424)) or (layer2_outputs(1023));
    layer3_outputs(1786) <= not(layer2_outputs(3089));
    layer3_outputs(1787) <= not((layer2_outputs(4786)) xor (layer2_outputs(7546)));
    layer3_outputs(1788) <= not(layer2_outputs(6468));
    layer3_outputs(1789) <= (layer2_outputs(6973)) and not (layer2_outputs(5797));
    layer3_outputs(1790) <= not(layer2_outputs(1742));
    layer3_outputs(1791) <= layer2_outputs(673);
    layer3_outputs(1792) <= not(layer2_outputs(6312));
    layer3_outputs(1793) <= (layer2_outputs(2761)) or (layer2_outputs(4860));
    layer3_outputs(1794) <= (layer2_outputs(5122)) and (layer2_outputs(3182));
    layer3_outputs(1795) <= not(layer2_outputs(4592)) or (layer2_outputs(2939));
    layer3_outputs(1796) <= (layer2_outputs(3469)) or (layer2_outputs(1930));
    layer3_outputs(1797) <= not((layer2_outputs(1577)) xor (layer2_outputs(1490)));
    layer3_outputs(1798) <= not((layer2_outputs(927)) xor (layer2_outputs(1188)));
    layer3_outputs(1799) <= (layer2_outputs(7654)) or (layer2_outputs(1795));
    layer3_outputs(1800) <= not((layer2_outputs(7635)) or (layer2_outputs(6999)));
    layer3_outputs(1801) <= not((layer2_outputs(94)) xor (layer2_outputs(3471)));
    layer3_outputs(1802) <= not(layer2_outputs(2280)) or (layer2_outputs(5138));
    layer3_outputs(1803) <= (layer2_outputs(5134)) and not (layer2_outputs(6985));
    layer3_outputs(1804) <= not(layer2_outputs(6684));
    layer3_outputs(1805) <= not(layer2_outputs(1699));
    layer3_outputs(1806) <= (layer2_outputs(3421)) and not (layer2_outputs(2023));
    layer3_outputs(1807) <= not(layer2_outputs(1359));
    layer3_outputs(1808) <= layer2_outputs(5486);
    layer3_outputs(1809) <= not(layer2_outputs(5670)) or (layer2_outputs(337));
    layer3_outputs(1810) <= layer2_outputs(7659);
    layer3_outputs(1811) <= layer2_outputs(2273);
    layer3_outputs(1812) <= layer2_outputs(4117);
    layer3_outputs(1813) <= not(layer2_outputs(6565)) or (layer2_outputs(1731));
    layer3_outputs(1814) <= not((layer2_outputs(7036)) xor (layer2_outputs(5663)));
    layer3_outputs(1815) <= not((layer2_outputs(3890)) and (layer2_outputs(5322)));
    layer3_outputs(1816) <= layer2_outputs(2621);
    layer3_outputs(1817) <= (layer2_outputs(1996)) or (layer2_outputs(2883));
    layer3_outputs(1818) <= layer2_outputs(131);
    layer3_outputs(1819) <= not(layer2_outputs(7232));
    layer3_outputs(1820) <= (layer2_outputs(3018)) and (layer2_outputs(7010));
    layer3_outputs(1821) <= (layer2_outputs(7000)) or (layer2_outputs(1361));
    layer3_outputs(1822) <= not(layer2_outputs(471)) or (layer2_outputs(5293));
    layer3_outputs(1823) <= layer2_outputs(3581);
    layer3_outputs(1824) <= not(layer2_outputs(2862)) or (layer2_outputs(2414));
    layer3_outputs(1825) <= (layer2_outputs(7208)) xor (layer2_outputs(2796));
    layer3_outputs(1826) <= layer2_outputs(3222);
    layer3_outputs(1827) <= (layer2_outputs(3280)) and not (layer2_outputs(2192));
    layer3_outputs(1828) <= layer2_outputs(2861);
    layer3_outputs(1829) <= not(layer2_outputs(6711));
    layer3_outputs(1830) <= (layer2_outputs(2179)) xor (layer2_outputs(2943));
    layer3_outputs(1831) <= not(layer2_outputs(3527));
    layer3_outputs(1832) <= not(layer2_outputs(3779));
    layer3_outputs(1833) <= not((layer2_outputs(2866)) xor (layer2_outputs(4043)));
    layer3_outputs(1834) <= layer2_outputs(1825);
    layer3_outputs(1835) <= not((layer2_outputs(452)) xor (layer2_outputs(4798)));
    layer3_outputs(1836) <= layer2_outputs(1002);
    layer3_outputs(1837) <= not((layer2_outputs(2589)) and (layer2_outputs(6983)));
    layer3_outputs(1838) <= not((layer2_outputs(1370)) xor (layer2_outputs(7591)));
    layer3_outputs(1839) <= layer2_outputs(4939);
    layer3_outputs(1840) <= not((layer2_outputs(241)) and (layer2_outputs(2188)));
    layer3_outputs(1841) <= (layer2_outputs(4722)) and (layer2_outputs(697));
    layer3_outputs(1842) <= (layer2_outputs(783)) xor (layer2_outputs(5909));
    layer3_outputs(1843) <= '1';
    layer3_outputs(1844) <= '0';
    layer3_outputs(1845) <= not(layer2_outputs(6002));
    layer3_outputs(1846) <= not(layer2_outputs(67)) or (layer2_outputs(3507));
    layer3_outputs(1847) <= layer2_outputs(753);
    layer3_outputs(1848) <= not(layer2_outputs(6623));
    layer3_outputs(1849) <= not(layer2_outputs(2330)) or (layer2_outputs(6117));
    layer3_outputs(1850) <= (layer2_outputs(2626)) and not (layer2_outputs(5854));
    layer3_outputs(1851) <= not(layer2_outputs(6582)) or (layer2_outputs(6369));
    layer3_outputs(1852) <= not(layer2_outputs(6327));
    layer3_outputs(1853) <= layer2_outputs(603);
    layer3_outputs(1854) <= not(layer2_outputs(3081)) or (layer2_outputs(3773));
    layer3_outputs(1855) <= (layer2_outputs(1721)) xor (layer2_outputs(6500));
    layer3_outputs(1856) <= layer2_outputs(968);
    layer3_outputs(1857) <= not(layer2_outputs(6847));
    layer3_outputs(1858) <= not(layer2_outputs(2942));
    layer3_outputs(1859) <= not(layer2_outputs(3670)) or (layer2_outputs(5369));
    layer3_outputs(1860) <= not(layer2_outputs(5867)) or (layer2_outputs(5246));
    layer3_outputs(1861) <= layer2_outputs(6169);
    layer3_outputs(1862) <= not((layer2_outputs(3850)) or (layer2_outputs(6853)));
    layer3_outputs(1863) <= not(layer2_outputs(3085)) or (layer2_outputs(2260));
    layer3_outputs(1864) <= (layer2_outputs(3033)) xor (layer2_outputs(433));
    layer3_outputs(1865) <= not(layer2_outputs(6699));
    layer3_outputs(1866) <= not(layer2_outputs(826));
    layer3_outputs(1867) <= (layer2_outputs(2944)) and not (layer2_outputs(5918));
    layer3_outputs(1868) <= (layer2_outputs(812)) xor (layer2_outputs(7640));
    layer3_outputs(1869) <= (layer2_outputs(3621)) xor (layer2_outputs(2564));
    layer3_outputs(1870) <= (layer2_outputs(6917)) and not (layer2_outputs(3082));
    layer3_outputs(1871) <= '0';
    layer3_outputs(1872) <= not((layer2_outputs(3978)) and (layer2_outputs(6770)));
    layer3_outputs(1873) <= (layer2_outputs(7167)) and not (layer2_outputs(129));
    layer3_outputs(1874) <= (layer2_outputs(2675)) and not (layer2_outputs(6976));
    layer3_outputs(1875) <= (layer2_outputs(2758)) xor (layer2_outputs(3021));
    layer3_outputs(1876) <= not(layer2_outputs(6436)) or (layer2_outputs(528));
    layer3_outputs(1877) <= layer2_outputs(3813);
    layer3_outputs(1878) <= not(layer2_outputs(2772));
    layer3_outputs(1879) <= not(layer2_outputs(6987));
    layer3_outputs(1880) <= layer2_outputs(1398);
    layer3_outputs(1881) <= not(layer2_outputs(4151)) or (layer2_outputs(5953));
    layer3_outputs(1882) <= not((layer2_outputs(4585)) xor (layer2_outputs(33)));
    layer3_outputs(1883) <= not(layer2_outputs(7539));
    layer3_outputs(1884) <= (layer2_outputs(328)) and not (layer2_outputs(366));
    layer3_outputs(1885) <= '1';
    layer3_outputs(1886) <= not(layer2_outputs(1909));
    layer3_outputs(1887) <= not(layer2_outputs(1461)) or (layer2_outputs(999));
    layer3_outputs(1888) <= layer2_outputs(4491);
    layer3_outputs(1889) <= not(layer2_outputs(1261));
    layer3_outputs(1890) <= not((layer2_outputs(2810)) xor (layer2_outputs(6842)));
    layer3_outputs(1891) <= layer2_outputs(6718);
    layer3_outputs(1892) <= not((layer2_outputs(3353)) xor (layer2_outputs(2835)));
    layer3_outputs(1893) <= not((layer2_outputs(7514)) or (layer2_outputs(388)));
    layer3_outputs(1894) <= not(layer2_outputs(2641));
    layer3_outputs(1895) <= '0';
    layer3_outputs(1896) <= not((layer2_outputs(1162)) and (layer2_outputs(5279)));
    layer3_outputs(1897) <= not((layer2_outputs(5753)) and (layer2_outputs(2779)));
    layer3_outputs(1898) <= layer2_outputs(587);
    layer3_outputs(1899) <= not((layer2_outputs(464)) xor (layer2_outputs(4515)));
    layer3_outputs(1900) <= not(layer2_outputs(3314));
    layer3_outputs(1901) <= (layer2_outputs(215)) xor (layer2_outputs(6004));
    layer3_outputs(1902) <= '1';
    layer3_outputs(1903) <= (layer2_outputs(6173)) or (layer2_outputs(3006));
    layer3_outputs(1904) <= '1';
    layer3_outputs(1905) <= layer2_outputs(6416);
    layer3_outputs(1906) <= layer2_outputs(149);
    layer3_outputs(1907) <= (layer2_outputs(1694)) or (layer2_outputs(4536));
    layer3_outputs(1908) <= (layer2_outputs(1078)) or (layer2_outputs(2213));
    layer3_outputs(1909) <= not(layer2_outputs(2119));
    layer3_outputs(1910) <= not(layer2_outputs(7377));
    layer3_outputs(1911) <= (layer2_outputs(5550)) and (layer2_outputs(1150));
    layer3_outputs(1912) <= not(layer2_outputs(397));
    layer3_outputs(1913) <= (layer2_outputs(3663)) and not (layer2_outputs(2600));
    layer3_outputs(1914) <= (layer2_outputs(1493)) or (layer2_outputs(1896));
    layer3_outputs(1915) <= not(layer2_outputs(1532));
    layer3_outputs(1916) <= not((layer2_outputs(7499)) or (layer2_outputs(1130)));
    layer3_outputs(1917) <= not(layer2_outputs(3291)) or (layer2_outputs(3050));
    layer3_outputs(1918) <= not((layer2_outputs(1579)) and (layer2_outputs(2923)));
    layer3_outputs(1919) <= layer2_outputs(4215);
    layer3_outputs(1920) <= not((layer2_outputs(2323)) or (layer2_outputs(1457)));
    layer3_outputs(1921) <= not(layer2_outputs(4908));
    layer3_outputs(1922) <= layer2_outputs(634);
    layer3_outputs(1923) <= layer2_outputs(6558);
    layer3_outputs(1924) <= not(layer2_outputs(2247));
    layer3_outputs(1925) <= not(layer2_outputs(2497));
    layer3_outputs(1926) <= layer2_outputs(4443);
    layer3_outputs(1927) <= layer2_outputs(3007);
    layer3_outputs(1928) <= not(layer2_outputs(4424));
    layer3_outputs(1929) <= not((layer2_outputs(7001)) or (layer2_outputs(6603)));
    layer3_outputs(1930) <= (layer2_outputs(4560)) and not (layer2_outputs(958));
    layer3_outputs(1931) <= (layer2_outputs(6782)) or (layer2_outputs(1244));
    layer3_outputs(1932) <= (layer2_outputs(2706)) and not (layer2_outputs(1203));
    layer3_outputs(1933) <= layer2_outputs(678);
    layer3_outputs(1934) <= not(layer2_outputs(775));
    layer3_outputs(1935) <= (layer2_outputs(4828)) and not (layer2_outputs(7420));
    layer3_outputs(1936) <= not(layer2_outputs(7339));
    layer3_outputs(1937) <= not(layer2_outputs(5624));
    layer3_outputs(1938) <= '1';
    layer3_outputs(1939) <= layer2_outputs(4133);
    layer3_outputs(1940) <= (layer2_outputs(5281)) and not (layer2_outputs(2310));
    layer3_outputs(1941) <= layer2_outputs(468);
    layer3_outputs(1942) <= (layer2_outputs(2450)) xor (layer2_outputs(1160));
    layer3_outputs(1943) <= (layer2_outputs(3558)) and not (layer2_outputs(6253));
    layer3_outputs(1944) <= layer2_outputs(1568);
    layer3_outputs(1945) <= not(layer2_outputs(5412));
    layer3_outputs(1946) <= not((layer2_outputs(2521)) xor (layer2_outputs(6485)));
    layer3_outputs(1947) <= not(layer2_outputs(930));
    layer3_outputs(1948) <= (layer2_outputs(277)) xor (layer2_outputs(2954));
    layer3_outputs(1949) <= not(layer2_outputs(41));
    layer3_outputs(1950) <= not(layer2_outputs(3943));
    layer3_outputs(1951) <= layer2_outputs(1505);
    layer3_outputs(1952) <= '1';
    layer3_outputs(1953) <= layer2_outputs(3609);
    layer3_outputs(1954) <= layer2_outputs(7406);
    layer3_outputs(1955) <= not((layer2_outputs(4545)) and (layer2_outputs(1077)));
    layer3_outputs(1956) <= layer2_outputs(7414);
    layer3_outputs(1957) <= layer2_outputs(1446);
    layer3_outputs(1958) <= layer2_outputs(6974);
    layer3_outputs(1959) <= not(layer2_outputs(2504)) or (layer2_outputs(592));
    layer3_outputs(1960) <= (layer2_outputs(6544)) xor (layer2_outputs(2562));
    layer3_outputs(1961) <= layer2_outputs(935);
    layer3_outputs(1962) <= not(layer2_outputs(4391));
    layer3_outputs(1963) <= not(layer2_outputs(5105));
    layer3_outputs(1964) <= (layer2_outputs(2402)) and not (layer2_outputs(3447));
    layer3_outputs(1965) <= not((layer2_outputs(6481)) and (layer2_outputs(6249)));
    layer3_outputs(1966) <= not((layer2_outputs(1296)) and (layer2_outputs(4479)));
    layer3_outputs(1967) <= layer2_outputs(3986);
    layer3_outputs(1968) <= layer2_outputs(674);
    layer3_outputs(1969) <= not(layer2_outputs(1895)) or (layer2_outputs(5070));
    layer3_outputs(1970) <= not(layer2_outputs(6293));
    layer3_outputs(1971) <= layer2_outputs(385);
    layer3_outputs(1972) <= '1';
    layer3_outputs(1973) <= not((layer2_outputs(2526)) and (layer2_outputs(4202)));
    layer3_outputs(1974) <= not(layer2_outputs(7027));
    layer3_outputs(1975) <= layer2_outputs(5647);
    layer3_outputs(1976) <= not((layer2_outputs(2322)) xor (layer2_outputs(2611)));
    layer3_outputs(1977) <= not((layer2_outputs(2532)) and (layer2_outputs(931)));
    layer3_outputs(1978) <= not(layer2_outputs(7104)) or (layer2_outputs(4705));
    layer3_outputs(1979) <= layer2_outputs(6356);
    layer3_outputs(1980) <= not((layer2_outputs(2073)) and (layer2_outputs(5797)));
    layer3_outputs(1981) <= not((layer2_outputs(4046)) or (layer2_outputs(2246)));
    layer3_outputs(1982) <= layer2_outputs(5039);
    layer3_outputs(1983) <= layer2_outputs(2603);
    layer3_outputs(1984) <= not(layer2_outputs(3458)) or (layer2_outputs(178));
    layer3_outputs(1985) <= (layer2_outputs(2239)) and (layer2_outputs(6508));
    layer3_outputs(1986) <= not(layer2_outputs(369));
    layer3_outputs(1987) <= layer2_outputs(6124);
    layer3_outputs(1988) <= not(layer2_outputs(3043)) or (layer2_outputs(5569));
    layer3_outputs(1989) <= (layer2_outputs(4252)) and not (layer2_outputs(4265));
    layer3_outputs(1990) <= (layer2_outputs(7121)) or (layer2_outputs(6830));
    layer3_outputs(1991) <= not(layer2_outputs(6391));
    layer3_outputs(1992) <= (layer2_outputs(1506)) and (layer2_outputs(5426));
    layer3_outputs(1993) <= layer2_outputs(1906);
    layer3_outputs(1994) <= not((layer2_outputs(7349)) or (layer2_outputs(154)));
    layer3_outputs(1995) <= '0';
    layer3_outputs(1996) <= not(layer2_outputs(3769));
    layer3_outputs(1997) <= '1';
    layer3_outputs(1998) <= (layer2_outputs(3347)) or (layer2_outputs(2392));
    layer3_outputs(1999) <= not(layer2_outputs(4881));
    layer3_outputs(2000) <= layer2_outputs(1783);
    layer3_outputs(2001) <= not(layer2_outputs(3713)) or (layer2_outputs(3651));
    layer3_outputs(2002) <= not((layer2_outputs(6216)) and (layer2_outputs(6882)));
    layer3_outputs(2003) <= layer2_outputs(1271);
    layer3_outputs(2004) <= not(layer2_outputs(2693));
    layer3_outputs(2005) <= not(layer2_outputs(3930));
    layer3_outputs(2006) <= not(layer2_outputs(2784)) or (layer2_outputs(2558));
    layer3_outputs(2007) <= (layer2_outputs(4580)) and (layer2_outputs(1073));
    layer3_outputs(2008) <= not(layer2_outputs(2048));
    layer3_outputs(2009) <= not(layer2_outputs(3281));
    layer3_outputs(2010) <= not(layer2_outputs(5747)) or (layer2_outputs(4523));
    layer3_outputs(2011) <= not(layer2_outputs(2534));
    layer3_outputs(2012) <= layer2_outputs(7668);
    layer3_outputs(2013) <= not((layer2_outputs(5605)) or (layer2_outputs(1474)));
    layer3_outputs(2014) <= layer2_outputs(1685);
    layer3_outputs(2015) <= not((layer2_outputs(722)) or (layer2_outputs(5992)));
    layer3_outputs(2016) <= not(layer2_outputs(2218));
    layer3_outputs(2017) <= not((layer2_outputs(1200)) or (layer2_outputs(2858)));
    layer3_outputs(2018) <= not(layer2_outputs(1112));
    layer3_outputs(2019) <= not((layer2_outputs(4508)) xor (layer2_outputs(4680)));
    layer3_outputs(2020) <= layer2_outputs(1617);
    layer3_outputs(2021) <= (layer2_outputs(7194)) or (layer2_outputs(7229));
    layer3_outputs(2022) <= not((layer2_outputs(1205)) or (layer2_outputs(1696)));
    layer3_outputs(2023) <= (layer2_outputs(1429)) or (layer2_outputs(4628));
    layer3_outputs(2024) <= (layer2_outputs(3900)) and (layer2_outputs(4157));
    layer3_outputs(2025) <= not(layer2_outputs(3382));
    layer3_outputs(2026) <= not((layer2_outputs(2917)) or (layer2_outputs(7120)));
    layer3_outputs(2027) <= (layer2_outputs(6234)) and (layer2_outputs(7085));
    layer3_outputs(2028) <= not(layer2_outputs(4150));
    layer3_outputs(2029) <= (layer2_outputs(2465)) or (layer2_outputs(15));
    layer3_outputs(2030) <= not((layer2_outputs(4361)) and (layer2_outputs(4842)));
    layer3_outputs(2031) <= layer2_outputs(3192);
    layer3_outputs(2032) <= (layer2_outputs(2194)) and (layer2_outputs(8));
    layer3_outputs(2033) <= layer2_outputs(5342);
    layer3_outputs(2034) <= layer2_outputs(2104);
    layer3_outputs(2035) <= not(layer2_outputs(3366));
    layer3_outputs(2036) <= not((layer2_outputs(192)) and (layer2_outputs(2227)));
    layer3_outputs(2037) <= layer2_outputs(6998);
    layer3_outputs(2038) <= (layer2_outputs(2497)) or (layer2_outputs(1717));
    layer3_outputs(2039) <= not((layer2_outputs(6342)) or (layer2_outputs(4242)));
    layer3_outputs(2040) <= not(layer2_outputs(4871)) or (layer2_outputs(4007));
    layer3_outputs(2041) <= (layer2_outputs(6719)) and not (layer2_outputs(4797));
    layer3_outputs(2042) <= (layer2_outputs(125)) and not (layer2_outputs(5548));
    layer3_outputs(2043) <= not(layer2_outputs(196));
    layer3_outputs(2044) <= not(layer2_outputs(3156));
    layer3_outputs(2045) <= not((layer2_outputs(6919)) or (layer2_outputs(5951)));
    layer3_outputs(2046) <= not(layer2_outputs(3686)) or (layer2_outputs(198));
    layer3_outputs(2047) <= layer2_outputs(652);
    layer3_outputs(2048) <= not(layer2_outputs(1817));
    layer3_outputs(2049) <= (layer2_outputs(5150)) or (layer2_outputs(3513));
    layer3_outputs(2050) <= (layer2_outputs(7614)) or (layer2_outputs(4069));
    layer3_outputs(2051) <= not(layer2_outputs(2097));
    layer3_outputs(2052) <= (layer2_outputs(6484)) and not (layer2_outputs(5131));
    layer3_outputs(2053) <= layer2_outputs(3943);
    layer3_outputs(2054) <= layer2_outputs(5346);
    layer3_outputs(2055) <= (layer2_outputs(7144)) and not (layer2_outputs(5749));
    layer3_outputs(2056) <= not(layer2_outputs(5682));
    layer3_outputs(2057) <= not(layer2_outputs(6432)) or (layer2_outputs(348));
    layer3_outputs(2058) <= not(layer2_outputs(6617)) or (layer2_outputs(1626));
    layer3_outputs(2059) <= not(layer2_outputs(2717));
    layer3_outputs(2060) <= not(layer2_outputs(831));
    layer3_outputs(2061) <= not(layer2_outputs(4799));
    layer3_outputs(2062) <= (layer2_outputs(1036)) and not (layer2_outputs(1452));
    layer3_outputs(2063) <= '0';
    layer3_outputs(2064) <= '1';
    layer3_outputs(2065) <= (layer2_outputs(1316)) and (layer2_outputs(7605));
    layer3_outputs(2066) <= layer2_outputs(6555);
    layer3_outputs(2067) <= not(layer2_outputs(2013));
    layer3_outputs(2068) <= (layer2_outputs(2467)) or (layer2_outputs(1979));
    layer3_outputs(2069) <= not(layer2_outputs(960));
    layer3_outputs(2070) <= layer2_outputs(4129);
    layer3_outputs(2071) <= (layer2_outputs(3926)) or (layer2_outputs(1177));
    layer3_outputs(2072) <= layer2_outputs(1837);
    layer3_outputs(2073) <= not((layer2_outputs(5325)) xor (layer2_outputs(2947)));
    layer3_outputs(2074) <= (layer2_outputs(482)) xor (layer2_outputs(3654));
    layer3_outputs(2075) <= not(layer2_outputs(5636));
    layer3_outputs(2076) <= not(layer2_outputs(768));
    layer3_outputs(2077) <= layer2_outputs(3533);
    layer3_outputs(2078) <= not((layer2_outputs(7059)) and (layer2_outputs(1709)));
    layer3_outputs(2079) <= not((layer2_outputs(2507)) xor (layer2_outputs(5141)));
    layer3_outputs(2080) <= not(layer2_outputs(2922)) or (layer2_outputs(7253));
    layer3_outputs(2081) <= not((layer2_outputs(1049)) and (layer2_outputs(2924)));
    layer3_outputs(2082) <= not(layer2_outputs(415));
    layer3_outputs(2083) <= not((layer2_outputs(7122)) or (layer2_outputs(2130)));
    layer3_outputs(2084) <= not((layer2_outputs(671)) or (layer2_outputs(2505)));
    layer3_outputs(2085) <= not(layer2_outputs(6883)) or (layer2_outputs(7214));
    layer3_outputs(2086) <= not(layer2_outputs(6582)) or (layer2_outputs(995));
    layer3_outputs(2087) <= not(layer2_outputs(6930));
    layer3_outputs(2088) <= not(layer2_outputs(1047));
    layer3_outputs(2089) <= not(layer2_outputs(4896)) or (layer2_outputs(5329));
    layer3_outputs(2090) <= layer2_outputs(4169);
    layer3_outputs(2091) <= layer2_outputs(141);
    layer3_outputs(2092) <= not((layer2_outputs(5344)) and (layer2_outputs(5117)));
    layer3_outputs(2093) <= not(layer2_outputs(1640));
    layer3_outputs(2094) <= (layer2_outputs(4455)) and (layer2_outputs(3646));
    layer3_outputs(2095) <= not((layer2_outputs(20)) and (layer2_outputs(7537)));
    layer3_outputs(2096) <= not(layer2_outputs(5494));
    layer3_outputs(2097) <= not(layer2_outputs(4091)) or (layer2_outputs(4942));
    layer3_outputs(2098) <= layer2_outputs(2172);
    layer3_outputs(2099) <= layer2_outputs(7464);
    layer3_outputs(2100) <= not(layer2_outputs(4894));
    layer3_outputs(2101) <= layer2_outputs(4373);
    layer3_outputs(2102) <= not((layer2_outputs(4572)) or (layer2_outputs(3094)));
    layer3_outputs(2103) <= not((layer2_outputs(1700)) or (layer2_outputs(3810)));
    layer3_outputs(2104) <= layer2_outputs(3959);
    layer3_outputs(2105) <= not(layer2_outputs(6077));
    layer3_outputs(2106) <= (layer2_outputs(365)) and not (layer2_outputs(3406));
    layer3_outputs(2107) <= layer2_outputs(5626);
    layer3_outputs(2108) <= (layer2_outputs(3785)) and not (layer2_outputs(472));
    layer3_outputs(2109) <= not((layer2_outputs(7677)) xor (layer2_outputs(2233)));
    layer3_outputs(2110) <= not(layer2_outputs(1482));
    layer3_outputs(2111) <= layer2_outputs(6723);
    layer3_outputs(2112) <= '1';
    layer3_outputs(2113) <= not(layer2_outputs(2171));
    layer3_outputs(2114) <= not(layer2_outputs(6038));
    layer3_outputs(2115) <= (layer2_outputs(1514)) or (layer2_outputs(3530));
    layer3_outputs(2116) <= '0';
    layer3_outputs(2117) <= not((layer2_outputs(7217)) or (layer2_outputs(3513)));
    layer3_outputs(2118) <= not(layer2_outputs(986)) or (layer2_outputs(1602));
    layer3_outputs(2119) <= not(layer2_outputs(7223)) or (layer2_outputs(88));
    layer3_outputs(2120) <= layer2_outputs(5136);
    layer3_outputs(2121) <= not((layer2_outputs(2941)) or (layer2_outputs(7320)));
    layer3_outputs(2122) <= layer2_outputs(1729);
    layer3_outputs(2123) <= (layer2_outputs(6268)) and (layer2_outputs(6219));
    layer3_outputs(2124) <= not(layer2_outputs(6993));
    layer3_outputs(2125) <= layer2_outputs(2770);
    layer3_outputs(2126) <= not(layer2_outputs(7450));
    layer3_outputs(2127) <= not(layer2_outputs(6173)) or (layer2_outputs(3961));
    layer3_outputs(2128) <= not(layer2_outputs(4685)) or (layer2_outputs(957));
    layer3_outputs(2129) <= layer2_outputs(6466);
    layer3_outputs(2130) <= not(layer2_outputs(6513));
    layer3_outputs(2131) <= (layer2_outputs(5220)) and not (layer2_outputs(3291));
    layer3_outputs(2132) <= not((layer2_outputs(5024)) and (layer2_outputs(1039)));
    layer3_outputs(2133) <= layer2_outputs(1126);
    layer3_outputs(2134) <= not((layer2_outputs(6052)) xor (layer2_outputs(4752)));
    layer3_outputs(2135) <= not(layer2_outputs(4658)) or (layer2_outputs(5068));
    layer3_outputs(2136) <= not((layer2_outputs(7660)) or (layer2_outputs(6701)));
    layer3_outputs(2137) <= not(layer2_outputs(1868));
    layer3_outputs(2138) <= not((layer2_outputs(5288)) or (layer2_outputs(1875)));
    layer3_outputs(2139) <= not(layer2_outputs(672)) or (layer2_outputs(5952));
    layer3_outputs(2140) <= layer2_outputs(6813);
    layer3_outputs(2141) <= not((layer2_outputs(7491)) or (layer2_outputs(4489)));
    layer3_outputs(2142) <= (layer2_outputs(6972)) and not (layer2_outputs(2101));
    layer3_outputs(2143) <= not(layer2_outputs(4837));
    layer3_outputs(2144) <= '1';
    layer3_outputs(2145) <= not(layer2_outputs(5194)) or (layer2_outputs(604));
    layer3_outputs(2146) <= (layer2_outputs(900)) and (layer2_outputs(1404));
    layer3_outputs(2147) <= not(layer2_outputs(6237));
    layer3_outputs(2148) <= (layer2_outputs(4141)) and (layer2_outputs(4379));
    layer3_outputs(2149) <= not((layer2_outputs(3498)) xor (layer2_outputs(2492)));
    layer3_outputs(2150) <= (layer2_outputs(6863)) and not (layer2_outputs(2526));
    layer3_outputs(2151) <= (layer2_outputs(6809)) and (layer2_outputs(3511));
    layer3_outputs(2152) <= not(layer2_outputs(1927)) or (layer2_outputs(2080));
    layer3_outputs(2153) <= (layer2_outputs(2528)) xor (layer2_outputs(2478));
    layer3_outputs(2154) <= not((layer2_outputs(7204)) or (layer2_outputs(4029)));
    layer3_outputs(2155) <= (layer2_outputs(1833)) and (layer2_outputs(3526));
    layer3_outputs(2156) <= not(layer2_outputs(1624));
    layer3_outputs(2157) <= not(layer2_outputs(1966));
    layer3_outputs(2158) <= not((layer2_outputs(7200)) xor (layer2_outputs(5299)));
    layer3_outputs(2159) <= not(layer2_outputs(1954));
    layer3_outputs(2160) <= (layer2_outputs(2276)) or (layer2_outputs(918));
    layer3_outputs(2161) <= not(layer2_outputs(3239)) or (layer2_outputs(4959));
    layer3_outputs(2162) <= not((layer2_outputs(124)) and (layer2_outputs(5076)));
    layer3_outputs(2163) <= not(layer2_outputs(4886));
    layer3_outputs(2164) <= not(layer2_outputs(6800)) or (layer2_outputs(7535));
    layer3_outputs(2165) <= (layer2_outputs(7578)) xor (layer2_outputs(1703));
    layer3_outputs(2166) <= not((layer2_outputs(5369)) or (layer2_outputs(2689)));
    layer3_outputs(2167) <= (layer2_outputs(4787)) or (layer2_outputs(7222));
    layer3_outputs(2168) <= not(layer2_outputs(2129));
    layer3_outputs(2169) <= not((layer2_outputs(7218)) xor (layer2_outputs(7068)));
    layer3_outputs(2170) <= (layer2_outputs(4212)) and not (layer2_outputs(840));
    layer3_outputs(2171) <= not((layer2_outputs(761)) xor (layer2_outputs(4897)));
    layer3_outputs(2172) <= (layer2_outputs(1574)) or (layer2_outputs(6977));
    layer3_outputs(2173) <= not(layer2_outputs(3435));
    layer3_outputs(2174) <= not((layer2_outputs(1367)) or (layer2_outputs(7554)));
    layer3_outputs(2175) <= not(layer2_outputs(5817));
    layer3_outputs(2176) <= layer2_outputs(3372);
    layer3_outputs(2177) <= not(layer2_outputs(1110));
    layer3_outputs(2178) <= layer2_outputs(2985);
    layer3_outputs(2179) <= '1';
    layer3_outputs(2180) <= not((layer2_outputs(890)) and (layer2_outputs(1692)));
    layer3_outputs(2181) <= (layer2_outputs(4727)) xor (layer2_outputs(4520));
    layer3_outputs(2182) <= (layer2_outputs(4439)) and (layer2_outputs(2222));
    layer3_outputs(2183) <= not(layer2_outputs(2005));
    layer3_outputs(2184) <= layer2_outputs(5556);
    layer3_outputs(2185) <= not((layer2_outputs(6745)) and (layer2_outputs(7296)));
    layer3_outputs(2186) <= (layer2_outputs(431)) and (layer2_outputs(965));
    layer3_outputs(2187) <= layer2_outputs(2580);
    layer3_outputs(2188) <= not((layer2_outputs(1442)) and (layer2_outputs(3563)));
    layer3_outputs(2189) <= (layer2_outputs(4640)) or (layer2_outputs(1157));
    layer3_outputs(2190) <= not((layer2_outputs(6658)) and (layer2_outputs(6170)));
    layer3_outputs(2191) <= (layer2_outputs(4417)) and not (layer2_outputs(5933));
    layer3_outputs(2192) <= layer2_outputs(134);
    layer3_outputs(2193) <= not(layer2_outputs(177));
    layer3_outputs(2194) <= not((layer2_outputs(2403)) and (layer2_outputs(92)));
    layer3_outputs(2195) <= not((layer2_outputs(2374)) or (layer2_outputs(5228)));
    layer3_outputs(2196) <= not(layer2_outputs(4976));
    layer3_outputs(2197) <= (layer2_outputs(2965)) and not (layer2_outputs(5296));
    layer3_outputs(2198) <= not((layer2_outputs(762)) and (layer2_outputs(4186)));
    layer3_outputs(2199) <= (layer2_outputs(6917)) and not (layer2_outputs(6508));
    layer3_outputs(2200) <= (layer2_outputs(7456)) and not (layer2_outputs(6266));
    layer3_outputs(2201) <= not(layer2_outputs(985)) or (layer2_outputs(6988));
    layer3_outputs(2202) <= layer2_outputs(4753);
    layer3_outputs(2203) <= not(layer2_outputs(4990));
    layer3_outputs(2204) <= not((layer2_outputs(1776)) or (layer2_outputs(4290)));
    layer3_outputs(2205) <= not(layer2_outputs(1257));
    layer3_outputs(2206) <= (layer2_outputs(7434)) and not (layer2_outputs(6269));
    layer3_outputs(2207) <= (layer2_outputs(4510)) and not (layer2_outputs(1305));
    layer3_outputs(2208) <= not(layer2_outputs(6567));
    layer3_outputs(2209) <= layer2_outputs(3644);
    layer3_outputs(2210) <= (layer2_outputs(2608)) and not (layer2_outputs(84));
    layer3_outputs(2211) <= (layer2_outputs(1812)) and not (layer2_outputs(2038));
    layer3_outputs(2212) <= (layer2_outputs(5941)) and not (layer2_outputs(6153));
    layer3_outputs(2213) <= not(layer2_outputs(593));
    layer3_outputs(2214) <= layer2_outputs(6948);
    layer3_outputs(2215) <= not(layer2_outputs(6758));
    layer3_outputs(2216) <= layer2_outputs(4446);
    layer3_outputs(2217) <= not((layer2_outputs(1985)) or (layer2_outputs(3142)));
    layer3_outputs(2218) <= layer2_outputs(6785);
    layer3_outputs(2219) <= (layer2_outputs(1333)) or (layer2_outputs(7262));
    layer3_outputs(2220) <= layer2_outputs(3795);
    layer3_outputs(2221) <= not((layer2_outputs(3456)) or (layer2_outputs(6891)));
    layer3_outputs(2222) <= (layer2_outputs(3251)) and (layer2_outputs(2436));
    layer3_outputs(2223) <= (layer2_outputs(5037)) or (layer2_outputs(6055));
    layer3_outputs(2224) <= layer2_outputs(6375);
    layer3_outputs(2225) <= layer2_outputs(5541);
    layer3_outputs(2226) <= not(layer2_outputs(1395)) or (layer2_outputs(1321));
    layer3_outputs(2227) <= layer2_outputs(5560);
    layer3_outputs(2228) <= not((layer2_outputs(853)) and (layer2_outputs(4453)));
    layer3_outputs(2229) <= not((layer2_outputs(3803)) and (layer2_outputs(4449)));
    layer3_outputs(2230) <= (layer2_outputs(7323)) and not (layer2_outputs(4032));
    layer3_outputs(2231) <= not(layer2_outputs(1647));
    layer3_outputs(2232) <= layer2_outputs(905);
    layer3_outputs(2233) <= layer2_outputs(4176);
    layer3_outputs(2234) <= layer2_outputs(3639);
    layer3_outputs(2235) <= not(layer2_outputs(51)) or (layer2_outputs(602));
    layer3_outputs(2236) <= layer2_outputs(3944);
    layer3_outputs(2237) <= not(layer2_outputs(1798));
    layer3_outputs(2238) <= not(layer2_outputs(1811));
    layer3_outputs(2239) <= '1';
    layer3_outputs(2240) <= (layer2_outputs(6661)) and (layer2_outputs(1879));
    layer3_outputs(2241) <= not(layer2_outputs(6446)) or (layer2_outputs(5649));
    layer3_outputs(2242) <= layer2_outputs(2782);
    layer3_outputs(2243) <= not((layer2_outputs(6093)) and (layer2_outputs(2177)));
    layer3_outputs(2244) <= (layer2_outputs(5717)) xor (layer2_outputs(7002));
    layer3_outputs(2245) <= (layer2_outputs(2019)) and (layer2_outputs(6346));
    layer3_outputs(2246) <= layer2_outputs(1632);
    layer3_outputs(2247) <= layer2_outputs(7565);
    layer3_outputs(2248) <= not(layer2_outputs(5331));
    layer3_outputs(2249) <= layer2_outputs(3892);
    layer3_outputs(2250) <= not((layer2_outputs(3882)) or (layer2_outputs(5248)));
    layer3_outputs(2251) <= not(layer2_outputs(855));
    layer3_outputs(2252) <= not(layer2_outputs(1586)) or (layer2_outputs(5549));
    layer3_outputs(2253) <= layer2_outputs(6906);
    layer3_outputs(2254) <= layer2_outputs(301);
    layer3_outputs(2255) <= not(layer2_outputs(4566));
    layer3_outputs(2256) <= not(layer2_outputs(2981));
    layer3_outputs(2257) <= (layer2_outputs(7150)) and not (layer2_outputs(2639));
    layer3_outputs(2258) <= not(layer2_outputs(1002));
    layer3_outputs(2259) <= (layer2_outputs(325)) and (layer2_outputs(5523));
    layer3_outputs(2260) <= not(layer2_outputs(3371));
    layer3_outputs(2261) <= not((layer2_outputs(1950)) and (layer2_outputs(3490)));
    layer3_outputs(2262) <= not(layer2_outputs(6493)) or (layer2_outputs(3071));
    layer3_outputs(2263) <= (layer2_outputs(6512)) and (layer2_outputs(4498));
    layer3_outputs(2264) <= layer2_outputs(6653);
    layer3_outputs(2265) <= not((layer2_outputs(3626)) and (layer2_outputs(4651)));
    layer3_outputs(2266) <= (layer2_outputs(6409)) xor (layer2_outputs(1160));
    layer3_outputs(2267) <= not(layer2_outputs(6384)) or (layer2_outputs(6694));
    layer3_outputs(2268) <= not(layer2_outputs(387));
    layer3_outputs(2269) <= not(layer2_outputs(3045));
    layer3_outputs(2270) <= not((layer2_outputs(1227)) or (layer2_outputs(1735)));
    layer3_outputs(2271) <= not(layer2_outputs(4550));
    layer3_outputs(2272) <= not((layer2_outputs(3348)) or (layer2_outputs(228)));
    layer3_outputs(2273) <= not(layer2_outputs(4776)) or (layer2_outputs(624));
    layer3_outputs(2274) <= not((layer2_outputs(5940)) or (layer2_outputs(2723)));
    layer3_outputs(2275) <= (layer2_outputs(92)) and (layer2_outputs(3877));
    layer3_outputs(2276) <= layer2_outputs(3017);
    layer3_outputs(2277) <= (layer2_outputs(3566)) and not (layer2_outputs(3243));
    layer3_outputs(2278) <= not((layer2_outputs(1352)) and (layer2_outputs(6050)));
    layer3_outputs(2279) <= (layer2_outputs(5354)) xor (layer2_outputs(119));
    layer3_outputs(2280) <= '1';
    layer3_outputs(2281) <= (layer2_outputs(1192)) and not (layer2_outputs(3123));
    layer3_outputs(2282) <= (layer2_outputs(7360)) or (layer2_outputs(1985));
    layer3_outputs(2283) <= (layer2_outputs(4581)) and not (layer2_outputs(2360));
    layer3_outputs(2284) <= '1';
    layer3_outputs(2285) <= layer2_outputs(3890);
    layer3_outputs(2286) <= not(layer2_outputs(2054));
    layer3_outputs(2287) <= not(layer2_outputs(5569));
    layer3_outputs(2288) <= (layer2_outputs(1802)) and (layer2_outputs(5252));
    layer3_outputs(2289) <= not(layer2_outputs(4412));
    layer3_outputs(2290) <= (layer2_outputs(5183)) and (layer2_outputs(3595));
    layer3_outputs(2291) <= not(layer2_outputs(6630));
    layer3_outputs(2292) <= layer2_outputs(6249);
    layer3_outputs(2293) <= not((layer2_outputs(5387)) and (layer2_outputs(4360)));
    layer3_outputs(2294) <= not(layer2_outputs(5696));
    layer3_outputs(2295) <= (layer2_outputs(4311)) and not (layer2_outputs(2170));
    layer3_outputs(2296) <= not(layer2_outputs(7117));
    layer3_outputs(2297) <= not((layer2_outputs(31)) xor (layer2_outputs(6843)));
    layer3_outputs(2298) <= layer2_outputs(3095);
    layer3_outputs(2299) <= not((layer2_outputs(2668)) and (layer2_outputs(5574)));
    layer3_outputs(2300) <= layer2_outputs(239);
    layer3_outputs(2301) <= not(layer2_outputs(5923)) or (layer2_outputs(5621));
    layer3_outputs(2302) <= (layer2_outputs(6557)) or (layer2_outputs(5671));
    layer3_outputs(2303) <= not(layer2_outputs(3039));
    layer3_outputs(2304) <= layer2_outputs(135);
    layer3_outputs(2305) <= (layer2_outputs(7254)) xor (layer2_outputs(6190));
    layer3_outputs(2306) <= (layer2_outputs(572)) and not (layer2_outputs(7312));
    layer3_outputs(2307) <= '0';
    layer3_outputs(2308) <= not(layer2_outputs(5222));
    layer3_outputs(2309) <= not(layer2_outputs(5072));
    layer3_outputs(2310) <= layer2_outputs(6864);
    layer3_outputs(2311) <= '0';
    layer3_outputs(2312) <= not(layer2_outputs(828));
    layer3_outputs(2313) <= layer2_outputs(4792);
    layer3_outputs(2314) <= (layer2_outputs(146)) and not (layer2_outputs(1303));
    layer3_outputs(2315) <= not((layer2_outputs(679)) and (layer2_outputs(7399)));
    layer3_outputs(2316) <= not((layer2_outputs(3173)) and (layer2_outputs(294)));
    layer3_outputs(2317) <= not((layer2_outputs(2325)) and (layer2_outputs(4359)));
    layer3_outputs(2318) <= not((layer2_outputs(6614)) xor (layer2_outputs(4899)));
    layer3_outputs(2319) <= (layer2_outputs(811)) and (layer2_outputs(4924));
    layer3_outputs(2320) <= (layer2_outputs(2167)) and not (layer2_outputs(5241));
    layer3_outputs(2321) <= not(layer2_outputs(1242));
    layer3_outputs(2322) <= (layer2_outputs(6876)) and not (layer2_outputs(6103));
    layer3_outputs(2323) <= not(layer2_outputs(2308));
    layer3_outputs(2324) <= layer2_outputs(1878);
    layer3_outputs(2325) <= not(layer2_outputs(6358)) or (layer2_outputs(1408));
    layer3_outputs(2326) <= not(layer2_outputs(6028)) or (layer2_outputs(3822));
    layer3_outputs(2327) <= layer2_outputs(7313);
    layer3_outputs(2328) <= layer2_outputs(1053);
    layer3_outputs(2329) <= not(layer2_outputs(704)) or (layer2_outputs(2656));
    layer3_outputs(2330) <= not(layer2_outputs(948));
    layer3_outputs(2331) <= not(layer2_outputs(6130)) or (layer2_outputs(2895));
    layer3_outputs(2332) <= not(layer2_outputs(4125));
    layer3_outputs(2333) <= (layer2_outputs(5995)) or (layer2_outputs(6265));
    layer3_outputs(2334) <= '1';
    layer3_outputs(2335) <= not((layer2_outputs(1591)) or (layer2_outputs(3859)));
    layer3_outputs(2336) <= (layer2_outputs(1972)) or (layer2_outputs(7486));
    layer3_outputs(2337) <= not((layer2_outputs(7374)) xor (layer2_outputs(5775)));
    layer3_outputs(2338) <= not((layer2_outputs(4555)) and (layer2_outputs(3052)));
    layer3_outputs(2339) <= layer2_outputs(1455);
    layer3_outputs(2340) <= (layer2_outputs(6692)) and (layer2_outputs(1191));
    layer3_outputs(2341) <= not((layer2_outputs(7163)) xor (layer2_outputs(3980)));
    layer3_outputs(2342) <= (layer2_outputs(2134)) and not (layer2_outputs(4638));
    layer3_outputs(2343) <= layer2_outputs(2133);
    layer3_outputs(2344) <= not(layer2_outputs(1456)) or (layer2_outputs(4067));
    layer3_outputs(2345) <= not((layer2_outputs(4397)) and (layer2_outputs(3918)));
    layer3_outputs(2346) <= not(layer2_outputs(4562));
    layer3_outputs(2347) <= not(layer2_outputs(6100));
    layer3_outputs(2348) <= layer2_outputs(7375);
    layer3_outputs(2349) <= not(layer2_outputs(2590)) or (layer2_outputs(3739));
    layer3_outputs(2350) <= (layer2_outputs(7131)) and not (layer2_outputs(1116));
    layer3_outputs(2351) <= (layer2_outputs(2798)) and not (layer2_outputs(223));
    layer3_outputs(2352) <= not((layer2_outputs(651)) or (layer2_outputs(1153)));
    layer3_outputs(2353) <= layer2_outputs(1960);
    layer3_outputs(2354) <= not(layer2_outputs(3632));
    layer3_outputs(2355) <= layer2_outputs(7013);
    layer3_outputs(2356) <= not(layer2_outputs(1192));
    layer3_outputs(2357) <= not((layer2_outputs(6784)) and (layer2_outputs(7007)));
    layer3_outputs(2358) <= not(layer2_outputs(3342));
    layer3_outputs(2359) <= not(layer2_outputs(15));
    layer3_outputs(2360) <= layer2_outputs(2790);
    layer3_outputs(2361) <= layer2_outputs(2151);
    layer3_outputs(2362) <= not(layer2_outputs(447)) or (layer2_outputs(6322));
    layer3_outputs(2363) <= layer2_outputs(2336);
    layer3_outputs(2364) <= (layer2_outputs(4540)) and not (layer2_outputs(3152));
    layer3_outputs(2365) <= not(layer2_outputs(2426));
    layer3_outputs(2366) <= '1';
    layer3_outputs(2367) <= (layer2_outputs(6528)) or (layer2_outputs(3614));
    layer3_outputs(2368) <= (layer2_outputs(326)) and not (layer2_outputs(7037));
    layer3_outputs(2369) <= not(layer2_outputs(5541));
    layer3_outputs(2370) <= (layer2_outputs(7095)) xor (layer2_outputs(4646));
    layer3_outputs(2371) <= (layer2_outputs(7569)) or (layer2_outputs(3695));
    layer3_outputs(2372) <= not(layer2_outputs(3183));
    layer3_outputs(2373) <= not(layer2_outputs(6600)) or (layer2_outputs(1991));
    layer3_outputs(2374) <= not(layer2_outputs(7607));
    layer3_outputs(2375) <= not(layer2_outputs(454));
    layer3_outputs(2376) <= (layer2_outputs(5931)) xor (layer2_outputs(5954));
    layer3_outputs(2377) <= layer2_outputs(4884);
    layer3_outputs(2378) <= layer2_outputs(32);
    layer3_outputs(2379) <= (layer2_outputs(5416)) xor (layer2_outputs(2618));
    layer3_outputs(2380) <= layer2_outputs(2795);
    layer3_outputs(2381) <= not(layer2_outputs(7566));
    layer3_outputs(2382) <= layer2_outputs(2018);
    layer3_outputs(2383) <= not(layer2_outputs(1084)) or (layer2_outputs(7593));
    layer3_outputs(2384) <= '0';
    layer3_outputs(2385) <= (layer2_outputs(6638)) and not (layer2_outputs(5817));
    layer3_outputs(2386) <= (layer2_outputs(5262)) and (layer2_outputs(402));
    layer3_outputs(2387) <= layer2_outputs(1380);
    layer3_outputs(2388) <= (layer2_outputs(371)) and not (layer2_outputs(1570));
    layer3_outputs(2389) <= not(layer2_outputs(2694));
    layer3_outputs(2390) <= layer2_outputs(7087);
    layer3_outputs(2391) <= layer2_outputs(1252);
    layer3_outputs(2392) <= not(layer2_outputs(7044));
    layer3_outputs(2393) <= layer2_outputs(1862);
    layer3_outputs(2394) <= (layer2_outputs(6267)) or (layer2_outputs(7372));
    layer3_outputs(2395) <= (layer2_outputs(6756)) and not (layer2_outputs(1376));
    layer3_outputs(2396) <= (layer2_outputs(3992)) and not (layer2_outputs(1437));
    layer3_outputs(2397) <= (layer2_outputs(6429)) or (layer2_outputs(612));
    layer3_outputs(2398) <= not(layer2_outputs(1646));
    layer3_outputs(2399) <= not(layer2_outputs(3964));
    layer3_outputs(2400) <= layer2_outputs(540);
    layer3_outputs(2401) <= not(layer2_outputs(1137));
    layer3_outputs(2402) <= not(layer2_outputs(6306));
    layer3_outputs(2403) <= not(layer2_outputs(5015));
    layer3_outputs(2404) <= not((layer2_outputs(3867)) or (layer2_outputs(6482)));
    layer3_outputs(2405) <= '0';
    layer3_outputs(2406) <= not((layer2_outputs(209)) or (layer2_outputs(3706)));
    layer3_outputs(2407) <= not((layer2_outputs(3520)) or (layer2_outputs(128)));
    layer3_outputs(2408) <= layer2_outputs(1816);
    layer3_outputs(2409) <= not((layer2_outputs(1488)) or (layer2_outputs(5645)));
    layer3_outputs(2410) <= (layer2_outputs(4544)) and not (layer2_outputs(7410));
    layer3_outputs(2411) <= layer2_outputs(4625);
    layer3_outputs(2412) <= (layer2_outputs(3532)) and (layer2_outputs(1495));
    layer3_outputs(2413) <= layer2_outputs(4462);
    layer3_outputs(2414) <= not((layer2_outputs(57)) xor (layer2_outputs(498)));
    layer3_outputs(2415) <= (layer2_outputs(5176)) and not (layer2_outputs(522));
    layer3_outputs(2416) <= layer2_outputs(4134);
    layer3_outputs(2417) <= layer2_outputs(2773);
    layer3_outputs(2418) <= not((layer2_outputs(1410)) xor (layer2_outputs(3693)));
    layer3_outputs(2419) <= not(layer2_outputs(4219)) or (layer2_outputs(1977));
    layer3_outputs(2420) <= layer2_outputs(6210);
    layer3_outputs(2421) <= not(layer2_outputs(6448)) or (layer2_outputs(2886));
    layer3_outputs(2422) <= not((layer2_outputs(6576)) or (layer2_outputs(3837)));
    layer3_outputs(2423) <= not((layer2_outputs(3041)) and (layer2_outputs(6067)));
    layer3_outputs(2424) <= layer2_outputs(7333);
    layer3_outputs(2425) <= (layer2_outputs(1563)) and not (layer2_outputs(6113));
    layer3_outputs(2426) <= (layer2_outputs(3455)) or (layer2_outputs(450));
    layer3_outputs(2427) <= not(layer2_outputs(4673));
    layer3_outputs(2428) <= not(layer2_outputs(3812)) or (layer2_outputs(616));
    layer3_outputs(2429) <= (layer2_outputs(1081)) and not (layer2_outputs(160));
    layer3_outputs(2430) <= not((layer2_outputs(803)) xor (layer2_outputs(2301)));
    layer3_outputs(2431) <= (layer2_outputs(2199)) or (layer2_outputs(5004));
    layer3_outputs(2432) <= not(layer2_outputs(3807));
    layer3_outputs(2433) <= '1';
    layer3_outputs(2434) <= (layer2_outputs(4679)) and not (layer2_outputs(645));
    layer3_outputs(2435) <= (layer2_outputs(7515)) and (layer2_outputs(2451));
    layer3_outputs(2436) <= layer2_outputs(5295);
    layer3_outputs(2437) <= layer2_outputs(6150);
    layer3_outputs(2438) <= '1';
    layer3_outputs(2439) <= not(layer2_outputs(3321)) or (layer2_outputs(1753));
    layer3_outputs(2440) <= not(layer2_outputs(4407));
    layer3_outputs(2441) <= layer2_outputs(1353);
    layer3_outputs(2442) <= (layer2_outputs(2425)) and not (layer2_outputs(276));
    layer3_outputs(2443) <= not(layer2_outputs(361));
    layer3_outputs(2444) <= layer2_outputs(6334);
    layer3_outputs(2445) <= '0';
    layer3_outputs(2446) <= not(layer2_outputs(666));
    layer3_outputs(2447) <= not(layer2_outputs(612));
    layer3_outputs(2448) <= (layer2_outputs(7568)) or (layer2_outputs(5931));
    layer3_outputs(2449) <= (layer2_outputs(2289)) or (layer2_outputs(6333));
    layer3_outputs(2450) <= layer2_outputs(416);
    layer3_outputs(2451) <= (layer2_outputs(4890)) or (layer2_outputs(302));
    layer3_outputs(2452) <= layer2_outputs(576);
    layer3_outputs(2453) <= not((layer2_outputs(2113)) or (layer2_outputs(6838)));
    layer3_outputs(2454) <= (layer2_outputs(1751)) or (layer2_outputs(3271));
    layer3_outputs(2455) <= not(layer2_outputs(3540)) or (layer2_outputs(3461));
    layer3_outputs(2456) <= (layer2_outputs(2705)) and (layer2_outputs(1936));
    layer3_outputs(2457) <= '1';
    layer3_outputs(2458) <= not((layer2_outputs(5708)) or (layer2_outputs(4634)));
    layer3_outputs(2459) <= (layer2_outputs(6677)) xor (layer2_outputs(4677));
    layer3_outputs(2460) <= not(layer2_outputs(1053));
    layer3_outputs(2461) <= (layer2_outputs(1778)) and not (layer2_outputs(5377));
    layer3_outputs(2462) <= not(layer2_outputs(11)) or (layer2_outputs(2968));
    layer3_outputs(2463) <= '0';
    layer3_outputs(2464) <= layer2_outputs(3415);
    layer3_outputs(2465) <= layer2_outputs(493);
    layer3_outputs(2466) <= '0';
    layer3_outputs(2467) <= not(layer2_outputs(1477));
    layer3_outputs(2468) <= not(layer2_outputs(5981));
    layer3_outputs(2469) <= not(layer2_outputs(7392));
    layer3_outputs(2470) <= not((layer2_outputs(7201)) xor (layer2_outputs(6424)));
    layer3_outputs(2471) <= (layer2_outputs(4085)) or (layer2_outputs(3394));
    layer3_outputs(2472) <= layer2_outputs(3091);
    layer3_outputs(2473) <= (layer2_outputs(2671)) and (layer2_outputs(519));
    layer3_outputs(2474) <= (layer2_outputs(5203)) and not (layer2_outputs(4367));
    layer3_outputs(2475) <= (layer2_outputs(2171)) and (layer2_outputs(6854));
    layer3_outputs(2476) <= (layer2_outputs(5320)) and not (layer2_outputs(2232));
    layer3_outputs(2477) <= not(layer2_outputs(7528)) or (layer2_outputs(670));
    layer3_outputs(2478) <= not(layer2_outputs(3409));
    layer3_outputs(2479) <= layer2_outputs(1496);
    layer3_outputs(2480) <= (layer2_outputs(891)) and (layer2_outputs(35));
    layer3_outputs(2481) <= (layer2_outputs(2035)) and (layer2_outputs(2447));
    layer3_outputs(2482) <= (layer2_outputs(6230)) and not (layer2_outputs(4310));
    layer3_outputs(2483) <= not((layer2_outputs(4368)) and (layer2_outputs(1877)));
    layer3_outputs(2484) <= not(layer2_outputs(60));
    layer3_outputs(2485) <= not((layer2_outputs(1561)) xor (layer2_outputs(2048)));
    layer3_outputs(2486) <= layer2_outputs(5366);
    layer3_outputs(2487) <= not(layer2_outputs(2850));
    layer3_outputs(2488) <= (layer2_outputs(5506)) or (layer2_outputs(4762));
    layer3_outputs(2489) <= '1';
    layer3_outputs(2490) <= (layer2_outputs(5772)) or (layer2_outputs(5889));
    layer3_outputs(2491) <= not((layer2_outputs(102)) and (layer2_outputs(6397)));
    layer3_outputs(2492) <= layer2_outputs(4417);
    layer3_outputs(2493) <= not(layer2_outputs(5102));
    layer3_outputs(2494) <= not(layer2_outputs(3966)) or (layer2_outputs(2058));
    layer3_outputs(2495) <= not((layer2_outputs(6291)) or (layer2_outputs(3842)));
    layer3_outputs(2496) <= not(layer2_outputs(6155));
    layer3_outputs(2497) <= not(layer2_outputs(2105)) or (layer2_outputs(6578));
    layer3_outputs(2498) <= layer2_outputs(2074);
    layer3_outputs(2499) <= layer2_outputs(5950);
    layer3_outputs(2500) <= (layer2_outputs(5592)) and not (layer2_outputs(6157));
    layer3_outputs(2501) <= layer2_outputs(2935);
    layer3_outputs(2502) <= layer2_outputs(2297);
    layer3_outputs(2503) <= not(layer2_outputs(6403)) or (layer2_outputs(348));
    layer3_outputs(2504) <= layer2_outputs(3681);
    layer3_outputs(2505) <= layer2_outputs(5232);
    layer3_outputs(2506) <= not(layer2_outputs(6862)) or (layer2_outputs(252));
    layer3_outputs(2507) <= not((layer2_outputs(3637)) or (layer2_outputs(6585)));
    layer3_outputs(2508) <= layer2_outputs(2753);
    layer3_outputs(2509) <= not(layer2_outputs(922));
    layer3_outputs(2510) <= not(layer2_outputs(708)) or (layer2_outputs(5346));
    layer3_outputs(2511) <= (layer2_outputs(6904)) and not (layer2_outputs(6168));
    layer3_outputs(2512) <= layer2_outputs(3442);
    layer3_outputs(2513) <= layer2_outputs(2164);
    layer3_outputs(2514) <= not(layer2_outputs(447));
    layer3_outputs(2515) <= (layer2_outputs(874)) and not (layer2_outputs(2150));
    layer3_outputs(2516) <= layer2_outputs(6839);
    layer3_outputs(2517) <= not((layer2_outputs(1481)) or (layer2_outputs(6019)));
    layer3_outputs(2518) <= not(layer2_outputs(6118));
    layer3_outputs(2519) <= not(layer2_outputs(4016)) or (layer2_outputs(1590));
    layer3_outputs(2520) <= not(layer2_outputs(1948)) or (layer2_outputs(279));
    layer3_outputs(2521) <= layer2_outputs(1766);
    layer3_outputs(2522) <= (layer2_outputs(4145)) xor (layer2_outputs(6713));
    layer3_outputs(2523) <= not(layer2_outputs(3773));
    layer3_outputs(2524) <= (layer2_outputs(4993)) xor (layer2_outputs(4880));
    layer3_outputs(2525) <= not((layer2_outputs(6105)) xor (layer2_outputs(62)));
    layer3_outputs(2526) <= not((layer2_outputs(608)) or (layer2_outputs(4641)));
    layer3_outputs(2527) <= not(layer2_outputs(3086));
    layer3_outputs(2528) <= '0';
    layer3_outputs(2529) <= (layer2_outputs(6126)) and (layer2_outputs(5488));
    layer3_outputs(2530) <= (layer2_outputs(2485)) and (layer2_outputs(7023));
    layer3_outputs(2531) <= layer2_outputs(4922);
    layer3_outputs(2532) <= layer2_outputs(4940);
    layer3_outputs(2533) <= not(layer2_outputs(6972));
    layer3_outputs(2534) <= (layer2_outputs(5035)) and (layer2_outputs(1071));
    layer3_outputs(2535) <= not(layer2_outputs(1579));
    layer3_outputs(2536) <= not(layer2_outputs(2873));
    layer3_outputs(2537) <= not(layer2_outputs(5629));
    layer3_outputs(2538) <= (layer2_outputs(5724)) and (layer2_outputs(1362));
    layer3_outputs(2539) <= layer2_outputs(6208);
    layer3_outputs(2540) <= not(layer2_outputs(498));
    layer3_outputs(2541) <= not((layer2_outputs(944)) and (layer2_outputs(7007)));
    layer3_outputs(2542) <= (layer2_outputs(6847)) and not (layer2_outputs(5679));
    layer3_outputs(2543) <= '0';
    layer3_outputs(2544) <= not(layer2_outputs(182));
    layer3_outputs(2545) <= '0';
    layer3_outputs(2546) <= '0';
    layer3_outputs(2547) <= not((layer2_outputs(335)) or (layer2_outputs(426)));
    layer3_outputs(2548) <= layer2_outputs(4101);
    layer3_outputs(2549) <= layer2_outputs(1757);
    layer3_outputs(2550) <= layer2_outputs(5594);
    layer3_outputs(2551) <= layer2_outputs(1955);
    layer3_outputs(2552) <= not((layer2_outputs(7329)) or (layer2_outputs(1890)));
    layer3_outputs(2553) <= layer2_outputs(1795);
    layer3_outputs(2554) <= not(layer2_outputs(5821));
    layer3_outputs(2555) <= not((layer2_outputs(5963)) or (layer2_outputs(1672)));
    layer3_outputs(2556) <= not(layer2_outputs(3308)) or (layer2_outputs(115));
    layer3_outputs(2557) <= (layer2_outputs(5333)) and not (layer2_outputs(7170));
    layer3_outputs(2558) <= layer2_outputs(95);
    layer3_outputs(2559) <= (layer2_outputs(7114)) and not (layer2_outputs(7624));
    layer3_outputs(2560) <= not((layer2_outputs(7221)) and (layer2_outputs(7334)));
    layer3_outputs(2561) <= not((layer2_outputs(1723)) or (layer2_outputs(3970)));
    layer3_outputs(2562) <= layer2_outputs(3810);
    layer3_outputs(2563) <= layer2_outputs(593);
    layer3_outputs(2564) <= not((layer2_outputs(466)) and (layer2_outputs(3875)));
    layer3_outputs(2565) <= layer2_outputs(6075);
    layer3_outputs(2566) <= not((layer2_outputs(293)) or (layer2_outputs(5391)));
    layer3_outputs(2567) <= not(layer2_outputs(5673)) or (layer2_outputs(2197));
    layer3_outputs(2568) <= not(layer2_outputs(3767)) or (layer2_outputs(1747));
    layer3_outputs(2569) <= layer2_outputs(2529);
    layer3_outputs(2570) <= not(layer2_outputs(1400));
    layer3_outputs(2571) <= not(layer2_outputs(1539));
    layer3_outputs(2572) <= not(layer2_outputs(3992)) or (layer2_outputs(1591));
    layer3_outputs(2573) <= not(layer2_outputs(5655));
    layer3_outputs(2574) <= layer2_outputs(4234);
    layer3_outputs(2575) <= layer2_outputs(266);
    layer3_outputs(2576) <= (layer2_outputs(5995)) and not (layer2_outputs(2162));
    layer3_outputs(2577) <= (layer2_outputs(2061)) xor (layer2_outputs(6604));
    layer3_outputs(2578) <= not((layer2_outputs(6588)) xor (layer2_outputs(1173)));
    layer3_outputs(2579) <= not(layer2_outputs(5519));
    layer3_outputs(2580) <= layer2_outputs(3637);
    layer3_outputs(2581) <= not(layer2_outputs(463)) or (layer2_outputs(839));
    layer3_outputs(2582) <= not(layer2_outputs(6194));
    layer3_outputs(2583) <= (layer2_outputs(5273)) and not (layer2_outputs(2653));
    layer3_outputs(2584) <= layer2_outputs(2358);
    layer3_outputs(2585) <= not(layer2_outputs(2391));
    layer3_outputs(2586) <= layer2_outputs(2491);
    layer3_outputs(2587) <= not((layer2_outputs(4311)) or (layer2_outputs(1519)));
    layer3_outputs(2588) <= (layer2_outputs(5331)) and not (layer2_outputs(883));
    layer3_outputs(2589) <= not(layer2_outputs(3856));
    layer3_outputs(2590) <= not((layer2_outputs(4659)) or (layer2_outputs(6953)));
    layer3_outputs(2591) <= (layer2_outputs(6255)) and (layer2_outputs(7533));
    layer3_outputs(2592) <= not((layer2_outputs(356)) xor (layer2_outputs(6588)));
    layer3_outputs(2593) <= '0';
    layer3_outputs(2594) <= layer2_outputs(1775);
    layer3_outputs(2595) <= not(layer2_outputs(6856));
    layer3_outputs(2596) <= layer2_outputs(3633);
    layer3_outputs(2597) <= (layer2_outputs(7610)) or (layer2_outputs(3089));
    layer3_outputs(2598) <= (layer2_outputs(2776)) and not (layer2_outputs(3815));
    layer3_outputs(2599) <= (layer2_outputs(7430)) and (layer2_outputs(4623));
    layer3_outputs(2600) <= (layer2_outputs(2624)) or (layer2_outputs(5267));
    layer3_outputs(2601) <= not(layer2_outputs(3066));
    layer3_outputs(2602) <= layer2_outputs(1250);
    layer3_outputs(2603) <= not(layer2_outputs(2544));
    layer3_outputs(2604) <= not((layer2_outputs(256)) or (layer2_outputs(1444)));
    layer3_outputs(2605) <= not(layer2_outputs(4941)) or (layer2_outputs(5237));
    layer3_outputs(2606) <= not(layer2_outputs(5871)) or (layer2_outputs(7066));
    layer3_outputs(2607) <= (layer2_outputs(5275)) and (layer2_outputs(2780));
    layer3_outputs(2608) <= not(layer2_outputs(2229));
    layer3_outputs(2609) <= not(layer2_outputs(216));
    layer3_outputs(2610) <= not(layer2_outputs(6166));
    layer3_outputs(2611) <= not(layer2_outputs(226));
    layer3_outputs(2612) <= not((layer2_outputs(307)) or (layer2_outputs(2328)));
    layer3_outputs(2613) <= '0';
    layer3_outputs(2614) <= (layer2_outputs(6270)) and not (layer2_outputs(7451));
    layer3_outputs(2615) <= not((layer2_outputs(6030)) and (layer2_outputs(3817)));
    layer3_outputs(2616) <= layer2_outputs(810);
    layer3_outputs(2617) <= not(layer2_outputs(5731));
    layer3_outputs(2618) <= not((layer2_outputs(472)) and (layer2_outputs(4072)));
    layer3_outputs(2619) <= not((layer2_outputs(2066)) xor (layer2_outputs(6592)));
    layer3_outputs(2620) <= layer2_outputs(2672);
    layer3_outputs(2621) <= not(layer2_outputs(5135));
    layer3_outputs(2622) <= not(layer2_outputs(632));
    layer3_outputs(2623) <= layer2_outputs(4082);
    layer3_outputs(2624) <= not(layer2_outputs(5716));
    layer3_outputs(2625) <= '0';
    layer3_outputs(2626) <= not((layer2_outputs(5997)) or (layer2_outputs(3560)));
    layer3_outputs(2627) <= layer2_outputs(4374);
    layer3_outputs(2628) <= layer2_outputs(4912);
    layer3_outputs(2629) <= layer2_outputs(150);
    layer3_outputs(2630) <= not((layer2_outputs(6867)) and (layer2_outputs(3170)));
    layer3_outputs(2631) <= not(layer2_outputs(5660)) or (layer2_outputs(633));
    layer3_outputs(2632) <= layer2_outputs(1219);
    layer3_outputs(2633) <= layer2_outputs(3611);
    layer3_outputs(2634) <= layer2_outputs(2266);
    layer3_outputs(2635) <= not((layer2_outputs(4211)) and (layer2_outputs(6347)));
    layer3_outputs(2636) <= layer2_outputs(2271);
    layer3_outputs(2637) <= '1';
    layer3_outputs(2638) <= not((layer2_outputs(6840)) and (layer2_outputs(4562)));
    layer3_outputs(2639) <= not(layer2_outputs(3184)) or (layer2_outputs(838));
    layer3_outputs(2640) <= layer2_outputs(3947);
    layer3_outputs(2641) <= layer2_outputs(6693);
    layer3_outputs(2642) <= not(layer2_outputs(7579));
    layer3_outputs(2643) <= not((layer2_outputs(6359)) or (layer2_outputs(35)));
    layer3_outputs(2644) <= not(layer2_outputs(745));
    layer3_outputs(2645) <= (layer2_outputs(4656)) and not (layer2_outputs(1809));
    layer3_outputs(2646) <= not(layer2_outputs(2931));
    layer3_outputs(2647) <= layer2_outputs(3847);
    layer3_outputs(2648) <= not(layer2_outputs(4088));
    layer3_outputs(2649) <= layer2_outputs(2006);
    layer3_outputs(2650) <= not(layer2_outputs(1040));
    layer3_outputs(2651) <= not(layer2_outputs(7266)) or (layer2_outputs(3376));
    layer3_outputs(2652) <= not(layer2_outputs(3758)) or (layer2_outputs(159));
    layer3_outputs(2653) <= (layer2_outputs(4754)) and not (layer2_outputs(5163));
    layer3_outputs(2654) <= not(layer2_outputs(5974));
    layer3_outputs(2655) <= layer2_outputs(290);
    layer3_outputs(2656) <= layer2_outputs(424);
    layer3_outputs(2657) <= (layer2_outputs(6739)) and not (layer2_outputs(6437));
    layer3_outputs(2658) <= layer2_outputs(6086);
    layer3_outputs(2659) <= not(layer2_outputs(3764));
    layer3_outputs(2660) <= not((layer2_outputs(3137)) and (layer2_outputs(5827)));
    layer3_outputs(2661) <= layer2_outputs(2546);
    layer3_outputs(2662) <= (layer2_outputs(5917)) and (layer2_outputs(2520));
    layer3_outputs(2663) <= (layer2_outputs(7090)) or (layer2_outputs(306));
    layer3_outputs(2664) <= (layer2_outputs(275)) xor (layer2_outputs(1674));
    layer3_outputs(2665) <= (layer2_outputs(4589)) and not (layer2_outputs(1788));
    layer3_outputs(2666) <= layer2_outputs(617);
    layer3_outputs(2667) <= (layer2_outputs(7415)) and (layer2_outputs(5501));
    layer3_outputs(2668) <= not(layer2_outputs(7494));
    layer3_outputs(2669) <= (layer2_outputs(4238)) and not (layer2_outputs(4464));
    layer3_outputs(2670) <= not(layer2_outputs(4289));
    layer3_outputs(2671) <= not(layer2_outputs(718)) or (layer2_outputs(6216));
    layer3_outputs(2672) <= (layer2_outputs(7623)) and not (layer2_outputs(5669));
    layer3_outputs(2673) <= (layer2_outputs(5811)) and (layer2_outputs(3720));
    layer3_outputs(2674) <= not(layer2_outputs(6728));
    layer3_outputs(2675) <= (layer2_outputs(303)) xor (layer2_outputs(2900));
    layer3_outputs(2676) <= (layer2_outputs(6680)) and not (layer2_outputs(5824));
    layer3_outputs(2677) <= layer2_outputs(5188);
    layer3_outputs(2678) <= not(layer2_outputs(5051)) or (layer2_outputs(2925));
    layer3_outputs(2679) <= not(layer2_outputs(2473));
    layer3_outputs(2680) <= not((layer2_outputs(2245)) and (layer2_outputs(1852)));
    layer3_outputs(2681) <= not((layer2_outputs(5721)) or (layer2_outputs(3851)));
    layer3_outputs(2682) <= layer2_outputs(1507);
    layer3_outputs(2683) <= not(layer2_outputs(5508)) or (layer2_outputs(1535));
    layer3_outputs(2684) <= not((layer2_outputs(547)) xor (layer2_outputs(4297)));
    layer3_outputs(2685) <= not(layer2_outputs(3112));
    layer3_outputs(2686) <= not((layer2_outputs(7015)) and (layer2_outputs(7004)));
    layer3_outputs(2687) <= not(layer2_outputs(7582));
    layer3_outputs(2688) <= not(layer2_outputs(1073));
    layer3_outputs(2689) <= (layer2_outputs(1219)) or (layer2_outputs(7162));
    layer3_outputs(2690) <= not((layer2_outputs(3687)) or (layer2_outputs(3508)));
    layer3_outputs(2691) <= not(layer2_outputs(6129)) or (layer2_outputs(6086));
    layer3_outputs(2692) <= layer2_outputs(4957);
    layer3_outputs(2693) <= not(layer2_outputs(6232));
    layer3_outputs(2694) <= not(layer2_outputs(3396)) or (layer2_outputs(3682));
    layer3_outputs(2695) <= (layer2_outputs(5189)) and (layer2_outputs(3521));
    layer3_outputs(2696) <= layer2_outputs(6458);
    layer3_outputs(2697) <= not(layer2_outputs(3793)) or (layer2_outputs(1020));
    layer3_outputs(2698) <= (layer2_outputs(2644)) and not (layer2_outputs(4731));
    layer3_outputs(2699) <= (layer2_outputs(4482)) or (layer2_outputs(6761));
    layer3_outputs(2700) <= (layer2_outputs(4057)) and not (layer2_outputs(2427));
    layer3_outputs(2701) <= '0';
    layer3_outputs(2702) <= not((layer2_outputs(5311)) or (layer2_outputs(580)));
    layer3_outputs(2703) <= (layer2_outputs(3891)) or (layer2_outputs(6896));
    layer3_outputs(2704) <= (layer2_outputs(3524)) xor (layer2_outputs(1410));
    layer3_outputs(2705) <= not((layer2_outputs(1426)) or (layer2_outputs(2146)));
    layer3_outputs(2706) <= layer2_outputs(6039);
    layer3_outputs(2707) <= not((layer2_outputs(5210)) and (layer2_outputs(3170)));
    layer3_outputs(2708) <= not(layer2_outputs(3334));
    layer3_outputs(2709) <= not((layer2_outputs(1174)) or (layer2_outputs(6154)));
    layer3_outputs(2710) <= not(layer2_outputs(6795));
    layer3_outputs(2711) <= (layer2_outputs(6457)) and not (layer2_outputs(205));
    layer3_outputs(2712) <= '0';
    layer3_outputs(2713) <= not(layer2_outputs(7313));
    layer3_outputs(2714) <= not((layer2_outputs(180)) and (layer2_outputs(6314)));
    layer3_outputs(2715) <= (layer2_outputs(4553)) or (layer2_outputs(3896));
    layer3_outputs(2716) <= layer2_outputs(5634);
    layer3_outputs(2717) <= (layer2_outputs(4257)) and not (layer2_outputs(6666));
    layer3_outputs(2718) <= not((layer2_outputs(5955)) and (layer2_outputs(6822)));
    layer3_outputs(2719) <= not(layer2_outputs(5395));
    layer3_outputs(2720) <= layer2_outputs(1578);
    layer3_outputs(2721) <= not(layer2_outputs(4919)) or (layer2_outputs(2632));
    layer3_outputs(2722) <= layer2_outputs(6315);
    layer3_outputs(2723) <= layer2_outputs(184);
    layer3_outputs(2724) <= not(layer2_outputs(1673)) or (layer2_outputs(1856));
    layer3_outputs(2725) <= (layer2_outputs(3385)) and not (layer2_outputs(1730));
    layer3_outputs(2726) <= '1';
    layer3_outputs(2727) <= not((layer2_outputs(2524)) or (layer2_outputs(1614)));
    layer3_outputs(2728) <= not(layer2_outputs(3270));
    layer3_outputs(2729) <= (layer2_outputs(6374)) and (layer2_outputs(3020));
    layer3_outputs(2730) <= not(layer2_outputs(262)) or (layer2_outputs(3311));
    layer3_outputs(2731) <= not(layer2_outputs(5129)) or (layer2_outputs(6526));
    layer3_outputs(2732) <= (layer2_outputs(5177)) and (layer2_outputs(3574));
    layer3_outputs(2733) <= not(layer2_outputs(2614));
    layer3_outputs(2734) <= not(layer2_outputs(3124));
    layer3_outputs(2735) <= not(layer2_outputs(1643));
    layer3_outputs(2736) <= (layer2_outputs(5520)) and (layer2_outputs(1719));
    layer3_outputs(2737) <= (layer2_outputs(1450)) and not (layer2_outputs(813));
    layer3_outputs(2738) <= layer2_outputs(2111);
    layer3_outputs(2739) <= (layer2_outputs(5718)) and (layer2_outputs(5698));
    layer3_outputs(2740) <= not(layer2_outputs(3885));
    layer3_outputs(2741) <= (layer2_outputs(2170)) and (layer2_outputs(5155));
    layer3_outputs(2742) <= (layer2_outputs(2312)) xor (layer2_outputs(3085));
    layer3_outputs(2743) <= layer2_outputs(4315);
    layer3_outputs(2744) <= not(layer2_outputs(3887));
    layer3_outputs(2745) <= not(layer2_outputs(3516)) or (layer2_outputs(6973));
    layer3_outputs(2746) <= (layer2_outputs(873)) and (layer2_outputs(5664));
    layer3_outputs(2747) <= not(layer2_outputs(5512));
    layer3_outputs(2748) <= not((layer2_outputs(1636)) or (layer2_outputs(5353)));
    layer3_outputs(2749) <= not(layer2_outputs(5536));
    layer3_outputs(2750) <= (layer2_outputs(4885)) and (layer2_outputs(2674));
    layer3_outputs(2751) <= not(layer2_outputs(4397));
    layer3_outputs(2752) <= not(layer2_outputs(6806));
    layer3_outputs(2753) <= (layer2_outputs(2556)) and not (layer2_outputs(6197));
    layer3_outputs(2754) <= not(layer2_outputs(6107)) or (layer2_outputs(6869));
    layer3_outputs(2755) <= layer2_outputs(6629);
    layer3_outputs(2756) <= layer2_outputs(3764);
    layer3_outputs(2757) <= not(layer2_outputs(2374)) or (layer2_outputs(4463));
    layer3_outputs(2758) <= not(layer2_outputs(3366));
    layer3_outputs(2759) <= (layer2_outputs(5349)) and (layer2_outputs(5975));
    layer3_outputs(2760) <= (layer2_outputs(3166)) xor (layer2_outputs(6400));
    layer3_outputs(2761) <= not(layer2_outputs(6538));
    layer3_outputs(2762) <= (layer2_outputs(2200)) and (layer2_outputs(5564));
    layer3_outputs(2763) <= layer2_outputs(1977);
    layer3_outputs(2764) <= (layer2_outputs(6451)) and not (layer2_outputs(243));
    layer3_outputs(2765) <= layer2_outputs(6790);
    layer3_outputs(2766) <= not(layer2_outputs(4861)) or (layer2_outputs(2226));
    layer3_outputs(2767) <= (layer2_outputs(4378)) and not (layer2_outputs(2088));
    layer3_outputs(2768) <= not((layer2_outputs(6961)) or (layer2_outputs(4923)));
    layer3_outputs(2769) <= not(layer2_outputs(3782));
    layer3_outputs(2770) <= (layer2_outputs(1451)) xor (layer2_outputs(4644));
    layer3_outputs(2771) <= layer2_outputs(5357);
    layer3_outputs(2772) <= (layer2_outputs(998)) and not (layer2_outputs(2548));
    layer3_outputs(2773) <= (layer2_outputs(7679)) or (layer2_outputs(1846));
    layer3_outputs(2774) <= layer2_outputs(5074);
    layer3_outputs(2775) <= not((layer2_outputs(7392)) and (layer2_outputs(7475)));
    layer3_outputs(2776) <= layer2_outputs(6552);
    layer3_outputs(2777) <= not(layer2_outputs(801)) or (layer2_outputs(2430));
    layer3_outputs(2778) <= (layer2_outputs(881)) xor (layer2_outputs(7367));
    layer3_outputs(2779) <= not(layer2_outputs(1923));
    layer3_outputs(2780) <= layer2_outputs(351);
    layer3_outputs(2781) <= not(layer2_outputs(1050));
    layer3_outputs(2782) <= (layer2_outputs(2636)) and not (layer2_outputs(2144));
    layer3_outputs(2783) <= '1';
    layer3_outputs(2784) <= not(layer2_outputs(3577));
    layer3_outputs(2785) <= (layer2_outputs(3008)) or (layer2_outputs(3157));
    layer3_outputs(2786) <= not(layer2_outputs(7387));
    layer3_outputs(2787) <= not(layer2_outputs(1566));
    layer3_outputs(2788) <= layer2_outputs(533);
    layer3_outputs(2789) <= not(layer2_outputs(4217));
    layer3_outputs(2790) <= (layer2_outputs(3084)) or (layer2_outputs(61));
    layer3_outputs(2791) <= (layer2_outputs(618)) xor (layer2_outputs(4564));
    layer3_outputs(2792) <= not(layer2_outputs(7363));
    layer3_outputs(2793) <= not(layer2_outputs(6154));
    layer3_outputs(2794) <= not(layer2_outputs(6549));
    layer3_outputs(2795) <= not(layer2_outputs(3957));
    layer3_outputs(2796) <= not((layer2_outputs(3731)) and (layer2_outputs(6052)));
    layer3_outputs(2797) <= not(layer2_outputs(1290)) or (layer2_outputs(6521));
    layer3_outputs(2798) <= '0';
    layer3_outputs(2799) <= not(layer2_outputs(3399));
    layer3_outputs(2800) <= not(layer2_outputs(5139)) or (layer2_outputs(3446));
    layer3_outputs(2801) <= not(layer2_outputs(2201));
    layer3_outputs(2802) <= not(layer2_outputs(5799));
    layer3_outputs(2803) <= (layer2_outputs(1897)) or (layer2_outputs(3030));
    layer3_outputs(2804) <= (layer2_outputs(316)) or (layer2_outputs(1258));
    layer3_outputs(2805) <= layer2_outputs(5313);
    layer3_outputs(2806) <= layer2_outputs(570);
    layer3_outputs(2807) <= layer2_outputs(2744);
    layer3_outputs(2808) <= not(layer2_outputs(3264));
    layer3_outputs(2809) <= layer2_outputs(3732);
    layer3_outputs(2810) <= layer2_outputs(5778);
    layer3_outputs(2811) <= not((layer2_outputs(5440)) or (layer2_outputs(607)));
    layer3_outputs(2812) <= not((layer2_outputs(6317)) or (layer2_outputs(1713)));
    layer3_outputs(2813) <= (layer2_outputs(4414)) and (layer2_outputs(414));
    layer3_outputs(2814) <= layer2_outputs(500);
    layer3_outputs(2815) <= not(layer2_outputs(843));
    layer3_outputs(2816) <= layer2_outputs(2498);
    layer3_outputs(2817) <= not(layer2_outputs(560));
    layer3_outputs(2818) <= not(layer2_outputs(5067)) or (layer2_outputs(5958));
    layer3_outputs(2819) <= not(layer2_outputs(4261));
    layer3_outputs(2820) <= layer2_outputs(852);
    layer3_outputs(2821) <= not(layer2_outputs(479));
    layer3_outputs(2822) <= not((layer2_outputs(7052)) and (layer2_outputs(4829)));
    layer3_outputs(2823) <= not((layer2_outputs(1094)) or (layer2_outputs(45)));
    layer3_outputs(2824) <= layer2_outputs(6714);
    layer3_outputs(2825) <= not(layer2_outputs(2622)) or (layer2_outputs(171));
    layer3_outputs(2826) <= layer2_outputs(4729);
    layer3_outputs(2827) <= (layer2_outputs(5652)) and (layer2_outputs(4678));
    layer3_outputs(2828) <= (layer2_outputs(3609)) and not (layer2_outputs(4698));
    layer3_outputs(2829) <= layer2_outputs(2323);
    layer3_outputs(2830) <= layer2_outputs(1164);
    layer3_outputs(2831) <= not(layer2_outputs(6593));
    layer3_outputs(2832) <= (layer2_outputs(1782)) and not (layer2_outputs(6222));
    layer3_outputs(2833) <= (layer2_outputs(2089)) and not (layer2_outputs(2720));
    layer3_outputs(2834) <= (layer2_outputs(1663)) or (layer2_outputs(2021));
    layer3_outputs(2835) <= (layer2_outputs(4645)) and (layer2_outputs(6576));
    layer3_outputs(2836) <= (layer2_outputs(397)) xor (layer2_outputs(4567));
    layer3_outputs(2837) <= layer2_outputs(7523);
    layer3_outputs(2838) <= layer2_outputs(6569);
    layer3_outputs(2839) <= not((layer2_outputs(5581)) and (layer2_outputs(5851)));
    layer3_outputs(2840) <= not(layer2_outputs(6262)) or (layer2_outputs(4419));
    layer3_outputs(2841) <= not((layer2_outputs(894)) or (layer2_outputs(3243)));
    layer3_outputs(2842) <= layer2_outputs(2379);
    layer3_outputs(2843) <= layer2_outputs(4106);
    layer3_outputs(2844) <= not((layer2_outputs(6271)) or (layer2_outputs(3721)));
    layer3_outputs(2845) <= (layer2_outputs(591)) and not (layer2_outputs(5876));
    layer3_outputs(2846) <= not((layer2_outputs(4830)) and (layer2_outputs(3699)));
    layer3_outputs(2847) <= (layer2_outputs(4844)) and not (layer2_outputs(1492));
    layer3_outputs(2848) <= not(layer2_outputs(5587)) or (layer2_outputs(6046));
    layer3_outputs(2849) <= not(layer2_outputs(6767));
    layer3_outputs(2850) <= not((layer2_outputs(1264)) and (layer2_outputs(3063)));
    layer3_outputs(2851) <= (layer2_outputs(7155)) and not (layer2_outputs(5672));
    layer3_outputs(2852) <= not(layer2_outputs(6183)) or (layer2_outputs(733));
    layer3_outputs(2853) <= '1';
    layer3_outputs(2854) <= not(layer2_outputs(3600)) or (layer2_outputs(304));
    layer3_outputs(2855) <= not(layer2_outputs(3435));
    layer3_outputs(2856) <= layer2_outputs(2451);
    layer3_outputs(2857) <= not((layer2_outputs(3282)) or (layer2_outputs(6766)));
    layer3_outputs(2858) <= layer2_outputs(5190);
    layer3_outputs(2859) <= not((layer2_outputs(5835)) xor (layer2_outputs(5554)));
    layer3_outputs(2860) <= (layer2_outputs(7525)) and not (layer2_outputs(1710));
    layer3_outputs(2861) <= (layer2_outputs(5600)) and not (layer2_outputs(641));
    layer3_outputs(2862) <= not((layer2_outputs(1660)) or (layer2_outputs(5725)));
    layer3_outputs(2863) <= (layer2_outputs(6337)) and not (layer2_outputs(662));
    layer3_outputs(2864) <= (layer2_outputs(5819)) and not (layer2_outputs(3104));
    layer3_outputs(2865) <= not(layer2_outputs(904));
    layer3_outputs(2866) <= layer2_outputs(6583);
    layer3_outputs(2867) <= not(layer2_outputs(47));
    layer3_outputs(2868) <= (layer2_outputs(6742)) and (layer2_outputs(6589));
    layer3_outputs(2869) <= not(layer2_outputs(810)) or (layer2_outputs(1413));
    layer3_outputs(2870) <= (layer2_outputs(6385)) or (layer2_outputs(7488));
    layer3_outputs(2871) <= not(layer2_outputs(6878));
    layer3_outputs(2872) <= not(layer2_outputs(7433));
    layer3_outputs(2873) <= not(layer2_outputs(6687));
    layer3_outputs(2874) <= (layer2_outputs(3059)) and not (layer2_outputs(6934));
    layer3_outputs(2875) <= not(layer2_outputs(6428));
    layer3_outputs(2876) <= (layer2_outputs(3032)) and not (layer2_outputs(1828));
    layer3_outputs(2877) <= layer2_outputs(5702);
    layer3_outputs(2878) <= not((layer2_outputs(5875)) and (layer2_outputs(6833)));
    layer3_outputs(2879) <= (layer2_outputs(1613)) and (layer2_outputs(944));
    layer3_outputs(2880) <= (layer2_outputs(5269)) and not (layer2_outputs(710));
    layer3_outputs(2881) <= not((layer2_outputs(7525)) and (layer2_outputs(7611)));
    layer3_outputs(2882) <= '1';
    layer3_outputs(2883) <= layer2_outputs(5433);
    layer3_outputs(2884) <= (layer2_outputs(1341)) and not (layer2_outputs(3941));
    layer3_outputs(2885) <= '0';
    layer3_outputs(2886) <= not(layer2_outputs(5706));
    layer3_outputs(2887) <= layer2_outputs(2903);
    layer3_outputs(2888) <= not(layer2_outputs(4724)) or (layer2_outputs(5904));
    layer3_outputs(2889) <= not(layer2_outputs(7608));
    layer3_outputs(2890) <= not(layer2_outputs(2063)) or (layer2_outputs(7276));
    layer3_outputs(2891) <= not(layer2_outputs(967));
    layer3_outputs(2892) <= not(layer2_outputs(3706));
    layer3_outputs(2893) <= not(layer2_outputs(4706));
    layer3_outputs(2894) <= '1';
    layer3_outputs(2895) <= not(layer2_outputs(5718));
    layer3_outputs(2896) <= not(layer2_outputs(765));
    layer3_outputs(2897) <= not((layer2_outputs(3960)) and (layer2_outputs(5545)));
    layer3_outputs(2898) <= layer2_outputs(3026);
    layer3_outputs(2899) <= not(layer2_outputs(6486));
    layer3_outputs(2900) <= not(layer2_outputs(214));
    layer3_outputs(2901) <= layer2_outputs(6900);
    layer3_outputs(2902) <= layer2_outputs(5033);
    layer3_outputs(2903) <= not(layer2_outputs(6818));
    layer3_outputs(2904) <= not(layer2_outputs(5001));
    layer3_outputs(2905) <= layer2_outputs(4741);
    layer3_outputs(2906) <= not(layer2_outputs(6789));
    layer3_outputs(2907) <= (layer2_outputs(3426)) and not (layer2_outputs(4128));
    layer3_outputs(2908) <= (layer2_outputs(6332)) and (layer2_outputs(5349));
    layer3_outputs(2909) <= (layer2_outputs(2822)) and (layer2_outputs(6483));
    layer3_outputs(2910) <= not((layer2_outputs(5915)) or (layer2_outputs(427)));
    layer3_outputs(2911) <= not(layer2_outputs(5073));
    layer3_outputs(2912) <= '1';
    layer3_outputs(2913) <= not(layer2_outputs(557)) or (layer2_outputs(6210));
    layer3_outputs(2914) <= (layer2_outputs(5487)) and (layer2_outputs(4992));
    layer3_outputs(2915) <= (layer2_outputs(3893)) or (layer2_outputs(3415));
    layer3_outputs(2916) <= not(layer2_outputs(933));
    layer3_outputs(2917) <= not(layer2_outputs(7482)) or (layer2_outputs(2899));
    layer3_outputs(2918) <= '1';
    layer3_outputs(2919) <= not(layer2_outputs(4597));
    layer3_outputs(2920) <= layer2_outputs(6984);
    layer3_outputs(2921) <= not(layer2_outputs(1476)) or (layer2_outputs(1868));
    layer3_outputs(2922) <= not(layer2_outputs(1373)) or (layer2_outputs(6247));
    layer3_outputs(2923) <= '1';
    layer3_outputs(2924) <= layer2_outputs(2411);
    layer3_outputs(2925) <= (layer2_outputs(7006)) or (layer2_outputs(3592));
    layer3_outputs(2926) <= '1';
    layer3_outputs(2927) <= layer2_outputs(7534);
    layer3_outputs(2928) <= not(layer2_outputs(7603));
    layer3_outputs(2929) <= (layer2_outputs(6732)) and not (layer2_outputs(526));
    layer3_outputs(2930) <= not((layer2_outputs(4840)) and (layer2_outputs(6296)));
    layer3_outputs(2931) <= not((layer2_outputs(6001)) and (layer2_outputs(3902)));
    layer3_outputs(2932) <= not((layer2_outputs(3478)) and (layer2_outputs(3551)));
    layer3_outputs(2933) <= (layer2_outputs(6754)) and not (layer2_outputs(3390));
    layer3_outputs(2934) <= not(layer2_outputs(4287)) or (layer2_outputs(5789));
    layer3_outputs(2935) <= not(layer2_outputs(2193)) or (layer2_outputs(3054));
    layer3_outputs(2936) <= not(layer2_outputs(866));
    layer3_outputs(2937) <= layer2_outputs(1901);
    layer3_outputs(2938) <= (layer2_outputs(2470)) xor (layer2_outputs(3738));
    layer3_outputs(2939) <= not((layer2_outputs(627)) and (layer2_outputs(6909)));
    layer3_outputs(2940) <= not(layer2_outputs(2851));
    layer3_outputs(2941) <= not(layer2_outputs(2940));
    layer3_outputs(2942) <= layer2_outputs(4949);
    layer3_outputs(2943) <= layer2_outputs(5263);
    layer3_outputs(2944) <= not(layer2_outputs(6189));
    layer3_outputs(2945) <= not((layer2_outputs(2259)) and (layer2_outputs(2962)));
    layer3_outputs(2946) <= layer2_outputs(2208);
    layer3_outputs(2947) <= (layer2_outputs(4037)) xor (layer2_outputs(1739));
    layer3_outputs(2948) <= layer2_outputs(6306);
    layer3_outputs(2949) <= (layer2_outputs(488)) xor (layer2_outputs(631));
    layer3_outputs(2950) <= layer2_outputs(5027);
    layer3_outputs(2951) <= not(layer2_outputs(4650)) or (layer2_outputs(3395));
    layer3_outputs(2952) <= not(layer2_outputs(1041));
    layer3_outputs(2953) <= not(layer2_outputs(2270));
    layer3_outputs(2954) <= not(layer2_outputs(7611));
    layer3_outputs(2955) <= (layer2_outputs(3244)) or (layer2_outputs(2472));
    layer3_outputs(2956) <= not((layer2_outputs(3207)) or (layer2_outputs(675)));
    layer3_outputs(2957) <= not(layer2_outputs(7622)) or (layer2_outputs(4278));
    layer3_outputs(2958) <= not(layer2_outputs(425)) or (layer2_outputs(7381));
    layer3_outputs(2959) <= not(layer2_outputs(1320));
    layer3_outputs(2960) <= layer2_outputs(3354);
    layer3_outputs(2961) <= (layer2_outputs(4730)) and not (layer2_outputs(3976));
    layer3_outputs(2962) <= (layer2_outputs(6417)) and not (layer2_outputs(6955));
    layer3_outputs(2963) <= not(layer2_outputs(6149));
    layer3_outputs(2964) <= layer2_outputs(5754);
    layer3_outputs(2965) <= not(layer2_outputs(5589));
    layer3_outputs(2966) <= (layer2_outputs(791)) or (layer2_outputs(2406));
    layer3_outputs(2967) <= '0';
    layer3_outputs(2968) <= not(layer2_outputs(5970));
    layer3_outputs(2969) <= '1';
    layer3_outputs(2970) <= not(layer2_outputs(3701));
    layer3_outputs(2971) <= (layer2_outputs(715)) and not (layer2_outputs(6118));
    layer3_outputs(2972) <= not(layer2_outputs(3044));
    layer3_outputs(2973) <= layer2_outputs(2106);
    layer3_outputs(2974) <= layer2_outputs(6686);
    layer3_outputs(2975) <= not((layer2_outputs(3489)) and (layer2_outputs(7539)));
    layer3_outputs(2976) <= not((layer2_outputs(1028)) and (layer2_outputs(6989)));
    layer3_outputs(2977) <= not(layer2_outputs(1869));
    layer3_outputs(2978) <= layer2_outputs(5738);
    layer3_outputs(2979) <= (layer2_outputs(5963)) xor (layer2_outputs(751));
    layer3_outputs(2980) <= not((layer2_outputs(1184)) xor (layer2_outputs(314)));
    layer3_outputs(2981) <= layer2_outputs(5689);
    layer3_outputs(2982) <= not(layer2_outputs(432)) or (layer2_outputs(5119));
    layer3_outputs(2983) <= not(layer2_outputs(4357));
    layer3_outputs(2984) <= '0';
    layer3_outputs(2985) <= layer2_outputs(7327);
    layer3_outputs(2986) <= (layer2_outputs(1693)) and not (layer2_outputs(4706));
    layer3_outputs(2987) <= not(layer2_outputs(6746));
    layer3_outputs(2988) <= not(layer2_outputs(353));
    layer3_outputs(2989) <= not(layer2_outputs(2838)) or (layer2_outputs(1113));
    layer3_outputs(2990) <= not((layer2_outputs(3118)) or (layer2_outputs(825)));
    layer3_outputs(2991) <= not(layer2_outputs(5284));
    layer3_outputs(2992) <= not(layer2_outputs(5928)) or (layer2_outputs(3765));
    layer3_outputs(2993) <= not(layer2_outputs(1098)) or (layer2_outputs(2019));
    layer3_outputs(2994) <= layer2_outputs(6220);
    layer3_outputs(2995) <= not(layer2_outputs(6954)) or (layer2_outputs(4464));
    layer3_outputs(2996) <= '1';
    layer3_outputs(2997) <= (layer2_outputs(4173)) and (layer2_outputs(6373));
    layer3_outputs(2998) <= layer2_outputs(1349);
    layer3_outputs(2999) <= layer2_outputs(4783);
    layer3_outputs(3000) <= (layer2_outputs(7251)) or (layer2_outputs(5473));
    layer3_outputs(3001) <= layer2_outputs(3770);
    layer3_outputs(3002) <= not(layer2_outputs(7463)) or (layer2_outputs(6068));
    layer3_outputs(3003) <= not(layer2_outputs(2491));
    layer3_outputs(3004) <= not(layer2_outputs(1730));
    layer3_outputs(3005) <= layer2_outputs(2881);
    layer3_outputs(3006) <= not((layer2_outputs(3806)) or (layer2_outputs(7377)));
    layer3_outputs(3007) <= not(layer2_outputs(4859));
    layer3_outputs(3008) <= not(layer2_outputs(2999));
    layer3_outputs(3009) <= not(layer2_outputs(6295));
    layer3_outputs(3010) <= '1';
    layer3_outputs(3011) <= (layer2_outputs(5459)) or (layer2_outputs(6431));
    layer3_outputs(3012) <= not(layer2_outputs(5091));
    layer3_outputs(3013) <= not(layer2_outputs(6557));
    layer3_outputs(3014) <= not(layer2_outputs(798)) or (layer2_outputs(5839));
    layer3_outputs(3015) <= not(layer2_outputs(6128));
    layer3_outputs(3016) <= not((layer2_outputs(4094)) xor (layer2_outputs(4611)));
    layer3_outputs(3017) <= not((layer2_outputs(2477)) xor (layer2_outputs(5097)));
    layer3_outputs(3018) <= not((layer2_outputs(4146)) or (layer2_outputs(2762)));
    layer3_outputs(3019) <= not(layer2_outputs(6139));
    layer3_outputs(3020) <= not(layer2_outputs(2407));
    layer3_outputs(3021) <= not(layer2_outputs(4639)) or (layer2_outputs(3922));
    layer3_outputs(3022) <= not(layer2_outputs(2885));
    layer3_outputs(3023) <= layer2_outputs(3004);
    layer3_outputs(3024) <= not((layer2_outputs(1605)) xor (layer2_outputs(2982)));
    layer3_outputs(3025) <= not(layer2_outputs(6058));
    layer3_outputs(3026) <= (layer2_outputs(913)) and not (layer2_outputs(1749));
    layer3_outputs(3027) <= not((layer2_outputs(4893)) and (layer2_outputs(542)));
    layer3_outputs(3028) <= (layer2_outputs(3517)) and not (layer2_outputs(1334));
    layer3_outputs(3029) <= (layer2_outputs(194)) and not (layer2_outputs(5278));
    layer3_outputs(3030) <= (layer2_outputs(2014)) xor (layer2_outputs(4865));
    layer3_outputs(3031) <= not(layer2_outputs(3651)) or (layer2_outputs(7132));
    layer3_outputs(3032) <= layer2_outputs(7559);
    layer3_outputs(3033) <= not((layer2_outputs(4270)) xor (layer2_outputs(6744)));
    layer3_outputs(3034) <= (layer2_outputs(47)) xor (layer2_outputs(7013));
    layer3_outputs(3035) <= (layer2_outputs(448)) and (layer2_outputs(6651));
    layer3_outputs(3036) <= not(layer2_outputs(1660)) or (layer2_outputs(7116));
    layer3_outputs(3037) <= (layer2_outputs(4353)) and (layer2_outputs(5176));
    layer3_outputs(3038) <= (layer2_outputs(1249)) and not (layer2_outputs(7174));
    layer3_outputs(3039) <= not(layer2_outputs(2722)) or (layer2_outputs(6445));
    layer3_outputs(3040) <= '1';
    layer3_outputs(3041) <= (layer2_outputs(6420)) and (layer2_outputs(2634));
    layer3_outputs(3042) <= (layer2_outputs(5661)) and not (layer2_outputs(3774));
    layer3_outputs(3043) <= layer2_outputs(1792);
    layer3_outputs(3044) <= (layer2_outputs(1246)) or (layer2_outputs(4955));
    layer3_outputs(3045) <= '0';
    layer3_outputs(3046) <= not(layer2_outputs(2127)) or (layer2_outputs(874));
    layer3_outputs(3047) <= not(layer2_outputs(5385)) or (layer2_outputs(432));
    layer3_outputs(3048) <= not((layer2_outputs(4966)) and (layer2_outputs(4285)));
    layer3_outputs(3049) <= not(layer2_outputs(5156));
    layer3_outputs(3050) <= layer2_outputs(1346);
    layer3_outputs(3051) <= (layer2_outputs(5052)) or (layer2_outputs(4328));
    layer3_outputs(3052) <= (layer2_outputs(3328)) or (layer2_outputs(7422));
    layer3_outputs(3053) <= not(layer2_outputs(1135));
    layer3_outputs(3054) <= layer2_outputs(5855);
    layer3_outputs(3055) <= layer2_outputs(6894);
    layer3_outputs(3056) <= (layer2_outputs(690)) and not (layer2_outputs(3029));
    layer3_outputs(3057) <= (layer2_outputs(6870)) xor (layer2_outputs(1186));
    layer3_outputs(3058) <= not((layer2_outputs(3148)) and (layer2_outputs(2531)));
    layer3_outputs(3059) <= not(layer2_outputs(939));
    layer3_outputs(3060) <= (layer2_outputs(2153)) and (layer2_outputs(448));
    layer3_outputs(3061) <= not((layer2_outputs(6554)) and (layer2_outputs(4866)));
    layer3_outputs(3062) <= not((layer2_outputs(1313)) and (layer2_outputs(4310)));
    layer3_outputs(3063) <= layer2_outputs(467);
    layer3_outputs(3064) <= not((layer2_outputs(660)) or (layer2_outputs(5993)));
    layer3_outputs(3065) <= layer2_outputs(5403);
    layer3_outputs(3066) <= (layer2_outputs(795)) and not (layer2_outputs(2606));
    layer3_outputs(3067) <= layer2_outputs(1544);
    layer3_outputs(3068) <= layer2_outputs(1554);
    layer3_outputs(3069) <= (layer2_outputs(6962)) xor (layer2_outputs(6966));
    layer3_outputs(3070) <= not(layer2_outputs(3115));
    layer3_outputs(3071) <= not((layer2_outputs(5713)) and (layer2_outputs(4307)));
    layer3_outputs(3072) <= (layer2_outputs(1569)) and not (layer2_outputs(4906));
    layer3_outputs(3073) <= not(layer2_outputs(5337));
    layer3_outputs(3074) <= layer2_outputs(7121);
    layer3_outputs(3075) <= '0';
    layer3_outputs(3076) <= layer2_outputs(2118);
    layer3_outputs(3077) <= not(layer2_outputs(4527));
    layer3_outputs(3078) <= (layer2_outputs(5245)) and not (layer2_outputs(6258));
    layer3_outputs(3079) <= not(layer2_outputs(1270));
    layer3_outputs(3080) <= (layer2_outputs(6374)) xor (layer2_outputs(3285));
    layer3_outputs(3081) <= layer2_outputs(4740);
    layer3_outputs(3082) <= layer2_outputs(3522);
    layer3_outputs(3083) <= not(layer2_outputs(5377));
    layer3_outputs(3084) <= not(layer2_outputs(3603));
    layer3_outputs(3085) <= not(layer2_outputs(4092));
    layer3_outputs(3086) <= not(layer2_outputs(6348)) or (layer2_outputs(706));
    layer3_outputs(3087) <= layer2_outputs(202);
    layer3_outputs(3088) <= layer2_outputs(5729);
    layer3_outputs(3089) <= not(layer2_outputs(1236)) or (layer2_outputs(7436));
    layer3_outputs(3090) <= not(layer2_outputs(1468));
    layer3_outputs(3091) <= not(layer2_outputs(565));
    layer3_outputs(3092) <= (layer2_outputs(1356)) and not (layer2_outputs(877));
    layer3_outputs(3093) <= '1';
    layer3_outputs(3094) <= not((layer2_outputs(4820)) and (layer2_outputs(222)));
    layer3_outputs(3095) <= not((layer2_outputs(2415)) or (layer2_outputs(1498)));
    layer3_outputs(3096) <= not(layer2_outputs(5017));
    layer3_outputs(3097) <= (layer2_outputs(7224)) and (layer2_outputs(4851));
    layer3_outputs(3098) <= (layer2_outputs(3288)) or (layer2_outputs(1309));
    layer3_outputs(3099) <= (layer2_outputs(4662)) or (layer2_outputs(3550));
    layer3_outputs(3100) <= (layer2_outputs(1417)) or (layer2_outputs(5184));
    layer3_outputs(3101) <= layer2_outputs(5077);
    layer3_outputs(3102) <= not((layer2_outputs(4972)) and (layer2_outputs(2109)));
    layer3_outputs(3103) <= (layer2_outputs(2936)) xor (layer2_outputs(3608));
    layer3_outputs(3104) <= not(layer2_outputs(6748));
    layer3_outputs(3105) <= layer2_outputs(6016);
    layer3_outputs(3106) <= (layer2_outputs(1176)) or (layer2_outputs(6311));
    layer3_outputs(3107) <= (layer2_outputs(3918)) and not (layer2_outputs(7634));
    layer3_outputs(3108) <= layer2_outputs(2920);
    layer3_outputs(3109) <= not((layer2_outputs(4182)) and (layer2_outputs(3280)));
    layer3_outputs(3110) <= not(layer2_outputs(3676));
    layer3_outputs(3111) <= layer2_outputs(7008);
    layer3_outputs(3112) <= (layer2_outputs(2725)) xor (layer2_outputs(7286));
    layer3_outputs(3113) <= (layer2_outputs(7060)) or (layer2_outputs(6494));
    layer3_outputs(3114) <= '0';
    layer3_outputs(3115) <= '1';
    layer3_outputs(3116) <= not(layer2_outputs(4142));
    layer3_outputs(3117) <= not(layer2_outputs(5086));
    layer3_outputs(3118) <= not((layer2_outputs(5986)) or (layer2_outputs(4549)));
    layer3_outputs(3119) <= '1';
    layer3_outputs(3120) <= not(layer2_outputs(5559));
    layer3_outputs(3121) <= (layer2_outputs(5358)) xor (layer2_outputs(5844));
    layer3_outputs(3122) <= not(layer2_outputs(2046));
    layer3_outputs(3123) <= layer2_outputs(3718);
    layer3_outputs(3124) <= not(layer2_outputs(4009)) or (layer2_outputs(2284));
    layer3_outputs(3125) <= not(layer2_outputs(1332));
    layer3_outputs(3126) <= (layer2_outputs(2304)) and not (layer2_outputs(3610));
    layer3_outputs(3127) <= (layer2_outputs(2175)) or (layer2_outputs(4644));
    layer3_outputs(3128) <= layer2_outputs(6550);
    layer3_outputs(3129) <= not((layer2_outputs(77)) and (layer2_outputs(6805)));
    layer3_outputs(3130) <= (layer2_outputs(931)) and not (layer2_outputs(6233));
    layer3_outputs(3131) <= not(layer2_outputs(4183));
    layer3_outputs(3132) <= not((layer2_outputs(5064)) or (layer2_outputs(7664)));
    layer3_outputs(3133) <= not(layer2_outputs(829)) or (layer2_outputs(5497));
    layer3_outputs(3134) <= (layer2_outputs(3777)) and not (layer2_outputs(1831));
    layer3_outputs(3135) <= not(layer2_outputs(6239));
    layer3_outputs(3136) <= (layer2_outputs(6830)) xor (layer2_outputs(2319));
    layer3_outputs(3137) <= not(layer2_outputs(6161));
    layer3_outputs(3138) <= layer2_outputs(551);
    layer3_outputs(3139) <= (layer2_outputs(887)) or (layer2_outputs(3276));
    layer3_outputs(3140) <= layer2_outputs(2722);
    layer3_outputs(3141) <= (layer2_outputs(5970)) or (layer2_outputs(1675));
    layer3_outputs(3142) <= not((layer2_outputs(3429)) and (layer2_outputs(2533)));
    layer3_outputs(3143) <= not(layer2_outputs(5146)) or (layer2_outputs(2759));
    layer3_outputs(3144) <= not((layer2_outputs(1289)) and (layer2_outputs(4284)));
    layer3_outputs(3145) <= not((layer2_outputs(7304)) or (layer2_outputs(6908)));
    layer3_outputs(3146) <= not(layer2_outputs(969));
    layer3_outputs(3147) <= layer2_outputs(3411);
    layer3_outputs(3148) <= (layer2_outputs(3348)) xor (layer2_outputs(6501));
    layer3_outputs(3149) <= not(layer2_outputs(5006)) or (layer2_outputs(2549));
    layer3_outputs(3150) <= layer2_outputs(2930);
    layer3_outputs(3151) <= layer2_outputs(7082);
    layer3_outputs(3152) <= layer2_outputs(6561);
    layer3_outputs(3153) <= layer2_outputs(3625);
    layer3_outputs(3154) <= '1';
    layer3_outputs(3155) <= (layer2_outputs(1454)) xor (layer2_outputs(137));
    layer3_outputs(3156) <= (layer2_outputs(7050)) and not (layer2_outputs(1295));
    layer3_outputs(3157) <= not((layer2_outputs(5920)) or (layer2_outputs(7245)));
    layer3_outputs(3158) <= layer2_outputs(405);
    layer3_outputs(3159) <= not((layer2_outputs(7209)) and (layer2_outputs(668)));
    layer3_outputs(3160) <= (layer2_outputs(2177)) and not (layer2_outputs(7514));
    layer3_outputs(3161) <= not(layer2_outputs(6938));
    layer3_outputs(3162) <= not((layer2_outputs(2963)) and (layer2_outputs(6774)));
    layer3_outputs(3163) <= not(layer2_outputs(6088));
    layer3_outputs(3164) <= (layer2_outputs(1287)) or (layer2_outputs(573));
    layer3_outputs(3165) <= (layer2_outputs(2906)) and not (layer2_outputs(5644));
    layer3_outputs(3166) <= (layer2_outputs(7063)) and not (layer2_outputs(2994));
    layer3_outputs(3167) <= not(layer2_outputs(3571)) or (layer2_outputs(3296));
    layer3_outputs(3168) <= layer2_outputs(6719);
    layer3_outputs(3169) <= layer2_outputs(7259);
    layer3_outputs(3170) <= not(layer2_outputs(263));
    layer3_outputs(3171) <= layer2_outputs(7012);
    layer3_outputs(3172) <= not(layer2_outputs(211));
    layer3_outputs(3173) <= layer2_outputs(1738);
    layer3_outputs(3174) <= not(layer2_outputs(871)) or (layer2_outputs(848));
    layer3_outputs(3175) <= not(layer2_outputs(902));
    layer3_outputs(3176) <= (layer2_outputs(4409)) and not (layer2_outputs(2279));
    layer3_outputs(3177) <= layer2_outputs(6811);
    layer3_outputs(3178) <= (layer2_outputs(5038)) or (layer2_outputs(1649));
    layer3_outputs(3179) <= layer2_outputs(5047);
    layer3_outputs(3180) <= (layer2_outputs(5882)) and not (layer2_outputs(2444));
    layer3_outputs(3181) <= not(layer2_outputs(4744)) or (layer2_outputs(3801));
    layer3_outputs(3182) <= (layer2_outputs(2310)) xor (layer2_outputs(94));
    layer3_outputs(3183) <= not(layer2_outputs(1476));
    layer3_outputs(3184) <= (layer2_outputs(1971)) and not (layer2_outputs(7368));
    layer3_outputs(3185) <= layer2_outputs(4659);
    layer3_outputs(3186) <= not(layer2_outputs(1344));
    layer3_outputs(3187) <= layer2_outputs(700);
    layer3_outputs(3188) <= not(layer2_outputs(326));
    layer3_outputs(3189) <= (layer2_outputs(1583)) or (layer2_outputs(4140));
    layer3_outputs(3190) <= layer2_outputs(4808);
    layer3_outputs(3191) <= (layer2_outputs(6497)) or (layer2_outputs(2571));
    layer3_outputs(3192) <= (layer2_outputs(4062)) and (layer2_outputs(2867));
    layer3_outputs(3193) <= (layer2_outputs(5800)) or (layer2_outputs(3563));
    layer3_outputs(3194) <= layer2_outputs(2288);
    layer3_outputs(3195) <= not(layer2_outputs(2595)) or (layer2_outputs(1146));
    layer3_outputs(3196) <= not(layer2_outputs(6598));
    layer3_outputs(3197) <= not((layer2_outputs(848)) and (layer2_outputs(1929)));
    layer3_outputs(3198) <= (layer2_outputs(4313)) and not (layer2_outputs(2293));
    layer3_outputs(3199) <= not((layer2_outputs(34)) xor (layer2_outputs(7364)));
    layer3_outputs(3200) <= not(layer2_outputs(2365));
    layer3_outputs(3201) <= (layer2_outputs(3013)) and not (layer2_outputs(3843));
    layer3_outputs(3202) <= (layer2_outputs(5204)) and (layer2_outputs(4687));
    layer3_outputs(3203) <= (layer2_outputs(4442)) and (layer2_outputs(1924));
    layer3_outputs(3204) <= not(layer2_outputs(4201));
    layer3_outputs(3205) <= layer2_outputs(1233);
    layer3_outputs(3206) <= layer2_outputs(912);
    layer3_outputs(3207) <= (layer2_outputs(4175)) and (layer2_outputs(6741));
    layer3_outputs(3208) <= layer2_outputs(771);
    layer3_outputs(3209) <= '0';
    layer3_outputs(3210) <= not((layer2_outputs(2675)) and (layer2_outputs(7136)));
    layer3_outputs(3211) <= not((layer2_outputs(2613)) xor (layer2_outputs(2003)));
    layer3_outputs(3212) <= (layer2_outputs(7448)) and (layer2_outputs(2020));
    layer3_outputs(3213) <= not(layer2_outputs(5471));
    layer3_outputs(3214) <= layer2_outputs(862);
    layer3_outputs(3215) <= '0';
    layer3_outputs(3216) <= (layer2_outputs(4121)) xor (layer2_outputs(673));
    layer3_outputs(3217) <= (layer2_outputs(3894)) xor (layer2_outputs(4799));
    layer3_outputs(3218) <= not((layer2_outputs(5828)) or (layer2_outputs(5783)));
    layer3_outputs(3219) <= (layer2_outputs(5714)) xor (layer2_outputs(2343));
    layer3_outputs(3220) <= not(layer2_outputs(7575));
    layer3_outputs(3221) <= (layer2_outputs(430)) xor (layer2_outputs(4387));
    layer3_outputs(3222) <= layer2_outputs(4445);
    layer3_outputs(3223) <= (layer2_outputs(1921)) and (layer2_outputs(7321));
    layer3_outputs(3224) <= not(layer2_outputs(128));
    layer3_outputs(3225) <= not(layer2_outputs(5530)) or (layer2_outputs(2279));
    layer3_outputs(3226) <= layer2_outputs(3432);
    layer3_outputs(3227) <= not(layer2_outputs(5386)) or (layer2_outputs(7048));
    layer3_outputs(3228) <= (layer2_outputs(3872)) and (layer2_outputs(6589));
    layer3_outputs(3229) <= (layer2_outputs(4269)) and (layer2_outputs(5010));
    layer3_outputs(3230) <= (layer2_outputs(6829)) or (layer2_outputs(273));
    layer3_outputs(3231) <= not(layer2_outputs(5180));
    layer3_outputs(3232) <= '1';
    layer3_outputs(3233) <= layer2_outputs(6349);
    layer3_outputs(3234) <= (layer2_outputs(1148)) and (layer2_outputs(4317));
    layer3_outputs(3235) <= not(layer2_outputs(518)) or (layer2_outputs(1011));
    layer3_outputs(3236) <= '1';
    layer3_outputs(3237) <= layer2_outputs(4249);
    layer3_outputs(3238) <= not(layer2_outputs(4613));
    layer3_outputs(3239) <= not((layer2_outputs(1920)) or (layer2_outputs(7405)));
    layer3_outputs(3240) <= layer2_outputs(5022);
    layer3_outputs(3241) <= (layer2_outputs(5109)) and (layer2_outputs(1351));
    layer3_outputs(3242) <= not((layer2_outputs(2929)) xor (layer2_outputs(4961)));
    layer3_outputs(3243) <= not((layer2_outputs(6963)) and (layer2_outputs(6884)));
    layer3_outputs(3244) <= not((layer2_outputs(3782)) or (layer2_outputs(1891)));
    layer3_outputs(3245) <= (layer2_outputs(315)) xor (layer2_outputs(7546));
    layer3_outputs(3246) <= layer2_outputs(6810);
    layer3_outputs(3247) <= not(layer2_outputs(3468));
    layer3_outputs(3248) <= layer2_outputs(4416);
    layer3_outputs(3249) <= not(layer2_outputs(3480)) or (layer2_outputs(2481));
    layer3_outputs(3250) <= not((layer2_outputs(7387)) or (layer2_outputs(7674)));
    layer3_outputs(3251) <= not(layer2_outputs(4067)) or (layer2_outputs(1836));
    layer3_outputs(3252) <= not(layer2_outputs(2202)) or (layer2_outputs(7146));
    layer3_outputs(3253) <= layer2_outputs(3797);
    layer3_outputs(3254) <= (layer2_outputs(5092)) or (layer2_outputs(4286));
    layer3_outputs(3255) <= layer2_outputs(6534);
    layer3_outputs(3256) <= layer2_outputs(1600);
    layer3_outputs(3257) <= (layer2_outputs(1171)) or (layer2_outputs(6347));
    layer3_outputs(3258) <= (layer2_outputs(562)) and (layer2_outputs(170));
    layer3_outputs(3259) <= not(layer2_outputs(7175));
    layer3_outputs(3260) <= not(layer2_outputs(2022));
    layer3_outputs(3261) <= not(layer2_outputs(4468));
    layer3_outputs(3262) <= layer2_outputs(11);
    layer3_outputs(3263) <= not(layer2_outputs(1321));
    layer3_outputs(3264) <= layer2_outputs(6246);
    layer3_outputs(3265) <= not(layer2_outputs(4822));
    layer3_outputs(3266) <= not(layer2_outputs(5297));
    layer3_outputs(3267) <= not(layer2_outputs(3012)) or (layer2_outputs(3284));
    layer3_outputs(3268) <= not(layer2_outputs(4781));
    layer3_outputs(3269) <= layer2_outputs(721);
    layer3_outputs(3270) <= layer2_outputs(4822);
    layer3_outputs(3271) <= not(layer2_outputs(863));
    layer3_outputs(3272) <= layer2_outputs(4047);
    layer3_outputs(3273) <= not(layer2_outputs(2418));
    layer3_outputs(3274) <= (layer2_outputs(7460)) and not (layer2_outputs(7429));
    layer3_outputs(3275) <= not(layer2_outputs(2511));
    layer3_outputs(3276) <= layer2_outputs(3074);
    layer3_outputs(3277) <= not(layer2_outputs(4328));
    layer3_outputs(3278) <= (layer2_outputs(4423)) and (layer2_outputs(6408));
    layer3_outputs(3279) <= not(layer2_outputs(5795)) or (layer2_outputs(3554));
    layer3_outputs(3280) <= '1';
    layer3_outputs(3281) <= not(layer2_outputs(5687));
    layer3_outputs(3282) <= (layer2_outputs(6040)) and (layer2_outputs(4343));
    layer3_outputs(3283) <= (layer2_outputs(5802)) and (layer2_outputs(5166));
    layer3_outputs(3284) <= not(layer2_outputs(6150)) or (layer2_outputs(6989));
    layer3_outputs(3285) <= (layer2_outputs(6932)) and not (layer2_outputs(3910));
    layer3_outputs(3286) <= not(layer2_outputs(7226));
    layer3_outputs(3287) <= layer2_outputs(5985);
    layer3_outputs(3288) <= not(layer2_outputs(228));
    layer3_outputs(3289) <= not(layer2_outputs(2925)) or (layer2_outputs(2186));
    layer3_outputs(3290) <= layer2_outputs(5452);
    layer3_outputs(3291) <= not(layer2_outputs(7636)) or (layer2_outputs(3451));
    layer3_outputs(3292) <= not((layer2_outputs(574)) or (layer2_outputs(610)));
    layer3_outputs(3293) <= (layer2_outputs(4981)) and (layer2_outputs(413));
    layer3_outputs(3294) <= layer2_outputs(1790);
    layer3_outputs(3295) <= not((layer2_outputs(7442)) xor (layer2_outputs(4875)));
    layer3_outputs(3296) <= (layer2_outputs(5460)) and not (layer2_outputs(6076));
    layer3_outputs(3297) <= layer2_outputs(2068);
    layer3_outputs(3298) <= not(layer2_outputs(3731));
    layer3_outputs(3299) <= (layer2_outputs(1425)) or (layer2_outputs(4971));
    layer3_outputs(3300) <= not(layer2_outputs(606)) or (layer2_outputs(798));
    layer3_outputs(3301) <= not(layer2_outputs(4642)) or (layer2_outputs(95));
    layer3_outputs(3302) <= not(layer2_outputs(4633)) or (layer2_outputs(3198));
    layer3_outputs(3303) <= layer2_outputs(3402);
    layer3_outputs(3304) <= (layer2_outputs(4487)) and not (layer2_outputs(2519));
    layer3_outputs(3305) <= not(layer2_outputs(2490));
    layer3_outputs(3306) <= layer2_outputs(5164);
    layer3_outputs(3307) <= layer2_outputs(6471);
    layer3_outputs(3308) <= not((layer2_outputs(3135)) or (layer2_outputs(642)));
    layer3_outputs(3309) <= (layer2_outputs(1392)) and not (layer2_outputs(3456));
    layer3_outputs(3310) <= not(layer2_outputs(4081));
    layer3_outputs(3311) <= (layer2_outputs(4914)) and not (layer2_outputs(3665));
    layer3_outputs(3312) <= layer2_outputs(5969);
    layer3_outputs(3313) <= not((layer2_outputs(841)) xor (layer2_outputs(6423)));
    layer3_outputs(3314) <= layer2_outputs(3407);
    layer3_outputs(3315) <= layer2_outputs(5111);
    layer3_outputs(3316) <= (layer2_outputs(1304)) and not (layer2_outputs(2315));
    layer3_outputs(3317) <= not(layer2_outputs(1441));
    layer3_outputs(3318) <= not(layer2_outputs(7597));
    layer3_outputs(3319) <= not((layer2_outputs(393)) and (layer2_outputs(2221)));
    layer3_outputs(3320) <= layer2_outputs(1615);
    layer3_outputs(3321) <= not(layer2_outputs(6479));
    layer3_outputs(3322) <= not(layer2_outputs(7555));
    layer3_outputs(3323) <= not(layer2_outputs(5885));
    layer3_outputs(3324) <= '0';
    layer3_outputs(3325) <= not(layer2_outputs(4210)) or (layer2_outputs(136));
    layer3_outputs(3326) <= (layer2_outputs(7035)) and not (layer2_outputs(2716));
    layer3_outputs(3327) <= not(layer2_outputs(721));
    layer3_outputs(3328) <= layer2_outputs(4113);
    layer3_outputs(3329) <= (layer2_outputs(5029)) and not (layer2_outputs(2007));
    layer3_outputs(3330) <= not(layer2_outputs(5465));
    layer3_outputs(3331) <= (layer2_outputs(2313)) and (layer2_outputs(3226));
    layer3_outputs(3332) <= not(layer2_outputs(6301)) or (layer2_outputs(3433));
    layer3_outputs(3333) <= not((layer2_outputs(7305)) or (layer2_outputs(85)));
    layer3_outputs(3334) <= layer2_outputs(5703);
    layer3_outputs(3335) <= (layer2_outputs(6415)) or (layer2_outputs(5258));
    layer3_outputs(3336) <= layer2_outputs(5213);
    layer3_outputs(3337) <= not(layer2_outputs(417));
    layer3_outputs(3338) <= layer2_outputs(6165);
    layer3_outputs(3339) <= layer2_outputs(5513);
    layer3_outputs(3340) <= (layer2_outputs(4607)) and not (layer2_outputs(2251));
    layer3_outputs(3341) <= not((layer2_outputs(6278)) or (layer2_outputs(139)));
    layer3_outputs(3342) <= not(layer2_outputs(2926));
    layer3_outputs(3343) <= not(layer2_outputs(2249));
    layer3_outputs(3344) <= (layer2_outputs(4947)) and not (layer2_outputs(3728));
    layer3_outputs(3345) <= layer2_outputs(6178);
    layer3_outputs(3346) <= (layer2_outputs(2253)) and not (layer2_outputs(24));
    layer3_outputs(3347) <= not(layer2_outputs(3901));
    layer3_outputs(3348) <= not(layer2_outputs(2077)) or (layer2_outputs(179));
    layer3_outputs(3349) <= (layer2_outputs(4862)) and (layer2_outputs(3692));
    layer3_outputs(3350) <= (layer2_outputs(286)) xor (layer2_outputs(168));
    layer3_outputs(3351) <= not(layer2_outputs(113)) or (layer2_outputs(7171));
    layer3_outputs(3352) <= layer2_outputs(5930);
    layer3_outputs(3353) <= not(layer2_outputs(1099)) or (layer2_outputs(729));
    layer3_outputs(3354) <= not((layer2_outputs(7602)) or (layer2_outputs(1593)));
    layer3_outputs(3355) <= not(layer2_outputs(7552)) or (layer2_outputs(2198));
    layer3_outputs(3356) <= not(layer2_outputs(5085));
    layer3_outputs(3357) <= not((layer2_outputs(2733)) and (layer2_outputs(4939)));
    layer3_outputs(3358) <= not(layer2_outputs(5431));
    layer3_outputs(3359) <= (layer2_outputs(1846)) or (layer2_outputs(1345));
    layer3_outputs(3360) <= layer2_outputs(3150);
    layer3_outputs(3361) <= not(layer2_outputs(2792));
    layer3_outputs(3362) <= layer2_outputs(1123);
    layer3_outputs(3363) <= layer2_outputs(3502);
    layer3_outputs(3364) <= not((layer2_outputs(1964)) or (layer2_outputs(1932)));
    layer3_outputs(3365) <= layer2_outputs(183);
    layer3_outputs(3366) <= layer2_outputs(4982);
    layer3_outputs(3367) <= layer2_outputs(3500);
    layer3_outputs(3368) <= not(layer2_outputs(5464)) or (layer2_outputs(685));
    layer3_outputs(3369) <= (layer2_outputs(4872)) and not (layer2_outputs(2597));
    layer3_outputs(3370) <= layer2_outputs(4663);
    layer3_outputs(3371) <= not((layer2_outputs(5206)) xor (layer2_outputs(6717)));
    layer3_outputs(3372) <= (layer2_outputs(7484)) xor (layer2_outputs(3969));
    layer3_outputs(3373) <= layer2_outputs(2231);
    layer3_outputs(3374) <= not(layer2_outputs(3011));
    layer3_outputs(3375) <= (layer2_outputs(6975)) and not (layer2_outputs(3038));
    layer3_outputs(3376) <= layer2_outputs(6370);
    layer3_outputs(3377) <= not((layer2_outputs(4075)) and (layer2_outputs(7101)));
    layer3_outputs(3378) <= layer2_outputs(3915);
    layer3_outputs(3379) <= not(layer2_outputs(5055));
    layer3_outputs(3380) <= not(layer2_outputs(6526)) or (layer2_outputs(4373));
    layer3_outputs(3381) <= not((layer2_outputs(2104)) and (layer2_outputs(590)));
    layer3_outputs(3382) <= not(layer2_outputs(2627));
    layer3_outputs(3383) <= not(layer2_outputs(2828)) or (layer2_outputs(7275));
    layer3_outputs(3384) <= (layer2_outputs(4690)) and not (layer2_outputs(6624));
    layer3_outputs(3385) <= (layer2_outputs(6881)) and not (layer2_outputs(5946));
    layer3_outputs(3386) <= layer2_outputs(6638);
    layer3_outputs(3387) <= layer2_outputs(7575);
    layer3_outputs(3388) <= not(layer2_outputs(1626));
    layer3_outputs(3389) <= not((layer2_outputs(1186)) or (layer2_outputs(6788)));
    layer3_outputs(3390) <= layer2_outputs(121);
    layer3_outputs(3391) <= layer2_outputs(1744);
    layer3_outputs(3392) <= layer2_outputs(3028);
    layer3_outputs(3393) <= layer2_outputs(3176);
    layer3_outputs(3394) <= not(layer2_outputs(3766));
    layer3_outputs(3395) <= layer2_outputs(4418);
    layer3_outputs(3396) <= not((layer2_outputs(2021)) or (layer2_outputs(1755)));
    layer3_outputs(3397) <= '1';
    layer3_outputs(3398) <= (layer2_outputs(6647)) and not (layer2_outputs(5832));
    layer3_outputs(3399) <= (layer2_outputs(3341)) or (layer2_outputs(3181));
    layer3_outputs(3400) <= not((layer2_outputs(6450)) and (layer2_outputs(3249)));
    layer3_outputs(3401) <= (layer2_outputs(1818)) and (layer2_outputs(4256));
    layer3_outputs(3402) <= not(layer2_outputs(5254)) or (layer2_outputs(7319));
    layer3_outputs(3403) <= layer2_outputs(1249);
    layer3_outputs(3404) <= '1';
    layer3_outputs(3405) <= not(layer2_outputs(3736)) or (layer2_outputs(2640));
    layer3_outputs(3406) <= (layer2_outputs(5796)) and (layer2_outputs(5812));
    layer3_outputs(3407) <= layer2_outputs(6571);
    layer3_outputs(3408) <= not(layer2_outputs(6257));
    layer3_outputs(3409) <= not(layer2_outputs(5063));
    layer3_outputs(3410) <= (layer2_outputs(548)) and (layer2_outputs(5704));
    layer3_outputs(3411) <= not(layer2_outputs(3202));
    layer3_outputs(3412) <= not(layer2_outputs(4345));
    layer3_outputs(3413) <= not(layer2_outputs(7471)) or (layer2_outputs(3775));
    layer3_outputs(3414) <= layer2_outputs(6673);
    layer3_outputs(3415) <= layer2_outputs(7485);
    layer3_outputs(3416) <= (layer2_outputs(5213)) or (layer2_outputs(3026));
    layer3_outputs(3417) <= (layer2_outputs(2999)) and not (layer2_outputs(341));
    layer3_outputs(3418) <= (layer2_outputs(6926)) xor (layer2_outputs(2123));
    layer3_outputs(3419) <= not(layer2_outputs(2377)) or (layer2_outputs(752));
    layer3_outputs(3420) <= not(layer2_outputs(2331));
    layer3_outputs(3421) <= not(layer2_outputs(5957)) or (layer2_outputs(6250));
    layer3_outputs(3422) <= layer2_outputs(338);
    layer3_outputs(3423) <= layer2_outputs(5201);
    layer3_outputs(3424) <= layer2_outputs(2863);
    layer3_outputs(3425) <= not(layer2_outputs(1992));
    layer3_outputs(3426) <= '0';
    layer3_outputs(3427) <= not(layer2_outputs(993));
    layer3_outputs(3428) <= layer2_outputs(5048);
    layer3_outputs(3429) <= layer2_outputs(3171);
    layer3_outputs(3430) <= (layer2_outputs(5110)) and not (layer2_outputs(4812));
    layer3_outputs(3431) <= not(layer2_outputs(4813)) or (layer2_outputs(4521));
    layer3_outputs(3432) <= (layer2_outputs(4424)) and not (layer2_outputs(962));
    layer3_outputs(3433) <= layer2_outputs(1018);
    layer3_outputs(3434) <= not(layer2_outputs(7466)) or (layer2_outputs(3762));
    layer3_outputs(3435) <= not((layer2_outputs(2887)) or (layer2_outputs(225)));
    layer3_outputs(3436) <= (layer2_outputs(2094)) and not (layer2_outputs(2830));
    layer3_outputs(3437) <= (layer2_outputs(4595)) xor (layer2_outputs(767));
    layer3_outputs(3438) <= layer2_outputs(7140);
    layer3_outputs(3439) <= '0';
    layer3_outputs(3440) <= not(layer2_outputs(6812)) or (layer2_outputs(650));
    layer3_outputs(3441) <= (layer2_outputs(6966)) and (layer2_outputs(1125));
    layer3_outputs(3442) <= not(layer2_outputs(1994));
    layer3_outputs(3443) <= (layer2_outputs(2831)) and not (layer2_outputs(1393));
    layer3_outputs(3444) <= not(layer2_outputs(7032));
    layer3_outputs(3445) <= (layer2_outputs(6496)) and not (layer2_outputs(1255));
    layer3_outputs(3446) <= layer2_outputs(941);
    layer3_outputs(3447) <= (layer2_outputs(1961)) and not (layer2_outputs(1654));
    layer3_outputs(3448) <= not((layer2_outputs(6793)) and (layer2_outputs(6283)));
    layer3_outputs(3449) <= layer2_outputs(1427);
    layer3_outputs(3450) <= (layer2_outputs(3227)) or (layer2_outputs(1665));
    layer3_outputs(3451) <= not(layer2_outputs(6482));
    layer3_outputs(3452) <= (layer2_outputs(6606)) and not (layer2_outputs(5316));
    layer3_outputs(3453) <= (layer2_outputs(2162)) and (layer2_outputs(422));
    layer3_outputs(3454) <= (layer2_outputs(3338)) and not (layer2_outputs(51));
    layer3_outputs(3455) <= (layer2_outputs(257)) xor (layer2_outputs(3839));
    layer3_outputs(3456) <= layer2_outputs(5895);
    layer3_outputs(3457) <= (layer2_outputs(5410)) xor (layer2_outputs(3136));
    layer3_outputs(3458) <= not(layer2_outputs(5943));
    layer3_outputs(3459) <= not(layer2_outputs(5564));
    layer3_outputs(3460) <= layer2_outputs(6704);
    layer3_outputs(3461) <= (layer2_outputs(7133)) or (layer2_outputs(1330));
    layer3_outputs(3462) <= layer2_outputs(849);
    layer3_outputs(3463) <= (layer2_outputs(2285)) and not (layer2_outputs(5147));
    layer3_outputs(3464) <= not(layer2_outputs(5560)) or (layer2_outputs(507));
    layer3_outputs(3465) <= (layer2_outputs(4191)) and not (layer2_outputs(5162));
    layer3_outputs(3466) <= layer2_outputs(906);
    layer3_outputs(3467) <= not(layer2_outputs(5118));
    layer3_outputs(3468) <= not(layer2_outputs(5263)) or (layer2_outputs(6514));
    layer3_outputs(3469) <= not(layer2_outputs(797));
    layer3_outputs(3470) <= (layer2_outputs(438)) and not (layer2_outputs(6763));
    layer3_outputs(3471) <= not(layer2_outputs(5329));
    layer3_outputs(3472) <= (layer2_outputs(1933)) and not (layer2_outputs(6075));
    layer3_outputs(3473) <= not(layer2_outputs(216));
    layer3_outputs(3474) <= (layer2_outputs(7298)) and (layer2_outputs(3345));
    layer3_outputs(3475) <= not(layer2_outputs(4022)) or (layer2_outputs(2725));
    layer3_outputs(3476) <= (layer2_outputs(3657)) and (layer2_outputs(1291));
    layer3_outputs(3477) <= layer2_outputs(1198);
    layer3_outputs(3478) <= not(layer2_outputs(6363));
    layer3_outputs(3479) <= layer2_outputs(6902);
    layer3_outputs(3480) <= (layer2_outputs(2308)) and not (layer2_outputs(398));
    layer3_outputs(3481) <= not((layer2_outputs(1267)) and (layer2_outputs(6493)));
    layer3_outputs(3482) <= '0';
    layer3_outputs(3483) <= layer2_outputs(3186);
    layer3_outputs(3484) <= layer2_outputs(6354);
    layer3_outputs(3485) <= not(layer2_outputs(1388));
    layer3_outputs(3486) <= (layer2_outputs(1158)) or (layer2_outputs(5941));
    layer3_outputs(3487) <= not(layer2_outputs(6372));
    layer3_outputs(3488) <= '1';
    layer3_outputs(3489) <= (layer2_outputs(2839)) and not (layer2_outputs(6997));
    layer3_outputs(3490) <= (layer2_outputs(558)) and not (layer2_outputs(7265));
    layer3_outputs(3491) <= layer2_outputs(3103);
    layer3_outputs(3492) <= not(layer2_outputs(7337));
    layer3_outputs(3493) <= not(layer2_outputs(271)) or (layer2_outputs(2110));
    layer3_outputs(3494) <= not((layer2_outputs(4907)) and (layer2_outputs(259)));
    layer3_outputs(3495) <= not((layer2_outputs(4916)) or (layer2_outputs(6247)));
    layer3_outputs(3496) <= not((layer2_outputs(5317)) xor (layer2_outputs(100)));
    layer3_outputs(3497) <= (layer2_outputs(2380)) and not (layer2_outputs(2071));
    layer3_outputs(3498) <= layer2_outputs(4116);
    layer3_outputs(3499) <= not(layer2_outputs(1221));
    layer3_outputs(3500) <= (layer2_outputs(4839)) and (layer2_outputs(3040));
    layer3_outputs(3501) <= layer2_outputs(3063);
    layer3_outputs(3502) <= not(layer2_outputs(7139));
    layer3_outputs(3503) <= (layer2_outputs(7254)) and not (layer2_outputs(1553));
    layer3_outputs(3504) <= not(layer2_outputs(4506));
    layer3_outputs(3505) <= layer2_outputs(5810);
    layer3_outputs(3506) <= not(layer2_outputs(6296));
    layer3_outputs(3507) <= (layer2_outputs(93)) or (layer2_outputs(742));
    layer3_outputs(3508) <= (layer2_outputs(5461)) and not (layer2_outputs(4911));
    layer3_outputs(3509) <= '1';
    layer3_outputs(3510) <= not(layer2_outputs(963));
    layer3_outputs(3511) <= not((layer2_outputs(6392)) and (layer2_outputs(3628)));
    layer3_outputs(3512) <= not((layer2_outputs(7643)) xor (layer2_outputs(3518)));
    layer3_outputs(3513) <= layer2_outputs(3060);
    layer3_outputs(3514) <= (layer2_outputs(5405)) and not (layer2_outputs(5758));
    layer3_outputs(3515) <= not(layer2_outputs(5235)) or (layer2_outputs(136));
    layer3_outputs(3516) <= not(layer2_outputs(600));
    layer3_outputs(3517) <= (layer2_outputs(7185)) and (layer2_outputs(1308));
    layer3_outputs(3518) <= layer2_outputs(6850);
    layer3_outputs(3519) <= (layer2_outputs(4735)) and (layer2_outputs(1705));
    layer3_outputs(3520) <= layer2_outputs(5728);
    layer3_outputs(3521) <= (layer2_outputs(4975)) and not (layer2_outputs(1087));
    layer3_outputs(3522) <= not((layer2_outputs(3262)) or (layer2_outputs(2683)));
    layer3_outputs(3523) <= (layer2_outputs(53)) and not (layer2_outputs(4322));
    layer3_outputs(3524) <= layer2_outputs(6336);
    layer3_outputs(3525) <= not((layer2_outputs(7325)) or (layer2_outputs(3146)));
    layer3_outputs(3526) <= not(layer2_outputs(5251));
    layer3_outputs(3527) <= not(layer2_outputs(4907));
    layer3_outputs(3528) <= not(layer2_outputs(6577)) or (layer2_outputs(7398));
    layer3_outputs(3529) <= layer2_outputs(2378);
    layer3_outputs(3530) <= not(layer2_outputs(6636));
    layer3_outputs(3531) <= layer2_outputs(4158);
    layer3_outputs(3532) <= not((layer2_outputs(1838)) and (layer2_outputs(5310)));
    layer3_outputs(3533) <= not((layer2_outputs(5587)) or (layer2_outputs(4524)));
    layer3_outputs(3534) <= (layer2_outputs(1860)) and not (layer2_outputs(3903));
    layer3_outputs(3535) <= (layer2_outputs(145)) xor (layer2_outputs(2007));
    layer3_outputs(3536) <= layer2_outputs(6738);
    layer3_outputs(3537) <= not((layer2_outputs(5893)) and (layer2_outputs(4218)));
    layer3_outputs(3538) <= '0';
    layer3_outputs(3539) <= not((layer2_outputs(499)) and (layer2_outputs(2950)));
    layer3_outputs(3540) <= not(layer2_outputs(1986));
    layer3_outputs(3541) <= not((layer2_outputs(1253)) or (layer2_outputs(5168)));
    layer3_outputs(3542) <= (layer2_outputs(4980)) xor (layer2_outputs(1518));
    layer3_outputs(3543) <= (layer2_outputs(7234)) and (layer2_outputs(5375));
    layer3_outputs(3544) <= not(layer2_outputs(7588));
    layer3_outputs(3545) <= (layer2_outputs(2943)) and (layer2_outputs(5796));
    layer3_outputs(3546) <= layer2_outputs(2846);
    layer3_outputs(3547) <= layer2_outputs(400);
    layer3_outputs(3548) <= not(layer2_outputs(4539)) or (layer2_outputs(1180));
    layer3_outputs(3549) <= not((layer2_outputs(3752)) and (layer2_outputs(1758)));
    layer3_outputs(3550) <= layer2_outputs(3483);
    layer3_outputs(3551) <= (layer2_outputs(1488)) and not (layer2_outputs(2712));
    layer3_outputs(3552) <= not(layer2_outputs(4752));
    layer3_outputs(3553) <= not(layer2_outputs(3093));
    layer3_outputs(3554) <= layer2_outputs(6940);
    layer3_outputs(3555) <= layer2_outputs(953);
    layer3_outputs(3556) <= not(layer2_outputs(4181));
    layer3_outputs(3557) <= not(layer2_outputs(4882));
    layer3_outputs(3558) <= (layer2_outputs(2159)) or (layer2_outputs(5807));
    layer3_outputs(3559) <= layer2_outputs(7402);
    layer3_outputs(3560) <= not(layer2_outputs(775)) or (layer2_outputs(1084));
    layer3_outputs(3561) <= not((layer2_outputs(2970)) and (layer2_outputs(6338)));
    layer3_outputs(3562) <= '1';
    layer3_outputs(3563) <= not(layer2_outputs(6686));
    layer3_outputs(3564) <= layer2_outputs(6925);
    layer3_outputs(3565) <= layer2_outputs(645);
    layer3_outputs(3566) <= not(layer2_outputs(685));
    layer3_outputs(3567) <= layer2_outputs(2095);
    layer3_outputs(3568) <= not(layer2_outputs(6470));
    layer3_outputs(3569) <= (layer2_outputs(5512)) and (layer2_outputs(117));
    layer3_outputs(3570) <= not((layer2_outputs(1876)) xor (layer2_outputs(3422)));
    layer3_outputs(3571) <= not(layer2_outputs(155));
    layer3_outputs(3572) <= '1';
    layer3_outputs(3573) <= (layer2_outputs(1486)) and not (layer2_outputs(2811));
    layer3_outputs(3574) <= layer2_outputs(4551);
    layer3_outputs(3575) <= not(layer2_outputs(2412));
    layer3_outputs(3576) <= not(layer2_outputs(1605));
    layer3_outputs(3577) <= not(layer2_outputs(1331));
    layer3_outputs(3578) <= not(layer2_outputs(3215)) or (layer2_outputs(5347));
    layer3_outputs(3579) <= not(layer2_outputs(3340));
    layer3_outputs(3580) <= layer2_outputs(836);
    layer3_outputs(3581) <= layer2_outputs(4902);
    layer3_outputs(3582) <= not(layer2_outputs(4288)) or (layer2_outputs(1858));
    layer3_outputs(3583) <= not(layer2_outputs(960));
    layer3_outputs(3584) <= not(layer2_outputs(478));
    layer3_outputs(3585) <= layer2_outputs(114);
    layer3_outputs(3586) <= not(layer2_outputs(1281));
    layer3_outputs(3587) <= not(layer2_outputs(4857));
    layer3_outputs(3588) <= layer2_outputs(565);
    layer3_outputs(3589) <= layer2_outputs(6422);
    layer3_outputs(3590) <= not(layer2_outputs(4073));
    layer3_outputs(3591) <= (layer2_outputs(3378)) and not (layer2_outputs(4723));
    layer3_outputs(3592) <= layer2_outputs(1212);
    layer3_outputs(3593) <= layer2_outputs(511);
    layer3_outputs(3594) <= (layer2_outputs(2224)) or (layer2_outputs(4756));
    layer3_outputs(3595) <= not(layer2_outputs(720));
    layer3_outputs(3596) <= not((layer2_outputs(4690)) and (layer2_outputs(5816)));
    layer3_outputs(3597) <= (layer2_outputs(3684)) xor (layer2_outputs(5499));
    layer3_outputs(3598) <= layer2_outputs(5398);
    layer3_outputs(3599) <= not((layer2_outputs(6763)) and (layer2_outputs(6814)));
    layer3_outputs(3600) <= not(layer2_outputs(559));
    layer3_outputs(3601) <= not(layer2_outputs(4041));
    layer3_outputs(3602) <= layer2_outputs(6092);
    layer3_outputs(3603) <= layer2_outputs(1770);
    layer3_outputs(3604) <= (layer2_outputs(4195)) and not (layer2_outputs(4655));
    layer3_outputs(3605) <= layer2_outputs(3193);
    layer3_outputs(3606) <= not(layer2_outputs(4231));
    layer3_outputs(3607) <= not((layer2_outputs(1391)) or (layer2_outputs(7444)));
    layer3_outputs(3608) <= layer2_outputs(6660);
    layer3_outputs(3609) <= not(layer2_outputs(2552));
    layer3_outputs(3610) <= layer2_outputs(6601);
    layer3_outputs(3611) <= not((layer2_outputs(628)) xor (layer2_outputs(3236)));
    layer3_outputs(3612) <= layer2_outputs(1732);
    layer3_outputs(3613) <= not((layer2_outputs(293)) and (layer2_outputs(4337)));
    layer3_outputs(3614) <= layer2_outputs(622);
    layer3_outputs(3615) <= not((layer2_outputs(2885)) and (layer2_outputs(6960)));
    layer3_outputs(3616) <= layer2_outputs(7228);
    layer3_outputs(3617) <= layer2_outputs(6414);
    layer3_outputs(3618) <= (layer2_outputs(3223)) and not (layer2_outputs(4290));
    layer3_outputs(3619) <= (layer2_outputs(4498)) and not (layer2_outputs(5253));
    layer3_outputs(3620) <= (layer2_outputs(268)) xor (layer2_outputs(4054));
    layer3_outputs(3621) <= not(layer2_outputs(7405));
    layer3_outputs(3622) <= not(layer2_outputs(1368)) or (layer2_outputs(2249));
    layer3_outputs(3623) <= not(layer2_outputs(5342));
    layer3_outputs(3624) <= not((layer2_outputs(4104)) and (layer2_outputs(2983)));
    layer3_outputs(3625) <= '1';
    layer3_outputs(3626) <= not((layer2_outputs(1617)) and (layer2_outputs(7287)));
    layer3_outputs(3627) <= layer2_outputs(1340);
    layer3_outputs(3628) <= not((layer2_outputs(3454)) xor (layer2_outputs(1138)));
    layer3_outputs(3629) <= not(layer2_outputs(908));
    layer3_outputs(3630) <= not(layer2_outputs(3115));
    layer3_outputs(3631) <= not(layer2_outputs(6193));
    layer3_outputs(3632) <= not(layer2_outputs(352));
    layer3_outputs(3633) <= (layer2_outputs(5005)) or (layer2_outputs(4493));
    layer3_outputs(3634) <= not(layer2_outputs(5360)) or (layer2_outputs(4575));
    layer3_outputs(3635) <= not(layer2_outputs(1232));
    layer3_outputs(3636) <= (layer2_outputs(5903)) and (layer2_outputs(1286));
    layer3_outputs(3637) <= '1';
    layer3_outputs(3638) <= (layer2_outputs(5823)) and (layer2_outputs(687));
    layer3_outputs(3639) <= not(layer2_outputs(5279)) or (layer2_outputs(3222));
    layer3_outputs(3640) <= not((layer2_outputs(6144)) and (layer2_outputs(4381)));
    layer3_outputs(3641) <= not((layer2_outputs(5514)) or (layer2_outputs(5866)));
    layer3_outputs(3642) <= (layer2_outputs(530)) xor (layer2_outputs(6783));
    layer3_outputs(3643) <= not(layer2_outputs(6090));
    layer3_outputs(3644) <= (layer2_outputs(4163)) and not (layer2_outputs(2237));
    layer3_outputs(3645) <= not(layer2_outputs(7538));
    layer3_outputs(3646) <= layer2_outputs(3892);
    layer3_outputs(3647) <= not(layer2_outputs(5243));
    layer3_outputs(3648) <= not(layer2_outputs(2044));
    layer3_outputs(3649) <= (layer2_outputs(1692)) and not (layer2_outputs(6586));
    layer3_outputs(3650) <= (layer2_outputs(3323)) and not (layer2_outputs(1644));
    layer3_outputs(3651) <= '1';
    layer3_outputs(3652) <= not(layer2_outputs(5552)) or (layer2_outputs(3410));
    layer3_outputs(3653) <= layer2_outputs(6914);
    layer3_outputs(3654) <= layer2_outputs(966);
    layer3_outputs(3655) <= layer2_outputs(3888);
    layer3_outputs(3656) <= layer2_outputs(3247);
    layer3_outputs(3657) <= (layer2_outputs(4693)) and not (layer2_outputs(2593));
    layer3_outputs(3658) <= not(layer2_outputs(3393)) or (layer2_outputs(3076));
    layer3_outputs(3659) <= layer2_outputs(2926);
    layer3_outputs(3660) <= (layer2_outputs(4941)) and (layer2_outputs(4595));
    layer3_outputs(3661) <= not(layer2_outputs(3356));
    layer3_outputs(3662) <= not((layer2_outputs(7246)) xor (layer2_outputs(5217)));
    layer3_outputs(3663) <= not(layer2_outputs(1644));
    layer3_outputs(3664) <= not((layer2_outputs(5627)) or (layer2_outputs(2536)));
    layer3_outputs(3665) <= (layer2_outputs(158)) and not (layer2_outputs(2724));
    layer3_outputs(3666) <= layer2_outputs(2837);
    layer3_outputs(3667) <= (layer2_outputs(321)) and (layer2_outputs(3168));
    layer3_outputs(3668) <= not(layer2_outputs(7249)) or (layer2_outputs(870));
    layer3_outputs(3669) <= not(layer2_outputs(325));
    layer3_outputs(3670) <= (layer2_outputs(6454)) and not (layer2_outputs(3709));
    layer3_outputs(3671) <= layer2_outputs(3997);
    layer3_outputs(3672) <= not((layer2_outputs(3184)) xor (layer2_outputs(470)));
    layer3_outputs(3673) <= not(layer2_outputs(2486)) or (layer2_outputs(5365));
    layer3_outputs(3674) <= not(layer2_outputs(1015));
    layer3_outputs(3675) <= not(layer2_outputs(5666)) or (layer2_outputs(3994));
    layer3_outputs(3676) <= not(layer2_outputs(6248));
    layer3_outputs(3677) <= not(layer2_outputs(517));
    layer3_outputs(3678) <= not((layer2_outputs(2932)) and (layer2_outputs(1429)));
    layer3_outputs(3679) <= layer2_outputs(5032);
    layer3_outputs(3680) <= not(layer2_outputs(4333));
    layer3_outputs(3681) <= (layer2_outputs(6355)) and (layer2_outputs(5837));
    layer3_outputs(3682) <= not(layer2_outputs(1887));
    layer3_outputs(3683) <= '1';
    layer3_outputs(3684) <= not(layer2_outputs(4777)) or (layer2_outputs(4070));
    layer3_outputs(3685) <= layer2_outputs(4938);
    layer3_outputs(3686) <= layer2_outputs(5404);
    layer3_outputs(3687) <= not(layer2_outputs(1411)) or (layer2_outputs(6980));
    layer3_outputs(3688) <= not((layer2_outputs(2699)) xor (layer2_outputs(1123)));
    layer3_outputs(3689) <= layer2_outputs(4615);
    layer3_outputs(3690) <= layer2_outputs(3724);
    layer3_outputs(3691) <= (layer2_outputs(3559)) and (layer2_outputs(6671));
    layer3_outputs(3692) <= (layer2_outputs(5762)) and not (layer2_outputs(2831));
    layer3_outputs(3693) <= (layer2_outputs(4990)) or (layer2_outputs(2584));
    layer3_outputs(3694) <= not(layer2_outputs(2854));
    layer3_outputs(3695) <= layer2_outputs(2206);
    layer3_outputs(3696) <= (layer2_outputs(3564)) or (layer2_outputs(1152));
    layer3_outputs(3697) <= (layer2_outputs(643)) or (layer2_outputs(2844));
    layer3_outputs(3698) <= (layer2_outputs(5568)) xor (layer2_outputs(3822));
    layer3_outputs(3699) <= (layer2_outputs(2845)) and not (layer2_outputs(4183));
    layer3_outputs(3700) <= (layer2_outputs(3746)) and (layer2_outputs(3025));
    layer3_outputs(3701) <= not(layer2_outputs(942));
    layer3_outputs(3702) <= (layer2_outputs(4326)) and (layer2_outputs(5199));
    layer3_outputs(3703) <= not((layer2_outputs(7043)) and (layer2_outputs(5290)));
    layer3_outputs(3704) <= not(layer2_outputs(3484));
    layer3_outputs(3705) <= not(layer2_outputs(5719)) or (layer2_outputs(3722));
    layer3_outputs(3706) <= '1';
    layer3_outputs(3707) <= '0';
    layer3_outputs(3708) <= not((layer2_outputs(6295)) and (layer2_outputs(2801)));
    layer3_outputs(3709) <= (layer2_outputs(5908)) and not (layer2_outputs(5509));
    layer3_outputs(3710) <= layer2_outputs(6166);
    layer3_outputs(3711) <= layer2_outputs(1531);
    layer3_outputs(3712) <= not(layer2_outputs(4747));
    layer3_outputs(3713) <= (layer2_outputs(5151)) xor (layer2_outputs(6995));
    layer3_outputs(3714) <= layer2_outputs(3274);
    layer3_outputs(3715) <= not(layer2_outputs(7187)) or (layer2_outputs(6530));
    layer3_outputs(3716) <= (layer2_outputs(476)) xor (layer2_outputs(2619));
    layer3_outputs(3717) <= not((layer2_outputs(5205)) or (layer2_outputs(3912)));
    layer3_outputs(3718) <= layer2_outputs(668);
    layer3_outputs(3719) <= (layer2_outputs(460)) or (layer2_outputs(460));
    layer3_outputs(3720) <= not(layer2_outputs(7167));
    layer3_outputs(3721) <= (layer2_outputs(4412)) or (layer2_outputs(7580));
    layer3_outputs(3722) <= not(layer2_outputs(3522));
    layer3_outputs(3723) <= '0';
    layer3_outputs(3724) <= (layer2_outputs(3111)) or (layer2_outputs(729));
    layer3_outputs(3725) <= not((layer2_outputs(7197)) or (layer2_outputs(7129)));
    layer3_outputs(3726) <= (layer2_outputs(5937)) and (layer2_outputs(5489));
    layer3_outputs(3727) <= not(layer2_outputs(5477)) or (layer2_outputs(2619));
    layer3_outputs(3728) <= not((layer2_outputs(1594)) xor (layer2_outputs(1238)));
    layer3_outputs(3729) <= layer2_outputs(2604);
    layer3_outputs(3730) <= layer2_outputs(2333);
    layer3_outputs(3731) <= (layer2_outputs(6007)) and not (layer2_outputs(4190));
    layer3_outputs(3732) <= not(layer2_outputs(4632));
    layer3_outputs(3733) <= (layer2_outputs(7309)) and not (layer2_outputs(1716));
    layer3_outputs(3734) <= layer2_outputs(2869);
    layer3_outputs(3735) <= (layer2_outputs(773)) or (layer2_outputs(3753));
    layer3_outputs(3736) <= layer2_outputs(2043);
    layer3_outputs(3737) <= (layer2_outputs(5035)) and not (layer2_outputs(2291));
    layer3_outputs(3738) <= not(layer2_outputs(3290)) or (layer2_outputs(5212));
    layer3_outputs(3739) <= not((layer2_outputs(4797)) and (layer2_outputs(6145)));
    layer3_outputs(3740) <= (layer2_outputs(2176)) or (layer2_outputs(531));
    layer3_outputs(3741) <= not(layer2_outputs(4376));
    layer3_outputs(3742) <= (layer2_outputs(4586)) and (layer2_outputs(2843));
    layer3_outputs(3743) <= layer2_outputs(2089);
    layer3_outputs(3744) <= not(layer2_outputs(44));
    layer3_outputs(3745) <= not(layer2_outputs(5688));
    layer3_outputs(3746) <= not(layer2_outputs(4697)) or (layer2_outputs(3162));
    layer3_outputs(3747) <= not(layer2_outputs(5186));
    layer3_outputs(3748) <= layer2_outputs(6906);
    layer3_outputs(3749) <= (layer2_outputs(4088)) and not (layer2_outputs(3367));
    layer3_outputs(3750) <= not(layer2_outputs(3065));
    layer3_outputs(3751) <= layer2_outputs(2965);
    layer3_outputs(3752) <= layer2_outputs(4558);
    layer3_outputs(3753) <= not(layer2_outputs(6926));
    layer3_outputs(3754) <= (layer2_outputs(2617)) xor (layer2_outputs(1634));
    layer3_outputs(3755) <= not((layer2_outputs(7496)) xor (layer2_outputs(842)));
    layer3_outputs(3756) <= not(layer2_outputs(1223)) or (layer2_outputs(1863));
    layer3_outputs(3757) <= layer2_outputs(182);
    layer3_outputs(3758) <= '1';
    layer3_outputs(3759) <= not(layer2_outputs(2361));
    layer3_outputs(3760) <= not((layer2_outputs(3102)) or (layer2_outputs(5822)));
    layer3_outputs(3761) <= (layer2_outputs(6808)) xor (layer2_outputs(3946));
    layer3_outputs(3762) <= not(layer2_outputs(4519));
    layer3_outputs(3763) <= not(layer2_outputs(5517));
    layer3_outputs(3764) <= (layer2_outputs(6994)) and (layer2_outputs(5169));
    layer3_outputs(3765) <= (layer2_outputs(126)) or (layer2_outputs(4391));
    layer3_outputs(3766) <= not((layer2_outputs(6156)) and (layer2_outputs(4139)));
    layer3_outputs(3767) <= not(layer2_outputs(7375)) or (layer2_outputs(4696));
    layer3_outputs(3768) <= (layer2_outputs(4262)) and not (layer2_outputs(5400));
    layer3_outputs(3769) <= not((layer2_outputs(2120)) or (layer2_outputs(6211)));
    layer3_outputs(3770) <= layer2_outputs(636);
    layer3_outputs(3771) <= layer2_outputs(3320);
    layer3_outputs(3772) <= (layer2_outputs(6182)) or (layer2_outputs(3860));
    layer3_outputs(3773) <= not(layer2_outputs(1844)) or (layer2_outputs(489));
    layer3_outputs(3774) <= (layer2_outputs(3991)) and not (layer2_outputs(7278));
    layer3_outputs(3775) <= not(layer2_outputs(1666));
    layer3_outputs(3776) <= (layer2_outputs(591)) and not (layer2_outputs(7481));
    layer3_outputs(3777) <= not(layer2_outputs(2179)) or (layer2_outputs(3022));
    layer3_outputs(3778) <= layer2_outputs(2513);
    layer3_outputs(3779) <= layer2_outputs(772);
    layer3_outputs(3780) <= not(layer2_outputs(6556));
    layer3_outputs(3781) <= not(layer2_outputs(697));
    layer3_outputs(3782) <= (layer2_outputs(2908)) and not (layer2_outputs(6116));
    layer3_outputs(3783) <= not((layer2_outputs(7457)) or (layer2_outputs(541)));
    layer3_outputs(3784) <= not(layer2_outputs(4859));
    layer3_outputs(3785) <= not(layer2_outputs(7053)) or (layer2_outputs(2404));
    layer3_outputs(3786) <= layer2_outputs(3499);
    layer3_outputs(3787) <= (layer2_outputs(5667)) or (layer2_outputs(2174));
    layer3_outputs(3788) <= (layer2_outputs(750)) and not (layer2_outputs(7018));
    layer3_outputs(3789) <= layer2_outputs(1396);
    layer3_outputs(3790) <= layer2_outputs(3770);
    layer3_outputs(3791) <= not(layer2_outputs(3191));
    layer3_outputs(3792) <= layer2_outputs(7081);
    layer3_outputs(3793) <= (layer2_outputs(2387)) and not (layer2_outputs(3254));
    layer3_outputs(3794) <= layer2_outputs(6299);
    layer3_outputs(3795) <= layer2_outputs(3498);
    layer3_outputs(3796) <= layer2_outputs(1116);
    layer3_outputs(3797) <= layer2_outputs(5926);
    layer3_outputs(3798) <= not(layer2_outputs(4454));
    layer3_outputs(3799) <= layer2_outputs(3464);
    layer3_outputs(3800) <= (layer2_outputs(2255)) and (layer2_outputs(4299));
    layer3_outputs(3801) <= not((layer2_outputs(5438)) and (layer2_outputs(3546)));
    layer3_outputs(3802) <= not((layer2_outputs(3758)) xor (layer2_outputs(7453)));
    layer3_outputs(3803) <= not(layer2_outputs(6927));
    layer3_outputs(3804) <= not(layer2_outputs(457)) or (layer2_outputs(4596));
    layer3_outputs(3805) <= not(layer2_outputs(5164)) or (layer2_outputs(226));
    layer3_outputs(3806) <= layer2_outputs(2172);
    layer3_outputs(3807) <= not(layer2_outputs(4516)) or (layer2_outputs(6954));
    layer3_outputs(3808) <= (layer2_outputs(3691)) and (layer2_outputs(6096));
    layer3_outputs(3809) <= layer2_outputs(5051);
    layer3_outputs(3810) <= not((layer2_outputs(5318)) and (layer2_outputs(3772)));
    layer3_outputs(3811) <= (layer2_outputs(3635)) xor (layer2_outputs(5987));
    layer3_outputs(3812) <= not((layer2_outputs(5401)) and (layer2_outputs(7474)));
    layer3_outputs(3813) <= (layer2_outputs(6682)) or (layer2_outputs(475));
    layer3_outputs(3814) <= not(layer2_outputs(5282)) or (layer2_outputs(3316));
    layer3_outputs(3815) <= layer2_outputs(4708);
    layer3_outputs(3816) <= not((layer2_outputs(3344)) xor (layer2_outputs(2252)));
    layer3_outputs(3817) <= (layer2_outputs(4018)) and not (layer2_outputs(5669));
    layer3_outputs(3818) <= not(layer2_outputs(6370));
    layer3_outputs(3819) <= not(layer2_outputs(7480)) or (layer2_outputs(4871));
    layer3_outputs(3820) <= (layer2_outputs(596)) and not (layer2_outputs(1725));
    layer3_outputs(3821) <= layer2_outputs(6517);
    layer3_outputs(3822) <= (layer2_outputs(1030)) or (layer2_outputs(615));
    layer3_outputs(3823) <= layer2_outputs(6935);
    layer3_outputs(3824) <= layer2_outputs(4591);
    layer3_outputs(3825) <= not(layer2_outputs(2880));
    layer3_outputs(3826) <= layer2_outputs(2945);
    layer3_outputs(3827) <= (layer2_outputs(7641)) and (layer2_outputs(3657));
    layer3_outputs(3828) <= (layer2_outputs(7091)) and not (layer2_outputs(6590));
    layer3_outputs(3829) <= not(layer2_outputs(4686)) or (layer2_outputs(4066));
    layer3_outputs(3830) <= not(layer2_outputs(6864));
    layer3_outputs(3831) <= (layer2_outputs(5487)) and not (layer2_outputs(3144));
    layer3_outputs(3832) <= (layer2_outputs(1050)) and not (layer2_outputs(6187));
    layer3_outputs(3833) <= not(layer2_outputs(1724));
    layer3_outputs(3834) <= not(layer2_outputs(1342));
    layer3_outputs(3835) <= layer2_outputs(473);
    layer3_outputs(3836) <= not(layer2_outputs(6048));
    layer3_outputs(3837) <= (layer2_outputs(1329)) and not (layer2_outputs(7188));
    layer3_outputs(3838) <= not(layer2_outputs(1218));
    layer3_outputs(3839) <= not(layer2_outputs(6565));
    layer3_outputs(3840) <= not(layer2_outputs(5258)) or (layer2_outputs(782));
    layer3_outputs(3841) <= not(layer2_outputs(6691)) or (layer2_outputs(3359));
    layer3_outputs(3842) <= layer2_outputs(3096);
    layer3_outputs(3843) <= not(layer2_outputs(3561)) or (layer2_outputs(6344));
    layer3_outputs(3844) <= not(layer2_outputs(3408));
    layer3_outputs(3845) <= not(layer2_outputs(3004));
    layer3_outputs(3846) <= not(layer2_outputs(2836)) or (layer2_outputs(5814));
    layer3_outputs(3847) <= not(layer2_outputs(162));
    layer3_outputs(3848) <= not(layer2_outputs(6045));
    layer3_outputs(3849) <= layer2_outputs(3002);
    layer3_outputs(3850) <= (layer2_outputs(1492)) and not (layer2_outputs(104));
    layer3_outputs(3851) <= not(layer2_outputs(6057));
    layer3_outputs(3852) <= layer2_outputs(2595);
    layer3_outputs(3853) <= layer2_outputs(501);
    layer3_outputs(3854) <= not(layer2_outputs(3399));
    layer3_outputs(3855) <= not((layer2_outputs(3698)) and (layer2_outputs(4670)));
    layer3_outputs(3856) <= (layer2_outputs(5432)) or (layer2_outputs(3866));
    layer3_outputs(3857) <= '1';
    layer3_outputs(3858) <= not(layer2_outputs(5897)) or (layer2_outputs(7662));
    layer3_outputs(3859) <= (layer2_outputs(569)) xor (layer2_outputs(6475));
    layer3_outputs(3860) <= layer2_outputs(5685);
    layer3_outputs(3861) <= layer2_outputs(4843);
    layer3_outputs(3862) <= (layer2_outputs(1095)) and (layer2_outputs(4543));
    layer3_outputs(3863) <= not((layer2_outputs(7031)) or (layer2_outputs(1227)));
    layer3_outputs(3864) <= not((layer2_outputs(355)) and (layer2_outputs(811)));
    layer3_outputs(3865) <= (layer2_outputs(756)) and (layer2_outputs(3725));
    layer3_outputs(3866) <= not((layer2_outputs(4020)) and (layer2_outputs(6496)));
    layer3_outputs(3867) <= not(layer2_outputs(2516));
    layer3_outputs(3868) <= not(layer2_outputs(7421));
    layer3_outputs(3869) <= not(layer2_outputs(733)) or (layer2_outputs(7212));
    layer3_outputs(3870) <= (layer2_outputs(3944)) or (layer2_outputs(3277));
    layer3_outputs(3871) <= (layer2_outputs(3671)) and (layer2_outputs(5014));
    layer3_outputs(3872) <= (layer2_outputs(589)) and not (layer2_outputs(6545));
    layer3_outputs(3873) <= not(layer2_outputs(695));
    layer3_outputs(3874) <= (layer2_outputs(2363)) or (layer2_outputs(524));
    layer3_outputs(3875) <= not(layer2_outputs(4671));
    layer3_outputs(3876) <= layer2_outputs(188);
    layer3_outputs(3877) <= layer2_outputs(7469);
    layer3_outputs(3878) <= (layer2_outputs(689)) and (layer2_outputs(6235));
    layer3_outputs(3879) <= not(layer2_outputs(6259));
    layer3_outputs(3880) <= (layer2_outputs(5744)) and (layer2_outputs(831));
    layer3_outputs(3881) <= not((layer2_outputs(6600)) and (layer2_outputs(2640)));
    layer3_outputs(3882) <= (layer2_outputs(1682)) or (layer2_outputs(2058));
    layer3_outputs(3883) <= not(layer2_outputs(1102));
    layer3_outputs(3884) <= layer2_outputs(3398);
    layer3_outputs(3885) <= not(layer2_outputs(204));
    layer3_outputs(3886) <= (layer2_outputs(605)) and (layer2_outputs(3392));
    layer3_outputs(3887) <= layer2_outputs(3194);
    layer3_outputs(3888) <= layer2_outputs(4891);
    layer3_outputs(3889) <= layer2_outputs(5634);
    layer3_outputs(3890) <= not((layer2_outputs(5630)) or (layer2_outputs(6418)));
    layer3_outputs(3891) <= layer2_outputs(4765);
    layer3_outputs(3892) <= not(layer2_outputs(5434)) or (layer2_outputs(3631));
    layer3_outputs(3893) <= not((layer2_outputs(1879)) or (layer2_outputs(3973)));
    layer3_outputs(3894) <= (layer2_outputs(6343)) or (layer2_outputs(5420));
    layer3_outputs(3895) <= not(layer2_outputs(6872));
    layer3_outputs(3896) <= not((layer2_outputs(7629)) or (layer2_outputs(268)));
    layer3_outputs(3897) <= (layer2_outputs(3245)) and (layer2_outputs(5764));
    layer3_outputs(3898) <= not(layer2_outputs(1538)) or (layer2_outputs(5566));
    layer3_outputs(3899) <= layer2_outputs(7304);
    layer3_outputs(3900) <= not(layer2_outputs(3533));
    layer3_outputs(3901) <= '0';
    layer3_outputs(3902) <= not(layer2_outputs(5675));
    layer3_outputs(3903) <= (layer2_outputs(6915)) and not (layer2_outputs(2166));
    layer3_outputs(3904) <= layer2_outputs(5447);
    layer3_outputs(3905) <= not(layer2_outputs(1248));
    layer3_outputs(3906) <= layer2_outputs(952);
    layer3_outputs(3907) <= (layer2_outputs(3216)) and (layer2_outputs(4657));
    layer3_outputs(3908) <= not((layer2_outputs(4607)) or (layer2_outputs(4950)));
    layer3_outputs(3909) <= not(layer2_outputs(7047));
    layer3_outputs(3910) <= (layer2_outputs(4142)) and not (layer2_outputs(87));
    layer3_outputs(3911) <= not((layer2_outputs(7413)) or (layer2_outputs(3112)));
    layer3_outputs(3912) <= (layer2_outputs(2706)) and not (layer2_outputs(3129));
    layer3_outputs(3913) <= not(layer2_outputs(1663));
    layer3_outputs(3914) <= layer2_outputs(903);
    layer3_outputs(3915) <= layer2_outputs(86);
    layer3_outputs(3916) <= not(layer2_outputs(284));
    layer3_outputs(3917) <= (layer2_outputs(7075)) and (layer2_outputs(6505));
    layer3_outputs(3918) <= layer2_outputs(5359);
    layer3_outputs(3919) <= (layer2_outputs(6200)) and not (layer2_outputs(7067));
    layer3_outputs(3920) <= not(layer2_outputs(2490)) or (layer2_outputs(3823));
    layer3_outputs(3921) <= layer2_outputs(424);
    layer3_outputs(3922) <= not(layer2_outputs(1900));
    layer3_outputs(3923) <= (layer2_outputs(5857)) and not (layer2_outputs(1758));
    layer3_outputs(3924) <= not(layer2_outputs(84));
    layer3_outputs(3925) <= not(layer2_outputs(1871));
    layer3_outputs(3926) <= not(layer2_outputs(4180));
    layer3_outputs(3927) <= (layer2_outputs(1834)) xor (layer2_outputs(1102));
    layer3_outputs(3928) <= not(layer2_outputs(3213));
    layer3_outputs(3929) <= not(layer2_outputs(6219)) or (layer2_outputs(2366));
    layer3_outputs(3930) <= (layer2_outputs(4258)) and (layer2_outputs(680));
    layer3_outputs(3931) <= layer2_outputs(3443);
    layer3_outputs(3932) <= (layer2_outputs(2015)) and (layer2_outputs(2181));
    layer3_outputs(3933) <= not(layer2_outputs(1519));
    layer3_outputs(3934) <= not((layer2_outputs(3826)) and (layer2_outputs(3274)));
    layer3_outputs(3935) <= (layer2_outputs(3120)) and not (layer2_outputs(7239));
    layer3_outputs(3936) <= layer2_outputs(1212);
    layer3_outputs(3937) <= not(layer2_outputs(766));
    layer3_outputs(3938) <= (layer2_outputs(7472)) xor (layer2_outputs(4726));
    layer3_outputs(3939) <= not(layer2_outputs(4195));
    layer3_outputs(3940) <= layer2_outputs(4418);
    layer3_outputs(3941) <= layer2_outputs(7311);
    layer3_outputs(3942) <= (layer2_outputs(2543)) and (layer2_outputs(6663));
    layer3_outputs(3943) <= not(layer2_outputs(1612));
    layer3_outputs(3944) <= (layer2_outputs(2214)) and (layer2_outputs(3666));
    layer3_outputs(3945) <= '0';
    layer3_outputs(3946) <= (layer2_outputs(4100)) xor (layer2_outputs(1883));
    layer3_outputs(3947) <= layer2_outputs(6963);
    layer3_outputs(3948) <= layer2_outputs(5998);
    layer3_outputs(3949) <= (layer2_outputs(3981)) and not (layer2_outputs(7394));
    layer3_outputs(3950) <= layer2_outputs(6655);
    layer3_outputs(3951) <= '0';
    layer3_outputs(3952) <= (layer2_outputs(7124)) and (layer2_outputs(1029));
    layer3_outputs(3953) <= not(layer2_outputs(431));
    layer3_outputs(3954) <= (layer2_outputs(6654)) and not (layer2_outputs(2688));
    layer3_outputs(3955) <= not(layer2_outputs(1864));
    layer3_outputs(3956) <= '0';
    layer3_outputs(3957) <= not((layer2_outputs(3474)) and (layer2_outputs(7249)));
    layer3_outputs(3958) <= layer2_outputs(1464);
    layer3_outputs(3959) <= not(layer2_outputs(3044)) or (layer2_outputs(6786));
    layer3_outputs(3960) <= (layer2_outputs(6890)) xor (layer2_outputs(4529));
    layer3_outputs(3961) <= layer2_outputs(4174);
    layer3_outputs(3962) <= not(layer2_outputs(6986));
    layer3_outputs(3963) <= (layer2_outputs(6364)) xor (layer2_outputs(3679));
    layer3_outputs(3964) <= not((layer2_outputs(724)) and (layer2_outputs(4643)));
    layer3_outputs(3965) <= not((layer2_outputs(7656)) and (layer2_outputs(2321)));
    layer3_outputs(3966) <= not(layer2_outputs(5739));
    layer3_outputs(3967) <= not(layer2_outputs(489));
    layer3_outputs(3968) <= not(layer2_outputs(7356));
    layer3_outputs(3969) <= not(layer2_outputs(629));
    layer3_outputs(3970) <= not((layer2_outputs(4)) or (layer2_outputs(803)));
    layer3_outputs(3971) <= (layer2_outputs(844)) xor (layer2_outputs(2408));
    layer3_outputs(3972) <= not(layer2_outputs(6125)) or (layer2_outputs(3674));
    layer3_outputs(3973) <= layer2_outputs(4323);
    layer3_outputs(3974) <= not(layer2_outputs(2602)) or (layer2_outputs(4852));
    layer3_outputs(3975) <= not((layer2_outputs(3631)) or (layer2_outputs(5490)));
    layer3_outputs(3976) <= not(layer2_outputs(6300));
    layer3_outputs(3977) <= not(layer2_outputs(6562));
    layer3_outputs(3978) <= not(layer2_outputs(6894)) or (layer2_outputs(1823));
    layer3_outputs(3979) <= not((layer2_outputs(2401)) or (layer2_outputs(2156)));
    layer3_outputs(3980) <= not(layer2_outputs(7445));
    layer3_outputs(3981) <= layer2_outputs(7058);
    layer3_outputs(3982) <= not(layer2_outputs(5957));
    layer3_outputs(3983) <= (layer2_outputs(1201)) and not (layer2_outputs(4963));
    layer3_outputs(3984) <= not((layer2_outputs(6404)) or (layer2_outputs(5123)));
    layer3_outputs(3985) <= not(layer2_outputs(6081));
    layer3_outputs(3986) <= (layer2_outputs(1907)) and not (layer2_outputs(5846));
    layer3_outputs(3987) <= layer2_outputs(2114);
    layer3_outputs(3988) <= not(layer2_outputs(1819)) or (layer2_outputs(3838));
    layer3_outputs(3989) <= (layer2_outputs(7079)) and (layer2_outputs(5467));
    layer3_outputs(3990) <= (layer2_outputs(1336)) and (layer2_outputs(5707));
    layer3_outputs(3991) <= not((layer2_outputs(1414)) and (layer2_outputs(6785)));
    layer3_outputs(3992) <= not(layer2_outputs(484));
    layer3_outputs(3993) <= (layer2_outputs(274)) and not (layer2_outputs(4561));
    layer3_outputs(3994) <= not(layer2_outputs(2860)) or (layer2_outputs(2275));
    layer3_outputs(3995) <= layer2_outputs(7314);
    layer3_outputs(3996) <= layer2_outputs(715);
    layer3_outputs(3997) <= not(layer2_outputs(5317)) or (layer2_outputs(3069));
    layer3_outputs(3998) <= layer2_outputs(282);
    layer3_outputs(3999) <= not(layer2_outputs(4361));
    layer3_outputs(4000) <= '1';
    layer3_outputs(4001) <= not(layer2_outputs(7625));
    layer3_outputs(4002) <= not(layer2_outputs(1296));
    layer3_outputs(4003) <= (layer2_outputs(7549)) and not (layer2_outputs(4382));
    layer3_outputs(4004) <= (layer2_outputs(1149)) and not (layer2_outputs(7553));
    layer3_outputs(4005) <= not(layer2_outputs(105));
    layer3_outputs(4006) <= not(layer2_outputs(6345)) or (layer2_outputs(6381));
    layer3_outputs(4007) <= layer2_outputs(1911);
    layer3_outputs(4008) <= layer2_outputs(6624);
    layer3_outputs(4009) <= (layer2_outputs(58)) and not (layer2_outputs(499));
    layer3_outputs(4010) <= '0';
    layer3_outputs(4011) <= not(layer2_outputs(3247));
    layer3_outputs(4012) <= layer2_outputs(1225);
    layer3_outputs(4013) <= not(layer2_outputs(6149));
    layer3_outputs(4014) <= layer2_outputs(4457);
    layer3_outputs(4015) <= not((layer2_outputs(1413)) or (layer2_outputs(4203)));
    layer3_outputs(4016) <= (layer2_outputs(6341)) and not (layer2_outputs(4898));
    layer3_outputs(4017) <= not((layer2_outputs(922)) and (layer2_outputs(6264)));
    layer3_outputs(4018) <= (layer2_outputs(6273)) and not (layer2_outputs(1311));
    layer3_outputs(4019) <= layer2_outputs(5079);
    layer3_outputs(4020) <= not((layer2_outputs(6190)) or (layer2_outputs(6417)));
    layer3_outputs(4021) <= not(layer2_outputs(2916));
    layer3_outputs(4022) <= not((layer2_outputs(690)) xor (layer2_outputs(3236)));
    layer3_outputs(4023) <= not(layer2_outputs(6303));
    layer3_outputs(4024) <= (layer2_outputs(5205)) and not (layer2_outputs(5145));
    layer3_outputs(4025) <= layer2_outputs(3228);
    layer3_outputs(4026) <= not(layer2_outputs(4774));
    layer3_outputs(4027) <= layer2_outputs(1432);
    layer3_outputs(4028) <= layer2_outputs(4323);
    layer3_outputs(4029) <= not(layer2_outputs(6082)) or (layer2_outputs(5012));
    layer3_outputs(4030) <= layer2_outputs(2893);
    layer3_outputs(4031) <= layer2_outputs(7322);
    layer3_outputs(4032) <= layer2_outputs(6611);
    layer3_outputs(4033) <= not(layer2_outputs(3010)) or (layer2_outputs(5792));
    layer3_outputs(4034) <= not(layer2_outputs(2898));
    layer3_outputs(4035) <= (layer2_outputs(6664)) and (layer2_outputs(5343));
    layer3_outputs(4036) <= not(layer2_outputs(5092));
    layer3_outputs(4037) <= layer2_outputs(2067);
    layer3_outputs(4038) <= layer2_outputs(7613);
    layer3_outputs(4039) <= (layer2_outputs(7448)) and not (layer2_outputs(7336));
    layer3_outputs(4040) <= not(layer2_outputs(5304));
    layer3_outputs(4041) <= (layer2_outputs(6845)) and not (layer2_outputs(2461));
    layer3_outputs(4042) <= not((layer2_outputs(4200)) xor (layer2_outputs(7072)));
    layer3_outputs(4043) <= not(layer2_outputs(2638)) or (layer2_outputs(2102));
    layer3_outputs(4044) <= not((layer2_outputs(2152)) and (layer2_outputs(6129)));
    layer3_outputs(4045) <= not(layer2_outputs(264));
    layer3_outputs(4046) <= not((layer2_outputs(40)) or (layer2_outputs(2243)));
    layer3_outputs(4047) <= not((layer2_outputs(7159)) and (layer2_outputs(1035)));
    layer3_outputs(4048) <= not(layer2_outputs(706));
    layer3_outputs(4049) <= not(layer2_outputs(6970));
    layer3_outputs(4050) <= layer2_outputs(3909);
    layer3_outputs(4051) <= (layer2_outputs(1680)) and not (layer2_outputs(5767));
    layer3_outputs(4052) <= not(layer2_outputs(6866)) or (layer2_outputs(6956));
    layer3_outputs(4053) <= not(layer2_outputs(974)) or (layer2_outputs(1060));
    layer3_outputs(4054) <= not((layer2_outputs(1931)) or (layer2_outputs(4770)));
    layer3_outputs(4055) <= layer2_outputs(4048);
    layer3_outputs(4056) <= not(layer2_outputs(6257));
    layer3_outputs(4057) <= layer2_outputs(3441);
    layer3_outputs(4058) <= not(layer2_outputs(764)) or (layer2_outputs(6610));
    layer3_outputs(4059) <= not(layer2_outputs(3688));
    layer3_outputs(4060) <= '1';
    layer3_outputs(4061) <= (layer2_outputs(4753)) and (layer2_outputs(7045));
    layer3_outputs(4062) <= not((layer2_outputs(7001)) and (layer2_outputs(5057)));
    layer3_outputs(4063) <= (layer2_outputs(7483)) or (layer2_outputs(2575));
    layer3_outputs(4064) <= layer2_outputs(6099);
    layer3_outputs(4065) <= (layer2_outputs(4017)) or (layer2_outputs(5719));
    layer3_outputs(4066) <= (layer2_outputs(1471)) or (layer2_outputs(3842));
    layer3_outputs(4067) <= not((layer2_outputs(1434)) and (layer2_outputs(2721)));
    layer3_outputs(4068) <= not(layer2_outputs(6951));
    layer3_outputs(4069) <= not(layer2_outputs(3744));
    layer3_outputs(4070) <= (layer2_outputs(3828)) and not (layer2_outputs(7328));
    layer3_outputs(4071) <= not(layer2_outputs(1364));
    layer3_outputs(4072) <= (layer2_outputs(19)) xor (layer2_outputs(7635));
    layer3_outputs(4073) <= (layer2_outputs(7585)) and not (layer2_outputs(7004));
    layer3_outputs(4074) <= layer2_outputs(2964);
    layer3_outputs(4075) <= not(layer2_outputs(563)) or (layer2_outputs(6063));
    layer3_outputs(4076) <= not((layer2_outputs(4325)) xor (layer2_outputs(42)));
    layer3_outputs(4077) <= (layer2_outputs(2810)) or (layer2_outputs(5441));
    layer3_outputs(4078) <= layer2_outputs(5140);
    layer3_outputs(4079) <= (layer2_outputs(6741)) and (layer2_outputs(2774));
    layer3_outputs(4080) <= (layer2_outputs(426)) or (layer2_outputs(6025));
    layer3_outputs(4081) <= (layer2_outputs(4908)) and (layer2_outputs(5191));
    layer3_outputs(4082) <= (layer2_outputs(7095)) and not (layer2_outputs(2542));
    layer3_outputs(4083) <= not(layer2_outputs(1168)) or (layer2_outputs(2633));
    layer3_outputs(4084) <= not(layer2_outputs(1969));
    layer3_outputs(4085) <= not(layer2_outputs(4631)) or (layer2_outputs(1263));
    layer3_outputs(4086) <= (layer2_outputs(5674)) or (layer2_outputs(4331));
    layer3_outputs(4087) <= not(layer2_outputs(5237)) or (layer2_outputs(5608));
    layer3_outputs(4088) <= (layer2_outputs(2016)) and (layer2_outputs(5288));
    layer3_outputs(4089) <= (layer2_outputs(4184)) and (layer2_outputs(2366));
    layer3_outputs(4090) <= (layer2_outputs(1750)) or (layer2_outputs(2669));
    layer3_outputs(4091) <= not(layer2_outputs(2903));
    layer3_outputs(4092) <= (layer2_outputs(6807)) and (layer2_outputs(5080));
    layer3_outputs(4093) <= (layer2_outputs(4609)) or (layer2_outputs(2917));
    layer3_outputs(4094) <= not(layer2_outputs(814)) or (layer2_outputs(4793));
    layer3_outputs(4095) <= (layer2_outputs(1454)) xor (layer2_outputs(6564));
    layer3_outputs(4096) <= (layer2_outputs(7390)) and not (layer2_outputs(7590));
    layer3_outputs(4097) <= layer2_outputs(7430);
    layer3_outputs(4098) <= (layer2_outputs(2389)) and (layer2_outputs(883));
    layer3_outputs(4099) <= not(layer2_outputs(4927)) or (layer2_outputs(2714));
    layer3_outputs(4100) <= not(layer2_outputs(3627));
    layer3_outputs(4101) <= (layer2_outputs(3497)) and (layer2_outputs(4552));
    layer3_outputs(4102) <= not(layer2_outputs(3691));
    layer3_outputs(4103) <= (layer2_outputs(1327)) or (layer2_outputs(4783));
    layer3_outputs(4104) <= not(layer2_outputs(6245)) or (layer2_outputs(3200));
    layer3_outputs(4105) <= layer2_outputs(4176);
    layer3_outputs(4106) <= not(layer2_outputs(389));
    layer3_outputs(4107) <= not((layer2_outputs(5082)) or (layer2_outputs(4327)));
    layer3_outputs(4108) <= (layer2_outputs(2905)) and not (layer2_outputs(1150));
    layer3_outputs(4109) <= not((layer2_outputs(3525)) or (layer2_outputs(1481)));
    layer3_outputs(4110) <= '0';
    layer3_outputs(4111) <= (layer2_outputs(7132)) or (layer2_outputs(5223));
    layer3_outputs(4112) <= (layer2_outputs(5786)) and (layer2_outputs(221));
    layer3_outputs(4113) <= (layer2_outputs(5940)) and not (layer2_outputs(7069));
    layer3_outputs(4114) <= layer2_outputs(5152);
    layer3_outputs(4115) <= not(layer2_outputs(6727));
    layer3_outputs(4116) <= layer2_outputs(611);
    layer3_outputs(4117) <= not((layer2_outputs(6196)) or (layer2_outputs(1098)));
    layer3_outputs(4118) <= not(layer2_outputs(3704));
    layer3_outputs(4119) <= not(layer2_outputs(1888));
    layer3_outputs(4120) <= not(layer2_outputs(3423));
    layer3_outputs(4121) <= not((layer2_outputs(3088)) or (layer2_outputs(3035)));
    layer3_outputs(4122) <= layer2_outputs(2558);
    layer3_outputs(4123) <= not(layer2_outputs(5444));
    layer3_outputs(4124) <= layer2_outputs(2538);
    layer3_outputs(4125) <= not(layer2_outputs(7102));
    layer3_outputs(4126) <= (layer2_outputs(1655)) and not (layer2_outputs(7343));
    layer3_outputs(4127) <= layer2_outputs(2954);
    layer3_outputs(4128) <= not((layer2_outputs(1766)) xor (layer2_outputs(661)));
    layer3_outputs(4129) <= not(layer2_outputs(832));
    layer3_outputs(4130) <= (layer2_outputs(6127)) xor (layer2_outputs(5916));
    layer3_outputs(4131) <= not(layer2_outputs(1420));
    layer3_outputs(4132) <= (layer2_outputs(1056)) and not (layer2_outputs(5947));
    layer3_outputs(4133) <= layer2_outputs(4588);
    layer3_outputs(4134) <= not(layer2_outputs(7535));
    layer3_outputs(4135) <= layer2_outputs(1693);
    layer3_outputs(4136) <= not(layer2_outputs(2643));
    layer3_outputs(4137) <= not(layer2_outputs(725));
    layer3_outputs(4138) <= not((layer2_outputs(1380)) or (layer2_outputs(4826)));
    layer3_outputs(4139) <= '0';
    layer3_outputs(4140) <= layer2_outputs(3818);
    layer3_outputs(4141) <= (layer2_outputs(4230)) xor (layer2_outputs(4337));
    layer3_outputs(4142) <= not((layer2_outputs(1266)) xor (layer2_outputs(2431)));
    layer3_outputs(4143) <= layer2_outputs(3431);
    layer3_outputs(4144) <= not(layer2_outputs(178));
    layer3_outputs(4145) <= not((layer2_outputs(5088)) or (layer2_outputs(7348)));
    layer3_outputs(4146) <= not(layer2_outputs(2591));
    layer3_outputs(4147) <= not(layer2_outputs(919));
    layer3_outputs(4148) <= not(layer2_outputs(2596)) or (layer2_outputs(5366));
    layer3_outputs(4149) <= not(layer2_outputs(5850)) or (layer2_outputs(3492));
    layer3_outputs(4150) <= layer2_outputs(566);
    layer3_outputs(4151) <= not(layer2_outputs(4523));
    layer3_outputs(4152) <= layer2_outputs(3195);
    layer3_outputs(4153) <= not(layer2_outputs(1261));
    layer3_outputs(4154) <= layer2_outputs(6900);
    layer3_outputs(4155) <= not(layer2_outputs(2981));
    layer3_outputs(4156) <= (layer2_outputs(5847)) and not (layer2_outputs(164));
    layer3_outputs(4157) <= not(layer2_outputs(3931)) or (layer2_outputs(438));
    layer3_outputs(4158) <= layer2_outputs(4125);
    layer3_outputs(4159) <= not(layer2_outputs(789));
    layer3_outputs(4160) <= not(layer2_outputs(1310));
    layer3_outputs(4161) <= layer2_outputs(4301);
    layer3_outputs(4162) <= layer2_outputs(1955);
    layer3_outputs(4163) <= (layer2_outputs(2551)) and (layer2_outputs(4591));
    layer3_outputs(4164) <= '0';
    layer3_outputs(4165) <= layer2_outputs(3622);
    layer3_outputs(4166) <= not((layer2_outputs(1813)) or (layer2_outputs(6930)));
    layer3_outputs(4167) <= layer2_outputs(6134);
    layer3_outputs(4168) <= layer2_outputs(3572);
    layer3_outputs(4169) <= not((layer2_outputs(3479)) or (layer2_outputs(2359)));
    layer3_outputs(4170) <= (layer2_outputs(6981)) or (layer2_outputs(304));
    layer3_outputs(4171) <= not((layer2_outputs(1445)) xor (layer2_outputs(4466)));
    layer3_outputs(4172) <= (layer2_outputs(2676)) and (layer2_outputs(7002));
    layer3_outputs(4173) <= layer2_outputs(3719);
    layer3_outputs(4174) <= not(layer2_outputs(6172)) or (layer2_outputs(770));
    layer3_outputs(4175) <= (layer2_outputs(4809)) and not (layer2_outputs(5044));
    layer3_outputs(4176) <= (layer2_outputs(4436)) and not (layer2_outputs(564));
    layer3_outputs(4177) <= not(layer2_outputs(4675)) or (layer2_outputs(3441));
    layer3_outputs(4178) <= not(layer2_outputs(3879));
    layer3_outputs(4179) <= not(layer2_outputs(6520));
    layer3_outputs(4180) <= not((layer2_outputs(1609)) or (layer2_outputs(7131)));
    layer3_outputs(4181) <= (layer2_outputs(466)) and not (layer2_outputs(6625));
    layer3_outputs(4182) <= not(layer2_outputs(3947));
    layer3_outputs(4183) <= not(layer2_outputs(1242));
    layer3_outputs(4184) <= layer2_outputs(2971);
    layer3_outputs(4185) <= (layer2_outputs(868)) and not (layer2_outputs(5294));
    layer3_outputs(4186) <= (layer2_outputs(279)) and not (layer2_outputs(1855));
    layer3_outputs(4187) <= (layer2_outputs(1718)) and not (layer2_outputs(4276));
    layer3_outputs(4188) <= not(layer2_outputs(1931));
    layer3_outputs(4189) <= layer2_outputs(3136);
    layer3_outputs(4190) <= not(layer2_outputs(1689));
    layer3_outputs(4191) <= '1';
    layer3_outputs(4192) <= layer2_outputs(5461);
    layer3_outputs(4193) <= not(layer2_outputs(6690));
    layer3_outputs(4194) <= not((layer2_outputs(5338)) and (layer2_outputs(955)));
    layer3_outputs(4195) <= (layer2_outputs(339)) and (layer2_outputs(6250));
    layer3_outputs(4196) <= not(layer2_outputs(4120));
    layer3_outputs(4197) <= (layer2_outputs(2050)) and not (layer2_outputs(4830));
    layer3_outputs(4198) <= layer2_outputs(1195);
    layer3_outputs(4199) <= (layer2_outputs(4375)) and not (layer2_outputs(243));
    layer3_outputs(4200) <= not(layer2_outputs(1648)) or (layer2_outputs(5613));
    layer3_outputs(4201) <= (layer2_outputs(6106)) and not (layer2_outputs(5972));
    layer3_outputs(4202) <= (layer2_outputs(6060)) or (layer2_outputs(2096));
    layer3_outputs(4203) <= layer2_outputs(3640);
    layer3_outputs(4204) <= not((layer2_outputs(124)) xor (layer2_outputs(3365)));
    layer3_outputs(4205) <= not(layer2_outputs(3942));
    layer3_outputs(4206) <= (layer2_outputs(2904)) or (layer2_outputs(7270));
    layer3_outputs(4207) <= '1';
    layer3_outputs(4208) <= not((layer2_outputs(6392)) xor (layer2_outputs(5335)));
    layer3_outputs(4209) <= (layer2_outputs(1981)) and not (layer2_outputs(5070));
    layer3_outputs(4210) <= not(layer2_outputs(1945)) or (layer2_outputs(5818));
    layer3_outputs(4211) <= not(layer2_outputs(2439)) or (layer2_outputs(6044));
    layer3_outputs(4212) <= not(layer2_outputs(1951));
    layer3_outputs(4213) <= (layer2_outputs(3793)) or (layer2_outputs(6358));
    layer3_outputs(4214) <= layer2_outputs(456);
    layer3_outputs(4215) <= (layer2_outputs(2440)) and not (layer2_outputs(818));
    layer3_outputs(4216) <= not(layer2_outputs(2208));
    layer3_outputs(4217) <= layer2_outputs(1259);
    layer3_outputs(4218) <= (layer2_outputs(1943)) and not (layer2_outputs(6208));
    layer3_outputs(4219) <= layer2_outputs(1773);
    layer3_outputs(4220) <= not(layer2_outputs(6114));
    layer3_outputs(4221) <= not(layer2_outputs(2092));
    layer3_outputs(4222) <= not(layer2_outputs(4087));
    layer3_outputs(4223) <= not(layer2_outputs(5314)) or (layer2_outputs(4053));
    layer3_outputs(4224) <= (layer2_outputs(7225)) and not (layer2_outputs(4935));
    layer3_outputs(4225) <= (layer2_outputs(3218)) xor (layer2_outputs(1381));
    layer3_outputs(4226) <= not(layer2_outputs(4810)) or (layer2_outputs(3753));
    layer3_outputs(4227) <= layer2_outputs(7103);
    layer3_outputs(4228) <= (layer2_outputs(1365)) or (layer2_outputs(2250));
    layer3_outputs(4229) <= not(layer2_outputs(5523)) or (layer2_outputs(6391));
    layer3_outputs(4230) <= layer2_outputs(66);
    layer3_outputs(4231) <= not((layer2_outputs(6183)) xor (layer2_outputs(6002)));
    layer3_outputs(4232) <= layer2_outputs(4229);
    layer3_outputs(4233) <= not(layer2_outputs(6924));
    layer3_outputs(4234) <= not(layer2_outputs(3669));
    layer3_outputs(4235) <= (layer2_outputs(96)) and (layer2_outputs(6000));
    layer3_outputs(4236) <= (layer2_outputs(345)) or (layer2_outputs(7663));
    layer3_outputs(4237) <= not(layer2_outputs(4093)) or (layer2_outputs(4964));
    layer3_outputs(4238) <= (layer2_outputs(5406)) and not (layer2_outputs(6619));
    layer3_outputs(4239) <= not(layer2_outputs(716));
    layer3_outputs(4240) <= (layer2_outputs(4755)) and (layer2_outputs(6823));
    layer3_outputs(4241) <= layer2_outputs(5513);
    layer3_outputs(4242) <= not(layer2_outputs(7550));
    layer3_outputs(4243) <= not((layer2_outputs(2443)) or (layer2_outputs(5416)));
    layer3_outputs(4244) <= layer2_outputs(269);
    layer3_outputs(4245) <= layer2_outputs(4793);
    layer3_outputs(4246) <= '0';
    layer3_outputs(4247) <= layer2_outputs(3548);
    layer3_outputs(4248) <= not(layer2_outputs(614)) or (layer2_outputs(3598));
    layer3_outputs(4249) <= not((layer2_outputs(3934)) and (layer2_outputs(7577)));
    layer3_outputs(4250) <= layer2_outputs(5888);
    layer3_outputs(4251) <= layer2_outputs(1647);
    layer3_outputs(4252) <= layer2_outputs(7383);
    layer3_outputs(4253) <= (layer2_outputs(3277)) xor (layer2_outputs(194));
    layer3_outputs(4254) <= layer2_outputs(1755);
    layer3_outputs(4255) <= not(layer2_outputs(1004));
    layer3_outputs(4256) <= not(layer2_outputs(7137));
    layer3_outputs(4257) <= (layer2_outputs(3218)) and (layer2_outputs(6938));
    layer3_outputs(4258) <= not(layer2_outputs(6507));
    layer3_outputs(4259) <= not(layer2_outputs(7570)) or (layer2_outputs(501));
    layer3_outputs(4260) <= (layer2_outputs(5304)) or (layer2_outputs(1105));
    layer3_outputs(4261) <= (layer2_outputs(875)) and not (layer2_outputs(2737));
    layer3_outputs(4262) <= not((layer2_outputs(5116)) or (layer2_outputs(5966)));
    layer3_outputs(4263) <= not(layer2_outputs(2583));
    layer3_outputs(4264) <= not(layer2_outputs(2288)) or (layer2_outputs(6537));
    layer3_outputs(4265) <= '1';
    layer3_outputs(4266) <= not(layer2_outputs(6814));
    layer3_outputs(4267) <= not(layer2_outputs(1694)) or (layer2_outputs(3389));
    layer3_outputs(4268) <= layer2_outputs(3901);
    layer3_outputs(4269) <= not(layer2_outputs(6276));
    layer3_outputs(4270) <= layer2_outputs(2748);
    layer3_outputs(4271) <= not(layer2_outputs(1314)) or (layer2_outputs(5005));
    layer3_outputs(4272) <= (layer2_outputs(7567)) or (layer2_outputs(4476));
    layer3_outputs(4273) <= not(layer2_outputs(5832));
    layer3_outputs(4274) <= (layer2_outputs(4855)) and (layer2_outputs(790));
    layer3_outputs(4275) <= not((layer2_outputs(5628)) or (layer2_outputs(7373)));
    layer3_outputs(4276) <= layer2_outputs(7109);
    layer3_outputs(4277) <= not(layer2_outputs(5493));
    layer3_outputs(4278) <= not((layer2_outputs(3346)) and (layer2_outputs(5702)));
    layer3_outputs(4279) <= not(layer2_outputs(885)) or (layer2_outputs(3496));
    layer3_outputs(4280) <= not(layer2_outputs(968)) or (layer2_outputs(5994));
    layer3_outputs(4281) <= not(layer2_outputs(5884));
    layer3_outputs(4282) <= (layer2_outputs(5618)) and not (layer2_outputs(3710));
    layer3_outputs(4283) <= not(layer2_outputs(5418));
    layer3_outputs(4284) <= (layer2_outputs(5944)) and not (layer2_outputs(915));
    layer3_outputs(4285) <= (layer2_outputs(4969)) and (layer2_outputs(3237));
    layer3_outputs(4286) <= (layer2_outputs(5535)) xor (layer2_outputs(6581));
    layer3_outputs(4287) <= (layer2_outputs(7231)) and (layer2_outputs(4565));
    layer3_outputs(4288) <= not(layer2_outputs(4486)) or (layer2_outputs(1898));
    layer3_outputs(4289) <= not(layer2_outputs(852));
    layer3_outputs(4290) <= '0';
    layer3_outputs(4291) <= not((layer2_outputs(7557)) xor (layer2_outputs(3473)));
    layer3_outputs(4292) <= not((layer2_outputs(888)) or (layer2_outputs(6060)));
    layer3_outputs(4293) <= (layer2_outputs(2816)) or (layer2_outputs(6117));
    layer3_outputs(4294) <= (layer2_outputs(6042)) or (layer2_outputs(6804));
    layer3_outputs(4295) <= layer2_outputs(1030);
    layer3_outputs(4296) <= not(layer2_outputs(2191));
    layer3_outputs(4297) <= not(layer2_outputs(4500));
    layer3_outputs(4298) <= not(layer2_outputs(1946));
    layer3_outputs(4299) <= not(layer2_outputs(5531));
    layer3_outputs(4300) <= layer2_outputs(6387);
    layer3_outputs(4301) <= (layer2_outputs(4127)) and not (layer2_outputs(7108));
    layer3_outputs(4302) <= not(layer2_outputs(657));
    layer3_outputs(4303) <= (layer2_outputs(4148)) and not (layer2_outputs(7268));
    layer3_outputs(4304) <= not(layer2_outputs(6887));
    layer3_outputs(4305) <= (layer2_outputs(4410)) and (layer2_outputs(6663));
    layer3_outputs(4306) <= not((layer2_outputs(6682)) xor (layer2_outputs(7600)));
    layer3_outputs(4307) <= layer2_outputs(109);
    layer3_outputs(4308) <= not(layer2_outputs(5356));
    layer3_outputs(4309) <= (layer2_outputs(5567)) and not (layer2_outputs(5710));
    layer3_outputs(4310) <= not((layer2_outputs(6650)) and (layer2_outputs(4026)));
    layer3_outputs(4311) <= not(layer2_outputs(3064));
    layer3_outputs(4312) <= '1';
    layer3_outputs(4313) <= (layer2_outputs(2928)) and (layer2_outputs(4352));
    layer3_outputs(4314) <= not(layer2_outputs(2307));
    layer3_outputs(4315) <= layer2_outputs(4703);
    layer3_outputs(4316) <= '1';
    layer3_outputs(4317) <= not(layer2_outputs(4864));
    layer3_outputs(4318) <= layer2_outputs(6194);
    layer3_outputs(4319) <= (layer2_outputs(1473)) and not (layer2_outputs(6221));
    layer3_outputs(4320) <= (layer2_outputs(1167)) and not (layer2_outputs(5596));
    layer3_outputs(4321) <= not(layer2_outputs(2047));
    layer3_outputs(4322) <= layer2_outputs(97);
    layer3_outputs(4323) <= layer2_outputs(4791);
    layer3_outputs(4324) <= (layer2_outputs(620)) and not (layer2_outputs(5605));
    layer3_outputs(4325) <= not(layer2_outputs(2714));
    layer3_outputs(4326) <= (layer2_outputs(3326)) and (layer2_outputs(5520));
    layer3_outputs(4327) <= layer2_outputs(6006);
    layer3_outputs(4328) <= (layer2_outputs(4617)) and not (layer2_outputs(5768));
    layer3_outputs(4329) <= not((layer2_outputs(3224)) xor (layer2_outputs(5903)));
    layer3_outputs(4330) <= not(layer2_outputs(6656));
    layer3_outputs(4331) <= layer2_outputs(6298);
    layer3_outputs(4332) <= not(layer2_outputs(4764));
    layer3_outputs(4333) <= (layer2_outputs(5006)) xor (layer2_outputs(6011));
    layer3_outputs(4334) <= (layer2_outputs(2647)) and (layer2_outputs(3874));
    layer3_outputs(4335) <= not(layer2_outputs(7247));
    layer3_outputs(4336) <= not(layer2_outputs(6385));
    layer3_outputs(4337) <= not(layer2_outputs(2130)) or (layer2_outputs(3338));
    layer3_outputs(4338) <= not(layer2_outputs(7043));
    layer3_outputs(4339) <= not((layer2_outputs(2569)) or (layer2_outputs(7006)));
    layer3_outputs(4340) <= not(layer2_outputs(2692));
    layer3_outputs(4341) <= not(layer2_outputs(2705)) or (layer2_outputs(2384));
    layer3_outputs(4342) <= (layer2_outputs(233)) or (layer2_outputs(929));
    layer3_outputs(4343) <= not((layer2_outputs(7331)) and (layer2_outputs(5570)));
    layer3_outputs(4344) <= not((layer2_outputs(1434)) and (layer2_outputs(5808)));
    layer3_outputs(4345) <= not(layer2_outputs(1512));
    layer3_outputs(4346) <= not(layer2_outputs(2649)) or (layer2_outputs(172));
    layer3_outputs(4347) <= not(layer2_outputs(3030));
    layer3_outputs(4348) <= not(layer2_outputs(3062));
    layer3_outputs(4349) <= (layer2_outputs(6207)) or (layer2_outputs(2302));
    layer3_outputs(4350) <= not((layer2_outputs(142)) and (layer2_outputs(3742)));
    layer3_outputs(4351) <= not(layer2_outputs(595)) or (layer2_outputs(7409));
    layer3_outputs(4352) <= not(layer2_outputs(4480));
    layer3_outputs(4353) <= not(layer2_outputs(1089)) or (layer2_outputs(3984));
    layer3_outputs(4354) <= not(layer2_outputs(1092));
    layer3_outputs(4355) <= not((layer2_outputs(788)) xor (layer2_outputs(6749)));
    layer3_outputs(4356) <= (layer2_outputs(2677)) and not (layer2_outputs(5573));
    layer3_outputs(4357) <= (layer2_outputs(1398)) or (layer2_outputs(2707));
    layer3_outputs(4358) <= not((layer2_outputs(7549)) and (layer2_outputs(2418)));
    layer3_outputs(4359) <= (layer2_outputs(3416)) xor (layer2_outputs(5484));
    layer3_outputs(4360) <= layer2_outputs(606);
    layer3_outputs(4361) <= layer2_outputs(5480);
    layer3_outputs(4362) <= (layer2_outputs(2137)) xor (layer2_outputs(4325));
    layer3_outputs(4363) <= layer2_outputs(4341);
    layer3_outputs(4364) <= not((layer2_outputs(4587)) or (layer2_outputs(6534)));
    layer3_outputs(4365) <= layer2_outputs(1389);
    layer3_outputs(4366) <= not((layer2_outputs(4430)) or (layer2_outputs(2383)));
    layer3_outputs(4367) <= not(layer2_outputs(4528));
    layer3_outputs(4368) <= not(layer2_outputs(2053));
    layer3_outputs(4369) <= (layer2_outputs(3743)) and not (layer2_outputs(4063));
    layer3_outputs(4370) <= layer2_outputs(7346);
    layer3_outputs(4371) <= layer2_outputs(6419);
    layer3_outputs(4372) <= layer2_outputs(4912);
    layer3_outputs(4373) <= (layer2_outputs(7003)) and not (layer2_outputs(2819));
    layer3_outputs(4374) <= not(layer2_outputs(7225));
    layer3_outputs(4375) <= layer2_outputs(7412);
    layer3_outputs(4376) <= not(layer2_outputs(4789)) or (layer2_outputs(7082));
    layer3_outputs(4377) <= '0';
    layer3_outputs(4378) <= layer2_outputs(4576);
    layer3_outputs(4379) <= (layer2_outputs(6904)) and not (layer2_outputs(4775));
    layer3_outputs(4380) <= not((layer2_outputs(2736)) or (layer2_outputs(6264)));
    layer3_outputs(4381) <= not(layer2_outputs(245));
    layer3_outputs(4382) <= (layer2_outputs(7035)) and (layer2_outputs(3833));
    layer3_outputs(4383) <= (layer2_outputs(1905)) and not (layer2_outputs(6553));
    layer3_outputs(4384) <= '0';
    layer3_outputs(4385) <= not(layer2_outputs(1630));
    layer3_outputs(4386) <= (layer2_outputs(1514)) and (layer2_outputs(6732));
    layer3_outputs(4387) <= not(layer2_outputs(249));
    layer3_outputs(4388) <= layer2_outputs(4367);
    layer3_outputs(4389) <= (layer2_outputs(3440)) or (layer2_outputs(6622));
    layer3_outputs(4390) <= '1';
    layer3_outputs(4391) <= not(layer2_outputs(6789));
    layer3_outputs(4392) <= not((layer2_outputs(6460)) and (layer2_outputs(965)));
    layer3_outputs(4393) <= layer2_outputs(6634);
    layer3_outputs(4394) <= (layer2_outputs(4447)) or (layer2_outputs(3038));
    layer3_outputs(4395) <= not(layer2_outputs(1780)) or (layer2_outputs(5301));
    layer3_outputs(4396) <= layer2_outputs(5411);
    layer3_outputs(4397) <= not(layer2_outputs(6133));
    layer3_outputs(4398) <= (layer2_outputs(4282)) or (layer2_outputs(3794));
    layer3_outputs(4399) <= (layer2_outputs(3732)) and not (layer2_outputs(6433));
    layer3_outputs(4400) <= '1';
    layer3_outputs(4401) <= not(layer2_outputs(3730));
    layer3_outputs(4402) <= layer2_outputs(5061);
    layer3_outputs(4403) <= layer2_outputs(1709);
    layer3_outputs(4404) <= layer2_outputs(297);
    layer3_outputs(4405) <= not(layer2_outputs(6319)) or (layer2_outputs(6107));
    layer3_outputs(4406) <= not(layer2_outputs(1328));
    layer3_outputs(4407) <= not((layer2_outputs(4396)) or (layer2_outputs(3820)));
    layer3_outputs(4408) <= not(layer2_outputs(6432));
    layer3_outputs(4409) <= (layer2_outputs(3016)) and not (layer2_outputs(2234));
    layer3_outputs(4410) <= layer2_outputs(6371);
    layer3_outputs(4411) <= (layer2_outputs(5090)) and (layer2_outputs(4214));
    layer3_outputs(4412) <= layer2_outputs(3432);
    layer3_outputs(4413) <= '1';
    layer3_outputs(4414) <= (layer2_outputs(849)) and not (layer2_outputs(6506));
    layer3_outputs(4415) <= not(layer2_outputs(5311));
    layer3_outputs(4416) <= not(layer2_outputs(1031)) or (layer2_outputs(5866));
    layer3_outputs(4417) <= not((layer2_outputs(1193)) or (layer2_outputs(6722)));
    layer3_outputs(4418) <= not(layer2_outputs(7062));
    layer3_outputs(4419) <= '1';
    layer3_outputs(4420) <= layer2_outputs(7376);
    layer3_outputs(4421) <= not(layer2_outputs(5406)) or (layer2_outputs(6116));
    layer3_outputs(4422) <= (layer2_outputs(4185)) and not (layer2_outputs(2651));
    layer3_outputs(4423) <= layer2_outputs(830);
    layer3_outputs(4424) <= not((layer2_outputs(4566)) xor (layer2_outputs(5732)));
    layer3_outputs(4425) <= (layer2_outputs(3065)) and (layer2_outputs(7432));
    layer3_outputs(4426) <= (layer2_outputs(6831)) and not (layer2_outputs(5536));
    layer3_outputs(4427) <= (layer2_outputs(7576)) and (layer2_outputs(7206));
    layer3_outputs(4428) <= (layer2_outputs(1256)) xor (layer2_outputs(5031));
    layer3_outputs(4429) <= not(layer2_outputs(629)) or (layer2_outputs(1662));
    layer3_outputs(4430) <= not(layer2_outputs(7596));
    layer3_outputs(4431) <= layer2_outputs(4342);
    layer3_outputs(4432) <= (layer2_outputs(5040)) or (layer2_outputs(1173));
    layer3_outputs(4433) <= (layer2_outputs(3400)) or (layer2_outputs(4178));
    layer3_outputs(4434) <= layer2_outputs(1874);
    layer3_outputs(4435) <= not((layer2_outputs(86)) or (layer2_outputs(4159)));
    layer3_outputs(4436) <= '0';
    layer3_outputs(4437) <= (layer2_outputs(6965)) and (layer2_outputs(5912));
    layer3_outputs(4438) <= layer2_outputs(3333);
    layer3_outputs(4439) <= not(layer2_outputs(1902));
    layer3_outputs(4440) <= layer2_outputs(6751);
    layer3_outputs(4441) <= (layer2_outputs(1576)) and (layer2_outputs(6179));
    layer3_outputs(4442) <= layer2_outputs(3159);
    layer3_outputs(4443) <= (layer2_outputs(3544)) and not (layer2_outputs(7000));
    layer3_outputs(4444) <= layer2_outputs(6890);
    layer3_outputs(4445) <= not(layer2_outputs(2700)) or (layer2_outputs(191));
    layer3_outputs(4446) <= (layer2_outputs(3097)) or (layer2_outputs(5815));
    layer3_outputs(4447) <= layer2_outputs(3724);
    layer3_outputs(4448) <= not((layer2_outputs(1025)) or (layer2_outputs(5952)));
    layer3_outputs(4449) <= (layer2_outputs(414)) xor (layer2_outputs(1781));
    layer3_outputs(4450) <= not(layer2_outputs(347)) or (layer2_outputs(6041));
    layer3_outputs(4451) <= '1';
    layer3_outputs(4452) <= layer2_outputs(5803);
    layer3_outputs(4453) <= layer2_outputs(6574);
    layer3_outputs(4454) <= not((layer2_outputs(4854)) and (layer2_outputs(2501)));
    layer3_outputs(4455) <= not(layer2_outputs(7431));
    layer3_outputs(4456) <= layer2_outputs(7335);
    layer3_outputs(4457) <= not(layer2_outputs(6892)) or (layer2_outputs(7288));
    layer3_outputs(4458) <= (layer2_outputs(7479)) and (layer2_outputs(3891));
    layer3_outputs(4459) <= not(layer2_outputs(7280)) or (layer2_outputs(630));
    layer3_outputs(4460) <= (layer2_outputs(4167)) and not (layer2_outputs(2119));
    layer3_outputs(4461) <= not(layer2_outputs(6955));
    layer3_outputs(4462) <= layer2_outputs(5466);
    layer3_outputs(4463) <= not(layer2_outputs(5099));
    layer3_outputs(4464) <= not(layer2_outputs(5355));
    layer3_outputs(4465) <= not(layer2_outputs(3183));
    layer3_outputs(4466) <= not((layer2_outputs(4317)) xor (layer2_outputs(2777)));
    layer3_outputs(4467) <= not(layer2_outputs(1496)) or (layer2_outputs(1785));
    layer3_outputs(4468) <= layer2_outputs(7236);
    layer3_outputs(4469) <= layer2_outputs(2961);
    layer3_outputs(4470) <= (layer2_outputs(4420)) and not (layer2_outputs(3487));
    layer3_outputs(4471) <= layer2_outputs(657);
    layer3_outputs(4472) <= not(layer2_outputs(1874));
    layer3_outputs(4473) <= not((layer2_outputs(4153)) and (layer2_outputs(1741)));
    layer3_outputs(4474) <= not(layer2_outputs(548)) or (layer2_outputs(7595));
    layer3_outputs(4475) <= (layer2_outputs(2234)) and (layer2_outputs(5880));
    layer3_outputs(4476) <= not((layer2_outputs(2900)) and (layer2_outputs(7652)));
    layer3_outputs(4477) <= (layer2_outputs(3134)) and not (layer2_outputs(2938));
    layer3_outputs(4478) <= not((layer2_outputs(1019)) or (layer2_outputs(1446)));
    layer3_outputs(4479) <= layer2_outputs(6615);
    layer3_outputs(4480) <= (layer2_outputs(1301)) xor (layer2_outputs(1756));
    layer3_outputs(4481) <= not(layer2_outputs(5580)) or (layer2_outputs(4474));
    layer3_outputs(4482) <= not(layer2_outputs(5186));
    layer3_outputs(4483) <= layer2_outputs(3037);
    layer3_outputs(4484) <= not(layer2_outputs(6227));
    layer3_outputs(4485) <= (layer2_outputs(5391)) and not (layer2_outputs(7300));
    layer3_outputs(4486) <= not(layer2_outputs(656)) or (layer2_outputs(1157));
    layer3_outputs(4487) <= '1';
    layer3_outputs(4488) <= not(layer2_outputs(1086));
    layer3_outputs(4489) <= layer2_outputs(2892);
    layer3_outputs(4490) <= (layer2_outputs(4480)) and not (layer2_outputs(2887));
    layer3_outputs(4491) <= not((layer2_outputs(860)) or (layer2_outputs(403)));
    layer3_outputs(4492) <= (layer2_outputs(5274)) or (layer2_outputs(3683));
    layer3_outputs(4493) <= not((layer2_outputs(7671)) and (layer2_outputs(5948)));
    layer3_outputs(4494) <= not((layer2_outputs(5981)) or (layer2_outputs(937)));
    layer3_outputs(4495) <= (layer2_outputs(6936)) and (layer2_outputs(4314));
    layer3_outputs(4496) <= layer2_outputs(5456);
    layer3_outputs(4497) <= (layer2_outputs(6127)) and (layer2_outputs(4463));
    layer3_outputs(4498) <= not((layer2_outputs(3196)) and (layer2_outputs(2056)));
    layer3_outputs(4499) <= not(layer2_outputs(6234));
    layer3_outputs(4500) <= not((layer2_outputs(7403)) and (layer2_outputs(1967)));
    layer3_outputs(4501) <= layer2_outputs(5793);
    layer3_outputs(4502) <= (layer2_outputs(4869)) and not (layer2_outputs(4865));
    layer3_outputs(4503) <= (layer2_outputs(5551)) or (layer2_outputs(131));
    layer3_outputs(4504) <= (layer2_outputs(7416)) and (layer2_outputs(1085));
    layer3_outputs(4505) <= not(layer2_outputs(510)) or (layer2_outputs(2098));
    layer3_outputs(4506) <= not(layer2_outputs(5801));
    layer3_outputs(4507) <= not((layer2_outputs(4879)) and (layer2_outputs(7432)));
    layer3_outputs(4508) <= (layer2_outputs(5146)) or (layer2_outputs(1100));
    layer3_outputs(4509) <= not(layer2_outputs(4334)) or (layer2_outputs(3913));
    layer3_outputs(4510) <= '1';
    layer3_outputs(4511) <= not(layer2_outputs(3783)) or (layer2_outputs(2695));
    layer3_outputs(4512) <= layer2_outputs(2184);
    layer3_outputs(4513) <= (layer2_outputs(5016)) and not (layer2_outputs(6774));
    layer3_outputs(4514) <= not(layer2_outputs(1713)) or (layer2_outputs(1764));
    layer3_outputs(4515) <= '1';
    layer3_outputs(4516) <= not(layer2_outputs(3309));
    layer3_outputs(4517) <= (layer2_outputs(473)) and not (layer2_outputs(327));
    layer3_outputs(4518) <= not((layer2_outputs(2467)) or (layer2_outputs(5126)));
    layer3_outputs(4519) <= not((layer2_outputs(1445)) xor (layer2_outputs(2023)));
    layer3_outputs(4520) <= not(layer2_outputs(4451)) or (layer2_outputs(4454));
    layer3_outputs(4521) <= (layer2_outputs(4833)) and not (layer2_outputs(2113));
    layer3_outputs(4522) <= not(layer2_outputs(2625));
    layer3_outputs(4523) <= layer2_outputs(820);
    layer3_outputs(4524) <= not(layer2_outputs(4759));
    layer3_outputs(4525) <= layer2_outputs(7017);
    layer3_outputs(4526) <= not(layer2_outputs(7653));
    layer3_outputs(4527) <= (layer2_outputs(767)) and not (layer2_outputs(5925));
    layer3_outputs(4528) <= not((layer2_outputs(7029)) and (layer2_outputs(4270)));
    layer3_outputs(4529) <= not(layer2_outputs(1299));
    layer3_outputs(4530) <= not(layer2_outputs(3363));
    layer3_outputs(4531) <= layer2_outputs(961);
    layer3_outputs(4532) <= layer2_outputs(2163);
    layer3_outputs(4533) <= (layer2_outputs(6791)) and not (layer2_outputs(7137));
    layer3_outputs(4534) <= not((layer2_outputs(681)) or (layer2_outputs(1897)));
    layer3_outputs(4535) <= not(layer2_outputs(75));
    layer3_outputs(4536) <= not(layer2_outputs(4509));
    layer3_outputs(4537) <= not(layer2_outputs(3154));
    layer3_outputs(4538) <= (layer2_outputs(814)) xor (layer2_outputs(7058));
    layer3_outputs(4539) <= layer2_outputs(5590);
    layer3_outputs(4540) <= not(layer2_outputs(240));
    layer3_outputs(4541) <= (layer2_outputs(454)) and not (layer2_outputs(3350));
    layer3_outputs(4542) <= layer2_outputs(7170);
    layer3_outputs(4543) <= not(layer2_outputs(516)) or (layer2_outputs(1529));
    layer3_outputs(4544) <= not(layer2_outputs(949));
    layer3_outputs(4545) <= (layer2_outputs(539)) and not (layer2_outputs(5446));
    layer3_outputs(4546) <= (layer2_outputs(3254)) and (layer2_outputs(1638));
    layer3_outputs(4547) <= layer2_outputs(6221);
    layer3_outputs(4548) <= not(layer2_outputs(1423));
    layer3_outputs(4549) <= not(layer2_outputs(4411));
    layer3_outputs(4550) <= (layer2_outputs(5543)) and not (layer2_outputs(6841));
    layer3_outputs(4551) <= layer2_outputs(7389);
    layer3_outputs(4552) <= layer2_outputs(2860);
    layer3_outputs(4553) <= not(layer2_outputs(5652)) or (layer2_outputs(5937));
    layer3_outputs(4554) <= (layer2_outputs(1439)) and (layer2_outputs(4224));
    layer3_outputs(4555) <= not((layer2_outputs(17)) or (layer2_outputs(3342)));
    layer3_outputs(4556) <= not((layer2_outputs(2026)) or (layer2_outputs(3205)));
    layer3_outputs(4557) <= layer2_outputs(880);
    layer3_outputs(4558) <= not(layer2_outputs(236));
    layer3_outputs(4559) <= not(layer2_outputs(4348)) or (layer2_outputs(5074));
    layer3_outputs(4560) <= not(layer2_outputs(552));
    layer3_outputs(4561) <= not(layer2_outputs(4404));
    layer3_outputs(4562) <= (layer2_outputs(2802)) or (layer2_outputs(7673));
    layer3_outputs(4563) <= (layer2_outputs(3469)) and (layer2_outputs(3552));
    layer3_outputs(4564) <= layer2_outputs(6549);
    layer3_outputs(4565) <= not((layer2_outputs(7194)) and (layer2_outputs(5126)));
    layer3_outputs(4566) <= not(layer2_outputs(5546));
    layer3_outputs(4567) <= not(layer2_outputs(2624));
    layer3_outputs(4568) <= layer2_outputs(6836);
    layer3_outputs(4569) <= not(layer2_outputs(2742));
    layer3_outputs(4570) <= not(layer2_outputs(708)) or (layer2_outputs(2257));
    layer3_outputs(4571) <= not(layer2_outputs(2202));
    layer3_outputs(4572) <= not(layer2_outputs(2727));
    layer3_outputs(4573) <= not(layer2_outputs(3887));
    layer3_outputs(4574) <= (layer2_outputs(4483)) and not (layer2_outputs(2644));
    layer3_outputs(4575) <= (layer2_outputs(5833)) and not (layer2_outputs(7578));
    layer3_outputs(4576) <= layer2_outputs(5868);
    layer3_outputs(4577) <= layer2_outputs(2407);
    layer3_outputs(4578) <= '0';
    layer3_outputs(4579) <= not((layer2_outputs(5683)) or (layer2_outputs(6720)));
    layer3_outputs(4580) <= not(layer2_outputs(3371)) or (layer2_outputs(939));
    layer3_outputs(4581) <= layer2_outputs(69);
    layer3_outputs(4582) <= (layer2_outputs(2879)) and (layer2_outputs(6712));
    layer3_outputs(4583) <= not((layer2_outputs(1631)) and (layer2_outputs(3983)));
    layer3_outputs(4584) <= not(layer2_outputs(53));
    layer3_outputs(4585) <= not(layer2_outputs(4055)) or (layer2_outputs(2196));
    layer3_outputs(4586) <= not((layer2_outputs(509)) or (layer2_outputs(2180)));
    layer3_outputs(4587) <= (layer2_outputs(5453)) and not (layer2_outputs(1433));
    layer3_outputs(4588) <= not((layer2_outputs(3636)) and (layer2_outputs(7196)));
    layer3_outputs(4589) <= (layer2_outputs(5415)) and not (layer2_outputs(7028));
    layer3_outputs(4590) <= not(layer2_outputs(7385));
    layer3_outputs(4591) <= not(layer2_outputs(6396)) or (layer2_outputs(2838));
    layer3_outputs(4592) <= (layer2_outputs(3655)) and not (layer2_outputs(2972));
    layer3_outputs(4593) <= not((layer2_outputs(967)) or (layer2_outputs(4484)));
    layer3_outputs(4594) <= (layer2_outputs(23)) or (layer2_outputs(5337));
    layer3_outputs(4595) <= (layer2_outputs(861)) and not (layer2_outputs(4541));
    layer3_outputs(4596) <= not(layer2_outputs(5580)) or (layer2_outputs(7016));
    layer3_outputs(4597) <= layer2_outputs(5332);
    layer3_outputs(4598) <= layer2_outputs(3240);
    layer3_outputs(4599) <= layer2_outputs(4435);
    layer3_outputs(4600) <= layer2_outputs(4005);
    layer3_outputs(4601) <= not((layer2_outputs(1205)) or (layer2_outputs(5770)));
    layer3_outputs(4602) <= not(layer2_outputs(2463));
    layer3_outputs(4603) <= not(layer2_outputs(4025)) or (layer2_outputs(6098));
    layer3_outputs(4604) <= not(layer2_outputs(4844));
    layer3_outputs(4605) <= (layer2_outputs(5524)) and (layer2_outputs(71));
    layer3_outputs(4606) <= (layer2_outputs(3679)) xor (layer2_outputs(6895));
    layer3_outputs(4607) <= layer2_outputs(1004);
    layer3_outputs(4608) <= not((layer2_outputs(6244)) or (layer2_outputs(2940)));
    layer3_outputs(4609) <= layer2_outputs(7127);
    layer3_outputs(4610) <= not(layer2_outputs(2967));
    layer3_outputs(4611) <= (layer2_outputs(857)) and not (layer2_outputs(4545));
    layer3_outputs(4612) <= not(layer2_outputs(3147)) or (layer2_outputs(4676));
    layer3_outputs(4613) <= layer2_outputs(866);
    layer3_outputs(4614) <= (layer2_outputs(5341)) and not (layer2_outputs(4406));
    layer3_outputs(4615) <= not(layer2_outputs(7583));
    layer3_outputs(4616) <= layer2_outputs(6235);
    layer3_outputs(4617) <= layer2_outputs(1371);
    layer3_outputs(4618) <= not(layer2_outputs(6658));
    layer3_outputs(4619) <= not((layer2_outputs(6152)) and (layer2_outputs(2825)));
    layer3_outputs(4620) <= not(layer2_outputs(6721));
    layer3_outputs(4621) <= (layer2_outputs(6981)) and not (layer2_outputs(2399));
    layer3_outputs(4622) <= layer2_outputs(368);
    layer3_outputs(4623) <= not(layer2_outputs(1988));
    layer3_outputs(4624) <= not(layer2_outputs(5881));
    layer3_outputs(4625) <= not((layer2_outputs(5101)) and (layer2_outputs(3246)));
    layer3_outputs(4626) <= layer2_outputs(3617);
    layer3_outputs(4627) <= not(layer2_outputs(5637));
    layer3_outputs(4628) <= layer2_outputs(7171);
    layer3_outputs(4629) <= not(layer2_outputs(1127)) or (layer2_outputs(2330));
    layer3_outputs(4630) <= not(layer2_outputs(6022)) or (layer2_outputs(4046));
    layer3_outputs(4631) <= not(layer2_outputs(6329));
    layer3_outputs(4632) <= layer2_outputs(3600);
    layer3_outputs(4633) <= not(layer2_outputs(2833));
    layer3_outputs(4634) <= not((layer2_outputs(5142)) or (layer2_outputs(5990)));
    layer3_outputs(4635) <= layer2_outputs(3685);
    layer3_outputs(4636) <= layer2_outputs(2355);
    layer3_outputs(4637) <= (layer2_outputs(6747)) xor (layer2_outputs(940));
    layer3_outputs(4638) <= layer2_outputs(1622);
    layer3_outputs(4639) <= not(layer2_outputs(2298));
    layer3_outputs(4640) <= not(layer2_outputs(761)) or (layer2_outputs(4561));
    layer3_outputs(4641) <= not(layer2_outputs(7051));
    layer3_outputs(4642) <= layer2_outputs(3133);
    layer3_outputs(4643) <= not(layer2_outputs(7477)) or (layer2_outputs(523));
    layer3_outputs(4644) <= not(layer2_outputs(7501));
    layer3_outputs(4645) <= (layer2_outputs(2317)) and not (layer2_outputs(3061));
    layer3_outputs(4646) <= not(layer2_outputs(6566));
    layer3_outputs(4647) <= layer2_outputs(6642);
    layer3_outputs(4648) <= not(layer2_outputs(4098));
    layer3_outputs(4649) <= layer2_outputs(7558);
    layer3_outputs(4650) <= not((layer2_outputs(1966)) or (layer2_outputs(6817)));
    layer3_outputs(4651) <= not(layer2_outputs(390)) or (layer2_outputs(2444));
    layer3_outputs(4652) <= layer2_outputs(3652);
    layer3_outputs(4653) <= not((layer2_outputs(1866)) and (layer2_outputs(3064)));
    layer3_outputs(4654) <= not(layer2_outputs(1542));
    layer3_outputs(4655) <= not(layer2_outputs(4222)) or (layer2_outputs(5983));
    layer3_outputs(4656) <= layer2_outputs(4239);
    layer3_outputs(4657) <= not(layer2_outputs(3070));
    layer3_outputs(4658) <= not(layer2_outputs(7504)) or (layer2_outputs(7644));
    layer3_outputs(4659) <= (layer2_outputs(5039)) or (layer2_outputs(2530));
    layer3_outputs(4660) <= not(layer2_outputs(5658)) or (layer2_outputs(4761));
    layer3_outputs(4661) <= not(layer2_outputs(7627));
    layer3_outputs(4662) <= not(layer2_outputs(4971));
    layer3_outputs(4663) <= (layer2_outputs(1545)) and not (layer2_outputs(1177));
    layer3_outputs(4664) <= not(layer2_outputs(4975));
    layer3_outputs(4665) <= not(layer2_outputs(3269));
    layer3_outputs(4666) <= (layer2_outputs(3629)) and (layer2_outputs(1091));
    layer3_outputs(4667) <= not(layer2_outputs(1091));
    layer3_outputs(4668) <= layer2_outputs(1719);
    layer3_outputs(4669) <= layer2_outputs(2937);
    layer3_outputs(4670) <= layer2_outputs(5854);
    layer3_outputs(4671) <= not((layer2_outputs(3122)) or (layer2_outputs(6266)));
    layer3_outputs(4672) <= (layer2_outputs(6978)) and (layer2_outputs(556));
    layer3_outputs(4673) <= not(layer2_outputs(4386));
    layer3_outputs(4674) <= not(layer2_outputs(2990)) or (layer2_outputs(3019));
    layer3_outputs(4675) <= not((layer2_outputs(4888)) and (layer2_outputs(667)));
    layer3_outputs(4676) <= (layer2_outputs(5308)) and not (layer2_outputs(898));
    layer3_outputs(4677) <= layer2_outputs(3622);
    layer3_outputs(4678) <= layer2_outputs(3957);
    layer3_outputs(4679) <= not(layer2_outputs(3171));
    layer3_outputs(4680) <= not(layer2_outputs(585)) or (layer2_outputs(2955));
    layer3_outputs(4681) <= (layer2_outputs(2352)) and not (layer2_outputs(6280));
    layer3_outputs(4682) <= not((layer2_outputs(261)) or (layer2_outputs(6443)));
    layer3_outputs(4683) <= not((layer2_outputs(4951)) or (layer2_outputs(714)));
    layer3_outputs(4684) <= not(layer2_outputs(4985)) or (layer2_outputs(134));
    layer3_outputs(4685) <= (layer2_outputs(2401)) and not (layer2_outputs(2367));
    layer3_outputs(4686) <= layer2_outputs(6516);
    layer3_outputs(4687) <= not(layer2_outputs(4385)) or (layer2_outputs(2869));
    layer3_outputs(4688) <= not(layer2_outputs(4027));
    layer3_outputs(4689) <= not(layer2_outputs(79));
    layer3_outputs(4690) <= layer2_outputs(1722);
    layer3_outputs(4691) <= not(layer2_outputs(4803)) or (layer2_outputs(177));
    layer3_outputs(4692) <= not(layer2_outputs(6833));
    layer3_outputs(4693) <= not(layer2_outputs(2338));
    layer3_outputs(4694) <= not(layer2_outputs(4238));
    layer3_outputs(4695) <= not((layer2_outputs(2381)) and (layer2_outputs(7469)));
    layer3_outputs(4696) <= not(layer2_outputs(461)) or (layer2_outputs(6158));
    layer3_outputs(4697) <= not(layer2_outputs(1538));
    layer3_outputs(4698) <= '0';
    layer3_outputs(4699) <= layer2_outputs(5372);
    layer3_outputs(4700) <= layer2_outputs(3723);
    layer3_outputs(4701) <= not((layer2_outputs(4306)) xor (layer2_outputs(2872)));
    layer3_outputs(4702) <= not(layer2_outputs(542)) or (layer2_outputs(7657));
    layer3_outputs(4703) <= layer2_outputs(7626);
    layer3_outputs(4704) <= layer2_outputs(952);
    layer3_outputs(4705) <= (layer2_outputs(6321)) and (layer2_outputs(5219));
    layer3_outputs(4706) <= (layer2_outputs(7283)) and not (layer2_outputs(1991));
    layer3_outputs(4707) <= (layer2_outputs(132)) and not (layer2_outputs(3459));
    layer3_outputs(4708) <= not(layer2_outputs(3455));
    layer3_outputs(4709) <= not(layer2_outputs(5405)) or (layer2_outputs(2915));
    layer3_outputs(4710) <= not((layer2_outputs(7176)) or (layer2_outputs(6405)));
    layer3_outputs(4711) <= layer2_outputs(406);
    layer3_outputs(4712) <= (layer2_outputs(4293)) and not (layer2_outputs(4008));
    layer3_outputs(4713) <= layer2_outputs(2443);
    layer3_outputs(4714) <= '0';
    layer3_outputs(4715) <= (layer2_outputs(497)) or (layer2_outputs(6676));
    layer3_outputs(4716) <= not(layer2_outputs(3377));
    layer3_outputs(4717) <= not(layer2_outputs(699));
    layer3_outputs(4718) <= layer2_outputs(2832);
    layer3_outputs(4719) <= not(layer2_outputs(864));
    layer3_outputs(4720) <= (layer2_outputs(1081)) and not (layer2_outputs(2902));
    layer3_outputs(4721) <= layer2_outputs(5518);
    layer3_outputs(4722) <= not((layer2_outputs(7461)) or (layer2_outputs(7149)));
    layer3_outputs(4723) <= (layer2_outputs(6591)) and not (layer2_outputs(1509));
    layer3_outputs(4724) <= not((layer2_outputs(3160)) xor (layer2_outputs(324)));
    layer3_outputs(4725) <= '0';
    layer3_outputs(4726) <= not((layer2_outputs(4867)) and (layer2_outputs(5870)));
    layer3_outputs(4727) <= not(layer2_outputs(854)) or (layer2_outputs(2876));
    layer3_outputs(4728) <= (layer2_outputs(1577)) or (layer2_outputs(4114));
    layer3_outputs(4729) <= (layer2_outputs(6398)) and (layer2_outputs(5350));
    layer3_outputs(4730) <= (layer2_outputs(2453)) and (layer2_outputs(4740));
    layer3_outputs(4731) <= layer2_outputs(5838);
    layer3_outputs(4732) <= not(layer2_outputs(6688));
    layer3_outputs(4733) <= (layer2_outputs(6111)) and not (layer2_outputs(6072));
    layer3_outputs(4734) <= not(layer2_outputs(55));
    layer3_outputs(4735) <= (layer2_outputs(1379)) or (layer2_outputs(6913));
    layer3_outputs(4736) <= layer2_outputs(6796);
    layer3_outputs(4737) <= '0';
    layer3_outputs(4738) <= layer2_outputs(2295);
    layer3_outputs(4739) <= (layer2_outputs(882)) xor (layer2_outputs(5950));
    layer3_outputs(4740) <= layer2_outputs(955);
    layer3_outputs(4741) <= layer2_outputs(6325);
    layer3_outputs(4742) <= (layer2_outputs(6463)) xor (layer2_outputs(4350));
    layer3_outputs(4743) <= not(layer2_outputs(3439));
    layer3_outputs(4744) <= not(layer2_outputs(7111)) or (layer2_outputs(3923));
    layer3_outputs(4745) <= not(layer2_outputs(1986)) or (layer2_outputs(163));
    layer3_outputs(4746) <= layer2_outputs(1562);
    layer3_outputs(4747) <= not(layer2_outputs(1997));
    layer3_outputs(4748) <= not(layer2_outputs(7290)) or (layer2_outputs(5169));
    layer3_outputs(4749) <= not((layer2_outputs(7129)) xor (layer2_outputs(2335)));
    layer3_outputs(4750) <= '0';
    layer3_outputs(4751) <= layer2_outputs(1239);
    layer3_outputs(4752) <= not(layer2_outputs(7073));
    layer3_outputs(4753) <= layer2_outputs(2300);
    layer3_outputs(4754) <= (layer2_outputs(2210)) and not (layer2_outputs(4127));
    layer3_outputs(4755) <= (layer2_outputs(1106)) or (layer2_outputs(2479));
    layer3_outputs(4756) <= layer2_outputs(759);
    layer3_outputs(4757) <= layer2_outputs(4622);
    layer3_outputs(4758) <= layer2_outputs(3771);
    layer3_outputs(4759) <= not(layer2_outputs(7491));
    layer3_outputs(4760) <= not(layer2_outputs(4535));
    layer3_outputs(4761) <= (layer2_outputs(2102)) or (layer2_outputs(2381));
    layer3_outputs(4762) <= '0';
    layer3_outputs(4763) <= not((layer2_outputs(3273)) xor (layer2_outputs(5932)));
    layer3_outputs(4764) <= not(layer2_outputs(890)) or (layer2_outputs(2512));
    layer3_outputs(4765) <= not((layer2_outputs(6421)) or (layer2_outputs(6568)));
    layer3_outputs(4766) <= layer2_outputs(4824);
    layer3_outputs(4767) <= not(layer2_outputs(6053));
    layer3_outputs(4768) <= not(layer2_outputs(1378)) or (layer2_outputs(5812));
    layer3_outputs(4769) <= (layer2_outputs(6865)) and not (layer2_outputs(7355));
    layer3_outputs(4770) <= layer2_outputs(1103);
    layer3_outputs(4771) <= not(layer2_outputs(6928)) or (layer2_outputs(1837));
    layer3_outputs(4772) <= layer2_outputs(2527);
    layer3_outputs(4773) <= not((layer2_outputs(4661)) or (layer2_outputs(3696)));
    layer3_outputs(4774) <= (layer2_outputs(3594)) or (layer2_outputs(609));
    layer3_outputs(4775) <= '1';
    layer3_outputs(4776) <= not(layer2_outputs(991)) or (layer2_outputs(755));
    layer3_outputs(4777) <= not(layer2_outputs(6985));
    layer3_outputs(4778) <= layer2_outputs(329);
    layer3_outputs(4779) <= (layer2_outputs(1228)) and (layer2_outputs(785));
    layer3_outputs(4780) <= layer2_outputs(1867);
    layer3_outputs(4781) <= not((layer2_outputs(2683)) xor (layer2_outputs(3067)));
    layer3_outputs(4782) <= (layer2_outputs(6108)) xor (layer2_outputs(5178));
    layer3_outputs(4783) <= not(layer2_outputs(3503));
    layer3_outputs(4784) <= not(layer2_outputs(3857));
    layer3_outputs(4785) <= not(layer2_outputs(5053));
    layer3_outputs(4786) <= not((layer2_outputs(528)) or (layer2_outputs(2203)));
    layer3_outputs(4787) <= (layer2_outputs(4388)) and not (layer2_outputs(5395));
    layer3_outputs(4788) <= not(layer2_outputs(2760));
    layer3_outputs(4789) <= layer2_outputs(4078);
    layer3_outputs(4790) <= not((layer2_outputs(1326)) and (layer2_outputs(5037)));
    layer3_outputs(4791) <= (layer2_outputs(5616)) and (layer2_outputs(7241));
    layer3_outputs(4792) <= not(layer2_outputs(4985)) or (layer2_outputs(4115));
    layer3_outputs(4793) <= not(layer2_outputs(7608)) or (layer2_outputs(7271));
    layer3_outputs(4794) <= not(layer2_outputs(1083));
    layer3_outputs(4795) <= not(layer2_outputs(46));
    layer3_outputs(4796) <= not(layer2_outputs(2122));
    layer3_outputs(4797) <= not(layer2_outputs(6503)) or (layer2_outputs(6928));
    layer3_outputs(4798) <= (layer2_outputs(2574)) and not (layer2_outputs(6320));
    layer3_outputs(4799) <= layer2_outputs(7330);
    layer3_outputs(4800) <= not(layer2_outputs(1691));
    layer3_outputs(4801) <= layer2_outputs(5350);
    layer3_outputs(4802) <= not(layer2_outputs(4870));
    layer3_outputs(4803) <= not((layer2_outputs(2928)) or (layer2_outputs(5195)));
    layer3_outputs(4804) <= not(layer2_outputs(3175));
    layer3_outputs(4805) <= (layer2_outputs(6091)) or (layer2_outputs(480));
    layer3_outputs(4806) <= not(layer2_outputs(7138));
    layer3_outputs(4807) <= (layer2_outputs(842)) and (layer2_outputs(2848));
    layer3_outputs(4808) <= not(layer2_outputs(2311)) or (layer2_outputs(80));
    layer3_outputs(4809) <= (layer2_outputs(4109)) and (layer2_outputs(1310));
    layer3_outputs(4810) <= (layer2_outputs(5419)) xor (layer2_outputs(2726));
    layer3_outputs(4811) <= not(layer2_outputs(6578)) or (layer2_outputs(1745));
    layer3_outputs(4812) <= not(layer2_outputs(682));
    layer3_outputs(4813) <= not(layer2_outputs(6702)) or (layer2_outputs(1956));
    layer3_outputs(4814) <= layer2_outputs(949);
    layer3_outputs(4815) <= (layer2_outputs(4263)) and (layer2_outputs(6238));
    layer3_outputs(4816) <= not(layer2_outputs(375)) or (layer2_outputs(5974));
    layer3_outputs(4817) <= '0';
    layer3_outputs(4818) <= not(layer2_outputs(5242));
    layer3_outputs(4819) <= layer2_outputs(720);
    layer3_outputs(4820) <= (layer2_outputs(6831)) and not (layer2_outputs(3425));
    layer3_outputs(4821) <= layer2_outputs(3828);
    layer3_outputs(4822) <= not((layer2_outputs(3116)) and (layer2_outputs(283)));
    layer3_outputs(4823) <= layer2_outputs(7036);
    layer3_outputs(4824) <= not(layer2_outputs(747));
    layer3_outputs(4825) <= not(layer2_outputs(2790)) or (layer2_outputs(7238));
    layer3_outputs(4826) <= layer2_outputs(1679);
    layer3_outputs(4827) <= layer2_outputs(4016);
    layer3_outputs(4828) <= (layer2_outputs(1248)) and not (layer2_outputs(4784));
    layer3_outputs(4829) <= not(layer2_outputs(6331));
    layer3_outputs(4830) <= not((layer2_outputs(1269)) xor (layer2_outputs(7032)));
    layer3_outputs(4831) <= (layer2_outputs(5883)) xor (layer2_outputs(7678));
    layer3_outputs(4832) <= layer2_outputs(5868);
    layer3_outputs(4833) <= layer2_outputs(1353);
    layer3_outputs(4834) <= not(layer2_outputs(1532)) or (layer2_outputs(1042));
    layer3_outputs(4835) <= not((layer2_outputs(6889)) and (layer2_outputs(6835)));
    layer3_outputs(4836) <= (layer2_outputs(4946)) and not (layer2_outputs(956));
    layer3_outputs(4837) <= '0';
    layer3_outputs(4838) <= (layer2_outputs(1338)) or (layer2_outputs(80));
    layer3_outputs(4839) <= not(layer2_outputs(3677));
    layer3_outputs(4840) <= '0';
    layer3_outputs(4841) <= not((layer2_outputs(4576)) and (layer2_outputs(712)));
    layer3_outputs(4842) <= not(layer2_outputs(1174)) or (layer2_outputs(146));
    layer3_outputs(4843) <= not(layer2_outputs(1314)) or (layer2_outputs(5897));
    layer3_outputs(4844) <= layer2_outputs(2934);
    layer3_outputs(4845) <= layer2_outputs(6313);
    layer3_outputs(4846) <= not(layer2_outputs(7271));
    layer3_outputs(4847) <= not(layer2_outputs(6555)) or (layer2_outputs(3502));
    layer3_outputs(4848) <= (layer2_outputs(3829)) and (layer2_outputs(5457));
    layer3_outputs(4849) <= (layer2_outputs(1188)) xor (layer2_outputs(3650));
    layer3_outputs(4850) <= layer2_outputs(4568);
    layer3_outputs(4851) <= '1';
    layer3_outputs(4852) <= not(layer2_outputs(2385));
    layer3_outputs(4853) <= (layer2_outputs(896)) xor (layer2_outputs(1805));
    layer3_outputs(4854) <= not(layer2_outputs(4894));
    layer3_outputs(4855) <= not(layer2_outputs(4309));
    layer3_outputs(4856) <= layer2_outputs(3628);
    layer3_outputs(4857) <= not((layer2_outputs(7630)) xor (layer2_outputs(4200)));
    layer3_outputs(4858) <= layer2_outputs(6140);
    layer3_outputs(4859) <= (layer2_outputs(2709)) and not (layer2_outputs(3692));
    layer3_outputs(4860) <= not(layer2_outputs(1015));
    layer3_outputs(4861) <= layer2_outputs(4997);
    layer3_outputs(4862) <= not(layer2_outputs(1619));
    layer3_outputs(4863) <= layer2_outputs(1260);
    layer3_outputs(4864) <= (layer2_outputs(692)) and (layer2_outputs(879));
    layer3_outputs(4865) <= layer2_outputs(4095);
    layer3_outputs(4866) <= (layer2_outputs(7028)) or (layer2_outputs(1604));
    layer3_outputs(4867) <= not(layer2_outputs(3429));
    layer3_outputs(4868) <= (layer2_outputs(5259)) and (layer2_outputs(4802));
    layer3_outputs(4869) <= not((layer2_outputs(7609)) xor (layer2_outputs(4943)));
    layer3_outputs(4870) <= layer2_outputs(3292);
    layer3_outputs(4871) <= (layer2_outputs(3711)) xor (layer2_outputs(458));
    layer3_outputs(4872) <= (layer2_outputs(2582)) and not (layer2_outputs(5383));
    layer3_outputs(4873) <= (layer2_outputs(7581)) and not (layer2_outputs(195));
    layer3_outputs(4874) <= (layer2_outputs(7415)) and not (layer2_outputs(3997));
    layer3_outputs(4875) <= '1';
    layer3_outputs(4876) <= not(layer2_outputs(3491));
    layer3_outputs(4877) <= not(layer2_outputs(7350));
    layer3_outputs(4878) <= not(layer2_outputs(1611));
    layer3_outputs(4879) <= not(layer2_outputs(4884));
    layer3_outputs(4880) <= not(layer2_outputs(3760));
    layer3_outputs(4881) <= not((layer2_outputs(2628)) or (layer2_outputs(6669)));
    layer3_outputs(4882) <= (layer2_outputs(3746)) or (layer2_outputs(495));
    layer3_outputs(4883) <= not(layer2_outputs(2779));
    layer3_outputs(4884) <= (layer2_outputs(5610)) or (layer2_outputs(2343));
    layer3_outputs(4885) <= not(layer2_outputs(3991)) or (layer2_outputs(6386));
    layer3_outputs(4886) <= not((layer2_outputs(2436)) or (layer2_outputs(4872)));
    layer3_outputs(4887) <= layer2_outputs(5445);
    layer3_outputs(4888) <= layer2_outputs(1945);
    layer3_outputs(4889) <= not(layer2_outputs(232));
    layer3_outputs(4890) <= (layer2_outputs(2859)) and not (layer2_outputs(7403));
    layer3_outputs(4891) <= layer2_outputs(839);
    layer3_outputs(4892) <= layer2_outputs(6760);
    layer3_outputs(4893) <= '0';
    layer3_outputs(4894) <= not((layer2_outputs(666)) or (layer2_outputs(7178)));
    layer3_outputs(4895) <= not(layer2_outputs(4768));
    layer3_outputs(4896) <= not(layer2_outputs(5291));
    layer3_outputs(4897) <= (layer2_outputs(5853)) or (layer2_outputs(1117));
    layer3_outputs(4898) <= '1';
    layer3_outputs(4899) <= not(layer2_outputs(4378));
    layer3_outputs(4900) <= '1';
    layer3_outputs(4901) <= not(layer2_outputs(4132));
    layer3_outputs(4902) <= layer2_outputs(4123);
    layer3_outputs(4903) <= (layer2_outputs(496)) and not (layer2_outputs(6621));
    layer3_outputs(4904) <= not(layer2_outputs(3344));
    layer3_outputs(4905) <= (layer2_outputs(2052)) and not (layer2_outputs(3198));
    layer3_outputs(4906) <= (layer2_outputs(5434)) and not (layer2_outputs(695));
    layer3_outputs(4907) <= layer2_outputs(4324);
    layer3_outputs(4908) <= (layer2_outputs(6684)) and not (layer2_outputs(362));
    layer3_outputs(4909) <= not(layer2_outputs(4957));
    layer3_outputs(4910) <= '0';
    layer3_outputs(4911) <= (layer2_outputs(3541)) and not (layer2_outputs(4396));
    layer3_outputs(4912) <= (layer2_outputs(4226)) and (layer2_outputs(1628));
    layer3_outputs(4913) <= not(layer2_outputs(5615));
    layer3_outputs(4914) <= (layer2_outputs(696)) or (layer2_outputs(2501));
    layer3_outputs(4915) <= layer2_outputs(6940);
    layer3_outputs(4916) <= layer2_outputs(7098);
    layer3_outputs(4917) <= (layer2_outputs(4781)) and not (layer2_outputs(7619));
    layer3_outputs(4918) <= not(layer2_outputs(4440));
    layer3_outputs(4919) <= (layer2_outputs(2902)) or (layer2_outputs(5045));
    layer3_outputs(4920) <= '1';
    layer3_outputs(4921) <= layer2_outputs(2919);
    layer3_outputs(4922) <= layer2_outputs(6859);
    layer3_outputs(4923) <= not(layer2_outputs(3053));
    layer3_outputs(4924) <= layer2_outputs(3113);
    layer3_outputs(4925) <= (layer2_outputs(4039)) xor (layer2_outputs(2351));
    layer3_outputs(4926) <= not((layer2_outputs(5046)) xor (layer2_outputs(4996)));
    layer3_outputs(4927) <= layer2_outputs(2973);
    layer3_outputs(4928) <= not((layer2_outputs(3780)) and (layer2_outputs(3980)));
    layer3_outputs(4929) <= not(layer2_outputs(1880)) or (layer2_outputs(6607));
    layer3_outputs(4930) <= layer2_outputs(1799);
    layer3_outputs(4931) <= '0';
    layer3_outputs(4932) <= layer2_outputs(5680);
    layer3_outputs(4933) <= layer2_outputs(6316);
    layer3_outputs(4934) <= layer2_outputs(1211);
    layer3_outputs(4935) <= not((layer2_outputs(6092)) or (layer2_outputs(496)));
    layer3_outputs(4936) <= not((layer2_outputs(6860)) or (layer2_outputs(3168)));
    layer3_outputs(4937) <= not((layer2_outputs(588)) or (layer2_outputs(646)));
    layer3_outputs(4938) <= not((layer2_outputs(5040)) and (layer2_outputs(5301)));
    layer3_outputs(4939) <= not((layer2_outputs(7347)) xor (layer2_outputs(7084)));
    layer3_outputs(4940) <= not((layer2_outputs(7581)) or (layer2_outputs(40)));
    layer3_outputs(4941) <= layer2_outputs(696);
    layer3_outputs(4942) <= layer2_outputs(1448);
    layer3_outputs(4943) <= not(layer2_outputs(26));
    layer3_outputs(4944) <= (layer2_outputs(6724)) and (layer2_outputs(6616));
    layer3_outputs(4945) <= not((layer2_outputs(1336)) or (layer2_outputs(4158)));
    layer3_outputs(4946) <= not(layer2_outputs(5284));
    layer3_outputs(4947) <= not((layer2_outputs(17)) or (layer2_outputs(5772)));
    layer3_outputs(4948) <= (layer2_outputs(6619)) and (layer2_outputs(1175));
    layer3_outputs(4949) <= (layer2_outputs(5972)) and not (layer2_outputs(4472));
    layer3_outputs(4950) <= (layer2_outputs(2568)) or (layer2_outputs(157));
    layer3_outputs(4951) <= not((layer2_outputs(2979)) or (layer2_outputs(6050)));
    layer3_outputs(4952) <= not((layer2_outputs(429)) xor (layer2_outputs(1431)));
    layer3_outputs(4953) <= layer2_outputs(6990);
    layer3_outputs(4954) <= layer2_outputs(5397);
    layer3_outputs(4955) <= layer2_outputs(105);
    layer3_outputs(4956) <= not((layer2_outputs(6429)) or (layer2_outputs(6667)));
    layer3_outputs(4957) <= layer2_outputs(7669);
    layer3_outputs(4958) <= not(layer2_outputs(1863)) or (layer2_outputs(1723));
    layer3_outputs(4959) <= layer2_outputs(4541);
    layer3_outputs(4960) <= not(layer2_outputs(207));
    layer3_outputs(4961) <= not((layer2_outputs(5463)) and (layer2_outputs(7593)));
    layer3_outputs(4962) <= not(layer2_outputs(4952));
    layer3_outputs(4963) <= (layer2_outputs(5244)) xor (layer2_outputs(2770));
    layer3_outputs(4964) <= not((layer2_outputs(1908)) or (layer2_outputs(599)));
    layer3_outputs(4965) <= (layer2_outputs(1742)) and (layer2_outputs(3792));
    layer3_outputs(4966) <= layer2_outputs(5631);
    layer3_outputs(4967) <= (layer2_outputs(3936)) and (layer2_outputs(76));
    layer3_outputs(4968) <= (layer2_outputs(6617)) and not (layer2_outputs(3862));
    layer3_outputs(4969) <= not(layer2_outputs(4631));
    layer3_outputs(4970) <= not((layer2_outputs(6058)) or (layer2_outputs(4080)));
    layer3_outputs(4971) <= (layer2_outputs(3950)) and (layer2_outputs(4305));
    layer3_outputs(4972) <= not(layer2_outputs(2397));
    layer3_outputs(4973) <= not(layer2_outputs(2612)) or (layer2_outputs(3844));
    layer3_outputs(4974) <= layer2_outputs(3131);
    layer3_outputs(4975) <= not((layer2_outputs(7556)) xor (layer2_outputs(2550)));
    layer3_outputs(4976) <= not(layer2_outputs(96));
    layer3_outputs(4977) <= not(layer2_outputs(7455));
    layer3_outputs(4978) <= (layer2_outputs(1695)) and not (layer2_outputs(7526));
    layer3_outputs(4979) <= layer2_outputs(4734);
    layer3_outputs(4980) <= layer2_outputs(6411);
    layer3_outputs(4981) <= not((layer2_outputs(2034)) and (layer2_outputs(3512)));
    layer3_outputs(4982) <= not(layer2_outputs(6203)) or (layer2_outputs(5219));
    layer3_outputs(4983) <= layer2_outputs(5999);
    layer3_outputs(4984) <= (layer2_outputs(5199)) and not (layer2_outputs(5439));
    layer3_outputs(4985) <= not(layer2_outputs(4513)) or (layer2_outputs(3270));
    layer3_outputs(4986) <= not(layer2_outputs(2263));
    layer3_outputs(4987) <= (layer2_outputs(5586)) and (layer2_outputs(3928));
    layer3_outputs(4988) <= '0';
    layer3_outputs(4989) <= layer2_outputs(7481);
    layer3_outputs(4990) <= layer2_outputs(121);
    layer3_outputs(4991) <= not((layer2_outputs(5139)) xor (layer2_outputs(7086)));
    layer3_outputs(4992) <= not(layer2_outputs(873));
    layer3_outputs(4993) <= (layer2_outputs(5715)) and not (layer2_outputs(3659));
    layer3_outputs(4994) <= (layer2_outputs(731)) and not (layer2_outputs(2938));
    layer3_outputs(4995) <= not(layer2_outputs(391));
    layer3_outputs(4996) <= '1';
    layer3_outputs(4997) <= layer2_outputs(7107);
    layer3_outputs(4998) <= (layer2_outputs(1438)) and not (layer2_outputs(2370));
    layer3_outputs(4999) <= (layer2_outputs(2607)) and not (layer2_outputs(4682));
    layer3_outputs(5000) <= not(layer2_outputs(2604));
    layer3_outputs(5001) <= not(layer2_outputs(5539));
    layer3_outputs(5002) <= not(layer2_outputs(160));
    layer3_outputs(5003) <= not((layer2_outputs(7479)) or (layer2_outputs(3705)));
    layer3_outputs(5004) <= layer2_outputs(3748);
    layer3_outputs(5005) <= (layer2_outputs(6863)) and not (layer2_outputs(6531));
    layer3_outputs(5006) <= layer2_outputs(4485);
    layer3_outputs(5007) <= not(layer2_outputs(756)) or (layer2_outputs(5639));
    layer3_outputs(5008) <= not(layer2_outputs(1032));
    layer3_outputs(5009) <= not((layer2_outputs(4393)) or (layer2_outputs(7465)));
    layer3_outputs(5010) <= not(layer2_outputs(2696));
    layer3_outputs(5011) <= not((layer2_outputs(2189)) or (layer2_outputs(52)));
    layer3_outputs(5012) <= not(layer2_outputs(4934));
    layer3_outputs(5013) <= not(layer2_outputs(6313)) or (layer2_outputs(678));
    layer3_outputs(5014) <= not(layer2_outputs(3279));
    layer3_outputs(5015) <= layer2_outputs(4380);
    layer3_outputs(5016) <= not(layer2_outputs(7620));
    layer3_outputs(5017) <= not(layer2_outputs(6275));
    layer3_outputs(5018) <= not((layer2_outputs(6708)) and (layer2_outputs(4110)));
    layer3_outputs(5019) <= not((layer2_outputs(5045)) xor (layer2_outputs(2260)));
    layer3_outputs(5020) <= (layer2_outputs(3466)) or (layer2_outputs(1845));
    layer3_outputs(5021) <= (layer2_outputs(3391)) and not (layer2_outputs(6626));
    layer3_outputs(5022) <= (layer2_outputs(108)) and not (layer2_outputs(574));
    layer3_outputs(5023) <= layer2_outputs(6005);
    layer3_outputs(5024) <= not((layer2_outputs(3052)) and (layer2_outputs(4006)));
    layer3_outputs(5025) <= '0';
    layer3_outputs(5026) <= not(layer2_outputs(4669));
    layer3_outputs(5027) <= (layer2_outputs(62)) and (layer2_outputs(5368));
    layer3_outputs(5028) <= layer2_outputs(3599);
    layer3_outputs(5029) <= not((layer2_outputs(4294)) or (layer2_outputs(2708)));
    layer3_outputs(5030) <= (layer2_outputs(3865)) xor (layer2_outputs(2541));
    layer3_outputs(5031) <= (layer2_outputs(1542)) and (layer2_outputs(3101));
    layer3_outputs(5032) <= '1';
    layer3_outputs(5033) <= '0';
    layer3_outputs(5034) <= not(layer2_outputs(2258));
    layer3_outputs(5035) <= not((layer2_outputs(3725)) xor (layer2_outputs(3354)));
    layer3_outputs(5036) <= (layer2_outputs(5598)) and not (layer2_outputs(3448));
    layer3_outputs(5037) <= (layer2_outputs(1115)) or (layer2_outputs(7661));
    layer3_outputs(5038) <= not(layer2_outputs(986)) or (layer2_outputs(683));
    layer3_outputs(5039) <= layer2_outputs(5231);
    layer3_outputs(5040) <= not((layer2_outputs(3257)) and (layer2_outputs(3145)));
    layer3_outputs(5041) <= not(layer2_outputs(5959));
    layer3_outputs(5042) <= (layer2_outputs(4841)) and not (layer2_outputs(6069));
    layer3_outputs(5043) <= layer2_outputs(6407);
    layer3_outputs(5044) <= not(layer2_outputs(1111));
    layer3_outputs(5045) <= (layer2_outputs(4318)) xor (layer2_outputs(1704));
    layer3_outputs(5046) <= not((layer2_outputs(180)) or (layer2_outputs(2025)));
    layer3_outputs(5047) <= not(layer2_outputs(28)) or (layer2_outputs(2537));
    layer3_outputs(5048) <= not(layer2_outputs(3206));
    layer3_outputs(5049) <= not(layer2_outputs(5385));
    layer3_outputs(5050) <= not((layer2_outputs(6148)) and (layer2_outputs(90)));
    layer3_outputs(5051) <= not(layer2_outputs(1082)) or (layer2_outputs(3438));
    layer3_outputs(5052) <= not((layer2_outputs(4128)) or (layer2_outputs(7639)));
    layer3_outputs(5053) <= not(layer2_outputs(7560));
    layer3_outputs(5054) <= layer2_outputs(7267);
    layer3_outputs(5055) <= layer2_outputs(6953);
    layer3_outputs(5056) <= layer2_outputs(2687);
    layer3_outputs(5057) <= (layer2_outputs(5627)) and not (layer2_outputs(3863));
    layer3_outputs(5058) <= not(layer2_outputs(7206));
    layer3_outputs(5059) <= layer2_outputs(2096);
    layer3_outputs(5060) <= not(layer2_outputs(6261));
    layer3_outputs(5061) <= layer2_outputs(4020);
    layer3_outputs(5062) <= layer2_outputs(1995);
    layer3_outputs(5063) <= (layer2_outputs(7629)) and (layer2_outputs(2332));
    layer3_outputs(5064) <= not(layer2_outputs(1769));
    layer3_outputs(5065) <= not(layer2_outputs(6456)) or (layer2_outputs(3339));
    layer3_outputs(5066) <= (layer2_outputs(463)) or (layer2_outputs(7401));
    layer3_outputs(5067) <= (layer2_outputs(3125)) or (layer2_outputs(37));
    layer3_outputs(5068) <= (layer2_outputs(5748)) and (layer2_outputs(3738));
    layer3_outputs(5069) <= not(layer2_outputs(5257)) or (layer2_outputs(1745));
    layer3_outputs(5070) <= not((layer2_outputs(3925)) or (layer2_outputs(5291)));
    layer3_outputs(5071) <= not(layer2_outputs(3255));
    layer3_outputs(5072) <= layer2_outputs(4072);
    layer3_outputs(5073) <= not(layer2_outputs(6891)) or (layer2_outputs(4039));
    layer3_outputs(5074) <= (layer2_outputs(6777)) and (layer2_outputs(824));
    layer3_outputs(5075) <= layer2_outputs(5289);
    layer3_outputs(5076) <= not(layer2_outputs(49)) or (layer2_outputs(2755));
    layer3_outputs(5077) <= (layer2_outputs(3319)) xor (layer2_outputs(6486));
    layer3_outputs(5078) <= not(layer2_outputs(1294));
    layer3_outputs(5079) <= not((layer2_outputs(6728)) and (layer2_outputs(4408)));
    layer3_outputs(5080) <= not(layer2_outputs(1221));
    layer3_outputs(5081) <= not(layer2_outputs(7014));
    layer3_outputs(5082) <= not(layer2_outputs(3255)) or (layer2_outputs(2050));
    layer3_outputs(5083) <= not((layer2_outputs(2267)) xor (layer2_outputs(984)));
    layer3_outputs(5084) <= not(layer2_outputs(1880));
    layer3_outputs(5085) <= not(layer2_outputs(5672));
    layer3_outputs(5086) <= (layer2_outputs(1936)) and not (layer2_outputs(3781));
    layer3_outputs(5087) <= layer2_outputs(2182);
    layer3_outputs(5088) <= not(layer2_outputs(2033));
    layer3_outputs(5089) <= not(layer2_outputs(3478)) or (layer2_outputs(6187));
    layer3_outputs(5090) <= not(layer2_outputs(2146)) or (layer2_outputs(625));
    layer3_outputs(5091) <= layer2_outputs(4157);
    layer3_outputs(5092) <= not((layer2_outputs(5845)) xor (layer2_outputs(2592)));
    layer3_outputs(5093) <= (layer2_outputs(5077)) and not (layer2_outputs(7227));
    layer3_outputs(5094) <= not(layer2_outputs(5528)) or (layer2_outputs(1849));
    layer3_outputs(5095) <= not(layer2_outputs(6223));
    layer3_outputs(5096) <= not(layer2_outputs(4622));
    layer3_outputs(5097) <= not(layer2_outputs(4124)) or (layer2_outputs(7599));
    layer3_outputs(5098) <= not(layer2_outputs(5878));
    layer3_outputs(5099) <= not(layer2_outputs(3620));
    layer3_outputs(5100) <= (layer2_outputs(5540)) and (layer2_outputs(2120));
    layer3_outputs(5101) <= not(layer2_outputs(7564)) or (layer2_outputs(153));
    layer3_outputs(5102) <= not(layer2_outputs(7417));
    layer3_outputs(5103) <= not(layer2_outputs(4097)) or (layer2_outputs(4354));
    layer3_outputs(5104) <= (layer2_outputs(5623)) xor (layer2_outputs(7347));
    layer3_outputs(5105) <= (layer2_outputs(4769)) or (layer2_outputs(7208));
    layer3_outputs(5106) <= (layer2_outputs(698)) and (layer2_outputs(4192));
    layer3_outputs(5107) <= not(layer2_outputs(6472));
    layer3_outputs(5108) <= not((layer2_outputs(2861)) xor (layer2_outputs(5069)));
    layer3_outputs(5109) <= not(layer2_outputs(5064));
    layer3_outputs(5110) <= layer2_outputs(3100);
    layer3_outputs(5111) <= not(layer2_outputs(7622));
    layer3_outputs(5112) <= not((layer2_outputs(2463)) and (layer2_outputs(4038)));
    layer3_outputs(5113) <= (layer2_outputs(1685)) and (layer2_outputs(381));
    layer3_outputs(5114) <= not((layer2_outputs(2496)) or (layer2_outputs(804)));
    layer3_outputs(5115) <= layer2_outputs(5023);
    layer3_outputs(5116) <= (layer2_outputs(4934)) and not (layer2_outputs(1529));
    layer3_outputs(5117) <= layer2_outputs(7081);
    layer3_outputs(5118) <= not((layer2_outputs(256)) xor (layer2_outputs(959)));
    layer3_outputs(5119) <= layer2_outputs(5778);
    layer3_outputs(5120) <= (layer2_outputs(1371)) and not (layer2_outputs(5000));
    layer3_outputs(5121) <= layer2_outputs(6018);
    layer3_outputs(5122) <= not(layer2_outputs(4169));
    layer3_outputs(5123) <= layer2_outputs(5853);
    layer3_outputs(5124) <= not(layer2_outputs(2750));
    layer3_outputs(5125) <= not(layer2_outputs(5555));
    layer3_outputs(5126) <= not(layer2_outputs(6676));
    layer3_outputs(5127) <= not(layer2_outputs(4756));
    layer3_outputs(5128) <= not(layer2_outputs(5603));
    layer3_outputs(5129) <= not(layer2_outputs(2661));
    layer3_outputs(5130) <= layer2_outputs(4829);
    layer3_outputs(5131) <= not(layer2_outputs(5831));
    layer3_outputs(5132) <= '0';
    layer3_outputs(5133) <= not((layer2_outputs(3593)) and (layer2_outputs(653)));
    layer3_outputs(5134) <= (layer2_outputs(5127)) and not (layer2_outputs(5973));
    layer3_outputs(5135) <= layer2_outputs(5201);
    layer3_outputs(5136) <= not((layer2_outputs(7650)) xor (layer2_outputs(3491)));
    layer3_outputs(5137) <= layer2_outputs(6857);
    layer3_outputs(5138) <= not(layer2_outputs(4035));
    layer3_outputs(5139) <= layer2_outputs(2647);
    layer3_outputs(5140) <= layer2_outputs(6908);
    layer3_outputs(5141) <= not(layer2_outputs(6409));
    layer3_outputs(5142) <= not(layer2_outputs(4221)) or (layer2_outputs(3870));
    layer3_outputs(5143) <= not(layer2_outputs(3945));
    layer3_outputs(5144) <= not(layer2_outputs(3840));
    layer3_outputs(5145) <= '1';
    layer3_outputs(5146) <= not(layer2_outputs(1125));
    layer3_outputs(5147) <= not((layer2_outputs(7410)) or (layer2_outputs(7503)));
    layer3_outputs(5148) <= '1';
    layer3_outputs(5149) <= layer2_outputs(1021);
    layer3_outputs(5150) <= (layer2_outputs(1630)) and not (layer2_outputs(5988));
    layer3_outputs(5151) <= layer2_outputs(3031);
    layer3_outputs(5152) <= not(layer2_outputs(7245));
    layer3_outputs(5153) <= layer2_outputs(7583);
    layer3_outputs(5154) <= not((layer2_outputs(7232)) or (layer2_outputs(3830)));
    layer3_outputs(5155) <= layer2_outputs(4647);
    layer3_outputs(5156) <= not(layer2_outputs(4312));
    layer3_outputs(5157) <= not(layer2_outputs(6625)) or (layer2_outputs(1171));
    layer3_outputs(5158) <= not(layer2_outputs(1367)) or (layer2_outputs(5072));
    layer3_outputs(5159) <= layer2_outputs(6868);
    layer3_outputs(5160) <= layer2_outputs(5546);
    layer3_outputs(5161) <= (layer2_outputs(1273)) and (layer2_outputs(7425));
    layer3_outputs(5162) <= not(layer2_outputs(2354));
    layer3_outputs(5163) <= (layer2_outputs(6167)) and not (layer2_outputs(1894));
    layer3_outputs(5164) <= not((layer2_outputs(7151)) and (layer2_outputs(616)));
    layer3_outputs(5165) <= (layer2_outputs(1687)) or (layer2_outputs(7511));
    layer3_outputs(5166) <= (layer2_outputs(4713)) or (layer2_outputs(1608));
    layer3_outputs(5167) <= layer2_outputs(1154);
    layer3_outputs(5168) <= (layer2_outputs(7288)) and not (layer2_outputs(758));
    layer3_outputs(5169) <= not(layer2_outputs(2442));
    layer3_outputs(5170) <= (layer2_outputs(3776)) or (layer2_outputs(4369));
    layer3_outputs(5171) <= not((layer2_outputs(3102)) or (layer2_outputs(3355)));
    layer3_outputs(5172) <= layer2_outputs(4181);
    layer3_outputs(5173) <= (layer2_outputs(1592)) and not (layer2_outputs(3337));
    layer3_outputs(5174) <= not(layer2_outputs(3127));
    layer3_outputs(5175) <= layer2_outputs(5321);
    layer3_outputs(5176) <= not(layer2_outputs(5043));
    layer3_outputs(5177) <= layer2_outputs(4661);
    layer3_outputs(5178) <= (layer2_outputs(2022)) and (layer2_outputs(2535));
    layer3_outputs(5179) <= layer2_outputs(2910);
    layer3_outputs(5180) <= (layer2_outputs(6039)) xor (layer2_outputs(300));
    layer3_outputs(5181) <= not(layer2_outputs(5245));
    layer3_outputs(5182) <= not(layer2_outputs(648));
    layer3_outputs(5183) <= layer2_outputs(2843);
    layer3_outputs(5184) <= (layer2_outputs(2628)) or (layer2_outputs(4684));
    layer3_outputs(5185) <= layer2_outputs(3368);
    layer3_outputs(5186) <= layer2_outputs(1149);
    layer3_outputs(5187) <= not(layer2_outputs(165)) or (layer2_outputs(6437));
    layer3_outputs(5188) <= layer2_outputs(4015);
    layer3_outputs(5189) <= (layer2_outputs(1851)) and not (layer2_outputs(2334));
    layer3_outputs(5190) <= '1';
    layer3_outputs(5191) <= (layer2_outputs(3969)) xor (layer2_outputs(5976));
    layer3_outputs(5192) <= not(layer2_outputs(7667));
    layer3_outputs(5193) <= not((layer2_outputs(2713)) xor (layer2_outputs(2975)));
    layer3_outputs(5194) <= layer2_outputs(3134);
    layer3_outputs(5195) <= '0';
    layer3_outputs(5196) <= (layer2_outputs(4050)) and not (layer2_outputs(3369));
    layer3_outputs(5197) <= not((layer2_outputs(5249)) or (layer2_outputs(6337)));
    layer3_outputs(5198) <= '1';
    layer3_outputs(5199) <= layer2_outputs(1418);
    layer3_outputs(5200) <= not(layer2_outputs(3590)) or (layer2_outputs(6851));
    layer3_outputs(5201) <= not(layer2_outputs(4532));
    layer3_outputs(5202) <= not((layer2_outputs(689)) xor (layer2_outputs(6750)));
    layer3_outputs(5203) <= not((layer2_outputs(5891)) or (layer2_outputs(6142)));
    layer3_outputs(5204) <= not(layer2_outputs(5323));
    layer3_outputs(5205) <= (layer2_outputs(3669)) and not (layer2_outputs(2204));
    layer3_outputs(5206) <= not(layer2_outputs(7596));
    layer3_outputs(5207) <= layer2_outputs(4213);
    layer3_outputs(5208) <= (layer2_outputs(3809)) or (layer2_outputs(6213));
    layer3_outputs(5209) <= layer2_outputs(2148);
    layer3_outputs(5210) <= not(layer2_outputs(1377));
    layer3_outputs(5211) <= not(layer2_outputs(265));
    layer3_outputs(5212) <= layer2_outputs(1899);
    layer3_outputs(5213) <= layer2_outputs(5935);
    layer3_outputs(5214) <= (layer2_outputs(3131)) and not (layer2_outputs(65));
    layer3_outputs(5215) <= (layer2_outputs(1541)) and not (layer2_outputs(3585));
    layer3_outputs(5216) <= not(layer2_outputs(2062)) or (layer2_outputs(5799));
    layer3_outputs(5217) <= not(layer2_outputs(7203));
    layer3_outputs(5218) <= not((layer2_outputs(2775)) or (layer2_outputs(3593)));
    layer3_outputs(5219) <= layer2_outputs(3401);
    layer3_outputs(5220) <= not(layer2_outputs(926));
    layer3_outputs(5221) <= not((layer2_outputs(6402)) or (layer2_outputs(3373)));
    layer3_outputs(5222) <= not(layer2_outputs(935));
    layer3_outputs(5223) <= layer2_outputs(2081);
    layer3_outputs(5224) <= layer2_outputs(7388);
    layer3_outputs(5225) <= not((layer2_outputs(3772)) or (layer2_outputs(210)));
    layer3_outputs(5226) <= layer2_outputs(1133);
    layer3_outputs(5227) <= not(layer2_outputs(7499));
    layer3_outputs(5228) <= (layer2_outputs(5138)) or (layer2_outputs(5655));
    layer3_outputs(5229) <= not(layer2_outputs(1120)) or (layer2_outputs(2620));
    layer3_outputs(5230) <= not(layer2_outputs(7357));
    layer3_outputs(5231) <= not(layer2_outputs(6175));
    layer3_outputs(5232) <= not(layer2_outputs(5623));
    layer3_outputs(5233) <= (layer2_outputs(6805)) xor (layer2_outputs(7365));
    layer3_outputs(5234) <= (layer2_outputs(7366)) and not (layer2_outputs(6872));
    layer3_outputs(5235) <= not(layer2_outputs(5870)) or (layer2_outputs(370));
    layer3_outputs(5236) <= layer2_outputs(5323);
    layer3_outputs(5237) <= (layer2_outputs(6537)) and not (layer2_outputs(4978));
    layer3_outputs(5238) <= (layer2_outputs(7220)) and not (layer2_outputs(3043));
    layer3_outputs(5239) <= not(layer2_outputs(1187)) or (layer2_outputs(2992));
    layer3_outputs(5240) <= layer2_outputs(5121);
    layer3_outputs(5241) <= layer2_outputs(2585);
    layer3_outputs(5242) <= (layer2_outputs(1585)) or (layer2_outputs(3547));
    layer3_outputs(5243) <= layer2_outputs(4743);
    layer3_outputs(5244) <= not(layer2_outputs(2200));
    layer3_outputs(5245) <= layer2_outputs(7646);
    layer3_outputs(5246) <= layer2_outputs(6274);
    layer3_outputs(5247) <= layer2_outputs(3025);
    layer3_outputs(5248) <= not(layer2_outputs(7402)) or (layer2_outputs(4292));
    layer3_outputs(5249) <= not(layer2_outputs(2422));
    layer3_outputs(5250) <= not(layer2_outputs(887)) or (layer2_outputs(1969));
    layer3_outputs(5251) <= '0';
    layer3_outputs(5252) <= not((layer2_outputs(3617)) or (layer2_outputs(5277)));
    layer3_outputs(5253) <= layer2_outputs(2697);
    layer3_outputs(5254) <= layer2_outputs(736);
    layer3_outputs(5255) <= (layer2_outputs(3357)) and not (layer2_outputs(7308));
    layer3_outputs(5256) <= not(layer2_outputs(5791)) or (layer2_outputs(2));
    layer3_outputs(5257) <= (layer2_outputs(3835)) xor (layer2_outputs(3322));
    layer3_outputs(5258) <= (layer2_outputs(6920)) or (layer2_outputs(605));
    layer3_outputs(5259) <= (layer2_outputs(1786)) and (layer2_outputs(5912));
    layer3_outputs(5260) <= not(layer2_outputs(5865)) or (layer2_outputs(5954));
    layer3_outputs(5261) <= not(layer2_outputs(2541));
    layer3_outputs(5262) <= (layer2_outputs(1832)) and (layer2_outputs(3265));
    layer3_outputs(5263) <= not((layer2_outputs(2732)) and (layer2_outputs(6859)));
    layer3_outputs(5264) <= not((layer2_outputs(2410)) or (layer2_outputs(5475)));
    layer3_outputs(5265) <= not((layer2_outputs(2485)) or (layer2_outputs(5745)));
    layer3_outputs(5266) <= (layer2_outputs(2017)) and not (layer2_outputs(6921));
    layer3_outputs(5267) <= (layer2_outputs(1430)) or (layer2_outputs(2525));
    layer3_outputs(5268) <= layer2_outputs(6726);
    layer3_outputs(5269) <= not(layer2_outputs(4557)) or (layer2_outputs(4717));
    layer3_outputs(5270) <= not(layer2_outputs(1484));
    layer3_outputs(5271) <= (layer2_outputs(1565)) and (layer2_outputs(4593));
    layer3_outputs(5272) <= (layer2_outputs(1962)) and not (layer2_outputs(7306));
    layer3_outputs(5273) <= '1';
    layer3_outputs(5274) <= layer2_outputs(1946);
    layer3_outputs(5275) <= layer2_outputs(1733);
    layer3_outputs(5276) <= not(layer2_outputs(1963)) or (layer2_outputs(5071));
    layer3_outputs(5277) <= (layer2_outputs(6546)) and (layer2_outputs(5444));
    layer3_outputs(5278) <= (layer2_outputs(82)) or (layer2_outputs(923));
    layer3_outputs(5279) <= not(layer2_outputs(3831)) or (layer2_outputs(2434));
    layer3_outputs(5280) <= (layer2_outputs(3569)) and not (layer2_outputs(6520));
    layer3_outputs(5281) <= not(layer2_outputs(4549)) or (layer2_outputs(6529));
    layer3_outputs(5282) <= not(layer2_outputs(6206));
    layer3_outputs(5283) <= not((layer2_outputs(752)) and (layer2_outputs(1426)));
    layer3_outputs(5284) <= not((layer2_outputs(3289)) or (layer2_outputs(3666)));
    layer3_outputs(5285) <= not(layer2_outputs(1677));
    layer3_outputs(5286) <= layer2_outputs(2651);
    layer3_outputs(5287) <= '1';
    layer3_outputs(5288) <= not(layer2_outputs(3625));
    layer3_outputs(5289) <= not(layer2_outputs(3217));
    layer3_outputs(5290) <= (layer2_outputs(6765)) or (layer2_outputs(582));
    layer3_outputs(5291) <= not(layer2_outputs(6764));
    layer3_outputs(5292) <= not((layer2_outputs(482)) or (layer2_outputs(1037)));
    layer3_outputs(5293) <= layer2_outputs(7280);
    layer3_outputs(5294) <= not((layer2_outputs(2583)) or (layer2_outputs(2132)));
    layer3_outputs(5295) <= not(layer2_outputs(104)) or (layer2_outputs(6368));
    layer3_outputs(5296) <= (layer2_outputs(7257)) and not (layer2_outputs(1112));
    layer3_outputs(5297) <= layer2_outputs(5423);
    layer3_outputs(5298) <= not(layer2_outputs(1710)) or (layer2_outputs(3682));
    layer3_outputs(5299) <= layer2_outputs(5296);
    layer3_outputs(5300) <= (layer2_outputs(700)) or (layer2_outputs(904));
    layer3_outputs(5301) <= (layer2_outputs(3972)) and not (layer2_outputs(7307));
    layer3_outputs(5302) <= layer2_outputs(3452);
    layer3_outputs(5303) <= (layer2_outputs(2303)) and not (layer2_outputs(4131));
    layer3_outputs(5304) <= not(layer2_outputs(4421));
    layer3_outputs(5305) <= not((layer2_outputs(5769)) or (layer2_outputs(2264)));
    layer3_outputs(5306) <= layer2_outputs(303);
    layer3_outputs(5307) <= (layer2_outputs(5071)) and not (layer2_outputs(3266));
    layer3_outputs(5308) <= not(layer2_outputs(2530));
    layer3_outputs(5309) <= (layer2_outputs(6495)) or (layer2_outputs(6835));
    layer3_outputs(5310) <= not(layer2_outputs(6635));
    layer3_outputs(5311) <= layer2_outputs(7473);
    layer3_outputs(5312) <= not((layer2_outputs(4488)) or (layer2_outputs(2110)));
    layer3_outputs(5313) <= (layer2_outputs(2139)) and not (layer2_outputs(1161));
    layer3_outputs(5314) <= not(layer2_outputs(5544)) or (layer2_outputs(4512));
    layer3_outputs(5315) <= '0';
    layer3_outputs(5316) <= not(layer2_outputs(3368));
    layer3_outputs(5317) <= (layer2_outputs(2598)) and not (layer2_outputs(5921));
    layer3_outputs(5318) <= not(layer2_outputs(6));
    layer3_outputs(5319) <= not((layer2_outputs(102)) or (layer2_outputs(151)));
    layer3_outputs(5320) <= layer2_outputs(383);
    layer3_outputs(5321) <= not(layer2_outputs(5762));
    layer3_outputs(5322) <= not(layer2_outputs(81));
    layer3_outputs(5323) <= layer2_outputs(4662);
    layer3_outputs(5324) <= (layer2_outputs(3022)) or (layer2_outputs(1915));
    layer3_outputs(5325) <= layer2_outputs(4255);
    layer3_outputs(5326) <= (layer2_outputs(6672)) and (layer2_outputs(6935));
    layer3_outputs(5327) <= not(layer2_outputs(5713));
    layer3_outputs(5328) <= not(layer2_outputs(7062));
    layer3_outputs(5329) <= not(layer2_outputs(812));
    layer3_outputs(5330) <= not((layer2_outputs(5187)) and (layer2_outputs(2554)));
    layer3_outputs(5331) <= not((layer2_outputs(857)) and (layer2_outputs(7657)));
    layer3_outputs(5332) <= layer2_outputs(6898);
    layer3_outputs(5333) <= (layer2_outputs(2749)) and not (layer2_outputs(3412));
    layer3_outputs(5334) <= not(layer2_outputs(1814));
    layer3_outputs(5335) <= layer2_outputs(1291);
    layer3_outputs(5336) <= layer2_outputs(4973);
    layer3_outputs(5337) <= (layer2_outputs(6794)) and not (layer2_outputs(2552));
    layer3_outputs(5338) <= not((layer2_outputs(4962)) or (layer2_outputs(2296)));
    layer3_outputs(5339) <= layer2_outputs(5586);
    layer3_outputs(5340) <= not(layer2_outputs(3984));
    layer3_outputs(5341) <= not((layer2_outputs(6042)) and (layer2_outputs(6714)));
    layer3_outputs(5342) <= not(layer2_outputs(664)) or (layer2_outputs(1293));
    layer3_outputs(5343) <= not(layer2_outputs(2637)) or (layer2_outputs(3694));
    layer3_outputs(5344) <= not(layer2_outputs(1080));
    layer3_outputs(5345) <= layer2_outputs(3353);
    layer3_outputs(5346) <= layer2_outputs(825);
    layer3_outputs(5347) <= layer2_outputs(5159);
    layer3_outputs(5348) <= layer2_outputs(5619);
    layer3_outputs(5349) <= layer2_outputs(5597);
    layer3_outputs(5350) <= not((layer2_outputs(2998)) xor (layer2_outputs(6637)));
    layer3_outputs(5351) <= '1';
    layer3_outputs(5352) <= layer2_outputs(4433);
    layer3_outputs(5353) <= not(layer2_outputs(6215)) or (layer2_outputs(3176));
    layer3_outputs(5354) <= (layer2_outputs(211)) xor (layer2_outputs(161));
    layer3_outputs(5355) <= '1';
    layer3_outputs(5356) <= not(layer2_outputs(6108));
    layer3_outputs(5357) <= not((layer2_outputs(133)) or (layer2_outputs(7116)));
    layer3_outputs(5358) <= layer2_outputs(3715);
    layer3_outputs(5359) <= not((layer2_outputs(2193)) and (layer2_outputs(4071)));
    layer3_outputs(5360) <= layer2_outputs(2424);
    layer3_outputs(5361) <= layer2_outputs(2977);
    layer3_outputs(5362) <= '1';
    layer3_outputs(5363) <= not((layer2_outputs(1528)) and (layer2_outputs(1258)));
    layer3_outputs(5364) <= not(layer2_outputs(3202));
    layer3_outputs(5365) <= (layer2_outputs(2599)) and not (layer2_outputs(1773));
    layer3_outputs(5366) <= (layer2_outputs(260)) and not (layer2_outputs(1385));
    layer3_outputs(5367) <= not(layer2_outputs(3939));
    layer3_outputs(5368) <= not(layer2_outputs(6843));
    layer3_outputs(5369) <= layer2_outputs(6467);
    layer3_outputs(5370) <= not(layer2_outputs(650));
    layer3_outputs(5371) <= layer2_outputs(3200);
    layer3_outputs(5372) <= layer2_outputs(2336);
    layer3_outputs(5373) <= not(layer2_outputs(4057));
    layer3_outputs(5374) <= not(layer2_outputs(6459)) or (layer2_outputs(2219));
    layer3_outputs(5375) <= not(layer2_outputs(7073));
    layer3_outputs(5376) <= not((layer2_outputs(4928)) and (layer2_outputs(6849)));
    layer3_outputs(5377) <= layer2_outputs(5273);
    layer3_outputs(5378) <= not(layer2_outputs(2458));
    layer3_outputs(5379) <= layer2_outputs(5036);
    layer3_outputs(5380) <= not(layer2_outputs(6931));
    layer3_outputs(5381) <= (layer2_outputs(3471)) and not (layer2_outputs(3873));
    layer3_outputs(5382) <= not(layer2_outputs(851)) or (layer2_outputs(2548));
    layer3_outputs(5383) <= not(layer2_outputs(6880));
    layer3_outputs(5384) <= (layer2_outputs(3643)) or (layer2_outputs(5643));
    layer3_outputs(5385) <= not(layer2_outputs(5774));
    layer3_outputs(5386) <= not((layer2_outputs(3940)) and (layer2_outputs(1274)));
    layer3_outputs(5387) <= (layer2_outputs(3485)) and not (layer2_outputs(7374));
    layer3_outputs(5388) <= (layer2_outputs(5489)) and (layer2_outputs(4387));
    layer3_outputs(5389) <= not(layer2_outputs(6215)) or (layer2_outputs(2198));
    layer3_outputs(5390) <= not(layer2_outputs(1284)) or (layer2_outputs(7107));
    layer3_outputs(5391) <= not(layer2_outputs(3966)) or (layer2_outputs(1546));
    layer3_outputs(5392) <= layer2_outputs(4165);
    layer3_outputs(5393) <= not(layer2_outputs(4281));
    layer3_outputs(5394) <= not((layer2_outputs(6307)) xor (layer2_outputs(4683)));
    layer3_outputs(5395) <= layer2_outputs(5352);
    layer3_outputs(5396) <= not((layer2_outputs(3260)) and (layer2_outputs(6425)));
    layer3_outputs(5397) <= layer2_outputs(4281);
    layer3_outputs(5398) <= not((layer2_outputs(2075)) and (layer2_outputs(4401)));
    layer3_outputs(5399) <= layer2_outputs(1760);
    layer3_outputs(5400) <= not(layer2_outputs(3307));
    layer3_outputs(5401) <= not(layer2_outputs(7388)) or (layer2_outputs(289));
    layer3_outputs(5402) <= not(layer2_outputs(2546));
    layer3_outputs(5403) <= not(layer2_outputs(72));
    layer3_outputs(5404) <= not((layer2_outputs(4578)) or (layer2_outputs(3090)));
    layer3_outputs(5405) <= not(layer2_outputs(6326));
    layer3_outputs(5406) <= not(layer2_outputs(7492));
    layer3_outputs(5407) <= not((layer2_outputs(522)) xor (layer2_outputs(5858)));
    layer3_outputs(5408) <= (layer2_outputs(6887)) and (layer2_outputs(5218));
    layer3_outputs(5409) <= not(layer2_outputs(787)) or (layer2_outputs(3139));
    layer3_outputs(5410) <= (layer2_outputs(313)) and not (layer2_outputs(4194));
    layer3_outputs(5411) <= not((layer2_outputs(354)) and (layer2_outputs(5575)));
    layer3_outputs(5412) <= not(layer2_outputs(2551));
    layer3_outputs(5413) <= '1';
    layer3_outputs(5414) <= (layer2_outputs(5696)) or (layer2_outputs(2997));
    layer3_outputs(5415) <= (layer2_outputs(1463)) xor (layer2_outputs(3755));
    layer3_outputs(5416) <= not(layer2_outputs(3303));
    layer3_outputs(5417) <= (layer2_outputs(4835)) or (layer2_outputs(774));
    layer3_outputs(5418) <= not(layer2_outputs(1989)) or (layer2_outputs(747));
    layer3_outputs(5419) <= not(layer2_outputs(110));
    layer3_outputs(5420) <= not((layer2_outputs(5805)) and (layer2_outputs(4554)));
    layer3_outputs(5421) <= layer2_outputs(5433);
    layer3_outputs(5422) <= (layer2_outputs(4291)) and not (layer2_outputs(3754));
    layer3_outputs(5423) <= not(layer2_outputs(2870)) or (layer2_outputs(484));
    layer3_outputs(5424) <= layer2_outputs(3140);
    layer3_outputs(5425) <= layer2_outputs(4948);
    layer3_outputs(5426) <= not(layer2_outputs(1387));
    layer3_outputs(5427) <= not(layer2_outputs(787));
    layer3_outputs(5428) <= layer2_outputs(6780);
    layer3_outputs(5429) <= not((layer2_outputs(4429)) and (layer2_outputs(5468)));
    layer3_outputs(5430) <= (layer2_outputs(1135)) or (layer2_outputs(6870));
    layer3_outputs(5431) <= (layer2_outputs(458)) and not (layer2_outputs(1337));
    layer3_outputs(5432) <= not(layer2_outputs(6225));
    layer3_outputs(5433) <= not(layer2_outputs(3514));
    layer3_outputs(5434) <= not(layer2_outputs(6029));
    layer3_outputs(5435) <= not(layer2_outputs(6423)) or (layer2_outputs(4767));
    layer3_outputs(5436) <= (layer2_outputs(1265)) or (layer2_outputs(2856));
    layer3_outputs(5437) <= not(layer2_outputs(2349));
    layer3_outputs(5438) <= not((layer2_outputs(4182)) or (layer2_outputs(1820)));
    layer3_outputs(5439) <= not(layer2_outputs(1592));
    layer3_outputs(5440) <= layer2_outputs(6510);
    layer3_outputs(5441) <= not(layer2_outputs(1138)) or (layer2_outputs(4297));
    layer3_outputs(5442) <= (layer2_outputs(2987)) xor (layer2_outputs(2319));
    layer3_outputs(5443) <= (layer2_outputs(3681)) and not (layer2_outputs(2009));
    layer3_outputs(5444) <= not(layer2_outputs(1959)) or (layer2_outputs(4438));
    layer3_outputs(5445) <= (layer2_outputs(4303)) and not (layer2_outputs(2169));
    layer3_outputs(5446) <= layer2_outputs(806);
    layer3_outputs(5447) <= not(layer2_outputs(4465)) or (layer2_outputs(3489));
    layer3_outputs(5448) <= (layer2_outputs(6612)) and not (layer2_outputs(2061));
    layer3_outputs(5449) <= not(layer2_outputs(193)) or (layer2_outputs(5609));
    layer3_outputs(5450) <= not((layer2_outputs(6936)) or (layer2_outputs(1714)));
    layer3_outputs(5451) <= not(layer2_outputs(3553)) or (layer2_outputs(2708));
    layer3_outputs(5452) <= not((layer2_outputs(4252)) xor (layer2_outputs(4958)));
    layer3_outputs(5453) <= layer2_outputs(6383);
    layer3_outputs(5454) <= not((layer2_outputs(1967)) xor (layer2_outputs(4267)));
    layer3_outputs(5455) <= (layer2_outputs(1729)) xor (layer2_outputs(6114));
    layer3_outputs(5456) <= not(layer2_outputs(5753));
    layer3_outputs(5457) <= layer2_outputs(7370);
    layer3_outputs(5458) <= layer2_outputs(4415);
    layer3_outputs(5459) <= (layer2_outputs(1182)) and not (layer2_outputs(2992));
    layer3_outputs(5460) <= not(layer2_outputs(6501));
    layer3_outputs(5461) <= '0';
    layer3_outputs(5462) <= (layer2_outputs(4177)) or (layer2_outputs(2691));
    layer3_outputs(5463) <= layer2_outputs(168);
    layer3_outputs(5464) <= (layer2_outputs(3608)) and not (layer2_outputs(140));
    layer3_outputs(5465) <= not((layer2_outputs(3049)) and (layer2_outputs(6059)));
    layer3_outputs(5466) <= layer2_outputs(6256);
    layer3_outputs(5467) <= not(layer2_outputs(4688));
    layer3_outputs(5468) <= layer2_outputs(4809);
    layer3_outputs(5469) <= layer2_outputs(1386);
    layer3_outputs(5470) <= (layer2_outputs(292)) and (layer2_outputs(6311));
    layer3_outputs(5471) <= layer2_outputs(6288);
    layer3_outputs(5472) <= not(layer2_outputs(2538)) or (layer2_outputs(5980));
    layer3_outputs(5473) <= layer2_outputs(4385);
    layer3_outputs(5474) <= layer2_outputs(583);
    layer3_outputs(5475) <= not(layer2_outputs(7545)) or (layer2_outputs(407));
    layer3_outputs(5476) <= layer2_outputs(5203);
    layer3_outputs(5477) <= (layer2_outputs(1007)) xor (layer2_outputs(6960));
    layer3_outputs(5478) <= not((layer2_outputs(5055)) xor (layer2_outputs(5511)));
    layer3_outputs(5479) <= (layer2_outputs(4522)) and not (layer2_outputs(4268));
    layer3_outputs(5480) <= not((layer2_outputs(6240)) xor (layer2_outputs(2601)));
    layer3_outputs(5481) <= not(layer2_outputs(5877));
    layer3_outputs(5482) <= not(layer2_outputs(3789));
    layer3_outputs(5483) <= (layer2_outputs(2962)) and not (layer2_outputs(3858));
    layer3_outputs(5484) <= not(layer2_outputs(1560)) or (layer2_outputs(3225));
    layer3_outputs(5485) <= not(layer2_outputs(347));
    layer3_outputs(5486) <= (layer2_outputs(2291)) and (layer2_outputs(5848));
    layer3_outputs(5487) <= not(layer2_outputs(6178)) or (layer2_outputs(5462));
    layer3_outputs(5488) <= not(layer2_outputs(4206));
    layer3_outputs(5489) <= (layer2_outputs(1898)) and not (layer2_outputs(4704));
    layer3_outputs(5490) <= not(layer2_outputs(2143));
    layer3_outputs(5491) <= layer2_outputs(915);
    layer3_outputs(5492) <= not((layer2_outputs(1892)) xor (layer2_outputs(2045)));
    layer3_outputs(5493) <= (layer2_outputs(4429)) and (layer2_outputs(3317));
    layer3_outputs(5494) <= (layer2_outputs(1424)) and not (layer2_outputs(6109));
    layer3_outputs(5495) <= not(layer2_outputs(475));
    layer3_outputs(5496) <= not((layer2_outputs(3834)) xor (layer2_outputs(2085)));
    layer3_outputs(5497) <= layer2_outputs(5133);
    layer3_outputs(5498) <= (layer2_outputs(6452)) or (layer2_outputs(2839));
    layer3_outputs(5499) <= layer2_outputs(4605);
    layer3_outputs(5500) <= layer2_outputs(5591);
    layer3_outputs(5501) <= not(layer2_outputs(2730));
    layer3_outputs(5502) <= not((layer2_outputs(3015)) and (layer2_outputs(1727)));
    layer3_outputs(5503) <= layer2_outputs(4495);
    layer3_outputs(5504) <= (layer2_outputs(6621)) and (layer2_outputs(1534));
    layer3_outputs(5505) <= layer2_outputs(6700);
    layer3_outputs(5506) <= (layer2_outputs(1987)) and (layer2_outputs(5232));
    layer3_outputs(5507) <= not(layer2_outputs(2380)) or (layer2_outputs(4546));
    layer3_outputs(5508) <= not((layer2_outputs(3360)) or (layer2_outputs(5314)));
    layer3_outputs(5509) <= (layer2_outputs(630)) xor (layer2_outputs(7184));
    layer3_outputs(5510) <= layer2_outputs(774);
    layer3_outputs(5511) <= not((layer2_outputs(2897)) and (layer2_outputs(7117)));
    layer3_outputs(5512) <= (layer2_outputs(845)) and not (layer2_outputs(5777));
    layer3_outputs(5513) <= not(layer2_outputs(1631));
    layer3_outputs(5514) <= (layer2_outputs(2457)) and (layer2_outputs(334));
    layer3_outputs(5515) <= (layer2_outputs(4827)) and (layer2_outputs(140));
    layer3_outputs(5516) <= (layer2_outputs(3690)) xor (layer2_outputs(3670));
    layer3_outputs(5517) <= not(layer2_outputs(7563));
    layer3_outputs(5518) <= layer2_outputs(4760);
    layer3_outputs(5519) <= layer2_outputs(1076);
    layer3_outputs(5520) <= not(layer2_outputs(3799));
    layer3_outputs(5521) <= (layer2_outputs(7439)) and not (layer2_outputs(5993));
    layer3_outputs(5522) <= layer2_outputs(4940);
    layer3_outputs(5523) <= layer2_outputs(1668);
    layer3_outputs(5524) <= (layer2_outputs(3370)) xor (layer2_outputs(2036));
    layer3_outputs(5525) <= (layer2_outputs(876)) and not (layer2_outputs(3362));
    layer3_outputs(5526) <= not(layer2_outputs(3888));
    layer3_outputs(5527) <= layer2_outputs(1657);
    layer3_outputs(5528) <= (layer2_outputs(7106)) or (layer2_outputs(4750));
    layer3_outputs(5529) <= (layer2_outputs(4636)) and not (layer2_outputs(2368));
    layer3_outputs(5530) <= not((layer2_outputs(2327)) or (layer2_outputs(1601)));
    layer3_outputs(5531) <= not(layer2_outputs(71));
    layer3_outputs(5532) <= layer2_outputs(1222);
    layer3_outputs(5533) <= (layer2_outputs(6301)) and not (layer2_outputs(2877));
    layer3_outputs(5534) <= not(layer2_outputs(3284)) or (layer2_outputs(5947));
    layer3_outputs(5535) <= not(layer2_outputs(7204));
    layer3_outputs(5536) <= (layer2_outputs(7264)) xor (layer2_outputs(646));
    layer3_outputs(5537) <= layer2_outputs(5752);
    layer3_outputs(5538) <= '1';
    layer3_outputs(5539) <= layer2_outputs(3125);
    layer3_outputs(5540) <= '0';
    layer3_outputs(5541) <= not(layer2_outputs(5813));
    layer3_outputs(5542) <= layer2_outputs(1063);
    layer3_outputs(5543) <= (layer2_outputs(1827)) and not (layer2_outputs(7319));
    layer3_outputs(5544) <= not(layer2_outputs(3470));
    layer3_outputs(5545) <= layer2_outputs(1736);
    layer3_outputs(5546) <= not(layer2_outputs(844)) or (layer2_outputs(4444));
    layer3_outputs(5547) <= layer2_outputs(5382);
    layer3_outputs(5548) <= (layer2_outputs(6923)) or (layer2_outputs(1798));
    layer3_outputs(5549) <= not((layer2_outputs(1852)) and (layer2_outputs(6969)));
    layer3_outputs(5550) <= not((layer2_outputs(7497)) or (layer2_outputs(3904)));
    layer3_outputs(5551) <= '0';
    layer3_outputs(5552) <= (layer2_outputs(5705)) and (layer2_outputs(4246));
    layer3_outputs(5553) <= not(layer2_outputs(2783));
    layer3_outputs(5554) <= (layer2_outputs(3262)) and not (layer2_outputs(4594));
    layer3_outputs(5555) <= layer2_outputs(5642);
    layer3_outputs(5556) <= not(layer2_outputs(3417));
    layer3_outputs(5557) <= layer2_outputs(4938);
    layer3_outputs(5558) <= layer2_outputs(5932);
    layer3_outputs(5559) <= layer2_outputs(2635);
    layer3_outputs(5560) <= layer2_outputs(4309);
    layer3_outputs(5561) <= not(layer2_outputs(153));
    layer3_outputs(5562) <= not((layer2_outputs(6787)) or (layer2_outputs(266)));
    layer3_outputs(5563) <= not(layer2_outputs(4248));
    layer3_outputs(5564) <= not(layer2_outputs(2978));
    layer3_outputs(5565) <= not((layer2_outputs(4003)) and (layer2_outputs(4717)));
    layer3_outputs(5566) <= not(layer2_outputs(5929)) or (layer2_outputs(218));
    layer3_outputs(5567) <= (layer2_outputs(5752)) or (layer2_outputs(6033));
    layer3_outputs(5568) <= '0';
    layer3_outputs(5569) <= not(layer2_outputs(4977));
    layer3_outputs(5570) <= not(layer2_outputs(7338));
    layer3_outputs(5571) <= '1';
    layer3_outputs(5572) <= not(layer2_outputs(7413));
    layer3_outputs(5573) <= (layer2_outputs(3977)) or (layer2_outputs(7585));
    layer3_outputs(5574) <= (layer2_outputs(4636)) and not (layer2_outputs(443));
    layer3_outputs(5575) <= not(layer2_outputs(1653));
    layer3_outputs(5576) <= not((layer2_outputs(1035)) and (layer2_outputs(925)));
    layer3_outputs(5577) <= not(layer2_outputs(65)) or (layer2_outputs(6396));
    layer3_outputs(5578) <= not((layer2_outputs(1767)) or (layer2_outputs(3272)));
    layer3_outputs(5579) <= not((layer2_outputs(2393)) xor (layer2_outputs(7293)));
    layer3_outputs(5580) <= layer2_outputs(4254);
    layer3_outputs(5581) <= not(layer2_outputs(488));
    layer3_outputs(5582) <= '1';
    layer3_outputs(5583) <= not(layer2_outputs(3308));
    layer3_outputs(5584) <= not(layer2_outputs(6896));
    layer3_outputs(5585) <= not(layer2_outputs(6949)) or (layer2_outputs(4979));
    layer3_outputs(5586) <= layer2_outputs(1603);
    layer3_outputs(5587) <= not(layer2_outputs(5996)) or (layer2_outputs(1107));
    layer3_outputs(5588) <= layer2_outputs(6475);
    layer3_outputs(5589) <= not(layer2_outputs(6045));
    layer3_outputs(5590) <= not((layer2_outputs(3960)) or (layer2_outputs(938)));
    layer3_outputs(5591) <= not((layer2_outputs(3404)) xor (layer2_outputs(3654)));
    layer3_outputs(5592) <= not(layer2_outputs(123));
    layer3_outputs(5593) <= not(layer2_outputs(3916)) or (layer2_outputs(5182));
    layer3_outputs(5594) <= (layer2_outputs(4241)) and not (layer2_outputs(1912));
    layer3_outputs(5595) <= not(layer2_outputs(4343)) or (layer2_outputs(6030));
    layer3_outputs(5596) <= not(layer2_outputs(6362));
    layer3_outputs(5597) <= not(layer2_outputs(3987));
    layer3_outputs(5598) <= (layer2_outputs(7326)) xor (layer2_outputs(7193));
    layer3_outputs(5599) <= (layer2_outputs(3106)) or (layer2_outputs(3412));
    layer3_outputs(5600) <= not(layer2_outputs(3401));
    layer3_outputs(5601) <= layer2_outputs(6141);
    layer3_outputs(5602) <= layer2_outputs(305);
    layer3_outputs(5603) <= not((layer2_outputs(4813)) and (layer2_outputs(2545)));
    layer3_outputs(5604) <= (layer2_outputs(5105)) and not (layer2_outputs(1390));
    layer3_outputs(5605) <= layer2_outputs(1474);
    layer3_outputs(5606) <= not(layer2_outputs(3156));
    layer3_outputs(5607) <= not(layer2_outputs(272)) or (layer2_outputs(409));
    layer3_outputs(5608) <= not(layer2_outputs(976));
    layer3_outputs(5609) <= (layer2_outputs(2)) xor (layer2_outputs(286));
    layer3_outputs(5610) <= layer2_outputs(4063);
    layer3_outputs(5611) <= not((layer2_outputs(2341)) or (layer2_outputs(2914)));
    layer3_outputs(5612) <= '0';
    layer3_outputs(5613) <= not(layer2_outputs(1397));
    layer3_outputs(5614) <= not(layer2_outputs(26));
    layer3_outputs(5615) <= not((layer2_outputs(1096)) xor (layer2_outputs(3537)));
    layer3_outputs(5616) <= layer2_outputs(3618);
    layer3_outputs(5617) <= not(layer2_outputs(4130)) or (layer2_outputs(1543));
    layer3_outputs(5618) <= (layer2_outputs(2615)) and not (layer2_outputs(1485));
    layer3_outputs(5619) <= not(layer2_outputs(6622));
    layer3_outputs(5620) <= layer2_outputs(185);
    layer3_outputs(5621) <= layer2_outputs(5618);
    layer3_outputs(5622) <= not(layer2_outputs(120));
    layer3_outputs(5623) <= layer2_outputs(6275);
    layer3_outputs(5624) <= not((layer2_outputs(3990)) xor (layer2_outputs(7598)));
    layer3_outputs(5625) <= layer2_outputs(5676);
    layer3_outputs(5626) <= (layer2_outputs(1900)) and (layer2_outputs(4672));
    layer3_outputs(5627) <= not(layer2_outputs(7038));
    layer3_outputs(5628) <= layer2_outputs(1666);
    layer3_outputs(5629) <= not(layer2_outputs(7378));
    layer3_outputs(5630) <= not(layer2_outputs(5351));
    layer3_outputs(5631) <= not(layer2_outputs(3434));
    layer3_outputs(5632) <= (layer2_outputs(4322)) or (layer2_outputs(2072));
    layer3_outputs(5633) <= not((layer2_outputs(5439)) or (layer2_outputs(2829)));
    layer3_outputs(5634) <= not(layer2_outputs(1728));
    layer3_outputs(5635) <= not((layer2_outputs(4472)) and (layer2_outputs(145)));
    layer3_outputs(5636) <= not((layer2_outputs(174)) or (layer2_outputs(1103)));
    layer3_outputs(5637) <= not((layer2_outputs(771)) and (layer2_outputs(1489)));
    layer3_outputs(5638) <= layer2_outputs(184);
    layer3_outputs(5639) <= layer2_outputs(3315);
    layer3_outputs(5640) <= not((layer2_outputs(3854)) and (layer2_outputs(1645)));
    layer3_outputs(5641) <= (layer2_outputs(1285)) and not (layer2_outputs(5401));
    layer3_outputs(5642) <= layer2_outputs(7363);
    layer3_outputs(5643) <= not(layer2_outputs(83));
    layer3_outputs(5644) <= (layer2_outputs(6545)) and not (layer2_outputs(4392));
    layer3_outputs(5645) <= (layer2_outputs(4028)) and not (layer2_outputs(622));
    layer3_outputs(5646) <= '1';
    layer3_outputs(5647) <= layer2_outputs(2079);
    layer3_outputs(5648) <= layer2_outputs(3232);
    layer3_outputs(5649) <= not((layer2_outputs(1338)) or (layer2_outputs(1246)));
    layer3_outputs(5650) <= not((layer2_outputs(4266)) and (layer2_outputs(3536)));
    layer3_outputs(5651) <= (layer2_outputs(633)) and not (layer2_outputs(7265));
    layer3_outputs(5652) <= (layer2_outputs(2792)) xor (layer2_outputs(5538));
    layer3_outputs(5653) <= not((layer2_outputs(6459)) and (layer2_outputs(3163)));
    layer3_outputs(5654) <= not(layer2_outputs(4005));
    layer3_outputs(5655) <= layer2_outputs(1051);
    layer3_outputs(5656) <= not(layer2_outputs(6822)) or (layer2_outputs(5462));
    layer3_outputs(5657) <= (layer2_outputs(893)) and not (layer2_outputs(5929));
    layer3_outputs(5658) <= layer2_outputs(5786);
    layer3_outputs(5659) <= not((layer2_outputs(3098)) and (layer2_outputs(4388)));
    layer3_outputs(5660) <= layer2_outputs(4782);
    layer3_outputs(5661) <= (layer2_outputs(1826)) and not (layer2_outputs(7257));
    layer3_outputs(5662) <= not((layer2_outputs(5935)) xor (layer2_outputs(2622)));
    layer3_outputs(5663) <= not(layer2_outputs(7071)) or (layer2_outputs(1128));
    layer3_outputs(5664) <= layer2_outputs(2715);
    layer3_outputs(5665) <= not((layer2_outputs(3643)) or (layer2_outputs(1850)));
    layer3_outputs(5666) <= not(layer2_outputs(382)) or (layer2_outputs(4663));
    layer3_outputs(5667) <= (layer2_outputs(3333)) or (layer2_outputs(3542));
    layer3_outputs(5668) <= '0';
    layer3_outputs(5669) <= (layer2_outputs(5631)) and (layer2_outputs(5767));
    layer3_outputs(5670) <= (layer2_outputs(3426)) xor (layer2_outputs(4276));
    layer3_outputs(5671) <= not(layer2_outputs(4477)) or (layer2_outputs(7646));
    layer3_outputs(5672) <= (layer2_outputs(6008)) and (layer2_outputs(3819));
    layer3_outputs(5673) <= (layer2_outputs(4968)) and (layer2_outputs(2840));
    layer3_outputs(5674) <= not(layer2_outputs(3339));
    layer3_outputs(5675) <= not(layer2_outputs(2684));
    layer3_outputs(5676) <= layer2_outputs(2636);
    layer3_outputs(5677) <= not(layer2_outputs(1458)) or (layer2_outputs(5503));
    layer3_outputs(5678) <= (layer2_outputs(3998)) and (layer2_outputs(567));
    layer3_outputs(5679) <= layer2_outputs(2944);
    layer3_outputs(5680) <= not((layer2_outputs(2524)) and (layer2_outputs(2362)));
    layer3_outputs(5681) <= not(layer2_outputs(73));
    layer3_outputs(5682) <= layer2_outputs(5726);
    layer3_outputs(5683) <= layer2_outputs(5027);
    layer3_outputs(5684) <= '0';
    layer3_outputs(5685) <= not(layer2_outputs(2684)) or (layer2_outputs(4959));
    layer3_outputs(5686) <= layer2_outputs(1909);
    layer3_outputs(5687) <= not(layer2_outputs(3734));
    layer3_outputs(5688) <= (layer2_outputs(4013)) and not (layer2_outputs(603));
    layer3_outputs(5689) <= (layer2_outputs(1896)) xor (layer2_outputs(4048));
    layer3_outputs(5690) <= (layer2_outputs(7272)) and not (layer2_outputs(757));
    layer3_outputs(5691) <= layer2_outputs(3646);
    layer3_outputs(5692) <= not(layer2_outputs(830));
    layer3_outputs(5693) <= (layer2_outputs(4618)) and not (layer2_outputs(6736));
    layer3_outputs(5694) <= not(layer2_outputs(2916));
    layer3_outputs(5695) <= layer2_outputs(5504);
    layer3_outputs(5696) <= (layer2_outputs(776)) and (layer2_outputs(4202));
    layer3_outputs(5697) <= not(layer2_outputs(1707)) or (layer2_outputs(6455));
    layer3_outputs(5698) <= layer2_outputs(2183);
    layer3_outputs(5699) <= not((layer2_outputs(4529)) or (layer2_outputs(2371)));
    layer3_outputs(5700) <= layer2_outputs(2494);
    layer3_outputs(5701) <= not(layer2_outputs(4970));
    layer3_outputs(5702) <= layer2_outputs(4508);
    layer3_outputs(5703) <= (layer2_outputs(2256)) and (layer2_outputs(5230));
    layer3_outputs(5704) <= layer2_outputs(2774);
    layer3_outputs(5705) <= layer2_outputs(1122);
    layer3_outputs(5706) <= not(layer2_outputs(7353)) or (layer2_outputs(2055));
    layer3_outputs(5707) <= not(layer2_outputs(1884));
    layer3_outputs(5708) <= layer2_outputs(6815);
    layer3_outputs(5709) <= not(layer2_outputs(1775));
    layer3_outputs(5710) <= not(layer2_outputs(3462));
    layer3_outputs(5711) <= not((layer2_outputs(4280)) or (layer2_outputs(6272)));
    layer3_outputs(5712) <= not((layer2_outputs(363)) xor (layer2_outputs(3148)));
    layer3_outputs(5713) <= (layer2_outputs(1789)) xor (layer2_outputs(7222));
    layer3_outputs(5714) <= not(layer2_outputs(6968)) or (layer2_outputs(3932));
    layer3_outputs(5715) <= (layer2_outputs(4349)) and not (layer2_outputs(2158));
    layer3_outputs(5716) <= layer2_outputs(604);
    layer3_outputs(5717) <= not((layer2_outputs(1366)) or (layer2_outputs(273)));
    layer3_outputs(5718) <= layer2_outputs(7483);
    layer3_outputs(5719) <= not(layer2_outputs(6775));
    layer3_outputs(5720) <= (layer2_outputs(5306)) or (layer2_outputs(3800));
    layer3_outputs(5721) <= '1';
    layer3_outputs(5722) <= not(layer2_outputs(1841));
    layer3_outputs(5723) <= '1';
    layer3_outputs(5724) <= (layer2_outputs(2613)) or (layer2_outputs(530));
    layer3_outputs(5725) <= (layer2_outputs(5924)) and (layer2_outputs(1633));
    layer3_outputs(5726) <= (layer2_outputs(3612)) and not (layer2_outputs(6343));
    layer3_outputs(5727) <= not(layer2_outputs(3314));
    layer3_outputs(5728) <= layer2_outputs(6193);
    layer3_outputs(5729) <= not(layer2_outputs(6280));
    layer3_outputs(5730) <= not((layer2_outputs(658)) or (layer2_outputs(5078)));
    layer3_outputs(5731) <= not((layer2_outputs(4499)) or (layer2_outputs(1154)));
    layer3_outputs(5732) <= not((layer2_outputs(203)) or (layer2_outputs(3928)));
    layer3_outputs(5733) <= layer2_outputs(7115);
    layer3_outputs(5734) <= (layer2_outputs(461)) xor (layer2_outputs(4553));
    layer3_outputs(5735) <= (layer2_outputs(63)) and not (layer2_outputs(4620));
    layer3_outputs(5736) <= layer2_outputs(494);
    layer3_outputs(5737) <= layer2_outputs(1984);
    layer3_outputs(5738) <= not((layer2_outputs(6568)) and (layer2_outputs(2516)));
    layer3_outputs(5739) <= (layer2_outputs(2076)) or (layer2_outputs(5388));
    layer3_outputs(5740) <= (layer2_outputs(3495)) xor (layer2_outputs(2662));
    layer3_outputs(5741) <= not(layer2_outputs(5908));
    layer3_outputs(5742) <= (layer2_outputs(7158)) and not (layer2_outputs(4533));
    layer3_outputs(5743) <= (layer2_outputs(6376)) and not (layer2_outputs(4927));
    layer3_outputs(5744) <= (layer2_outputs(4724)) or (layer2_outputs(1272));
    layer3_outputs(5745) <= (layer2_outputs(3624)) or (layer2_outputs(1447));
    layer3_outputs(5746) <= (layer2_outputs(3194)) xor (layer2_outputs(7069));
    layer3_outputs(5747) <= layer2_outputs(5871);
    layer3_outputs(5748) <= not(layer2_outputs(6424));
    layer3_outputs(5749) <= not((layer2_outputs(6967)) or (layer2_outputs(6406)));
    layer3_outputs(5750) <= not(layer2_outputs(4873));
    layer3_outputs(5751) <= not(layer2_outputs(4987));
    layer3_outputs(5752) <= not(layer2_outputs(6387)) or (layer2_outputs(1343));
    layer3_outputs(5753) <= (layer2_outputs(2075)) or (layer2_outputs(2865));
    layer3_outputs(5754) <= not((layer2_outputs(1636)) xor (layer2_outputs(3235)));
    layer3_outputs(5755) <= not(layer2_outputs(387));
    layer3_outputs(5756) <= (layer2_outputs(4763)) and not (layer2_outputs(278));
    layer3_outputs(5757) <= not(layer2_outputs(6800)) or (layer2_outputs(4249));
    layer3_outputs(5758) <= (layer2_outputs(1524)) and not (layer2_outputs(3398));
    layer3_outputs(5759) <= not(layer2_outputs(7467));
    layer3_outputs(5760) <= not(layer2_outputs(344));
    layer3_outputs(5761) <= not(layer2_outputs(5550)) or (layer2_outputs(5054));
    layer3_outputs(5762) <= layer2_outputs(4450);
    layer3_outputs(5763) <= not(layer2_outputs(2984));
    layer3_outputs(5764) <= layer2_outputs(2655);
    layer3_outputs(5765) <= layer2_outputs(3963);
    layer3_outputs(5766) <= layer2_outputs(122);
    layer3_outputs(5767) <= not(layer2_outputs(2051));
    layer3_outputs(5768) <= (layer2_outputs(6796)) and not (layer2_outputs(3558));
    layer3_outputs(5769) <= layer2_outputs(5726);
    layer3_outputs(5770) <= not((layer2_outputs(1317)) or (layer2_outputs(6816)));
    layer3_outputs(5771) <= (layer2_outputs(2598)) or (layer2_outputs(870));
    layer3_outputs(5772) <= layer2_outputs(6490);
    layer3_outputs(5773) <= (layer2_outputs(5511)) or (layer2_outputs(4384));
    layer3_outputs(5774) <= (layer2_outputs(7316)) xor (layer2_outputs(2002));
    layer3_outputs(5775) <= layer2_outputs(4245);
    layer3_outputs(5776) <= (layer2_outputs(3703)) or (layer2_outputs(3197));
    layer3_outputs(5777) <= not(layer2_outputs(4801));
    layer3_outputs(5778) <= (layer2_outputs(1857)) and not (layer2_outputs(3603));
    layer3_outputs(5779) <= '0';
    layer3_outputs(5780) <= layer2_outputs(993);
    layer3_outputs(5781) <= not(layer2_outputs(1250));
    layer3_outputs(5782) <= not((layer2_outputs(4627)) or (layer2_outputs(2666)));
    layer3_outputs(5783) <= not((layer2_outputs(2176)) or (layer2_outputs(3211)));
    layer3_outputs(5784) <= not(layer2_outputs(2858));
    layer3_outputs(5785) <= layer2_outputs(3996);
    layer3_outputs(5786) <= (layer2_outputs(4956)) xor (layer2_outputs(978));
    layer3_outputs(5787) <= layer2_outputs(4803);
    layer3_outputs(5788) <= not(layer2_outputs(5344));
    layer3_outputs(5789) <= not(layer2_outputs(2517));
    layer3_outputs(5790) <= (layer2_outputs(442)) and not (layer2_outputs(5407));
    layer3_outputs(5791) <= (layer2_outputs(477)) and not (layer2_outputs(12));
    layer3_outputs(5792) <= not(layer2_outputs(1340));
    layer3_outputs(5793) <= layer2_outputs(4038);
    layer3_outputs(5794) <= not(layer2_outputs(1972)) or (layer2_outputs(1263));
    layer3_outputs(5795) <= '1';
    layer3_outputs(5796) <= not((layer2_outputs(161)) and (layer2_outputs(3634)));
    layer3_outputs(5797) <= not(layer2_outputs(5149));
    layer3_outputs(5798) <= not(layer2_outputs(4079)) or (layer2_outputs(2312));
    layer3_outputs(5799) <= '0';
    layer3_outputs(5800) <= layer2_outputs(1301);
    layer3_outputs(5801) <= layer2_outputs(1599);
    layer3_outputs(5802) <= not((layer2_outputs(4285)) or (layer2_outputs(1478)));
    layer3_outputs(5803) <= not(layer2_outputs(982)) or (layer2_outputs(4306));
    layer3_outputs(5804) <= not(layer2_outputs(846)) or (layer2_outputs(2615));
    layer3_outputs(5805) <= not(layer2_outputs(2123));
    layer3_outputs(5806) <= not(layer2_outputs(462));
    layer3_outputs(5807) <= not(layer2_outputs(1958));
    layer3_outputs(5808) <= not(layer2_outputs(2522)) or (layer2_outputs(5196));
    layer3_outputs(5809) <= (layer2_outputs(248)) and (layer2_outputs(3384));
    layer3_outputs(5810) <= not(layer2_outputs(2195)) or (layer2_outputs(4522));
    layer3_outputs(5811) <= not((layer2_outputs(928)) or (layer2_outputs(5891)));
    layer3_outputs(5812) <= not(layer2_outputs(4045)) or (layer2_outputs(1736));
    layer3_outputs(5813) <= layer2_outputs(254);
    layer3_outputs(5814) <= layer2_outputs(2051);
    layer3_outputs(5815) <= layer2_outputs(5594);
    layer3_outputs(5816) <= layer2_outputs(2052);
    layer3_outputs(5817) <= layer2_outputs(2672);
    layer3_outputs(5818) <= '1';
    layer3_outputs(5819) <= (layer2_outputs(5265)) and not (layer2_outputs(3973));
    layer3_outputs(5820) <= not((layer2_outputs(3107)) and (layer2_outputs(1589)));
    layer3_outputs(5821) <= not(layer2_outputs(1886)) or (layer2_outputs(2923));
    layer3_outputs(5822) <= (layer2_outputs(6176)) and (layer2_outputs(7371));
    layer3_outputs(5823) <= (layer2_outputs(4852)) and (layer2_outputs(954));
    layer3_outputs(5824) <= not(layer2_outputs(5046));
    layer3_outputs(5825) <= not(layer2_outputs(2665));
    layer3_outputs(5826) <= (layer2_outputs(994)) and not (layer2_outputs(5171));
    layer3_outputs(5827) <= not(layer2_outputs(516)) or (layer2_outputs(4421));
    layer3_outputs(5828) <= (layer2_outputs(165)) and (layer2_outputs(3897));
    layer3_outputs(5829) <= '0';
    layer3_outputs(5830) <= (layer2_outputs(4564)) xor (layer2_outputs(4049));
    layer3_outputs(5831) <= not(layer2_outputs(2892)) or (layer2_outputs(421));
    layer3_outputs(5832) <= layer2_outputs(138);
    layer3_outputs(5833) <= not(layer2_outputs(3735)) or (layer2_outputs(4076));
    layer3_outputs(5834) <= (layer2_outputs(1268)) and not (layer2_outputs(3246));
    layer3_outputs(5835) <= (layer2_outputs(4621)) or (layer2_outputs(4162));
    layer3_outputs(5836) <= not(layer2_outputs(2863));
    layer3_outputs(5837) <= not(layer2_outputs(1916)) or (layer2_outputs(1862));
    layer3_outputs(5838) <= not(layer2_outputs(3967));
    layer3_outputs(5839) <= (layer2_outputs(4858)) xor (layer2_outputs(6243));
    layer3_outputs(5840) <= (layer2_outputs(5730)) xor (layer2_outputs(5545));
    layer3_outputs(5841) <= not(layer2_outputs(6969));
    layer3_outputs(5842) <= not(layer2_outputs(995)) or (layer2_outputs(7277));
    layer3_outputs(5843) <= not(layer2_outputs(2961));
    layer3_outputs(5844) <= not(layer2_outputs(2221));
    layer3_outputs(5845) <= not((layer2_outputs(7502)) or (layer2_outputs(795)));
    layer3_outputs(5846) <= '1';
    layer3_outputs(5847) <= not(layer2_outputs(3528));
    layer3_outputs(5848) <= layer2_outputs(4882);
    layer3_outputs(5849) <= not(layer2_outputs(1744)) or (layer2_outputs(5473));
    layer3_outputs(5850) <= '1';
    layer3_outputs(5851) <= not((layer2_outputs(1359)) and (layer2_outputs(5939)));
    layer3_outputs(5852) <= '0';
    layer3_outputs(5853) <= layer2_outputs(5336);
    layer3_outputs(5854) <= not((layer2_outputs(7344)) or (layer2_outputs(6057)));
    layer3_outputs(5855) <= (layer2_outputs(3459)) and not (layer2_outputs(5687));
    layer3_outputs(5856) <= (layer2_outputs(3114)) and not (layer2_outputs(863));
    layer3_outputs(5857) <= (layer2_outputs(2688)) xor (layer2_outputs(7381));
    layer3_outputs(5858) <= not(layer2_outputs(649)) or (layer2_outputs(2069));
    layer3_outputs(5859) <= layer2_outputs(2832);
    layer3_outputs(5860) <= not((layer2_outputs(1792)) or (layer2_outputs(2617)));
    layer3_outputs(5861) <= not((layer2_outputs(3083)) or (layer2_outputs(1525)));
    layer3_outputs(5862) <= (layer2_outputs(5558)) or (layer2_outputs(1472));
    layer3_outputs(5863) <= layer2_outputs(941);
    layer3_outputs(5864) <= layer2_outputs(4785);
    layer3_outputs(5865) <= layer2_outputs(2841);
    layer3_outputs(5866) <= (layer2_outputs(4983)) and not (layer2_outputs(5229));
    layer3_outputs(5867) <= (layer2_outputs(6794)) and (layer2_outputs(3573));
    layer3_outputs(5868) <= not(layer2_outputs(1484));
    layer3_outputs(5869) <= (layer2_outputs(3153)) and not (layer2_outputs(517));
    layer3_outputs(5870) <= not(layer2_outputs(2013));
    layer3_outputs(5871) <= not(layer2_outputs(3834));
    layer3_outputs(5872) <= (layer2_outputs(1322)) and not (layer2_outputs(4428));
    layer3_outputs(5873) <= not(layer2_outputs(7393)) or (layer2_outputs(3985));
    layer3_outputs(5874) <= layer2_outputs(191);
    layer3_outputs(5875) <= not((layer2_outputs(7318)) and (layer2_outputs(2985)));
    layer3_outputs(5876) <= not((layer2_outputs(4329)) or (layer2_outputs(462)));
    layer3_outputs(5877) <= not(layer2_outputs(4573)) or (layer2_outputs(2331));
    layer3_outputs(5878) <= layer2_outputs(578);
    layer3_outputs(5879) <= layer2_outputs(2703);
    layer3_outputs(5880) <= not(layer2_outputs(568));
    layer3_outputs(5881) <= (layer2_outputs(4064)) and (layer2_outputs(5510));
    layer3_outputs(5882) <= not(layer2_outputs(2909)) or (layer2_outputs(6415));
    layer3_outputs(5883) <= layer2_outputs(5178);
    layer3_outputs(5884) <= not(layer2_outputs(1003));
    layer3_outputs(5885) <= not(layer2_outputs(1074)) or (layer2_outputs(6971));
    layer3_outputs(5886) <= not((layer2_outputs(494)) or (layer2_outputs(1737)));
    layer3_outputs(5887) <= not(layer2_outputs(3005));
    layer3_outputs(5888) <= layer2_outputs(3570);
    layer3_outputs(5889) <= not((layer2_outputs(5195)) or (layer2_outputs(4404)));
    layer3_outputs(5890) <= (layer2_outputs(4093)) or (layer2_outputs(7679));
    layer3_outputs(5891) <= (layer2_outputs(5260)) and not (layer2_outputs(6474));
    layer3_outputs(5892) <= (layer2_outputs(7220)) xor (layer2_outputs(1017));
    layer3_outputs(5893) <= (layer2_outputs(6535)) and (layer2_outputs(3169));
    layer3_outputs(5894) <= (layer2_outputs(4710)) xor (layer2_outputs(6885));
    layer3_outputs(5895) <= (layer2_outputs(6260)) and not (layer2_outputs(3139));
    layer3_outputs(5896) <= layer2_outputs(3130);
    layer3_outputs(5897) <= not(layer2_outputs(6185)) or (layer2_outputs(4903));
    layer3_outputs(5898) <= layer2_outputs(386);
    layer3_outputs(5899) <= not(layer2_outputs(0));
    layer3_outputs(5900) <= layer2_outputs(6821);
    layer3_outputs(5901) <= (layer2_outputs(4188)) and (layer2_outputs(3261));
    layer3_outputs(5902) <= (layer2_outputs(932)) or (layer2_outputs(3204));
    layer3_outputs(5903) <= not(layer2_outputs(4474));
    layer3_outputs(5904) <= not(layer2_outputs(3467));
    layer3_outputs(5905) <= not(layer2_outputs(816)) or (layer2_outputs(4858));
    layer3_outputs(5906) <= (layer2_outputs(3788)) and (layer2_outputs(1940));
    layer3_outputs(5907) <= layer2_outputs(3020);
    layer3_outputs(5908) <= not(layer2_outputs(4061)) or (layer2_outputs(4606));
    layer3_outputs(5909) <= not(layer2_outputs(3598));
    layer3_outputs(5910) <= (layer2_outputs(323)) and not (layer2_outputs(99));
    layer3_outputs(5911) <= not(layer2_outputs(1166));
    layer3_outputs(5912) <= not((layer2_outputs(1206)) or (layer2_outputs(4901)));
    layer3_outputs(5913) <= not((layer2_outputs(1088)) or (layer2_outputs(1119)));
    layer3_outputs(5914) <= (layer2_outputs(4782)) or (layer2_outputs(1806));
    layer3_outputs(5915) <= (layer2_outputs(5938)) and not (layer2_outputs(5004));
    layer3_outputs(5916) <= (layer2_outputs(7660)) xor (layer2_outputs(3832));
    layer3_outputs(5917) <= (layer2_outputs(98)) and not (layer2_outputs(5498));
    layer3_outputs(5918) <= '1';
    layer3_outputs(5919) <= (layer2_outputs(6654)) and not (layer2_outputs(6586));
    layer3_outputs(5920) <= layer2_outputs(4634);
    layer3_outputs(5921) <= layer2_outputs(441);
    layer3_outputs(5922) <= (layer2_outputs(1970)) and not (layer2_outputs(2920));
    layer3_outputs(5923) <= layer2_outputs(5049);
    layer3_outputs(5924) <= not(layer2_outputs(2199));
    layer3_outputs(5925) <= layer2_outputs(6290);
    layer3_outputs(5926) <= layer2_outputs(5021);
    layer3_outputs(5927) <= (layer2_outputs(3080)) and (layer2_outputs(5785));
    layer3_outputs(5928) <= (layer2_outputs(1323)) and (layer2_outputs(439));
    layer3_outputs(5929) <= (layer2_outputs(4983)) and not (layer2_outputs(3948));
    layer3_outputs(5930) <= not((layer2_outputs(4402)) or (layer2_outputs(2631)));
    layer3_outputs(5931) <= not(layer2_outputs(977)) or (layer2_outputs(1616));
    layer3_outputs(5932) <= not(layer2_outputs(6384));
    layer3_outputs(5933) <= not(layer2_outputs(6849)) or (layer2_outputs(1238));
    layer3_outputs(5934) <= layer2_outputs(3576);
    layer3_outputs(5935) <= not(layer2_outputs(212));
    layer3_outputs(5936) <= '0';
    layer3_outputs(5937) <= layer2_outputs(2630);
    layer3_outputs(5938) <= (layer2_outputs(7667)) and not (layer2_outputs(3328));
    layer3_outputs(5939) <= (layer2_outputs(3965)) and (layer2_outputs(2341));
    layer3_outputs(5940) <= not(layer2_outputs(5606)) or (layer2_outputs(6013));
    layer3_outputs(5941) <= not(layer2_outputs(7350)) or (layer2_outputs(5525));
    layer3_outputs(5942) <= not(layer2_outputs(6288));
    layer3_outputs(5943) <= not((layer2_outputs(6293)) and (layer2_outputs(6995)));
    layer3_outputs(5944) <= not(layer2_outputs(7098));
    layer3_outputs(5945) <= (layer2_outputs(7373)) and not (layer2_outputs(5029));
    layer3_outputs(5946) <= not((layer2_outputs(6220)) or (layer2_outputs(6063)));
    layer3_outputs(5947) <= '0';
    layer3_outputs(5948) <= layer2_outputs(701);
    layer3_outputs(5949) <= not(layer2_outputs(3177));
    layer3_outputs(5950) <= not(layer2_outputs(7113));
    layer3_outputs(5951) <= not((layer2_outputs(1010)) or (layer2_outputs(6792)));
    layer3_outputs(5952) <= not(layer2_outputs(3402));
    layer3_outputs(5953) <= not(layer2_outputs(3540)) or (layer2_outputs(2511));
    layer3_outputs(5954) <= '1';
    layer3_outputs(5955) <= (layer2_outputs(5295)) and not (layer2_outputs(4022));
    layer3_outputs(5956) <= layer2_outputs(4847);
    layer3_outputs(5957) <= not((layer2_outputs(7621)) and (layer2_outputs(263)));
    layer3_outputs(5958) <= layer2_outputs(3683);
    layer3_outputs(5959) <= layer2_outputs(7071);
    layer3_outputs(5960) <= not(layer2_outputs(6330));
    layer3_outputs(5961) <= layer2_outputs(534);
    layer3_outputs(5962) <= layer2_outputs(5890);
    layer3_outputs(5963) <= (layer2_outputs(1152)) and (layer2_outputs(6837));
    layer3_outputs(5964) <= layer2_outputs(4230);
    layer3_outputs(5965) <= not(layer2_outputs(6037)) or (layer2_outputs(1289));
    layer3_outputs(5966) <= not((layer2_outputs(2070)) and (layer2_outputs(3390)));
    layer3_outputs(5967) <= not((layer2_outputs(3267)) xor (layer2_outputs(4571)));
    layer3_outputs(5968) <= layer2_outputs(78);
    layer3_outputs(5969) <= not(layer2_outputs(5182));
    layer3_outputs(5970) <= layer2_outputs(3323);
    layer3_outputs(5971) <= not((layer2_outputs(5901)) or (layer2_outputs(2241)));
    layer3_outputs(5972) <= (layer2_outputs(6990)) and (layer2_outputs(4713));
    layer3_outputs(5973) <= not(layer2_outputs(4624));
    layer3_outputs(5974) <= not(layer2_outputs(4163)) or (layer2_outputs(6203));
    layer3_outputs(5975) <= layer2_outputs(4316);
    layer3_outputs(5976) <= not(layer2_outputs(624));
    layer3_outputs(5977) <= (layer2_outputs(2678)) and (layer2_outputs(6826));
    layer3_outputs(5978) <= not(layer2_outputs(4588)) or (layer2_outputs(1071));
    layer3_outputs(5979) <= (layer2_outputs(3693)) and (layer2_outputs(4507));
    layer3_outputs(5980) <= not((layer2_outputs(2765)) and (layer2_outputs(560)));
    layer3_outputs(5981) <= not(layer2_outputs(5934)) or (layer2_outputs(3114));
    layer3_outputs(5982) <= layer2_outputs(5712);
    layer3_outputs(5983) <= (layer2_outputs(6146)) and not (layer2_outputs(3975));
    layer3_outputs(5984) <= not(layer2_outputs(5562)) or (layer2_outputs(860));
    layer3_outputs(5985) <= (layer2_outputs(6657)) or (layer2_outputs(6213));
    layer3_outputs(5986) <= not(layer2_outputs(4946));
    layer3_outputs(5987) <= (layer2_outputs(330)) and not (layer2_outputs(4696));
    layer3_outputs(5988) <= layer2_outputs(436);
    layer3_outputs(5989) <= layer2_outputs(2259);
    layer3_outputs(5990) <= (layer2_outputs(5602)) and not (layer2_outputs(5521));
    layer3_outputs(5991) <= not(layer2_outputs(3971)) or (layer2_outputs(1000));
    layer3_outputs(5992) <= not(layer2_outputs(4569)) or (layer2_outputs(2187));
    layer3_outputs(5993) <= not(layer2_outputs(5207)) or (layer2_outputs(1952));
    layer3_outputs(5994) <= (layer2_outputs(590)) and not (layer2_outputs(1233));
    layer3_outputs(5995) <= not(layer2_outputs(374));
    layer3_outputs(5996) <= (layer2_outputs(6021)) and (layer2_outputs(6819));
    layer3_outputs(5997) <= not(layer2_outputs(3037));
    layer3_outputs(5998) <= (layer2_outputs(5565)) or (layer2_outputs(465));
    layer3_outputs(5999) <= not(layer2_outputs(5104)) or (layer2_outputs(3714));
    layer3_outputs(6000) <= not(layer2_outputs(925)) or (layer2_outputs(3899));
    layer3_outputs(6001) <= layer2_outputs(372);
    layer3_outputs(6002) <= (layer2_outputs(2416)) and (layer2_outputs(7371));
    layer3_outputs(6003) <= (layer2_outputs(5372)) and not (layer2_outputs(4329));
    layer3_outputs(6004) <= (layer2_outputs(227)) and not (layer2_outputs(6245));
    layer3_outputs(6005) <= not(layer2_outputs(7380)) or (layer2_outputs(260));
    layer3_outputs(6006) <= layer2_outputs(978);
    layer3_outputs(6007) <= not((layer2_outputs(1166)) or (layer2_outputs(2460)));
    layer3_outputs(6008) <= not((layer2_outputs(5493)) or (layer2_outputs(2355)));
    layer3_outputs(6009) <= not(layer2_outputs(5259));
    layer3_outputs(6010) <= (layer2_outputs(4170)) and not (layer2_outputs(2095));
    layer3_outputs(6011) <= (layer2_outputs(1079)) and (layer2_outputs(2547));
    layer3_outputs(6012) <= not(layer2_outputs(4495)) or (layer2_outputs(5100));
    layer3_outputs(6013) <= (layer2_outputs(5208)) or (layer2_outputs(4351));
    layer3_outputs(6014) <= (layer2_outputs(1811)) and not (layer2_outputs(2212));
    layer3_outputs(6015) <= layer2_outputs(5711);
    layer3_outputs(6016) <= (layer2_outputs(725)) and (layer2_outputs(2645));
    layer3_outputs(6017) <= not(layer2_outputs(1443));
    layer3_outputs(6018) <= not((layer2_outputs(3674)) and (layer2_outputs(5902)));
    layer3_outputs(6019) <= layer2_outputs(5577);
    layer3_outputs(6020) <= (layer2_outputs(4950)) xor (layer2_outputs(7458));
    layer3_outputs(6021) <= not(layer2_outputs(1679));
    layer3_outputs(6022) <= (layer2_outputs(1447)) and not (layer2_outputs(5826));
    layer3_outputs(6023) <= layer2_outputs(6670);
    layer3_outputs(6024) <= not((layer2_outputs(3146)) or (layer2_outputs(5268)));
    layer3_outputs(6025) <= not(layer2_outputs(2566));
    layer3_outputs(6026) <= not((layer2_outputs(2184)) xor (layer2_outputs(3447)));
    layer3_outputs(6027) <= layer2_outputs(3539);
    layer3_outputs(6028) <= (layer2_outputs(1325)) or (layer2_outputs(6035));
    layer3_outputs(6029) <= (layer2_outputs(5415)) and not (layer2_outputs(1299));
    layer3_outputs(6030) <= not(layer2_outputs(1223));
    layer3_outputs(6031) <= (layer2_outputs(4190)) and (layer2_outputs(3827));
    layer3_outputs(6032) <= layer2_outputs(5725);
    layer3_outputs(6033) <= not((layer2_outputs(7661)) or (layer2_outputs(4536)));
    layer3_outputs(6034) <= layer2_outputs(5651);
    layer3_outputs(6035) <= (layer2_outputs(5200)) and not (layer2_outputs(6595));
    layer3_outputs(6036) <= not((layer2_outputs(7398)) and (layer2_outputs(1372)));
    layer3_outputs(6037) <= not(layer2_outputs(3909));
    layer3_outputs(6038) <= not((layer2_outputs(6883)) and (layer2_outputs(1522)));
    layer3_outputs(6039) <= not(layer2_outputs(3304));
    layer3_outputs(6040) <= (layer2_outputs(4489)) xor (layer2_outputs(4869));
    layer3_outputs(6041) <= not(layer2_outputs(1973));
    layer3_outputs(6042) <= (layer2_outputs(3481)) and (layer2_outputs(1196));
    layer3_outputs(6043) <= layer2_outputs(8);
    layer3_outputs(6044) <= layer2_outputs(1435);
    layer3_outputs(6045) <= not(layer2_outputs(4745));
    layer3_outputs(6046) <= not(layer2_outputs(2956));
    layer3_outputs(6047) <= (layer2_outputs(3405)) xor (layer2_outputs(3749));
    layer3_outputs(6048) <= not((layer2_outputs(6698)) xor (layer2_outputs(2417)));
    layer3_outputs(6049) <= not((layer2_outputs(1541)) and (layer2_outputs(4439)));
    layer3_outputs(6050) <= not(layer2_outputs(4185)) or (layer2_outputs(3546));
    layer3_outputs(6051) <= not((layer2_outputs(794)) or (layer2_outputs(2150)));
    layer3_outputs(6052) <= layer2_outputs(3974);
    layer3_outputs(6053) <= (layer2_outputs(3079)) xor (layer2_outputs(4548));
    layer3_outputs(6054) <= not(layer2_outputs(2076));
    layer3_outputs(6055) <= (layer2_outputs(3448)) and (layer2_outputs(5851));
    layer3_outputs(6056) <= layer2_outputs(2563);
    layer3_outputs(6057) <= (layer2_outputs(4336)) and (layer2_outputs(3543));
    layer3_outputs(6058) <= layer2_outputs(3407);
    layer3_outputs(6059) <= '1';
    layer3_outputs(6060) <= layer2_outputs(5788);
    layer3_outputs(6061) <= not((layer2_outputs(4689)) and (layer2_outputs(1783)));
    layer3_outputs(6062) <= layer2_outputs(5781);
    layer3_outputs(6063) <= (layer2_outputs(4065)) and not (layer2_outputs(5030));
    layer3_outputs(6064) <= not((layer2_outputs(3000)) xor (layer2_outputs(1032)));
    layer3_outputs(6065) <= not(layer2_outputs(277));
    layer3_outputs(6066) <= not(layer2_outputs(4274));
    layer3_outputs(6067) <= not(layer2_outputs(1369));
    layer3_outputs(6068) <= not(layer2_outputs(336));
    layer3_outputs(6069) <= not((layer2_outputs(129)) and (layer2_outputs(1107)));
    layer3_outputs(6070) <= (layer2_outputs(5212)) or (layer2_outputs(2024));
    layer3_outputs(6071) <= (layer2_outputs(500)) and not (layer2_outputs(6354));
    layer3_outputs(6072) <= layer2_outputs(5579);
    layer3_outputs(6073) <= layer2_outputs(1024);
    layer3_outputs(6074) <= not((layer2_outputs(101)) or (layer2_outputs(6688)));
    layer3_outputs(6075) <= (layer2_outputs(1452)) and not (layer2_outputs(6639));
    layer3_outputs(6076) <= not(layer2_outputs(508));
    layer3_outputs(6077) <= not(layer2_outputs(5162));
    layer3_outputs(6078) <= (layer2_outputs(4448)) xor (layer2_outputs(2420));
    layer3_outputs(6079) <= (layer2_outputs(1639)) and not (layer2_outputs(5980));
    layer3_outputs(6080) <= not((layer2_outputs(1867)) xor (layer2_outputs(1859)));
    layer3_outputs(6081) <= not(layer2_outputs(1580));
    layer3_outputs(6082) <= (layer2_outputs(772)) and not (layer2_outputs(7303));
    layer3_outputs(6083) <= layer2_outputs(1057);
    layer3_outputs(6084) <= layer2_outputs(1033);
    layer3_outputs(6085) <= not(layer2_outputs(398)) or (layer2_outputs(3509));
    layer3_outputs(6086) <= layer2_outputs(3234);
    layer3_outputs(6087) <= '1';
    layer3_outputs(6088) <= not((layer2_outputs(7141)) or (layer2_outputs(3870)));
    layer3_outputs(6089) <= not(layer2_outputs(7192));
    layer3_outputs(6090) <= layer2_outputs(4401);
    layer3_outputs(6091) <= not(layer2_outputs(2901));
    layer3_outputs(6092) <= not(layer2_outputs(2412)) or (layer2_outputs(5281));
    layer3_outputs(6093) <= not((layer2_outputs(5414)) or (layer2_outputs(3380)));
    layer3_outputs(6094) <= not(layer2_outputs(1178));
    layer3_outputs(6095) <= not(layer2_outputs(156));
    layer3_outputs(6096) <= (layer2_outputs(4484)) or (layer2_outputs(2394));
    layer3_outputs(6097) <= (layer2_outputs(2083)) or (layer2_outputs(6138));
    layer3_outputs(6098) <= (layer2_outputs(4973)) and not (layer2_outputs(6773));
    layer3_outputs(6099) <= not(layer2_outputs(6782));
    layer3_outputs(6100) <= layer2_outputs(4867);
    layer3_outputs(6101) <= (layer2_outputs(3449)) or (layer2_outputs(3734));
    layer3_outputs(6102) <= layer2_outputs(7083);
    layer3_outputs(6103) <= (layer2_outputs(6119)) and not (layer2_outputs(3413));
    layer3_outputs(6104) <= not(layer2_outputs(5737)) or (layer2_outputs(2346));
    layer3_outputs(6105) <= not(layer2_outputs(3955)) or (layer2_outputs(4002));
    layer3_outputs(6106) <= '0';
    layer3_outputs(6107) <= not(layer2_outputs(1784)) or (layer2_outputs(1377));
    layer3_outputs(6108) <= not((layer2_outputs(5619)) and (layer2_outputs(6350)));
    layer3_outputs(6109) <= layer2_outputs(3809);
    layer3_outputs(6110) <= not(layer2_outputs(5399));
    layer3_outputs(6111) <= not(layer2_outputs(6304));
    layer3_outputs(6112) <= not(layer2_outputs(6603));
    layer3_outputs(6113) <= not(layer2_outputs(5009));
    layer3_outputs(6114) <= (layer2_outputs(2871)) or (layer2_outputs(6181));
    layer3_outputs(6115) <= layer2_outputs(5755);
    layer3_outputs(6116) <= layer2_outputs(3596);
    layer3_outputs(6117) <= not((layer2_outputs(3663)) and (layer2_outputs(5747)));
    layer3_outputs(6118) <= '1';
    layer3_outputs(6119) <= layer2_outputs(247);
    layer3_outputs(6120) <= layer2_outputs(7027);
    layer3_outputs(6121) <= layer2_outputs(6304);
    layer3_outputs(6122) <= (layer2_outputs(1297)) and not (layer2_outputs(349));
    layer3_outputs(6123) <= not(layer2_outputs(5088));
    layer3_outputs(6124) <= not(layer2_outputs(5089)) or (layer2_outputs(6134));
    layer3_outputs(6125) <= not(layer2_outputs(6633));
    layer3_outputs(6126) <= layer2_outputs(4845);
    layer3_outputs(6127) <= (layer2_outputs(3453)) and not (layer2_outputs(3335));
    layer3_outputs(6128) <= '0';
    layer3_outputs(6129) <= layer2_outputs(6660);
    layer3_outputs(6130) <= (layer2_outputs(2000)) and (layer2_outputs(3560));
    layer3_outputs(6131) <= layer2_outputs(4972);
    layer3_outputs(6132) <= not((layer2_outputs(3582)) and (layer2_outputs(1857)));
    layer3_outputs(6133) <= layer2_outputs(4348);
    layer3_outputs(6134) <= not(layer2_outputs(4718)) or (layer2_outputs(614));
    layer3_outputs(6135) <= layer2_outputs(5481);
    layer3_outputs(6136) <= not(layer2_outputs(186)) or (layer2_outputs(6510));
    layer3_outputs(6137) <= (layer2_outputs(3066)) or (layer2_outputs(2032));
    layer3_outputs(6138) <= not(layer2_outputs(5361));
    layer3_outputs(6139) <= not((layer2_outputs(573)) or (layer2_outputs(3167)));
    layer3_outputs(6140) <= not((layer2_outputs(2976)) or (layer2_outputs(2879)));
    layer3_outputs(6141) <= not(layer2_outputs(691));
    layer3_outputs(6142) <= not(layer2_outputs(5896));
    layer3_outputs(6143) <= layer2_outputs(3919);
    layer3_outputs(6144) <= not(layer2_outputs(7252));
    layer3_outputs(6145) <= not(layer2_outputs(743));
    layer3_outputs(6146) <= layer2_outputs(714);
    layer3_outputs(6147) <= not(layer2_outputs(4108));
    layer3_outputs(6148) <= layer2_outputs(5825);
    layer3_outputs(6149) <= (layer2_outputs(5333)) xor (layer2_outputs(1812));
    layer3_outputs(6150) <= not(layer2_outputs(6695));
    layer3_outputs(6151) <= (layer2_outputs(315)) and (layer2_outputs(5125));
    layer3_outputs(6152) <= not(layer2_outputs(3579));
    layer3_outputs(6153) <= layer2_outputs(4105);
    layer3_outputs(6154) <= layer2_outputs(2335);
    layer3_outputs(6155) <= layer2_outputs(5242);
    layer3_outputs(6156) <= not(layer2_outputs(5795)) or (layer2_outputs(4582));
    layer3_outputs(6157) <= layer2_outputs(2605);
    layer3_outputs(6158) <= layer2_outputs(2580);
    layer3_outputs(6159) <= layer2_outputs(4667);
    layer3_outputs(6160) <= not(layer2_outputs(635));
    layer3_outputs(6161) <= layer2_outputs(618);
    layer3_outputs(6162) <= not(layer2_outputs(5283));
    layer3_outputs(6163) <= (layer2_outputs(3054)) or (layer2_outputs(4086));
    layer3_outputs(6164) <= layer2_outputs(1001);
    layer3_outputs(6165) <= layer2_outputs(6662);
    layer3_outputs(6166) <= (layer2_outputs(1067)) and (layer2_outputs(3400));
    layer3_outputs(6167) <= layer2_outputs(327);
    layer3_outputs(6168) <= layer2_outputs(525);
    layer3_outputs(6169) <= not(layer2_outputs(1790));
    layer3_outputs(6170) <= (layer2_outputs(5100)) and (layer2_outputs(7532));
    layer3_outputs(6171) <= not((layer2_outputs(1941)) or (layer2_outputs(1598)));
    layer3_outputs(6172) <= '1';
    layer3_outputs(6173) <= (layer2_outputs(4219)) or (layer2_outputs(5031));
    layer3_outputs(6174) <= not(layer2_outputs(7380));
    layer3_outputs(6175) <= layer2_outputs(4433);
    layer3_outputs(6176) <= (layer2_outputs(3585)) and not (layer2_outputs(1022));
    layer3_outputs(6177) <= (layer2_outputs(5154)) and not (layer2_outputs(1306));
    layer3_outputs(6178) <= layer2_outputs(2011);
    layer3_outputs(6179) <= (layer2_outputs(5876)) and not (layer2_outputs(4188));
    layer3_outputs(6180) <= not((layer2_outputs(2836)) xor (layer2_outputs(2209)));
    layer3_outputs(6181) <= (layer2_outputs(3256)) and not (layer2_outputs(3437));
    layer3_outputs(6182) <= layer2_outputs(97);
    layer3_outputs(6183) <= layer2_outputs(1777);
    layer3_outputs(6184) <= not((layer2_outputs(5223)) or (layer2_outputs(5888)));
    layer3_outputs(6185) <= not(layer2_outputs(5751));
    layer3_outputs(6186) <= not(layer2_outputs(4954)) or (layer2_outputs(7186));
    layer3_outputs(6187) <= layer2_outputs(5582);
    layer3_outputs(6188) <= layer2_outputs(1601);
    layer3_outputs(6189) <= not((layer2_outputs(4849)) and (layer2_outputs(2878)));
    layer3_outputs(6190) <= layer2_outputs(3009);
    layer3_outputs(6191) <= (layer2_outputs(5684)) and not (layer2_outputs(1254));
    layer3_outputs(6192) <= '0';
    layer3_outputs(6193) <= not(layer2_outputs(1052));
    layer3_outputs(6194) <= (layer2_outputs(7533)) and (layer2_outputs(449));
    layer3_outputs(6195) <= not(layer2_outputs(5303));
    layer3_outputs(6196) <= not(layer2_outputs(2958));
    layer3_outputs(6197) <= '0';
    layer3_outputs(6198) <= (layer2_outputs(4638)) and not (layer2_outputs(1456));
    layer3_outputs(6199) <= layer2_outputs(5691);
    layer3_outputs(6200) <= not((layer2_outputs(2313)) or (layer2_outputs(703)));
    layer3_outputs(6201) <= not(layer2_outputs(5370)) or (layer2_outputs(5998));
    layer3_outputs(6202) <= not(layer2_outputs(2337));
    layer3_outputs(6203) <= not((layer2_outputs(2913)) or (layer2_outputs(5308)));
    layer3_outputs(6204) <= layer2_outputs(6080);
    layer3_outputs(6205) <= layer2_outputs(4194);
    layer3_outputs(6206) <= (layer2_outputs(4406)) and (layer2_outputs(1131));
    layer3_outputs(6207) <= not((layer2_outputs(7438)) or (layer2_outputs(5326)));
    layer3_outputs(6208) <= layer2_outputs(3330);
    layer3_outputs(6209) <= (layer2_outputs(3465)) or (layer2_outputs(1092));
    layer3_outputs(6210) <= (layer2_outputs(5174)) xor (layer2_outputs(5859));
    layer3_outputs(6211) <= not(layer2_outputs(4587)) or (layer2_outputs(6073));
    layer3_outputs(6212) <= not(layer2_outputs(2217)) or (layer2_outputs(5241));
    layer3_outputs(6213) <= (layer2_outputs(446)) xor (layer2_outputs(5677));
    layer3_outputs(6214) <= (layer2_outputs(7176)) and (layer2_outputs(7443));
    layer3_outputs(6215) <= layer2_outputs(3159);
    layer3_outputs(6216) <= layer2_outputs(1172);
    layer3_outputs(6217) <= not((layer2_outputs(5813)) and (layer2_outputs(4353)));
    layer3_outputs(6218) <= not((layer2_outputs(88)) and (layer2_outputs(4748)));
    layer3_outputs(6219) <= not(layer2_outputs(1335)) or (layer2_outputs(441));
    layer3_outputs(6220) <= not(layer2_outputs(2054));
    layer3_outputs(6221) <= '1';
    layer3_outputs(6222) <= not(layer2_outputs(3215));
    layer3_outputs(6223) <= (layer2_outputs(5211)) and (layer2_outputs(1543));
    layer3_outputs(6224) <= (layer2_outputs(7024)) and not (layer2_outputs(3294));
    layer3_outputs(6225) <= not(layer2_outputs(383));
    layer3_outputs(6226) <= '0';
    layer3_outputs(6227) <= (layer2_outputs(3467)) and (layer2_outputs(4554));
    layer3_outputs(6228) <= not((layer2_outputs(208)) and (layer2_outputs(1588)));
    layer3_outputs(6229) <= layer2_outputs(3137);
    layer3_outputs(6230) <= (layer2_outputs(5828)) and (layer2_outputs(2339));
    layer3_outputs(6231) <= (layer2_outputs(7162)) and not (layer2_outputs(2951));
    layer3_outputs(6232) <= not(layer2_outputs(483));
    layer3_outputs(6233) <= not((layer2_outputs(4000)) or (layer2_outputs(1914)));
    layer3_outputs(6234) <= layer2_outputs(4921);
    layer3_outputs(6235) <= not((layer2_outputs(3007)) xor (layer2_outputs(6674)));
    layer3_outputs(6236) <= not((layer2_outputs(7279)) and (layer2_outputs(1673)));
    layer3_outputs(6237) <= (layer2_outputs(6300)) and not (layer2_outputs(4349));
    layer3_outputs(6238) <= not(layer2_outputs(3450)) or (layer2_outputs(322));
    layer3_outputs(6239) <= not((layer2_outputs(3067)) or (layer2_outputs(3111)));
    layer3_outputs(6240) <= layer2_outputs(471);
    layer3_outputs(6241) <= not(layer2_outputs(5196)) or (layer2_outputs(1471));
    layer3_outputs(6242) <= layer2_outputs(1521);
    layer3_outputs(6243) <= (layer2_outputs(7120)) or (layer2_outputs(4243));
    layer3_outputs(6244) <= (layer2_outputs(2577)) and not (layer2_outputs(5679));
    layer3_outputs(6245) <= not((layer2_outputs(2077)) xor (layer2_outputs(2402)));
    layer3_outputs(6246) <= not(layer2_outputs(2136));
    layer3_outputs(6247) <= not((layer2_outputs(394)) and (layer2_outputs(2144)));
    layer3_outputs(6248) <= not(layer2_outputs(2559)) or (layer2_outputs(2220));
    layer3_outputs(6249) <= not(layer2_outputs(7020)) or (layer2_outputs(5964));
    layer3_outputs(6250) <= not(layer2_outputs(3763));
    layer3_outputs(6251) <= (layer2_outputs(2421)) and not (layer2_outputs(5319));
    layer3_outputs(6252) <= not(layer2_outputs(2230));
    layer3_outputs(6253) <= not(layer2_outputs(4465));
    layer3_outputs(6254) <= layer2_outputs(1137);
    layer3_outputs(6255) <= layer2_outputs(2344);
    layer3_outputs(6256) <= layer2_outputs(3662);
    layer3_outputs(6257) <= '0';
    layer3_outputs(6258) <= layer2_outputs(2837);
    layer3_outputs(6259) <= (layer2_outputs(492)) and (layer2_outputs(532));
    layer3_outputs(6260) <= layer2_outputs(7391);
    layer3_outputs(6261) <= not(layer2_outputs(6353));
    layer3_outputs(6262) <= layer2_outputs(3881);
    layer3_outputs(6263) <= not(layer2_outputs(1650));
    layer3_outputs(6264) <= not((layer2_outputs(2345)) or (layer2_outputs(2059)));
    layer3_outputs(6265) <= (layer2_outputs(4056)) and not (layer2_outputs(1355));
    layer3_outputs(6266) <= not(layer2_outputs(5255));
    layer3_outputs(6267) <= '1';
    layer3_outputs(6268) <= (layer2_outputs(2510)) and (layer2_outputs(3300));
    layer3_outputs(6269) <= not((layer2_outputs(7490)) xor (layer2_outputs(7285)));
    layer3_outputs(6270) <= not((layer2_outputs(961)) and (layer2_outputs(1215)));
    layer3_outputs(6271) <= layer2_outputs(7501);
    layer3_outputs(6272) <= layer2_outputs(7024);
    layer3_outputs(6273) <= not(layer2_outputs(3851));
    layer3_outputs(6274) <= layer2_outputs(7038);
    layer3_outputs(6275) <= (layer2_outputs(4003)) and not (layer2_outputs(6145));
    layer3_outputs(6276) <= not((layer2_outputs(5305)) xor (layer2_outputs(4921)));
    layer3_outputs(6277) <= not(layer2_outputs(4794));
    layer3_outputs(6278) <= not(layer2_outputs(3934)) or (layer2_outputs(3300));
    layer3_outputs(6279) <= (layer2_outputs(2862)) or (layer2_outputs(5879));
    layer3_outputs(6280) <= not(layer2_outputs(1722)) or (layer2_outputs(2852));
    layer3_outputs(6281) <= not(layer2_outputs(2441));
    layer3_outputs(6282) <= not(layer2_outputs(4878)) or (layer2_outputs(5644));
    layer3_outputs(6283) <= '0';
    layer3_outputs(6284) <= not(layer2_outputs(1304)) or (layer2_outputs(2847));
    layer3_outputs(6285) <= layer2_outputs(1048);
    layer3_outputs(6286) <= layer2_outputs(5791);
    layer3_outputs(6287) <= (layer2_outputs(3082)) and (layer2_outputs(6270));
    layer3_outputs(6288) <= (layer2_outputs(6382)) and not (layer2_outputs(2797));
    layer3_outputs(6289) <= not(layer2_outputs(2513));
    layer3_outputs(6290) <= layer2_outputs(1273);
    layer3_outputs(6291) <= layer2_outputs(5915);
    layer3_outputs(6292) <= not((layer2_outputs(7644)) or (layer2_outputs(5740)));
    layer3_outputs(6293) <= layer2_outputs(3727);
    layer3_outputs(6294) <= layer2_outputs(6112);
    layer3_outputs(6295) <= not(layer2_outputs(6997));
    layer3_outputs(6296) <= layer2_outputs(540);
    layer3_outputs(6297) <= layer2_outputs(5911);
    layer3_outputs(6298) <= not(layer2_outputs(6655)) or (layer2_outputs(3179));
    layer3_outputs(6299) <= (layer2_outputs(1518)) and (layer2_outputs(554));
    layer3_outputs(6300) <= not(layer2_outputs(907)) or (layer2_outputs(2952));
    layer3_outputs(6301) <= '1';
    layer3_outputs(6302) <= not(layer2_outputs(6412)) or (layer2_outputs(2145));
    layer3_outputs(6303) <= not(layer2_outputs(2236)) or (layer2_outputs(6876));
    layer3_outputs(6304) <= (layer2_outputs(2086)) or (layer2_outputs(5332));
    layer3_outputs(6305) <= layer2_outputs(4247);
    layer3_outputs(6306) <= layer2_outputs(3228);
    layer3_outputs(6307) <= (layer2_outputs(1197)) or (layer2_outputs(2766));
    layer3_outputs(6308) <= layer2_outputs(5606);
    layer3_outputs(6309) <= not(layer2_outputs(6781));
    layer3_outputs(6310) <= not(layer2_outputs(174)) or (layer2_outputs(1328));
    layer3_outputs(6311) <= (layer2_outputs(1691)) and not (layer2_outputs(4344));
    layer3_outputs(6312) <= not(layer2_outputs(3580)) or (layer2_outputs(4932));
    layer3_outputs(6313) <= layer2_outputs(4774);
    layer3_outputs(6314) <= not(layer2_outputs(294));
    layer3_outputs(6315) <= not(layer2_outputs(1423));
    layer3_outputs(6316) <= layer2_outputs(361);
    layer3_outputs(6317) <= layer2_outputs(1763);
    layer3_outputs(6318) <= '1';
    layer3_outputs(6319) <= layer2_outputs(6447);
    layer3_outputs(6320) <= layer2_outputs(3419);
    layer3_outputs(6321) <= not(layer2_outputs(4896));
    layer3_outputs(6322) <= not(layer2_outputs(7384));
    layer3_outputs(6323) <= not(layer2_outputs(4377));
    layer3_outputs(6324) <= not(layer2_outputs(3823));
    layer3_outputs(6325) <= (layer2_outputs(6554)) or (layer2_outputs(5453));
    layer3_outputs(6326) <= (layer2_outputs(1214)) and not (layer2_outputs(6632));
    layer3_outputs(6327) <= (layer2_outputs(1143)) or (layer2_outputs(6227));
    layer3_outputs(6328) <= (layer2_outputs(5087)) and not (layer2_outputs(3072));
    layer3_outputs(6329) <= layer2_outputs(6760);
    layer3_outputs(6330) <= not(layer2_outputs(7417)) or (layer2_outputs(5628));
    layer3_outputs(6331) <= (layer2_outputs(5639)) or (layer2_outputs(5388));
    layer3_outputs(6332) <= not((layer2_outputs(3722)) xor (layer2_outputs(3488)));
    layer3_outputs(6333) <= not(layer2_outputs(2149));
    layer3_outputs(6334) <= layer2_outputs(4010);
    layer3_outputs(6335) <= not((layer2_outputs(5860)) xor (layer2_outputs(7348)));
    layer3_outputs(6336) <= (layer2_outputs(6065)) and not (layer2_outputs(1278));
    layer3_outputs(6337) <= (layer2_outputs(6945)) and not (layer2_outputs(1218));
    layer3_outputs(6338) <= not(layer2_outputs(349));
    layer3_outputs(6339) <= not((layer2_outputs(202)) or (layer2_outputs(983)));
    layer3_outputs(6340) <= layer2_outputs(3509);
    layer3_outputs(6341) <= not(layer2_outputs(5454));
    layer3_outputs(6342) <= '0';
    layer3_outputs(6343) <= not(layer2_outputs(5739));
    layer3_outputs(6344) <= (layer2_outputs(2269)) or (layer2_outputs(1332));
    layer3_outputs(6345) <= '0';
    layer3_outputs(6346) <= (layer2_outputs(732)) and not (layer2_outputs(2789));
    layer3_outputs(6347) <= layer2_outputs(301);
    layer3_outputs(6348) <= not(layer2_outputs(5877));
    layer3_outputs(6349) <= (layer2_outputs(855)) or (layer2_outputs(2406));
    layer3_outputs(6350) <= (layer2_outputs(2446)) or (layer2_outputs(6062));
    layer3_outputs(6351) <= layer2_outputs(703);
    layer3_outputs(6352) <= not(layer2_outputs(5111));
    layer3_outputs(6353) <= (layer2_outputs(2112)) and (layer2_outputs(4818));
    layer3_outputs(6354) <= (layer2_outputs(4883)) and not (layer2_outputs(988));
    layer3_outputs(6355) <= (layer2_outputs(4698)) and (layer2_outputs(1225));
    layer3_outputs(6356) <= layer2_outputs(5907);
    layer3_outputs(6357) <= not((layer2_outputs(5640)) and (layer2_outputs(1616)));
    layer3_outputs(6358) <= (layer2_outputs(3216)) and not (layer2_outputs(251));
    layer3_outputs(6359) <= not(layer2_outputs(1521));
    layer3_outputs(6360) <= layer2_outputs(7243);
    layer3_outputs(6361) <= not(layer2_outputs(126));
    layer3_outputs(6362) <= not(layer2_outputs(1027)) or (layer2_outputs(1530));
    layer3_outputs(6363) <= not((layer2_outputs(3105)) or (layer2_outputs(2164)));
    layer3_outputs(6364) <= not((layer2_outputs(7420)) or (layer2_outputs(4904)));
    layer3_outputs(6365) <= not(layer2_outputs(7088));
    layer3_outputs(6366) <= not((layer2_outputs(6933)) xor (layer2_outputs(7351)));
    layer3_outputs(6367) <= (layer2_outputs(596)) and not (layer2_outputs(6360));
    layer3_outputs(6368) <= not(layer2_outputs(4892));
    layer3_outputs(6369) <= not((layer2_outputs(6608)) and (layer2_outputs(2702)));
    layer3_outputs(6370) <= (layer2_outputs(2483)) or (layer2_outputs(837));
    layer3_outputs(6371) <= not(layer2_outputs(5922));
    layer3_outputs(6372) <= layer2_outputs(3824);
    layer3_outputs(6373) <= layer2_outputs(6871);
    layer3_outputs(6374) <= not((layer2_outputs(1953)) or (layer2_outputs(6120)));
    layer3_outputs(6375) <= layer2_outputs(2752);
    layer3_outputs(6376) <= not((layer2_outputs(722)) and (layer2_outputs(4840)));
    layer3_outputs(6377) <= layer2_outputs(4118);
    layer3_outputs(6378) <= (layer2_outputs(2020)) and (layer2_outputs(2855));
    layer3_outputs(6379) <= not((layer2_outputs(3587)) and (layer2_outputs(6102)));
    layer3_outputs(6380) <= not(layer2_outputs(4293)) or (layer2_outputs(6408));
    layer3_outputs(6381) <= not((layer2_outputs(4626)) or (layer2_outputs(5478)));
    layer3_outputs(6382) <= (layer2_outputs(3110)) and not (layer2_outputs(4560));
    layer3_outputs(6383) <= '1';
    layer3_outputs(6384) <= layer2_outputs(1109);
    layer3_outputs(6385) <= (layer2_outputs(983)) and not (layer2_outputs(661));
    layer3_outputs(6386) <= layer2_outputs(3180);
    layer3_outputs(6387) <= not(layer2_outputs(5247)) or (layer2_outputs(372));
    layer3_outputs(6388) <= not(layer2_outputs(7516));
    layer3_outputs(6389) <= layer2_outputs(1036);
    layer3_outputs(6390) <= layer2_outputs(4160);
    layer3_outputs(6391) <= not(layer2_outputs(4759)) or (layer2_outputs(800));
    layer3_outputs(6392) <= not(layer2_outputs(5324));
    layer3_outputs(6393) <= not((layer2_outputs(3149)) or (layer2_outputs(7026)));
    layer3_outputs(6394) <= not(layer2_outputs(5821));
    layer3_outputs(6395) <= (layer2_outputs(2478)) xor (layer2_outputs(5789));
    layer3_outputs(6396) <= layer2_outputs(3305);
    layer3_outputs(6397) <= layer2_outputs(7378);
    layer3_outputs(6398) <= (layer2_outputs(837)) xor (layer2_outputs(655));
    layer3_outputs(6399) <= '1';
    layer3_outputs(6400) <= (layer2_outputs(3269)) or (layer2_outputs(7301));
    layer3_outputs(6401) <= not((layer2_outputs(6023)) or (layer2_outputs(4727)));
    layer3_outputs(6402) <= not(layer2_outputs(1164));
    layer3_outputs(6403) <= layer2_outputs(5910);
    layer3_outputs(6404) <= not(layer2_outputs(6074)) or (layer2_outputs(36));
    layer3_outputs(6405) <= layer2_outputs(6056);
    layer3_outputs(6406) <= layer2_outputs(1873);
    layer3_outputs(6407) <= (layer2_outputs(2440)) and (layer2_outputs(5482));
    layer3_outputs(6408) <= layer2_outputs(7077);
    layer3_outputs(6409) <= layer2_outputs(3418);
    layer3_outputs(6410) <= (layer2_outputs(5120)) and not (layer2_outputs(5109));
    layer3_outputs(6411) <= not(layer2_outputs(2214));
    layer3_outputs(6412) <= layer2_outputs(6759);
    layer3_outputs(6413) <= not(layer2_outputs(2609));
    layer3_outputs(6414) <= not(layer2_outputs(1070)) or (layer2_outputs(6528));
    layer3_outputs(6415) <= layer2_outputs(7618);
    layer3_outputs(6416) <= not((layer2_outputs(515)) and (layer2_outputs(4271)));
    layer3_outputs(6417) <= (layer2_outputs(175)) and (layer2_outputs(116));
    layer3_outputs(6418) <= not(layer2_outputs(5049)) or (layer2_outputs(4260));
    layer3_outputs(6419) <= not(layer2_outputs(6443));
    layer3_outputs(6420) <= not((layer2_outputs(4172)) or (layer2_outputs(6862)));
    layer3_outputs(6421) <= not(layer2_outputs(1556));
    layer3_outputs(6422) <= layer2_outputs(1524);
    layer3_outputs(6423) <= (layer2_outputs(3059)) or (layer2_outputs(332));
    layer3_outputs(6424) <= (layer2_outputs(2435)) and not (layer2_outputs(2793));
    layer3_outputs(6425) <= not(layer2_outputs(4222));
    layer3_outputs(6426) <= not((layer2_outputs(4936)) and (layer2_outputs(3717)));
    layer3_outputs(6427) <= not(layer2_outputs(4814)) or (layer2_outputs(5766));
    layer3_outputs(6428) <= layer2_outputs(2299);
    layer3_outputs(6429) <= not(layer2_outputs(5612));
    layer3_outputs(6430) <= not((layer2_outputs(1602)) and (layer2_outputs(2742)));
    layer3_outputs(6431) <= not((layer2_outputs(4115)) xor (layer2_outputs(3138)));
    layer3_outputs(6432) <= layer2_outputs(1830);
    layer3_outputs(6433) <= not((layer2_outputs(5641)) or (layer2_outputs(3241)));
    layer3_outputs(6434) <= layer2_outputs(4123);
    layer3_outputs(6435) <= not((layer2_outputs(4044)) xor (layer2_outputs(1236)));
    layer3_outputs(6436) <= not((layer2_outputs(3959)) xor (layer2_outputs(6291)));
    layer3_outputs(6437) <= not(layer2_outputs(5699));
    layer3_outputs(6438) <= (layer2_outputs(7334)) xor (layer2_outputs(7553));
    layer3_outputs(6439) <= not((layer2_outputs(502)) or (layer2_outputs(7182)));
    layer3_outputs(6440) <= layer2_outputs(2475);
    layer3_outputs(6441) <= not(layer2_outputs(446));
    layer3_outputs(6442) <= not(layer2_outputs(6123)) or (layer2_outputs(6734));
    layer3_outputs(6443) <= layer2_outputs(7190);
    layer3_outputs(6444) <= (layer2_outputs(3874)) or (layer2_outputs(2766));
    layer3_outputs(6445) <= (layer2_outputs(7537)) and not (layer2_outputs(2386));
    layer3_outputs(6446) <= not(layer2_outputs(3591));
    layer3_outputs(6447) <= layer2_outputs(2811);
    layer3_outputs(6448) <= (layer2_outputs(2987)) and (layer2_outputs(2274));
    layer3_outputs(6449) <= not(layer2_outputs(1213));
    layer3_outputs(6450) <= (layer2_outputs(5408)) or (layer2_outputs(2759));
    layer3_outputs(6451) <= layer2_outputs(634);
    layer3_outputs(6452) <= (layer2_outputs(1711)) and not (layer2_outputs(4965));
    layer3_outputs(6453) <= layer2_outputs(7437);
    layer3_outputs(6454) <= (layer2_outputs(6046)) xor (layer2_outputs(2346));
    layer3_outputs(6455) <= '0';
    layer3_outputs(6456) <= (layer2_outputs(77)) and not (layer2_outputs(6968));
    layer3_outputs(6457) <= layer2_outputs(1216);
    layer3_outputs(6458) <= (layer2_outputs(1999)) and not (layer2_outputs(4916));
    layer3_outputs(6459) <= layer2_outputs(7163);
    layer3_outputs(6460) <= (layer2_outputs(2001)) and not (layer2_outputs(7183));
    layer3_outputs(6461) <= not(layer2_outputs(7498));
    layer3_outputs(6462) <= (layer2_outputs(7299)) and not (layer2_outputs(411));
    layer3_outputs(6463) <= (layer2_outputs(1688)) and not (layer2_outputs(7436));
    layer3_outputs(6464) <= layer2_outputs(5021);
    layer3_outputs(6465) <= (layer2_outputs(746)) and not (layer2_outputs(4650));
    layer3_outputs(6466) <= not((layer2_outputs(5250)) and (layer2_outputs(5345)));
    layer3_outputs(6467) <= not(layer2_outputs(6505));
    layer3_outputs(6468) <= layer2_outputs(3517);
    layer3_outputs(6469) <= not(layer2_outputs(264)) or (layer2_outputs(2160));
    layer3_outputs(6470) <= not((layer2_outputs(5656)) or (layer2_outputs(5025)));
    layer3_outputs(6471) <= (layer2_outputs(3129)) and not (layer2_outputs(1309));
    layer3_outputs(6472) <= (layer2_outputs(3393)) or (layer2_outputs(10));
    layer3_outputs(6473) <= not(layer2_outputs(50));
    layer3_outputs(6474) <= not((layer2_outputs(6498)) xor (layer2_outputs(405)));
    layer3_outputs(6475) <= (layer2_outputs(2125)) and not (layer2_outputs(7212));
    layer3_outputs(6476) <= not(layer2_outputs(6748)) or (layer2_outputs(319));
    layer3_outputs(6477) <= not(layer2_outputs(1405));
    layer3_outputs(6478) <= '1';
    layer3_outputs(6479) <= (layer2_outputs(6180)) and not (layer2_outputs(984));
    layer3_outputs(6480) <= layer2_outputs(1421);
    layer3_outputs(6481) <= (layer2_outputs(6160)) and not (layer2_outputs(1569));
    layer3_outputs(6482) <= not(layer2_outputs(6879));
    layer3_outputs(6483) <= not((layer2_outputs(1074)) and (layer2_outputs(6478)));
    layer3_outputs(6484) <= not(layer2_outputs(1910)) or (layer2_outputs(2616));
    layer3_outputs(6485) <= not(layer2_outputs(6476));
    layer3_outputs(6486) <= not(layer2_outputs(2880));
    layer3_outputs(6487) <= not(layer2_outputs(977));
    layer3_outputs(6488) <= layer2_outputs(5582);
    layer3_outputs(6489) <= (layer2_outputs(6547)) xor (layer2_outputs(167));
    layer3_outputs(6490) <= (layer2_outputs(6979)) and not (layer2_outputs(3768));
    layer3_outputs(6491) <= not(layer2_outputs(791));
    layer3_outputs(6492) <= not(layer2_outputs(2060)) or (layer2_outputs(3942));
    layer3_outputs(6493) <= layer2_outputs(5);
    layer3_outputs(6494) <= (layer2_outputs(3144)) and (layer2_outputs(6888));
    layer3_outputs(6495) <= not(layer2_outputs(2354)) or (layer2_outputs(2518));
    layer3_outputs(6496) <= not(layer2_outputs(7620));
    layer3_outputs(6497) <= (layer2_outputs(5056)) or (layer2_outputs(5983));
    layer3_outputs(6498) <= not(layer2_outputs(1468));
    layer3_outputs(6499) <= (layer2_outputs(63)) and not (layer2_outputs(2115));
    layer3_outputs(6500) <= (layer2_outputs(2449)) and not (layer2_outputs(4514));
    layer3_outputs(6501) <= not(layer2_outputs(5226)) or (layer2_outputs(7218));
    layer3_outputs(6502) <= not(layer2_outputs(4031));
    layer3_outputs(6503) <= '0';
    layer3_outputs(6504) <= not((layer2_outputs(6130)) and (layer2_outputs(336)));
    layer3_outputs(6505) <= layer2_outputs(6202);
    layer3_outputs(6506) <= '1';
    layer3_outputs(6507) <= not(layer2_outputs(5567)) or (layer2_outputs(2610));
    layer3_outputs(6508) <= layer2_outputs(3808);
    layer3_outputs(6509) <= (layer2_outputs(5251)) or (layer2_outputs(1903));
    layer3_outputs(6510) <= not(layer2_outputs(7096)) or (layer2_outputs(3310));
    layer3_outputs(6511) <= not(layer2_outputs(2711));
    layer3_outputs(6512) <= '0';
    layer3_outputs(6513) <= (layer2_outputs(6615)) and not (layer2_outputs(5902));
    layer3_outputs(6514) <= not(layer2_outputs(2388));
    layer3_outputs(6515) <= not((layer2_outputs(7588)) or (layer2_outputs(44)));
    layer3_outputs(6516) <= not(layer2_outputs(2966));
    layer3_outputs(6517) <= (layer2_outputs(5558)) xor (layer2_outputs(3312));
    layer3_outputs(6518) <= not(layer2_outputs(3756));
    layer3_outputs(6519) <= (layer2_outputs(2347)) or (layer2_outputs(5239));
    layer3_outputs(6520) <= (layer2_outputs(4134)) xor (layer2_outputs(4796));
    layer3_outputs(6521) <= not(layer2_outputs(3965)) or (layer2_outputs(2274));
    layer3_outputs(6522) <= '0';
    layer3_outputs(6523) <= not(layer2_outputs(5516));
    layer3_outputs(6524) <= layer2_outputs(1300);
    layer3_outputs(6525) <= not(layer2_outputs(4217));
    layer3_outputs(6526) <= not(layer2_outputs(5637));
    layer3_outputs(6527) <= not((layer2_outputs(7379)) xor (layer2_outputs(2309)));
    layer3_outputs(6528) <= not((layer2_outputs(249)) or (layer2_outputs(3912)));
    layer3_outputs(6529) <= not(layer2_outputs(4023)) or (layer2_outputs(2728));
    layer3_outputs(6530) <= not((layer2_outputs(4570)) xor (layer2_outputs(4691)));
    layer3_outputs(6531) <= layer2_outputs(3008);
    layer3_outputs(6532) <= layer2_outputs(6180);
    layer3_outputs(6533) <= not((layer2_outputs(2448)) xor (layer2_outputs(5576)));
    layer3_outputs(6534) <= not(layer2_outputs(6462));
    layer3_outputs(6535) <= (layer2_outputs(2396)) or (layer2_outputs(2495));
    layer3_outputs(6536) <= not(layer2_outputs(6988));
    layer3_outputs(6537) <= not(layer2_outputs(5324));
    layer3_outputs(6538) <= not(layer2_outputs(1382));
    layer3_outputs(6539) <= not(layer2_outputs(5986));
    layer3_outputs(6540) <= not(layer2_outputs(2037));
    layer3_outputs(6541) <= layer2_outputs(1010);
    layer3_outputs(6542) <= layer2_outputs(4746);
    layer3_outputs(6543) <= not(layer2_outputs(3481));
    layer3_outputs(6544) <= not((layer2_outputs(7447)) or (layer2_outputs(4481)));
    layer3_outputs(6545) <= layer2_outputs(5103);
    layer3_outputs(6546) <= layer2_outputs(4526);
    layer3_outputs(6547) <= not(layer2_outputs(7628));
    layer3_outputs(6548) <= (layer2_outputs(5992)) and not (layer2_outputs(6640));
    layer3_outputs(6549) <= not(layer2_outputs(4518)) or (layer2_outputs(1882));
    layer3_outputs(6550) <= not((layer2_outputs(1274)) or (layer2_outputs(5827)));
    layer3_outputs(6551) <= layer2_outputs(878);
    layer3_outputs(6552) <= not(layer2_outputs(7459));
    layer3_outputs(6553) <= layer2_outputs(4614);
    layer3_outputs(6554) <= (layer2_outputs(306)) or (layer2_outputs(3207));
    layer3_outputs(6555) <= not(layer2_outputs(6106)) or (layer2_outputs(3192));
    layer3_outputs(6556) <= not(layer2_outputs(2219));
    layer3_outputs(6557) <= layer2_outputs(7520);
    layer3_outputs(6558) <= (layer2_outputs(7197)) and not (layer2_outputs(2151));
    layer3_outputs(6559) <= layer2_outputs(2643);
    layer3_outputs(6560) <= not(layer2_outputs(6745));
    layer3_outputs(6561) <= not(layer2_outputs(2682)) or (layer2_outputs(4024));
    layer3_outputs(6562) <= layer2_outputs(2338);
    layer3_outputs(6563) <= not(layer2_outputs(6323)) or (layer2_outputs(1628));
    layer3_outputs(6564) <= layer2_outputs(7281);
    layer3_outputs(6565) <= (layer2_outputs(30)) xor (layer2_outputs(3761));
    layer3_outputs(6566) <= layer2_outputs(5018);
    layer3_outputs(6567) <= not(layer2_outputs(6065));
    layer3_outputs(6568) <= layer2_outputs(5510);
    layer3_outputs(6569) <= (layer2_outputs(7345)) and (layer2_outputs(3846));
    layer3_outputs(6570) <= layer2_outputs(3559);
    layer3_outputs(6571) <= layer2_outputs(5693);
    layer3_outputs(6572) <= (layer2_outputs(4137)) and not (layer2_outputs(3687));
    layer3_outputs(6573) <= (layer2_outputs(6880)) xor (layer2_outputs(5804));
    layer3_outputs(6574) <= (layer2_outputs(1003)) and not (layer2_outputs(1511));
    layer3_outputs(6575) <= (layer2_outputs(2574)) and (layer2_outputs(1145));
    layer3_outputs(6576) <= not(layer2_outputs(6918));
    layer3_outputs(6577) <= (layer2_outputs(5530)) and not (layer2_outputs(252));
    layer3_outputs(6578) <= (layer2_outputs(7068)) or (layer2_outputs(5588));
    layer3_outputs(6579) <= (layer2_outputs(4103)) and not (layer2_outputs(2495));
    layer3_outputs(6580) <= not(layer2_outputs(726));
    layer3_outputs(6581) <= not(layer2_outputs(3974));
    layer3_outputs(6582) <= layer2_outputs(1469);
    layer3_outputs(6583) <= (layer2_outputs(6585)) or (layer2_outputs(6946));
    layer3_outputs(6584) <= not((layer2_outputs(5892)) and (layer2_outputs(4805)));
    layer3_outputs(6585) <= not((layer2_outputs(6365)) and (layer2_outputs(6730)));
    layer3_outputs(6586) <= not((layer2_outputs(5889)) or (layer2_outputs(642)));
    layer3_outputs(6587) <= not(layer2_outputs(7495));
    layer3_outputs(6588) <= not(layer2_outputs(1253)) or (layer2_outputs(1803));
    layer3_outputs(6589) <= not((layer2_outputs(2864)) or (layer2_outputs(6276)));
    layer3_outputs(6590) <= (layer2_outputs(7060)) and not (layer2_outputs(195));
    layer3_outputs(6591) <= (layer2_outputs(7286)) and not (layer2_outputs(2877));
    layer3_outputs(6592) <= '0';
    layer3_outputs(6593) <= layer2_outputs(4153);
    layer3_outputs(6594) <= not((layer2_outputs(4060)) xor (layer2_outputs(4383)));
    layer3_outputs(6595) <= layer2_outputs(4654);
    layer3_outputs(6596) <= not((layer2_outputs(3496)) and (layer2_outputs(4483)));
    layer3_outputs(6597) <= not(layer2_outputs(3208));
    layer3_outputs(6598) <= '0';
    layer3_outputs(6599) <= not((layer2_outputs(3742)) or (layer2_outputs(2307)));
    layer3_outputs(6600) <= not(layer2_outputs(1169)) or (layer2_outputs(3777));
    layer3_outputs(6601) <= (layer2_outputs(5989)) xor (layer2_outputs(4400));
    layer3_outputs(6602) <= not(layer2_outputs(4239)) or (layer2_outputs(3741));
    layer3_outputs(6603) <= not(layer2_outputs(3329));
    layer3_outputs(6604) <= not((layer2_outputs(784)) and (layer2_outputs(7597)));
    layer3_outputs(6605) <= (layer2_outputs(5110)) and (layer2_outputs(699));
    layer3_outputs(6606) <= (layer2_outputs(1185)) xor (layer2_outputs(2782));
    layer3_outputs(6607) <= layer2_outputs(7078);
    layer3_outputs(6608) <= layer2_outputs(4398);
    layer3_outputs(6609) <= not(layer2_outputs(7651));
    layer3_outputs(6610) <= not(layer2_outputs(920));
    layer3_outputs(6611) <= not(layer2_outputs(2481)) or (layer2_outputs(6824));
    layer3_outputs(6612) <= not(layer2_outputs(2190));
    layer3_outputs(6613) <= (layer2_outputs(2446)) or (layer2_outputs(6334));
    layer3_outputs(6614) <= (layer2_outputs(6762)) xor (layer2_outputs(6074));
    layer3_outputs(6615) <= not((layer2_outputs(6559)) or (layer2_outputs(3707)));
    layer3_outputs(6616) <= not(layer2_outputs(2158));
    layer3_outputs(6617) <= layer2_outputs(4664);
    layer3_outputs(6618) <= not(layer2_outputs(3808)) or (layer2_outputs(4766));
    layer3_outputs(6619) <= not(layer2_outputs(3009));
    layer3_outputs(6620) <= (layer2_outputs(2621)) and not (layer2_outputs(6083));
    layer3_outputs(6621) <= (layer2_outputs(4335)) and not (layer2_outputs(3128));
    layer3_outputs(6622) <= not(layer2_outputs(4542));
    layer3_outputs(6623) <= (layer2_outputs(7017)) and not (layer2_outputs(3396));
    layer3_outputs(6624) <= (layer2_outputs(3645)) and not (layer2_outputs(4919));
    layer3_outputs(6625) <= not((layer2_outputs(5563)) and (layer2_outputs(5968)));
    layer3_outputs(6626) <= not(layer2_outputs(1696)) or (layer2_outputs(5646));
    layer3_outputs(6627) <= (layer2_outputs(56)) and (layer2_outputs(5479));
    layer3_outputs(6628) <= not(layer2_outputs(3854));
    layer3_outputs(6629) <= not(layer2_outputs(3739));
    layer3_outputs(6630) <= not(layer2_outputs(4682));
    layer3_outputs(6631) <= layer2_outputs(975);
    layer3_outputs(6632) <= layer2_outputs(6488);
    layer3_outputs(6633) <= (layer2_outputs(2868)) and (layer2_outputs(14));
    layer3_outputs(6634) <= layer2_outputs(3514);
    layer3_outputs(6635) <= not(layer2_outputs(551));
    layer3_outputs(6636) <= (layer2_outputs(4241)) or (layer2_outputs(2899));
    layer3_outputs(6637) <= not(layer2_outputs(3387));
    layer3_outputs(6638) <= not(layer2_outputs(320)) or (layer2_outputs(483));
    layer3_outputs(6639) <= layer2_outputs(6851);
    layer3_outputs(6640) <= not((layer2_outputs(4876)) and (layer2_outputs(5249)));
    layer3_outputs(6641) <= not(layer2_outputs(2508)) or (layer2_outputs(670));
    layer3_outputs(6642) <= not((layer2_outputs(6697)) or (layer2_outputs(5079)));
    layer3_outputs(6643) <= layer2_outputs(459);
    layer3_outputs(6644) <= not((layer2_outputs(4305)) or (layer2_outputs(3861)));
    layer3_outputs(6645) <= not(layer2_outputs(5116));
    layer3_outputs(6646) <= '0';
    layer3_outputs(6647) <= (layer2_outputs(1865)) and not (layer2_outputs(2658));
    layer3_outputs(6648) <= layer2_outputs(1169);
    layer3_outputs(6649) <= (layer2_outputs(205)) or (layer2_outputs(6112));
    layer3_outputs(6650) <= layer2_outputs(3789);
    layer3_outputs(6651) <= not(layer2_outputs(2493)) or (layer2_outputs(5810));
    layer3_outputs(6652) <= not((layer2_outputs(2459)) xor (layer2_outputs(4988)));
    layer3_outputs(6653) <= layer2_outputs(1409);
    layer3_outputs(6654) <= (layer2_outputs(2498)) or (layer2_outputs(2824));
    layer3_outputs(6655) <= (layer2_outputs(7476)) and not (layer2_outputs(5392));
    layer3_outputs(6656) <= not((layer2_outputs(7)) or (layer2_outputs(6839)));
    layer3_outputs(6657) <= layer2_outputs(7464);
    layer3_outputs(6658) <= not(layer2_outputs(4685)) or (layer2_outputs(4552));
    layer3_outputs(6659) <= (layer2_outputs(886)) and not (layer2_outputs(6605));
    layer3_outputs(6660) <= not(layer2_outputs(2318));
    layer3_outputs(6661) <= not(layer2_outputs(3953)) or (layer2_outputs(3055));
    layer3_outputs(6662) <= (layer2_outputs(2271)) or (layer2_outputs(7324));
    layer3_outputs(6663) <= not((layer2_outputs(380)) xor (layer2_outputs(980)));
    layer3_outputs(6664) <= not((layer2_outputs(5474)) and (layer2_outputs(3201)));
    layer3_outputs(6665) <= not(layer2_outputs(4371)) or (layer2_outputs(6430));
    layer3_outputs(6666) <= layer2_outputs(879);
    layer3_outputs(6667) <= not(layer2_outputs(7356));
    layer3_outputs(6668) <= (layer2_outputs(1344)) and not (layer2_outputs(7459));
    layer3_outputs(6669) <= not(layer2_outputs(6159));
    layer3_outputs(6670) <= not(layer2_outputs(1843));
    layer3_outputs(6671) <= (layer2_outputs(1829)) and (layer2_outputs(2356));
    layer3_outputs(6672) <= not(layer2_outputs(5816));
    layer3_outputs(6673) <= not((layer2_outputs(5746)) and (layer2_outputs(6436)));
    layer3_outputs(6674) <= not((layer2_outputs(513)) or (layer2_outputs(280)));
    layer3_outputs(6675) <= (layer2_outputs(143)) and (layer2_outputs(2966));
    layer3_outputs(6676) <= not(layer2_outputs(5428));
    layer3_outputs(6677) <= layer2_outputs(5689);
    layer3_outputs(6678) <= not(layer2_outputs(1956)) or (layer2_outputs(261));
    layer3_outputs(6679) <= not(layer2_outputs(5841)) or (layer2_outputs(3177));
    layer3_outputs(6680) <= layer2_outputs(5157);
    layer3_outputs(6681) <= '0';
    layer3_outputs(6682) <= not((layer2_outputs(1136)) xor (layer2_outputs(7428)));
    layer3_outputs(6683) <= not(layer2_outputs(3145));
    layer3_outputs(6684) <= (layer2_outputs(840)) and (layer2_outputs(3359));
    layer3_outputs(6685) <= layer2_outputs(3430);
    layer3_outputs(6686) <= layer2_outputs(4410);
    layer3_outputs(6687) <= layer2_outputs(4811);
    layer3_outputs(6688) <= not(layer2_outputs(1552));
    layer3_outputs(6689) <= (layer2_outputs(2799)) or (layer2_outputs(4767));
    layer3_outputs(6690) <= (layer2_outputs(4966)) or (layer2_outputs(1283));
    layer3_outputs(6691) <= not(layer2_outputs(3055));
    layer3_outputs(6692) <= (layer2_outputs(3214)) or (layer2_outputs(3097));
    layer3_outputs(6693) <= not((layer2_outputs(74)) and (layer2_outputs(6533)));
    layer3_outputs(6694) <= not((layer2_outputs(1747)) or (layer2_outputs(3158)));
    layer3_outputs(6695) <= (layer2_outputs(686)) and not (layer2_outputs(3142));
    layer3_outputs(6696) <= not(layer2_outputs(4513)) or (layer2_outputs(417));
    layer3_outputs(6697) <= not(layer2_outputs(4491));
    layer3_outputs(6698) <= (layer2_outputs(6502)) and (layer2_outputs(6866));
    layer3_outputs(6699) <= not(layer2_outputs(404));
    layer3_outputs(6700) <= layer2_outputs(4414);
    layer3_outputs(6701) <= not((layer2_outputs(3704)) or (layer2_outputs(5371)));
    layer3_outputs(6702) <= (layer2_outputs(6478)) and (layer2_outputs(3949));
    layer3_outputs(6703) <= (layer2_outputs(5919)) and (layer2_outputs(1656));
    layer3_outputs(6704) <= (layer2_outputs(7396)) and (layer2_outputs(2324));
    layer3_outputs(6705) <= not(layer2_outputs(4278));
    layer3_outputs(6706) <= (layer2_outputs(4808)) and not (layer2_outputs(1887));
    layer3_outputs(6707) <= layer2_outputs(1388);
    layer3_outputs(6708) <= '0';
    layer3_outputs(6709) <= not(layer2_outputs(319));
    layer3_outputs(6710) <= layer2_outputs(3964);
    layer3_outputs(6711) <= not((layer2_outputs(2474)) or (layer2_outputs(2090)));
    layer3_outputs(6712) <= not((layer2_outputs(1288)) or (layer2_outputs(2449)));
    layer3_outputs(6713) <= layer2_outputs(6764);
    layer3_outputs(6714) <= layer2_outputs(1329);
    layer3_outputs(6715) <= layer2_outputs(5603);
    layer3_outputs(6716) <= not(layer2_outputs(1087));
    layer3_outputs(6717) <= (layer2_outputs(3989)) and not (layer2_outputs(7659));
    layer3_outputs(6718) <= layer2_outputs(5638);
    layer3_outputs(6719) <= not(layer2_outputs(4624));
    layer3_outputs(6720) <= not((layer2_outputs(7179)) xor (layer2_outputs(22)));
    layer3_outputs(6721) <= layer2_outputs(821);
    layer3_outputs(6722) <= not(layer2_outputs(5041));
    layer3_outputs(6723) <= not(layer2_outputs(4936)) or (layer2_outputs(688));
    layer3_outputs(6724) <= layer2_outputs(1108);
    layer3_outputs(6725) <= not(layer2_outputs(1415)) or (layer2_outputs(3825));
    layer3_outputs(6726) <= (layer2_outputs(169)) or (layer2_outputs(1128));
    layer3_outputs(6727) <= (layer2_outputs(6560)) xor (layer2_outputs(6254));
    layer3_outputs(6728) <= (layer2_outputs(5650)) and not (layer2_outputs(6768));
    layer3_outputs(6729) <= not((layer2_outputs(1918)) xor (layer2_outputs(6389)));
    layer3_outputs(6730) <= '0';
    layer3_outputs(6731) <= not((layer2_outputs(2015)) or (layer2_outputs(2136)));
    layer3_outputs(6732) <= layer2_outputs(6158);
    layer3_outputs(6733) <= layer2_outputs(3820);
    layer3_outputs(6734) <= (layer2_outputs(7409)) xor (layer2_outputs(401));
    layer3_outputs(6735) <= layer2_outputs(4915);
    layer3_outputs(6736) <= not((layer2_outputs(6594)) xor (layer2_outputs(5082)));
    layer3_outputs(6737) <= not((layer2_outputs(3312)) and (layer2_outputs(5951)));
    layer3_outputs(6738) <= not(layer2_outputs(2267));
    layer3_outputs(6739) <= not(layer2_outputs(2768)) or (layer2_outputs(6710));
    layer3_outputs(6740) <= (layer2_outputs(7443)) and not (layer2_outputs(2423));
    layer3_outputs(6741) <= layer2_outputs(7085);
    layer3_outputs(6742) <= (layer2_outputs(2911)) xor (layer2_outputs(6806));
    layer3_outputs(6743) <= not(layer2_outputs(1403));
    layer3_outputs(6744) <= layer2_outputs(4845);
    layer3_outputs(6745) <= not((layer2_outputs(2635)) or (layer2_outputs(1361)));
    layer3_outputs(6746) <= not(layer2_outputs(1712)) or (layer2_outputs(1333));
    layer3_outputs(6747) <= (layer2_outputs(1584)) and not (layer2_outputs(5969));
    layer3_outputs(6748) <= layer2_outputs(5264);
    layer3_outputs(6749) <= layer2_outputs(1618);
    layer3_outputs(6750) <= layer2_outputs(3361);
    layer3_outputs(6751) <= (layer2_outputs(1181)) and not (layer2_outputs(4933));
    layer3_outputs(6752) <= (layer2_outputs(1927)) and not (layer2_outputs(746));
    layer3_outputs(6753) <= not(layer2_outputs(6631));
    layer3_outputs(6754) <= layer2_outputs(7665);
    layer3_outputs(6755) <= not(layer2_outputs(7344));
    layer3_outputs(6756) <= not(layer2_outputs(4265));
    layer3_outputs(6757) <= '1';
    layer3_outputs(6758) <= not(layer2_outputs(2506));
    layer3_outputs(6759) <= layer2_outputs(5335);
    layer3_outputs(6760) <= not(layer2_outputs(3618));
    layer3_outputs(6761) <= (layer2_outputs(6942)) and not (layer2_outputs(7591));
    layer3_outputs(6762) <= layer2_outputs(6620);
    layer3_outputs(6763) <= not((layer2_outputs(3740)) and (layer2_outputs(2894)));
    layer3_outputs(6764) <= layer2_outputs(4083);
    layer3_outputs(6765) <= not((layer2_outputs(7338)) xor (layer2_outputs(4469)));
    layer3_outputs(6766) <= (layer2_outputs(5635)) and (layer2_outputs(6529));
    layer3_outputs(6767) <= not((layer2_outputs(2430)) and (layer2_outputs(3248)));
    layer3_outputs(6768) <= layer2_outputs(3075);
    layer3_outputs(6769) <= '0';
    layer3_outputs(6770) <= layer2_outputs(2844);
    layer3_outputs(6771) <= layer2_outputs(5917);
    layer3_outputs(6772) <= (layer2_outputs(6253)) and not (layer2_outputs(951));
    layer3_outputs(6773) <= not(layer2_outputs(2918)) or (layer2_outputs(6630));
    layer3_outputs(6774) <= (layer2_outputs(7424)) and (layer2_outputs(4837));
    layer3_outputs(6775) <= not((layer2_outputs(1881)) or (layer2_outputs(6027)));
    layer3_outputs(6776) <= layer2_outputs(5488);
    layer3_outputs(6777) <= layer2_outputs(768);
    layer3_outputs(6778) <= not((layer2_outputs(711)) or (layer2_outputs(5158)));
    layer3_outputs(6779) <= not(layer2_outputs(4606));
    layer3_outputs(6780) <= not(layer2_outputs(4930)) or (layer2_outputs(2734));
    layer3_outputs(6781) <= layer2_outputs(5735);
    layer3_outputs(6782) <= not(layer2_outputs(212));
    layer3_outputs(6783) <= not(layer2_outputs(7240));
    layer3_outputs(6784) <= (layer2_outputs(5180)) and not (layer2_outputs(369));
    layer3_outputs(6785) <= layer2_outputs(6919);
    layer3_outputs(6786) <= not(layer2_outputs(7393));
    layer3_outputs(6787) <= not((layer2_outputs(324)) or (layer2_outputs(4951)));
    layer3_outputs(6788) <= not((layer2_outputs(5458)) xor (layer2_outputs(6450)));
    layer3_outputs(6789) <= (layer2_outputs(5716)) and not (layer2_outputs(305));
    layer3_outputs(6790) <= (layer2_outputs(5691)) or (layer2_outputs(5899));
    layer3_outputs(6791) <= '0';
    layer3_outputs(6792) <= not((layer2_outputs(5916)) and (layer2_outputs(2731)));
    layer3_outputs(6793) <= not(layer2_outputs(3519));
    layer3_outputs(6794) <= not(layer2_outputs(7579));
    layer3_outputs(6795) <= not((layer2_outputs(1319)) or (layer2_outputs(3094)));
    layer3_outputs(6796) <= not(layer2_outputs(760));
    layer3_outputs(6797) <= not(layer2_outputs(6119)) or (layer2_outputs(2701));
    layer3_outputs(6798) <= not((layer2_outputs(5326)) and (layer2_outputs(2764)));
    layer3_outputs(6799) <= not(layer2_outputs(218)) or (layer2_outputs(4649));
    layer3_outputs(6800) <= (layer2_outputs(5140)) and not (layer2_outputs(876));
    layer3_outputs(6801) <= not((layer2_outputs(6229)) and (layer2_outputs(2950)));
    layer3_outputs(6802) <= not(layer2_outputs(3903));
    layer3_outputs(6803) <= not(layer2_outputs(5300)) or (layer2_outputs(7543));
    layer3_outputs(6804) <= not(layer2_outputs(5757)) or (layer2_outputs(2873));
    layer3_outputs(6805) <= layer2_outputs(2417);
    layer3_outputs(6806) <= (layer2_outputs(5188)) and not (layer2_outputs(1117));
    layer3_outputs(6807) <= (layer2_outputs(5809)) and (layer2_outputs(3860));
    layer3_outputs(6808) <= not(layer2_outputs(911));
    layer3_outputs(6809) <= not(layer2_outputs(5782));
    layer3_outputs(6810) <= not((layer2_outputs(1267)) xor (layer2_outputs(6481)));
    layer3_outputs(6811) <= layer2_outputs(2063);
    layer3_outputs(6812) <= (layer2_outputs(220)) and not (layer2_outputs(2817));
    layer3_outputs(6813) <= (layer2_outputs(2370)) or (layer2_outputs(2147));
    layer3_outputs(6814) <= not((layer2_outputs(3334)) and (layer2_outputs(730)));
    layer3_outputs(6815) <= not(layer2_outputs(6064));
    layer3_outputs(6816) <= not(layer2_outputs(2100));
    layer3_outputs(6817) <= not(layer2_outputs(6570));
    layer3_outputs(6818) <= not(layer2_outputs(5160)) or (layer2_outputs(1483));
    layer3_outputs(6819) <= not(layer2_outputs(531));
    layer3_outputs(6820) <= (layer2_outputs(858)) and not (layer2_outputs(7615));
    layer3_outputs(6821) <= (layer2_outputs(2464)) and not (layer2_outputs(3804));
    layer3_outputs(6822) <= not(layer2_outputs(4379));
    layer3_outputs(6823) <= '0';
    layer3_outputs(6824) <= '1';
    layer3_outputs(6825) <= layer2_outputs(6310);
    layer3_outputs(6826) <= not(layer2_outputs(5629));
    layer3_outputs(6827) <= not(layer2_outputs(225)) or (layer2_outputs(3703));
    layer3_outputs(6828) <= not((layer2_outputs(4279)) and (layer2_outputs(1162)));
    layer3_outputs(6829) <= (layer2_outputs(5985)) or (layer2_outputs(6093));
    layer3_outputs(6830) <= not(layer2_outputs(3197));
    layer3_outputs(6831) <= (layer2_outputs(254)) and not (layer2_outputs(2042));
    layer3_outputs(6832) <= not((layer2_outputs(5604)) or (layer2_outputs(2732)));
    layer3_outputs(6833) <= not(layer2_outputs(5910));
    layer3_outputs(6834) <= not(layer2_outputs(575));
    layer3_outputs(6835) <= not(layer2_outputs(5481));
    layer3_outputs(6836) <= not(layer2_outputs(6753));
    layer3_outputs(6837) <= (layer2_outputs(758)) and (layer2_outputs(3306));
    layer3_outputs(6838) <= (layer2_outputs(7281)) or (layer2_outputs(235));
    layer3_outputs(6839) <= not(layer2_outputs(3268));
    layer3_outputs(6840) <= not(layer2_outputs(3649)) or (layer2_outputs(702));
    layer3_outputs(6841) <= (layer2_outputs(3574)) and (layer2_outputs(313));
    layer3_outputs(6842) <= not(layer2_outputs(1751));
    layer3_outputs(6843) <= not(layer2_outputs(4702));
    layer3_outputs(6844) <= not(layer2_outputs(1935));
    layer3_outputs(6845) <= (layer2_outputs(3050)) and not (layer2_outputs(4889));
    layer3_outputs(6846) <= (layer2_outputs(1720)) and (layer2_outputs(13));
    layer3_outputs(6847) <= (layer2_outputs(3938)) and not (layer2_outputs(3832));
    layer3_outputs(6848) <= not(layer2_outputs(2689)) or (layer2_outputs(4160));
    layer3_outputs(6849) <= layer2_outputs(5872);
    layer3_outputs(6850) <= not((layer2_outputs(6665)) and (layer2_outputs(6317)));
    layer3_outputs(6851) <= (layer2_outputs(519)) and (layer2_outputs(1749));
    layer3_outputs(6852) <= not((layer2_outputs(3648)) xor (layer2_outputs(1510)));
    layer3_outputs(6853) <= layer2_outputs(2318);
    layer3_outputs(6854) <= not(layer2_outputs(2382));
    layer3_outputs(6855) <= not((layer2_outputs(5220)) xor (layer2_outputs(513)));
    layer3_outputs(6856) <= not((layer2_outputs(1033)) or (layer2_outputs(2765)));
    layer3_outputs(6857) <= layer2_outputs(395);
    layer3_outputs(6858) <= (layer2_outputs(3790)) and (layer2_outputs(5662));
    layer3_outputs(6859) <= not((layer2_outputs(2768)) or (layer2_outputs(910)));
    layer3_outputs(6860) <= layer2_outputs(6679);
    layer3_outputs(6861) <= not(layer2_outputs(1406)) or (layer2_outputs(6321));
    layer3_outputs(6862) <= not(layer2_outputs(7145));
    layer3_outputs(6863) <= (layer2_outputs(4014)) and not (layer2_outputs(899));
    layer3_outputs(6864) <= (layer2_outputs(4945)) and not (layer2_outputs(3316));
    layer3_outputs(6865) <= not(layer2_outputs(6262));
    layer3_outputs(6866) <= (layer2_outputs(6772)) xor (layer2_outputs(2907));
    layer3_outputs(6867) <= not(layer2_outputs(6323));
    layer3_outputs(6868) <= layer2_outputs(6402);
    layer3_outputs(6869) <= not(layer2_outputs(2660)) or (layer2_outputs(3878));
    layer3_outputs(6870) <= (layer2_outputs(7497)) and not (layer2_outputs(4497));
    layer3_outputs(6871) <= not((layer2_outputs(2988)) xor (layer2_outputs(1910)));
    layer3_outputs(6872) <= not((layer2_outputs(3655)) and (layer2_outputs(740)));
    layer3_outputs(6873) <= layer2_outputs(1608);
    layer3_outputs(6874) <= (layer2_outputs(2586)) and not (layer2_outputs(3716));
    layer3_outputs(6875) <= not(layer2_outputs(5728));
    layer3_outputs(6876) <= (layer2_outputs(442)) and (layer2_outputs(5991));
    layer3_outputs(6877) <= (layer2_outputs(3814)) or (layer2_outputs(2128));
    layer3_outputs(6878) <= not(layer2_outputs(6584));
    layer3_outputs(6879) <= layer2_outputs(1163);
    layer3_outputs(6880) <= (layer2_outputs(3814)) and not (layer2_outputs(1733));
    layer3_outputs(6881) <= layer2_outputs(6096);
    layer3_outputs(6882) <= not(layer2_outputs(1384));
    layer3_outputs(6883) <= (layer2_outputs(7339)) and not (layer2_outputs(2667));
    layer3_outputs(6884) <= layer2_outputs(2357);
    layer3_outputs(6885) <= not(layer2_outputs(3796));
    layer3_outputs(6886) <= not(layer2_outputs(6451));
    layer3_outputs(6887) <= not(layer2_outputs(3539));
    layer3_outputs(6888) <= not(layer2_outputs(3933));
    layer3_outputs(6889) <= layer2_outputs(3906);
    layer3_outputs(6890) <= layer2_outputs(3383);
    layer3_outputs(6891) <= layer2_outputs(794);
    layer3_outputs(6892) <= not(layer2_outputs(6212));
    layer3_outputs(6893) <= not(layer2_outputs(5641));
    layer3_outputs(6894) <= layer2_outputs(2261);
    layer3_outputs(6895) <= not(layer2_outputs(4216)) or (layer2_outputs(5298));
    layer3_outputs(6896) <= (layer2_outputs(3375)) and (layer2_outputs(7054));
    layer3_outputs(6897) <= (layer2_outputs(7196)) and not (layer2_outputs(7181));
    layer3_outputs(6898) <= (layer2_outputs(2057)) xor (layer2_outputs(6147));
    layer3_outputs(6899) <= not((layer2_outputs(7066)) and (layer2_outputs(571)));
    layer3_outputs(6900) <= not((layer2_outputs(3961)) and (layer2_outputs(1064)));
    layer3_outputs(6901) <= (layer2_outputs(7590)) and not (layer2_outputs(1669));
    layer3_outputs(6902) <= layer2_outputs(1189);
    layer3_outputs(6903) <= (layer2_outputs(6079)) xor (layer2_outputs(6916));
    layer3_outputs(6904) <= not(layer2_outputs(5087));
    layer3_outputs(6905) <= not(layer2_outputs(2744));
    layer3_outputs(6906) <= not(layer2_outputs(5160));
    layer3_outputs(6907) <= (layer2_outputs(5427)) and (layer2_outputs(3420));
    layer3_outputs(6908) <= not(layer2_outputs(25));
    layer3_outputs(6909) <= not(layer2_outputs(1394));
    layer3_outputs(6910) <= layer2_outputs(7541);
    layer3_outputs(6911) <= (layer2_outputs(6000)) and not (layer2_outputs(171));
    layer3_outputs(6912) <= layer2_outputs(85);
    layer3_outputs(6913) <= layer2_outputs(6121);
    layer3_outputs(6914) <= not(layer2_outputs(7314));
    layer3_outputs(6915) <= (layer2_outputs(3386)) and not (layer2_outputs(1480));
    layer3_outputs(6916) <= not(layer2_outputs(10));
    layer3_outputs(6917) <= not(layer2_outputs(6957)) or (layer2_outputs(2471));
    layer3_outputs(6918) <= not((layer2_outputs(440)) or (layer2_outputs(1833)));
    layer3_outputs(6919) <= (layer2_outputs(2602)) and not (layer2_outputs(5403));
    layer3_outputs(6920) <= layer2_outputs(4035);
    layer3_outputs(6921) <= not(layer2_outputs(6879));
    layer3_outputs(6922) <= (layer2_outputs(297)) xor (layer2_outputs(7089));
    layer3_outputs(6923) <= not(layer2_outputs(1190));
    layer3_outputs(6924) <= not((layer2_outputs(799)) or (layer2_outputs(581)));
    layer3_outputs(6925) <= not(layer2_outputs(6212)) or (layer2_outputs(5892));
    layer3_outputs(6926) <= not((layer2_outputs(3427)) xor (layer2_outputs(6633)));
    layer3_outputs(6927) <= not(layer2_outputs(3906));
    layer3_outputs(6928) <= not(layer2_outputs(1844));
    layer3_outputs(6929) <= not((layer2_outputs(6309)) xor (layer2_outputs(2286)));
    layer3_outputs(6930) <= not(layer2_outputs(4304)) or (layer2_outputs(4999));
    layer3_outputs(6931) <= not((layer2_outputs(7649)) xor (layer2_outputs(469)));
    layer3_outputs(6932) <= not(layer2_outputs(2835)) or (layer2_outputs(6551));
    layer3_outputs(6933) <= (layer2_outputs(5645)) and not (layer2_outputs(6845));
    layer3_outputs(6934) <= layer2_outputs(765);
    layer3_outputs(6935) <= not(layer2_outputs(2555)) or (layer2_outputs(964));
    layer3_outputs(6936) <= not(layer2_outputs(5234)) or (layer2_outputs(1489));
    layer3_outputs(6937) <= not(layer2_outputs(4364));
    layer3_outputs(6938) <= (layer2_outputs(1561)) and (layer2_outputs(2092));
    layer3_outputs(6939) <= not(layer2_outputs(2878));
    layer3_outputs(6940) <= not(layer2_outputs(7305));
    layer3_outputs(6941) <= layer2_outputs(7662);
    layer3_outputs(6942) <= layer2_outputs(4233);
    layer3_outputs(6943) <= not((layer2_outputs(2834)) or (layer2_outputs(5225)));
    layer3_outputs(6944) <= not(layer2_outputs(46));
    layer3_outputs(6945) <= not(layer2_outputs(310));
    layer3_outputs(6946) <= not(layer2_outputs(5515));
    layer3_outputs(6947) <= not(layer2_outputs(4001));
    layer3_outputs(6948) <= not(layer2_outputs(7423)) or (layer2_outputs(1383));
    layer3_outputs(6949) <= (layer2_outputs(7030)) and (layer2_outputs(7025));
    layer3_outputs(6950) <= not(layer2_outputs(6499));
    layer3_outputs(6951) <= (layer2_outputs(6197)) and not (layer2_outputs(1633));
    layer3_outputs(6952) <= (layer2_outputs(289)) and (layer2_outputs(379));
    layer3_outputs(6953) <= not(layer2_outputs(5297));
    layer3_outputs(6954) <= not((layer2_outputs(2690)) and (layer2_outputs(287)));
    layer3_outputs(6955) <= not(layer2_outputs(2566)) or (layer2_outputs(1590));
    layer3_outputs(6956) <= layer2_outputs(1044);
    layer3_outputs(6957) <= not((layer2_outputs(3229)) or (layer2_outputs(5801)));
    layer3_outputs(6958) <= '0';
    layer3_outputs(6959) <= not(layer2_outputs(7086));
    layer3_outputs(6960) <= layer2_outputs(4460);
    layer3_outputs(6961) <= (layer2_outputs(5423)) xor (layer2_outputs(586));
    layer3_outputs(6962) <= '0';
    layer3_outputs(6963) <= (layer2_outputs(5228)) xor (layer2_outputs(2874));
    layer3_outputs(6964) <= layer2_outputs(7065);
    layer3_outputs(6965) <= not((layer2_outputs(750)) xor (layer2_outputs(2662)));
    layer3_outputs(6966) <= (layer2_outputs(5190)) and (layer2_outputs(2273));
    layer3_outputs(6967) <= not(layer2_outputs(3283));
    layer3_outputs(6968) <= not(layer2_outputs(1042)) or (layer2_outputs(675));
    layer3_outputs(6969) <= not(layer2_outputs(3750));
    layer3_outputs(6970) <= (layer2_outputs(1786)) and (layer2_outputs(2342));
    layer3_outputs(6971) <= (layer2_outputs(4626)) or (layer2_outputs(3261));
    layer3_outputs(6972) <= (layer2_outputs(2083)) and not (layer2_outputs(1141));
    layer3_outputs(6973) <= not((layer2_outputs(3705)) and (layer2_outputs(4711)));
    layer3_outputs(6974) <= not(layer2_outputs(4280));
    layer3_outputs(6975) <= (layer2_outputs(1814)) xor (layer2_outputs(3827));
    layer3_outputs(6976) <= '1';
    layer3_outputs(6977) <= not((layer2_outputs(156)) and (layer2_outputs(4205)));
    layer3_outputs(6978) <= (layer2_outputs(6842)) or (layer2_outputs(4459));
    layer3_outputs(6979) <= layer2_outputs(7645);
    layer3_outputs(6980) <= not(layer2_outputs(2556));
    layer3_outputs(6981) <= not(layer2_outputs(2608)) or (layer2_outputs(3876));
    layer3_outputs(6982) <= layer2_outputs(5790);
    layer3_outputs(6983) <= not(layer2_outputs(4743));
    layer3_outputs(6984) <= (layer2_outputs(7112)) and not (layer2_outputs(5869));
    layer3_outputs(6985) <= not((layer2_outputs(3588)) xor (layer2_outputs(1494)));
    layer3_outputs(6986) <= (layer2_outputs(3982)) and not (layer2_outputs(1938));
    layer3_outputs(6987) <= layer2_outputs(1420);
    layer3_outputs(6988) <= not(layer2_outputs(1502));
    layer3_outputs(6989) <= not(layer2_outputs(3017));
    layer3_outputs(6990) <= (layer2_outputs(2115)) or (layer2_outputs(7242));
    layer3_outputs(6991) <= layer2_outputs(2447);
    layer3_outputs(6992) <= not((layer2_outputs(5058)) and (layer2_outputs(2068)));
    layer3_outputs(6993) <= (layer2_outputs(7472)) xor (layer2_outputs(3128));
    layer3_outputs(6994) <= (layer2_outputs(1043)) and not (layer2_outputs(7507));
    layer3_outputs(6995) <= not((layer2_outputs(4499)) xor (layer2_outputs(5522)));
    layer3_outputs(6996) <= not(layer2_outputs(2072)) or (layer2_outputs(6015));
    layer3_outputs(6997) <= not(layer2_outputs(2348));
    layer3_outputs(6998) <= (layer2_outputs(362)) and (layer2_outputs(5837));
    layer3_outputs(6999) <= layer2_outputs(3287);
    layer3_outputs(7000) <= (layer2_outputs(7592)) and not (layer2_outputs(1575));
    layer3_outputs(7001) <= (layer2_outputs(4567)) and not (layer2_outputs(7565));
    layer3_outputs(7002) <= not(layer2_outputs(3324));
    layer3_outputs(7003) <= layer2_outputs(5266);
    layer3_outputs(7004) <= layer2_outputs(5820);
    layer3_outputs(7005) <= '0';
    layer3_outputs(7006) <= not(layer2_outputs(2474));
    layer3_outputs(7007) <= not(layer2_outputs(932)) or (layer2_outputs(3397));
    layer3_outputs(7008) <= not(layer2_outputs(4356));
    layer3_outputs(7009) <= (layer2_outputs(889)) and not (layer2_outputs(2710));
    layer3_outputs(7010) <= layer2_outputs(5881);
    layer3_outputs(7011) <= (layer2_outputs(1906)) xor (layer2_outputs(6884));
    layer3_outputs(7012) <= (layer2_outputs(1508)) and (layer2_outputs(3343));
    layer3_outputs(7013) <= not(layer2_outputs(2508));
    layer3_outputs(7014) <= (layer2_outputs(4009)) or (layer2_outputs(7008));
    layer3_outputs(7015) <= '0';
    layer3_outputs(7016) <= not(layer2_outputs(3458));
    layer3_outputs(7017) <= not((layer2_outputs(4122)) and (layer2_outputs(469)));
    layer3_outputs(7018) <= (layer2_outputs(1895)) or (layer2_outputs(111));
    layer3_outputs(7019) <= not(layer2_outputs(3801));
    layer3_outputs(7020) <= not(layer2_outputs(5958));
    layer3_outputs(7021) <= layer2_outputs(5761);
    layer3_outputs(7022) <= not((layer2_outputs(2248)) or (layer2_outputs(1068)));
    layer3_outputs(7023) <= not(layer2_outputs(199));
    layer3_outputs(7024) <= (layer2_outputs(407)) and not (layer2_outputs(566));
    layer3_outputs(7025) <= not(layer2_outputs(1237)) or (layer2_outputs(7039));
    layer3_outputs(7026) <= layer2_outputs(2410);
    layer3_outputs(7027) <= '1';
    layer3_outputs(7028) <= (layer2_outputs(2540)) and not (layer2_outputs(760));
    layer3_outputs(7029) <= (layer2_outputs(5659)) and (layer2_outputs(905));
    layer3_outputs(7030) <= (layer2_outputs(6218)) xor (layer2_outputs(2365));
    layer3_outputs(7031) <= (layer2_outputs(2898)) or (layer2_outputs(5938));
    layer3_outputs(7032) <= not(layer2_outputs(6827));
    layer3_outputs(7033) <= not((layer2_outputs(7110)) or (layer2_outputs(1290)));
    layer3_outputs(7034) <= (layer2_outputs(5960)) xor (layer2_outputs(6394));
    layer3_outputs(7035) <= (layer2_outputs(2550)) and not (layer2_outputs(38));
    layer3_outputs(7036) <= not(layer2_outputs(2093)) or (layer2_outputs(3034));
    layer3_outputs(7037) <= not(layer2_outputs(4389));
    layer3_outputs(7038) <= layer2_outputs(2264);
    layer3_outputs(7039) <= layer2_outputs(6834);
    layer3_outputs(7040) <= layer2_outputs(6627);
    layer3_outputs(7041) <= not(layer2_outputs(5081)) or (layer2_outputs(479));
    layer3_outputs(7042) <= not(layer2_outputs(2433)) or (layer2_outputs(4066));
    layer3_outputs(7043) <= not((layer2_outputs(5543)) or (layer2_outputs(5779)));
    layer3_outputs(7044) <= not((layer2_outputs(2142)) or (layer2_outputs(4718)));
    layer3_outputs(7045) <= '0';
    layer3_outputs(7046) <= (layer2_outputs(7034)) and not (layer2_outputs(5852));
    layer3_outputs(7047) <= (layer2_outputs(2342)) or (layer2_outputs(3816));
    layer3_outputs(7048) <= not(layer2_outputs(6609));
    layer3_outputs(7049) <= not(layer2_outputs(6803));
    layer3_outputs(7050) <= '1';
    layer3_outputs(7051) <= layer2_outputs(880);
    layer3_outputs(7052) <= layer2_outputs(6362);
    layer3_outputs(7053) <= not((layer2_outputs(1374)) or (layer2_outputs(6611)));
    layer3_outputs(7054) <= not(layer2_outputs(7391));
    layer3_outputs(7055) <= (layer2_outputs(5617)) and not (layer2_outputs(5163));
    layer3_outputs(7056) <= '0';
    layer3_outputs(7057) <= not(layer2_outputs(684));
    layer3_outputs(7058) <= not((layer2_outputs(253)) or (layer2_outputs(2741)));
    layer3_outputs(7059) <= (layer2_outputs(4411)) and (layer2_outputs(2626));
    layer3_outputs(7060) <= layer2_outputs(5136);
    layer3_outputs(7061) <= (layer2_outputs(3882)) and not (layer2_outputs(89));
    layer3_outputs(7062) <= not(layer2_outputs(5149));
    layer3_outputs(7063) <= not(layer2_outputs(3972));
    layer3_outputs(7064) <= (layer2_outputs(1911)) xor (layer2_outputs(4617));
    layer3_outputs(7065) <= (layer2_outputs(6899)) or (layer2_outputs(1230));
    layer3_outputs(7066) <= (layer2_outputs(6690)) and (layer2_outputs(503));
    layer3_outputs(7067) <= not((layer2_outputs(5469)) and (layer2_outputs(5749)));
    layer3_outputs(7068) <= not((layer2_outputs(2466)) or (layer2_outputs(7087)));
    layer3_outputs(7069) <= layer2_outputs(4697);
    layer3_outputs(7070) <= (layer2_outputs(2750)) and not (layer2_outputs(1997));
    layer3_outputs(7071) <= layer2_outputs(5011);
    layer3_outputs(7072) <= not(layer2_outputs(1001)) or (layer2_outputs(5804));
    layer3_outputs(7073) <= (layer2_outputs(381)) xor (layer2_outputs(7164));
    layer3_outputs(7074) <= '0';
    layer3_outputs(7075) <= layer2_outputs(1312);
    layer3_outputs(7076) <= not(layer2_outputs(6575)) or (layer2_outputs(1082));
    layer3_outputs(7077) <= not(layer2_outputs(2505));
    layer3_outputs(7078) <= not((layer2_outputs(6079)) and (layer2_outputs(2437)));
    layer3_outputs(7079) <= layer2_outputs(3786);
    layer3_outputs(7080) <= not((layer2_outputs(262)) or (layer2_outputs(1701)));
    layer3_outputs(7081) <= layer2_outputs(1479);
    layer3_outputs(7082) <= layer2_outputs(2833);
    layer3_outputs(7083) <= not((layer2_outputs(6932)) or (layer2_outputs(2953)));
    layer3_outputs(7084) <= not((layer2_outputs(117)) and (layer2_outputs(5122)));
    layer3_outputs(7085) <= (layer2_outputs(4751)) and not (layer2_outputs(867));
    layer3_outputs(7086) <= layer2_outputs(5003);
    layer3_outputs(7087) <= not((layer2_outputs(6325)) and (layer2_outputs(2439)));
    layer3_outputs(7088) <= not(layer2_outputs(2124)) or (layer2_outputs(3232));
    layer3_outputs(7089) <= (layer2_outputs(4413)) and (layer2_outputs(3036));
    layer3_outputs(7090) <= not(layer2_outputs(5393));
    layer3_outputs(7091) <= (layer2_outputs(4186)) and (layer2_outputs(6157));
    layer3_outputs(7092) <= not(layer2_outputs(7166)) or (layer2_outputs(5482));
    layer3_outputs(7093) <= not((layer2_outputs(506)) and (layer2_outputs(5840)));
    layer3_outputs(7094) <= not(layer2_outputs(7146));
    layer3_outputs(7095) <= not(layer2_outputs(5901)) or (layer2_outputs(3480));
    layer3_outputs(7096) <= not(layer2_outputs(834));
    layer3_outputs(7097) <= (layer2_outputs(3278)) or (layer2_outputs(3534));
    layer3_outputs(7098) <= layer2_outputs(5736);
    layer3_outputs(7099) <= not(layer2_outputs(2305));
    layer3_outputs(7100) <= (layer2_outputs(4677)) and (layer2_outputs(4247));
    layer3_outputs(7101) <= layer2_outputs(3350);
    layer3_outputs(7102) <= not(layer2_outputs(267));
    layer3_outputs(7103) <= (layer2_outputs(7606)) and not (layer2_outputs(2131));
    layer3_outputs(7104) <= not((layer2_outputs(1597)) and (layer2_outputs(786)));
    layer3_outputs(7105) <= not((layer2_outputs(3380)) and (layer2_outputs(583)));
    layer3_outputs(7106) <= not((layer2_outputs(4923)) or (layer2_outputs(437)));
    layer3_outputs(7107) <= (layer2_outputs(1501)) and not (layer2_outputs(1954));
    layer3_outputs(7108) <= not((layer2_outputs(1127)) or (layer2_outputs(7336)));
    layer3_outputs(7109) <= (layer2_outputs(5152)) or (layer2_outputs(1341));
    layer3_outputs(7110) <= not(layer2_outputs(4225));
    layer3_outputs(7111) <= layer2_outputs(1360);
    layer3_outputs(7112) <= (layer2_outputs(3981)) and (layer2_outputs(4640));
    layer3_outputs(7113) <= not(layer2_outputs(6707));
    layer3_outputs(7114) <= (layer2_outputs(5456)) xor (layer2_outputs(4024));
    layer3_outputs(7115) <= (layer2_outputs(1241)) and (layer2_outputs(5028));
    layer3_outputs(7116) <= layer2_outputs(5764);
    layer3_outputs(7117) <= layer2_outputs(6177);
    layer3_outputs(7118) <= layer2_outputs(5741);
    layer3_outputs(7119) <= layer2_outputs(4729);
    layer3_outputs(7120) <= layer2_outputs(7358);
    layer3_outputs(7121) <= (layer2_outputs(4413)) or (layer2_outputs(6581));
    layer3_outputs(7122) <= not((layer2_outputs(1603)) or (layer2_outputs(7612)));
    layer3_outputs(7123) <= (layer2_outputs(827)) or (layer2_outputs(1510));
    layer3_outputs(7124) <= layer2_outputs(5364);
    layer3_outputs(7125) <= (layer2_outputs(1228)) and not (layer2_outputs(2311));
    layer3_outputs(7126) <= (layer2_outputs(7505)) or (layer2_outputs(575));
    layer3_outputs(7127) <= layer2_outputs(5360);
    layer3_outputs(7128) <= not(layer2_outputs(5899));
    layer3_outputs(7129) <= not(layer2_outputs(154));
    layer3_outputs(7130) <= (layer2_outputs(1635)) and not (layer2_outputs(4082));
    layer3_outputs(7131) <= (layer2_outputs(7292)) and (layer2_outputs(1473));
    layer3_outputs(7132) <= layer2_outputs(815);
    layer3_outputs(7133) <= (layer2_outputs(1187)) and (layer2_outputs(1530));
    layer3_outputs(7134) <= not(layer2_outputs(1392));
    layer3_outputs(7135) <= not(layer2_outputs(5956)) or (layer2_outputs(6277));
    layer3_outputs(7136) <= not((layer2_outputs(4143)) or (layer2_outputs(4259)));
    layer3_outputs(7137) <= not(layer2_outputs(5556));
    layer3_outputs(7138) <= (layer2_outputs(1061)) and (layer2_outputs(3640));
    layer3_outputs(7139) <= (layer2_outputs(2499)) or (layer2_outputs(1978));
    layer3_outputs(7140) <= (layer2_outputs(5026)) xor (layer2_outputs(5521));
    layer3_outputs(7141) <= not(layer2_outputs(7386));
    layer3_outputs(7142) <= not(layer2_outputs(7108));
    layer3_outputs(7143) <= not(layer2_outputs(3675)) or (layer2_outputs(7134));
    layer3_outputs(7144) <= layer2_outputs(2106);
    layer3_outputs(7145) <= not(layer2_outputs(7586)) or (layer2_outputs(4481));
    layer3_outputs(7146) <= not(layer2_outputs(3647)) or (layer2_outputs(2456));
    layer3_outputs(7147) <= not(layer2_outputs(1558)) or (layer2_outputs(4237));
    layer3_outputs(7148) <= not(layer2_outputs(6527)) or (layer2_outputs(1487));
    layer3_outputs(7149) <= layer2_outputs(6570);
    layer3_outputs(7150) <= (layer2_outputs(526)) and (layer2_outputs(6477));
    layer3_outputs(7151) <= not(layer2_outputs(1886));
    layer3_outputs(7152) <= (layer2_outputs(1072)) xor (layer2_outputs(6771));
    layer3_outputs(7153) <= layer2_outputs(1614);
    layer3_outputs(7154) <= layer2_outputs(1397);
    layer3_outputs(7155) <= not(layer2_outputs(5292));
    layer3_outputs(7156) <= '0';
    layer3_outputs(7157) <= (layer2_outputs(4800)) or (layer2_outputs(2918));
    layer3_outputs(7158) <= not((layer2_outputs(4556)) xor (layer2_outputs(6948)));
    layer3_outputs(7159) <= layer2_outputs(6945);
    layer3_outputs(7160) <= layer2_outputs(451);
    layer3_outputs(7161) <= (layer2_outputs(5922)) or (layer2_outputs(6258));
    layer3_outputs(7162) <= layer2_outputs(4061);
    layer3_outputs(7163) <= not(layer2_outputs(4892));
    layer3_outputs(7164) <= (layer2_outputs(4028)) and not (layer2_outputs(357));
    layer3_outputs(7165) <= layer2_outputs(5167);
    layer3_outputs(7166) <= layer2_outputs(4150);
    layer3_outputs(7167) <= (layer2_outputs(5437)) and (layer2_outputs(2555));
    layer3_outputs(7168) <= not((layer2_outputs(529)) xor (layer2_outputs(1918)));
    layer3_outputs(7169) <= layer2_outputs(5502);
    layer3_outputs(7170) <= not(layer2_outputs(118)) or (layer2_outputs(490));
    layer3_outputs(7171) <= (layer2_outputs(2178)) and (layer2_outputs(1247));
    layer3_outputs(7172) <= layer2_outputs(2462);
    layer3_outputs(7173) <= not(layer2_outputs(141));
    layer3_outputs(7174) <= (layer2_outputs(5080)) and not (layer2_outputs(4319));
    layer3_outputs(7175) <= not(layer2_outputs(7276));
    layer3_outputs(7176) <= not((layer2_outputs(7672)) and (layer2_outputs(4807)));
    layer3_outputs(7177) <= layer2_outputs(4436);
    layer3_outputs(7178) <= (layer2_outputs(1621)) and not (layer2_outputs(4770));
    layer3_outputs(7179) <= (layer2_outputs(7538)) and (layer2_outputs(6054));
    layer3_outputs(7180) <= not(layer2_outputs(2245));
    layer3_outputs(7181) <= layer2_outputs(394);
    layer3_outputs(7182) <= layer2_outputs(6005);
    layer3_outputs(7183) <= (layer2_outputs(5826)) and not (layer2_outputs(5114));
    layer3_outputs(7184) <= (layer2_outputs(1941)) xor (layer2_outputs(5987));
    layer3_outputs(7185) <= '1';
    layer3_outputs(7186) <= not(layer2_outputs(1100));
    layer3_outputs(7187) <= not((layer2_outputs(2933)) xor (layer2_outputs(5336)));
    layer3_outputs(7188) <= (layer2_outputs(6848)) or (layer2_outputs(7508));
    layer3_outputs(7189) <= not(layer2_outputs(4850));
    layer3_outputs(7190) <= (layer2_outputs(5544)) xor (layer2_outputs(1853));
    layer3_outputs(7191) <= not(layer2_outputs(6893)) or (layer2_outputs(6303));
    layer3_outputs(7192) <= layer2_outputs(4944);
    layer3_outputs(7193) <= not(layer2_outputs(1511));
    layer3_outputs(7194) <= layer2_outputs(2108);
    layer3_outputs(7195) <= not(layer2_outputs(7513));
    layer3_outputs(7196) <= (layer2_outputs(2268)) and not (layer2_outputs(5551));
    layer3_outputs(7197) <= not(layer2_outputs(4548));
    layer3_outputs(7198) <= layer2_outputs(1600);
    layer3_outputs(7199) <= not(layer2_outputs(1866));
    layer3_outputs(7200) <= not(layer2_outputs(1838));
    layer3_outputs(7201) <= layer2_outputs(3047);
    layer3_outputs(7202) <= not(layer2_outputs(4888));
    layer3_outputs(7203) <= layer2_outputs(5504);
    layer3_outputs(7204) <= layer2_outputs(6780);
    layer3_outputs(7205) <= (layer2_outputs(5705)) or (layer2_outputs(5690));
    layer3_outputs(7206) <= not(layer2_outputs(1523)) or (layer2_outputs(4231));
    layer3_outputs(7207) <= not(layer2_outputs(6322)) or (layer2_outputs(3602));
    layer3_outputs(7208) <= not(layer2_outputs(1324)) or (layer2_outputs(4473));
    layer3_outputs(7209) <= not(layer2_outputs(5018));
    layer3_outputs(7210) <= (layer2_outputs(5227)) and not (layer2_outputs(3867));
    layer3_outputs(7211) <= not(layer2_outputs(6121));
    layer3_outputs(7212) <= not(layer2_outputs(559));
    layer3_outputs(7213) <= not(layer2_outputs(3862));
    layer3_outputs(7214) <= not(layer2_outputs(822));
    layer3_outputs(7215) <= not(layer2_outputs(7462));
    layer3_outputs(7216) <= not(layer2_outputs(6583));
    layer3_outputs(7217) <= (layer2_outputs(2666)) and not (layer2_outputs(6641));
    layer3_outputs(7218) <= not(layer2_outputs(7674));
    layer3_outputs(7219) <= layer2_outputs(288);
    layer3_outputs(7220) <= '1';
    layer3_outputs(7221) <= not((layer2_outputs(3740)) and (layer2_outputs(3212)));
    layer3_outputs(7222) <= (layer2_outputs(295)) and (layer2_outputs(7211));
    layer3_outputs(7223) <= not(layer2_outputs(7216));
    layer3_outputs(7224) <= not(layer2_outputs(1416)) or (layer2_outputs(7070));
    layer3_outputs(7225) <= layer2_outputs(5017);
    layer3_outputs(7226) <= not(layer2_outputs(400));
    layer3_outputs(7227) <= not(layer2_outputs(824));
    layer3_outputs(7228) <= not(layer2_outputs(4766));
    layer3_outputs(7229) <= layer2_outputs(170);
    layer3_outputs(7230) <= not((layer2_outputs(5692)) or (layer2_outputs(5882)));
    layer3_outputs(7231) <= not(layer2_outputs(3935));
    layer3_outputs(7232) <= not(layer2_outputs(4648));
    layer3_outputs(7233) <= not(layer2_outputs(7366));
    layer3_outputs(7234) <= not((layer2_outputs(3364)) or (layer2_outputs(1327)));
    layer3_outputs(7235) <= not((layer2_outputs(2471)) xor (layer2_outputs(6858)));
    layer3_outputs(7236) <= (layer2_outputs(7309)) or (layer2_outputs(6612));
    layer3_outputs(7237) <= '1';
    layer3_outputs(7238) <= not(layer2_outputs(6543));
    layer3_outputs(7239) <= not((layer2_outputs(6297)) or (layer2_outputs(5738)));
    layer3_outputs(7240) <= (layer2_outputs(4632)) and (layer2_outputs(7351));
    layer3_outputs(7241) <= (layer2_outputs(2989)) and not (layer2_outputs(6195));
    layer3_outputs(7242) <= not((layer2_outputs(3392)) or (layer2_outputs(1402)));
    layer3_outputs(7243) <= (layer2_outputs(677)) and (layer2_outputs(4517));
    layer3_outputs(7244) <= not(layer2_outputs(6115));
    layer3_outputs(7245) <= (layer2_outputs(5601)) and not (layer2_outputs(3615));
    layer3_outputs(7246) <= not(layer2_outputs(728)) or (layer2_outputs(4291));
    layer3_outputs(7247) <= not(layer2_outputs(982));
    layer3_outputs(7248) <= not(layer2_outputs(3451));
    layer3_outputs(7249) <= not((layer2_outputs(6577)) or (layer2_outputs(3836)));
    layer3_outputs(7250) <= not(layer2_outputs(5525)) or (layer2_outputs(5537));
    layer3_outputs(7251) <= (layer2_outputs(6895)) and not (layer2_outputs(4974));
    layer3_outputs(7252) <= (layer2_outputs(2718)) and (layer2_outputs(4708));
    layer3_outputs(7253) <= not((layer2_outputs(1661)) and (layer2_outputs(537)));
    layer3_outputs(7254) <= layer2_outputs(3135);
    layer3_outputs(7255) <= not(layer2_outputs(6066));
    layer3_outputs(7256) <= not(layer2_outputs(3039));
    layer3_outputs(7257) <= not(layer2_outputs(7478));
    layer3_outputs(7258) <= not(layer2_outputs(1512));
    layer3_outputs(7259) <= not((layer2_outputs(1892)) and (layer2_outputs(4785)));
    layer3_outputs(7260) <= not(layer2_outputs(4608));
    layer3_outputs(7261) <= (layer2_outputs(5640)) and (layer2_outputs(6656));
    layer3_outputs(7262) <= layer2_outputs(1121);
    layer3_outputs(7263) <= not(layer2_outputs(6685));
    layer3_outputs(7264) <= (layer2_outputs(4447)) and (layer2_outputs(278));
    layer3_outputs(7265) <= (layer2_outputs(5500)) xor (layer2_outputs(7325));
    layer3_outputs(7266) <= (layer2_outputs(5770)) and not (layer2_outputs(4672));
    layer3_outputs(7267) <= not(layer2_outputs(7563));
    layer3_outputs(7268) <= '0';
    layer3_outputs(7269) <= layer2_outputs(4090);
    layer3_outputs(7270) <= not(layer2_outputs(4836)) or (layer2_outputs(6315));
    layer3_outputs(7271) <= layer2_outputs(4398);
    layer3_outputs(7272) <= (layer2_outputs(2760)) and (layer2_outputs(6548));
    layer3_outputs(7273) <= not((layer2_outputs(5448)) or (layer2_outputs(1407)));
    layer3_outputs(7274) <= (layer2_outputs(6718)) xor (layer2_outputs(1697));
    layer3_outputs(7275) <= not(layer2_outputs(3352)) or (layer2_outputs(2896));
    layer3_outputs(7276) <= '1';
    layer3_outputs(7277) <= layer2_outputs(7421);
    layer3_outputs(7278) <= not(layer2_outputs(7527)) or (layer2_outputs(395));
    layer3_outputs(7279) <= not(layer2_outputs(5568));
    layer3_outputs(7280) <= not(layer2_outputs(4494));
    layer3_outputs(7281) <= layer2_outputs(3083);
    layer3_outputs(7282) <= layer2_outputs(1008);
    layer3_outputs(7283) <= not(layer2_outputs(4504));
    layer3_outputs(7284) <= not(layer2_outputs(492)) or (layer2_outputs(3988));
    layer3_outputs(7285) <= layer2_outputs(4802);
    layer3_outputs(7286) <= not((layer2_outputs(222)) or (layer2_outputs(2064)));
    layer3_outputs(7287) <= not(layer2_outputs(2082));
    layer3_outputs(7288) <= layer2_outputs(3931);
    layer3_outputs(7289) <= not(layer2_outputs(2532));
    layer3_outputs(7290) <= (layer2_outputs(18)) and not (layer2_outputs(2101));
    layer3_outputs(7291) <= (layer2_outputs(6668)) and (layer2_outputs(2387));
    layer3_outputs(7292) <= '1';
    layer3_outputs(7293) <= not((layer2_outputs(3051)) and (layer2_outputs(3358)));
    layer3_outputs(7294) <= layer2_outputs(6998);
    layer3_outputs(7295) <= layer2_outputs(2191);
    layer3_outputs(7296) <= not(layer2_outputs(1262));
    layer3_outputs(7297) <= '1';
    layer3_outputs(7298) <= '0';
    layer3_outputs(7299) <= not(layer2_outputs(5555)) or (layer2_outputs(7279));
    layer3_outputs(7300) <= not((layer2_outputs(4068)) or (layer2_outputs(3258)));
    layer3_outputs(7301) <= not(layer2_outputs(3100));
    layer3_outputs(7302) <= not(layer2_outputs(1810));
    layer3_outputs(7303) <= not(layer2_outputs(6179));
    layer3_outputs(7304) <= not((layer2_outputs(3908)) and (layer2_outputs(6082)));
    layer3_outputs(7305) <= layer2_outputs(166);
    layer3_outputs(7306) <= not(layer2_outputs(4794)) or (layer2_outputs(4776));
    layer3_outputs(7307) <= layer2_outputs(2971);
    layer3_outputs(7308) <= not(layer2_outputs(6487));
    layer3_outputs(7309) <= not((layer2_outputs(966)) and (layer2_outputs(3556)));
    layer3_outputs(7310) <= not(layer2_outputs(6224));
    layer3_outputs(7311) <= (layer2_outputs(3710)) and not (layer2_outputs(2282));
    layer3_outputs(7312) <= not((layer2_outputs(3589)) and (layer2_outputs(6206)));
    layer3_outputs(7313) <= (layer2_outputs(3632)) and not (layer2_outputs(3490));
    layer3_outputs(7314) <= layer2_outputs(5707);
    layer3_outputs(7315) <= not(layer2_outputs(4084));
    layer3_outputs(7316) <= not(layer2_outputs(3641));
    layer3_outputs(7317) <= layer2_outputs(4193);
    layer3_outputs(7318) <= layer2_outputs(5455);
    layer3_outputs(7319) <= not(layer2_outputs(6804)) or (layer2_outputs(4905));
    layer3_outputs(7320) <= (layer2_outputs(1682)) and (layer2_outputs(3147));
    layer3_outputs(7321) <= (layer2_outputs(1109)) or (layer2_outputs(2040));
    layer3_outputs(7322) <= not((layer2_outputs(2982)) and (layer2_outputs(1060)));
    layer3_outputs(7323) <= not(layer2_outputs(7552));
    layer3_outputs(7324) <= '0';
    layer3_outputs(7325) <= '1';
    layer3_outputs(7326) <= (layer2_outputs(4692)) and not (layer2_outputs(5448));
    layer3_outputs(7327) <= not(layer2_outputs(4338)) or (layer2_outputs(6705));
    layer3_outputs(7328) <= not((layer2_outputs(5222)) and (layer2_outputs(1170)));
    layer3_outputs(7329) <= not(layer2_outputs(1516));
    layer3_outputs(7330) <= not(layer2_outputs(106));
    layer3_outputs(7331) <= not(layer2_outputs(2749));
    layer3_outputs(7332) <= not(layer2_outputs(2347));
    layer3_outputs(7333) <= layer2_outputs(6673);
    layer3_outputs(7334) <= layer2_outputs(6504);
    layer3_outputs(7335) <= (layer2_outputs(4098)) or (layer2_outputs(406));
    layer3_outputs(7336) <= not(layer2_outputs(196));
    layer3_outputs(7337) <= not(layer2_outputs(6492)) or (layer2_outputs(4758));
    layer3_outputs(7338) <= layer2_outputs(1379);
    layer3_outputs(7339) <= not((layer2_outputs(1421)) and (layer2_outputs(6941)));
    layer3_outputs(7340) <= layer2_outputs(2578);
    layer3_outputs(7341) <= (layer2_outputs(2514)) xor (layer2_outputs(7140));
    layer3_outputs(7342) <= layer2_outputs(2921);
    layer3_outputs(7343) <= (layer2_outputs(5671)) or (layer2_outputs(5927));
    layer3_outputs(7344) <= not((layer2_outputs(3227)) or (layer2_outputs(3336)));
    layer3_outputs(7345) <= not(layer2_outputs(4866));
    layer3_outputs(7346) <= not((layer2_outputs(111)) xor (layer2_outputs(1646)));
    layer3_outputs(7347) <= not((layer2_outputs(1564)) and (layer2_outputs(4723)));
    layer3_outputs(7348) <= not(layer2_outputs(4146));
    layer3_outputs(7349) <= layer2_outputs(137);
    layer3_outputs(7350) <= not((layer2_outputs(3853)) and (layer2_outputs(7547)));
    layer3_outputs(7351) <= (layer2_outputs(1347)) and not (layer2_outputs(2468));
    layer3_outputs(7352) <= (layer2_outputs(7416)) and (layer2_outputs(3121));
    layer3_outputs(7353) <= not(layer2_outputs(1610));
    layer3_outputs(7354) <= not(layer2_outputs(5788));
    layer3_outputs(7355) <= layer2_outputs(7317);
    layer3_outputs(7356) <= not(layer2_outputs(4654)) or (layer2_outputs(2678));
    layer3_outputs(7357) <= '0';
    layer3_outputs(7358) <= layer2_outputs(3676);
    layer3_outputs(7359) <= not(layer2_outputs(1580));
    layer3_outputs(7360) <= (layer2_outputs(103)) and not (layer2_outputs(1576));
    layer3_outputs(7361) <= (layer2_outputs(7243)) or (layer2_outputs(3571));
    layer3_outputs(7362) <= not(layer2_outputs(2361));
    layer3_outputs(7363) <= not(layer2_outputs(6546)) or (layer2_outputs(6494));
    layer3_outputs(7364) <= layer2_outputs(3077);
    layer3_outputs(7365) <= layer2_outputs(4405);
    layer3_outputs(7366) <= layer2_outputs(3837);
    layer3_outputs(7367) <= not((layer2_outputs(4577)) and (layer2_outputs(5616)));
    layer3_outputs(7368) <= layer2_outputs(2884);
    layer3_outputs(7369) <= not(layer2_outputs(3604));
    layer3_outputs(7370) <= (layer2_outputs(6131)) or (layer2_outputs(934));
    layer3_outputs(7371) <= (layer2_outputs(6461)) and not (layer2_outputs(3275));
    layer3_outputs(7372) <= (layer2_outputs(1759)) or (layer2_outputs(788));
    layer3_outputs(7373) <= layer2_outputs(4572);
    layer3_outputs(7374) <= layer2_outputs(3436);
    layer3_outputs(7375) <= layer2_outputs(2891);
    layer3_outputs(7376) <= (layer2_outputs(1113)) or (layer2_outputs(7544));
    layer3_outputs(7377) <= layer2_outputs(76);
    layer3_outputs(7378) <= layer2_outputs(2207);
    layer3_outputs(7379) <= not(layer2_outputs(6511));
    layer3_outputs(7380) <= not((layer2_outputs(6530)) xor (layer2_outputs(2108)));
    layer3_outputs(7381) <= layer2_outputs(7486);
    layer3_outputs(7382) <= '0';
    layer3_outputs(7383) <= layer2_outputs(4993);
    layer3_outputs(7384) <= not(layer2_outputs(5607));
    layer3_outputs(7385) <= layer2_outputs(1206);
    layer3_outputs(7386) <= (layer2_outputs(7238)) and not (layer2_outputs(2306));
    layer3_outputs(7387) <= not((layer2_outputs(6110)) xor (layer2_outputs(5765)));
    layer3_outputs(7388) <= not(layer2_outputs(707)) or (layer2_outputs(6435));
    layer3_outputs(7389) <= not(layer2_outputs(5303)) or (layer2_outputs(5120));
    layer3_outputs(7390) <= not(layer2_outputs(1681));
    layer3_outputs(7391) <= not((layer2_outputs(3561)) xor (layer2_outputs(1746)));
    layer3_outputs(7392) <= layer2_outputs(5211);
    layer3_outputs(7393) <= not(layer2_outputs(2655));
    layer3_outputs(7394) <= not(layer2_outputs(4078)) or (layer2_outputs(1016));
    layer3_outputs(7395) <= not(layer2_outputs(7589)) or (layer2_outputs(858));
    layer3_outputs(7396) <= (layer2_outputs(5781)) xor (layer2_outputs(4232));
    layer3_outputs(7397) <= layer2_outputs(6139);
    layer3_outputs(7398) <= not(layer2_outputs(2795));
    layer3_outputs(7399) <= layer2_outputs(6236);
    layer3_outputs(7400) <= not(layer2_outputs(693));
    layer3_outputs(7401) <= layer2_outputs(5648);
    layer3_outputs(7402) <= (layer2_outputs(4695)) and not (layer2_outputs(7473));
    layer3_outputs(7403) <= not((layer2_outputs(404)) and (layer2_outputs(7467)));
    layer3_outputs(7404) <= layer2_outputs(3927);
    layer3_outputs(7405) <= (layer2_outputs(3638)) and not (layer2_outputs(5485));
    layer3_outputs(7406) <= (layer2_outputs(1217)) xor (layer2_outputs(2991));
    layer3_outputs(7407) <= (layer2_outputs(1403)) and (layer2_outputs(5458));
    layer3_outputs(7408) <= not(layer2_outputs(3678));
    layer3_outputs(7409) <= layer2_outputs(5898);
    layer3_outputs(7410) <= (layer2_outputs(2396)) and (layer2_outputs(7470));
    layer3_outputs(7411) <= (layer2_outputs(4087)) and (layer2_outputs(5966));
    layer3_outputs(7412) <= layer2_outputs(4243);
    layer3_outputs(7413) <= not(layer2_outputs(4795));
    layer3_outputs(7414) <= layer2_outputs(4982);
    layer3_outputs(7415) <= '0';
    layer3_outputs(7416) <= not(layer2_outputs(2409));
    layer3_outputs(7417) <= layer2_outputs(2730);
    layer3_outputs(7418) <= layer2_outputs(2175);
    layer3_outputs(7419) <= '0';
    layer3_outputs(7420) <= (layer2_outputs(2391)) and not (layer2_outputs(6231));
    layer3_outputs(7421) <= not((layer2_outputs(1483)) and (layer2_outputs(701)));
    layer3_outputs(7422) <= (layer2_outputs(1063)) and (layer2_outputs(2287));
    layer3_outputs(7423) <= not(layer2_outputs(3949));
    layer3_outputs(7424) <= not(layer2_outputs(410)) or (layer2_outputs(4033));
    layer3_outputs(7425) <= layer2_outputs(2686);
    layer3_outputs(7426) <= not((layer2_outputs(6519)) or (layer2_outputs(7019)));
    layer3_outputs(7427) <= layer2_outputs(2649);
    layer3_outputs(7428) <= layer2_outputs(7118);
    layer3_outputs(7429) <= (layer2_outputs(1040)) or (layer2_outputs(1139));
    layer3_outputs(7430) <= layer2_outputs(1612);
    layer3_outputs(7431) <= layer2_outputs(3204);
    layer3_outputs(7432) <= not(layer2_outputs(106));
    layer3_outputs(7433) <= (layer2_outputs(244)) and (layer2_outputs(4703));
    layer3_outputs(7434) <= (layer2_outputs(4430)) xor (layer2_outputs(3248));
    layer3_outputs(7435) <= not((layer2_outputs(1975)) or (layer2_outputs(2178)));
    layer3_outputs(7436) <= not(layer2_outputs(2582));
    layer3_outputs(7437) <= (layer2_outputs(4133)) and (layer2_outputs(6798));
    layer3_outputs(7438) <= not(layer2_outputs(1358));
    layer3_outputs(7439) <= layer2_outputs(2650);
    layer3_outputs(7440) <= not(layer2_outputs(1976)) or (layer2_outputs(2739));
    layer3_outputs(7441) <= not((layer2_outputs(6689)) or (layer2_outputs(3452)));
    layer3_outputs(7442) <= (layer2_outputs(790)) or (layer2_outputs(7106));
    layer3_outputs(7443) <= not(layer2_outputs(4671)) or (layer2_outputs(3213));
    layer3_outputs(7444) <= not((layer2_outputs(2597)) or (layer2_outputs(238)));
    layer3_outputs(7445) <= (layer2_outputs(987)) or (layer2_outputs(4669));
    layer3_outputs(7446) <= not((layer2_outputs(969)) and (layer2_outputs(5313)));
    layer3_outputs(7447) <= (layer2_outputs(7536)) and (layer2_outputs(98));
    layer3_outputs(7448) <= (layer2_outputs(4721)) and (layer2_outputs(3575));
    layer3_outputs(7449) <= layer2_outputs(7261);
    layer3_outputs(7450) <= not(layer2_outputs(2939));
    layer3_outputs(7451) <= layer2_outputs(1706);
    layer3_outputs(7452) <= layer2_outputs(1350);
    layer3_outputs(7453) <= layer2_outputs(5561);
    layer3_outputs(7454) <= '0';
    layer3_outputs(7455) <= layer2_outputs(7260);
    layer3_outputs(7456) <= not((layer2_outputs(3727)) and (layer2_outputs(6616)));
    layer3_outputs(7457) <= not(layer2_outputs(5078));
    layer3_outputs(7458) <= not((layer2_outputs(6151)) xor (layer2_outputs(3505)));
    layer3_outputs(7459) <= not(layer2_outputs(175));
    layer3_outputs(7460) <= not((layer2_outputs(1014)) and (layer2_outputs(4838)));
    layer3_outputs(7461) <= (layer2_outputs(5460)) xor (layer2_outputs(6016));
    layer3_outputs(7462) <= not(layer2_outputs(3298));
    layer3_outputs(7463) <= not((layer2_outputs(5084)) or (layer2_outputs(894)));
    layer3_outputs(7464) <= not(layer2_outputs(6314)) or (layer2_outputs(3250));
    layer3_outputs(7465) <= not(layer2_outputs(3856));
    layer3_outputs(7466) <= not(layer2_outputs(7566));
    layer3_outputs(7467) <= layer2_outputs(7310);
    layer3_outputs(7468) <= not(layer2_outputs(3516));
    layer3_outputs(7469) <= not((layer2_outputs(6053)) or (layer2_outputs(5218)));
    layer3_outputs(7470) <= (layer2_outputs(5794)) and not (layer2_outputs(6328));
    layer3_outputs(7471) <= layer2_outputs(2087);
    layer3_outputs(7472) <= (layer2_outputs(419)) and (layer2_outputs(3109));
    layer3_outputs(7473) <= '1';
    layer3_outputs(7474) <= not((layer2_outputs(2596)) and (layer2_outputs(4895)));
    layer3_outputs(7475) <= not(layer2_outputs(2842)) or (layer2_outputs(6465));
    layer3_outputs(7476) <= not((layer2_outputs(1933)) and (layer2_outputs(4356)));
    layer3_outputs(7477) <= layer2_outputs(555);
    layer3_outputs(7478) <= not(layer2_outputs(2901));
    layer3_outputs(7479) <= not(layer2_outputs(68)) or (layer2_outputs(3283));
    layer3_outputs(7480) <= (layer2_outputs(3607)) and (layer2_outputs(4207));
    layer3_outputs(7481) <= not(layer2_outputs(763));
    layer3_outputs(7482) <= not((layer2_outputs(5328)) xor (layer2_outputs(6769)));
    layer3_outputs(7483) <= (layer2_outputs(3749)) and not (layer2_outputs(7465));
    layer3_outputs(7484) <= layer2_outputs(3219);
    layer3_outputs(7485) <= not(layer2_outputs(4394));
    layer3_outputs(7486) <= not((layer2_outputs(189)) and (layer2_outputs(3624)));
    layer3_outputs(7487) <= not(layer2_outputs(1347)) or (layer2_outputs(5327));
    layer3_outputs(7488) <= layer2_outputs(529);
    layer3_outputs(7489) <= (layer2_outputs(7042)) and not (layer2_outputs(4656));
    layer3_outputs(7490) <= not((layer2_outputs(1090)) xor (layer2_outputs(1942)));
    layer3_outputs(7491) <= (layer2_outputs(3309)) and not (layer2_outputs(3952));
    layer3_outputs(7492) <= '0';
    layer3_outputs(7493) <= not(layer2_outputs(2438));
    layer3_outputs(7494) <= layer2_outputs(2419);
    layer3_outputs(7495) <= not(layer2_outputs(231));
    layer3_outputs(7496) <= not(layer2_outputs(1627));
    layer3_outputs(7497) <= not(layer2_outputs(3726)) or (layer2_outputs(4051));
    layer3_outputs(7498) <= not(layer2_outputs(4879)) or (layer2_outputs(2854));
    layer3_outputs(7499) <= not((layer2_outputs(4136)) or (layer2_outputs(2405)));
    layer3_outputs(7500) <= not(layer2_outputs(1260));
    layer3_outputs(7501) <= layer2_outputs(7632);
    layer3_outputs(7502) <= layer2_outputs(619);
    layer3_outputs(7503) <= not(layer2_outputs(1302)) or (layer2_outputs(2254));
    layer3_outputs(7504) <= not(layer2_outputs(7207));
    layer3_outputs(7505) <= not((layer2_outputs(900)) and (layer2_outputs(114)));
    layer3_outputs(7506) <= (layer2_outputs(2579)) xor (layer2_outputs(6162));
    layer3_outputs(7507) <= not((layer2_outputs(2812)) xor (layer2_outputs(6983)));
    layer3_outputs(7508) <= layer2_outputs(328);
    layer3_outputs(7509) <= (layer2_outputs(4490)) and not (layer2_outputs(6238));
    layer3_outputs(7510) <= (layer2_outputs(5334)) and (layer2_outputs(3586));
    layer3_outputs(7511) <= (layer2_outputs(6618)) xor (layer2_outputs(5165));
    layer3_outputs(7512) <= not((layer2_outputs(7536)) or (layer2_outputs(6022)));
    layer3_outputs(7513) <= not(layer2_outputs(6043)) or (layer2_outputs(940));
    layer3_outputs(7514) <= not(layer2_outputs(5984));
    layer3_outputs(7515) <= layer2_outputs(3953);
    layer3_outputs(7516) <= not((layer2_outputs(6298)) or (layer2_outputs(5928)));
    layer3_outputs(7517) <= not(layer2_outputs(5746)) or (layer2_outputs(1777));
    layer3_outputs(7518) <= layer2_outputs(5411);
    layer3_outputs(7519) <= layer2_outputs(367);
    layer3_outputs(7520) <= layer2_outputs(4779);
    layer3_outputs(7521) <= not(layer2_outputs(4757)) or (layer2_outputs(2594));
    layer3_outputs(7522) <= layer2_outputs(5066);
    layer3_outputs(7523) <= layer2_outputs(1929);
    layer3_outputs(7524) <= not((layer2_outputs(3886)) or (layer2_outputs(5069)));
    layer3_outputs(7525) <= '1';
    layer3_outputs(7526) <= layer2_outputs(7287);
    layer3_outputs(7527) <= not(layer2_outputs(5909));
    layer3_outputs(7528) <= layer2_outputs(3588);
    layer3_outputs(7529) <= (layer2_outputs(7450)) and not (layer2_outputs(5622));
    layer3_outputs(7530) <= not((layer2_outputs(4375)) xor (layer2_outputs(6799)));
    layer3_outputs(7531) <= (layer2_outputs(7343)) and (layer2_outputs(3048));
    layer3_outputs(7532) <= not(layer2_outputs(2088));
    layer3_outputs(7533) <= not((layer2_outputs(5712)) and (layer2_outputs(7231)));
    layer3_outputs(7534) <= not(layer2_outputs(7298));
    layer3_outputs(7535) <= not(layer2_outputs(1362));
    layer3_outputs(7536) <= (layer2_outputs(4558)) or (layer2_outputs(3639));
    layer3_outputs(7537) <= not(layer2_outputs(3036)) or (layer2_outputs(2257));
    layer3_outputs(7538) <= not(layer2_outputs(4321));
    layer3_outputs(7539) <= (layer2_outputs(719)) and not (layer2_outputs(1144));
    layer3_outputs(7540) <= layer2_outputs(1093);
    layer3_outputs(7541) <= not((layer2_outputs(7638)) or (layer2_outputs(474)));
    layer3_outputs(7542) <= not(layer2_outputs(5050));
    layer3_outputs(7543) <= layer2_outputs(2646);
    layer3_outputs(7544) <= not((layer2_outputs(886)) or (layer2_outputs(3365)));
    layer3_outputs(7545) <= not(layer2_outputs(6367)) or (layer2_outputs(3902));
    layer3_outputs(7546) <= not((layer2_outputs(827)) or (layer2_outputs(193)));
    layer3_outputs(7547) <= (layer2_outputs(7234)) and not (layer2_outputs(3580));
    layer3_outputs(7548) <= (layer2_outputs(1701)) and not (layer2_outputs(3483));
    layer3_outputs(7549) <= not(layer2_outputs(4687)) or (layer2_outputs(7183));
    layer3_outputs(7550) <= not(layer2_outputs(5733)) or (layer2_outputs(2301));
    layer3_outputs(7551) <= not(layer2_outputs(6378));
    layer3_outputs(7552) <= (layer2_outputs(7394)) or (layer2_outputs(3557));
    layer3_outputs(7553) <= '1';
    layer3_outputs(7554) <= (layer2_outputs(6999)) and not (layer2_outputs(3));
    layer3_outputs(7555) <= not(layer2_outputs(6099));
    layer3_outputs(7556) <= layer2_outputs(5002);
    layer3_outputs(7557) <= (layer2_outputs(6584)) xor (layer2_outputs(1526));
    layer3_outputs(7558) <= not(layer2_outputs(6226));
    layer3_outputs(7559) <= not((layer2_outputs(3409)) or (layer2_outputs(5942)));
    layer3_outputs(7560) <= not(layer2_outputs(643)) or (layer2_outputs(5838));
    layer3_outputs(7561) <= layer2_outputs(6596);
    layer3_outputs(7562) <= (layer2_outputs(1235)) xor (layer2_outputs(4074));
    layer3_outputs(7563) <= not(layer2_outputs(5115));
    layer3_outputs(7564) <= (layer2_outputs(4374)) and (layer2_outputs(1286));
    layer3_outputs(7565) <= layer2_outputs(4136);
    layer3_outputs(7566) <= '1';
    layer3_outputs(7567) <= not((layer2_outputs(3881)) and (layer2_outputs(1516)));
    layer3_outputs(7568) <= not(layer2_outputs(6922)) or (layer2_outputs(418));
    layer3_outputs(7569) <= (layer2_outputs(2360)) xor (layer2_outputs(3696));
    layer3_outputs(7570) <= layer2_outputs(4878);
    layer3_outputs(7571) <= not(layer2_outputs(621));
    layer3_outputs(7572) <= '1';
    layer3_outputs(7573) <= not(layer2_outputs(1027)) or (layer2_outputs(5422));
    layer3_outputs(7574) <= not((layer2_outputs(6441)) and (layer2_outputs(2977)));
    layer3_outputs(7575) <= (layer2_outputs(6470)) and not (layer2_outputs(1843));
    layer3_outputs(7576) <= not(layer2_outputs(4461));
    layer3_outputs(7577) <= not(layer2_outputs(5161)) or (layer2_outputs(6977));
    layer3_outputs(7578) <= (layer2_outputs(5272)) and not (layer2_outputs(6339));
    layer3_outputs(7579) <= layer2_outputs(2785);
    layer3_outputs(7580) <= not(layer2_outputs(5485));
    layer3_outputs(7581) <= layer2_outputs(954);
    layer3_outputs(7582) <= not(layer2_outputs(6330)) or (layer2_outputs(1980));
    layer3_outputs(7583) <= layer2_outputs(2317);
    layer3_outputs(7584) <= layer2_outputs(4709);
    layer3_outputs(7585) <= not(layer2_outputs(7115)) or (layer2_outputs(1754));
    layer3_outputs(7586) <= not(layer2_outputs(3564));
    layer3_outputs(7587) <= layer2_outputs(534);
    layer3_outputs(7588) <= not(layer2_outputs(1281));
    layer3_outputs(7589) <= not(layer2_outputs(3475)) or (layer2_outputs(536));
    layer3_outputs(7590) <= layer2_outputs(6047);
    layer3_outputs(7591) <= not(layer2_outputs(4479));
    layer3_outputs(7592) <= layer2_outputs(6380);
    layer3_outputs(7593) <= not((layer2_outputs(600)) and (layer2_outputs(1229)));
    layer3_outputs(7594) <= not((layer2_outputs(902)) or (layer2_outputs(2911)));
    layer3_outputs(7595) <= not(layer2_outputs(1114));
    layer3_outputs(7596) <= layer2_outputs(1607);
    layer3_outputs(7597) <= (layer2_outputs(5617)) and not (layer2_outputs(2281));
    layer3_outputs(7598) <= not(layer2_outputs(1893));
    layer3_outputs(7599) <= not(layer2_outputs(6103));
    layer3_outputs(7600) <= not((layer2_outputs(898)) xor (layer2_outputs(3420)));
    layer3_outputs(7601) <= not(layer2_outputs(859));
    layer3_outputs(7602) <= layer2_outputs(139);
    layer3_outputs(7603) <= not((layer2_outputs(7274)) or (layer2_outputs(2757)));
    layer3_outputs(7604) <= not(layer2_outputs(6200));
    layer3_outputs(7605) <= (layer2_outputs(2806)) xor (layer2_outputs(1239));
    layer3_outputs(7606) <= (layer2_outputs(3579)) and not (layer2_outputs(527));
    layer3_outputs(7607) <= layer2_outputs(2375);
    layer3_outputs(7608) <= not(layer2_outputs(933));
    layer3_outputs(7609) <= layer2_outputs(7180);
    layer3_outputs(7610) <= (layer2_outputs(0)) and not (layer2_outputs(2223));
    layer3_outputs(7611) <= layer2_outputs(6798);
    layer3_outputs(7612) <= not(layer2_outputs(2716)) or (layer2_outputs(5019));
    layer3_outputs(7613) <= layer2_outputs(410);
    layer3_outputs(7614) <= not(layer2_outputs(4533));
    layer3_outputs(7615) <= layer2_outputs(2452);
    layer3_outputs(7616) <= layer2_outputs(1683);
    layer3_outputs(7617) <= layer2_outputs(3619);
    layer3_outputs(7618) <= not(layer2_outputs(4910));
    layer3_outputs(7619) <= (layer2_outputs(6551)) or (layer2_outputs(3664));
    layer3_outputs(7620) <= layer2_outputs(449);
    layer3_outputs(7621) <= not(layer2_outputs(4154)) or (layer2_outputs(901));
    layer3_outputs(7622) <= (layer2_outputs(144)) and (layer2_outputs(1059));
    layer3_outputs(7623) <= layer2_outputs(704);
    layer3_outputs(7624) <= layer2_outputs(5155);
    layer3_outputs(7625) <= layer2_outputs(5780);
    layer3_outputs(7626) <= '1';
    layer3_outputs(7627) <= layer2_outputs(4155);
    layer3_outputs(7628) <= not(layer2_outputs(5590));
    layer3_outputs(7629) <= (layer2_outputs(183)) xor (layer2_outputs(4129));
    layer3_outputs(7630) <= layer2_outputs(1563);
    layer3_outputs(7631) <= layer2_outputs(3597);
    layer3_outputs(7632) <= layer2_outputs(1650);
    layer3_outputs(7633) <= layer2_outputs(1959);
    layer3_outputs(7634) <= layer2_outputs(7151);
    layer3_outputs(7635) <= layer2_outputs(173);
    layer3_outputs(7636) <= layer2_outputs(1105);
    layer3_outputs(7637) <= not((layer2_outputs(793)) and (layer2_outputs(6671)));
    layer3_outputs(7638) <= layer2_outputs(3895);
    layer3_outputs(7639) <= not(layer2_outputs(1829));
    layer3_outputs(7640) <= (layer2_outputs(6731)) xor (layer2_outputs(207));
    layer3_outputs(7641) <= layer2_outputs(544);
    layer3_outputs(7642) <= not((layer2_outputs(4906)) and (layer2_outputs(6393)));
    layer3_outputs(7643) <= not(layer2_outputs(6410));
    layer3_outputs(7644) <= layer2_outputs(5839);
    layer3_outputs(7645) <= not((layer2_outputs(5114)) xor (layer2_outputs(3166)));
    layer3_outputs(7646) <= not(layer2_outputs(6964)) or (layer2_outputs(4502));
    layer3_outputs(7647) <= not(layer2_outputs(990)) or (layer2_outputs(2329));
    layer3_outputs(7648) <= not(layer2_outputs(7492));
    layer3_outputs(7649) <= (layer2_outputs(6241)) xor (layer2_outputs(5319));
    layer3_outputs(7650) <= not(layer2_outputs(5695));
    layer3_outputs(7651) <= layer2_outputs(2186);
    layer3_outputs(7652) <= (layer2_outputs(6040)) or (layer2_outputs(2745));
    layer3_outputs(7653) <= not(layer2_outputs(5945));
    layer3_outputs(7654) <= '0';
    layer3_outputs(7655) <= not(layer2_outputs(549));
    layer3_outputs(7656) <= layer2_outputs(143);
    layer3_outputs(7657) <= layer2_outputs(2561);
    layer3_outputs(7658) <= layer2_outputs(6645);
    layer3_outputs(7659) <= not(layer2_outputs(2489));
    layer3_outputs(7660) <= layer2_outputs(7315);
    layer3_outputs(7661) <= not(layer2_outputs(2998));
    layer3_outputs(7662) <= '1';
    layer3_outputs(7663) <= not(layer2_outputs(4155));
    layer3_outputs(7664) <= layer2_outputs(6579);
    layer3_outputs(7665) <= not(layer2_outputs(3476)) or (layer2_outputs(478));
    layer3_outputs(7666) <= layer2_outputs(2953);
    layer3_outputs(7667) <= (layer2_outputs(113)) xor (layer2_outputs(5779));
    layer3_outputs(7668) <= layer2_outputs(4108);
    layer3_outputs(7669) <= (layer2_outputs(1641)) and not (layer2_outputs(6944));
    layer3_outputs(7670) <= layer2_outputs(5202);
    layer3_outputs(7671) <= not(layer2_outputs(6009)) or (layer2_outputs(5584));
    layer3_outputs(7672) <= (layer2_outputs(4984)) and not (layer2_outputs(4694));
    layer3_outputs(7673) <= not(layer2_outputs(4269));
    layer3_outputs(7674) <= layer2_outputs(3499);
    layer3_outputs(7675) <= not(layer2_outputs(2842));
    layer3_outputs(7676) <= not((layer2_outputs(5973)) xor (layer2_outputs(4893)));
    layer3_outputs(7677) <= layer2_outputs(1350);
    layer3_outputs(7678) <= not(layer2_outputs(7434)) or (layer2_outputs(959));
    layer3_outputs(7679) <= '0';
    layer4_outputs(0) <= not(layer3_outputs(593));
    layer4_outputs(1) <= not(layer3_outputs(1173));
    layer4_outputs(2) <= layer3_outputs(7580);
    layer4_outputs(3) <= not(layer3_outputs(1910)) or (layer3_outputs(3408));
    layer4_outputs(4) <= not(layer3_outputs(4606));
    layer4_outputs(5) <= (layer3_outputs(667)) xor (layer3_outputs(1482));
    layer4_outputs(6) <= not(layer3_outputs(2863));
    layer4_outputs(7) <= not((layer3_outputs(5753)) or (layer3_outputs(7467)));
    layer4_outputs(8) <= '1';
    layer4_outputs(9) <= not(layer3_outputs(6801));
    layer4_outputs(10) <= not(layer3_outputs(1386));
    layer4_outputs(11) <= not(layer3_outputs(6565));
    layer4_outputs(12) <= not(layer3_outputs(2641));
    layer4_outputs(13) <= layer3_outputs(5086);
    layer4_outputs(14) <= not(layer3_outputs(1160));
    layer4_outputs(15) <= not((layer3_outputs(7529)) or (layer3_outputs(4179)));
    layer4_outputs(16) <= layer3_outputs(5009);
    layer4_outputs(17) <= layer3_outputs(6259);
    layer4_outputs(18) <= not(layer3_outputs(3919));
    layer4_outputs(19) <= (layer3_outputs(5607)) and not (layer3_outputs(6305));
    layer4_outputs(20) <= (layer3_outputs(6672)) or (layer3_outputs(5358));
    layer4_outputs(21) <= not((layer3_outputs(3321)) xor (layer3_outputs(5763)));
    layer4_outputs(22) <= layer3_outputs(7042);
    layer4_outputs(23) <= layer3_outputs(1471);
    layer4_outputs(24) <= not(layer3_outputs(1515));
    layer4_outputs(25) <= (layer3_outputs(575)) and not (layer3_outputs(4242));
    layer4_outputs(26) <= not(layer3_outputs(6266));
    layer4_outputs(27) <= not(layer3_outputs(4767));
    layer4_outputs(28) <= (layer3_outputs(3941)) xor (layer3_outputs(2243));
    layer4_outputs(29) <= not(layer3_outputs(3661));
    layer4_outputs(30) <= not(layer3_outputs(92)) or (layer3_outputs(4302));
    layer4_outputs(31) <= layer3_outputs(7597);
    layer4_outputs(32) <= not((layer3_outputs(1710)) xor (layer3_outputs(3705)));
    layer4_outputs(33) <= not(layer3_outputs(6133));
    layer4_outputs(34) <= not((layer3_outputs(1663)) and (layer3_outputs(915)));
    layer4_outputs(35) <= not(layer3_outputs(4167));
    layer4_outputs(36) <= (layer3_outputs(5625)) and not (layer3_outputs(2355));
    layer4_outputs(37) <= layer3_outputs(4921);
    layer4_outputs(38) <= not((layer3_outputs(4706)) or (layer3_outputs(3395)));
    layer4_outputs(39) <= (layer3_outputs(7405)) and (layer3_outputs(6430));
    layer4_outputs(40) <= (layer3_outputs(1792)) and not (layer3_outputs(3392));
    layer4_outputs(41) <= not((layer3_outputs(5933)) and (layer3_outputs(5157)));
    layer4_outputs(42) <= (layer3_outputs(1084)) and (layer3_outputs(1618));
    layer4_outputs(43) <= layer3_outputs(4929);
    layer4_outputs(44) <= layer3_outputs(3474);
    layer4_outputs(45) <= not(layer3_outputs(66));
    layer4_outputs(46) <= layer3_outputs(5639);
    layer4_outputs(47) <= (layer3_outputs(3037)) and not (layer3_outputs(4117));
    layer4_outputs(48) <= (layer3_outputs(1079)) and not (layer3_outputs(3755));
    layer4_outputs(49) <= not(layer3_outputs(4572));
    layer4_outputs(50) <= (layer3_outputs(2433)) and not (layer3_outputs(4781));
    layer4_outputs(51) <= not((layer3_outputs(6651)) xor (layer3_outputs(1657)));
    layer4_outputs(52) <= not((layer3_outputs(1915)) and (layer3_outputs(666)));
    layer4_outputs(53) <= layer3_outputs(2964);
    layer4_outputs(54) <= layer3_outputs(1797);
    layer4_outputs(55) <= not(layer3_outputs(1337)) or (layer3_outputs(6883));
    layer4_outputs(56) <= (layer3_outputs(217)) or (layer3_outputs(2471));
    layer4_outputs(57) <= not(layer3_outputs(2493));
    layer4_outputs(58) <= (layer3_outputs(5572)) and not (layer3_outputs(6633));
    layer4_outputs(59) <= not(layer3_outputs(97)) or (layer3_outputs(5883));
    layer4_outputs(60) <= not(layer3_outputs(3860)) or (layer3_outputs(6918));
    layer4_outputs(61) <= layer3_outputs(672);
    layer4_outputs(62) <= (layer3_outputs(5041)) or (layer3_outputs(7611));
    layer4_outputs(63) <= (layer3_outputs(7333)) and not (layer3_outputs(40));
    layer4_outputs(64) <= not(layer3_outputs(247));
    layer4_outputs(65) <= (layer3_outputs(2724)) xor (layer3_outputs(6500));
    layer4_outputs(66) <= layer3_outputs(1691);
    layer4_outputs(67) <= not(layer3_outputs(3200)) or (layer3_outputs(2122));
    layer4_outputs(68) <= layer3_outputs(1549);
    layer4_outputs(69) <= not(layer3_outputs(989));
    layer4_outputs(70) <= (layer3_outputs(6133)) and not (layer3_outputs(4229));
    layer4_outputs(71) <= not(layer3_outputs(6712));
    layer4_outputs(72) <= not((layer3_outputs(2411)) and (layer3_outputs(2496)));
    layer4_outputs(73) <= not((layer3_outputs(4322)) and (layer3_outputs(3021)));
    layer4_outputs(74) <= (layer3_outputs(6900)) and (layer3_outputs(3180));
    layer4_outputs(75) <= not(layer3_outputs(3258));
    layer4_outputs(76) <= not((layer3_outputs(471)) or (layer3_outputs(392)));
    layer4_outputs(77) <= not(layer3_outputs(6809)) or (layer3_outputs(2990));
    layer4_outputs(78) <= layer3_outputs(2266);
    layer4_outputs(79) <= not(layer3_outputs(2605));
    layer4_outputs(80) <= layer3_outputs(3750);
    layer4_outputs(81) <= not(layer3_outputs(4785));
    layer4_outputs(82) <= not(layer3_outputs(592));
    layer4_outputs(83) <= not(layer3_outputs(5202));
    layer4_outputs(84) <= (layer3_outputs(7509)) xor (layer3_outputs(3714));
    layer4_outputs(85) <= not(layer3_outputs(808));
    layer4_outputs(86) <= (layer3_outputs(6320)) and (layer3_outputs(696));
    layer4_outputs(87) <= not((layer3_outputs(2709)) and (layer3_outputs(1858)));
    layer4_outputs(88) <= not(layer3_outputs(4043));
    layer4_outputs(89) <= not(layer3_outputs(1320));
    layer4_outputs(90) <= (layer3_outputs(6961)) and not (layer3_outputs(3698));
    layer4_outputs(91) <= not(layer3_outputs(2418));
    layer4_outputs(92) <= not(layer3_outputs(6875)) or (layer3_outputs(4997));
    layer4_outputs(93) <= layer3_outputs(7122);
    layer4_outputs(94) <= not((layer3_outputs(4767)) and (layer3_outputs(5088)));
    layer4_outputs(95) <= layer3_outputs(6601);
    layer4_outputs(96) <= layer3_outputs(1709);
    layer4_outputs(97) <= layer3_outputs(2550);
    layer4_outputs(98) <= layer3_outputs(5329);
    layer4_outputs(99) <= not(layer3_outputs(1260));
    layer4_outputs(100) <= layer3_outputs(5269);
    layer4_outputs(101) <= not(layer3_outputs(360)) or (layer3_outputs(5528));
    layer4_outputs(102) <= (layer3_outputs(1416)) or (layer3_outputs(6732));
    layer4_outputs(103) <= layer3_outputs(1356);
    layer4_outputs(104) <= not((layer3_outputs(7414)) or (layer3_outputs(6010)));
    layer4_outputs(105) <= not(layer3_outputs(4819));
    layer4_outputs(106) <= '1';
    layer4_outputs(107) <= not(layer3_outputs(4623)) or (layer3_outputs(6461));
    layer4_outputs(108) <= (layer3_outputs(7644)) and not (layer3_outputs(1053));
    layer4_outputs(109) <= layer3_outputs(4337);
    layer4_outputs(110) <= not(layer3_outputs(6793));
    layer4_outputs(111) <= layer3_outputs(7048);
    layer4_outputs(112) <= not(layer3_outputs(4283));
    layer4_outputs(113) <= layer3_outputs(7139);
    layer4_outputs(114) <= not((layer3_outputs(880)) or (layer3_outputs(4091)));
    layer4_outputs(115) <= not((layer3_outputs(6846)) xor (layer3_outputs(1502)));
    layer4_outputs(116) <= layer3_outputs(2101);
    layer4_outputs(117) <= layer3_outputs(7372);
    layer4_outputs(118) <= layer3_outputs(6550);
    layer4_outputs(119) <= not(layer3_outputs(2431));
    layer4_outputs(120) <= not((layer3_outputs(6284)) xor (layer3_outputs(6151)));
    layer4_outputs(121) <= (layer3_outputs(6313)) or (layer3_outputs(145));
    layer4_outputs(122) <= (layer3_outputs(7083)) or (layer3_outputs(7378));
    layer4_outputs(123) <= '0';
    layer4_outputs(124) <= (layer3_outputs(665)) and not (layer3_outputs(4258));
    layer4_outputs(125) <= not(layer3_outputs(2970));
    layer4_outputs(126) <= not(layer3_outputs(7349));
    layer4_outputs(127) <= layer3_outputs(4247);
    layer4_outputs(128) <= (layer3_outputs(5306)) and not (layer3_outputs(4582));
    layer4_outputs(129) <= layer3_outputs(2627);
    layer4_outputs(130) <= (layer3_outputs(4111)) and (layer3_outputs(1353));
    layer4_outputs(131) <= (layer3_outputs(3450)) and (layer3_outputs(1790));
    layer4_outputs(132) <= not(layer3_outputs(3060));
    layer4_outputs(133) <= layer3_outputs(5786);
    layer4_outputs(134) <= layer3_outputs(5910);
    layer4_outputs(135) <= not((layer3_outputs(7634)) or (layer3_outputs(4702)));
    layer4_outputs(136) <= (layer3_outputs(2021)) xor (layer3_outputs(1167));
    layer4_outputs(137) <= layer3_outputs(6685);
    layer4_outputs(138) <= '1';
    layer4_outputs(139) <= layer3_outputs(2343);
    layer4_outputs(140) <= (layer3_outputs(6191)) and (layer3_outputs(1270));
    layer4_outputs(141) <= not(layer3_outputs(7493));
    layer4_outputs(142) <= (layer3_outputs(3227)) and not (layer3_outputs(3377));
    layer4_outputs(143) <= not((layer3_outputs(3960)) xor (layer3_outputs(6448)));
    layer4_outputs(144) <= not(layer3_outputs(478)) or (layer3_outputs(1422));
    layer4_outputs(145) <= layer3_outputs(871);
    layer4_outputs(146) <= not(layer3_outputs(112));
    layer4_outputs(147) <= not((layer3_outputs(6469)) xor (layer3_outputs(6214)));
    layer4_outputs(148) <= (layer3_outputs(5582)) xor (layer3_outputs(2707));
    layer4_outputs(149) <= layer3_outputs(5542);
    layer4_outputs(150) <= (layer3_outputs(678)) and not (layer3_outputs(4143));
    layer4_outputs(151) <= not(layer3_outputs(6815));
    layer4_outputs(152) <= (layer3_outputs(1756)) xor (layer3_outputs(581));
    layer4_outputs(153) <= layer3_outputs(903);
    layer4_outputs(154) <= (layer3_outputs(7617)) xor (layer3_outputs(5595));
    layer4_outputs(155) <= not(layer3_outputs(4651));
    layer4_outputs(156) <= layer3_outputs(4847);
    layer4_outputs(157) <= not((layer3_outputs(2644)) xor (layer3_outputs(6416)));
    layer4_outputs(158) <= not((layer3_outputs(6694)) xor (layer3_outputs(6280)));
    layer4_outputs(159) <= not(layer3_outputs(4608));
    layer4_outputs(160) <= not(layer3_outputs(5416));
    layer4_outputs(161) <= '0';
    layer4_outputs(162) <= (layer3_outputs(4564)) or (layer3_outputs(879));
    layer4_outputs(163) <= (layer3_outputs(6985)) or (layer3_outputs(252));
    layer4_outputs(164) <= not(layer3_outputs(4049));
    layer4_outputs(165) <= not((layer3_outputs(3561)) or (layer3_outputs(7557)));
    layer4_outputs(166) <= (layer3_outputs(462)) or (layer3_outputs(6200));
    layer4_outputs(167) <= (layer3_outputs(5095)) or (layer3_outputs(5365));
    layer4_outputs(168) <= not((layer3_outputs(6907)) and (layer3_outputs(5164)));
    layer4_outputs(169) <= not(layer3_outputs(1368)) or (layer3_outputs(5812));
    layer4_outputs(170) <= (layer3_outputs(3113)) and (layer3_outputs(122));
    layer4_outputs(171) <= (layer3_outputs(154)) and not (layer3_outputs(4294));
    layer4_outputs(172) <= not((layer3_outputs(1352)) and (layer3_outputs(10)));
    layer4_outputs(173) <= layer3_outputs(2005);
    layer4_outputs(174) <= layer3_outputs(4733);
    layer4_outputs(175) <= not(layer3_outputs(22)) or (layer3_outputs(1534));
    layer4_outputs(176) <= (layer3_outputs(5986)) and (layer3_outputs(1480));
    layer4_outputs(177) <= not((layer3_outputs(510)) or (layer3_outputs(4222)));
    layer4_outputs(178) <= layer3_outputs(4992);
    layer4_outputs(179) <= not(layer3_outputs(7250));
    layer4_outputs(180) <= (layer3_outputs(5978)) xor (layer3_outputs(2068));
    layer4_outputs(181) <= '0';
    layer4_outputs(182) <= not(layer3_outputs(6138));
    layer4_outputs(183) <= not(layer3_outputs(6003));
    layer4_outputs(184) <= layer3_outputs(4845);
    layer4_outputs(185) <= layer3_outputs(5239);
    layer4_outputs(186) <= layer3_outputs(3368);
    layer4_outputs(187) <= (layer3_outputs(4836)) and not (layer3_outputs(6247));
    layer4_outputs(188) <= layer3_outputs(6981);
    layer4_outputs(189) <= layer3_outputs(3094);
    layer4_outputs(190) <= layer3_outputs(4041);
    layer4_outputs(191) <= layer3_outputs(1438);
    layer4_outputs(192) <= layer3_outputs(4948);
    layer4_outputs(193) <= (layer3_outputs(1861)) and not (layer3_outputs(3237));
    layer4_outputs(194) <= not(layer3_outputs(6046)) or (layer3_outputs(6976));
    layer4_outputs(195) <= not(layer3_outputs(4884));
    layer4_outputs(196) <= not(layer3_outputs(6017)) or (layer3_outputs(537));
    layer4_outputs(197) <= not(layer3_outputs(5907));
    layer4_outputs(198) <= not((layer3_outputs(391)) xor (layer3_outputs(481)));
    layer4_outputs(199) <= not(layer3_outputs(5414));
    layer4_outputs(200) <= layer3_outputs(133);
    layer4_outputs(201) <= (layer3_outputs(4398)) and not (layer3_outputs(5141));
    layer4_outputs(202) <= not(layer3_outputs(5683)) or (layer3_outputs(162));
    layer4_outputs(203) <= not((layer3_outputs(5770)) or (layer3_outputs(5903)));
    layer4_outputs(204) <= (layer3_outputs(5834)) xor (layer3_outputs(3492));
    layer4_outputs(205) <= not(layer3_outputs(1838)) or (layer3_outputs(5714));
    layer4_outputs(206) <= not(layer3_outputs(7114));
    layer4_outputs(207) <= not(layer3_outputs(1426));
    layer4_outputs(208) <= not((layer3_outputs(7030)) or (layer3_outputs(7461)));
    layer4_outputs(209) <= not((layer3_outputs(6424)) or (layer3_outputs(2558)));
    layer4_outputs(210) <= not(layer3_outputs(3856));
    layer4_outputs(211) <= (layer3_outputs(1679)) and (layer3_outputs(5001));
    layer4_outputs(212) <= layer3_outputs(1189);
    layer4_outputs(213) <= not(layer3_outputs(4151)) or (layer3_outputs(4679));
    layer4_outputs(214) <= not(layer3_outputs(146));
    layer4_outputs(215) <= (layer3_outputs(2506)) or (layer3_outputs(7589));
    layer4_outputs(216) <= layer3_outputs(3196);
    layer4_outputs(217) <= not(layer3_outputs(958));
    layer4_outputs(218) <= not((layer3_outputs(6422)) xor (layer3_outputs(6756)));
    layer4_outputs(219) <= not(layer3_outputs(6630));
    layer4_outputs(220) <= (layer3_outputs(5871)) xor (layer3_outputs(6154));
    layer4_outputs(221) <= not(layer3_outputs(6782)) or (layer3_outputs(3263));
    layer4_outputs(222) <= layer3_outputs(1770);
    layer4_outputs(223) <= not((layer3_outputs(4152)) and (layer3_outputs(2766)));
    layer4_outputs(224) <= not((layer3_outputs(2888)) or (layer3_outputs(1298)));
    layer4_outputs(225) <= (layer3_outputs(1812)) or (layer3_outputs(3584));
    layer4_outputs(226) <= not((layer3_outputs(3199)) or (layer3_outputs(3604)));
    layer4_outputs(227) <= not(layer3_outputs(7508));
    layer4_outputs(228) <= not((layer3_outputs(6082)) xor (layer3_outputs(5723)));
    layer4_outputs(229) <= layer3_outputs(7060);
    layer4_outputs(230) <= not(layer3_outputs(3557));
    layer4_outputs(231) <= not(layer3_outputs(4165));
    layer4_outputs(232) <= not(layer3_outputs(515));
    layer4_outputs(233) <= not(layer3_outputs(874));
    layer4_outputs(234) <= not(layer3_outputs(596)) or (layer3_outputs(4171));
    layer4_outputs(235) <= not((layer3_outputs(4722)) or (layer3_outputs(6729)));
    layer4_outputs(236) <= not((layer3_outputs(7178)) or (layer3_outputs(7310)));
    layer4_outputs(237) <= (layer3_outputs(432)) and not (layer3_outputs(2397));
    layer4_outputs(238) <= not(layer3_outputs(6888));
    layer4_outputs(239) <= (layer3_outputs(2193)) and (layer3_outputs(2318));
    layer4_outputs(240) <= not(layer3_outputs(283)) or (layer3_outputs(5760));
    layer4_outputs(241) <= (layer3_outputs(3916)) xor (layer3_outputs(7402));
    layer4_outputs(242) <= (layer3_outputs(3827)) xor (layer3_outputs(5545));
    layer4_outputs(243) <= not(layer3_outputs(6241));
    layer4_outputs(244) <= not((layer3_outputs(102)) or (layer3_outputs(1749)));
    layer4_outputs(245) <= layer3_outputs(1845);
    layer4_outputs(246) <= (layer3_outputs(1078)) xor (layer3_outputs(2044));
    layer4_outputs(247) <= not(layer3_outputs(1889));
    layer4_outputs(248) <= not(layer3_outputs(1279)) or (layer3_outputs(6735));
    layer4_outputs(249) <= not(layer3_outputs(5873)) or (layer3_outputs(1582));
    layer4_outputs(250) <= not(layer3_outputs(5557));
    layer4_outputs(251) <= not((layer3_outputs(3623)) xor (layer3_outputs(2993)));
    layer4_outputs(252) <= not(layer3_outputs(3077)) or (layer3_outputs(231));
    layer4_outputs(253) <= not((layer3_outputs(1423)) xor (layer3_outputs(5998)));
    layer4_outputs(254) <= not(layer3_outputs(7616));
    layer4_outputs(255) <= (layer3_outputs(5656)) xor (layer3_outputs(2077));
    layer4_outputs(256) <= not((layer3_outputs(569)) and (layer3_outputs(5668)));
    layer4_outputs(257) <= layer3_outputs(4758);
    layer4_outputs(258) <= not((layer3_outputs(3649)) xor (layer3_outputs(6668)));
    layer4_outputs(259) <= not(layer3_outputs(1222));
    layer4_outputs(260) <= layer3_outputs(6061);
    layer4_outputs(261) <= not(layer3_outputs(144));
    layer4_outputs(262) <= (layer3_outputs(19)) and not (layer3_outputs(5138));
    layer4_outputs(263) <= not((layer3_outputs(6307)) or (layer3_outputs(5218)));
    layer4_outputs(264) <= not(layer3_outputs(1745));
    layer4_outputs(265) <= not(layer3_outputs(471));
    layer4_outputs(266) <= layer3_outputs(689);
    layer4_outputs(267) <= not(layer3_outputs(5460));
    layer4_outputs(268) <= layer3_outputs(7468);
    layer4_outputs(269) <= not((layer3_outputs(3359)) and (layer3_outputs(3193)));
    layer4_outputs(270) <= (layer3_outputs(3795)) xor (layer3_outputs(2715));
    layer4_outputs(271) <= not(layer3_outputs(71));
    layer4_outputs(272) <= layer3_outputs(5524);
    layer4_outputs(273) <= not((layer3_outputs(3949)) or (layer3_outputs(72)));
    layer4_outputs(274) <= not((layer3_outputs(1773)) or (layer3_outputs(6926)));
    layer4_outputs(275) <= not((layer3_outputs(2362)) and (layer3_outputs(4365)));
    layer4_outputs(276) <= not((layer3_outputs(489)) xor (layer3_outputs(2611)));
    layer4_outputs(277) <= layer3_outputs(175);
    layer4_outputs(278) <= not(layer3_outputs(6720)) or (layer3_outputs(2013));
    layer4_outputs(279) <= (layer3_outputs(4068)) xor (layer3_outputs(4543));
    layer4_outputs(280) <= (layer3_outputs(4175)) or (layer3_outputs(5673));
    layer4_outputs(281) <= not(layer3_outputs(5783)) or (layer3_outputs(5493));
    layer4_outputs(282) <= not(layer3_outputs(1490));
    layer4_outputs(283) <= not(layer3_outputs(186));
    layer4_outputs(284) <= not((layer3_outputs(5068)) xor (layer3_outputs(1499)));
    layer4_outputs(285) <= not(layer3_outputs(5401));
    layer4_outputs(286) <= not(layer3_outputs(6920));
    layer4_outputs(287) <= (layer3_outputs(4376)) and (layer3_outputs(1447));
    layer4_outputs(288) <= (layer3_outputs(6255)) and not (layer3_outputs(1906));
    layer4_outputs(289) <= not(layer3_outputs(3042));
    layer4_outputs(290) <= not(layer3_outputs(1648)) or (layer3_outputs(4987));
    layer4_outputs(291) <= not(layer3_outputs(6121));
    layer4_outputs(292) <= not((layer3_outputs(7310)) and (layer3_outputs(6663)));
    layer4_outputs(293) <= not(layer3_outputs(1334));
    layer4_outputs(294) <= (layer3_outputs(6953)) and not (layer3_outputs(4070));
    layer4_outputs(295) <= layer3_outputs(2905);
    layer4_outputs(296) <= not((layer3_outputs(49)) and (layer3_outputs(1647)));
    layer4_outputs(297) <= (layer3_outputs(2292)) xor (layer3_outputs(4107));
    layer4_outputs(298) <= not(layer3_outputs(6257));
    layer4_outputs(299) <= (layer3_outputs(3397)) or (layer3_outputs(2806));
    layer4_outputs(300) <= (layer3_outputs(5087)) xor (layer3_outputs(5328));
    layer4_outputs(301) <= not(layer3_outputs(4573)) or (layer3_outputs(1483));
    layer4_outputs(302) <= not((layer3_outputs(2436)) or (layer3_outputs(1539)));
    layer4_outputs(303) <= (layer3_outputs(7119)) and not (layer3_outputs(3929));
    layer4_outputs(304) <= not(layer3_outputs(3230));
    layer4_outputs(305) <= not(layer3_outputs(3823));
    layer4_outputs(306) <= (layer3_outputs(5250)) and not (layer3_outputs(4292));
    layer4_outputs(307) <= layer3_outputs(2513);
    layer4_outputs(308) <= layer3_outputs(489);
    layer4_outputs(309) <= not((layer3_outputs(5602)) xor (layer3_outputs(1873)));
    layer4_outputs(310) <= layer3_outputs(3222);
    layer4_outputs(311) <= (layer3_outputs(2019)) and not (layer3_outputs(2776));
    layer4_outputs(312) <= '0';
    layer4_outputs(313) <= (layer3_outputs(3440)) and (layer3_outputs(4351));
    layer4_outputs(314) <= not(layer3_outputs(2387));
    layer4_outputs(315) <= (layer3_outputs(5506)) or (layer3_outputs(5647));
    layer4_outputs(316) <= layer3_outputs(1849);
    layer4_outputs(317) <= layer3_outputs(706);
    layer4_outputs(318) <= not(layer3_outputs(3159));
    layer4_outputs(319) <= not(layer3_outputs(7588));
    layer4_outputs(320) <= not((layer3_outputs(1785)) and (layer3_outputs(5986)));
    layer4_outputs(321) <= not(layer3_outputs(1695)) or (layer3_outputs(4363));
    layer4_outputs(322) <= (layer3_outputs(1788)) and not (layer3_outputs(6269));
    layer4_outputs(323) <= not(layer3_outputs(3274));
    layer4_outputs(324) <= not((layer3_outputs(5070)) or (layer3_outputs(4793)));
    layer4_outputs(325) <= (layer3_outputs(1775)) or (layer3_outputs(845));
    layer4_outputs(326) <= not(layer3_outputs(6864));
    layer4_outputs(327) <= not(layer3_outputs(3058));
    layer4_outputs(328) <= (layer3_outputs(7642)) xor (layer3_outputs(1271));
    layer4_outputs(329) <= (layer3_outputs(7323)) and not (layer3_outputs(928));
    layer4_outputs(330) <= not(layer3_outputs(2997));
    layer4_outputs(331) <= (layer3_outputs(3904)) xor (layer3_outputs(1294));
    layer4_outputs(332) <= (layer3_outputs(7325)) xor (layer3_outputs(6893));
    layer4_outputs(333) <= layer3_outputs(7149);
    layer4_outputs(334) <= not(layer3_outputs(6314));
    layer4_outputs(335) <= layer3_outputs(6423);
    layer4_outputs(336) <= layer3_outputs(4367);
    layer4_outputs(337) <= not((layer3_outputs(3585)) and (layer3_outputs(3741)));
    layer4_outputs(338) <= layer3_outputs(6076);
    layer4_outputs(339) <= not(layer3_outputs(630));
    layer4_outputs(340) <= not(layer3_outputs(2584));
    layer4_outputs(341) <= not(layer3_outputs(6054)) or (layer3_outputs(4445));
    layer4_outputs(342) <= layer3_outputs(2055);
    layer4_outputs(343) <= (layer3_outputs(5964)) and not (layer3_outputs(431));
    layer4_outputs(344) <= layer3_outputs(7114);
    layer4_outputs(345) <= not(layer3_outputs(21));
    layer4_outputs(346) <= not((layer3_outputs(280)) xor (layer3_outputs(1627)));
    layer4_outputs(347) <= not(layer3_outputs(6738)) or (layer3_outputs(6710));
    layer4_outputs(348) <= not(layer3_outputs(5339));
    layer4_outputs(349) <= layer3_outputs(2377);
    layer4_outputs(350) <= not(layer3_outputs(2237));
    layer4_outputs(351) <= layer3_outputs(5117);
    layer4_outputs(352) <= not((layer3_outputs(5502)) xor (layer3_outputs(3220)));
    layer4_outputs(353) <= not(layer3_outputs(1269));
    layer4_outputs(354) <= layer3_outputs(6332);
    layer4_outputs(355) <= layer3_outputs(4586);
    layer4_outputs(356) <= not(layer3_outputs(456));
    layer4_outputs(357) <= layer3_outputs(631);
    layer4_outputs(358) <= layer3_outputs(1890);
    layer4_outputs(359) <= not(layer3_outputs(7265));
    layer4_outputs(360) <= layer3_outputs(6808);
    layer4_outputs(361) <= layer3_outputs(5728);
    layer4_outputs(362) <= not(layer3_outputs(5780));
    layer4_outputs(363) <= layer3_outputs(2634);
    layer4_outputs(364) <= not(layer3_outputs(6770));
    layer4_outputs(365) <= not(layer3_outputs(1303));
    layer4_outputs(366) <= not(layer3_outputs(7361));
    layer4_outputs(367) <= not(layer3_outputs(2696));
    layer4_outputs(368) <= layer3_outputs(3871);
    layer4_outputs(369) <= '1';
    layer4_outputs(370) <= not((layer3_outputs(4425)) and (layer3_outputs(218)));
    layer4_outputs(371) <= (layer3_outputs(2450)) and (layer3_outputs(3276));
    layer4_outputs(372) <= not((layer3_outputs(982)) or (layer3_outputs(1042)));
    layer4_outputs(373) <= layer3_outputs(1632);
    layer4_outputs(374) <= not((layer3_outputs(2439)) or (layer3_outputs(2377)));
    layer4_outputs(375) <= (layer3_outputs(3176)) and (layer3_outputs(4822));
    layer4_outputs(376) <= layer3_outputs(214);
    layer4_outputs(377) <= (layer3_outputs(2104)) xor (layer3_outputs(3334));
    layer4_outputs(378) <= (layer3_outputs(1702)) and not (layer3_outputs(7364));
    layer4_outputs(379) <= not(layer3_outputs(1954));
    layer4_outputs(380) <= not(layer3_outputs(5099));
    layer4_outputs(381) <= (layer3_outputs(7164)) and not (layer3_outputs(2916));
    layer4_outputs(382) <= (layer3_outputs(2614)) or (layer3_outputs(1286));
    layer4_outputs(383) <= (layer3_outputs(6574)) and not (layer3_outputs(5691));
    layer4_outputs(384) <= not(layer3_outputs(4902));
    layer4_outputs(385) <= (layer3_outputs(3883)) xor (layer3_outputs(1831));
    layer4_outputs(386) <= layer3_outputs(7425);
    layer4_outputs(387) <= layer3_outputs(2829);
    layer4_outputs(388) <= layer3_outputs(1794);
    layer4_outputs(389) <= not(layer3_outputs(6175));
    layer4_outputs(390) <= layer3_outputs(2645);
    layer4_outputs(391) <= not(layer3_outputs(5988));
    layer4_outputs(392) <= not(layer3_outputs(7316));
    layer4_outputs(393) <= (layer3_outputs(5386)) and (layer3_outputs(179));
    layer4_outputs(394) <= not(layer3_outputs(6518));
    layer4_outputs(395) <= layer3_outputs(5540);
    layer4_outputs(396) <= not(layer3_outputs(366));
    layer4_outputs(397) <= (layer3_outputs(4012)) and not (layer3_outputs(3848));
    layer4_outputs(398) <= (layer3_outputs(5348)) and not (layer3_outputs(2811));
    layer4_outputs(399) <= layer3_outputs(1426);
    layer4_outputs(400) <= not(layer3_outputs(4944));
    layer4_outputs(401) <= (layer3_outputs(6252)) and (layer3_outputs(4851));
    layer4_outputs(402) <= '1';
    layer4_outputs(403) <= not(layer3_outputs(2176)) or (layer3_outputs(1022));
    layer4_outputs(404) <= layer3_outputs(1399);
    layer4_outputs(405) <= layer3_outputs(470);
    layer4_outputs(406) <= not((layer3_outputs(7340)) xor (layer3_outputs(2123)));
    layer4_outputs(407) <= not(layer3_outputs(7254));
    layer4_outputs(408) <= not((layer3_outputs(5517)) xor (layer3_outputs(5604)));
    layer4_outputs(409) <= not(layer3_outputs(4001)) or (layer3_outputs(2278));
    layer4_outputs(410) <= not(layer3_outputs(2140)) or (layer3_outputs(4203));
    layer4_outputs(411) <= not((layer3_outputs(579)) xor (layer3_outputs(4667)));
    layer4_outputs(412) <= not((layer3_outputs(6228)) and (layer3_outputs(2362)));
    layer4_outputs(413) <= layer3_outputs(6852);
    layer4_outputs(414) <= layer3_outputs(967);
    layer4_outputs(415) <= (layer3_outputs(5834)) and (layer3_outputs(350));
    layer4_outputs(416) <= (layer3_outputs(4080)) xor (layer3_outputs(2924));
    layer4_outputs(417) <= (layer3_outputs(5355)) and not (layer3_outputs(5127));
    layer4_outputs(418) <= not(layer3_outputs(1441));
    layer4_outputs(419) <= not((layer3_outputs(3973)) and (layer3_outputs(2852)));
    layer4_outputs(420) <= not(layer3_outputs(4184)) or (layer3_outputs(1190));
    layer4_outputs(421) <= (layer3_outputs(1717)) xor (layer3_outputs(1049));
    layer4_outputs(422) <= layer3_outputs(3116);
    layer4_outputs(423) <= (layer3_outputs(6597)) and not (layer3_outputs(3720));
    layer4_outputs(424) <= (layer3_outputs(3486)) xor (layer3_outputs(4498));
    layer4_outputs(425) <= not(layer3_outputs(7475));
    layer4_outputs(426) <= layer3_outputs(2725);
    layer4_outputs(427) <= layer3_outputs(7413);
    layer4_outputs(428) <= layer3_outputs(2883);
    layer4_outputs(429) <= not(layer3_outputs(6021));
    layer4_outputs(430) <= layer3_outputs(3511);
    layer4_outputs(431) <= not(layer3_outputs(6719)) or (layer3_outputs(3005));
    layer4_outputs(432) <= not(layer3_outputs(227));
    layer4_outputs(433) <= not(layer3_outputs(6153));
    layer4_outputs(434) <= (layer3_outputs(4325)) and not (layer3_outputs(4452));
    layer4_outputs(435) <= layer3_outputs(5876);
    layer4_outputs(436) <= not(layer3_outputs(750)) or (layer3_outputs(7069));
    layer4_outputs(437) <= not(layer3_outputs(6316));
    layer4_outputs(438) <= (layer3_outputs(6619)) or (layer3_outputs(5215));
    layer4_outputs(439) <= not(layer3_outputs(6237));
    layer4_outputs(440) <= not(layer3_outputs(2597));
    layer4_outputs(441) <= (layer3_outputs(7246)) and not (layer3_outputs(5138));
    layer4_outputs(442) <= layer3_outputs(3278);
    layer4_outputs(443) <= not((layer3_outputs(6779)) and (layer3_outputs(4314)));
    layer4_outputs(444) <= not(layer3_outputs(4149)) or (layer3_outputs(7506));
    layer4_outputs(445) <= not(layer3_outputs(7034));
    layer4_outputs(446) <= not(layer3_outputs(3092));
    layer4_outputs(447) <= not(layer3_outputs(3694));
    layer4_outputs(448) <= not(layer3_outputs(5181));
    layer4_outputs(449) <= layer3_outputs(4560);
    layer4_outputs(450) <= (layer3_outputs(1460)) or (layer3_outputs(6088));
    layer4_outputs(451) <= not((layer3_outputs(2661)) xor (layer3_outputs(2826)));
    layer4_outputs(452) <= not(layer3_outputs(6343));
    layer4_outputs(453) <= (layer3_outputs(6315)) and not (layer3_outputs(1585));
    layer4_outputs(454) <= not((layer3_outputs(7170)) or (layer3_outputs(1923)));
    layer4_outputs(455) <= not((layer3_outputs(5639)) xor (layer3_outputs(725)));
    layer4_outputs(456) <= (layer3_outputs(3639)) xor (layer3_outputs(4331));
    layer4_outputs(457) <= (layer3_outputs(3031)) and (layer3_outputs(3866));
    layer4_outputs(458) <= not(layer3_outputs(7556));
    layer4_outputs(459) <= layer3_outputs(3374);
    layer4_outputs(460) <= (layer3_outputs(3792)) or (layer3_outputs(5605));
    layer4_outputs(461) <= not((layer3_outputs(5094)) or (layer3_outputs(104)));
    layer4_outputs(462) <= layer3_outputs(6831);
    layer4_outputs(463) <= layer3_outputs(7280);
    layer4_outputs(464) <= layer3_outputs(1563);
    layer4_outputs(465) <= not(layer3_outputs(719));
    layer4_outputs(466) <= (layer3_outputs(1200)) and not (layer3_outputs(6237));
    layer4_outputs(467) <= not(layer3_outputs(2150));
    layer4_outputs(468) <= layer3_outputs(529);
    layer4_outputs(469) <= layer3_outputs(3840);
    layer4_outputs(470) <= layer3_outputs(1310);
    layer4_outputs(471) <= not(layer3_outputs(7363));
    layer4_outputs(472) <= not((layer3_outputs(3583)) or (layer3_outputs(7217)));
    layer4_outputs(473) <= layer3_outputs(2109);
    layer4_outputs(474) <= layer3_outputs(742);
    layer4_outputs(475) <= (layer3_outputs(2022)) and (layer3_outputs(5746));
    layer4_outputs(476) <= not(layer3_outputs(3980));
    layer4_outputs(477) <= layer3_outputs(6231);
    layer4_outputs(478) <= not((layer3_outputs(796)) and (layer3_outputs(5139)));
    layer4_outputs(479) <= not((layer3_outputs(5442)) or (layer3_outputs(2592)));
    layer4_outputs(480) <= not((layer3_outputs(3072)) and (layer3_outputs(6453)));
    layer4_outputs(481) <= not((layer3_outputs(1082)) and (layer3_outputs(6344)));
    layer4_outputs(482) <= not((layer3_outputs(350)) and (layer3_outputs(1715)));
    layer4_outputs(483) <= not(layer3_outputs(638));
    layer4_outputs(484) <= not(layer3_outputs(2794)) or (layer3_outputs(6570));
    layer4_outputs(485) <= (layer3_outputs(6065)) and not (layer3_outputs(6106));
    layer4_outputs(486) <= not(layer3_outputs(6246));
    layer4_outputs(487) <= (layer3_outputs(1829)) or (layer3_outputs(6163));
    layer4_outputs(488) <= (layer3_outputs(1320)) xor (layer3_outputs(4339));
    layer4_outputs(489) <= layer3_outputs(5169);
    layer4_outputs(490) <= (layer3_outputs(2483)) and not (layer3_outputs(4787));
    layer4_outputs(491) <= not((layer3_outputs(6740)) xor (layer3_outputs(3544)));
    layer4_outputs(492) <= not(layer3_outputs(6023));
    layer4_outputs(493) <= (layer3_outputs(5599)) xor (layer3_outputs(3294));
    layer4_outputs(494) <= not(layer3_outputs(3401));
    layer4_outputs(495) <= not(layer3_outputs(92)) or (layer3_outputs(5350));
    layer4_outputs(496) <= layer3_outputs(3871);
    layer4_outputs(497) <= layer3_outputs(750);
    layer4_outputs(498) <= not(layer3_outputs(5047));
    layer4_outputs(499) <= layer3_outputs(7601);
    layer4_outputs(500) <= not(layer3_outputs(2548));
    layer4_outputs(501) <= not((layer3_outputs(2577)) or (layer3_outputs(4283)));
    layer4_outputs(502) <= (layer3_outputs(3685)) xor (layer3_outputs(708));
    layer4_outputs(503) <= not(layer3_outputs(7383)) or (layer3_outputs(3170));
    layer4_outputs(504) <= not(layer3_outputs(818)) or (layer3_outputs(3313));
    layer4_outputs(505) <= not((layer3_outputs(1536)) and (layer3_outputs(3059)));
    layer4_outputs(506) <= layer3_outputs(604);
    layer4_outputs(507) <= not(layer3_outputs(5520));
    layer4_outputs(508) <= not((layer3_outputs(5771)) xor (layer3_outputs(4920)));
    layer4_outputs(509) <= (layer3_outputs(5727)) and (layer3_outputs(6762));
    layer4_outputs(510) <= not(layer3_outputs(2337));
    layer4_outputs(511) <= layer3_outputs(3248);
    layer4_outputs(512) <= not((layer3_outputs(398)) or (layer3_outputs(4507)));
    layer4_outputs(513) <= not(layer3_outputs(5443));
    layer4_outputs(514) <= (layer3_outputs(4954)) or (layer3_outputs(816));
    layer4_outputs(515) <= layer3_outputs(6679);
    layer4_outputs(516) <= (layer3_outputs(1330)) and not (layer3_outputs(5325));
    layer4_outputs(517) <= not(layer3_outputs(4401));
    layer4_outputs(518) <= layer3_outputs(1019);
    layer4_outputs(519) <= layer3_outputs(1152);
    layer4_outputs(520) <= layer3_outputs(4402);
    layer4_outputs(521) <= (layer3_outputs(7672)) or (layer3_outputs(7028));
    layer4_outputs(522) <= not((layer3_outputs(1843)) xor (layer3_outputs(6658)));
    layer4_outputs(523) <= not((layer3_outputs(3197)) xor (layer3_outputs(1827)));
    layer4_outputs(524) <= not((layer3_outputs(3487)) or (layer3_outputs(3088)));
    layer4_outputs(525) <= not(layer3_outputs(6434));
    layer4_outputs(526) <= not(layer3_outputs(3178)) or (layer3_outputs(3778));
    layer4_outputs(527) <= not(layer3_outputs(1554));
    layer4_outputs(528) <= not((layer3_outputs(1058)) xor (layer3_outputs(7492)));
    layer4_outputs(529) <= layer3_outputs(3582);
    layer4_outputs(530) <= (layer3_outputs(5896)) and (layer3_outputs(7287));
    layer4_outputs(531) <= not(layer3_outputs(747));
    layer4_outputs(532) <= (layer3_outputs(4995)) or (layer3_outputs(5982));
    layer4_outputs(533) <= not((layer3_outputs(7360)) and (layer3_outputs(658)));
    layer4_outputs(534) <= (layer3_outputs(2896)) and (layer3_outputs(3300));
    layer4_outputs(535) <= not(layer3_outputs(1667));
    layer4_outputs(536) <= not((layer3_outputs(882)) xor (layer3_outputs(2495)));
    layer4_outputs(537) <= not((layer3_outputs(1916)) or (layer3_outputs(2211)));
    layer4_outputs(538) <= (layer3_outputs(5214)) and not (layer3_outputs(2984));
    layer4_outputs(539) <= not((layer3_outputs(1707)) and (layer3_outputs(596)));
    layer4_outputs(540) <= layer3_outputs(3875);
    layer4_outputs(541) <= (layer3_outputs(6807)) xor (layer3_outputs(7354));
    layer4_outputs(542) <= not((layer3_outputs(5678)) and (layer3_outputs(3373)));
    layer4_outputs(543) <= (layer3_outputs(7274)) or (layer3_outputs(1600));
    layer4_outputs(544) <= layer3_outputs(2655);
    layer4_outputs(545) <= (layer3_outputs(3479)) and (layer3_outputs(748));
    layer4_outputs(546) <= (layer3_outputs(3473)) and (layer3_outputs(3356));
    layer4_outputs(547) <= (layer3_outputs(7487)) and (layer3_outputs(1214));
    layer4_outputs(548) <= layer3_outputs(2249);
    layer4_outputs(549) <= not(layer3_outputs(1347));
    layer4_outputs(550) <= not((layer3_outputs(974)) or (layer3_outputs(3014)));
    layer4_outputs(551) <= (layer3_outputs(3791)) and (layer3_outputs(605));
    layer4_outputs(552) <= layer3_outputs(5940);
    layer4_outputs(553) <= layer3_outputs(1473);
    layer4_outputs(554) <= not((layer3_outputs(1400)) or (layer3_outputs(2081)));
    layer4_outputs(555) <= not(layer3_outputs(5126));
    layer4_outputs(556) <= not((layer3_outputs(4981)) xor (layer3_outputs(2948)));
    layer4_outputs(557) <= (layer3_outputs(1162)) and not (layer3_outputs(4958));
    layer4_outputs(558) <= not(layer3_outputs(176)) or (layer3_outputs(2933));
    layer4_outputs(559) <= not(layer3_outputs(6043));
    layer4_outputs(560) <= not((layer3_outputs(1969)) or (layer3_outputs(3725)));
    layer4_outputs(561) <= layer3_outputs(3616);
    layer4_outputs(562) <= (layer3_outputs(6159)) or (layer3_outputs(805));
    layer4_outputs(563) <= layer3_outputs(7219);
    layer4_outputs(564) <= layer3_outputs(2980);
    layer4_outputs(565) <= layer3_outputs(3820);
    layer4_outputs(566) <= not(layer3_outputs(2699));
    layer4_outputs(567) <= layer3_outputs(6604);
    layer4_outputs(568) <= not(layer3_outputs(1332));
    layer4_outputs(569) <= not(layer3_outputs(5856)) or (layer3_outputs(6542));
    layer4_outputs(570) <= not((layer3_outputs(3321)) and (layer3_outputs(7073)));
    layer4_outputs(571) <= not(layer3_outputs(5038));
    layer4_outputs(572) <= not(layer3_outputs(2825));
    layer4_outputs(573) <= not(layer3_outputs(3889));
    layer4_outputs(574) <= not(layer3_outputs(2730));
    layer4_outputs(575) <= not(layer3_outputs(1830));
    layer4_outputs(576) <= layer3_outputs(3817);
    layer4_outputs(577) <= (layer3_outputs(5718)) or (layer3_outputs(6810));
    layer4_outputs(578) <= not(layer3_outputs(5046));
    layer4_outputs(579) <= not(layer3_outputs(346)) or (layer3_outputs(4011));
    layer4_outputs(580) <= not((layer3_outputs(277)) xor (layer3_outputs(7313)));
    layer4_outputs(581) <= (layer3_outputs(6890)) and not (layer3_outputs(2995));
    layer4_outputs(582) <= not(layer3_outputs(5492));
    layer4_outputs(583) <= layer3_outputs(6624);
    layer4_outputs(584) <= not(layer3_outputs(6185));
    layer4_outputs(585) <= not((layer3_outputs(5202)) or (layer3_outputs(5230)));
    layer4_outputs(586) <= layer3_outputs(4100);
    layer4_outputs(587) <= layer3_outputs(3473);
    layer4_outputs(588) <= layer3_outputs(587);
    layer4_outputs(589) <= (layer3_outputs(2339)) and not (layer3_outputs(100));
    layer4_outputs(590) <= not(layer3_outputs(327));
    layer4_outputs(591) <= not(layer3_outputs(6432));
    layer4_outputs(592) <= not(layer3_outputs(4497));
    layer4_outputs(593) <= not(layer3_outputs(4141));
    layer4_outputs(594) <= not(layer3_outputs(5468));
    layer4_outputs(595) <= (layer3_outputs(1206)) xor (layer3_outputs(5577));
    layer4_outputs(596) <= (layer3_outputs(7248)) and not (layer3_outputs(4910));
    layer4_outputs(597) <= not(layer3_outputs(2648));
    layer4_outputs(598) <= layer3_outputs(827);
    layer4_outputs(599) <= not(layer3_outputs(5300)) or (layer3_outputs(988));
    layer4_outputs(600) <= not(layer3_outputs(1086));
    layer4_outputs(601) <= (layer3_outputs(3621)) and not (layer3_outputs(1126));
    layer4_outputs(602) <= (layer3_outputs(4400)) xor (layer3_outputs(1605));
    layer4_outputs(603) <= layer3_outputs(6956);
    layer4_outputs(604) <= layer3_outputs(2886);
    layer4_outputs(605) <= not(layer3_outputs(5651));
    layer4_outputs(606) <= layer3_outputs(4768);
    layer4_outputs(607) <= not((layer3_outputs(1277)) or (layer3_outputs(1111)));
    layer4_outputs(608) <= (layer3_outputs(6501)) and not (layer3_outputs(6002));
    layer4_outputs(609) <= (layer3_outputs(6404)) and not (layer3_outputs(3085));
    layer4_outputs(610) <= layer3_outputs(5188);
    layer4_outputs(611) <= (layer3_outputs(2571)) xor (layer3_outputs(7270));
    layer4_outputs(612) <= layer3_outputs(4461);
    layer4_outputs(613) <= not(layer3_outputs(1194)) or (layer3_outputs(7182));
    layer4_outputs(614) <= not(layer3_outputs(1619)) or (layer3_outputs(268));
    layer4_outputs(615) <= not(layer3_outputs(549)) or (layer3_outputs(6936));
    layer4_outputs(616) <= not(layer3_outputs(4548)) or (layer3_outputs(4600));
    layer4_outputs(617) <= layer3_outputs(7443);
    layer4_outputs(618) <= layer3_outputs(741);
    layer4_outputs(619) <= layer3_outputs(1771);
    layer4_outputs(620) <= not(layer3_outputs(7619));
    layer4_outputs(621) <= layer3_outputs(157);
    layer4_outputs(622) <= (layer3_outputs(6375)) and (layer3_outputs(2800));
    layer4_outputs(623) <= layer3_outputs(1019);
    layer4_outputs(624) <= not(layer3_outputs(6699));
    layer4_outputs(625) <= layer3_outputs(4341);
    layer4_outputs(626) <= (layer3_outputs(3925)) xor (layer3_outputs(7165));
    layer4_outputs(627) <= not(layer3_outputs(5383));
    layer4_outputs(628) <= '1';
    layer4_outputs(629) <= not(layer3_outputs(7238));
    layer4_outputs(630) <= (layer3_outputs(2448)) and (layer3_outputs(7172));
    layer4_outputs(631) <= layer3_outputs(7079);
    layer4_outputs(632) <= not(layer3_outputs(7009));
    layer4_outputs(633) <= layer3_outputs(2830);
    layer4_outputs(634) <= (layer3_outputs(3442)) xor (layer3_outputs(5279));
    layer4_outputs(635) <= layer3_outputs(4916);
    layer4_outputs(636) <= (layer3_outputs(6537)) xor (layer3_outputs(2663));
    layer4_outputs(637) <= layer3_outputs(5569);
    layer4_outputs(638) <= layer3_outputs(2583);
    layer4_outputs(639) <= (layer3_outputs(6459)) or (layer3_outputs(5245));
    layer4_outputs(640) <= layer3_outputs(15);
    layer4_outputs(641) <= layer3_outputs(4253);
    layer4_outputs(642) <= (layer3_outputs(2904)) xor (layer3_outputs(130));
    layer4_outputs(643) <= not(layer3_outputs(3456));
    layer4_outputs(644) <= not((layer3_outputs(6602)) xor (layer3_outputs(1176)));
    layer4_outputs(645) <= not(layer3_outputs(5353));
    layer4_outputs(646) <= (layer3_outputs(1111)) or (layer3_outputs(7665));
    layer4_outputs(647) <= layer3_outputs(3591);
    layer4_outputs(648) <= not((layer3_outputs(7411)) and (layer3_outputs(6090)));
    layer4_outputs(649) <= not(layer3_outputs(3366));
    layer4_outputs(650) <= not((layer3_outputs(112)) and (layer3_outputs(1544)));
    layer4_outputs(651) <= layer3_outputs(5211);
    layer4_outputs(652) <= (layer3_outputs(5418)) or (layer3_outputs(3907));
    layer4_outputs(653) <= layer3_outputs(5645);
    layer4_outputs(654) <= layer3_outputs(248);
    layer4_outputs(655) <= layer3_outputs(3309);
    layer4_outputs(656) <= not(layer3_outputs(5706)) or (layer3_outputs(3166));
    layer4_outputs(657) <= layer3_outputs(332);
    layer4_outputs(658) <= (layer3_outputs(7629)) and not (layer3_outputs(5912));
    layer4_outputs(659) <= not(layer3_outputs(3416));
    layer4_outputs(660) <= not((layer3_outputs(5277)) and (layer3_outputs(5298)));
    layer4_outputs(661) <= '0';
    layer4_outputs(662) <= layer3_outputs(321);
    layer4_outputs(663) <= not((layer3_outputs(1474)) xor (layer3_outputs(4106)));
    layer4_outputs(664) <= not(layer3_outputs(7444));
    layer4_outputs(665) <= layer3_outputs(5994);
    layer4_outputs(666) <= layer3_outputs(7107);
    layer4_outputs(667) <= not(layer3_outputs(6210)) or (layer3_outputs(1355));
    layer4_outputs(668) <= layer3_outputs(5420);
    layer4_outputs(669) <= (layer3_outputs(2860)) and not (layer3_outputs(2466));
    layer4_outputs(670) <= layer3_outputs(2572);
    layer4_outputs(671) <= not(layer3_outputs(1786));
    layer4_outputs(672) <= not(layer3_outputs(3667));
    layer4_outputs(673) <= layer3_outputs(5885);
    layer4_outputs(674) <= layer3_outputs(7582);
    layer4_outputs(675) <= '0';
    layer4_outputs(676) <= not(layer3_outputs(7637)) or (layer3_outputs(523));
    layer4_outputs(677) <= '0';
    layer4_outputs(678) <= not(layer3_outputs(3788));
    layer4_outputs(679) <= not((layer3_outputs(3988)) and (layer3_outputs(4205)));
    layer4_outputs(680) <= not(layer3_outputs(5128));
    layer4_outputs(681) <= layer3_outputs(5165);
    layer4_outputs(682) <= not(layer3_outputs(6873));
    layer4_outputs(683) <= (layer3_outputs(2606)) and not (layer3_outputs(4119));
    layer4_outputs(684) <= (layer3_outputs(2743)) and not (layer3_outputs(4633));
    layer4_outputs(685) <= not(layer3_outputs(3959));
    layer4_outputs(686) <= not(layer3_outputs(1011));
    layer4_outputs(687) <= (layer3_outputs(1964)) and not (layer3_outputs(6849));
    layer4_outputs(688) <= not(layer3_outputs(617));
    layer4_outputs(689) <= layer3_outputs(2009);
    layer4_outputs(690) <= (layer3_outputs(3078)) or (layer3_outputs(2355));
    layer4_outputs(691) <= not(layer3_outputs(7374));
    layer4_outputs(692) <= not(layer3_outputs(1809));
    layer4_outputs(693) <= layer3_outputs(4467);
    layer4_outputs(694) <= layer3_outputs(5958);
    layer4_outputs(695) <= not((layer3_outputs(4833)) xor (layer3_outputs(64)));
    layer4_outputs(696) <= not(layer3_outputs(4540));
    layer4_outputs(697) <= layer3_outputs(6119);
    layer4_outputs(698) <= not(layer3_outputs(3048));
    layer4_outputs(699) <= (layer3_outputs(5337)) and (layer3_outputs(4269));
    layer4_outputs(700) <= (layer3_outputs(4037)) and (layer3_outputs(984));
    layer4_outputs(701) <= not(layer3_outputs(5541)) or (layer3_outputs(5722));
    layer4_outputs(702) <= not((layer3_outputs(2541)) xor (layer3_outputs(3758)));
    layer4_outputs(703) <= (layer3_outputs(4589)) and not (layer3_outputs(48));
    layer4_outputs(704) <= (layer3_outputs(3579)) or (layer3_outputs(6647));
    layer4_outputs(705) <= not(layer3_outputs(1041));
    layer4_outputs(706) <= not(layer3_outputs(6810));
    layer4_outputs(707) <= layer3_outputs(5973);
    layer4_outputs(708) <= not(layer3_outputs(4875)) or (layer3_outputs(5886));
    layer4_outputs(709) <= not((layer3_outputs(2600)) xor (layer3_outputs(4212)));
    layer4_outputs(710) <= not((layer3_outputs(2347)) xor (layer3_outputs(5155)));
    layer4_outputs(711) <= (layer3_outputs(2008)) and not (layer3_outputs(2962));
    layer4_outputs(712) <= (layer3_outputs(244)) and (layer3_outputs(3710));
    layer4_outputs(713) <= not(layer3_outputs(6769));
    layer4_outputs(714) <= layer3_outputs(7162);
    layer4_outputs(715) <= layer3_outputs(368);
    layer4_outputs(716) <= not((layer3_outputs(4672)) and (layer3_outputs(2579)));
    layer4_outputs(717) <= (layer3_outputs(6094)) and (layer3_outputs(4817));
    layer4_outputs(718) <= layer3_outputs(1800);
    layer4_outputs(719) <= layer3_outputs(6115);
    layer4_outputs(720) <= not(layer3_outputs(6169));
    layer4_outputs(721) <= layer3_outputs(7640);
    layer4_outputs(722) <= (layer3_outputs(1951)) or (layer3_outputs(6462));
    layer4_outputs(723) <= not(layer3_outputs(6559));
    layer4_outputs(724) <= (layer3_outputs(5366)) or (layer3_outputs(2804));
    layer4_outputs(725) <= layer3_outputs(1529);
    layer4_outputs(726) <= not(layer3_outputs(3268));
    layer4_outputs(727) <= not(layer3_outputs(3091));
    layer4_outputs(728) <= not(layer3_outputs(893));
    layer4_outputs(729) <= layer3_outputs(6148);
    layer4_outputs(730) <= not((layer3_outputs(4170)) and (layer3_outputs(6121)));
    layer4_outputs(731) <= (layer3_outputs(57)) or (layer3_outputs(5376));
    layer4_outputs(732) <= not((layer3_outputs(4236)) and (layer3_outputs(2472)));
    layer4_outputs(733) <= not(layer3_outputs(6020));
    layer4_outputs(734) <= (layer3_outputs(5890)) and not (layer3_outputs(3894));
    layer4_outputs(735) <= not(layer3_outputs(5924));
    layer4_outputs(736) <= layer3_outputs(7506);
    layer4_outputs(737) <= not(layer3_outputs(178));
    layer4_outputs(738) <= (layer3_outputs(1223)) xor (layer3_outputs(6653));
    layer4_outputs(739) <= layer3_outputs(6481);
    layer4_outputs(740) <= not(layer3_outputs(1524)) or (layer3_outputs(2475));
    layer4_outputs(741) <= (layer3_outputs(14)) and not (layer3_outputs(4605));
    layer4_outputs(742) <= not(layer3_outputs(3278));
    layer4_outputs(743) <= not(layer3_outputs(1028)) or (layer3_outputs(5960));
    layer4_outputs(744) <= not(layer3_outputs(7517));
    layer4_outputs(745) <= not((layer3_outputs(6070)) or (layer3_outputs(4305)));
    layer4_outputs(746) <= not(layer3_outputs(4853)) or (layer3_outputs(3861));
    layer4_outputs(747) <= (layer3_outputs(5019)) or (layer3_outputs(5306));
    layer4_outputs(748) <= '0';
    layer4_outputs(749) <= not((layer3_outputs(659)) xor (layer3_outputs(7186)));
    layer4_outputs(750) <= not((layer3_outputs(942)) xor (layer3_outputs(4431)));
    layer4_outputs(751) <= (layer3_outputs(5361)) xor (layer3_outputs(6828));
    layer4_outputs(752) <= layer3_outputs(4163);
    layer4_outputs(753) <= not((layer3_outputs(1778)) and (layer3_outputs(6083)));
    layer4_outputs(754) <= (layer3_outputs(3138)) and not (layer3_outputs(2864));
    layer4_outputs(755) <= layer3_outputs(421);
    layer4_outputs(756) <= not(layer3_outputs(583));
    layer4_outputs(757) <= (layer3_outputs(7561)) and not (layer3_outputs(4460));
    layer4_outputs(758) <= layer3_outputs(6001);
    layer4_outputs(759) <= not(layer3_outputs(3300));
    layer4_outputs(760) <= (layer3_outputs(5829)) and not (layer3_outputs(3724));
    layer4_outputs(761) <= layer3_outputs(7674);
    layer4_outputs(762) <= (layer3_outputs(1519)) and (layer3_outputs(6627));
    layer4_outputs(763) <= (layer3_outputs(1187)) and (layer3_outputs(7633));
    layer4_outputs(764) <= (layer3_outputs(1070)) xor (layer3_outputs(191));
    layer4_outputs(765) <= not(layer3_outputs(568)) or (layer3_outputs(7524));
    layer4_outputs(766) <= not(layer3_outputs(5400));
    layer4_outputs(767) <= (layer3_outputs(379)) and not (layer3_outputs(1920));
    layer4_outputs(768) <= layer3_outputs(6874);
    layer4_outputs(769) <= (layer3_outputs(5520)) and not (layer3_outputs(5053));
    layer4_outputs(770) <= (layer3_outputs(552)) and (layer3_outputs(3994));
    layer4_outputs(771) <= layer3_outputs(3292);
    layer4_outputs(772) <= layer3_outputs(4015);
    layer4_outputs(773) <= not(layer3_outputs(7567));
    layer4_outputs(774) <= not(layer3_outputs(3010)) or (layer3_outputs(2890));
    layer4_outputs(775) <= not(layer3_outputs(3559)) or (layer3_outputs(842));
    layer4_outputs(776) <= layer3_outputs(5638);
    layer4_outputs(777) <= not((layer3_outputs(5118)) and (layer3_outputs(3770)));
    layer4_outputs(778) <= '1';
    layer4_outputs(779) <= not(layer3_outputs(2482));
    layer4_outputs(780) <= not(layer3_outputs(5537)) or (layer3_outputs(3293));
    layer4_outputs(781) <= layer3_outputs(2071);
    layer4_outputs(782) <= not(layer3_outputs(5058));
    layer4_outputs(783) <= not(layer3_outputs(7596)) or (layer3_outputs(4039));
    layer4_outputs(784) <= not(layer3_outputs(317));
    layer4_outputs(785) <= not(layer3_outputs(5281)) or (layer3_outputs(3544));
    layer4_outputs(786) <= (layer3_outputs(4047)) or (layer3_outputs(1245));
    layer4_outputs(787) <= (layer3_outputs(1316)) or (layer3_outputs(1944));
    layer4_outputs(788) <= layer3_outputs(3928);
    layer4_outputs(789) <= not(layer3_outputs(6771));
    layer4_outputs(790) <= layer3_outputs(6111);
    layer4_outputs(791) <= not(layer3_outputs(6777)) or (layer3_outputs(646));
    layer4_outputs(792) <= layer3_outputs(182);
    layer4_outputs(793) <= not(layer3_outputs(4173));
    layer4_outputs(794) <= layer3_outputs(4286);
    layer4_outputs(795) <= not(layer3_outputs(6619));
    layer4_outputs(796) <= (layer3_outputs(4894)) and (layer3_outputs(6649));
    layer4_outputs(797) <= (layer3_outputs(3900)) and not (layer3_outputs(4022));
    layer4_outputs(798) <= not(layer3_outputs(5231));
    layer4_outputs(799) <= not(layer3_outputs(7066));
    layer4_outputs(800) <= not(layer3_outputs(6070));
    layer4_outputs(801) <= (layer3_outputs(2694)) and not (layer3_outputs(314));
    layer4_outputs(802) <= not(layer3_outputs(6709));
    layer4_outputs(803) <= layer3_outputs(428);
    layer4_outputs(804) <= not(layer3_outputs(3164)) or (layer3_outputs(6632));
    layer4_outputs(805) <= not((layer3_outputs(2076)) xor (layer3_outputs(4611)));
    layer4_outputs(806) <= not(layer3_outputs(4884));
    layer4_outputs(807) <= not(layer3_outputs(2233));
    layer4_outputs(808) <= layer3_outputs(6703);
    layer4_outputs(809) <= (layer3_outputs(354)) and not (layer3_outputs(4588));
    layer4_outputs(810) <= not(layer3_outputs(7023)) or (layer3_outputs(3985));
    layer4_outputs(811) <= not(layer3_outputs(560)) or (layer3_outputs(880));
    layer4_outputs(812) <= not((layer3_outputs(319)) or (layer3_outputs(3917)));
    layer4_outputs(813) <= not((layer3_outputs(7532)) xor (layer3_outputs(5227)));
    layer4_outputs(814) <= not((layer3_outputs(3946)) xor (layer3_outputs(3737)));
    layer4_outputs(815) <= not(layer3_outputs(6488));
    layer4_outputs(816) <= (layer3_outputs(54)) and (layer3_outputs(6408));
    layer4_outputs(817) <= (layer3_outputs(2112)) and (layer3_outputs(1270));
    layer4_outputs(818) <= not(layer3_outputs(3036));
    layer4_outputs(819) <= not(layer3_outputs(4428));
    layer4_outputs(820) <= layer3_outputs(1173);
    layer4_outputs(821) <= not(layer3_outputs(4003)) or (layer3_outputs(1132));
    layer4_outputs(822) <= layer3_outputs(109);
    layer4_outputs(823) <= (layer3_outputs(5457)) and not (layer3_outputs(6929));
    layer4_outputs(824) <= layer3_outputs(5318);
    layer4_outputs(825) <= layer3_outputs(7641);
    layer4_outputs(826) <= not(layer3_outputs(906));
    layer4_outputs(827) <= not(layer3_outputs(2610));
    layer4_outputs(828) <= not((layer3_outputs(5604)) or (layer3_outputs(7233)));
    layer4_outputs(829) <= not(layer3_outputs(6477)) or (layer3_outputs(5791));
    layer4_outputs(830) <= not(layer3_outputs(1909));
    layer4_outputs(831) <= not(layer3_outputs(1640));
    layer4_outputs(832) <= not((layer3_outputs(4669)) or (layer3_outputs(844)));
    layer4_outputs(833) <= layer3_outputs(557);
    layer4_outputs(834) <= layer3_outputs(4915);
    layer4_outputs(835) <= (layer3_outputs(863)) and not (layer3_outputs(4935));
    layer4_outputs(836) <= not(layer3_outputs(4064));
    layer4_outputs(837) <= not(layer3_outputs(6739)) or (layer3_outputs(4758));
    layer4_outputs(838) <= (layer3_outputs(2269)) xor (layer3_outputs(5675));
    layer4_outputs(839) <= layer3_outputs(6251);
    layer4_outputs(840) <= not(layer3_outputs(233));
    layer4_outputs(841) <= layer3_outputs(4656);
    layer4_outputs(842) <= not(layer3_outputs(6955)) or (layer3_outputs(3347));
    layer4_outputs(843) <= (layer3_outputs(7032)) and not (layer3_outputs(535));
    layer4_outputs(844) <= not((layer3_outputs(3481)) and (layer3_outputs(5859)));
    layer4_outputs(845) <= not((layer3_outputs(7596)) xor (layer3_outputs(7108)));
    layer4_outputs(846) <= not(layer3_outputs(1051)) or (layer3_outputs(1091));
    layer4_outputs(847) <= layer3_outputs(7520);
    layer4_outputs(848) <= (layer3_outputs(5370)) and (layer3_outputs(1565));
    layer4_outputs(849) <= not(layer3_outputs(2703));
    layer4_outputs(850) <= not(layer3_outputs(109));
    layer4_outputs(851) <= not((layer3_outputs(4236)) or (layer3_outputs(2045)));
    layer4_outputs(852) <= not(layer3_outputs(2679));
    layer4_outputs(853) <= not(layer3_outputs(759));
    layer4_outputs(854) <= layer3_outputs(2361);
    layer4_outputs(855) <= not(layer3_outputs(2208));
    layer4_outputs(856) <= not((layer3_outputs(6263)) and (layer3_outputs(5395)));
    layer4_outputs(857) <= (layer3_outputs(2147)) and (layer3_outputs(5389));
    layer4_outputs(858) <= layer3_outputs(5497);
    layer4_outputs(859) <= (layer3_outputs(4036)) and not (layer3_outputs(1445));
    layer4_outputs(860) <= not((layer3_outputs(914)) and (layer3_outputs(3919)));
    layer4_outputs(861) <= not(layer3_outputs(5212)) or (layer3_outputs(5895));
    layer4_outputs(862) <= not(layer3_outputs(5373));
    layer4_outputs(863) <= (layer3_outputs(4651)) and not (layer3_outputs(5504));
    layer4_outputs(864) <= (layer3_outputs(4206)) and not (layer3_outputs(6702));
    layer4_outputs(865) <= not(layer3_outputs(3516));
    layer4_outputs(866) <= not(layer3_outputs(2490));
    layer4_outputs(867) <= (layer3_outputs(3439)) and not (layer3_outputs(7292));
    layer4_outputs(868) <= layer3_outputs(933);
    layer4_outputs(869) <= layer3_outputs(2172);
    layer4_outputs(870) <= not(layer3_outputs(5523)) or (layer3_outputs(6551));
    layer4_outputs(871) <= layer3_outputs(3169);
    layer4_outputs(872) <= layer3_outputs(4386);
    layer4_outputs(873) <= (layer3_outputs(3724)) xor (layer3_outputs(2695));
    layer4_outputs(874) <= not((layer3_outputs(4291)) or (layer3_outputs(7146)));
    layer4_outputs(875) <= not(layer3_outputs(6240));
    layer4_outputs(876) <= (layer3_outputs(3940)) and not (layer3_outputs(479));
    layer4_outputs(877) <= not(layer3_outputs(7601));
    layer4_outputs(878) <= layer3_outputs(7361);
    layer4_outputs(879) <= layer3_outputs(6103);
    layer4_outputs(880) <= layer3_outputs(4489);
    layer4_outputs(881) <= (layer3_outputs(2307)) and (layer3_outputs(6014));
    layer4_outputs(882) <= not((layer3_outputs(4720)) xor (layer3_outputs(2108)));
    layer4_outputs(883) <= (layer3_outputs(3683)) or (layer3_outputs(209));
    layer4_outputs(884) <= layer3_outputs(3859);
    layer4_outputs(885) <= layer3_outputs(6555);
    layer4_outputs(886) <= layer3_outputs(7650);
    layer4_outputs(887) <= layer3_outputs(2294);
    layer4_outputs(888) <= (layer3_outputs(1232)) and not (layer3_outputs(4861));
    layer4_outputs(889) <= not(layer3_outputs(2274));
    layer4_outputs(890) <= layer3_outputs(2369);
    layer4_outputs(891) <= (layer3_outputs(857)) and not (layer3_outputs(7113));
    layer4_outputs(892) <= (layer3_outputs(3411)) and not (layer3_outputs(7561));
    layer4_outputs(893) <= layer3_outputs(5857);
    layer4_outputs(894) <= not((layer3_outputs(4537)) or (layer3_outputs(4539)));
    layer4_outputs(895) <= layer3_outputs(103);
    layer4_outputs(896) <= not(layer3_outputs(4020));
    layer4_outputs(897) <= layer3_outputs(6298);
    layer4_outputs(898) <= not(layer3_outputs(1321));
    layer4_outputs(899) <= not(layer3_outputs(4330));
    layer4_outputs(900) <= not((layer3_outputs(3705)) and (layer3_outputs(3818)));
    layer4_outputs(901) <= (layer3_outputs(5884)) and not (layer3_outputs(2841));
    layer4_outputs(902) <= not(layer3_outputs(2133)) or (layer3_outputs(5626));
    layer4_outputs(903) <= not((layer3_outputs(1242)) xor (layer3_outputs(5033)));
    layer4_outputs(904) <= (layer3_outputs(1493)) and not (layer3_outputs(5176));
    layer4_outputs(905) <= layer3_outputs(2136);
    layer4_outputs(906) <= not((layer3_outputs(4371)) or (layer3_outputs(7069)));
    layer4_outputs(907) <= (layer3_outputs(3668)) and not (layer3_outputs(2873));
    layer4_outputs(908) <= layer3_outputs(6249);
    layer4_outputs(909) <= '0';
    layer4_outputs(910) <= layer3_outputs(6129);
    layer4_outputs(911) <= (layer3_outputs(2011)) and not (layer3_outputs(4972));
    layer4_outputs(912) <= (layer3_outputs(7404)) and not (layer3_outputs(2084));
    layer4_outputs(913) <= not(layer3_outputs(2049));
    layer4_outputs(914) <= '0';
    layer4_outputs(915) <= layer3_outputs(5657);
    layer4_outputs(916) <= layer3_outputs(5862);
    layer4_outputs(917) <= not(layer3_outputs(7014));
    layer4_outputs(918) <= not((layer3_outputs(6425)) xor (layer3_outputs(6757)));
    layer4_outputs(919) <= (layer3_outputs(1927)) and not (layer3_outputs(5527));
    layer4_outputs(920) <= not(layer3_outputs(1943));
    layer4_outputs(921) <= not(layer3_outputs(7279));
    layer4_outputs(922) <= not(layer3_outputs(5316));
    layer4_outputs(923) <= layer3_outputs(764);
    layer4_outputs(924) <= (layer3_outputs(1016)) xor (layer3_outputs(6764));
    layer4_outputs(925) <= (layer3_outputs(4820)) and not (layer3_outputs(6195));
    layer4_outputs(926) <= '1';
    layer4_outputs(927) <= layer3_outputs(6585);
    layer4_outputs(928) <= not((layer3_outputs(2088)) or (layer3_outputs(4913)));
    layer4_outputs(929) <= not((layer3_outputs(7371)) and (layer3_outputs(5629)));
    layer4_outputs(930) <= layer3_outputs(3966);
    layer4_outputs(931) <= layer3_outputs(3369);
    layer4_outputs(932) <= layer3_outputs(1367);
    layer4_outputs(933) <= not(layer3_outputs(5043));
    layer4_outputs(934) <= not(layer3_outputs(2720));
    layer4_outputs(935) <= not(layer3_outputs(6894)) or (layer3_outputs(6454));
    layer4_outputs(936) <= layer3_outputs(5179);
    layer4_outputs(937) <= (layer3_outputs(6239)) and (layer3_outputs(2294));
    layer4_outputs(938) <= not((layer3_outputs(4324)) and (layer3_outputs(4054)));
    layer4_outputs(939) <= not(layer3_outputs(3995));
    layer4_outputs(940) <= not((layer3_outputs(7215)) xor (layer3_outputs(2503)));
    layer4_outputs(941) <= (layer3_outputs(6823)) xor (layer3_outputs(4192));
    layer4_outputs(942) <= not((layer3_outputs(5149)) and (layer3_outputs(4434)));
    layer4_outputs(943) <= not(layer3_outputs(3567));
    layer4_outputs(944) <= layer3_outputs(4569);
    layer4_outputs(945) <= not(layer3_outputs(1419));
    layer4_outputs(946) <= not(layer3_outputs(6534));
    layer4_outputs(947) <= not(layer3_outputs(5302));
    layer4_outputs(948) <= not(layer3_outputs(6182));
    layer4_outputs(949) <= layer3_outputs(4955);
    layer4_outputs(950) <= '1';
    layer4_outputs(951) <= '0';
    layer4_outputs(952) <= (layer3_outputs(5963)) and not (layer3_outputs(5108));
    layer4_outputs(953) <= (layer3_outputs(4653)) and not (layer3_outputs(6429));
    layer4_outputs(954) <= (layer3_outputs(2604)) and (layer3_outputs(60));
    layer4_outputs(955) <= (layer3_outputs(5732)) and not (layer3_outputs(3451));
    layer4_outputs(956) <= layer3_outputs(493);
    layer4_outputs(957) <= not(layer3_outputs(6554));
    layer4_outputs(958) <= layer3_outputs(6388);
    layer4_outputs(959) <= (layer3_outputs(1067)) and (layer3_outputs(3457));
    layer4_outputs(960) <= (layer3_outputs(2719)) or (layer3_outputs(6439));
    layer4_outputs(961) <= not(layer3_outputs(6013));
    layer4_outputs(962) <= not(layer3_outputs(3192));
    layer4_outputs(963) <= layer3_outputs(5344);
    layer4_outputs(964) <= layer3_outputs(1021);
    layer4_outputs(965) <= not((layer3_outputs(6021)) and (layer3_outputs(3336)));
    layer4_outputs(966) <= layer3_outputs(1479);
    layer4_outputs(967) <= layer3_outputs(5636);
    layer4_outputs(968) <= not(layer3_outputs(3303)) or (layer3_outputs(3653));
    layer4_outputs(969) <= (layer3_outputs(4389)) or (layer3_outputs(3013));
    layer4_outputs(970) <= layer3_outputs(1446);
    layer4_outputs(971) <= not(layer3_outputs(7046));
    layer4_outputs(972) <= (layer3_outputs(5652)) xor (layer3_outputs(4556));
    layer4_outputs(973) <= (layer3_outputs(6900)) and (layer3_outputs(3355));
    layer4_outputs(974) <= (layer3_outputs(4792)) and (layer3_outputs(7480));
    layer4_outputs(975) <= layer3_outputs(5549);
    layer4_outputs(976) <= not(layer3_outputs(5970)) or (layer3_outputs(6738));
    layer4_outputs(977) <= not(layer3_outputs(3948));
    layer4_outputs(978) <= not(layer3_outputs(4186));
    layer4_outputs(979) <= layer3_outputs(1630);
    layer4_outputs(980) <= not(layer3_outputs(5007));
    layer4_outputs(981) <= layer3_outputs(5954);
    layer4_outputs(982) <= not(layer3_outputs(6219));
    layer4_outputs(983) <= layer3_outputs(964);
    layer4_outputs(984) <= not((layer3_outputs(6432)) xor (layer3_outputs(4676)));
    layer4_outputs(985) <= not((layer3_outputs(1562)) or (layer3_outputs(2727)));
    layer4_outputs(986) <= not((layer3_outputs(4944)) or (layer3_outputs(1844)));
    layer4_outputs(987) <= layer3_outputs(410);
    layer4_outputs(988) <= (layer3_outputs(6131)) and not (layer3_outputs(7205));
    layer4_outputs(989) <= not(layer3_outputs(3942)) or (layer3_outputs(2609));
    layer4_outputs(990) <= layer3_outputs(6915);
    layer4_outputs(991) <= not(layer3_outputs(1415));
    layer4_outputs(992) <= layer3_outputs(5005);
    layer4_outputs(993) <= (layer3_outputs(6260)) and not (layer3_outputs(230));
    layer4_outputs(994) <= (layer3_outputs(7208)) xor (layer3_outputs(2461));
    layer4_outputs(995) <= layer3_outputs(7624);
    layer4_outputs(996) <= (layer3_outputs(2877)) and not (layer3_outputs(2346));
    layer4_outputs(997) <= not(layer3_outputs(3006));
    layer4_outputs(998) <= layer3_outputs(978);
    layer4_outputs(999) <= (layer3_outputs(7598)) or (layer3_outputs(1617));
    layer4_outputs(1000) <= (layer3_outputs(6173)) and (layer3_outputs(58));
    layer4_outputs(1001) <= (layer3_outputs(7165)) xor (layer3_outputs(6803));
    layer4_outputs(1002) <= layer3_outputs(6999);
    layer4_outputs(1003) <= layer3_outputs(6287);
    layer4_outputs(1004) <= not(layer3_outputs(643));
    layer4_outputs(1005) <= not(layer3_outputs(2314));
    layer4_outputs(1006) <= not(layer3_outputs(6351));
    layer4_outputs(1007) <= not(layer3_outputs(5281));
    layer4_outputs(1008) <= not(layer3_outputs(1994));
    layer4_outputs(1009) <= (layer3_outputs(5337)) and not (layer3_outputs(5778));
    layer4_outputs(1010) <= layer3_outputs(3895);
    layer4_outputs(1011) <= not((layer3_outputs(4097)) and (layer3_outputs(632)));
    layer4_outputs(1012) <= not((layer3_outputs(7496)) and (layer3_outputs(4251)));
    layer4_outputs(1013) <= not(layer3_outputs(6330)) or (layer3_outputs(1836));
    layer4_outputs(1014) <= (layer3_outputs(960)) and not (layer3_outputs(966));
    layer4_outputs(1015) <= not((layer3_outputs(3708)) xor (layer3_outputs(7428)));
    layer4_outputs(1016) <= (layer3_outputs(2305)) and not (layer3_outputs(4607));
    layer4_outputs(1017) <= not(layer3_outputs(5990)) or (layer3_outputs(3052));
    layer4_outputs(1018) <= layer3_outputs(1910);
    layer4_outputs(1019) <= layer3_outputs(4120);
    layer4_outputs(1020) <= not((layer3_outputs(1995)) and (layer3_outputs(3404)));
    layer4_outputs(1021) <= (layer3_outputs(6019)) xor (layer3_outputs(3173));
    layer4_outputs(1022) <= not(layer3_outputs(2722));
    layer4_outputs(1023) <= layer3_outputs(7061);
    layer4_outputs(1024) <= not(layer3_outputs(4807));
    layer4_outputs(1025) <= not(layer3_outputs(4052));
    layer4_outputs(1026) <= not(layer3_outputs(2222));
    layer4_outputs(1027) <= layer3_outputs(5309);
    layer4_outputs(1028) <= layer3_outputs(6023);
    layer4_outputs(1029) <= not(layer3_outputs(7024));
    layer4_outputs(1030) <= not(layer3_outputs(7546)) or (layer3_outputs(3897));
    layer4_outputs(1031) <= layer3_outputs(5038);
    layer4_outputs(1032) <= (layer3_outputs(3505)) xor (layer3_outputs(7477));
    layer4_outputs(1033) <= not(layer3_outputs(1417)) or (layer3_outputs(4412));
    layer4_outputs(1034) <= not(layer3_outputs(5002)) or (layer3_outputs(613));
    layer4_outputs(1035) <= not(layer3_outputs(1782));
    layer4_outputs(1036) <= layer3_outputs(2530);
    layer4_outputs(1037) <= layer3_outputs(7104);
    layer4_outputs(1038) <= not(layer3_outputs(6986));
    layer4_outputs(1039) <= (layer3_outputs(1532)) xor (layer3_outputs(1272));
    layer4_outputs(1040) <= (layer3_outputs(1938)) or (layer3_outputs(232));
    layer4_outputs(1041) <= not(layer3_outputs(854));
    layer4_outputs(1042) <= layer3_outputs(652);
    layer4_outputs(1043) <= not(layer3_outputs(7486));
    layer4_outputs(1044) <= (layer3_outputs(4194)) and (layer3_outputs(4761));
    layer4_outputs(1045) <= layer3_outputs(4203);
    layer4_outputs(1046) <= layer3_outputs(6883);
    layer4_outputs(1047) <= (layer3_outputs(7268)) xor (layer3_outputs(433));
    layer4_outputs(1048) <= (layer3_outputs(6387)) or (layer3_outputs(6548));
    layer4_outputs(1049) <= not(layer3_outputs(2770));
    layer4_outputs(1050) <= (layer3_outputs(6067)) xor (layer3_outputs(597));
    layer4_outputs(1051) <= not(layer3_outputs(5369));
    layer4_outputs(1052) <= (layer3_outputs(7209)) and not (layer3_outputs(6223));
    layer4_outputs(1053) <= (layer3_outputs(1361)) xor (layer3_outputs(5292));
    layer4_outputs(1054) <= layer3_outputs(5943);
    layer4_outputs(1055) <= not(layer3_outputs(4417));
    layer4_outputs(1056) <= not((layer3_outputs(2865)) xor (layer3_outputs(2581)));
    layer4_outputs(1057) <= (layer3_outputs(3273)) and not (layer3_outputs(6890));
    layer4_outputs(1058) <= (layer3_outputs(2430)) xor (layer3_outputs(2321));
    layer4_outputs(1059) <= (layer3_outputs(1543)) and not (layer3_outputs(623));
    layer4_outputs(1060) <= layer3_outputs(1595);
    layer4_outputs(1061) <= not((layer3_outputs(2061)) or (layer3_outputs(395)));
    layer4_outputs(1062) <= not(layer3_outputs(1520));
    layer4_outputs(1063) <= not((layer3_outputs(3820)) or (layer3_outputs(2322)));
    layer4_outputs(1064) <= (layer3_outputs(3027)) and not (layer3_outputs(362));
    layer4_outputs(1065) <= (layer3_outputs(3900)) and (layer3_outputs(2055));
    layer4_outputs(1066) <= not(layer3_outputs(2335));
    layer4_outputs(1067) <= not(layer3_outputs(3514));
    layer4_outputs(1068) <= not((layer3_outputs(5612)) xor (layer3_outputs(2558)));
    layer4_outputs(1069) <= layer3_outputs(931);
    layer4_outputs(1070) <= layer3_outputs(7571);
    layer4_outputs(1071) <= layer3_outputs(3477);
    layer4_outputs(1072) <= not(layer3_outputs(6760));
    layer4_outputs(1073) <= (layer3_outputs(6392)) and not (layer3_outputs(4696));
    layer4_outputs(1074) <= not(layer3_outputs(5459)) or (layer3_outputs(6465));
    layer4_outputs(1075) <= not(layer3_outputs(5565)) or (layer3_outputs(2324));
    layer4_outputs(1076) <= not(layer3_outputs(469));
    layer4_outputs(1077) <= layer3_outputs(3746);
    layer4_outputs(1078) <= not(layer3_outputs(3687));
    layer4_outputs(1079) <= (layer3_outputs(82)) and (layer3_outputs(6174));
    layer4_outputs(1080) <= not(layer3_outputs(4491));
    layer4_outputs(1081) <= not(layer3_outputs(3898));
    layer4_outputs(1082) <= not(layer3_outputs(3332)) or (layer3_outputs(3234));
    layer4_outputs(1083) <= layer3_outputs(111);
    layer4_outputs(1084) <= (layer3_outputs(1825)) xor (layer3_outputs(100));
    layer4_outputs(1085) <= layer3_outputs(3444);
    layer4_outputs(1086) <= layer3_outputs(2075);
    layer4_outputs(1087) <= layer3_outputs(3227);
    layer4_outputs(1088) <= not(layer3_outputs(1796));
    layer4_outputs(1089) <= not(layer3_outputs(4050));
    layer4_outputs(1090) <= not((layer3_outputs(128)) and (layer3_outputs(2888)));
    layer4_outputs(1091) <= (layer3_outputs(4545)) xor (layer3_outputs(1780));
    layer4_outputs(1092) <= (layer3_outputs(1463)) and not (layer3_outputs(5336));
    layer4_outputs(1093) <= layer3_outputs(7290);
    layer4_outputs(1094) <= (layer3_outputs(2594)) xor (layer3_outputs(5355));
    layer4_outputs(1095) <= not(layer3_outputs(3381));
    layer4_outputs(1096) <= not((layer3_outputs(5213)) and (layer3_outputs(6116)));
    layer4_outputs(1097) <= (layer3_outputs(6027)) or (layer3_outputs(3993));
    layer4_outputs(1098) <= not(layer3_outputs(6400));
    layer4_outputs(1099) <= not(layer3_outputs(3160));
    layer4_outputs(1100) <= (layer3_outputs(6191)) xor (layer3_outputs(6931));
    layer4_outputs(1101) <= not(layer3_outputs(3423));
    layer4_outputs(1102) <= not(layer3_outputs(7542)) or (layer3_outputs(6557));
    layer4_outputs(1103) <= not((layer3_outputs(1065)) or (layer3_outputs(6060)));
    layer4_outputs(1104) <= not((layer3_outputs(5553)) xor (layer3_outputs(1201)));
    layer4_outputs(1105) <= layer3_outputs(7159);
    layer4_outputs(1106) <= not(layer3_outputs(829));
    layer4_outputs(1107) <= not(layer3_outputs(5283));
    layer4_outputs(1108) <= (layer3_outputs(734)) and not (layer3_outputs(7548));
    layer4_outputs(1109) <= not(layer3_outputs(6675));
    layer4_outputs(1110) <= not(layer3_outputs(7014));
    layer4_outputs(1111) <= not(layer3_outputs(7029));
    layer4_outputs(1112) <= (layer3_outputs(2840)) and not (layer3_outputs(6366));
    layer4_outputs(1113) <= not((layer3_outputs(4338)) xor (layer3_outputs(4383)));
    layer4_outputs(1114) <= (layer3_outputs(3961)) and not (layer3_outputs(1324));
    layer4_outputs(1115) <= (layer3_outputs(3211)) xor (layer3_outputs(4976));
    layer4_outputs(1116) <= (layer3_outputs(2365)) or (layer3_outputs(1217));
    layer4_outputs(1117) <= not(layer3_outputs(4355));
    layer4_outputs(1118) <= not(layer3_outputs(1057));
    layer4_outputs(1119) <= not(layer3_outputs(2553)) or (layer3_outputs(4609));
    layer4_outputs(1120) <= not((layer3_outputs(5425)) and (layer3_outputs(661)));
    layer4_outputs(1121) <= not((layer3_outputs(5550)) and (layer3_outputs(4698)));
    layer4_outputs(1122) <= (layer3_outputs(413)) and not (layer3_outputs(5342));
    layer4_outputs(1123) <= not(layer3_outputs(6937));
    layer4_outputs(1124) <= not(layer3_outputs(2570));
    layer4_outputs(1125) <= not((layer3_outputs(3393)) xor (layer3_outputs(2042)));
    layer4_outputs(1126) <= layer3_outputs(15);
    layer4_outputs(1127) <= (layer3_outputs(4513)) and not (layer3_outputs(1080));
    layer4_outputs(1128) <= not((layer3_outputs(3579)) or (layer3_outputs(1873)));
    layer4_outputs(1129) <= not(layer3_outputs(5844));
    layer4_outputs(1130) <= (layer3_outputs(1404)) and not (layer3_outputs(704));
    layer4_outputs(1131) <= not(layer3_outputs(961));
    layer4_outputs(1132) <= not(layer3_outputs(585));
    layer4_outputs(1133) <= layer3_outputs(4928);
    layer4_outputs(1134) <= not(layer3_outputs(6822));
    layer4_outputs(1135) <= not(layer3_outputs(2470));
    layer4_outputs(1136) <= layer3_outputs(4280);
    layer4_outputs(1137) <= not(layer3_outputs(5044)) or (layer3_outputs(2790));
    layer4_outputs(1138) <= layer3_outputs(1180);
    layer4_outputs(1139) <= not(layer3_outputs(204));
    layer4_outputs(1140) <= not((layer3_outputs(7394)) and (layer3_outputs(4733)));
    layer4_outputs(1141) <= not(layer3_outputs(7413));
    layer4_outputs(1142) <= not(layer3_outputs(1513)) or (layer3_outputs(3679));
    layer4_outputs(1143) <= layer3_outputs(2954);
    layer4_outputs(1144) <= '1';
    layer4_outputs(1145) <= not(layer3_outputs(5804)) or (layer3_outputs(1766));
    layer4_outputs(1146) <= not(layer3_outputs(2304));
    layer4_outputs(1147) <= not(layer3_outputs(1983));
    layer4_outputs(1148) <= not(layer3_outputs(2803));
    layer4_outputs(1149) <= not((layer3_outputs(3587)) xor (layer3_outputs(1983)));
    layer4_outputs(1150) <= (layer3_outputs(6310)) xor (layer3_outputs(4109));
    layer4_outputs(1151) <= not((layer3_outputs(6005)) or (layer3_outputs(3949)));
    layer4_outputs(1152) <= (layer3_outputs(5848)) and not (layer3_outputs(5219));
    layer4_outputs(1153) <= not((layer3_outputs(159)) or (layer3_outputs(3264)));
    layer4_outputs(1154) <= not((layer3_outputs(344)) and (layer3_outputs(7123)));
    layer4_outputs(1155) <= (layer3_outputs(343)) xor (layer3_outputs(4399));
    layer4_outputs(1156) <= (layer3_outputs(3166)) or (layer3_outputs(7453));
    layer4_outputs(1157) <= not(layer3_outputs(4287));
    layer4_outputs(1158) <= layer3_outputs(2575);
    layer4_outputs(1159) <= not((layer3_outputs(6124)) and (layer3_outputs(5067)));
    layer4_outputs(1160) <= layer3_outputs(6561);
    layer4_outputs(1161) <= not((layer3_outputs(2578)) or (layer3_outputs(4033)));
    layer4_outputs(1162) <= (layer3_outputs(1806)) xor (layer3_outputs(3793));
    layer4_outputs(1163) <= not(layer3_outputs(4091)) or (layer3_outputs(1500));
    layer4_outputs(1164) <= layer3_outputs(7116);
    layer4_outputs(1165) <= layer3_outputs(920);
    layer4_outputs(1166) <= not(layer3_outputs(7439));
    layer4_outputs(1167) <= '0';
    layer4_outputs(1168) <= not(layer3_outputs(5121));
    layer4_outputs(1169) <= not(layer3_outputs(5869));
    layer4_outputs(1170) <= not(layer3_outputs(4393));
    layer4_outputs(1171) <= layer3_outputs(1338);
    layer4_outputs(1172) <= not(layer3_outputs(1879));
    layer4_outputs(1173) <= layer3_outputs(5535);
    layer4_outputs(1174) <= not((layer3_outputs(2299)) xor (layer3_outputs(1592)));
    layer4_outputs(1175) <= not(layer3_outputs(3082));
    layer4_outputs(1176) <= not((layer3_outputs(3086)) xor (layer3_outputs(6416)));
    layer4_outputs(1177) <= (layer3_outputs(7133)) xor (layer3_outputs(2410));
    layer4_outputs(1178) <= (layer3_outputs(2746)) and not (layer3_outputs(6187));
    layer4_outputs(1179) <= layer3_outputs(4653);
    layer4_outputs(1180) <= not(layer3_outputs(659));
    layer4_outputs(1181) <= not((layer3_outputs(4356)) xor (layer3_outputs(4918)));
    layer4_outputs(1182) <= layer3_outputs(2141);
    layer4_outputs(1183) <= (layer3_outputs(1601)) and not (layer3_outputs(3534));
    layer4_outputs(1184) <= not((layer3_outputs(3018)) or (layer3_outputs(7015)));
    layer4_outputs(1185) <= not(layer3_outputs(3664));
    layer4_outputs(1186) <= not((layer3_outputs(4140)) xor (layer3_outputs(1864)));
    layer4_outputs(1187) <= not((layer3_outputs(7098)) and (layer3_outputs(6528)));
    layer4_outputs(1188) <= not(layer3_outputs(5302));
    layer4_outputs(1189) <= (layer3_outputs(4964)) and (layer3_outputs(4339));
    layer4_outputs(1190) <= layer3_outputs(563);
    layer4_outputs(1191) <= not(layer3_outputs(1857)) or (layer3_outputs(3193));
    layer4_outputs(1192) <= not((layer3_outputs(2479)) or (layer3_outputs(7447)));
    layer4_outputs(1193) <= not(layer3_outputs(2589)) or (layer3_outputs(2082));
    layer4_outputs(1194) <= not(layer3_outputs(3163));
    layer4_outputs(1195) <= layer3_outputs(881);
    layer4_outputs(1196) <= layer3_outputs(1753);
    layer4_outputs(1197) <= layer3_outputs(3067);
    layer4_outputs(1198) <= not(layer3_outputs(1682));
    layer4_outputs(1199) <= (layer3_outputs(7463)) and (layer3_outputs(5501));
    layer4_outputs(1200) <= not((layer3_outputs(6086)) xor (layer3_outputs(74)));
    layer4_outputs(1201) <= (layer3_outputs(2732)) and not (layer3_outputs(3666));
    layer4_outputs(1202) <= layer3_outputs(1810);
    layer4_outputs(1203) <= layer3_outputs(2074);
    layer4_outputs(1204) <= not((layer3_outputs(3522)) or (layer3_outputs(4183)));
    layer4_outputs(1205) <= layer3_outputs(2765);
    layer4_outputs(1206) <= (layer3_outputs(2147)) xor (layer3_outputs(3821));
    layer4_outputs(1207) <= not(layer3_outputs(5133));
    layer4_outputs(1208) <= not(layer3_outputs(3999));
    layer4_outputs(1209) <= layer3_outputs(5375);
    layer4_outputs(1210) <= (layer3_outputs(6383)) xor (layer3_outputs(500));
    layer4_outputs(1211) <= not(layer3_outputs(2502));
    layer4_outputs(1212) <= not((layer3_outputs(4713)) xor (layer3_outputs(2876)));
    layer4_outputs(1213) <= (layer3_outputs(2016)) and not (layer3_outputs(5515));
    layer4_outputs(1214) <= (layer3_outputs(1285)) and not (layer3_outputs(2121));
    layer4_outputs(1215) <= not((layer3_outputs(210)) xor (layer3_outputs(599)));
    layer4_outputs(1216) <= (layer3_outputs(7410)) and (layer3_outputs(3866));
    layer4_outputs(1217) <= layer3_outputs(2965);
    layer4_outputs(1218) <= not((layer3_outputs(3431)) and (layer3_outputs(2854)));
    layer4_outputs(1219) <= layer3_outputs(3112);
    layer4_outputs(1220) <= layer3_outputs(4504);
    layer4_outputs(1221) <= not(layer3_outputs(5432)) or (layer3_outputs(5103));
    layer4_outputs(1222) <= (layer3_outputs(160)) and not (layer3_outputs(2712));
    layer4_outputs(1223) <= not(layer3_outputs(859));
    layer4_outputs(1224) <= layer3_outputs(6878);
    layer4_outputs(1225) <= (layer3_outputs(4246)) or (layer3_outputs(1540));
    layer4_outputs(1226) <= not(layer3_outputs(2859)) or (layer3_outputs(2308));
    layer4_outputs(1227) <= (layer3_outputs(3625)) or (layer3_outputs(183));
    layer4_outputs(1228) <= not((layer3_outputs(1153)) and (layer3_outputs(3394)));
    layer4_outputs(1229) <= layer3_outputs(3003);
    layer4_outputs(1230) <= not(layer3_outputs(1469));
    layer4_outputs(1231) <= not((layer3_outputs(1504)) and (layer3_outputs(1934)));
    layer4_outputs(1232) <= layer3_outputs(125);
    layer4_outputs(1233) <= '0';
    layer4_outputs(1234) <= not(layer3_outputs(6185));
    layer4_outputs(1235) <= (layer3_outputs(261)) xor (layer3_outputs(2697));
    layer4_outputs(1236) <= not((layer3_outputs(1854)) xor (layer3_outputs(6599)));
    layer4_outputs(1237) <= layer3_outputs(4666);
    layer4_outputs(1238) <= not(layer3_outputs(2472));
    layer4_outputs(1239) <= not(layer3_outputs(3990));
    layer4_outputs(1240) <= (layer3_outputs(2094)) or (layer3_outputs(5915));
    layer4_outputs(1241) <= not(layer3_outputs(6281));
    layer4_outputs(1242) <= layer3_outputs(2996);
    layer4_outputs(1243) <= not(layer3_outputs(878));
    layer4_outputs(1244) <= '1';
    layer4_outputs(1245) <= (layer3_outputs(6144)) or (layer3_outputs(594));
    layer4_outputs(1246) <= not((layer3_outputs(5433)) and (layer3_outputs(829)));
    layer4_outputs(1247) <= not(layer3_outputs(4031));
    layer4_outputs(1248) <= layer3_outputs(6337);
    layer4_outputs(1249) <= layer3_outputs(2711);
    layer4_outputs(1250) <= not(layer3_outputs(5458)) or (layer3_outputs(6041));
    layer4_outputs(1251) <= '1';
    layer4_outputs(1252) <= not((layer3_outputs(6563)) xor (layer3_outputs(2673)));
    layer4_outputs(1253) <= (layer3_outputs(7181)) and not (layer3_outputs(7457));
    layer4_outputs(1254) <= (layer3_outputs(5085)) and not (layer3_outputs(1349));
    layer4_outputs(1255) <= layer3_outputs(3171);
    layer4_outputs(1256) <= layer3_outputs(5335);
    layer4_outputs(1257) <= '1';
    layer4_outputs(1258) <= (layer3_outputs(1806)) and not (layer3_outputs(2435));
    layer4_outputs(1259) <= not(layer3_outputs(2864)) or (layer3_outputs(4369));
    layer4_outputs(1260) <= not((layer3_outputs(5830)) or (layer3_outputs(1779)));
    layer4_outputs(1261) <= '0';
    layer4_outputs(1262) <= (layer3_outputs(6303)) and (layer3_outputs(5469));
    layer4_outputs(1263) <= layer3_outputs(5949);
    layer4_outputs(1264) <= not(layer3_outputs(3434)) or (layer3_outputs(5409));
    layer4_outputs(1265) <= not(layer3_outputs(3301));
    layer4_outputs(1266) <= (layer3_outputs(5025)) and not (layer3_outputs(2973));
    layer4_outputs(1267) <= layer3_outputs(2640);
    layer4_outputs(1268) <= (layer3_outputs(4408)) and not (layer3_outputs(7643));
    layer4_outputs(1269) <= layer3_outputs(5414);
    layer4_outputs(1270) <= (layer3_outputs(6374)) xor (layer3_outputs(5885));
    layer4_outputs(1271) <= layer3_outputs(3996);
    layer4_outputs(1272) <= not(layer3_outputs(251));
    layer4_outputs(1273) <= not(layer3_outputs(1648));
    layer4_outputs(1274) <= not((layer3_outputs(3037)) or (layer3_outputs(3930)));
    layer4_outputs(1275) <= not((layer3_outputs(3719)) xor (layer3_outputs(312)));
    layer4_outputs(1276) <= not(layer3_outputs(7354));
    layer4_outputs(1277) <= (layer3_outputs(5051)) and (layer3_outputs(7435));
    layer4_outputs(1278) <= layer3_outputs(7266);
    layer4_outputs(1279) <= not(layer3_outputs(5516));
    layer4_outputs(1280) <= (layer3_outputs(629)) or (layer3_outputs(3719));
    layer4_outputs(1281) <= not(layer3_outputs(4879));
    layer4_outputs(1282) <= (layer3_outputs(6476)) or (layer3_outputs(5073));
    layer4_outputs(1283) <= layer3_outputs(1903);
    layer4_outputs(1284) <= not(layer3_outputs(4081));
    layer4_outputs(1285) <= (layer3_outputs(6170)) and not (layer3_outputs(4074));
    layer4_outputs(1286) <= not((layer3_outputs(3523)) and (layer3_outputs(4159)));
    layer4_outputs(1287) <= layer3_outputs(7196);
    layer4_outputs(1288) <= layer3_outputs(1584);
    layer4_outputs(1289) <= not(layer3_outputs(4375));
    layer4_outputs(1290) <= (layer3_outputs(1119)) xor (layer3_outputs(6373));
    layer4_outputs(1291) <= not(layer3_outputs(971)) or (layer3_outputs(3666));
    layer4_outputs(1292) <= layer3_outputs(3269);
    layer4_outputs(1293) <= layer3_outputs(7646);
    layer4_outputs(1294) <= (layer3_outputs(7082)) and not (layer3_outputs(1017));
    layer4_outputs(1295) <= not((layer3_outputs(5003)) or (layer3_outputs(5508)));
    layer4_outputs(1296) <= (layer3_outputs(2320)) or (layer3_outputs(6089));
    layer4_outputs(1297) <= not(layer3_outputs(3695)) or (layer3_outputs(575));
    layer4_outputs(1298) <= not(layer3_outputs(5706));
    layer4_outputs(1299) <= not(layer3_outputs(1205));
    layer4_outputs(1300) <= not(layer3_outputs(5701));
    layer4_outputs(1301) <= (layer3_outputs(7643)) and (layer3_outputs(1814));
    layer4_outputs(1302) <= layer3_outputs(244);
    layer4_outputs(1303) <= '0';
    layer4_outputs(1304) <= not(layer3_outputs(6033)) or (layer3_outputs(6562));
    layer4_outputs(1305) <= not((layer3_outputs(2454)) or (layer3_outputs(29)));
    layer4_outputs(1306) <= not((layer3_outputs(6921)) or (layer3_outputs(737)));
    layer4_outputs(1307) <= (layer3_outputs(473)) or (layer3_outputs(4769));
    layer4_outputs(1308) <= not((layer3_outputs(7432)) xor (layer3_outputs(5954)));
    layer4_outputs(1309) <= layer3_outputs(5796);
    layer4_outputs(1310) <= not(layer3_outputs(5497));
    layer4_outputs(1311) <= layer3_outputs(2210);
    layer4_outputs(1312) <= not(layer3_outputs(5519)) or (layer3_outputs(3497));
    layer4_outputs(1313) <= (layer3_outputs(4164)) and not (layer3_outputs(977));
    layer4_outputs(1314) <= not((layer3_outputs(4353)) and (layer3_outputs(3063)));
    layer4_outputs(1315) <= (layer3_outputs(4529)) xor (layer3_outputs(6767));
    layer4_outputs(1316) <= not((layer3_outputs(6429)) xor (layer3_outputs(2177)));
    layer4_outputs(1317) <= not(layer3_outputs(6044));
    layer4_outputs(1318) <= not(layer3_outputs(4619));
    layer4_outputs(1319) <= (layer3_outputs(1533)) xor (layer3_outputs(5482));
    layer4_outputs(1320) <= not(layer3_outputs(6468));
    layer4_outputs(1321) <= not(layer3_outputs(5249));
    layer4_outputs(1322) <= not(layer3_outputs(5803));
    layer4_outputs(1323) <= (layer3_outputs(5413)) or (layer3_outputs(3532));
    layer4_outputs(1324) <= not(layer3_outputs(3909));
    layer4_outputs(1325) <= not((layer3_outputs(582)) or (layer3_outputs(5477)));
    layer4_outputs(1326) <= (layer3_outputs(4990)) and (layer3_outputs(3823));
    layer4_outputs(1327) <= '1';
    layer4_outputs(1328) <= not(layer3_outputs(6928));
    layer4_outputs(1329) <= not(layer3_outputs(6116));
    layer4_outputs(1330) <= not((layer3_outputs(7377)) or (layer3_outputs(1744)));
    layer4_outputs(1331) <= not((layer3_outputs(3513)) xor (layer3_outputs(447)));
    layer4_outputs(1332) <= (layer3_outputs(2230)) and not (layer3_outputs(7189));
    layer4_outputs(1333) <= (layer3_outputs(2028)) or (layer3_outputs(1580));
    layer4_outputs(1334) <= not(layer3_outputs(7280));
    layer4_outputs(1335) <= not(layer3_outputs(2646));
    layer4_outputs(1336) <= layer3_outputs(4420);
    layer4_outputs(1337) <= layer3_outputs(4310);
    layer4_outputs(1338) <= not((layer3_outputs(1360)) and (layer3_outputs(3721)));
    layer4_outputs(1339) <= not((layer3_outputs(5402)) xor (layer3_outputs(7416)));
    layer4_outputs(1340) <= layer3_outputs(52);
    layer4_outputs(1341) <= layer3_outputs(5384);
    layer4_outputs(1342) <= (layer3_outputs(2485)) or (layer3_outputs(3054));
    layer4_outputs(1343) <= not(layer3_outputs(3461)) or (layer3_outputs(3565));
    layer4_outputs(1344) <= not((layer3_outputs(2087)) or (layer3_outputs(1615)));
    layer4_outputs(1345) <= (layer3_outputs(509)) or (layer3_outputs(4998));
    layer4_outputs(1346) <= layer3_outputs(359);
    layer4_outputs(1347) <= (layer3_outputs(3552)) and not (layer3_outputs(3118));
    layer4_outputs(1348) <= (layer3_outputs(3965)) or (layer3_outputs(2899));
    layer4_outputs(1349) <= layer3_outputs(6653);
    layer4_outputs(1350) <= not(layer3_outputs(7534));
    layer4_outputs(1351) <= (layer3_outputs(6330)) or (layer3_outputs(4881));
    layer4_outputs(1352) <= layer3_outputs(3012);
    layer4_outputs(1353) <= not(layer3_outputs(7583));
    layer4_outputs(1354) <= (layer3_outputs(7562)) and (layer3_outputs(6637));
    layer4_outputs(1355) <= not(layer3_outputs(7421));
    layer4_outputs(1356) <= not(layer3_outputs(783));
    layer4_outputs(1357) <= layer3_outputs(7600);
    layer4_outputs(1358) <= not(layer3_outputs(3418));
    layer4_outputs(1359) <= not(layer3_outputs(4456));
    layer4_outputs(1360) <= layer3_outputs(5719);
    layer4_outputs(1361) <= layer3_outputs(5200);
    layer4_outputs(1362) <= not((layer3_outputs(7327)) or (layer3_outputs(237)));
    layer4_outputs(1363) <= layer3_outputs(230);
    layer4_outputs(1364) <= not(layer3_outputs(4454)) or (layer3_outputs(2708));
    layer4_outputs(1365) <= layer3_outputs(2767);
    layer4_outputs(1366) <= layer3_outputs(1865);
    layer4_outputs(1367) <= not(layer3_outputs(5623));
    layer4_outputs(1368) <= (layer3_outputs(337)) or (layer3_outputs(793));
    layer4_outputs(1369) <= not((layer3_outputs(864)) xor (layer3_outputs(5684)));
    layer4_outputs(1370) <= not(layer3_outputs(3669));
    layer4_outputs(1371) <= not(layer3_outputs(6011));
    layer4_outputs(1372) <= layer3_outputs(4063);
    layer4_outputs(1373) <= layer3_outputs(3768);
    layer4_outputs(1374) <= not((layer3_outputs(3671)) or (layer3_outputs(2170)));
    layer4_outputs(1375) <= not(layer3_outputs(1013)) or (layer3_outputs(5491));
    layer4_outputs(1376) <= not((layer3_outputs(3470)) and (layer3_outputs(2338)));
    layer4_outputs(1377) <= not((layer3_outputs(126)) or (layer3_outputs(1306)));
    layer4_outputs(1378) <= (layer3_outputs(6747)) xor (layer3_outputs(391));
    layer4_outputs(1379) <= (layer3_outputs(54)) xor (layer3_outputs(2410));
    layer4_outputs(1380) <= not(layer3_outputs(6356));
    layer4_outputs(1381) <= not(layer3_outputs(1882));
    layer4_outputs(1382) <= not(layer3_outputs(236));
    layer4_outputs(1383) <= not(layer3_outputs(6527)) or (layer3_outputs(1296));
    layer4_outputs(1384) <= not(layer3_outputs(5689));
    layer4_outputs(1385) <= layer3_outputs(1352);
    layer4_outputs(1386) <= not((layer3_outputs(3972)) and (layer3_outputs(5290)));
    layer4_outputs(1387) <= not(layer3_outputs(6098)) or (layer3_outputs(4472));
    layer4_outputs(1388) <= not(layer3_outputs(4022));
    layer4_outputs(1389) <= (layer3_outputs(6680)) and not (layer3_outputs(2702));
    layer4_outputs(1390) <= layer3_outputs(4288);
    layer4_outputs(1391) <= not((layer3_outputs(6785)) xor (layer3_outputs(7157)));
    layer4_outputs(1392) <= (layer3_outputs(252)) and (layer3_outputs(1475));
    layer4_outputs(1393) <= not((layer3_outputs(1266)) xor (layer3_outputs(7444)));
    layer4_outputs(1394) <= not(layer3_outputs(6461)) or (layer3_outputs(1906));
    layer4_outputs(1395) <= not(layer3_outputs(18));
    layer4_outputs(1396) <= layer3_outputs(7530);
    layer4_outputs(1397) <= not((layer3_outputs(6874)) and (layer3_outputs(1572)));
    layer4_outputs(1398) <= not(layer3_outputs(2580));
    layer4_outputs(1399) <= not((layer3_outputs(2503)) and (layer3_outputs(980)));
    layer4_outputs(1400) <= not(layer3_outputs(3754)) or (layer3_outputs(4915));
    layer4_outputs(1401) <= not(layer3_outputs(795));
    layer4_outputs(1402) <= not((layer3_outputs(2132)) or (layer3_outputs(5717)));
    layer4_outputs(1403) <= not(layer3_outputs(1491));
    layer4_outputs(1404) <= (layer3_outputs(4204)) and not (layer3_outputs(3479));
    layer4_outputs(1405) <= not((layer3_outputs(4491)) and (layer3_outputs(1699)));
    layer4_outputs(1406) <= (layer3_outputs(1671)) and not (layer3_outputs(5898));
    layer4_outputs(1407) <= (layer3_outputs(2674)) and not (layer3_outputs(2120));
    layer4_outputs(1408) <= not(layer3_outputs(6745));
    layer4_outputs(1409) <= not(layer3_outputs(5151));
    layer4_outputs(1410) <= (layer3_outputs(1493)) and (layer3_outputs(1043));
    layer4_outputs(1411) <= layer3_outputs(7184);
    layer4_outputs(1412) <= (layer3_outputs(2152)) and (layer3_outputs(4708));
    layer4_outputs(1413) <= not(layer3_outputs(293));
    layer4_outputs(1414) <= not(layer3_outputs(3936));
    layer4_outputs(1415) <= layer3_outputs(3243);
    layer4_outputs(1416) <= not(layer3_outputs(2399));
    layer4_outputs(1417) <= not(layer3_outputs(6308));
    layer4_outputs(1418) <= not(layer3_outputs(738)) or (layer3_outputs(4702));
    layer4_outputs(1419) <= (layer3_outputs(4094)) and not (layer3_outputs(3888));
    layer4_outputs(1420) <= layer3_outputs(5451);
    layer4_outputs(1421) <= not((layer3_outputs(2505)) xor (layer3_outputs(2950)));
    layer4_outputs(1422) <= layer3_outputs(6611);
    layer4_outputs(1423) <= not(layer3_outputs(4660));
    layer4_outputs(1424) <= not((layer3_outputs(947)) and (layer3_outputs(898)));
    layer4_outputs(1425) <= not(layer3_outputs(3534));
    layer4_outputs(1426) <= '0';
    layer4_outputs(1427) <= layer3_outputs(1979);
    layer4_outputs(1428) <= (layer3_outputs(3563)) xor (layer3_outputs(1110));
    layer4_outputs(1429) <= (layer3_outputs(4796)) or (layer3_outputs(7542));
    layer4_outputs(1430) <= not((layer3_outputs(1898)) or (layer3_outputs(7083)));
    layer4_outputs(1431) <= not(layer3_outputs(4021));
    layer4_outputs(1432) <= (layer3_outputs(3398)) and not (layer3_outputs(1745));
    layer4_outputs(1433) <= not(layer3_outputs(6380));
    layer4_outputs(1434) <= (layer3_outputs(5873)) or (layer3_outputs(692));
    layer4_outputs(1435) <= not((layer3_outputs(5181)) and (layer3_outputs(594)));
    layer4_outputs(1436) <= not(layer3_outputs(6433));
    layer4_outputs(1437) <= layer3_outputs(7296);
    layer4_outputs(1438) <= (layer3_outputs(3279)) and not (layer3_outputs(833));
    layer4_outputs(1439) <= not((layer3_outputs(3684)) and (layer3_outputs(2675)));
    layer4_outputs(1440) <= not(layer3_outputs(2306));
    layer4_outputs(1441) <= layer3_outputs(2515);
    layer4_outputs(1442) <= not(layer3_outputs(4632));
    layer4_outputs(1443) <= not((layer3_outputs(6743)) and (layer3_outputs(1195)));
    layer4_outputs(1444) <= (layer3_outputs(349)) or (layer3_outputs(5766));
    layer4_outputs(1445) <= not(layer3_outputs(1497)) or (layer3_outputs(4218));
    layer4_outputs(1446) <= not(layer3_outputs(2631));
    layer4_outputs(1447) <= (layer3_outputs(5817)) and not (layer3_outputs(3946));
    layer4_outputs(1448) <= not(layer3_outputs(4168)) or (layer3_outputs(5704));
    layer4_outputs(1449) <= not((layer3_outputs(2981)) or (layer3_outputs(7625)));
    layer4_outputs(1450) <= not(layer3_outputs(7199));
    layer4_outputs(1451) <= not((layer3_outputs(2031)) and (layer3_outputs(4980)));
    layer4_outputs(1452) <= not((layer3_outputs(5674)) xor (layer3_outputs(5729)));
    layer4_outputs(1453) <= not(layer3_outputs(4394)) or (layer3_outputs(2345));
    layer4_outputs(1454) <= layer3_outputs(6019);
    layer4_outputs(1455) <= (layer3_outputs(1431)) and not (layer3_outputs(4490));
    layer4_outputs(1456) <= not(layer3_outputs(1149));
    layer4_outputs(1457) <= not((layer3_outputs(5364)) xor (layer3_outputs(5730)));
    layer4_outputs(1458) <= (layer3_outputs(1349)) or (layer3_outputs(2834));
    layer4_outputs(1459) <= not((layer3_outputs(3053)) or (layer3_outputs(4179)));
    layer4_outputs(1460) <= not((layer3_outputs(2443)) xor (layer3_outputs(6887)));
    layer4_outputs(1461) <= not(layer3_outputs(2747));
    layer4_outputs(1462) <= not((layer3_outputs(1834)) or (layer3_outputs(105)));
    layer4_outputs(1463) <= (layer3_outputs(2451)) and not (layer3_outputs(805));
    layer4_outputs(1464) <= (layer3_outputs(4860)) and not (layer3_outputs(6745));
    layer4_outputs(1465) <= not(layer3_outputs(1641)) or (layer3_outputs(28));
    layer4_outputs(1466) <= layer3_outputs(6081);
    layer4_outputs(1467) <= not(layer3_outputs(76)) or (layer3_outputs(115));
    layer4_outputs(1468) <= not(layer3_outputs(2745));
    layer4_outputs(1469) <= not(layer3_outputs(3781)) or (layer3_outputs(1231));
    layer4_outputs(1470) <= (layer3_outputs(6886)) or (layer3_outputs(868));
    layer4_outputs(1471) <= (layer3_outputs(394)) or (layer3_outputs(3508));
    layer4_outputs(1472) <= not((layer3_outputs(4602)) or (layer3_outputs(479)));
    layer4_outputs(1473) <= layer3_outputs(3882);
    layer4_outputs(1474) <= (layer3_outputs(1202)) or (layer3_outputs(2887));
    layer4_outputs(1475) <= (layer3_outputs(7116)) or (layer3_outputs(6761));
    layer4_outputs(1476) <= not(layer3_outputs(6471));
    layer4_outputs(1477) <= (layer3_outputs(1095)) or (layer3_outputs(2754));
    layer4_outputs(1478) <= not(layer3_outputs(2758));
    layer4_outputs(1479) <= not((layer3_outputs(4142)) and (layer3_outputs(6338)));
    layer4_outputs(1480) <= not(layer3_outputs(998));
    layer4_outputs(1481) <= not((layer3_outputs(1375)) or (layer3_outputs(1921)));
    layer4_outputs(1482) <= not(layer3_outputs(5865)) or (layer3_outputs(3325));
    layer4_outputs(1483) <= (layer3_outputs(6227)) xor (layer3_outputs(841));
    layer4_outputs(1484) <= (layer3_outputs(5187)) and not (layer3_outputs(7311));
    layer4_outputs(1485) <= not(layer3_outputs(5956)) or (layer3_outputs(7584));
    layer4_outputs(1486) <= not(layer3_outputs(1143));
    layer4_outputs(1487) <= (layer3_outputs(5402)) and not (layer3_outputs(2778));
    layer4_outputs(1488) <= not((layer3_outputs(6714)) and (layer3_outputs(3453)));
    layer4_outputs(1489) <= not((layer3_outputs(5322)) or (layer3_outputs(4126)));
    layer4_outputs(1490) <= (layer3_outputs(745)) and not (layer3_outputs(2870));
    layer4_outputs(1491) <= layer3_outputs(5259);
    layer4_outputs(1492) <= layer3_outputs(4049);
    layer4_outputs(1493) <= not((layer3_outputs(2363)) and (layer3_outputs(3305)));
    layer4_outputs(1494) <= layer3_outputs(7040);
    layer4_outputs(1495) <= not(layer3_outputs(5429));
    layer4_outputs(1496) <= layer3_outputs(5400);
    layer4_outputs(1497) <= layer3_outputs(2298);
    layer4_outputs(1498) <= (layer3_outputs(4030)) or (layer3_outputs(2220));
    layer4_outputs(1499) <= not((layer3_outputs(3760)) xor (layer3_outputs(2910)));
    layer4_outputs(1500) <= layer3_outputs(7499);
    layer4_outputs(1501) <= (layer3_outputs(6350)) or (layer3_outputs(7103));
    layer4_outputs(1502) <= '0';
    layer4_outputs(1503) <= (layer3_outputs(6097)) and not (layer3_outputs(1291));
    layer4_outputs(1504) <= not((layer3_outputs(5698)) or (layer3_outputs(2867)));
    layer4_outputs(1505) <= (layer3_outputs(664)) or (layer3_outputs(122));
    layer4_outputs(1506) <= (layer3_outputs(557)) and not (layer3_outputs(5710));
    layer4_outputs(1507) <= layer3_outputs(7510);
    layer4_outputs(1508) <= not(layer3_outputs(99));
    layer4_outputs(1509) <= (layer3_outputs(3917)) or (layer3_outputs(644));
    layer4_outputs(1510) <= not(layer3_outputs(703));
    layer4_outputs(1511) <= layer3_outputs(5767);
    layer4_outputs(1512) <= layer3_outputs(1980);
    layer4_outputs(1513) <= not((layer3_outputs(4689)) xor (layer3_outputs(2212)));
    layer4_outputs(1514) <= not(layer3_outputs(6234));
    layer4_outputs(1515) <= not(layer3_outputs(5320));
    layer4_outputs(1516) <= (layer3_outputs(4263)) and (layer3_outputs(6039));
    layer4_outputs(1517) <= (layer3_outputs(1881)) and not (layer3_outputs(7511));
    layer4_outputs(1518) <= not(layer3_outputs(3652)) or (layer3_outputs(3730));
    layer4_outputs(1519) <= not(layer3_outputs(2660));
    layer4_outputs(1520) <= layer3_outputs(965);
    layer4_outputs(1521) <= not(layer3_outputs(63));
    layer4_outputs(1522) <= not((layer3_outputs(4909)) or (layer3_outputs(3372)));
    layer4_outputs(1523) <= (layer3_outputs(2206)) and not (layer3_outputs(5872));
    layer4_outputs(1524) <= (layer3_outputs(1052)) or (layer3_outputs(4593));
    layer4_outputs(1525) <= not((layer3_outputs(2417)) xor (layer3_outputs(1535)));
    layer4_outputs(1526) <= not(layer3_outputs(7505));
    layer4_outputs(1527) <= not(layer3_outputs(830)) or (layer3_outputs(1530));
    layer4_outputs(1528) <= layer3_outputs(7180);
    layer4_outputs(1529) <= (layer3_outputs(6158)) or (layer3_outputs(3518));
    layer4_outputs(1530) <= (layer3_outputs(5408)) xor (layer3_outputs(7535));
    layer4_outputs(1531) <= (layer3_outputs(45)) and not (layer3_outputs(3596));
    layer4_outputs(1532) <= (layer3_outputs(516)) and not (layer3_outputs(4337));
    layer4_outputs(1533) <= not(layer3_outputs(7533));
    layer4_outputs(1534) <= not(layer3_outputs(4084));
    layer4_outputs(1535) <= (layer3_outputs(7255)) and not (layer3_outputs(870));
    layer4_outputs(1536) <= (layer3_outputs(4047)) and not (layer3_outputs(3146));
    layer4_outputs(1537) <= layer3_outputs(2536);
    layer4_outputs(1538) <= not((layer3_outputs(3186)) xor (layer3_outputs(5634)));
    layer4_outputs(1539) <= not((layer3_outputs(937)) xor (layer3_outputs(1628)));
    layer4_outputs(1540) <= (layer3_outputs(5091)) and not (layer3_outputs(673));
    layer4_outputs(1541) <= layer3_outputs(5309);
    layer4_outputs(1542) <= layer3_outputs(298);
    layer4_outputs(1543) <= not(layer3_outputs(5157));
    layer4_outputs(1544) <= layer3_outputs(1097);
    layer4_outputs(1545) <= layer3_outputs(4397);
    layer4_outputs(1546) <= not(layer3_outputs(7335));
    layer4_outputs(1547) <= not(layer3_outputs(322));
    layer4_outputs(1548) <= not(layer3_outputs(7102)) or (layer3_outputs(3510));
    layer4_outputs(1549) <= layer3_outputs(5465);
    layer4_outputs(1550) <= layer3_outputs(1813);
    layer4_outputs(1551) <= (layer3_outputs(5357)) or (layer3_outputs(1703));
    layer4_outputs(1552) <= not(layer3_outputs(3407));
    layer4_outputs(1553) <= not(layer3_outputs(340));
    layer4_outputs(1554) <= not(layer3_outputs(2555)) or (layer3_outputs(3317));
    layer4_outputs(1555) <= not(layer3_outputs(320));
    layer4_outputs(1556) <= (layer3_outputs(281)) and not (layer3_outputs(1491));
    layer4_outputs(1557) <= (layer3_outputs(1069)) or (layer3_outputs(6035));
    layer4_outputs(1558) <= layer3_outputs(4190);
    layer4_outputs(1559) <= '0';
    layer4_outputs(1560) <= (layer3_outputs(1834)) xor (layer3_outputs(3527));
    layer4_outputs(1561) <= (layer3_outputs(6987)) and (layer3_outputs(5630));
    layer4_outputs(1562) <= (layer3_outputs(6543)) and not (layer3_outputs(3160));
    layer4_outputs(1563) <= layer3_outputs(5197);
    layer4_outputs(1564) <= not(layer3_outputs(3950));
    layer4_outputs(1565) <= (layer3_outputs(6248)) and (layer3_outputs(2039));
    layer4_outputs(1566) <= (layer3_outputs(1301)) and not (layer3_outputs(4664));
    layer4_outputs(1567) <= not(layer3_outputs(6339));
    layer4_outputs(1568) <= layer3_outputs(1171);
    layer4_outputs(1569) <= not((layer3_outputs(7556)) or (layer3_outputs(4593)));
    layer4_outputs(1570) <= not(layer3_outputs(6835));
    layer4_outputs(1571) <= not(layer3_outputs(5174)) or (layer3_outputs(1453));
    layer4_outputs(1572) <= not(layer3_outputs(5223)) or (layer3_outputs(4317));
    layer4_outputs(1573) <= (layer3_outputs(1213)) and not (layer3_outputs(3846));
    layer4_outputs(1574) <= layer3_outputs(5693);
    layer4_outputs(1575) <= (layer3_outputs(2029)) and (layer3_outputs(3235));
    layer4_outputs(1576) <= (layer3_outputs(7573)) and (layer3_outputs(257));
    layer4_outputs(1577) <= layer3_outputs(416);
    layer4_outputs(1578) <= (layer3_outputs(6480)) and (layer3_outputs(248));
    layer4_outputs(1579) <= '0';
    layer4_outputs(1580) <= layer3_outputs(179);
    layer4_outputs(1581) <= not((layer3_outputs(886)) xor (layer3_outputs(115)));
    layer4_outputs(1582) <= not(layer3_outputs(5013)) or (layer3_outputs(7007));
    layer4_outputs(1583) <= (layer3_outputs(4148)) xor (layer3_outputs(4439));
    layer4_outputs(1584) <= not(layer3_outputs(6366)) or (layer3_outputs(2789));
    layer4_outputs(1585) <= not(layer3_outputs(5570));
    layer4_outputs(1586) <= (layer3_outputs(6340)) or (layer3_outputs(3024));
    layer4_outputs(1587) <= (layer3_outputs(3272)) and not (layer3_outputs(3392));
    layer4_outputs(1588) <= not(layer3_outputs(5942));
    layer4_outputs(1589) <= (layer3_outputs(2556)) and not (layer3_outputs(890));
    layer4_outputs(1590) <= not(layer3_outputs(4589));
    layer4_outputs(1591) <= not(layer3_outputs(1494));
    layer4_outputs(1592) <= (layer3_outputs(1083)) xor (layer3_outputs(3934));
    layer4_outputs(1593) <= (layer3_outputs(5813)) and not (layer3_outputs(4000));
    layer4_outputs(1594) <= not(layer3_outputs(1631));
    layer4_outputs(1595) <= not((layer3_outputs(4524)) or (layer3_outputs(6449)));
    layer4_outputs(1596) <= not(layer3_outputs(6792)) or (layer3_outputs(7291));
    layer4_outputs(1597) <= not((layer3_outputs(743)) xor (layer3_outputs(2467)));
    layer4_outputs(1598) <= not(layer3_outputs(3417));
    layer4_outputs(1599) <= layer3_outputs(6827);
    layer4_outputs(1600) <= layer3_outputs(4286);
    layer4_outputs(1601) <= not((layer3_outputs(7609)) xor (layer3_outputs(1024)));
    layer4_outputs(1602) <= (layer3_outputs(1558)) xor (layer3_outputs(4379));
    layer4_outputs(1603) <= not(layer3_outputs(5062));
    layer4_outputs(1604) <= not((layer3_outputs(1467)) and (layer3_outputs(6328)));
    layer4_outputs(1605) <= not(layer3_outputs(6994));
    layer4_outputs(1606) <= (layer3_outputs(104)) and not (layer3_outputs(1109));
    layer4_outputs(1607) <= not(layer3_outputs(5575));
    layer4_outputs(1608) <= layer3_outputs(703);
    layer4_outputs(1609) <= not((layer3_outputs(6412)) and (layer3_outputs(2285)));
    layer4_outputs(1610) <= not(layer3_outputs(5699)) or (layer3_outputs(3244));
    layer4_outputs(1611) <= layer3_outputs(465);
    layer4_outputs(1612) <= not((layer3_outputs(4064)) or (layer3_outputs(820)));
    layer4_outputs(1613) <= not((layer3_outputs(6722)) and (layer3_outputs(6504)));
    layer4_outputs(1614) <= (layer3_outputs(1363)) xor (layer3_outputs(5947));
    layer4_outputs(1615) <= layer3_outputs(7674);
    layer4_outputs(1616) <= not(layer3_outputs(7013));
    layer4_outputs(1617) <= (layer3_outputs(3650)) and not (layer3_outputs(4058));
    layer4_outputs(1618) <= (layer3_outputs(4243)) and not (layer3_outputs(3463));
    layer4_outputs(1619) <= not((layer3_outputs(6256)) xor (layer3_outputs(4668)));
    layer4_outputs(1620) <= not(layer3_outputs(1616));
    layer4_outputs(1621) <= (layer3_outputs(5199)) xor (layer3_outputs(2283));
    layer4_outputs(1622) <= layer3_outputs(234);
    layer4_outputs(1623) <= (layer3_outputs(1538)) and not (layer3_outputs(553));
    layer4_outputs(1624) <= (layer3_outputs(4247)) xor (layer3_outputs(3213));
    layer4_outputs(1625) <= not(layer3_outputs(4188));
    layer4_outputs(1626) <= not(layer3_outputs(6792));
    layer4_outputs(1627) <= layer3_outputs(702);
    layer4_outputs(1628) <= not(layer3_outputs(2034));
    layer4_outputs(1629) <= not((layer3_outputs(4112)) and (layer3_outputs(807)));
    layer4_outputs(1630) <= '1';
    layer4_outputs(1631) <= layer3_outputs(6262);
    layer4_outputs(1632) <= not(layer3_outputs(4567));
    layer4_outputs(1633) <= not(layer3_outputs(6517));
    layer4_outputs(1634) <= layer3_outputs(1083);
    layer4_outputs(1635) <= not(layer3_outputs(4819));
    layer4_outputs(1636) <= (layer3_outputs(5192)) or (layer3_outputs(3498));
    layer4_outputs(1637) <= layer3_outputs(335);
    layer4_outputs(1638) <= not(layer3_outputs(1598)) or (layer3_outputs(7026));
    layer4_outputs(1639) <= layer3_outputs(5399);
    layer4_outputs(1640) <= not((layer3_outputs(4073)) xor (layer3_outputs(6135)));
    layer4_outputs(1641) <= (layer3_outputs(2252)) xor (layer3_outputs(4358));
    layer4_outputs(1642) <= (layer3_outputs(1182)) and (layer3_outputs(1146));
    layer4_outputs(1643) <= not(layer3_outputs(1466));
    layer4_outputs(1644) <= not((layer3_outputs(4682)) and (layer3_outputs(836)));
    layer4_outputs(1645) <= '0';
    layer4_outputs(1646) <= (layer3_outputs(6815)) xor (layer3_outputs(3568));
    layer4_outputs(1647) <= layer3_outputs(6821);
    layer4_outputs(1648) <= (layer3_outputs(6420)) and not (layer3_outputs(4791));
    layer4_outputs(1649) <= (layer3_outputs(1796)) xor (layer3_outputs(3134));
    layer4_outputs(1650) <= not(layer3_outputs(1108));
    layer4_outputs(1651) <= not(layer3_outputs(4416)) or (layer3_outputs(716));
    layer4_outputs(1652) <= not(layer3_outputs(1188));
    layer4_outputs(1653) <= (layer3_outputs(4473)) and not (layer3_outputs(3692));
    layer4_outputs(1654) <= layer3_outputs(5907);
    layer4_outputs(1655) <= layer3_outputs(2452);
    layer4_outputs(1656) <= (layer3_outputs(6311)) or (layer3_outputs(6812));
    layer4_outputs(1657) <= not(layer3_outputs(483));
    layer4_outputs(1658) <= not(layer3_outputs(1005)) or (layer3_outputs(2501));
    layer4_outputs(1659) <= (layer3_outputs(399)) and (layer3_outputs(5846));
    layer4_outputs(1660) <= not(layer3_outputs(4302)) or (layer3_outputs(5901));
    layer4_outputs(1661) <= layer3_outputs(5774);
    layer4_outputs(1662) <= not(layer3_outputs(2779));
    layer4_outputs(1663) <= not(layer3_outputs(7543)) or (layer3_outputs(2667));
    layer4_outputs(1664) <= (layer3_outputs(5734)) and not (layer3_outputs(5930));
    layer4_outputs(1665) <= layer3_outputs(6963);
    layer4_outputs(1666) <= (layer3_outputs(4789)) and not (layer3_outputs(1842));
    layer4_outputs(1667) <= layer3_outputs(4882);
    layer4_outputs(1668) <= (layer3_outputs(7490)) and not (layer3_outputs(3254));
    layer4_outputs(1669) <= not(layer3_outputs(5153));
    layer4_outputs(1670) <= not(layer3_outputs(4728)) or (layer3_outputs(2979));
    layer4_outputs(1671) <= (layer3_outputs(7021)) and (layer3_outputs(6092));
    layer4_outputs(1672) <= layer3_outputs(7393);
    layer4_outputs(1673) <= not((layer3_outputs(3439)) or (layer3_outputs(3414)));
    layer4_outputs(1674) <= not(layer3_outputs(1403));
    layer4_outputs(1675) <= (layer3_outputs(1164)) or (layer3_outputs(2199));
    layer4_outputs(1676) <= (layer3_outputs(3187)) and not (layer3_outputs(2017));
    layer4_outputs(1677) <= not((layer3_outputs(5094)) and (layer3_outputs(765)));
    layer4_outputs(1678) <= (layer3_outputs(5824)) and (layer3_outputs(5010));
    layer4_outputs(1679) <= not(layer3_outputs(4849)) or (layer3_outputs(5496));
    layer4_outputs(1680) <= layer3_outputs(1485);
    layer4_outputs(1681) <= not(layer3_outputs(2710));
    layer4_outputs(1682) <= layer3_outputs(723);
    layer4_outputs(1683) <= (layer3_outputs(6713)) and (layer3_outputs(3379));
    layer4_outputs(1684) <= layer3_outputs(397);
    layer4_outputs(1685) <= not(layer3_outputs(7448));
    layer4_outputs(1686) <= layer3_outputs(3828);
    layer4_outputs(1687) <= not((layer3_outputs(474)) xor (layer3_outputs(6784)));
    layer4_outputs(1688) <= not(layer3_outputs(4446));
    layer4_outputs(1689) <= not((layer3_outputs(180)) and (layer3_outputs(861)));
    layer4_outputs(1690) <= not(layer3_outputs(1362)) or (layer3_outputs(5532));
    layer4_outputs(1691) <= (layer3_outputs(3168)) and not (layer3_outputs(3681));
    layer4_outputs(1692) <= (layer3_outputs(2908)) or (layer3_outputs(5916));
    layer4_outputs(1693) <= not(layer3_outputs(2065));
    layer4_outputs(1694) <= not(layer3_outputs(5989));
    layer4_outputs(1695) <= layer3_outputs(7675);
    layer4_outputs(1696) <= not(layer3_outputs(2994));
    layer4_outputs(1697) <= layer3_outputs(7149);
    layer4_outputs(1698) <= not(layer3_outputs(2934));
    layer4_outputs(1699) <= (layer3_outputs(5448)) and not (layer3_outputs(7237));
    layer4_outputs(1700) <= not(layer3_outputs(6306));
    layer4_outputs(1701) <= not(layer3_outputs(508));
    layer4_outputs(1702) <= layer3_outputs(955);
    layer4_outputs(1703) <= not(layer3_outputs(5893));
    layer4_outputs(1704) <= not(layer3_outputs(6192)) or (layer3_outputs(3595));
    layer4_outputs(1705) <= layer3_outputs(1963);
    layer4_outputs(1706) <= layer3_outputs(3351);
    layer4_outputs(1707) <= not(layer3_outputs(2915)) or (layer3_outputs(5251));
    layer4_outputs(1708) <= not(layer3_outputs(3286));
    layer4_outputs(1709) <= layer3_outputs(7036);
    layer4_outputs(1710) <= layer3_outputs(3576);
    layer4_outputs(1711) <= not(layer3_outputs(2562));
    layer4_outputs(1712) <= (layer3_outputs(2219)) and not (layer3_outputs(5538));
    layer4_outputs(1713) <= not(layer3_outputs(851));
    layer4_outputs(1714) <= not((layer3_outputs(3137)) xor (layer3_outputs(2205)));
    layer4_outputs(1715) <= not(layer3_outputs(7499));
    layer4_outputs(1716) <= not(layer3_outputs(6296));
    layer4_outputs(1717) <= (layer3_outputs(5048)) or (layer3_outputs(5074));
    layer4_outputs(1718) <= not(layer3_outputs(286));
    layer4_outputs(1719) <= not((layer3_outputs(5045)) or (layer3_outputs(5555)));
    layer4_outputs(1720) <= layer3_outputs(6385);
    layer4_outputs(1721) <= (layer3_outputs(4229)) and not (layer3_outputs(1711));
    layer4_outputs(1722) <= not(layer3_outputs(2381));
    layer4_outputs(1723) <= not((layer3_outputs(7656)) or (layer3_outputs(3554)));
    layer4_outputs(1724) <= (layer3_outputs(7430)) and not (layer3_outputs(7677));
    layer4_outputs(1725) <= not((layer3_outputs(4647)) and (layer3_outputs(150)));
    layer4_outputs(1726) <= not(layer3_outputs(3128));
    layer4_outputs(1727) <= not((layer3_outputs(3191)) and (layer3_outputs(5655)));
    layer4_outputs(1728) <= (layer3_outputs(158)) and not (layer3_outputs(6130));
    layer4_outputs(1729) <= not((layer3_outputs(1226)) or (layer3_outputs(4308)));
    layer4_outputs(1730) <= '0';
    layer4_outputs(1731) <= not((layer3_outputs(1380)) or (layer3_outputs(5106)));
    layer4_outputs(1732) <= not(layer3_outputs(6442));
    layer4_outputs(1733) <= layer3_outputs(600);
    layer4_outputs(1734) <= (layer3_outputs(2337)) and not (layer3_outputs(5538));
    layer4_outputs(1735) <= (layer3_outputs(62)) or (layer3_outputs(5211));
    layer4_outputs(1736) <= not((layer3_outputs(5819)) or (layer3_outputs(1632)));
    layer4_outputs(1737) <= not((layer3_outputs(6659)) xor (layer3_outputs(2225)));
    layer4_outputs(1738) <= not(layer3_outputs(4239));
    layer4_outputs(1739) <= not((layer3_outputs(1976)) xor (layer3_outputs(6492)));
    layer4_outputs(1740) <= not(layer3_outputs(2762));
    layer4_outputs(1741) <= not(layer3_outputs(1768)) or (layer3_outputs(883));
    layer4_outputs(1742) <= (layer3_outputs(2977)) and not (layer3_outputs(3428));
    layer4_outputs(1743) <= (layer3_outputs(592)) or (layer3_outputs(3819));
    layer4_outputs(1744) <= not(layer3_outputs(7436));
    layer4_outputs(1745) <= not(layer3_outputs(7329));
    layer4_outputs(1746) <= '1';
    layer4_outputs(1747) <= (layer3_outputs(4989)) and not (layer3_outputs(6118));
    layer4_outputs(1748) <= layer3_outputs(5216);
    layer4_outputs(1749) <= not(layer3_outputs(3626));
    layer4_outputs(1750) <= not(layer3_outputs(583));
    layer4_outputs(1751) <= not(layer3_outputs(2793));
    layer4_outputs(1752) <= layer3_outputs(6435);
    layer4_outputs(1753) <= '1';
    layer4_outputs(1754) <= '0';
    layer4_outputs(1755) <= not(layer3_outputs(5887));
    layer4_outputs(1756) <= not(layer3_outputs(597)) or (layer3_outputs(4116));
    layer4_outputs(1757) <= not(layer3_outputs(1455));
    layer4_outputs(1758) <= (layer3_outputs(968)) and not (layer3_outputs(822));
    layer4_outputs(1759) <= (layer3_outputs(203)) and not (layer3_outputs(731));
    layer4_outputs(1760) <= not(layer3_outputs(3359));
    layer4_outputs(1761) <= not(layer3_outputs(3923));
    layer4_outputs(1762) <= not(layer3_outputs(5081));
    layer4_outputs(1763) <= not(layer3_outputs(828));
    layer4_outputs(1764) <= not((layer3_outputs(2374)) and (layer3_outputs(1984)));
    layer4_outputs(1765) <= not(layer3_outputs(3794)) or (layer3_outputs(4705));
    layer4_outputs(1766) <= layer3_outputs(2960);
    layer4_outputs(1767) <= not((layer3_outputs(77)) xor (layer3_outputs(7426)));
    layer4_outputs(1768) <= layer3_outputs(5304);
    layer4_outputs(1769) <= (layer3_outputs(5263)) and not (layer3_outputs(6055));
    layer4_outputs(1770) <= not(layer3_outputs(7101)) or (layer3_outputs(6301));
    layer4_outputs(1771) <= layer3_outputs(6291);
    layer4_outputs(1772) <= not((layer3_outputs(728)) or (layer3_outputs(508)));
    layer4_outputs(1773) <= (layer3_outputs(1505)) xor (layer3_outputs(3713));
    layer4_outputs(1774) <= layer3_outputs(3346);
    layer4_outputs(1775) <= layer3_outputs(1618);
    layer4_outputs(1776) <= (layer3_outputs(1134)) or (layer3_outputs(7631));
    layer4_outputs(1777) <= not(layer3_outputs(4374));
    layer4_outputs(1778) <= not(layer3_outputs(3694));
    layer4_outputs(1779) <= not(layer3_outputs(6975));
    layer4_outputs(1780) <= (layer3_outputs(4226)) and not (layer3_outputs(5203));
    layer4_outputs(1781) <= layer3_outputs(3225);
    layer4_outputs(1782) <= not(layer3_outputs(5498)) or (layer3_outputs(1283));
    layer4_outputs(1783) <= not(layer3_outputs(387));
    layer4_outputs(1784) <= not(layer3_outputs(7505));
    layer4_outputs(1785) <= not(layer3_outputs(6081));
    layer4_outputs(1786) <= '0';
    layer4_outputs(1787) <= (layer3_outputs(7052)) and not (layer3_outputs(2376));
    layer4_outputs(1788) <= not(layer3_outputs(7472));
    layer4_outputs(1789) <= layer3_outputs(3845);
    layer4_outputs(1790) <= not(layer3_outputs(6017));
    layer4_outputs(1791) <= not(layer3_outputs(7253));
    layer4_outputs(1792) <= layer3_outputs(1342);
    layer4_outputs(1793) <= not(layer3_outputs(3460)) or (layer3_outputs(3848));
    layer4_outputs(1794) <= not(layer3_outputs(4778));
    layer4_outputs(1795) <= layer3_outputs(2559);
    layer4_outputs(1796) <= not(layer3_outputs(7331));
    layer4_outputs(1797) <= not(layer3_outputs(3597));
    layer4_outputs(1798) <= layer3_outputs(7062);
    layer4_outputs(1799) <= layer3_outputs(6693);
    layer4_outputs(1800) <= layer3_outputs(6095);
    layer4_outputs(1801) <= '0';
    layer4_outputs(1802) <= not(layer3_outputs(5480));
    layer4_outputs(1803) <= layer3_outputs(7339);
    layer4_outputs(1804) <= (layer3_outputs(6346)) or (layer3_outputs(683));
    layer4_outputs(1805) <= layer3_outputs(2093);
    layer4_outputs(1806) <= (layer3_outputs(2124)) or (layer3_outputs(1931));
    layer4_outputs(1807) <= layer3_outputs(2394);
    layer4_outputs(1808) <= not(layer3_outputs(965)) or (layer3_outputs(2560));
    layer4_outputs(1809) <= not(layer3_outputs(5319));
    layer4_outputs(1810) <= not(layer3_outputs(5361));
    layer4_outputs(1811) <= (layer3_outputs(3727)) or (layer3_outputs(3825));
    layer4_outputs(1812) <= (layer3_outputs(2464)) and not (layer3_outputs(7478));
    layer4_outputs(1813) <= not((layer3_outputs(5125)) or (layer3_outputs(527)));
    layer4_outputs(1814) <= not(layer3_outputs(4346));
    layer4_outputs(1815) <= (layer3_outputs(5077)) and (layer3_outputs(6062));
    layer4_outputs(1816) <= layer3_outputs(1635);
    layer4_outputs(1817) <= not((layer3_outputs(2764)) or (layer3_outputs(3931)));
    layer4_outputs(1818) <= layer3_outputs(4680);
    layer4_outputs(1819) <= (layer3_outputs(57)) xor (layer3_outputs(2705));
    layer4_outputs(1820) <= not(layer3_outputs(94));
    layer4_outputs(1821) <= not((layer3_outputs(7639)) and (layer3_outputs(69)));
    layer4_outputs(1822) <= not((layer3_outputs(5343)) or (layer3_outputs(1357)));
    layer4_outputs(1823) <= not(layer3_outputs(1327));
    layer4_outputs(1824) <= not(layer3_outputs(6949));
    layer4_outputs(1825) <= not((layer3_outputs(6903)) or (layer3_outputs(5950)));
    layer4_outputs(1826) <= (layer3_outputs(2778)) or (layer3_outputs(4421));
    layer4_outputs(1827) <= (layer3_outputs(2325)) xor (layer3_outputs(6419));
    layer4_outputs(1828) <= not(layer3_outputs(4212));
    layer4_outputs(1829) <= (layer3_outputs(4812)) or (layer3_outputs(2059));
    layer4_outputs(1830) <= layer3_outputs(5807);
    layer4_outputs(1831) <= layer3_outputs(1326);
    layer4_outputs(1832) <= layer3_outputs(1018);
    layer4_outputs(1833) <= not(layer3_outputs(3814));
    layer4_outputs(1834) <= not(layer3_outputs(1732));
    layer4_outputs(1835) <= (layer3_outputs(7427)) and not (layer3_outputs(270));
    layer4_outputs(1836) <= layer3_outputs(2818);
    layer4_outputs(1837) <= layer3_outputs(1939);
    layer4_outputs(1838) <= not((layer3_outputs(4850)) xor (layer3_outputs(4137)));
    layer4_outputs(1839) <= layer3_outputs(2913);
    layer4_outputs(1840) <= '0';
    layer4_outputs(1841) <= layer3_outputs(5759);
    layer4_outputs(1842) <= not((layer3_outputs(480)) and (layer3_outputs(2532)));
    layer4_outputs(1843) <= layer3_outputs(6475);
    layer4_outputs(1844) <= not((layer3_outputs(1793)) xor (layer3_outputs(7560)));
    layer4_outputs(1845) <= (layer3_outputs(5500)) and not (layer3_outputs(7101));
    layer4_outputs(1846) <= not(layer3_outputs(5962));
    layer4_outputs(1847) <= layer3_outputs(586);
    layer4_outputs(1848) <= not(layer3_outputs(421));
    layer4_outputs(1849) <= layer3_outputs(4360);
    layer4_outputs(1850) <= layer3_outputs(3354);
    layer4_outputs(1851) <= not((layer3_outputs(4038)) xor (layer3_outputs(5069)));
    layer4_outputs(1852) <= layer3_outputs(5299);
    layer4_outputs(1853) <= '1';
    layer4_outputs(1854) <= layer3_outputs(4026);
    layer4_outputs(1855) <= layer3_outputs(6319);
    layer4_outputs(1856) <= layer3_outputs(6912);
    layer4_outputs(1857) <= (layer3_outputs(4559)) and (layer3_outputs(284));
    layer4_outputs(1858) <= not(layer3_outputs(6477)) or (layer3_outputs(6502));
    layer4_outputs(1859) <= (layer3_outputs(6100)) and (layer3_outputs(5439));
    layer4_outputs(1860) <= not(layer3_outputs(3596));
    layer4_outputs(1861) <= not(layer3_outputs(7377)) or (layer3_outputs(449));
    layer4_outputs(1862) <= layer3_outputs(537);
    layer4_outputs(1863) <= (layer3_outputs(5083)) or (layer3_outputs(1069));
    layer4_outputs(1864) <= layer3_outputs(2469);
    layer4_outputs(1865) <= not(layer3_outputs(3266));
    layer4_outputs(1866) <= (layer3_outputs(5931)) and (layer3_outputs(4906));
    layer4_outputs(1867) <= (layer3_outputs(2175)) and not (layer3_outputs(2484));
    layer4_outputs(1868) <= (layer3_outputs(2782)) xor (layer3_outputs(6201));
    layer4_outputs(1869) <= not(layer3_outputs(6574)) or (layer3_outputs(4453));
    layer4_outputs(1870) <= not(layer3_outputs(404));
    layer4_outputs(1871) <= not(layer3_outputs(451));
    layer4_outputs(1872) <= (layer3_outputs(2357)) or (layer3_outputs(1449));
    layer4_outputs(1873) <= (layer3_outputs(76)) and not (layer3_outputs(5509));
    layer4_outputs(1874) <= not((layer3_outputs(5671)) xor (layer3_outputs(396)));
    layer4_outputs(1875) <= not(layer3_outputs(1533));
    layer4_outputs(1876) <= layer3_outputs(612);
    layer4_outputs(1877) <= layer3_outputs(2170);
    layer4_outputs(1878) <= not(layer3_outputs(7054));
    layer4_outputs(1879) <= layer3_outputs(7070);
    layer4_outputs(1880) <= (layer3_outputs(4121)) xor (layer3_outputs(6278));
    layer4_outputs(1881) <= layer3_outputs(4296);
    layer4_outputs(1882) <= layer3_outputs(1381);
    layer4_outputs(1883) <= not((layer3_outputs(6555)) and (layer3_outputs(3438)));
    layer4_outputs(1884) <= (layer3_outputs(3780)) and not (layer3_outputs(2265));
    layer4_outputs(1885) <= (layer3_outputs(1791)) or (layer3_outputs(3029));
    layer4_outputs(1886) <= layer3_outputs(6716);
    layer4_outputs(1887) <= not(layer3_outputs(3339));
    layer4_outputs(1888) <= (layer3_outputs(5072)) and not (layer3_outputs(5029));
    layer4_outputs(1889) <= not(layer3_outputs(3958));
    layer4_outputs(1890) <= not(layer3_outputs(3939)) or (layer3_outputs(3909));
    layer4_outputs(1891) <= (layer3_outputs(4193)) or (layer3_outputs(860));
    layer4_outputs(1892) <= (layer3_outputs(1688)) and (layer3_outputs(724));
    layer4_outputs(1893) <= not((layer3_outputs(1896)) xor (layer3_outputs(4686)));
    layer4_outputs(1894) <= not(layer3_outputs(6963));
    layer4_outputs(1895) <= layer3_outputs(161);
    layer4_outputs(1896) <= not((layer3_outputs(6676)) xor (layer3_outputs(4451)));
    layer4_outputs(1897) <= layer3_outputs(3151);
    layer4_outputs(1898) <= not((layer3_outputs(6194)) or (layer3_outputs(4685)));
    layer4_outputs(1899) <= not(layer3_outputs(2957)) or (layer3_outputs(7632));
    layer4_outputs(1900) <= layer3_outputs(1246);
    layer4_outputs(1901) <= not(layer3_outputs(699)) or (layer3_outputs(5186));
    layer4_outputs(1902) <= layer3_outputs(1692);
    layer4_outputs(1903) <= not((layer3_outputs(2272)) xor (layer3_outputs(1461)));
    layer4_outputs(1904) <= not(layer3_outputs(4826));
    layer4_outputs(1905) <= layer3_outputs(300);
    layer4_outputs(1906) <= layer3_outputs(1712);
    layer4_outputs(1907) <= not(layer3_outputs(5647)) or (layer3_outputs(2698));
    layer4_outputs(1908) <= not((layer3_outputs(4399)) and (layer3_outputs(7260)));
    layer4_outputs(1909) <= layer3_outputs(3963);
    layer4_outputs(1910) <= (layer3_outputs(171)) and (layer3_outputs(2666));
    layer4_outputs(1911) <= '1';
    layer4_outputs(1912) <= layer3_outputs(3873);
    layer4_outputs(1913) <= not((layer3_outputs(3331)) and (layer3_outputs(1828)));
    layer4_outputs(1914) <= (layer3_outputs(6335)) and not (layer3_outputs(6880));
    layer4_outputs(1915) <= not(layer3_outputs(1135));
    layer4_outputs(1916) <= layer3_outputs(4481);
    layer4_outputs(1917) <= (layer3_outputs(3129)) and not (layer3_outputs(7296));
    layer4_outputs(1918) <= not((layer3_outputs(3345)) and (layer3_outputs(1603)));
    layer4_outputs(1919) <= not(layer3_outputs(5452));
    layer4_outputs(1920) <= layer3_outputs(823);
    layer4_outputs(1921) <= not((layer3_outputs(4234)) and (layer3_outputs(4927)));
    layer4_outputs(1922) <= not(layer3_outputs(1169));
    layer4_outputs(1923) <= not((layer3_outputs(7060)) xor (layer3_outputs(5860)));
    layer4_outputs(1924) <= not(layer3_outputs(7113));
    layer4_outputs(1925) <= layer3_outputs(760);
    layer4_outputs(1926) <= not(layer3_outputs(4830)) or (layer3_outputs(6865));
    layer4_outputs(1927) <= (layer3_outputs(6666)) and not (layer3_outputs(3799));
    layer4_outputs(1928) <= layer3_outputs(7396);
    layer4_outputs(1929) <= (layer3_outputs(5953)) and not (layer3_outputs(7294));
    layer4_outputs(1930) <= not(layer3_outputs(3635));
    layer4_outputs(1931) <= layer3_outputs(4969);
    layer4_outputs(1932) <= not((layer3_outputs(5555)) xor (layer3_outputs(4983)));
    layer4_outputs(1933) <= not(layer3_outputs(4307)) or (layer3_outputs(2866));
    layer4_outputs(1934) <= not(layer3_outputs(7581));
    layer4_outputs(1935) <= not((layer3_outputs(3332)) xor (layer3_outputs(5918)));
    layer4_outputs(1936) <= not(layer3_outputs(4782)) or (layer3_outputs(3161));
    layer4_outputs(1937) <= (layer3_outputs(1336)) and not (layer3_outputs(6269));
    layer4_outputs(1938) <= layer3_outputs(4327);
    layer4_outputs(1939) <= not(layer3_outputs(1524));
    layer4_outputs(1940) <= not(layer3_outputs(6683));
    layer4_outputs(1941) <= not(layer3_outputs(5566)) or (layer3_outputs(1865));
    layer4_outputs(1942) <= (layer3_outputs(5049)) and not (layer3_outputs(1872));
    layer4_outputs(1943) <= not(layer3_outputs(2330)) or (layer3_outputs(4658));
    layer4_outputs(1944) <= (layer3_outputs(528)) and not (layer3_outputs(656));
    layer4_outputs(1945) <= layer3_outputs(332);
    layer4_outputs(1946) <= not((layer3_outputs(2179)) or (layer3_outputs(7488)));
    layer4_outputs(1947) <= not((layer3_outputs(1114)) or (layer3_outputs(1780)));
    layer4_outputs(1948) <= (layer3_outputs(430)) xor (layer3_outputs(4472));
    layer4_outputs(1949) <= layer3_outputs(7605);
    layer4_outputs(1950) <= not((layer3_outputs(4440)) and (layer3_outputs(5897)));
    layer4_outputs(1951) <= not(layer3_outputs(1816));
    layer4_outputs(1952) <= layer3_outputs(2818);
    layer4_outputs(1953) <= layer3_outputs(4505);
    layer4_outputs(1954) <= (layer3_outputs(3982)) and not (layer3_outputs(3144));
    layer4_outputs(1955) <= (layer3_outputs(2460)) or (layer3_outputs(536));
    layer4_outputs(1956) <= not((layer3_outputs(7333)) and (layer3_outputs(3050)));
    layer4_outputs(1957) <= layer3_outputs(2676);
    layer4_outputs(1958) <= not(layer3_outputs(2542));
    layer4_outputs(1959) <= not(layer3_outputs(2394));
    layer4_outputs(1960) <= (layer3_outputs(5903)) or (layer3_outputs(2616));
    layer4_outputs(1961) <= not(layer3_outputs(1408));
    layer4_outputs(1962) <= layer3_outputs(4349);
    layer4_outputs(1963) <= (layer3_outputs(1290)) and (layer3_outputs(2909));
    layer4_outputs(1964) <= layer3_outputs(378);
    layer4_outputs(1965) <= not(layer3_outputs(2378));
    layer4_outputs(1966) <= layer3_outputs(6398);
    layer4_outputs(1967) <= not(layer3_outputs(3806));
    layer4_outputs(1968) <= layer3_outputs(349);
    layer4_outputs(1969) <= (layer3_outputs(2667)) or (layer3_outputs(5372));
    layer4_outputs(1970) <= not((layer3_outputs(4803)) or (layer3_outputs(3327)));
    layer4_outputs(1971) <= not(layer3_outputs(1960));
    layer4_outputs(1972) <= not(layer3_outputs(1306));
    layer4_outputs(1973) <= not((layer3_outputs(3369)) or (layer3_outputs(4250)));
    layer4_outputs(1974) <= not(layer3_outputs(5847));
    layer4_outputs(1975) <= not(layer3_outputs(6561));
    layer4_outputs(1976) <= layer3_outputs(5665);
    layer4_outputs(1977) <= layer3_outputs(3704);
    layer4_outputs(1978) <= not(layer3_outputs(5870)) or (layer3_outputs(7068));
    layer4_outputs(1979) <= layer3_outputs(1434);
    layer4_outputs(1980) <= layer3_outputs(1002);
    layer4_outputs(1981) <= layer3_outputs(4129);
    layer4_outputs(1982) <= layer3_outputs(2151);
    layer4_outputs(1983) <= layer3_outputs(4233);
    layer4_outputs(1984) <= (layer3_outputs(1289)) or (layer3_outputs(532));
    layer4_outputs(1985) <= (layer3_outputs(222)) and (layer3_outputs(3838));
    layer4_outputs(1986) <= (layer3_outputs(4786)) and (layer3_outputs(4907));
    layer4_outputs(1987) <= layer3_outputs(5207);
    layer4_outputs(1988) <= layer3_outputs(1074);
    layer4_outputs(1989) <= layer3_outputs(3001);
    layer4_outputs(1990) <= not(layer3_outputs(4105));
    layer4_outputs(1991) <= (layer3_outputs(2560)) and not (layer3_outputs(5477));
    layer4_outputs(1992) <= layer3_outputs(4888);
    layer4_outputs(1993) <= not(layer3_outputs(3838)) or (layer3_outputs(1041));
    layer4_outputs(1994) <= (layer3_outputs(6540)) and (layer3_outputs(4519));
    layer4_outputs(1995) <= not(layer3_outputs(4200)) or (layer3_outputs(5664));
    layer4_outputs(1996) <= (layer3_outputs(7539)) or (layer3_outputs(139));
    layer4_outputs(1997) <= not(layer3_outputs(148));
    layer4_outputs(1998) <= not(layer3_outputs(203)) or (layer3_outputs(5920));
    layer4_outputs(1999) <= not(layer3_outputs(5197));
    layer4_outputs(2000) <= layer3_outputs(7294);
    layer4_outputs(2001) <= not(layer3_outputs(5793));
    layer4_outputs(2002) <= layer3_outputs(3804);
    layer4_outputs(2003) <= '0';
    layer4_outputs(2004) <= layer3_outputs(3162);
    layer4_outputs(2005) <= layer3_outputs(6203);
    layer4_outputs(2006) <= layer3_outputs(5631);
    layer4_outputs(2007) <= (layer3_outputs(5288)) or (layer3_outputs(2232));
    layer4_outputs(2008) <= not(layer3_outputs(2422));
    layer4_outputs(2009) <= (layer3_outputs(2841)) or (layer3_outputs(7651));
    layer4_outputs(2010) <= not(layer3_outputs(2175));
    layer4_outputs(2011) <= layer3_outputs(4626);
    layer4_outputs(2012) <= (layer3_outputs(4921)) or (layer3_outputs(4522));
    layer4_outputs(2013) <= '1';
    layer4_outputs(2014) <= not(layer3_outputs(1354));
    layer4_outputs(2015) <= layer3_outputs(6844);
    layer4_outputs(2016) <= not(layer3_outputs(3598));
    layer4_outputs(2017) <= (layer3_outputs(6503)) and not (layer3_outputs(6901));
    layer4_outputs(2018) <= (layer3_outputs(796)) and not (layer3_outputs(3969));
    layer4_outputs(2019) <= not((layer3_outputs(325)) or (layer3_outputs(68)));
    layer4_outputs(2020) <= (layer3_outputs(1765)) xor (layer3_outputs(6031));
    layer4_outputs(2021) <= not(layer3_outputs(178));
    layer4_outputs(2022) <= layer3_outputs(2025);
    layer4_outputs(2023) <= not(layer3_outputs(457));
    layer4_outputs(2024) <= (layer3_outputs(1046)) and not (layer3_outputs(7488));
    layer4_outputs(2025) <= not((layer3_outputs(355)) or (layer3_outputs(7072)));
    layer4_outputs(2026) <= (layer3_outputs(5391)) and (layer3_outputs(6771));
    layer4_outputs(2027) <= not(layer3_outputs(1868)) or (layer3_outputs(4700));
    layer4_outputs(2028) <= not(layer3_outputs(5096));
    layer4_outputs(2029) <= (layer3_outputs(2116)) xor (layer3_outputs(2520));
    layer4_outputs(2030) <= (layer3_outputs(4187)) or (layer3_outputs(5690));
    layer4_outputs(2031) <= (layer3_outputs(7203)) and (layer3_outputs(6156));
    layer4_outputs(2032) <= (layer3_outputs(761)) and not (layer3_outputs(162));
    layer4_outputs(2033) <= not(layer3_outputs(93)) or (layer3_outputs(7679));
    layer4_outputs(2034) <= layer3_outputs(3568);
    layer4_outputs(2035) <= (layer3_outputs(720)) and (layer3_outputs(5289));
    layer4_outputs(2036) <= not((layer3_outputs(1341)) xor (layer3_outputs(2209)));
    layer4_outputs(2037) <= not(layer3_outputs(625));
    layer4_outputs(2038) <= layer3_outputs(4663);
    layer4_outputs(2039) <= not((layer3_outputs(46)) or (layer3_outputs(633)));
    layer4_outputs(2040) <= not((layer3_outputs(5866)) xor (layer3_outputs(4544)));
    layer4_outputs(2041) <= not(layer3_outputs(563));
    layer4_outputs(2042) <= not(layer3_outputs(4066));
    layer4_outputs(2043) <= layer3_outputs(7317);
    layer4_outputs(2044) <= not(layer3_outputs(4793));
    layer4_outputs(2045) <= layer3_outputs(6650);
    layer4_outputs(2046) <= layer3_outputs(6950);
    layer4_outputs(2047) <= layer3_outputs(3858);
    layer4_outputs(2048) <= (layer3_outputs(6971)) and not (layer3_outputs(4824));
    layer4_outputs(2049) <= not(layer3_outputs(5608));
    layer4_outputs(2050) <= (layer3_outputs(5256)) and (layer3_outputs(3734));
    layer4_outputs(2051) <= layer3_outputs(5733);
    layer4_outputs(2052) <= (layer3_outputs(4309)) and (layer3_outputs(1922));
    layer4_outputs(2053) <= not(layer3_outputs(4223)) or (layer3_outputs(5929));
    layer4_outputs(2054) <= not(layer3_outputs(7433));
    layer4_outputs(2055) <= not((layer3_outputs(7591)) or (layer3_outputs(3716)));
    layer4_outputs(2056) <= layer3_outputs(2881);
    layer4_outputs(2057) <= '0';
    layer4_outputs(2058) <= not(layer3_outputs(5968));
    layer4_outputs(2059) <= not((layer3_outputs(5633)) and (layer3_outputs(3580)));
    layer4_outputs(2060) <= layer3_outputs(1578);
    layer4_outputs(2061) <= layer3_outputs(3572);
    layer4_outputs(2062) <= not((layer3_outputs(3049)) or (layer3_outputs(1787)));
    layer4_outputs(2063) <= not(layer3_outputs(3449));
    layer4_outputs(2064) <= not(layer3_outputs(1318)) or (layer3_outputs(3455));
    layer4_outputs(2065) <= not(layer3_outputs(591));
    layer4_outputs(2066) <= not((layer3_outputs(1984)) and (layer3_outputs(2726)));
    layer4_outputs(2067) <= layer3_outputs(1307);
    layer4_outputs(2068) <= layer3_outputs(1284);
    layer4_outputs(2069) <= layer3_outputs(2473);
    layer4_outputs(2070) <= not(layer3_outputs(3444));
    layer4_outputs(2071) <= not(layer3_outputs(1963));
    layer4_outputs(2072) <= layer3_outputs(2120);
    layer4_outputs(2073) <= layer3_outputs(7324);
    layer4_outputs(2074) <= (layer3_outputs(273)) xor (layer3_outputs(3121));
    layer4_outputs(2075) <= layer3_outputs(6828);
    layer4_outputs(2076) <= (layer3_outputs(4418)) and not (layer3_outputs(3141));
    layer4_outputs(2077) <= layer3_outputs(4095);
    layer4_outputs(2078) <= (layer3_outputs(3217)) and (layer3_outputs(4199));
    layer4_outputs(2079) <= '0';
    layer4_outputs(2080) <= layer3_outputs(5750);
    layer4_outputs(2081) <= not(layer3_outputs(7161));
    layer4_outputs(2082) <= (layer3_outputs(5752)) and (layer3_outputs(3520));
    layer4_outputs(2083) <= not(layer3_outputs(3302));
    layer4_outputs(2084) <= not((layer3_outputs(278)) and (layer3_outputs(4846)));
    layer4_outputs(2085) <= (layer3_outputs(6869)) xor (layer3_outputs(4439));
    layer4_outputs(2086) <= (layer3_outputs(6088)) or (layer3_outputs(4307));
    layer4_outputs(2087) <= not(layer3_outputs(1859));
    layer4_outputs(2088) <= (layer3_outputs(6124)) and not (layer3_outputs(7256));
    layer4_outputs(2089) <= not(layer3_outputs(548)) or (layer3_outputs(998));
    layer4_outputs(2090) <= (layer3_outputs(589)) and not (layer3_outputs(2138));
    layer4_outputs(2091) <= layer3_outputs(7412);
    layer4_outputs(2092) <= not(layer3_outputs(1303));
    layer4_outputs(2093) <= not(layer3_outputs(3203)) or (layer3_outputs(1032));
    layer4_outputs(2094) <= not(layer3_outputs(5122));
    layer4_outputs(2095) <= (layer3_outputs(3188)) xor (layer3_outputs(6788));
    layer4_outputs(2096) <= layer3_outputs(7593);
    layer4_outputs(2097) <= not(layer3_outputs(6270));
    layer4_outputs(2098) <= not(layer3_outputs(1552));
    layer4_outputs(2099) <= (layer3_outputs(6819)) and not (layer3_outputs(674));
    layer4_outputs(2100) <= not((layer3_outputs(4072)) and (layer3_outputs(235)));
    layer4_outputs(2101) <= (layer3_outputs(7356)) and not (layer3_outputs(875));
    layer4_outputs(2102) <= not(layer3_outputs(3833));
    layer4_outputs(2103) <= layer3_outputs(2001);
    layer4_outputs(2104) <= (layer3_outputs(5536)) xor (layer3_outputs(2512));
    layer4_outputs(2105) <= not(layer3_outputs(2356));
    layer4_outputs(2106) <= (layer3_outputs(5054)) xor (layer3_outputs(5346));
    layer4_outputs(2107) <= not(layer3_outputs(1958));
    layer4_outputs(2108) <= not(layer3_outputs(1942));
    layer4_outputs(2109) <= not(layer3_outputs(499));
    layer4_outputs(2110) <= layer3_outputs(4180);
    layer4_outputs(2111) <= layer3_outputs(6038);
    layer4_outputs(2112) <= not((layer3_outputs(2875)) and (layer3_outputs(5580)));
    layer4_outputs(2113) <= not(layer3_outputs(61)) or (layer3_outputs(1723));
    layer4_outputs(2114) <= layer3_outputs(3214);
    layer4_outputs(2115) <= not(layer3_outputs(1936)) or (layer3_outputs(5131));
    layer4_outputs(2116) <= layer3_outputs(5598);
    layer4_outputs(2117) <= (layer3_outputs(2988)) and not (layer3_outputs(1042));
    layer4_outputs(2118) <= not(layer3_outputs(7656)) or (layer3_outputs(5864));
    layer4_outputs(2119) <= (layer3_outputs(4661)) and not (layer3_outputs(655));
    layer4_outputs(2120) <= (layer3_outputs(521)) and not (layer3_outputs(2474));
    layer4_outputs(2121) <= layer3_outputs(5878);
    layer4_outputs(2122) <= layer3_outputs(3910);
    layer4_outputs(2123) <= not(layer3_outputs(6149));
    layer4_outputs(2124) <= layer3_outputs(2244);
    layer4_outputs(2125) <= not(layer3_outputs(2625));
    layer4_outputs(2126) <= not(layer3_outputs(1307));
    layer4_outputs(2127) <= layer3_outputs(5407);
    layer4_outputs(2128) <= not(layer3_outputs(3252)) or (layer3_outputs(3361));
    layer4_outputs(2129) <= not(layer3_outputs(2168)) or (layer3_outputs(3711));
    layer4_outputs(2130) <= (layer3_outputs(88)) or (layer3_outputs(4730));
    layer4_outputs(2131) <= not(layer3_outputs(2481));
    layer4_outputs(2132) <= not(layer3_outputs(6594)) or (layer3_outputs(909));
    layer4_outputs(2133) <= not(layer3_outputs(267));
    layer4_outputs(2134) <= not(layer3_outputs(5123));
    layer4_outputs(2135) <= (layer3_outputs(5680)) xor (layer3_outputs(1747));
    layer4_outputs(2136) <= not((layer3_outputs(3503)) or (layer3_outputs(3229)));
    layer4_outputs(2137) <= (layer3_outputs(2060)) xor (layer3_outputs(4527));
    layer4_outputs(2138) <= layer3_outputs(1431);
    layer4_outputs(2139) <= not(layer3_outputs(541)) or (layer3_outputs(5809));
    layer4_outputs(2140) <= not((layer3_outputs(4014)) xor (layer3_outputs(6743)));
    layer4_outputs(2141) <= '0';
    layer4_outputs(2142) <= layer3_outputs(4966);
    layer4_outputs(2143) <= (layer3_outputs(6488)) and not (layer3_outputs(1317));
    layer4_outputs(2144) <= not((layer3_outputs(5851)) xor (layer3_outputs(1527)));
    layer4_outputs(2145) <= layer3_outputs(12);
    layer4_outputs(2146) <= layer3_outputs(6327);
    layer4_outputs(2147) <= layer3_outputs(7380);
    layer4_outputs(2148) <= not(layer3_outputs(794));
    layer4_outputs(2149) <= not((layer3_outputs(688)) xor (layer3_outputs(2122)));
    layer4_outputs(2150) <= layer3_outputs(7336);
    layer4_outputs(2151) <= not(layer3_outputs(2886));
    layer4_outputs(2152) <= layer3_outputs(6290);
    layer4_outputs(2153) <= layer3_outputs(3588);
    layer4_outputs(2154) <= not((layer3_outputs(3372)) xor (layer3_outputs(3845)));
    layer4_outputs(2155) <= not(layer3_outputs(1975));
    layer4_outputs(2156) <= layer3_outputs(7094);
    layer4_outputs(2157) <= layer3_outputs(5994);
    layer4_outputs(2158) <= layer3_outputs(2680);
    layer4_outputs(2159) <= not(layer3_outputs(5267)) or (layer3_outputs(74));
    layer4_outputs(2160) <= layer3_outputs(5841);
    layer4_outputs(2161) <= layer3_outputs(1095);
    layer4_outputs(2162) <= layer3_outputs(6057);
    layer4_outputs(2163) <= not(layer3_outputs(991));
    layer4_outputs(2164) <= layer3_outputs(5584);
    layer4_outputs(2165) <= not((layer3_outputs(5846)) or (layer3_outputs(5233)));
    layer4_outputs(2166) <= not(layer3_outputs(1945));
    layer4_outputs(2167) <= (layer3_outputs(6859)) or (layer3_outputs(3308));
    layer4_outputs(2168) <= not(layer3_outputs(5957));
    layer4_outputs(2169) <= (layer3_outputs(5016)) and (layer3_outputs(3539));
    layer4_outputs(2170) <= layer3_outputs(2774);
    layer4_outputs(2171) <= (layer3_outputs(1661)) or (layer3_outputs(4549));
    layer4_outputs(2172) <= not(layer3_outputs(6615));
    layer4_outputs(2173) <= layer3_outputs(3068);
    layer4_outputs(2174) <= not(layer3_outputs(3429)) or (layer3_outputs(2884));
    layer4_outputs(2175) <= layer3_outputs(5748);
    layer4_outputs(2176) <= (layer3_outputs(4194)) and not (layer3_outputs(6740));
    layer4_outputs(2177) <= not(layer3_outputs(2636)) or (layer3_outputs(3933));
    layer4_outputs(2178) <= layer3_outputs(1077);
    layer4_outputs(2179) <= (layer3_outputs(642)) and not (layer3_outputs(1487));
    layer4_outputs(2180) <= (layer3_outputs(2843)) and not (layer3_outputs(5648));
    layer4_outputs(2181) <= not((layer3_outputs(2529)) xor (layer3_outputs(5243)));
    layer4_outputs(2182) <= layer3_outputs(5382);
    layer4_outputs(2183) <= not((layer3_outputs(681)) or (layer3_outputs(7265)));
    layer4_outputs(2184) <= (layer3_outputs(2091)) and not (layer3_outputs(191));
    layer4_outputs(2185) <= not((layer3_outputs(726)) xor (layer3_outputs(3385)));
    layer4_outputs(2186) <= not(layer3_outputs(2953));
    layer4_outputs(2187) <= layer3_outputs(1815);
    layer4_outputs(2188) <= not(layer3_outputs(3589));
    layer4_outputs(2189) <= layer3_outputs(2017);
    layer4_outputs(2190) <= not(layer3_outputs(7056)) or (layer3_outputs(5148));
    layer4_outputs(2191) <= not(layer3_outputs(7214));
    layer4_outputs(2192) <= layer3_outputs(6877);
    layer4_outputs(2193) <= layer3_outputs(5670);
    layer4_outputs(2194) <= not((layer3_outputs(3734)) or (layer3_outputs(5253)));
    layer4_outputs(2195) <= (layer3_outputs(7145)) and not (layer3_outputs(993));
    layer4_outputs(2196) <= (layer3_outputs(7173)) xor (layer3_outputs(826));
    layer4_outputs(2197) <= (layer3_outputs(488)) and not (layer3_outputs(3665));
    layer4_outputs(2198) <= layer3_outputs(6073);
    layer4_outputs(2199) <= layer3_outputs(3910);
    layer4_outputs(2200) <= not(layer3_outputs(2092)) or (layer3_outputs(1478));
    layer4_outputs(2201) <= layer3_outputs(2655);
    layer4_outputs(2202) <= layer3_outputs(3178);
    layer4_outputs(2203) <= not(layer3_outputs(3757));
    layer4_outputs(2204) <= layer3_outputs(3179);
    layer4_outputs(2205) <= not(layer3_outputs(3914));
    layer4_outputs(2206) <= not(layer3_outputs(4)) or (layer3_outputs(7481));
    layer4_outputs(2207) <= layer3_outputs(4321);
    layer4_outputs(2208) <= layer3_outputs(6203);
    layer4_outputs(2209) <= layer3_outputs(7169);
    layer4_outputs(2210) <= layer3_outputs(5747);
    layer4_outputs(2211) <= '0';
    layer4_outputs(2212) <= (layer3_outputs(3480)) and not (layer3_outputs(7263));
    layer4_outputs(2213) <= (layer3_outputs(6609)) or (layer3_outputs(776));
    layer4_outputs(2214) <= not(layer3_outputs(1784));
    layer4_outputs(2215) <= (layer3_outputs(7538)) xor (layer3_outputs(5403));
    layer4_outputs(2216) <= not((layer3_outputs(7381)) xor (layer3_outputs(2336)));
    layer4_outputs(2217) <= (layer3_outputs(3800)) and not (layer3_outputs(2188));
    layer4_outputs(2218) <= not(layer3_outputs(221));
    layer4_outputs(2219) <= not(layer3_outputs(7266));
    layer4_outputs(2220) <= (layer3_outputs(939)) and not (layer3_outputs(4097));
    layer4_outputs(2221) <= layer3_outputs(3133);
    layer4_outputs(2222) <= not(layer3_outputs(3831));
    layer4_outputs(2223) <= layer3_outputs(3535);
    layer4_outputs(2224) <= layer3_outputs(5039);
    layer4_outputs(2225) <= not(layer3_outputs(3133));
    layer4_outputs(2226) <= (layer3_outputs(3745)) or (layer3_outputs(3986));
    layer4_outputs(2227) <= (layer3_outputs(2426)) and not (layer3_outputs(2353));
    layer4_outputs(2228) <= not(layer3_outputs(515));
    layer4_outputs(2229) <= layer3_outputs(6085);
    layer4_outputs(2230) <= layer3_outputs(1771);
    layer4_outputs(2231) <= layer3_outputs(6000);
    layer4_outputs(2232) <= layer3_outputs(5415);
    layer4_outputs(2233) <= not(layer3_outputs(4938));
    layer4_outputs(2234) <= layer3_outputs(3338);
    layer4_outputs(2235) <= not(layer3_outputs(7604));
    layer4_outputs(2236) <= (layer3_outputs(2296)) xor (layer3_outputs(2142));
    layer4_outputs(2237) <= not(layer3_outputs(1550));
    layer4_outputs(2238) <= not((layer3_outputs(1561)) or (layer3_outputs(7392)));
    layer4_outputs(2239) <= layer3_outputs(710);
    layer4_outputs(2240) <= layer3_outputs(6303);
    layer4_outputs(2241) <= (layer3_outputs(2926)) xor (layer3_outputs(2744));
    layer4_outputs(2242) <= layer3_outputs(810);
    layer4_outputs(2243) <= layer3_outputs(5811);
    layer4_outputs(2244) <= not(layer3_outputs(4597));
    layer4_outputs(2245) <= not(layer3_outputs(4381));
    layer4_outputs(2246) <= layer3_outputs(3459);
    layer4_outputs(2247) <= layer3_outputs(4671);
    layer4_outputs(2248) <= (layer3_outputs(5498)) and (layer3_outputs(2750));
    layer4_outputs(2249) <= not(layer3_outputs(1953));
    layer4_outputs(2250) <= not(layer3_outputs(298));
    layer4_outputs(2251) <= layer3_outputs(5467);
    layer4_outputs(2252) <= layer3_outputs(5875);
    layer4_outputs(2253) <= not(layer3_outputs(7562));
    layer4_outputs(2254) <= (layer3_outputs(148)) and not (layer3_outputs(2790));
    layer4_outputs(2255) <= layer3_outputs(1986);
    layer4_outputs(2256) <= not((layer3_outputs(737)) xor (layer3_outputs(601)));
    layer4_outputs(2257) <= layer3_outputs(4469);
    layer4_outputs(2258) <= layer3_outputs(4956);
    layer4_outputs(2259) <= (layer3_outputs(118)) and not (layer3_outputs(7518));
    layer4_outputs(2260) <= not(layer3_outputs(706));
    layer4_outputs(2261) <= (layer3_outputs(2051)) and (layer3_outputs(1282));
    layer4_outputs(2262) <= (layer3_outputs(3515)) and (layer3_outputs(5572));
    layer4_outputs(2263) <= (layer3_outputs(4485)) and (layer3_outputs(5050));
    layer4_outputs(2264) <= not((layer3_outputs(6568)) or (layer3_outputs(6291)));
    layer4_outputs(2265) <= (layer3_outputs(6194)) or (layer3_outputs(1082));
    layer4_outputs(2266) <= layer3_outputs(3468);
    layer4_outputs(2267) <= layer3_outputs(4244);
    layer4_outputs(2268) <= (layer3_outputs(1237)) or (layer3_outputs(3504));
    layer4_outputs(2269) <= (layer3_outputs(7304)) or (layer3_outputs(3777));
    layer4_outputs(2270) <= not(layer3_outputs(6922));
    layer4_outputs(2271) <= '1';
    layer4_outputs(2272) <= not(layer3_outputs(5648));
    layer4_outputs(2273) <= not((layer3_outputs(2942)) and (layer3_outputs(4146)));
    layer4_outputs(2274) <= layer3_outputs(2861);
    layer4_outputs(2275) <= (layer3_outputs(4643)) and not (layer3_outputs(1192));
    layer4_outputs(2276) <= (layer3_outputs(5058)) xor (layer3_outputs(643));
    layer4_outputs(2277) <= layer3_outputs(5649);
    layer4_outputs(2278) <= not((layer3_outputs(725)) or (layer3_outputs(3351)));
    layer4_outputs(2279) <= layer3_outputs(6044);
    layer4_outputs(2280) <= not(layer3_outputs(6984));
    layer4_outputs(2281) <= (layer3_outputs(613)) xor (layer3_outputs(990));
    layer4_outputs(2282) <= not(layer3_outputs(7200));
    layer4_outputs(2283) <= not((layer3_outputs(3849)) and (layer3_outputs(4929)));
    layer4_outputs(2284) <= not((layer3_outputs(3115)) and (layer3_outputs(3976)));
    layer4_outputs(2285) <= not((layer3_outputs(3647)) or (layer3_outputs(3506)));
    layer4_outputs(2286) <= (layer3_outputs(85)) or (layer3_outputs(3269));
    layer4_outputs(2287) <= (layer3_outputs(1170)) and not (layer3_outputs(5789));
    layer4_outputs(2288) <= not(layer3_outputs(5661));
    layer4_outputs(2289) <= layer3_outputs(5526);
    layer4_outputs(2290) <= layer3_outputs(4579);
    layer4_outputs(2291) <= not(layer3_outputs(7222));
    layer4_outputs(2292) <= (layer3_outputs(1033)) xor (layer3_outputs(6090));
    layer4_outputs(2293) <= (layer3_outputs(6733)) and (layer3_outputs(4695));
    layer4_outputs(2294) <= layer3_outputs(7373);
    layer4_outputs(2295) <= not(layer3_outputs(2379));
    layer4_outputs(2296) <= not(layer3_outputs(3047));
    layer4_outputs(2297) <= not((layer3_outputs(5806)) and (layer3_outputs(2919)));
    layer4_outputs(2298) <= (layer3_outputs(6042)) and (layer3_outputs(830));
    layer4_outputs(2299) <= not(layer3_outputs(352));
    layer4_outputs(2300) <= not(layer3_outputs(383));
    layer4_outputs(2301) <= layer3_outputs(2441);
    layer4_outputs(2302) <= not(layer3_outputs(2498)) or (layer3_outputs(5446));
    layer4_outputs(2303) <= layer3_outputs(3427);
    layer4_outputs(2304) <= (layer3_outputs(6052)) and not (layer3_outputs(4132));
    layer4_outputs(2305) <= not(layer3_outputs(3542)) or (layer3_outputs(3676));
    layer4_outputs(2306) <= not((layer3_outputs(1884)) or (layer3_outputs(3366)));
    layer4_outputs(2307) <= (layer3_outputs(2516)) or (layer3_outputs(1125));
    layer4_outputs(2308) <= layer3_outputs(6711);
    layer4_outputs(2309) <= (layer3_outputs(2064)) or (layer3_outputs(338));
    layer4_outputs(2310) <= not((layer3_outputs(4573)) and (layer3_outputs(6689)));
    layer4_outputs(2311) <= layer3_outputs(2524);
    layer4_outputs(2312) <= (layer3_outputs(4604)) and (layer3_outputs(6117));
    layer4_outputs(2313) <= (layer3_outputs(2962)) or (layer3_outputs(6306));
    layer4_outputs(2314) <= (layer3_outputs(3696)) and (layer3_outputs(1768));
    layer4_outputs(2315) <= (layer3_outputs(3256)) or (layer3_outputs(1044));
    layer4_outputs(2316) <= not((layer3_outputs(5085)) or (layer3_outputs(7178)));
    layer4_outputs(2317) <= layer3_outputs(6884);
    layer4_outputs(2318) <= not(layer3_outputs(1878));
    layer4_outputs(2319) <= not(layer3_outputs(5529));
    layer4_outputs(2320) <= not(layer3_outputs(3700));
    layer4_outputs(2321) <= (layer3_outputs(2189)) and not (layer3_outputs(7458));
    layer4_outputs(2322) <= not(layer3_outputs(2309));
    layer4_outputs(2323) <= (layer3_outputs(4424)) and (layer3_outputs(519));
    layer4_outputs(2324) <= not(layer3_outputs(1438));
    layer4_outputs(2325) <= (layer3_outputs(7220)) xor (layer3_outputs(6447));
    layer4_outputs(2326) <= layer3_outputs(689);
    layer4_outputs(2327) <= layer3_outputs(3125);
    layer4_outputs(2328) <= not((layer3_outputs(4265)) or (layer3_outputs(4498)));
    layer4_outputs(2329) <= not(layer3_outputs(17));
    layer4_outputs(2330) <= layer3_outputs(893);
    layer4_outputs(2331) <= not(layer3_outputs(2766));
    layer4_outputs(2332) <= (layer3_outputs(4085)) and not (layer3_outputs(6386));
    layer4_outputs(2333) <= not(layer3_outputs(6274)) or (layer3_outputs(6251));
    layer4_outputs(2334) <= (layer3_outputs(841)) and not (layer3_outputs(2591));
    layer4_outputs(2335) <= layer3_outputs(5042);
    layer4_outputs(2336) <= '1';
    layer4_outputs(2337) <= not((layer3_outputs(950)) and (layer3_outputs(789)));
    layer4_outputs(2338) <= layer3_outputs(2628);
    layer4_outputs(2339) <= not(layer3_outputs(2653));
    layer4_outputs(2340) <= layer3_outputs(6062);
    layer4_outputs(2341) <= layer3_outputs(6932);
    layer4_outputs(2342) <= not((layer3_outputs(2810)) and (layer3_outputs(7007)));
    layer4_outputs(2343) <= layer3_outputs(2968);
    layer4_outputs(2344) <= (layer3_outputs(4268)) and not (layer3_outputs(2412));
    layer4_outputs(2345) <= (layer3_outputs(5076)) and not (layer3_outputs(388));
    layer4_outputs(2346) <= not(layer3_outputs(5581));
    layer4_outputs(2347) <= not(layer3_outputs(967));
    layer4_outputs(2348) <= not(layer3_outputs(3428));
    layer4_outputs(2349) <= not((layer3_outputs(6050)) xor (layer3_outputs(5787)));
    layer4_outputs(2350) <= not(layer3_outputs(5452));
    layer4_outputs(2351) <= layer3_outputs(5645);
    layer4_outputs(2352) <= (layer3_outputs(2279)) and (layer3_outputs(6022));
    layer4_outputs(2353) <= not(layer3_outputs(2460));
    layer4_outputs(2354) <= not((layer3_outputs(2855)) xor (layer3_outputs(6639)));
    layer4_outputs(2355) <= (layer3_outputs(3393)) and (layer3_outputs(3472));
    layer4_outputs(2356) <= not(layer3_outputs(6051));
    layer4_outputs(2357) <= layer3_outputs(311);
    layer4_outputs(2358) <= not(layer3_outputs(10));
    layer4_outputs(2359) <= not(layer3_outputs(4747));
    layer4_outputs(2360) <= not((layer3_outputs(7628)) xor (layer3_outputs(7179)));
    layer4_outputs(2361) <= (layer3_outputs(7147)) or (layer3_outputs(4716));
    layer4_outputs(2362) <= not(layer3_outputs(3658));
    layer4_outputs(2363) <= layer3_outputs(2257);
    layer4_outputs(2364) <= (layer3_outputs(4923)) xor (layer3_outputs(7234));
    layer4_outputs(2365) <= '0';
    layer4_outputs(2366) <= not(layer3_outputs(313)) or (layer3_outputs(3340));
    layer4_outputs(2367) <= (layer3_outputs(6495)) xor (layer3_outputs(3822));
    layer4_outputs(2368) <= not(layer3_outputs(3110));
    layer4_outputs(2369) <= (layer3_outputs(4978)) and not (layer3_outputs(7246));
    layer4_outputs(2370) <= not((layer3_outputs(4870)) or (layer3_outputs(3304)));
    layer4_outputs(2371) <= (layer3_outputs(3096)) and not (layer3_outputs(5915));
    layer4_outputs(2372) <= not((layer3_outputs(475)) and (layer3_outputs(3603)));
    layer4_outputs(2373) <= not((layer3_outputs(3953)) xor (layer3_outputs(4862)));
    layer4_outputs(2374) <= layer3_outputs(621);
    layer4_outputs(2375) <= (layer3_outputs(6284)) xor (layer3_outputs(809));
    layer4_outputs(2376) <= (layer3_outputs(5101)) and not (layer3_outputs(3064));
    layer4_outputs(2377) <= layer3_outputs(6882);
    layer4_outputs(2378) <= layer3_outputs(2703);
    layer4_outputs(2379) <= not(layer3_outputs(4968));
    layer4_outputs(2380) <= not(layer3_outputs(3908)) or (layer3_outputs(944));
    layer4_outputs(2381) <= '1';
    layer4_outputs(2382) <= layer3_outputs(5874);
    layer4_outputs(2383) <= layer3_outputs(2718);
    layer4_outputs(2384) <= not(layer3_outputs(3798));
    layer4_outputs(2385) <= not(layer3_outputs(6857));
    layer4_outputs(2386) <= layer3_outputs(4189);
    layer4_outputs(2387) <= (layer3_outputs(6388)) and (layer3_outputs(6957));
    layer4_outputs(2388) <= layer3_outputs(5709);
    layer4_outputs(2389) <= not(layer3_outputs(3414)) or (layer3_outputs(4372));
    layer4_outputs(2390) <= not((layer3_outputs(3134)) or (layer3_outputs(359)));
    layer4_outputs(2391) <= not(layer3_outputs(7193));
    layer4_outputs(2392) <= (layer3_outputs(3538)) and not (layer3_outputs(6584));
    layer4_outputs(2393) <= (layer3_outputs(3772)) and (layer3_outputs(7577));
    layer4_outputs(2394) <= not((layer3_outputs(2575)) and (layer3_outputs(2806)));
    layer4_outputs(2395) <= (layer3_outputs(4520)) and not (layer3_outputs(77));
    layer4_outputs(2396) <= layer3_outputs(6869);
    layer4_outputs(2397) <= layer3_outputs(4547);
    layer4_outputs(2398) <= layer3_outputs(5012);
    layer4_outputs(2399) <= (layer3_outputs(5356)) xor (layer3_outputs(7228));
    layer4_outputs(2400) <= not(layer3_outputs(5809)) or (layer3_outputs(6996));
    layer4_outputs(2401) <= not((layer3_outputs(1959)) and (layer3_outputs(6948)));
    layer4_outputs(2402) <= not(layer3_outputs(1267)) or (layer3_outputs(7496));
    layer4_outputs(2403) <= (layer3_outputs(910)) or (layer3_outputs(2599));
    layer4_outputs(2404) <= layer3_outputs(881);
    layer4_outputs(2405) <= not(layer3_outputs(1011));
    layer4_outputs(2406) <= (layer3_outputs(6944)) xor (layer3_outputs(979));
    layer4_outputs(2407) <= not((layer3_outputs(6129)) xor (layer3_outputs(4377)));
    layer4_outputs(2408) <= not((layer3_outputs(4403)) and (layer3_outputs(4446)));
    layer4_outputs(2409) <= not(layer3_outputs(5011));
    layer4_outputs(2410) <= not(layer3_outputs(2317));
    layer4_outputs(2411) <= not(layer3_outputs(5471));
    layer4_outputs(2412) <= not(layer3_outputs(2726));
    layer4_outputs(2413) <= (layer3_outputs(446)) and not (layer3_outputs(1944));
    layer4_outputs(2414) <= (layer3_outputs(7284)) and not (layer3_outputs(4092));
    layer4_outputs(2415) <= not(layer3_outputs(588));
    layer4_outputs(2416) <= not(layer3_outputs(7515));
    layer4_outputs(2417) <= layer3_outputs(4423);
    layer4_outputs(2418) <= (layer3_outputs(5160)) and (layer3_outputs(3802));
    layer4_outputs(2419) <= (layer3_outputs(1175)) and (layer3_outputs(1554));
    layer4_outputs(2420) <= not(layer3_outputs(6390));
    layer4_outputs(2421) <= (layer3_outputs(4640)) or (layer3_outputs(7110));
    layer4_outputs(2422) <= not(layer3_outputs(1424));
    layer4_outputs(2423) <= not((layer3_outputs(1847)) and (layer3_outputs(7252)));
    layer4_outputs(2424) <= layer3_outputs(5671);
    layer4_outputs(2425) <= (layer3_outputs(1300)) or (layer3_outputs(5517));
    layer4_outputs(2426) <= not(layer3_outputs(6508)) or (layer3_outputs(6216));
    layer4_outputs(2427) <= (layer3_outputs(6028)) or (layer3_outputs(5398));
    layer4_outputs(2428) <= not((layer3_outputs(7250)) and (layer3_outputs(4388)));
    layer4_outputs(2429) <= not((layer3_outputs(2491)) and (layer3_outputs(4681)));
    layer4_outputs(2430) <= not((layer3_outputs(4622)) xor (layer3_outputs(3472)));
    layer4_outputs(2431) <= layer3_outputs(4249);
    layer4_outputs(2432) <= '0';
    layer4_outputs(2433) <= layer3_outputs(1911);
    layer4_outputs(2434) <= not(layer3_outputs(5431));
    layer4_outputs(2435) <= layer3_outputs(1614);
    layer4_outputs(2436) <= layer3_outputs(3315);
    layer4_outputs(2437) <= layer3_outputs(2308);
    layer4_outputs(2438) <= not(layer3_outputs(6180));
    layer4_outputs(2439) <= not(layer3_outputs(6108)) or (layer3_outputs(7399));
    layer4_outputs(2440) <= (layer3_outputs(4817)) and not (layer3_outputs(3304));
    layer4_outputs(2441) <= not(layer3_outputs(2911));
    layer4_outputs(2442) <= layer3_outputs(3728);
    layer4_outputs(2443) <= not(layer3_outputs(7543)) or (layer3_outputs(3282));
    layer4_outputs(2444) <= (layer3_outputs(5821)) and not (layer3_outputs(7414));
    layer4_outputs(2445) <= (layer3_outputs(3617)) xor (layer3_outputs(6198));
    layer4_outputs(2446) <= (layer3_outputs(510)) or (layer3_outputs(1911));
    layer4_outputs(2447) <= (layer3_outputs(2267)) xor (layer3_outputs(6730));
    layer4_outputs(2448) <= not(layer3_outputs(3928));
    layer4_outputs(2449) <= not(layer3_outputs(7041)) or (layer3_outputs(3126));
    layer4_outputs(2450) <= not(layer3_outputs(3582)) or (layer3_outputs(6523));
    layer4_outputs(2451) <= layer3_outputs(5407);
    layer4_outputs(2452) <= not(layer3_outputs(2287)) or (layer3_outputs(5611));
    layer4_outputs(2453) <= not(layer3_outputs(2668));
    layer4_outputs(2454) <= (layer3_outputs(4665)) or (layer3_outputs(382));
    layer4_outputs(2455) <= not(layer3_outputs(4799));
    layer4_outputs(2456) <= not(layer3_outputs(756));
    layer4_outputs(2457) <= not((layer3_outputs(7406)) or (layer3_outputs(2603)));
    layer4_outputs(2458) <= not(layer3_outputs(2358)) or (layer3_outputs(439));
    layer4_outputs(2459) <= (layer3_outputs(862)) or (layer3_outputs(3002));
    layer4_outputs(2460) <= not(layer3_outputs(4310));
    layer4_outputs(2461) <= (layer3_outputs(3069)) and not (layer3_outputs(3423));
    layer4_outputs(2462) <= (layer3_outputs(1596)) and not (layer3_outputs(6363));
    layer4_outputs(2463) <= not(layer3_outputs(3754));
    layer4_outputs(2464) <= not(layer3_outputs(1279));
    layer4_outputs(2465) <= not((layer3_outputs(4603)) or (layer3_outputs(7081)));
    layer4_outputs(2466) <= (layer3_outputs(1076)) xor (layer3_outputs(7195));
    layer4_outputs(2467) <= (layer3_outputs(1740)) xor (layer3_outputs(3636));
    layer4_outputs(2468) <= (layer3_outputs(5303)) or (layer3_outputs(4280));
    layer4_outputs(2469) <= not(layer3_outputs(180));
    layer4_outputs(2470) <= (layer3_outputs(5818)) and not (layer3_outputs(3872));
    layer4_outputs(2471) <= layer3_outputs(6736);
    layer4_outputs(2472) <= not(layer3_outputs(5079));
    layer4_outputs(2473) <= layer3_outputs(2225);
    layer4_outputs(2474) <= not(layer3_outputs(6514));
    layer4_outputs(2475) <= layer3_outputs(2492);
    layer4_outputs(2476) <= layer3_outputs(3821);
    layer4_outputs(2477) <= layer3_outputs(1495);
    layer4_outputs(2478) <= not(layer3_outputs(5464));
    layer4_outputs(2479) <= layer3_outputs(129);
    layer4_outputs(2480) <= '1';
    layer4_outputs(2481) <= layer3_outputs(5630);
    layer4_outputs(2482) <= layer3_outputs(2442);
    layer4_outputs(2483) <= (layer3_outputs(856)) and (layer3_outputs(7388));
    layer4_outputs(2484) <= layer3_outputs(6513);
    layer4_outputs(2485) <= not(layer3_outputs(4315));
    layer4_outputs(2486) <= not(layer3_outputs(3521));
    layer4_outputs(2487) <= not((layer3_outputs(3012)) and (layer3_outputs(5487)));
    layer4_outputs(2488) <= not((layer3_outputs(3370)) xor (layer3_outputs(7096)));
    layer4_outputs(2489) <= (layer3_outputs(3965)) and not (layer3_outputs(2236));
    layer4_outputs(2490) <= not((layer3_outputs(7666)) or (layer3_outputs(1895)));
    layer4_outputs(2491) <= not((layer3_outputs(6723)) or (layer3_outputs(1853)));
    layer4_outputs(2492) <= (layer3_outputs(4230)) xor (layer3_outputs(2441));
    layer4_outputs(2493) <= not((layer3_outputs(7242)) or (layer3_outputs(3732)));
    layer4_outputs(2494) <= layer3_outputs(1385);
    layer4_outputs(2495) <= layer3_outputs(6535);
    layer4_outputs(2496) <= not((layer3_outputs(2070)) and (layer3_outputs(4998)));
    layer4_outputs(2497) <= (layer3_outputs(3249)) xor (layer3_outputs(2447));
    layer4_outputs(2498) <= layer3_outputs(3092);
    layer4_outputs(2499) <= not(layer3_outputs(7610));
    layer4_outputs(2500) <= not(layer3_outputs(275));
    layer4_outputs(2501) <= layer3_outputs(6687);
    layer4_outputs(2502) <= not(layer3_outputs(6244));
    layer4_outputs(2503) <= (layer3_outputs(5998)) and not (layer3_outputs(105));
    layer4_outputs(2504) <= not(layer3_outputs(6235));
    layer4_outputs(2505) <= (layer3_outputs(6517)) and (layer3_outputs(735));
    layer4_outputs(2506) <= layer3_outputs(2931);
    layer4_outputs(2507) <= (layer3_outputs(5322)) or (layer3_outputs(2598));
    layer4_outputs(2508) <= not((layer3_outputs(1719)) or (layer3_outputs(6032)));
    layer4_outputs(2509) <= (layer3_outputs(3768)) and (layer3_outputs(1044));
    layer4_outputs(2510) <= (layer3_outputs(6640)) and not (layer3_outputs(4880));
    layer4_outputs(2511) <= not(layer3_outputs(7611));
    layer4_outputs(2512) <= (layer3_outputs(2850)) and not (layer3_outputs(4035));
    layer4_outputs(2513) <= not(layer3_outputs(5745));
    layer4_outputs(2514) <= not(layer3_outputs(4008));
    layer4_outputs(2515) <= (layer3_outputs(4076)) and not (layer3_outputs(2559));
    layer4_outputs(2516) <= not(layer3_outputs(4783));
    layer4_outputs(2517) <= (layer3_outputs(4166)) and (layer3_outputs(6358));
    layer4_outputs(2518) <= not(layer3_outputs(6979)) or (layer3_outputs(4801));
    layer4_outputs(2519) <= (layer3_outputs(684)) and not (layer3_outputs(6661));
    layer4_outputs(2520) <= (layer3_outputs(193)) xor (layer3_outputs(3205));
    layer4_outputs(2521) <= not(layer3_outputs(4896)) or (layer3_outputs(1923));
    layer4_outputs(2522) <= (layer3_outputs(6482)) and not (layer3_outputs(7231));
    layer4_outputs(2523) <= not((layer3_outputs(4263)) xor (layer3_outputs(4080)));
    layer4_outputs(2524) <= layer3_outputs(4040);
    layer4_outputs(2525) <= (layer3_outputs(2695)) xor (layer3_outputs(4953));
    layer4_outputs(2526) <= layer3_outputs(4237);
    layer4_outputs(2527) <= not(layer3_outputs(7150));
    layer4_outputs(2528) <= layer3_outputs(1157);
    layer4_outputs(2529) <= not(layer3_outputs(4823));
    layer4_outputs(2530) <= layer3_outputs(6843);
    layer4_outputs(2531) <= not(layer3_outputs(2381));
    layer4_outputs(2532) <= layer3_outputs(806);
    layer4_outputs(2533) <= not((layer3_outputs(4219)) and (layer3_outputs(1280)));
    layer4_outputs(2534) <= (layer3_outputs(5011)) xor (layer3_outputs(797));
    layer4_outputs(2535) <= not(layer3_outputs(5431));
    layer4_outputs(2536) <= not(layer3_outputs(1568));
    layer4_outputs(2537) <= layer3_outputs(1149);
    layer4_outputs(2538) <= not(layer3_outputs(879));
    layer4_outputs(2539) <= (layer3_outputs(6584)) or (layer3_outputs(3913));
    layer4_outputs(2540) <= (layer3_outputs(4622)) or (layer3_outputs(1955));
    layer4_outputs(2541) <= not(layer3_outputs(436)) or (layer3_outputs(434));
    layer4_outputs(2542) <= not(layer3_outputs(4604)) or (layer3_outputs(1744));
    layer4_outputs(2543) <= layer3_outputs(6632);
    layer4_outputs(2544) <= not((layer3_outputs(7551)) xor (layer3_outputs(6924)));
    layer4_outputs(2545) <= layer3_outputs(7408);
    layer4_outputs(2546) <= layer3_outputs(1472);
    layer4_outputs(2547) <= layer3_outputs(5113);
    layer4_outputs(2548) <= (layer3_outputs(1990)) and (layer3_outputs(2026));
    layer4_outputs(2549) <= not(layer3_outputs(7240)) or (layer3_outputs(3545));
    layer4_outputs(2550) <= (layer3_outputs(2129)) and (layer3_outputs(3422));
    layer4_outputs(2551) <= (layer3_outputs(5419)) and not (layer3_outputs(4093));
    layer4_outputs(2552) <= not(layer3_outputs(7494));
    layer4_outputs(2553) <= not(layer3_outputs(6656));
    layer4_outputs(2554) <= (layer3_outputs(846)) xor (layer3_outputs(4748));
    layer4_outputs(2555) <= (layer3_outputs(957)) or (layer3_outputs(1751));
    layer4_outputs(2556) <= not(layer3_outputs(5634));
    layer4_outputs(2557) <= (layer3_outputs(7001)) or (layer3_outputs(3053));
    layer4_outputs(2558) <= layer3_outputs(380);
    layer4_outputs(2559) <= not(layer3_outputs(7508));
    layer4_outputs(2560) <= not(layer3_outputs(1681)) or (layer3_outputs(2854));
    layer4_outputs(2561) <= (layer3_outputs(3945)) xor (layer3_outputs(3155));
    layer4_outputs(2562) <= (layer3_outputs(4781)) or (layer3_outputs(3951));
    layer4_outputs(2563) <= not(layer3_outputs(654));
    layer4_outputs(2564) <= layer3_outputs(6538);
    layer4_outputs(2565) <= not(layer3_outputs(6285));
    layer4_outputs(2566) <= (layer3_outputs(308)) and (layer3_outputs(2268));
    layer4_outputs(2567) <= not(layer3_outputs(2967));
    layer4_outputs(2568) <= not(layer3_outputs(4741));
    layer4_outputs(2569) <= layer3_outputs(3171);
    layer4_outputs(2570) <= (layer3_outputs(819)) and not (layer3_outputs(905));
    layer4_outputs(2571) <= (layer3_outputs(4571)) or (layer3_outputs(5595));
    layer4_outputs(2572) <= not((layer3_outputs(1180)) xor (layer3_outputs(425)));
    layer4_outputs(2573) <= layer3_outputs(4005);
    layer4_outputs(2574) <= not(layer3_outputs(2360));
    layer4_outputs(2575) <= (layer3_outputs(4160)) or (layer3_outputs(6156));
    layer4_outputs(2576) <= not((layer3_outputs(7407)) or (layer3_outputs(6464)));
    layer4_outputs(2577) <= not((layer3_outputs(260)) or (layer3_outputs(2697)));
    layer4_outputs(2578) <= not(layer3_outputs(1356));
    layer4_outputs(2579) <= (layer3_outputs(3100)) and (layer3_outputs(3539));
    layer4_outputs(2580) <= layer3_outputs(1201);
    layer4_outputs(2581) <= (layer3_outputs(4824)) and not (layer3_outputs(7667));
    layer4_outputs(2582) <= (layer3_outputs(1449)) xor (layer3_outputs(6612));
    layer4_outputs(2583) <= not(layer3_outputs(4276));
    layer4_outputs(2584) <= (layer3_outputs(2903)) xor (layer3_outputs(1007));
    layer4_outputs(2585) <= not(layer3_outputs(7609));
    layer4_outputs(2586) <= layer3_outputs(2574);
    layer4_outputs(2587) <= layer3_outputs(5162);
    layer4_outputs(2588) <= (layer3_outputs(1971)) and not (layer3_outputs(6479));
    layer4_outputs(2589) <= layer3_outputs(5673);
    layer4_outputs(2590) <= layer3_outputs(2425);
    layer4_outputs(2591) <= layer3_outputs(6835);
    layer4_outputs(2592) <= not(layer3_outputs(4172));
    layer4_outputs(2593) <= '0';
    layer4_outputs(2594) <= not(layer3_outputs(3772));
    layer4_outputs(2595) <= layer3_outputs(6105);
    layer4_outputs(2596) <= layer3_outputs(5406);
    layer4_outputs(2597) <= (layer3_outputs(7034)) and not (layer3_outputs(6127));
    layer4_outputs(2598) <= not(layer3_outputs(7058));
    layer4_outputs(2599) <= not(layer3_outputs(2192));
    layer4_outputs(2600) <= (layer3_outputs(3242)) and not (layer3_outputs(2939));
    layer4_outputs(2601) <= not((layer3_outputs(4450)) and (layer3_outputs(1351)));
    layer4_outputs(2602) <= not(layer3_outputs(2392));
    layer4_outputs(2603) <= (layer3_outputs(5939)) or (layer3_outputs(5830));
    layer4_outputs(2604) <= not(layer3_outputs(6707)) or (layer3_outputs(1189));
    layer4_outputs(2605) <= not(layer3_outputs(3585));
    layer4_outputs(2606) <= layer3_outputs(4966);
    layer4_outputs(2607) <= layer3_outputs(1762);
    layer4_outputs(2608) <= (layer3_outputs(6798)) or (layer3_outputs(2617));
    layer4_outputs(2609) <= not(layer3_outputs(2900));
    layer4_outputs(2610) <= layer3_outputs(926);
    layer4_outputs(2611) <= layer3_outputs(3762);
    layer4_outputs(2612) <= not(layer3_outputs(272));
    layer4_outputs(2613) <= not(layer3_outputs(3458));
    layer4_outputs(2614) <= not((layer3_outputs(2912)) and (layer3_outputs(5270)));
    layer4_outputs(2615) <= not(layer3_outputs(1988));
    layer4_outputs(2616) <= layer3_outputs(2797);
    layer4_outputs(2617) <= not(layer3_outputs(4638));
    layer4_outputs(2618) <= (layer3_outputs(1330)) and not (layer3_outputs(7331));
    layer4_outputs(2619) <= not((layer3_outputs(6236)) xor (layer3_outputs(3002)));
    layer4_outputs(2620) <= not(layer3_outputs(5862));
    layer4_outputs(2621) <= not(layer3_outputs(588)) or (layer3_outputs(6527));
    layer4_outputs(2622) <= not(layer3_outputs(4285));
    layer4_outputs(2623) <= not((layer3_outputs(7519)) and (layer3_outputs(1803)));
    layer4_outputs(2624) <= not(layer3_outputs(3235));
    layer4_outputs(2625) <= layer3_outputs(955);
    layer4_outputs(2626) <= not((layer3_outputs(5459)) and (layer3_outputs(2916)));
    layer4_outputs(2627) <= layer3_outputs(1398);
    layer4_outputs(2628) <= (layer3_outputs(5098)) and (layer3_outputs(3605));
    layer4_outputs(2629) <= layer3_outputs(7432);
    layer4_outputs(2630) <= not(layer3_outputs(1386)) or (layer3_outputs(3468));
    layer4_outputs(2631) <= layer3_outputs(4447);
    layer4_outputs(2632) <= not(layer3_outputs(4580)) or (layer3_outputs(3314));
    layer4_outputs(2633) <= layer3_outputs(4);
    layer4_outputs(2634) <= (layer3_outputs(3802)) and (layer3_outputs(570));
    layer4_outputs(2635) <= layer3_outputs(5633);
    layer4_outputs(2636) <= not(layer3_outputs(2943));
    layer4_outputs(2637) <= not(layer3_outputs(6068)) or (layer3_outputs(6986));
    layer4_outputs(2638) <= layer3_outputs(552);
    layer4_outputs(2639) <= not(layer3_outputs(1611));
    layer4_outputs(2640) <= (layer3_outputs(1548)) xor (layer3_outputs(4003));
    layer4_outputs(2641) <= '1';
    layer4_outputs(2642) <= not(layer3_outputs(2249)) or (layer3_outputs(6800));
    layer4_outputs(2643) <= (layer3_outputs(3207)) or (layer3_outputs(5982));
    layer4_outputs(2644) <= layer3_outputs(1255);
    layer4_outputs(2645) <= layer3_outputs(2587);
    layer4_outputs(2646) <= not((layer3_outputs(861)) xor (layer3_outputs(1262)));
    layer4_outputs(2647) <= not((layer3_outputs(1132)) xor (layer3_outputs(6078)));
    layer4_outputs(2648) <= not(layer3_outputs(2053));
    layer4_outputs(2649) <= not(layer3_outputs(339));
    layer4_outputs(2650) <= not(layer3_outputs(5140));
    layer4_outputs(2651) <= layer3_outputs(5456);
    layer4_outputs(2652) <= not(layer3_outputs(4065));
    layer4_outputs(2653) <= layer3_outputs(6731);
    layer4_outputs(2654) <= layer3_outputs(6783);
    layer4_outputs(2655) <= (layer3_outputs(3424)) and (layer3_outputs(4494));
    layer4_outputs(2656) <= not((layer3_outputs(6179)) or (layer3_outputs(7268)));
    layer4_outputs(2657) <= (layer3_outputs(3065)) xor (layer3_outputs(4913));
    layer4_outputs(2658) <= layer3_outputs(2414);
    layer4_outputs(2659) <= layer3_outputs(3761);
    layer4_outputs(2660) <= not(layer3_outputs(6913));
    layer4_outputs(2661) <= (layer3_outputs(6973)) xor (layer3_outputs(5251));
    layer4_outputs(2662) <= not(layer3_outputs(3208)) or (layer3_outputs(5447));
    layer4_outputs(2663) <= not(layer3_outputs(3583));
    layer4_outputs(2664) <= not(layer3_outputs(2535));
    layer4_outputs(2665) <= not((layer3_outputs(2267)) and (layer3_outputs(5474)));
    layer4_outputs(2666) <= (layer3_outputs(4533)) or (layer3_outputs(3435));
    layer4_outputs(2667) <= not(layer3_outputs(185)) or (layer3_outputs(1735));
    layer4_outputs(2668) <= not((layer3_outputs(5485)) xor (layer3_outputs(3884)));
    layer4_outputs(2669) <= layer3_outputs(6755);
    layer4_outputs(2670) <= not(layer3_outputs(5345));
    layer4_outputs(2671) <= layer3_outputs(99);
    layer4_outputs(2672) <= (layer3_outputs(1039)) and (layer3_outputs(2187));
    layer4_outputs(2673) <= (layer3_outputs(5340)) and not (layer3_outputs(5));
    layer4_outputs(2674) <= not((layer3_outputs(456)) or (layer3_outputs(1159)));
    layer4_outputs(2675) <= not(layer3_outputs(2186));
    layer4_outputs(2676) <= not((layer3_outputs(4246)) or (layer3_outputs(1912)));
    layer4_outputs(2677) <= not((layer3_outputs(1696)) or (layer3_outputs(4628)));
    layer4_outputs(2678) <= (layer3_outputs(6012)) xor (layer3_outputs(5628));
    layer4_outputs(2679) <= not(layer3_outputs(7227)) or (layer3_outputs(1718));
    layer4_outputs(2680) <= layer3_outputs(5220);
    layer4_outputs(2681) <= (layer3_outputs(1232)) or (layer3_outputs(2253));
    layer4_outputs(2682) <= not(layer3_outputs(5582));
    layer4_outputs(2683) <= not(layer3_outputs(799));
    layer4_outputs(2684) <= layer3_outputs(5115);
    layer4_outputs(2685) <= not(layer3_outputs(2850)) or (layer3_outputs(1762));
    layer4_outputs(2686) <= (layer3_outputs(2002)) and (layer3_outputs(1338));
    layer4_outputs(2687) <= layer3_outputs(6028);
    layer4_outputs(2688) <= not(layer3_outputs(962));
    layer4_outputs(2689) <= not(layer3_outputs(4668));
    layer4_outputs(2690) <= not(layer3_outputs(5618));
    layer4_outputs(2691) <= not(layer3_outputs(4128)) or (layer3_outputs(6753));
    layer4_outputs(2692) <= layer3_outputs(4338);
    layer4_outputs(2693) <= not(layer3_outputs(1244));
    layer4_outputs(2694) <= (layer3_outputs(3167)) xor (layer3_outputs(6093));
    layer4_outputs(2695) <= not(layer3_outputs(1050));
    layer4_outputs(2696) <= (layer3_outputs(1161)) or (layer3_outputs(4990));
    layer4_outputs(2697) <= (layer3_outputs(6242)) and (layer3_outputs(5722));
    layer4_outputs(2698) <= not(layer3_outputs(6545));
    layer4_outputs(2699) <= layer3_outputs(2675);
    layer4_outputs(2700) <= layer3_outputs(7166);
    layer4_outputs(2701) <= layer3_outputs(3079);
    layer4_outputs(2702) <= not(layer3_outputs(5587));
    layer4_outputs(2703) <= not(layer3_outputs(2761));
    layer4_outputs(2704) <= (layer3_outputs(6789)) and not (layer3_outputs(3932));
    layer4_outputs(2705) <= layer3_outputs(7262);
    layer4_outputs(2706) <= layer3_outputs(7017);
    layer4_outputs(2707) <= not(layer3_outputs(3221));
    layer4_outputs(2708) <= layer3_outputs(2595);
    layer4_outputs(2709) <= (layer3_outputs(3267)) and not (layer3_outputs(7627));
    layer4_outputs(2710) <= not(layer3_outputs(5533)) or (layer3_outputs(4871));
    layer4_outputs(2711) <= layer3_outputs(6829);
    layer4_outputs(2712) <= not((layer3_outputs(440)) or (layer3_outputs(6433)));
    layer4_outputs(2713) <= (layer3_outputs(2986)) and not (layer3_outputs(1393));
    layer4_outputs(2714) <= not((layer3_outputs(3906)) and (layer3_outputs(7424)));
    layer4_outputs(2715) <= layer3_outputs(774);
    layer4_outputs(2716) <= not(layer3_outputs(5360));
    layer4_outputs(2717) <= not((layer3_outputs(1925)) and (layer3_outputs(2730)));
    layer4_outputs(2718) <= layer3_outputs(6805);
    layer4_outputs(2719) <= layer3_outputs(189);
    layer4_outputs(2720) <= layer3_outputs(4811);
    layer4_outputs(2721) <= not(layer3_outputs(2051));
    layer4_outputs(2722) <= layer3_outputs(5586);
    layer4_outputs(2723) <= (layer3_outputs(565)) or (layer3_outputs(5254));
    layer4_outputs(2724) <= not(layer3_outputs(235));
    layer4_outputs(2725) <= layer3_outputs(7107);
    layer4_outputs(2726) <= (layer3_outputs(484)) xor (layer3_outputs(7487));
    layer4_outputs(2727) <= layer3_outputs(5387);
    layer4_outputs(2728) <= (layer3_outputs(1073)) xor (layer3_outputs(2595));
    layer4_outputs(2729) <= layer3_outputs(4550);
    layer4_outputs(2730) <= not(layer3_outputs(1364));
    layer4_outputs(2731) <= (layer3_outputs(1881)) and not (layer3_outputs(5482));
    layer4_outputs(2732) <= layer3_outputs(2135);
    layer4_outputs(2733) <= not(layer3_outputs(1644));
    layer4_outputs(2734) <= not((layer3_outputs(4694)) or (layer3_outputs(2904)));
    layer4_outputs(2735) <= not(layer3_outputs(3198)) or (layer3_outputs(7580));
    layer4_outputs(2736) <= (layer3_outputs(50)) and not (layer3_outputs(223));
    layer4_outputs(2737) <= not(layer3_outputs(6343));
    layer4_outputs(2738) <= (layer3_outputs(3497)) and (layer3_outputs(2866));
    layer4_outputs(2739) <= not(layer3_outputs(5576));
    layer4_outputs(2740) <= layer3_outputs(7434);
    layer4_outputs(2741) <= (layer3_outputs(2707)) or (layer3_outputs(492));
    layer4_outputs(2742) <= (layer3_outputs(7117)) and not (layer3_outputs(345));
    layer4_outputs(2743) <= not((layer3_outputs(3051)) or (layer3_outputs(6766)));
    layer4_outputs(2744) <= (layer3_outputs(315)) xor (layer3_outputs(7426));
    layer4_outputs(2745) <= not((layer3_outputs(7142)) or (layer3_outputs(2541)));
    layer4_outputs(2746) <= '0';
    layer4_outputs(2747) <= (layer3_outputs(3567)) xor (layer3_outputs(1729));
    layer4_outputs(2748) <= not(layer3_outputs(1534));
    layer4_outputs(2749) <= not((layer3_outputs(7162)) or (layer3_outputs(5825)));
    layer4_outputs(2750) <= not(layer3_outputs(5374));
    layer4_outputs(2751) <= (layer3_outputs(2277)) and not (layer3_outputs(403));
    layer4_outputs(2752) <= not(layer3_outputs(4772));
    layer4_outputs(2753) <= not((layer3_outputs(2836)) xor (layer3_outputs(1358)));
    layer4_outputs(2754) <= layer3_outputs(6547);
    layer4_outputs(2755) <= not(layer3_outputs(7330)) or (layer3_outputs(6996));
    layer4_outputs(2756) <= not(layer3_outputs(4057)) or (layer3_outputs(506));
    layer4_outputs(2757) <= not(layer3_outputs(3095));
    layer4_outputs(2758) <= not((layer3_outputs(785)) or (layer3_outputs(6243)));
    layer4_outputs(2759) <= not((layer3_outputs(6694)) and (layer3_outputs(6616)));
    layer4_outputs(2760) <= not(layer3_outputs(3524));
    layer4_outputs(2761) <= (layer3_outputs(1973)) xor (layer3_outputs(669));
    layer4_outputs(2762) <= (layer3_outputs(1207)) xor (layer3_outputs(5502));
    layer4_outputs(2763) <= (layer3_outputs(6345)) and not (layer3_outputs(2228));
    layer4_outputs(2764) <= not(layer3_outputs(4849));
    layer4_outputs(2765) <= (layer3_outputs(6688)) xor (layer3_outputs(4073));
    layer4_outputs(2766) <= layer3_outputs(637);
    layer4_outputs(2767) <= (layer3_outputs(2780)) or (layer3_outputs(4185));
    layer4_outputs(2768) <= (layer3_outputs(2945)) xor (layer3_outputs(1776));
    layer4_outputs(2769) <= not(layer3_outputs(2050));
    layer4_outputs(2770) <= (layer3_outputs(1337)) xor (layer3_outputs(4538));
    layer4_outputs(2771) <= layer3_outputs(5232);
    layer4_outputs(2772) <= not((layer3_outputs(4143)) or (layer3_outputs(2832)));
    layer4_outputs(2773) <= layer3_outputs(6667);
    layer4_outputs(2774) <= not(layer3_outputs(1130)) or (layer3_outputs(6656));
    layer4_outputs(2775) <= layer3_outputs(6459);
    layer4_outputs(2776) <= layer3_outputs(3496);
    layer4_outputs(2777) <= layer3_outputs(1213);
    layer4_outputs(2778) <= not(layer3_outputs(4568));
    layer4_outputs(2779) <= (layer3_outputs(119)) and not (layer3_outputs(6781));
    layer4_outputs(2780) <= not((layer3_outputs(6299)) xor (layer3_outputs(763)));
    layer4_outputs(2781) <= layer3_outputs(3613);
    layer4_outputs(2782) <= (layer3_outputs(3146)) and not (layer3_outputs(3317));
    layer4_outputs(2783) <= not(layer3_outputs(569));
    layer4_outputs(2784) <= not(layer3_outputs(1490));
    layer4_outputs(2785) <= (layer3_outputs(3115)) xor (layer3_outputs(2258));
    layer4_outputs(2786) <= (layer3_outputs(4517)) and (layer3_outputs(1568));
    layer4_outputs(2787) <= (layer3_outputs(410)) and not (layer3_outputs(4618));
    layer4_outputs(2788) <= layer3_outputs(7012);
    layer4_outputs(2789) <= not(layer3_outputs(3718)) or (layer3_outputs(3675));
    layer4_outputs(2790) <= not((layer3_outputs(6135)) or (layer3_outputs(5744)));
    layer4_outputs(2791) <= layer3_outputs(4169);
    layer4_outputs(2792) <= (layer3_outputs(7254)) and (layer3_outputs(976));
    layer4_outputs(2793) <= layer3_outputs(3437);
    layer4_outputs(2794) <= (layer3_outputs(1841)) or (layer3_outputs(174));
    layer4_outputs(2795) <= not(layer3_outputs(7098));
    layer4_outputs(2796) <= not((layer3_outputs(5075)) and (layer3_outputs(4444)));
    layer4_outputs(2797) <= not((layer3_outputs(7062)) xor (layer3_outputs(7148)));
    layer4_outputs(2798) <= layer3_outputs(3897);
    layer4_outputs(2799) <= layer3_outputs(5252);
    layer4_outputs(2800) <= not(layer3_outputs(1714));
    layer4_outputs(2801) <= not((layer3_outputs(1660)) and (layer3_outputs(307)));
    layer4_outputs(2802) <= (layer3_outputs(365)) and (layer3_outputs(5904));
    layer4_outputs(2803) <= not((layer3_outputs(11)) and (layer3_outputs(2869)));
    layer4_outputs(2804) <= not((layer3_outputs(4991)) or (layer3_outputs(3207)));
    layer4_outputs(2805) <= not((layer3_outputs(1127)) or (layer3_outputs(169)));
    layer4_outputs(2806) <= not(layer3_outputs(1737)) or (layer3_outputs(336));
    layer4_outputs(2807) <= not((layer3_outputs(4969)) or (layer3_outputs(2974)));
    layer4_outputs(2808) <= (layer3_outputs(1439)) or (layer3_outputs(3188));
    layer4_outputs(2809) <= layer3_outputs(229);
    layer4_outputs(2810) <= not(layer3_outputs(4610));
    layer4_outputs(2811) <= layer3_outputs(5028);
    layer4_outputs(2812) <= layer3_outputs(6749);
    layer4_outputs(2813) <= not((layer3_outputs(7226)) or (layer3_outputs(4024)));
    layer4_outputs(2814) <= not((layer3_outputs(73)) xor (layer3_outputs(6318)));
    layer4_outputs(2815) <= (layer3_outputs(4410)) and not (layer3_outputs(1436));
    layer4_outputs(2816) <= not(layer3_outputs(2416)) or (layer3_outputs(4705));
    layer4_outputs(2817) <= (layer3_outputs(1154)) or (layer3_outputs(889));
    layer4_outputs(2818) <= (layer3_outputs(1165)) xor (layer3_outputs(1124));
    layer4_outputs(2819) <= layer3_outputs(4821);
    layer4_outputs(2820) <= '1';
    layer4_outputs(2821) <= (layer3_outputs(5816)) or (layer3_outputs(1874));
    layer4_outputs(2822) <= not(layer3_outputs(3438));
    layer4_outputs(2823) <= (layer3_outputs(4463)) and not (layer3_outputs(6719));
    layer4_outputs(2824) <= layer3_outputs(2328);
    layer4_outputs(2825) <= not((layer3_outputs(4746)) xor (layer3_outputs(5701)));
    layer4_outputs(2826) <= not(layer3_outputs(605));
    layer4_outputs(2827) <= not((layer3_outputs(186)) or (layer3_outputs(3330)));
    layer4_outputs(2828) <= not(layer3_outputs(4016));
    layer4_outputs(2829) <= layer3_outputs(2810);
    layer4_outputs(2830) <= layer3_outputs(4982);
    layer4_outputs(2831) <= not(layer3_outputs(4994));
    layer4_outputs(2832) <= not(layer3_outputs(1447));
    layer4_outputs(2833) <= (layer3_outputs(6664)) and not (layer3_outputs(5175));
    layer4_outputs(2834) <= (layer3_outputs(4211)) and (layer3_outputs(7600));
    layer4_outputs(2835) <= not(layer3_outputs(3674));
    layer4_outputs(2836) <= not((layer3_outputs(214)) xor (layer3_outputs(7391)));
    layer4_outputs(2837) <= not(layer3_outputs(1004));
    layer4_outputs(2838) <= not((layer3_outputs(3271)) and (layer3_outputs(4586)));
    layer4_outputs(2839) <= not((layer3_outputs(5568)) xor (layer3_outputs(4270)));
    layer4_outputs(2840) <= not(layer3_outputs(251));
    layer4_outputs(2841) <= not(layer3_outputs(4958));
    layer4_outputs(2842) <= layer3_outputs(6377);
    layer4_outputs(2843) <= layer3_outputs(6316);
    layer4_outputs(2844) <= not((layer3_outputs(3717)) or (layer3_outputs(7365)));
    layer4_outputs(2845) <= not((layer3_outputs(4090)) and (layer3_outputs(2858)));
    layer4_outputs(2846) <= (layer3_outputs(1390)) and not (layer3_outputs(3969));
    layer4_outputs(2847) <= layer3_outputs(983);
    layer4_outputs(2848) <= (layer3_outputs(2809)) and not (layer3_outputs(6453));
    layer4_outputs(2849) <= not(layer3_outputs(1571));
    layer4_outputs(2850) <= layer3_outputs(5220);
    layer4_outputs(2851) <= layer3_outputs(3469);
    layer4_outputs(2852) <= layer3_outputs(621);
    layer4_outputs(2853) <= (layer3_outputs(4261)) xor (layer3_outputs(5845));
    layer4_outputs(2854) <= not(layer3_outputs(3143)) or (layer3_outputs(1288));
    layer4_outputs(2855) <= not(layer3_outputs(3240));
    layer4_outputs(2856) <= (layer3_outputs(1085)) or (layer3_outputs(3449));
    layer4_outputs(2857) <= (layer3_outputs(4506)) and not (layer3_outputs(1089));
    layer4_outputs(2858) <= layer3_outputs(754);
    layer4_outputs(2859) <= (layer3_outputs(6752)) or (layer3_outputs(5371));
    layer4_outputs(2860) <= not(layer3_outputs(4648));
    layer4_outputs(2861) <= not(layer3_outputs(2871));
    layer4_outputs(2862) <= not((layer3_outputs(1502)) or (layer3_outputs(1)));
    layer4_outputs(2863) <= not(layer3_outputs(2389)) or (layer3_outputs(3215));
    layer4_outputs(2864) <= not(layer3_outputs(6022));
    layer4_outputs(2865) <= (layer3_outputs(6412)) and (layer3_outputs(6365));
    layer4_outputs(2866) <= not(layer3_outputs(4657)) or (layer3_outputs(3128));
    layer4_outputs(2867) <= layer3_outputs(1365);
    layer4_outputs(2868) <= '1';
    layer4_outputs(2869) <= layer3_outputs(792);
    layer4_outputs(2870) <= layer3_outputs(798);
    layer4_outputs(2871) <= not((layer3_outputs(6146)) or (layer3_outputs(5800)));
    layer4_outputs(2872) <= layer3_outputs(7155);
    layer4_outputs(2873) <= not(layer3_outputs(7141));
    layer4_outputs(2874) <= not(layer3_outputs(1612));
    layer4_outputs(2875) <= layer3_outputs(5643);
    layer4_outputs(2876) <= layer3_outputs(4986);
    layer4_outputs(2877) <= layer3_outputs(4572);
    layer4_outputs(2878) <= not((layer3_outputs(4092)) or (layer3_outputs(3800)));
    layer4_outputs(2879) <= not(layer3_outputs(6305));
    layer4_outputs(2880) <= layer3_outputs(6581);
    layer4_outputs(2881) <= layer3_outputs(6927);
    layer4_outputs(2882) <= layer3_outputs(7076);
    layer4_outputs(2883) <= not((layer3_outputs(3125)) xor (layer3_outputs(4409)));
    layer4_outputs(2884) <= layer3_outputs(4479);
    layer4_outputs(2885) <= not(layer3_outputs(4637));
    layer4_outputs(2886) <= not((layer3_outputs(3348)) and (layer3_outputs(5904)));
    layer4_outputs(2887) <= (layer3_outputs(2657)) xor (layer3_outputs(5638));
    layer4_outputs(2888) <= (layer3_outputs(4552)) and not (layer3_outputs(4858));
    layer4_outputs(2889) <= (layer3_outputs(2185)) or (layer3_outputs(5995));
    layer4_outputs(2890) <= not((layer3_outputs(3202)) or (layer3_outputs(6772)));
    layer4_outputs(2891) <= not((layer3_outputs(3215)) xor (layer3_outputs(7522)));
    layer4_outputs(2892) <= layer3_outputs(1626);
    layer4_outputs(2893) <= not(layer3_outputs(7054));
    layer4_outputs(2894) <= (layer3_outputs(6497)) xor (layer3_outputs(6635));
    layer4_outputs(2895) <= not(layer3_outputs(6566));
    layer4_outputs(2896) <= layer3_outputs(3402);
    layer4_outputs(2897) <= not(layer3_outputs(5353));
    layer4_outputs(2898) <= layer3_outputs(1212);
    layer4_outputs(2899) <= layer3_outputs(6894);
    layer4_outputs(2900) <= (layer3_outputs(3556)) and not (layer3_outputs(3112));
    layer4_outputs(2901) <= not(layer3_outputs(1950));
    layer4_outputs(2902) <= (layer3_outputs(765)) and not (layer3_outputs(7084));
    layer4_outputs(2903) <= layer3_outputs(6600);
    layer4_outputs(2904) <= not(layer3_outputs(4514));
    layer4_outputs(2905) <= (layer3_outputs(1382)) and not (layer3_outputs(1665));
    layer4_outputs(2906) <= not((layer3_outputs(6814)) xor (layer3_outputs(4100)));
    layer4_outputs(2907) <= layer3_outputs(4359);
    layer4_outputs(2908) <= layer3_outputs(6892);
    layer4_outputs(2909) <= layer3_outputs(3761);
    layer4_outputs(2910) <= (layer3_outputs(4255)) xor (layer3_outputs(3228));
    layer4_outputs(2911) <= (layer3_outputs(3270)) xor (layer3_outputs(534));
    layer4_outputs(2912) <= layer3_outputs(4061);
    layer4_outputs(2913) <= not(layer3_outputs(4331));
    layer4_outputs(2914) <= not(layer3_outputs(1559));
    layer4_outputs(2915) <= (layer3_outputs(5490)) or (layer3_outputs(2991));
    layer4_outputs(2916) <= layer3_outputs(4094);
    layer4_outputs(2917) <= layer3_outputs(1264);
    layer4_outputs(2918) <= not(layer3_outputs(7406));
    layer4_outputs(2919) <= not(layer3_outputs(2549));
    layer4_outputs(2920) <= layer3_outputs(1693);
    layer4_outputs(2921) <= (layer3_outputs(979)) and not (layer3_outputs(2359));
    layer4_outputs(2922) <= not((layer3_outputs(4256)) xor (layer3_outputs(3108)));
    layer4_outputs(2923) <= layer3_outputs(992);
    layer4_outputs(2924) <= layer3_outputs(4437);
    layer4_outputs(2925) <= (layer3_outputs(4946)) or (layer3_outputs(4779));
    layer4_outputs(2926) <= layer3_outputs(1819);
    layer4_outputs(2927) <= (layer3_outputs(3465)) and not (layer3_outputs(7289));
    layer4_outputs(2928) <= not((layer3_outputs(7297)) xor (layer3_outputs(5017)));
    layer4_outputs(2929) <= not(layer3_outputs(3182));
    layer4_outputs(2930) <= not((layer3_outputs(5344)) and (layer3_outputs(4967)));
    layer4_outputs(2931) <= (layer3_outputs(2046)) or (layer3_outputs(3221));
    layer4_outputs(2932) <= (layer3_outputs(5444)) and not (layer3_outputs(1071));
    layer4_outputs(2933) <= (layer3_outputs(4117)) and not (layer3_outputs(4487));
    layer4_outputs(2934) <= not(layer3_outputs(2758));
    layer4_outputs(2935) <= not((layer3_outputs(2874)) and (layer3_outputs(5773)));
    layer4_outputs(2936) <= not(layer3_outputs(4453));
    layer4_outputs(2937) <= not(layer3_outputs(7623));
    layer4_outputs(2938) <= (layer3_outputs(5089)) xor (layer3_outputs(2807));
    layer4_outputs(2939) <= not(layer3_outputs(5276)) or (layer3_outputs(6096));
    layer4_outputs(2940) <= (layer3_outputs(4301)) and (layer3_outputs(3061));
    layer4_outputs(2941) <= (layer3_outputs(3684)) and not (layer3_outputs(6181));
    layer4_outputs(2942) <= layer3_outputs(641);
    layer4_outputs(2943) <= not(layer3_outputs(5177));
    layer4_outputs(2944) <= (layer3_outputs(6701)) and not (layer3_outputs(3335));
    layer4_outputs(2945) <= not(layer3_outputs(3877)) or (layer3_outputs(2342));
    layer4_outputs(2946) <= layer3_outputs(1629);
    layer4_outputs(2947) <= not(layer3_outputs(716));
    layer4_outputs(2948) <= not(layer3_outputs(5757));
    layer4_outputs(2949) <= not((layer3_outputs(6449)) or (layer3_outputs(4354)));
    layer4_outputs(2950) <= layer3_outputs(3217);
    layer4_outputs(2951) <= layer3_outputs(6037);
    layer4_outputs(2952) <= not((layer3_outputs(6352)) xor (layer3_outputs(2976)));
    layer4_outputs(2953) <= (layer3_outputs(3054)) xor (layer3_outputs(2552));
    layer4_outputs(2954) <= (layer3_outputs(3951)) and not (layer3_outputs(7433));
    layer4_outputs(2955) <= not(layer3_outputs(7419));
    layer4_outputs(2956) <= not(layer3_outputs(7257));
    layer4_outputs(2957) <= not(layer3_outputs(3868));
    layer4_outputs(2958) <= not(layer3_outputs(852));
    layer4_outputs(2959) <= (layer3_outputs(7566)) xor (layer3_outputs(5317));
    layer4_outputs(2960) <= (layer3_outputs(5111)) and not (layer3_outputs(430));
    layer4_outputs(2961) <= not(layer3_outputs(1115));
    layer4_outputs(2962) <= not(layer3_outputs(3337));
    layer4_outputs(2963) <= not(layer3_outputs(6763));
    layer4_outputs(2964) <= layer3_outputs(2215);
    layer4_outputs(2965) <= layer3_outputs(4780);
    layer4_outputs(2966) <= not((layer3_outputs(2364)) or (layer3_outputs(1872)));
    layer4_outputs(2967) <= layer3_outputs(7445);
    layer4_outputs(2968) <= not(layer3_outputs(4942));
    layer4_outputs(2969) <= (layer3_outputs(7323)) or (layer3_outputs(5983));
    layer4_outputs(2970) <= (layer3_outputs(5558)) xor (layer3_outputs(4233));
    layer4_outputs(2971) <= layer3_outputs(539);
    layer4_outputs(2972) <= not(layer3_outputs(5835)) or (layer3_outputs(2211));
    layer4_outputs(2973) <= not(layer3_outputs(2796));
    layer4_outputs(2974) <= not(layer3_outputs(2022));
    layer4_outputs(2975) <= layer3_outputs(4535);
    layer4_outputs(2976) <= not(layer3_outputs(1860));
    layer4_outputs(2977) <= not((layer3_outputs(120)) and (layer3_outputs(1163)));
    layer4_outputs(2978) <= (layer3_outputs(571)) xor (layer3_outputs(1012));
    layer4_outputs(2979) <= (layer3_outputs(1421)) or (layer3_outputs(5264));
    layer4_outputs(2980) <= (layer3_outputs(7633)) or (layer3_outputs(5225));
    layer4_outputs(2981) <= not((layer3_outputs(6414)) or (layer3_outputs(7179)));
    layer4_outputs(2982) <= not(layer3_outputs(1274));
    layer4_outputs(2983) <= not((layer3_outputs(4594)) and (layer3_outputs(6800)));
    layer4_outputs(2984) <= layer3_outputs(1826);
    layer4_outputs(2985) <= not(layer3_outputs(1779));
    layer4_outputs(2986) <= (layer3_outputs(5020)) xor (layer3_outputs(3762));
    layer4_outputs(2987) <= not(layer3_outputs(438));
    layer4_outputs(2988) <= layer3_outputs(7450);
    layer4_outputs(2989) <= not(layer3_outputs(4950)) or (layer3_outputs(6652));
    layer4_outputs(2990) <= layer3_outputs(103);
    layer4_outputs(2991) <= not((layer3_outputs(301)) or (layer3_outputs(3981)));
    layer4_outputs(2992) <= not((layer3_outputs(4232)) and (layer3_outputs(449)));
    layer4_outputs(2993) <= not(layer3_outputs(1658)) or (layer3_outputs(4574));
    layer4_outputs(2994) <= not((layer3_outputs(2963)) xor (layer3_outputs(2098)));
    layer4_outputs(2995) <= layer3_outputs(6199);
    layer4_outputs(2996) <= not(layer3_outputs(4581));
    layer4_outputs(2997) <= (layer3_outputs(2351)) xor (layer3_outputs(7332));
    layer4_outputs(2998) <= not(layer3_outputs(6626));
    layer4_outputs(2999) <= (layer3_outputs(6053)) xor (layer3_outputs(405));
    layer4_outputs(3000) <= (layer3_outputs(1844)) xor (layer3_outputs(6520));
    layer4_outputs(3001) <= not(layer3_outputs(5247));
    layer4_outputs(3002) <= not(layer3_outputs(7468));
    layer4_outputs(3003) <= not(layer3_outputs(218));
    layer4_outputs(3004) <= not((layer3_outputs(7369)) xor (layer3_outputs(1610)));
    layer4_outputs(3005) <= layer3_outputs(4196);
    layer4_outputs(3006) <= layer3_outputs(3292);
    layer4_outputs(3007) <= not(layer3_outputs(1947));
    layer4_outputs(3008) <= layer3_outputs(6235);
    layer4_outputs(3009) <= (layer3_outputs(3957)) and not (layer3_outputs(396));
    layer4_outputs(3010) <= not((layer3_outputs(1156)) and (layer3_outputs(545)));
    layer4_outputs(3011) <= (layer3_outputs(5683)) and not (layer3_outputs(1922));
    layer4_outputs(3012) <= layer3_outputs(6376);
    layer4_outputs(3013) <= layer3_outputs(3518);
    layer4_outputs(3014) <= layer3_outputs(667);
    layer4_outputs(3015) <= not(layer3_outputs(4896)) or (layer3_outputs(3703));
    layer4_outputs(3016) <= (layer3_outputs(4704)) or (layer3_outputs(295));
    layer4_outputs(3017) <= (layer3_outputs(409)) xor (layer3_outputs(1654));
    layer4_outputs(3018) <= not(layer3_outputs(5712));
    layer4_outputs(3019) <= not(layer3_outputs(3336));
    layer4_outputs(3020) <= layer3_outputs(1760);
    layer4_outputs(3021) <= not(layer3_outputs(2038));
    layer4_outputs(3022) <= not((layer3_outputs(472)) and (layer3_outputs(5594)));
    layer4_outputs(3023) <= not(layer3_outputs(3388));
    layer4_outputs(3024) <= (layer3_outputs(624)) or (layer3_outputs(4598));
    layer4_outputs(3025) <= not(layer3_outputs(2519)) or (layer3_outputs(5195));
    layer4_outputs(3026) <= not((layer3_outputs(5415)) or (layer3_outputs(466)));
    layer4_outputs(3027) <= not((layer3_outputs(1261)) xor (layer3_outputs(3035)));
    layer4_outputs(3028) <= (layer3_outputs(3646)) and (layer3_outputs(389));
    layer4_outputs(3029) <= not(layer3_outputs(7134));
    layer4_outputs(3030) <= not((layer3_outputs(2626)) and (layer3_outputs(3830)));
    layer4_outputs(3031) <= not(layer3_outputs(2983));
    layer4_outputs(3032) <= (layer3_outputs(234)) and not (layer3_outputs(3750));
    layer4_outputs(3033) <= (layer3_outputs(2639)) or (layer3_outputs(4519));
    layer4_outputs(3034) <= layer3_outputs(3578);
    layer4_outputs(3035) <= not((layer3_outputs(4382)) xor (layer3_outputs(7257)));
    layer4_outputs(3036) <= not(layer3_outputs(196)) or (layer3_outputs(4193));
    layer4_outputs(3037) <= layer3_outputs(522);
    layer4_outputs(3038) <= (layer3_outputs(29)) xor (layer3_outputs(6773));
    layer4_outputs(3039) <= (layer3_outputs(5653)) or (layer3_outputs(7026));
    layer4_outputs(3040) <= layer3_outputs(2607);
    layer4_outputs(3041) <= (layer3_outputs(5054)) and not (layer3_outputs(27));
    layer4_outputs(3042) <= not((layer3_outputs(2205)) or (layer3_outputs(2546)));
    layer4_outputs(3043) <= not(layer3_outputs(1064)) or (layer3_outputs(3218));
    layer4_outputs(3044) <= (layer3_outputs(953)) and not (layer3_outputs(7513));
    layer4_outputs(3045) <= not(layer3_outputs(6289));
    layer4_outputs(3046) <= not(layer3_outputs(3818));
    layer4_outputs(3047) <= layer3_outputs(3339);
    layer4_outputs(3048) <= not((layer3_outputs(3370)) xor (layer3_outputs(5102)));
    layer4_outputs(3049) <= not(layer3_outputs(5616));
    layer4_outputs(3050) <= not(layer3_outputs(3574));
    layer4_outputs(3051) <= (layer3_outputs(520)) xor (layer3_outputs(5357));
    layer4_outputs(3052) <= layer3_outputs(1335);
    layer4_outputs(3053) <= (layer3_outputs(4113)) or (layer3_outputs(3041));
    layer4_outputs(3054) <= layer3_outputs(1035);
    layer4_outputs(3055) <= not(layer3_outputs(6420));
    layer4_outputs(3056) <= not(layer3_outputs(4429)) or (layer3_outputs(7470));
    layer4_outputs(3057) <= not(layer3_outputs(2023)) or (layer3_outputs(6313));
    layer4_outputs(3058) <= not(layer3_outputs(5589)) or (layer3_outputs(2169));
    layer4_outputs(3059) <= not(layer3_outputs(850));
    layer4_outputs(3060) <= layer3_outputs(7346);
    layer4_outputs(3061) <= layer3_outputs(1613);
    layer4_outputs(3062) <= not(layer3_outputs(2756)) or (layer3_outputs(7084));
    layer4_outputs(3063) <= not(layer3_outputs(2346));
    layer4_outputs(3064) <= layer3_outputs(3903);
    layer4_outputs(3065) <= layer3_outputs(6091);
    layer4_outputs(3066) <= not(layer3_outputs(2146)) or (layer3_outputs(4192));
    layer4_outputs(3067) <= not(layer3_outputs(1677)) or (layer3_outputs(3520));
    layer4_outputs(3068) <= layer3_outputs(6732);
    layer4_outputs(3069) <= not((layer3_outputs(5575)) and (layer3_outputs(5144)));
    layer4_outputs(3070) <= not((layer3_outputs(5241)) xor (layer3_outputs(6325)));
    layer4_outputs(3071) <= (layer3_outputs(5476)) and not (layer3_outputs(2000));
    layer4_outputs(3072) <= layer3_outputs(6298);
    layer4_outputs(3073) <= layer3_outputs(4899);
    layer4_outputs(3074) <= not(layer3_outputs(1912));
    layer4_outputs(3075) <= (layer3_outputs(2140)) and not (layer3_outputs(6292));
    layer4_outputs(3076) <= not(layer3_outputs(7042)) or (layer3_outputs(2665));
    layer4_outputs(3077) <= layer3_outputs(3139);
    layer4_outputs(3078) <= (layer3_outputs(6564)) and (layer3_outputs(3663));
    layer4_outputs(3079) <= layer3_outputs(3556);
    layer4_outputs(3080) <= not(layer3_outputs(5392));
    layer4_outputs(3081) <= (layer3_outputs(7064)) xor (layer3_outputs(4505));
    layer4_outputs(3082) <= (layer3_outputs(800)) and not (layer3_outputs(3537));
    layer4_outputs(3083) <= not((layer3_outputs(2622)) and (layer3_outputs(5065)));
    layer4_outputs(3084) <= not(layer3_outputs(4320));
    layer4_outputs(3085) <= not(layer3_outputs(759));
    layer4_outputs(3086) <= not(layer3_outputs(803));
    layer4_outputs(3087) <= layer3_outputs(4392);
    layer4_outputs(3088) <= (layer3_outputs(3499)) and not (layer3_outputs(4741));
    layer4_outputs(3089) <= (layer3_outputs(2592)) xor (layer3_outputs(690));
    layer4_outputs(3090) <= not((layer3_outputs(2035)) or (layer3_outputs(5922)));
    layer4_outputs(3091) <= layer3_outputs(3550);
    layer4_outputs(3092) <= not((layer3_outputs(5624)) or (layer3_outputs(2691)));
    layer4_outputs(3093) <= not(layer3_outputs(2919));
    layer4_outputs(3094) <= not(layer3_outputs(5919));
    layer4_outputs(3095) <= not((layer3_outputs(2281)) or (layer3_outputs(1403)));
    layer4_outputs(3096) <= not((layer3_outputs(4874)) and (layer3_outputs(5654)));
    layer4_outputs(3097) <= not(layer3_outputs(1802)) or (layer3_outputs(807));
    layer4_outputs(3098) <= not(layer3_outputs(5758)) or (layer3_outputs(428));
    layer4_outputs(3099) <= not(layer3_outputs(6709));
    layer4_outputs(3100) <= layer3_outputs(811);
    layer4_outputs(3101) <= not(layer3_outputs(3998));
    layer4_outputs(3102) <= not(layer3_outputs(6838));
    layer4_outputs(3103) <= not((layer3_outputs(2971)) and (layer3_outputs(7233)));
    layer4_outputs(3104) <= not(layer3_outputs(2097)) or (layer3_outputs(1103));
    layer4_outputs(3105) <= not((layer3_outputs(4249)) or (layer3_outputs(3504)));
    layer4_outputs(3106) <= layer3_outputs(2421);
    layer4_outputs(3107) <= not(layer3_outputs(7202));
    layer4_outputs(3108) <= layer3_outputs(4499);
    layer4_outputs(3109) <= (layer3_outputs(1642)) or (layer3_outputs(3382));
    layer4_outputs(3110) <= not((layer3_outputs(5490)) and (layer3_outputs(4719)));
    layer4_outputs(3111) <= not(layer3_outputs(2223));
    layer4_outputs(3112) <= not(layer3_outputs(5231)) or (layer3_outputs(1916));
    layer4_outputs(3113) <= (layer3_outputs(1617)) or (layer3_outputs(2579));
    layer4_outputs(3114) <= layer3_outputs(3277);
    layer4_outputs(3115) <= not(layer3_outputs(3061));
    layer4_outputs(3116) <= layer3_outputs(4327);
    layer4_outputs(3117) <= (layer3_outputs(2853)) xor (layer3_outputs(6211));
    layer4_outputs(3118) <= (layer3_outputs(4157)) and not (layer3_outputs(2688));
    layer4_outputs(3119) <= layer3_outputs(3431);
    layer4_outputs(3120) <= layer3_outputs(718);
    layer4_outputs(3121) <= layer3_outputs(3656);
    layer4_outputs(3122) <= not(layer3_outputs(7651));
    layer4_outputs(3123) <= layer3_outputs(4828);
    layer4_outputs(3124) <= not(layer3_outputs(3026));
    layer4_outputs(3125) <= layer3_outputs(6550);
    layer4_outputs(3126) <= (layer3_outputs(5341)) and not (layer3_outputs(2959));
    layer4_outputs(3127) <= (layer3_outputs(5815)) and not (layer3_outputs(6347));
    layer4_outputs(3128) <= not(layer3_outputs(2114));
    layer4_outputs(3129) <= (layer3_outputs(4582)) or (layer3_outputs(2698));
    layer4_outputs(3130) <= (layer3_outputs(6871)) and (layer3_outputs(2613));
    layer4_outputs(3131) <= (layer3_outputs(7357)) or (layer3_outputs(6794));
    layer4_outputs(3132) <= (layer3_outputs(1248)) xor (layer3_outputs(616));
    layer4_outputs(3133) <= not((layer3_outputs(7002)) xor (layer3_outputs(2334)));
    layer4_outputs(3134) <= (layer3_outputs(827)) and (layer3_outputs(7424));
    layer4_outputs(3135) <= not(layer3_outputs(7649)) or (layer3_outputs(1031));
    layer4_outputs(3136) <= not((layer3_outputs(7647)) and (layer3_outputs(1715)));
    layer4_outputs(3137) <= layer3_outputs(2696);
    layer4_outputs(3138) <= layer3_outputs(3447);
    layer4_outputs(3139) <= layer3_outputs(656);
    layer4_outputs(3140) <= '0';
    layer4_outputs(3141) <= layer3_outputs(2293);
    layer4_outputs(3142) <= not(layer3_outputs(3881)) or (layer3_outputs(3610));
    layer4_outputs(3143) <= not(layer3_outputs(1192));
    layer4_outputs(3144) <= (layer3_outputs(4910)) and not (layer3_outputs(5158));
    layer4_outputs(3145) <= not(layer3_outputs(5727));
    layer4_outputs(3146) <= not(layer3_outputs(1634)) or (layer3_outputs(5188));
    layer4_outputs(3147) <= not(layer3_outputs(7086));
    layer4_outputs(3148) <= not(layer3_outputs(2031));
    layer4_outputs(3149) <= (layer3_outputs(2993)) and not (layer3_outputs(615));
    layer4_outputs(3150) <= layer3_outputs(5174);
    layer4_outputs(3151) <= not(layer3_outputs(5554));
    layer4_outputs(3152) <= (layer3_outputs(6971)) and (layer3_outputs(761));
    layer4_outputs(3153) <= not(layer3_outputs(200));
    layer4_outputs(3154) <= not(layer3_outputs(997));
    layer4_outputs(3155) <= not((layer3_outputs(402)) xor (layer3_outputs(4274)));
    layer4_outputs(3156) <= not(layer3_outputs(4783));
    layer4_outputs(3157) <= (layer3_outputs(2649)) xor (layer3_outputs(7307));
    layer4_outputs(3158) <= layer3_outputs(6189);
    layer4_outputs(3159) <= (layer3_outputs(5736)) and not (layer3_outputs(5172));
    layer4_outputs(3160) <= '0';
    layer4_outputs(3161) <= layer3_outputs(5620);
    layer4_outputs(3162) <= not(layer3_outputs(7368));
    layer4_outputs(3163) <= not((layer3_outputs(1413)) xor (layer3_outputs(6504)));
    layer4_outputs(3164) <= (layer3_outputs(2164)) xor (layer3_outputs(1989));
    layer4_outputs(3165) <= (layer3_outputs(1336)) or (layer3_outputs(4523));
    layer4_outputs(3166) <= (layer3_outputs(3753)) and not (layer3_outputs(2805));
    layer4_outputs(3167) <= layer3_outputs(5505);
    layer4_outputs(3168) <= layer3_outputs(4839);
    layer4_outputs(3169) <= layer3_outputs(3328);
    layer4_outputs(3170) <= not(layer3_outputs(917)) or (layer3_outputs(7259));
    layer4_outputs(3171) <= layer3_outputs(1731);
    layer4_outputs(3172) <= not((layer3_outputs(1898)) or (layer3_outputs(2877)));
    layer4_outputs(3173) <= (layer3_outputs(293)) xor (layer3_outputs(4252));
    layer4_outputs(3174) <= layer3_outputs(3460);
    layer4_outputs(3175) <= not(layer3_outputs(7208));
    layer4_outputs(3176) <= (layer3_outputs(1577)) xor (layer3_outputs(902));
    layer4_outputs(3177) <= not(layer3_outputs(2535));
    layer4_outputs(3178) <= not(layer3_outputs(222));
    layer4_outputs(3179) <= (layer3_outputs(726)) and not (layer3_outputs(168));
    layer4_outputs(3180) <= (layer3_outputs(408)) and not (layer3_outputs(4753));
    layer4_outputs(3181) <= not(layer3_outputs(3677));
    layer4_outputs(3182) <= not((layer3_outputs(101)) or (layer3_outputs(4607)));
    layer4_outputs(3183) <= not(layer3_outputs(3982));
    layer4_outputs(3184) <= not((layer3_outputs(5822)) or (layer3_outputs(6036)));
    layer4_outputs(3185) <= (layer3_outputs(6534)) and (layer3_outputs(6666));
    layer4_outputs(3186) <= not(layer3_outputs(7537));
    layer4_outputs(3187) <= layer3_outputs(3142);
    layer4_outputs(3188) <= (layer3_outputs(264)) or (layer3_outputs(3697));
    layer4_outputs(3189) <= (layer3_outputs(4844)) and not (layer3_outputs(4222));
    layer4_outputs(3190) <= layer3_outputs(407);
    layer4_outputs(3191) <= (layer3_outputs(5491)) and (layer3_outputs(6140));
    layer4_outputs(3192) <= layer3_outputs(7615);
    layer4_outputs(3193) <= not((layer3_outputs(1574)) or (layer3_outputs(2306)));
    layer4_outputs(3194) <= not(layer3_outputs(4591)) or (layer3_outputs(83));
    layer4_outputs(3195) <= (layer3_outputs(4032)) or (layer3_outputs(2949));
    layer4_outputs(3196) <= (layer3_outputs(1757)) and not (layer3_outputs(5134));
    layer4_outputs(3197) <= layer3_outputs(5894);
    layer4_outputs(3198) <= not((layer3_outputs(4688)) and (layer3_outputs(3803)));
    layer4_outputs(3199) <= not(layer3_outputs(6573));
    layer4_outputs(3200) <= layer3_outputs(4539);
    layer4_outputs(3201) <= layer3_outputs(2693);
    layer4_outputs(3202) <= layer3_outputs(1915);
    layer4_outputs(3203) <= (layer3_outputs(3862)) and not (layer3_outputs(40));
    layer4_outputs(3204) <= layer3_outputs(2519);
    layer4_outputs(3205) <= not(layer3_outputs(1613));
    layer4_outputs(3206) <= not(layer3_outputs(1485));
    layer4_outputs(3207) <= (layer3_outputs(6765)) and not (layer3_outputs(3892));
    layer4_outputs(3208) <= layer3_outputs(6624);
    layer4_outputs(3209) <= (layer3_outputs(3809)) and not (layer3_outputs(407));
    layer4_outputs(3210) <= not((layer3_outputs(4928)) or (layer3_outputs(2600)));
    layer4_outputs(3211) <= (layer3_outputs(1959)) and not (layer3_outputs(7653));
    layer4_outputs(3212) <= not(layer3_outputs(4191));
    layer4_outputs(3213) <= not(layer3_outputs(3686)) or (layer3_outputs(7067));
    layer4_outputs(3214) <= not((layer3_outputs(1842)) xor (layer3_outputs(6321)));
    layer4_outputs(3215) <= layer3_outputs(2634);
    layer4_outputs(3216) <= layer3_outputs(4946);
    layer4_outputs(3217) <= (layer3_outputs(1941)) and (layer3_outputs(853));
    layer4_outputs(3218) <= not(layer3_outputs(6902));
    layer4_outputs(3219) <= (layer3_outputs(4627)) and (layer3_outputs(279));
    layer4_outputs(3220) <= layer3_outputs(6024);
    layer4_outputs(3221) <= (layer3_outputs(6483)) and (layer3_outputs(2439));
    layer4_outputs(3222) <= layer3_outputs(4735);
    layer4_outputs(3223) <= layer3_outputs(3808);
    layer4_outputs(3224) <= (layer3_outputs(2285)) and not (layer3_outputs(1526));
    layer4_outputs(3225) <= layer3_outputs(6268);
    layer4_outputs(3226) <= (layer3_outputs(5185)) or (layer3_outputs(6228));
    layer4_outputs(3227) <= not(layer3_outputs(239));
    layer4_outputs(3228) <= not((layer3_outputs(1324)) xor (layer3_outputs(6897)));
    layer4_outputs(3229) <= not(layer3_outputs(6333));
    layer4_outputs(3230) <= layer3_outputs(2125);
    layer4_outputs(3231) <= not(layer3_outputs(1624));
    layer4_outputs(3232) <= (layer3_outputs(2219)) or (layer3_outputs(3833));
    layer4_outputs(3233) <= (layer3_outputs(6297)) and (layer3_outputs(3576));
    layer4_outputs(3234) <= (layer3_outputs(2584)) and (layer3_outputs(5752));
    layer4_outputs(3235) <= not(layer3_outputs(2903));
    layer4_outputs(3236) <= (layer3_outputs(1966)) and not (layer3_outputs(1668));
    layer4_outputs(3237) <= not(layer3_outputs(7602)) or (layer3_outputs(1377));
    layer4_outputs(3238) <= not((layer3_outputs(1112)) xor (layer3_outputs(6379)));
    layer4_outputs(3239) <= not(layer3_outputs(4689)) or (layer3_outputs(4044));
    layer4_outputs(3240) <= layer3_outputs(5036);
    layer4_outputs(3241) <= not(layer3_outputs(5278));
    layer4_outputs(3242) <= (layer3_outputs(1143)) and (layer3_outputs(102));
    layer4_outputs(3243) <= not(layer3_outputs(1809)) or (layer3_outputs(7272));
    layer4_outputs(3244) <= not(layer3_outputs(1716));
    layer4_outputs(3245) <= layer3_outputs(1936);
    layer4_outputs(3246) <= layer3_outputs(3008);
    layer4_outputs(3247) <= (layer3_outputs(5066)) and (layer3_outputs(2677));
    layer4_outputs(3248) <= not((layer3_outputs(2890)) and (layer3_outputs(7059)));
    layer4_outputs(3249) <= layer3_outputs(7125);
    layer4_outputs(3250) <= not((layer3_outputs(6507)) xor (layer3_outputs(3952)));
    layer4_outputs(3251) <= layer3_outputs(7431);
    layer4_outputs(3252) <= not((layer3_outputs(7636)) or (layer3_outputs(1518)));
    layer4_outputs(3253) <= (layer3_outputs(6395)) xor (layer3_outputs(2329));
    layer4_outputs(3254) <= not(layer3_outputs(6816));
    layer4_outputs(3255) <= layer3_outputs(6319);
    layer4_outputs(3256) <= not(layer3_outputs(744));
    layer4_outputs(3257) <= (layer3_outputs(734)) or (layer3_outputs(5239));
    layer4_outputs(3258) <= not(layer3_outputs(5397));
    layer4_outputs(3259) <= not(layer3_outputs(2901));
    layer4_outputs(3260) <= (layer3_outputs(3835)) xor (layer3_outputs(5924));
    layer4_outputs(3261) <= (layer3_outputs(5078)) xor (layer3_outputs(3997));
    layer4_outputs(3262) <= not(layer3_outputs(7209));
    layer4_outputs(3263) <= layer3_outputs(3365);
    layer4_outputs(3264) <= layer3_outputs(1549);
    layer4_outputs(3265) <= not(layer3_outputs(1142)) or (layer3_outputs(4421));
    layer4_outputs(3266) <= not(layer3_outputs(2218));
    layer4_outputs(3267) <= (layer3_outputs(6570)) xor (layer3_outputs(6652));
    layer4_outputs(3268) <= layer3_outputs(3070);
    layer4_outputs(3269) <= not(layer3_outputs(7096));
    layer4_outputs(3270) <= not(layer3_outputs(89));
    layer4_outputs(3271) <= not(layer3_outputs(7630));
    layer4_outputs(3272) <= layer3_outputs(2340);
    layer4_outputs(3273) <= (layer3_outputs(5761)) and (layer3_outputs(6933));
    layer4_outputs(3274) <= layer3_outputs(1343);
    layer4_outputs(3275) <= layer3_outputs(1183);
    layer4_outputs(3276) <= layer3_outputs(6925);
    layer4_outputs(3277) <= not((layer3_outputs(41)) xor (layer3_outputs(4784)));
    layer4_outputs(3278) <= not((layer3_outputs(3604)) xor (layer3_outputs(833)));
    layer4_outputs(3279) <= not(layer3_outputs(156)) or (layer3_outputs(2415));
    layer4_outputs(3280) <= (layer3_outputs(5965)) and not (layer3_outputs(4979));
    layer4_outputs(3281) <= layer3_outputs(1588);
    layer4_outputs(3282) <= not(layer3_outputs(941));
    layer4_outputs(3283) <= not(layer3_outputs(6142));
    layer4_outputs(3284) <= (layer3_outputs(6112)) and not (layer3_outputs(3570));
    layer4_outputs(3285) <= (layer3_outputs(2887)) or (layer3_outputs(3620));
    layer4_outputs(3286) <= layer3_outputs(1692);
    layer4_outputs(3287) <= layer3_outputs(4975);
    layer4_outputs(3288) <= not(layer3_outputs(5826));
    layer4_outputs(3289) <= layer3_outputs(7516);
    layer4_outputs(3290) <= (layer3_outputs(1249)) and not (layer3_outputs(5481));
    layer4_outputs(3291) <= (layer3_outputs(2501)) or (layer3_outputs(4039));
    layer4_outputs(3292) <= not(layer3_outputs(5952));
    layer4_outputs(3293) <= (layer3_outputs(296)) xor (layer3_outputs(821));
    layer4_outputs(3294) <= layer3_outputs(2273);
    layer4_outputs(3295) <= not(layer3_outputs(4971));
    layer4_outputs(3296) <= not(layer3_outputs(846));
    layer4_outputs(3297) <= not(layer3_outputs(1772));
    layer4_outputs(3298) <= layer3_outputs(1370);
    layer4_outputs(3299) <= (layer3_outputs(3733)) and not (layer3_outputs(4122));
    layer4_outputs(3300) <= not((layer3_outputs(5376)) and (layer3_outputs(1391)));
    layer4_outputs(3301) <= layer3_outputs(1454);
    layer4_outputs(3302) <= (layer3_outputs(4706)) and (layer3_outputs(386));
    layer4_outputs(3303) <= (layer3_outputs(4909)) or (layer3_outputs(197));
    layer4_outputs(3304) <= (layer3_outputs(2133)) and (layer3_outputs(2754));
    layer4_outputs(3305) <= not(layer3_outputs(6398));
    layer4_outputs(3306) <= layer3_outputs(3141);
    layer4_outputs(3307) <= (layer3_outputs(4129)) or (layer3_outputs(7442));
    layer4_outputs(3308) <= not(layer3_outputs(5152)) or (layer3_outputs(4820));
    layer4_outputs(3309) <= layer3_outputs(4292);
    layer4_outputs(3310) <= (layer3_outputs(337)) and not (layer3_outputs(3643));
    layer4_outputs(3311) <= not((layer3_outputs(1456)) xor (layer3_outputs(4209)));
    layer4_outputs(3312) <= layer3_outputs(562);
    layer4_outputs(3313) <= not(layer3_outputs(4214));
    layer4_outputs(3314) <= (layer3_outputs(4609)) and (layer3_outputs(3972));
    layer4_outputs(3315) <= (layer3_outputs(5368)) and (layer3_outputs(3464));
    layer4_outputs(3316) <= layer3_outputs(1961);
    layer4_outputs(3317) <= (layer3_outputs(1854)) and not (layer3_outputs(4602));
    layer4_outputs(3318) <= (layer3_outputs(618)) and not (layer3_outputs(925));
    layer4_outputs(3319) <= not(layer3_outputs(5134));
    layer4_outputs(3320) <= (layer3_outputs(3307)) and (layer3_outputs(3839));
    layer4_outputs(3321) <= not(layer3_outputs(7075));
    layer4_outputs(3322) <= not(layer3_outputs(11));
    layer4_outputs(3323) <= (layer3_outputs(5041)) or (layer3_outputs(6039));
    layer4_outputs(3324) <= not(layer3_outputs(385));
    layer4_outputs(3325) <= layer3_outputs(6148);
    layer4_outputs(3326) <= (layer3_outputs(5808)) xor (layer3_outputs(5112));
    layer4_outputs(3327) <= not(layer3_outputs(6143)) or (layer3_outputs(732));
    layer4_outputs(3328) <= not(layer3_outputs(3059));
    layer4_outputs(3329) <= (layer3_outputs(5672)) and not (layer3_outputs(3569));
    layer4_outputs(3330) <= layer3_outputs(6744);
    layer4_outputs(3331) <= (layer3_outputs(5240)) and not (layer3_outputs(7300));
    layer4_outputs(3332) <= (layer3_outputs(6508)) and not (layer3_outputs(832));
    layer4_outputs(3333) <= (layer3_outputs(1281)) and (layer3_outputs(6706));
    layer4_outputs(3334) <= '0';
    layer4_outputs(3335) <= not(layer3_outputs(81)) or (layer3_outputs(6969));
    layer4_outputs(3336) <= layer3_outputs(1564);
    layer4_outputs(3337) <= (layer3_outputs(6769)) xor (layer3_outputs(4226));
    layer4_outputs(3338) <= not((layer3_outputs(3425)) and (layer3_outputs(1954)));
    layer4_outputs(3339) <= layer3_outputs(5926);
    layer4_outputs(3340) <= (layer3_outputs(5655)) xor (layer3_outputs(1355));
    layer4_outputs(3341) <= layer3_outputs(4934);
    layer4_outputs(3342) <= not(layer3_outputs(3383));
    layer4_outputs(3343) <= (layer3_outputs(7306)) or (layer3_outputs(7549));
    layer4_outputs(3344) <= layer3_outputs(5637);
    layer4_outputs(3345) <= layer3_outputs(442);
    layer4_outputs(3346) <= layer3_outputs(545);
    layer4_outputs(3347) <= not(layer3_outputs(3267));
    layer4_outputs(3348) <= (layer3_outputs(1120)) and not (layer3_outputs(930));
    layer4_outputs(3349) <= layer3_outputs(680);
    layer4_outputs(3350) <= not((layer3_outputs(6710)) or (layer3_outputs(3614)));
    layer4_outputs(3351) <= not(layer3_outputs(3936)) or (layer3_outputs(3698));
    layer4_outputs(3352) <= (layer3_outputs(6080)) and not (layer3_outputs(2496));
    layer4_outputs(3353) <= not(layer3_outputs(6940));
    layer4_outputs(3354) <= not(layer3_outputs(2130));
    layer4_outputs(3355) <= not(layer3_outputs(6071)) or (layer3_outputs(3922));
    layer4_outputs(3356) <= layer3_outputs(317);
    layer4_outputs(3357) <= (layer3_outputs(4872)) or (layer3_outputs(1929));
    layer4_outputs(3358) <= not(layer3_outputs(6141)) or (layer3_outputs(1297));
    layer4_outputs(3359) <= not(layer3_outputs(5015));
    layer4_outputs(3360) <= layer3_outputs(3353);
    layer4_outputs(3361) <= layer3_outputs(744);
    layer4_outputs(3362) <= layer3_outputs(3532);
    layer4_outputs(3363) <= not(layer3_outputs(7362));
    layer4_outputs(3364) <= layer3_outputs(5332);
    layer4_outputs(3365) <= '1';
    layer4_outputs(3366) <= layer3_outputs(5686);
    layer4_outputs(3367) <= not(layer3_outputs(1176));
    layer4_outputs(3368) <= not(layer3_outputs(4756)) or (layer3_outputs(4667));
    layer4_outputs(3369) <= not(layer3_outputs(2392));
    layer4_outputs(3370) <= not(layer3_outputs(1437)) or (layer3_outputs(5286));
    layer4_outputs(3371) <= not(layer3_outputs(4845));
    layer4_outputs(3372) <= not((layer3_outputs(2618)) and (layer3_outputs(3364)));
    layer4_outputs(3373) <= not(layer3_outputs(6526));
    layer4_outputs(3374) <= not((layer3_outputs(5004)) and (layer3_outputs(6588)));
    layer4_outputs(3375) <= (layer3_outputs(1808)) and not (layer3_outputs(3737));
    layer4_outputs(3376) <= not(layer3_outputs(1150));
    layer4_outputs(3377) <= not(layer3_outputs(1400)) or (layer3_outputs(4721));
    layer4_outputs(3378) <= layer3_outputs(1517);
    layer4_outputs(3379) <= (layer3_outputs(1981)) and not (layer3_outputs(1497));
    layer4_outputs(3380) <= (layer3_outputs(2020)) and (layer3_outputs(2567));
    layer4_outputs(3381) <= layer3_outputs(5379);
    layer4_outputs(3382) <= layer3_outputs(5736);
    layer4_outputs(3383) <= layer3_outputs(4239);
    layer4_outputs(3384) <= not(layer3_outputs(161));
    layer4_outputs(3385) <= layer3_outputs(4925);
    layer4_outputs(3386) <= (layer3_outputs(3785)) and (layer3_outputs(393));
    layer4_outputs(3387) <= not((layer3_outputs(6423)) and (layer3_outputs(5663)));
    layer4_outputs(3388) <= layer3_outputs(1924);
    layer4_outputs(3389) <= '0';
    layer4_outputs(3390) <= not(layer3_outputs(147));
    layer4_outputs(3391) <= layer3_outputs(826);
    layer4_outputs(3392) <= not((layer3_outputs(3839)) and (layer3_outputs(4852)));
    layer4_outputs(3393) <= not(layer3_outputs(6992));
    layer4_outputs(3394) <= not(layer3_outputs(937));
    layer4_outputs(3395) <= layer3_outputs(6498);
    layer4_outputs(3396) <= (layer3_outputs(3495)) or (layer3_outputs(45));
    layer4_outputs(3397) <= not(layer3_outputs(1918));
    layer4_outputs(3398) <= not(layer3_outputs(7123));
    layer4_outputs(3399) <= not(layer3_outputs(3483)) or (layer3_outputs(5151));
    layer4_outputs(3400) <= layer3_outputs(5536);
    layer4_outputs(3401) <= not(layer3_outputs(5914)) or (layer3_outputs(5168));
    layer4_outputs(3402) <= not((layer3_outputs(561)) xor (layer3_outputs(4640)));
    layer4_outputs(3403) <= layer3_outputs(2259);
    layer4_outputs(3404) <= layer3_outputs(2468);
    layer4_outputs(3405) <= '1';
    layer4_outputs(3406) <= (layer3_outputs(7450)) or (layer3_outputs(7289));
    layer4_outputs(3407) <= layer3_outputs(4329);
    layer4_outputs(3408) <= (layer3_outputs(721)) and not (layer3_outputs(5656));
    layer4_outputs(3409) <= not((layer3_outputs(223)) xor (layer3_outputs(6443)));
    layer4_outputs(3410) <= not(layer3_outputs(2228)) or (layer3_outputs(5690));
    layer4_outputs(3411) <= not(layer3_outputs(4461));
    layer4_outputs(3412) <= (layer3_outputs(6011)) and (layer3_outputs(3722));
    layer4_outputs(3413) <= (layer3_outputs(4484)) and not (layer3_outputs(2555));
    layer4_outputs(3414) <= layer3_outputs(2373);
    layer4_outputs(3415) <= (layer3_outputs(2836)) and (layer3_outputs(4455));
    layer4_outputs(3416) <= layer3_outputs(2481);
    layer4_outputs(3417) <= layer3_outputs(6961);
    layer4_outputs(3418) <= (layer3_outputs(2493)) or (layer3_outputs(2546));
    layer4_outputs(3419) <= (layer3_outputs(7033)) xor (layer3_outputs(4562));
    layer4_outputs(3420) <= not(layer3_outputs(6932));
    layer4_outputs(3421) <= not((layer3_outputs(6790)) xor (layer3_outputs(2354)));
    layer4_outputs(3422) <= (layer3_outputs(6975)) or (layer3_outputs(1682));
    layer4_outputs(3423) <= layer3_outputs(3253);
    layer4_outputs(3424) <= not(layer3_outputs(4967)) or (layer3_outputs(7081));
    layer4_outputs(3425) <= (layer3_outputs(86)) or (layer3_outputs(6846));
    layer4_outputs(3426) <= layer3_outputs(5039);
    layer4_outputs(3427) <= not(layer3_outputs(6889)) or (layer3_outputs(270));
    layer4_outputs(3428) <= (layer3_outputs(143)) and (layer3_outputs(4912));
    layer4_outputs(3429) <= layer3_outputs(4975);
    layer4_outputs(3430) <= not(layer3_outputs(4407)) or (layer3_outputs(3947));
    layer4_outputs(3431) <= layer3_outputs(5859);
    layer4_outputs(3432) <= not((layer3_outputs(3488)) and (layer3_outputs(3066)));
    layer4_outputs(3433) <= layer3_outputs(4259);
    layer4_outputs(3434) <= not(layer3_outputs(4675));
    layer4_outputs(3435) <= not(layer3_outputs(2958));
    layer4_outputs(3436) <= not(layer3_outputs(3933));
    layer4_outputs(3437) <= not((layer3_outputs(5868)) xor (layer3_outputs(1419)));
    layer4_outputs(3438) <= not(layer3_outputs(5208));
    layer4_outputs(3439) <= layer3_outputs(628);
    layer4_outputs(3440) <= not((layer3_outputs(578)) xor (layer3_outputs(6898)));
    layer4_outputs(3441) <= not(layer3_outputs(2012)) or (layer3_outputs(4363));
    layer4_outputs(3442) <= (layer3_outputs(5625)) and (layer3_outputs(65));
    layer4_outputs(3443) <= layer3_outputs(5879);
    layer4_outputs(3444) <= layer3_outputs(2586);
    layer4_outputs(3445) <= not(layer3_outputs(5269));
    layer4_outputs(3446) <= not(layer3_outputs(6190));
    layer4_outputs(3447) <= not(layer3_outputs(6276));
    layer4_outputs(3448) <= not(layer3_outputs(912));
    layer4_outputs(3449) <= '0';
    layer4_outputs(3450) <= not(layer3_outputs(7364));
    layer4_outputs(3451) <= not(layer3_outputs(6617));
    layer4_outputs(3452) <= (layer3_outputs(6456)) and not (layer3_outputs(534));
    layer4_outputs(3453) <= (layer3_outputs(67)) and (layer3_outputs(6329));
    layer4_outputs(3454) <= not(layer3_outputs(3345)) or (layer3_outputs(5917));
    layer4_outputs(3455) <= not((layer3_outputs(7160)) or (layer3_outputs(1743)));
    layer4_outputs(3456) <= (layer3_outputs(7210)) or (layer3_outputs(5026));
    layer4_outputs(3457) <= layer3_outputs(2301);
    layer4_outputs(3458) <= layer3_outputs(1607);
    layer4_outputs(3459) <= (layer3_outputs(6359)) and not (layer3_outputs(4367));
    layer4_outputs(3460) <= layer3_outputs(723);
    layer4_outputs(3461) <= (layer3_outputs(3368)) and not (layer3_outputs(7521));
    layer4_outputs(3462) <= layer3_outputs(6682);
    layer4_outputs(3463) <= (layer3_outputs(2918)) and not (layer3_outputs(2000));
    layer4_outputs(3464) <= '0';
    layer4_outputs(3465) <= not((layer3_outputs(4099)) and (layer3_outputs(6760)));
    layer4_outputs(3466) <= not(layer3_outputs(2649));
    layer4_outputs(3467) <= not(layer3_outputs(2467)) or (layer3_outputs(266));
    layer4_outputs(3468) <= layer3_outputs(3107);
    layer4_outputs(3469) <= not(layer3_outputs(4537)) or (layer3_outputs(724));
    layer4_outputs(3470) <= not(layer3_outputs(6553));
    layer4_outputs(3471) <= layer3_outputs(3058);
    layer4_outputs(3472) <= not(layer3_outputs(3896));
    layer4_outputs(3473) <= layer3_outputs(7485);
    layer4_outputs(3474) <= not((layer3_outputs(6791)) xor (layer3_outputs(4030)));
    layer4_outputs(3475) <= layer3_outputs(3653);
    layer4_outputs(3476) <= not(layer3_outputs(3967));
    layer4_outputs(3477) <= not((layer3_outputs(1937)) or (layer3_outputs(3157)));
    layer4_outputs(3478) <= layer3_outputs(5437);
    layer4_outputs(3479) <= layer3_outputs(6577);
    layer4_outputs(3480) <= not(layer3_outputs(2261)) or (layer3_outputs(2430));
    layer4_outputs(3481) <= layer3_outputs(7676);
    layer4_outputs(3482) <= (layer3_outputs(7560)) and not (layer3_outputs(2288));
    layer4_outputs(3483) <= (layer3_outputs(2870)) xor (layer3_outputs(5692));
    layer4_outputs(3484) <= (layer3_outputs(2610)) and not (layer3_outputs(1123));
    layer4_outputs(3485) <= layer3_outputs(3612);
    layer4_outputs(3486) <= layer3_outputs(7417);
    layer4_outputs(3487) <= not(layer3_outputs(4924)) or (layer3_outputs(4548));
    layer4_outputs(3488) <= not(layer3_outputs(849));
    layer4_outputs(3489) <= (layer3_outputs(662)) and not (layer3_outputs(5393));
    layer4_outputs(3490) <= not(layer3_outputs(5734));
    layer4_outputs(3491) <= layer3_outputs(4424);
    layer4_outputs(3492) <= not(layer3_outputs(6625)) or (layer3_outputs(3643));
    layer4_outputs(3493) <= not(layer3_outputs(3682));
    layer4_outputs(3494) <= layer3_outputs(5716);
    layer4_outputs(3495) <= (layer3_outputs(4575)) or (layer3_outputs(3500));
    layer4_outputs(3496) <= layer3_outputs(6387);
    layer4_outputs(3497) <= (layer3_outputs(1930)) and not (layer3_outputs(6580));
    layer4_outputs(3498) <= not(layer3_outputs(1031));
    layer4_outputs(3499) <= not((layer3_outputs(1299)) or (layer3_outputs(1241)));
    layer4_outputs(3500) <= layer3_outputs(3070);
    layer4_outputs(3501) <= not((layer3_outputs(4886)) or (layer3_outputs(1305)));
    layer4_outputs(3502) <= not(layer3_outputs(5628));
    layer4_outputs(3503) <= (layer3_outputs(2232)) and not (layer3_outputs(4465));
    layer4_outputs(3504) <= not(layer3_outputs(7020));
    layer4_outputs(3505) <= not(layer3_outputs(7470));
    layer4_outputs(3506) <= not((layer3_outputs(957)) xor (layer3_outputs(6597)));
    layer4_outputs(3507) <= layer3_outputs(6509);
    layer4_outputs(3508) <= (layer3_outputs(1783)) or (layer3_outputs(7063));
    layer4_outputs(3509) <= (layer3_outputs(2188)) or (layer3_outputs(3850));
    layer4_outputs(3510) <= not(layer3_outputs(386)) or (layer3_outputs(2918));
    layer4_outputs(3511) <= (layer3_outputs(2090)) and not (layer3_outputs(4754));
    layer4_outputs(3512) <= not((layer3_outputs(2251)) and (layer3_outputs(2194)));
    layer4_outputs(3513) <= (layer3_outputs(6339)) and not (layer3_outputs(6692));
    layer4_outputs(3514) <= (layer3_outputs(5838)) and not (layer3_outputs(5827));
    layer4_outputs(3515) <= not(layer3_outputs(362));
    layer4_outputs(3516) <= (layer3_outputs(2037)) and (layer3_outputs(5558));
    layer4_outputs(3517) <= (layer3_outputs(4028)) and not (layer3_outputs(4979));
    layer4_outputs(3518) <= not(layer3_outputs(2194));
    layer4_outputs(3519) <= not(layer3_outputs(4319)) or (layer3_outputs(2845));
    layer4_outputs(3520) <= not((layer3_outputs(739)) or (layer3_outputs(3893)));
    layer4_outputs(3521) <= (layer3_outputs(3531)) and not (layer3_outputs(5238));
    layer4_outputs(3522) <= layer3_outputs(6852);
    layer4_outputs(3523) <= '1';
    layer4_outputs(3524) <= layer3_outputs(4832);
    layer4_outputs(3525) <= layer3_outputs(4187);
    layer4_outputs(3526) <= not(layer3_outputs(6636));
    layer4_outputs(3527) <= (layer3_outputs(6168)) and (layer3_outputs(5546));
    layer4_outputs(3528) <= not(layer3_outputs(6029)) or (layer3_outputs(3741));
    layer4_outputs(3529) <= not(layer3_outputs(1956)) or (layer3_outputs(4815));
    layer4_outputs(3530) <= not(layer3_outputs(6218)) or (layer3_outputs(5496));
    layer4_outputs(3531) <= layer3_outputs(1649);
    layer4_outputs(3532) <= (layer3_outputs(896)) xor (layer3_outputs(5976));
    layer4_outputs(3533) <= (layer3_outputs(4792)) and not (layer3_outputs(7134));
    layer4_outputs(3534) <= '0';
    layer4_outputs(3535) <= not(layer3_outputs(804));
    layer4_outputs(3536) <= not((layer3_outputs(452)) xor (layer3_outputs(7275)));
    layer4_outputs(3537) <= (layer3_outputs(6737)) and not (layer3_outputs(6286));
    layer4_outputs(3538) <= not((layer3_outputs(4656)) and (layer3_outputs(6000)));
    layer4_outputs(3539) <= not(layer3_outputs(7130));
    layer4_outputs(3540) <= not((layer3_outputs(2257)) or (layer3_outputs(648)));
    layer4_outputs(3541) <= not((layer3_outputs(2952)) or (layer3_outputs(6069)));
    layer4_outputs(3542) <= not(layer3_outputs(2892));
    layer4_outputs(3543) <= layer3_outputs(289);
    layer4_outputs(3544) <= not(layer3_outputs(2530)) or (layer3_outputs(6628));
    layer4_outputs(3545) <= not(layer3_outputs(6413)) or (layer3_outputs(4729));
    layer4_outputs(3546) <= layer3_outputs(2911);
    layer4_outputs(3547) <= layer3_outputs(7320);
    layer4_outputs(3548) <= layer3_outputs(7592);
    layer4_outputs(3549) <= (layer3_outputs(55)) or (layer3_outputs(6167));
    layer4_outputs(3550) <= not(layer3_outputs(137));
    layer4_outputs(3551) <= layer3_outputs(5136);
    layer4_outputs(3552) <= not(layer3_outputs(4836));
    layer4_outputs(3553) <= (layer3_outputs(5392)) and (layer3_outputs(209));
    layer4_outputs(3554) <= layer3_outputs(6741);
    layer4_outputs(3555) <= (layer3_outputs(2297)) and not (layer3_outputs(5740));
    layer4_outputs(3556) <= (layer3_outputs(601)) and not (layer3_outputs(3644));
    layer4_outputs(3557) <= (layer3_outputs(7422)) xor (layer3_outputs(376));
    layer4_outputs(3558) <= layer3_outputs(6764);
    layer4_outputs(3559) <= not((layer3_outputs(1928)) or (layer3_outputs(2863)));
    layer4_outputs(3560) <= layer3_outputs(5574);
    layer4_outputs(3561) <= layer3_outputs(1553);
    layer4_outputs(3562) <= layer3_outputs(393);
    layer4_outputs(3563) <= not((layer3_outputs(860)) or (layer3_outputs(6988)));
    layer4_outputs(3564) <= layer3_outputs(4438);
    layer4_outputs(3565) <= not(layer3_outputs(2668));
    layer4_outputs(3566) <= not(layer3_outputs(6344));
    layer4_outputs(3567) <= not(layer3_outputs(855));
    layer4_outputs(3568) <= not(layer3_outputs(7000));
    layer4_outputs(3569) <= not(layer3_outputs(3558));
    layer4_outputs(3570) <= (layer3_outputs(7635)) or (layer3_outputs(1690));
    layer4_outputs(3571) <= not(layer3_outputs(6084));
    layer4_outputs(3572) <= not((layer3_outputs(4293)) and (layer3_outputs(1266)));
    layer4_outputs(3573) <= (layer3_outputs(5632)) and not (layer3_outputs(3508));
    layer4_outputs(3574) <= layer3_outputs(4261);
    layer4_outputs(3575) <= layer3_outputs(3862);
    layer4_outputs(3576) <= not(layer3_outputs(1198));
    layer4_outputs(3577) <= not(layer3_outputs(5341));
    layer4_outputs(3578) <= (layer3_outputs(1313)) and (layer3_outputs(6726));
    layer4_outputs(3579) <= layer3_outputs(2717);
    layer4_outputs(3580) <= not(layer3_outputs(4311));
    layer4_outputs(3581) <= (layer3_outputs(6157)) or (layer3_outputs(6863));
    layer4_outputs(3582) <= not(layer3_outputs(5801));
    layer4_outputs(3583) <= (layer3_outputs(6428)) and (layer3_outputs(1012));
    layer4_outputs(3584) <= layer3_outputs(4521);
    layer4_outputs(3585) <= not(layer3_outputs(6510));
    layer4_outputs(3586) <= not((layer3_outputs(2652)) or (layer3_outputs(4288)));
    layer4_outputs(3587) <= layer3_outputs(1537);
    layer4_outputs(3588) <= layer3_outputs(272);
    layer4_outputs(3589) <= layer3_outputs(32);
    layer4_outputs(3590) <= layer3_outputs(4679);
    layer4_outputs(3591) <= not(layer3_outputs(1900));
    layer4_outputs(3592) <= layer3_outputs(1974);
    layer4_outputs(3593) <= not(layer3_outputs(6955));
    layer4_outputs(3594) <= not((layer3_outputs(3566)) or (layer3_outputs(1030)));
    layer4_outputs(3595) <= (layer3_outputs(1448)) and (layer3_outputs(2477));
    layer4_outputs(3596) <= layer3_outputs(2490);
    layer4_outputs(3597) <= not(layer3_outputs(5013));
    layer4_outputs(3598) <= layer3_outputs(3902);
    layer4_outputs(3599) <= not((layer3_outputs(483)) or (layer3_outputs(593)));
    layer4_outputs(3600) <= (layer3_outputs(4211)) xor (layer3_outputs(1328));
    layer4_outputs(3601) <= layer3_outputs(183);
    layer4_outputs(3602) <= not(layer3_outputs(789));
    layer4_outputs(3603) <= not(layer3_outputs(4019));
    layer4_outputs(3604) <= not(layer3_outputs(3169));
    layer4_outputs(3605) <= not(layer3_outputs(6402));
    layer4_outputs(3606) <= not(layer3_outputs(5513));
    layer4_outputs(3607) <= not((layer3_outputs(2030)) or (layer3_outputs(5980)));
    layer4_outputs(3608) <= (layer3_outputs(7319)) and not (layer3_outputs(5741));
    layer4_outputs(3609) <= (layer3_outputs(3573)) and not (layer3_outputs(5291));
    layer4_outputs(3610) <= layer3_outputs(5410);
    layer4_outputs(3611) <= not((layer3_outputs(187)) or (layer3_outputs(2426)));
    layer4_outputs(3612) <= not(layer3_outputs(3189)) or (layer3_outputs(4391));
    layer4_outputs(3613) <= not(layer3_outputs(5259)) or (layer3_outputs(4275));
    layer4_outputs(3614) <= not((layer3_outputs(2738)) or (layer3_outputs(3123)));
    layer4_outputs(3615) <= (layer3_outputs(5877)) and (layer3_outputs(3066));
    layer4_outputs(3616) <= not(layer3_outputs(6493));
    layer4_outputs(3617) <= (layer3_outputs(4482)) and not (layer3_outputs(5596));
    layer4_outputs(3618) <= layer3_outputs(7032);
    layer4_outputs(3619) <= (layer3_outputs(1704)) and not (layer3_outputs(2612));
    layer4_outputs(3620) <= not((layer3_outputs(4953)) and (layer3_outputs(2106)));
    layer4_outputs(3621) <= not(layer3_outputs(1737));
    layer4_outputs(3622) <= '1';
    layer4_outputs(3623) <= layer3_outputs(5313);
    layer4_outputs(3624) <= not(layer3_outputs(6288));
    layer4_outputs(3625) <= not(layer3_outputs(6164)) or (layer3_outputs(7646));
    layer4_outputs(3626) <= layer3_outputs(1429);
    layer4_outputs(3627) <= not(layer3_outputs(254)) or (layer3_outputs(581));
    layer4_outputs(3628) <= not(layer3_outputs(6640));
    layer4_outputs(3629) <= not(layer3_outputs(584));
    layer4_outputs(3630) <= not(layer3_outputs(1929));
    layer4_outputs(3631) <= not(layer3_outputs(5034));
    layer4_outputs(3632) <= (layer3_outputs(2448)) xor (layer3_outputs(4732));
    layer4_outputs(3633) <= (layer3_outputs(4694)) or (layer3_outputs(4914));
    layer4_outputs(3634) <= (layer3_outputs(907)) and (layer3_outputs(4407));
    layer4_outputs(3635) <= (layer3_outputs(7620)) xor (layer3_outputs(5925));
    layer4_outputs(3636) <= (layer3_outputs(2186)) xor (layer3_outputs(7172));
    layer4_outputs(3637) <= layer3_outputs(2891);
    layer4_outputs(3638) <= layer3_outputs(2275);
    layer4_outputs(3639) <= layer3_outputs(763);
    layer4_outputs(3640) <= not(layer3_outputs(2451));
    layer4_outputs(3641) <= not((layer3_outputs(4209)) and (layer3_outputs(276)));
    layer4_outputs(3642) <= (layer3_outputs(1981)) or (layer3_outputs(6941));
    layer4_outputs(3643) <= not((layer3_outputs(4328)) or (layer3_outputs(4905)));
    layer4_outputs(3644) <= not(layer3_outputs(2083));
    layer4_outputs(3645) <= (layer3_outputs(2033)) and not (layer3_outputs(2327));
    layer4_outputs(3646) <= layer3_outputs(4131);
    layer4_outputs(3647) <= (layer3_outputs(1820)) or (layer3_outputs(3165));
    layer4_outputs(3648) <= (layer3_outputs(982)) xor (layer3_outputs(3892));
    layer4_outputs(3649) <= layer3_outputs(4492);
    layer4_outputs(3650) <= layer3_outputs(1607);
    layer4_outputs(3651) <= layer3_outputs(573);
    layer4_outputs(3652) <= not(layer3_outputs(4672));
    layer4_outputs(3653) <= not(layer3_outputs(3943));
    layer4_outputs(3654) <= not((layer3_outputs(7038)) xor (layer3_outputs(6455)));
    layer4_outputs(3655) <= not((layer3_outputs(4441)) or (layer3_outputs(7338)));
    layer4_outputs(3656) <= not((layer3_outputs(3756)) and (layer3_outputs(660)));
    layer4_outputs(3657) <= layer3_outputs(3136);
    layer4_outputs(3658) <= layer3_outputs(5854);
    layer4_outputs(3659) <= not(layer3_outputs(6209)) or (layer3_outputs(2066));
    layer4_outputs(3660) <= (layer3_outputs(213)) xor (layer3_outputs(6049));
    layer4_outputs(3661) <= (layer3_outputs(884)) and not (layer3_outputs(3777));
    layer4_outputs(3662) <= (layer3_outputs(1076)) xor (layer3_outputs(6566));
    layer4_outputs(3663) <= not((layer3_outputs(1784)) and (layer3_outputs(4037)));
    layer4_outputs(3664) <= not(layer3_outputs(1747));
    layer4_outputs(3665) <= (layer3_outputs(3628)) and not (layer3_outputs(1833));
    layer4_outputs(3666) <= layer3_outputs(3314);
    layer4_outputs(3667) <= not(layer3_outputs(5462));
    layer4_outputs(3668) <= (layer3_outputs(5427)) or (layer3_outputs(4483));
    layer4_outputs(3669) <= not((layer3_outputs(490)) and (layer3_outputs(4595)));
    layer4_outputs(3670) <= (layer3_outputs(4493)) and not (layer3_outputs(4146));
    layer4_outputs(3671) <= not(layer3_outputs(1676));
    layer4_outputs(3672) <= not(layer3_outputs(3766));
    layer4_outputs(3673) <= (layer3_outputs(2495)) and (layer3_outputs(546));
    layer4_outputs(3674) <= (layer3_outputs(773)) and (layer3_outputs(1435));
    layer4_outputs(3675) <= layer3_outputs(1713);
    layer4_outputs(3676) <= (layer3_outputs(6255)) and (layer3_outputs(4134));
    layer4_outputs(3677) <= (layer3_outputs(2638)) and not (layer3_outputs(2102));
    layer4_outputs(3678) <= (layer3_outputs(1940)) and (layer3_outputs(2150));
    layer4_outputs(3679) <= (layer3_outputs(7016)) or (layer3_outputs(3780));
    layer4_outputs(3680) <= layer3_outputs(2459);
    layer4_outputs(3681) <= not(layer3_outputs(7097)) or (layer3_outputs(2093));
    layer4_outputs(3682) <= (layer3_outputs(3016)) and not (layer3_outputs(2690));
    layer4_outputs(3683) <= not(layer3_outputs(353));
    layer4_outputs(3684) <= not(layer3_outputs(6178)) or (layer3_outputs(6847));
    layer4_outputs(3685) <= '1';
    layer4_outputs(3686) <= not(layer3_outputs(1406)) or (layer3_outputs(51));
    layer4_outputs(3687) <= layer3_outputs(4415);
    layer4_outputs(3688) <= not((layer3_outputs(5511)) and (layer3_outputs(1302)));
    layer4_outputs(3689) <= (layer3_outputs(2688)) and (layer3_outputs(131));
    layer4_outputs(3690) <= (layer3_outputs(4111)) and (layer3_outputs(3106));
    layer4_outputs(3691) <= not(layer3_outputs(4196));
    layer4_outputs(3692) <= not(layer3_outputs(4703));
    layer4_outputs(3693) <= not(layer3_outputs(1551));
    layer4_outputs(3694) <= layer3_outputs(4048);
    layer4_outputs(3695) <= layer3_outputs(1479);
    layer4_outputs(3696) <= not(layer3_outputs(4669));
    layer4_outputs(3697) <= layer3_outputs(3646);
    layer4_outputs(3698) <= (layer3_outputs(6935)) and not (layer3_outputs(4466));
    layer4_outputs(3699) <= not((layer3_outputs(4152)) or (layer3_outputs(3310)));
    layer4_outputs(3700) <= not((layer3_outputs(1209)) or (layer3_outputs(5149)));
    layer4_outputs(3701) <= not(layer3_outputs(3851)) or (layer3_outputs(6162));
    layer4_outputs(3702) <= layer3_outputs(4907);
    layer4_outputs(3703) <= layer3_outputs(6043);
    layer4_outputs(3704) <= not(layer3_outputs(2956));
    layer4_outputs(3705) <= (layer3_outputs(4255)) and not (layer3_outputs(3664));
    layer4_outputs(3706) <= not(layer3_outputs(5762));
    layer4_outputs(3707) <= layer3_outputs(1209);
    layer4_outputs(3708) <= layer3_outputs(5580);
    layer4_outputs(3709) <= not(layer3_outputs(4624));
    layer4_outputs(3710) <= not(layer3_outputs(4300));
    layer4_outputs(3711) <= not((layer3_outputs(7242)) or (layer3_outputs(903)));
    layer4_outputs(3712) <= layer3_outputs(3752);
    layer4_outputs(3713) <= layer3_outputs(7008);
    layer4_outputs(3714) <= '0';
    layer4_outputs(3715) <= not((layer3_outputs(2699)) xor (layer3_outputs(2072)));
    layer4_outputs(3716) <= layer3_outputs(2920);
    layer4_outputs(3717) <= not(layer3_outputs(3756));
    layer4_outputs(3718) <= layer3_outputs(2449);
    layer4_outputs(3719) <= layer3_outputs(4865);
    layer4_outputs(3720) <= layer3_outputs(4627);
    layer4_outputs(3721) <= not(layer3_outputs(4148)) or (layer3_outputs(1866));
    layer4_outputs(3722) <= not((layer3_outputs(3843)) xor (layer3_outputs(4079)));
    layer4_outputs(3723) <= (layer3_outputs(2685)) or (layer3_outputs(4401));
    layer4_outputs(3724) <= layer3_outputs(3172);
    layer4_outputs(3725) <= layer3_outputs(2517);
    layer4_outputs(3726) <= not((layer3_outputs(2686)) or (layer3_outputs(2846)));
    layer4_outputs(3727) <= (layer3_outputs(5297)) or (layer3_outputs(2429));
    layer4_outputs(3728) <= not((layer3_outputs(2737)) or (layer3_outputs(6358)));
    layer4_outputs(3729) <= not(layer3_outputs(5035)) or (layer3_outputs(1802));
    layer4_outputs(3730) <= (layer3_outputs(2557)) and not (layer3_outputs(525));
    layer4_outputs(3731) <= not(layer3_outputs(657));
    layer4_outputs(3732) <= (layer3_outputs(173)) xor (layer3_outputs(3197));
    layer4_outputs(3733) <= not(layer3_outputs(4067)) or (layer3_outputs(5792));
    layer4_outputs(3734) <= (layer3_outputs(3419)) and not (layer3_outputs(5064));
    layer4_outputs(3735) <= not((layer3_outputs(4738)) xor (layer3_outputs(6457)));
    layer4_outputs(3736) <= not(layer3_outputs(4323));
    layer4_outputs(3737) <= not(layer3_outputs(6611)) or (layer3_outputs(3220));
    layer4_outputs(3738) <= not(layer3_outputs(1134));
    layer4_outputs(3739) <= not((layer3_outputs(117)) or (layer3_outputs(7198)));
    layer4_outputs(3740) <= (layer3_outputs(3288)) and not (layer3_outputs(4826));
    layer4_outputs(3741) <= not((layer3_outputs(6048)) and (layer3_outputs(7152)));
    layer4_outputs(3742) <= not(layer3_outputs(4140)) or (layer3_outputs(1350));
    layer4_outputs(3743) <= (layer3_outputs(3427)) and not (layer3_outputs(3634));
    layer4_outputs(3744) <= not(layer3_outputs(5688));
    layer4_outputs(3745) <= layer3_outputs(2723);
    layer4_outputs(3746) <= not(layer3_outputs(1099));
    layer4_outputs(3747) <= layer3_outputs(7369);
    layer4_outputs(3748) <= (layer3_outputs(3828)) and not (layer3_outputs(5984));
    layer4_outputs(3749) <= layer3_outputs(7223);
    layer4_outputs(3750) <= not((layer3_outputs(7528)) xor (layer3_outputs(3586)));
    layer4_outputs(3751) <= layer3_outputs(1748);
    layer4_outputs(3752) <= layer3_outputs(5807);
    layer4_outputs(3753) <= layer3_outputs(7478);
    layer4_outputs(3754) <= not(layer3_outputs(4693));
    layer4_outputs(3755) <= not(layer3_outputs(1174));
    layer4_outputs(3756) <= not(layer3_outputs(12));
    layer4_outputs(3757) <= not((layer3_outputs(2290)) or (layer3_outputs(6947)));
    layer4_outputs(3758) <= layer3_outputs(2476);
    layer4_outputs(3759) <= not(layer3_outputs(4477)) or (layer3_outputs(1068));
    layer4_outputs(3760) <= (layer3_outputs(2582)) and not (layer3_outputs(6460));
    layer4_outputs(3761) <= not(layer3_outputs(1510));
    layer4_outputs(3762) <= (layer3_outputs(5213)) xor (layer3_outputs(3648));
    layer4_outputs(3763) <= layer3_outputs(2309);
    layer4_outputs(3764) <= not((layer3_outputs(5120)) or (layer3_outputs(5591)));
    layer4_outputs(3765) <= not(layer3_outputs(1247)) or (layer3_outputs(4848));
    layer4_outputs(3766) <= (layer3_outputs(3966)) and (layer3_outputs(3566));
    layer4_outputs(3767) <= layer3_outputs(7108);
    layer4_outputs(3768) <= layer3_outputs(2605);
    layer4_outputs(3769) <= '1';
    layer4_outputs(3770) <= (layer3_outputs(4177)) and not (layer3_outputs(6389));
    layer4_outputs(3771) <= not(layer3_outputs(6465)) or (layer3_outputs(7258));
    layer4_outputs(3772) <= not(layer3_outputs(6585));
    layer4_outputs(3773) <= not((layer3_outputs(6126)) and (layer3_outputs(6678)));
    layer4_outputs(3774) <= not((layer3_outputs(2819)) and (layer3_outputs(2624)));
    layer4_outputs(3775) <= not(layer3_outputs(2932)) or (layer3_outputs(5242));
    layer4_outputs(3776) <= not(layer3_outputs(6662)) or (layer3_outputs(2661));
    layer4_outputs(3777) <= not(layer3_outputs(3275));
    layer4_outputs(3778) <= layer3_outputs(7277);
    layer4_outputs(3779) <= (layer3_outputs(2388)) or (layer3_outputs(4437));
    layer4_outputs(3780) <= layer3_outputs(6349);
    layer4_outputs(3781) <= (layer3_outputs(2720)) and (layer3_outputs(2048));
    layer4_outputs(3782) <= not((layer3_outputs(4846)) and (layer3_outputs(5694)));
    layer4_outputs(3783) <= layer3_outputs(491);
    layer4_outputs(3784) <= not((layer3_outputs(4708)) and (layer3_outputs(1148)));
    layer4_outputs(3785) <= (layer3_outputs(6101)) and not (layer3_outputs(4190));
    layer4_outputs(3786) <= layer3_outputs(5987);
    layer4_outputs(3787) <= (layer3_outputs(1799)) and not (layer3_outputs(771));
    layer4_outputs(3788) <= not((layer3_outputs(5311)) and (layer3_outputs(3108)));
    layer4_outputs(3789) <= (layer3_outputs(2736)) and not (layer3_outputs(918));
    layer4_outputs(3790) <= not((layer3_outputs(6836)) and (layer3_outputs(715)));
    layer4_outputs(3791) <= layer3_outputs(661);
    layer4_outputs(3792) <= (layer3_outputs(367)) and (layer3_outputs(7430));
    layer4_outputs(3793) <= not(layer3_outputs(2851));
    layer4_outputs(3794) <= not(layer3_outputs(3499));
    layer4_outputs(3795) <= layer3_outputs(2571);
    layer4_outputs(3796) <= (layer3_outputs(7077)) and not (layer3_outputs(2644));
    layer4_outputs(3797) <= not(layer3_outputs(7091));
    layer4_outputs(3798) <= not((layer3_outputs(3531)) or (layer3_outputs(1146)));
    layer4_outputs(3799) <= layer3_outputs(6108);
    layer4_outputs(3800) <= not((layer3_outputs(2534)) xor (layer3_outputs(2831)));
    layer4_outputs(3801) <= (layer3_outputs(1370)) and not (layer3_outputs(6722));
    layer4_outputs(3802) <= layer3_outputs(4343);
    layer4_outputs(3803) <= (layer3_outputs(2263)) xor (layer3_outputs(729));
    layer4_outputs(3804) <= not(layer3_outputs(1388));
    layer4_outputs(3805) <= not(layer3_outputs(3627)) or (layer3_outputs(1754));
    layer4_outputs(3806) <= not(layer3_outputs(6132));
    layer4_outputs(3807) <= (layer3_outputs(5124)) or (layer3_outputs(198));
    layer4_outputs(3808) <= (layer3_outputs(6428)) and not (layer3_outputs(7213));
    layer4_outputs(3809) <= not(layer3_outputs(3622));
    layer4_outputs(3810) <= (layer3_outputs(660)) and (layer3_outputs(7343));
    layer4_outputs(3811) <= (layer3_outputs(5256)) and (layer3_outputs(5472));
    layer4_outputs(3812) <= (layer3_outputs(4348)) and not (layer3_outputs(6825));
    layer4_outputs(3813) <= (layer3_outputs(3142)) and not (layer3_outputs(3163));
    layer4_outputs(3814) <= (layer3_outputs(6798)) and not (layer3_outputs(3260));
    layer4_outputs(3815) <= (layer3_outputs(6806)) or (layer3_outputs(6691));
    layer4_outputs(3816) <= (layer3_outputs(3262)) and not (layer3_outputs(1036));
    layer4_outputs(3817) <= layer3_outputs(5978);
    layer4_outputs(3818) <= not(layer3_outputs(836)) or (layer3_outputs(6110));
    layer4_outputs(3819) <= not(layer3_outputs(6049));
    layer4_outputs(3820) <= (layer3_outputs(6436)) and not (layer3_outputs(6542));
    layer4_outputs(3821) <= layer3_outputs(1726);
    layer4_outputs(3822) <= '0';
    layer4_outputs(3823) <= not((layer3_outputs(6111)) xor (layer3_outputs(1294)));
    layer4_outputs(3824) <= not(layer3_outputs(1640)) or (layer3_outputs(1443));
    layer4_outputs(3825) <= not((layer3_outputs(225)) or (layer3_outputs(5768)));
    layer4_outputs(3826) <= not(layer3_outputs(2619)) or (layer3_outputs(518));
    layer4_outputs(3827) <= (layer3_outputs(6120)) and not (layer3_outputs(6622));
    layer4_outputs(3828) <= not((layer3_outputs(2847)) or (layer3_outputs(1117)));
    layer4_outputs(3829) <= (layer3_outputs(845)) xor (layer3_outputs(1137));
    layer4_outputs(3830) <= layer3_outputs(3850);
    layer4_outputs(3831) <= layer3_outputs(7213);
    layer4_outputs(3832) <= not(layer3_outputs(6144));
    layer4_outputs(3833) <= not(layer3_outputs(604));
    layer4_outputs(3834) <= layer3_outputs(1482);
    layer4_outputs(3835) <= not(layer3_outputs(7479)) or (layer3_outputs(142));
    layer4_outputs(3836) <= (layer3_outputs(3944)) and not (layer3_outputs(6802));
    layer4_outputs(3837) <= layer3_outputs(6009);
    layer4_outputs(3838) <= layer3_outputs(5783);
    layer4_outputs(3839) <= (layer3_outputs(4469)) and (layer3_outputs(2100));
    layer4_outputs(3840) <= not(layer3_outputs(4332));
    layer4_outputs(3841) <= layer3_outputs(4227);
    layer4_outputs(3842) <= (layer3_outputs(811)) and (layer3_outputs(3104));
    layer4_outputs(3843) <= not(layer3_outputs(2603));
    layer4_outputs(3844) <= (layer3_outputs(2817)) and not (layer3_outputs(5465));
    layer4_outputs(3845) <= (layer3_outputs(2009)) and not (layer3_outputs(6847));
    layer4_outputs(3846) <= layer3_outputs(2110);
    layer4_outputs(3847) <= layer3_outputs(7120);
    layer4_outputs(3848) <= (layer3_outputs(5810)) and not (layer3_outputs(3888));
    layer4_outputs(3849) <= layer3_outputs(1892);
    layer4_outputs(3850) <= not((layer3_outputs(2126)) and (layer3_outputs(6467)));
    layer4_outputs(3851) <= layer3_outputs(1275);
    layer4_outputs(3852) <= layer3_outputs(6208);
    layer4_outputs(3853) <= not(layer3_outputs(6254));
    layer4_outputs(3854) <= layer3_outputs(6892);
    layer4_outputs(3855) <= layer3_outputs(1558);
    layer4_outputs(3856) <= (layer3_outputs(5861)) and (layer3_outputs(2238));
    layer4_outputs(3857) <= (layer3_outputs(4182)) and (layer3_outputs(6002));
    layer4_outputs(3858) <= layer3_outputs(6916);
    layer4_outputs(3859) <= layer3_outputs(1283);
    layer4_outputs(3860) <= layer3_outputs(6699);
    layer4_outputs(3861) <= not((layer3_outputs(4906)) xor (layer3_outputs(1090)));
    layer4_outputs(3862) <= not((layer3_outputs(7320)) xor (layer3_outputs(757)));
    layer4_outputs(3863) <= (layer3_outputs(4608)) xor (layer3_outputs(4995));
    layer4_outputs(3864) <= not(layer3_outputs(3478));
    layer4_outputs(3865) <= not((layer3_outputs(4804)) xor (layer3_outputs(2182)));
    layer4_outputs(3866) <= not((layer3_outputs(612)) or (layer3_outputs(3390)));
    layer4_outputs(3867) <= layer3_outputs(2796);
    layer4_outputs(3868) <= not((layer3_outputs(1539)) xor (layer3_outputs(2280)));
    layer4_outputs(3869) <= (layer3_outputs(7044)) and (layer3_outputs(6448));
    layer4_outputs(3870) <= not((layer3_outputs(5635)) xor (layer3_outputs(2045)));
    layer4_outputs(3871) <= not(layer3_outputs(6400));
    layer4_outputs(3872) <= not(layer3_outputs(4369));
    layer4_outputs(3873) <= (layer3_outputs(4395)) and not (layer3_outputs(1633));
    layer4_outputs(3874) <= layer3_outputs(4943);
    layer4_outputs(3875) <= layer3_outputs(4531);
    layer4_outputs(3876) <= not(layer3_outputs(3945)) or (layer3_outputs(5543));
    layer4_outputs(3877) <= not(layer3_outputs(2358));
    layer4_outputs(3878) <= (layer3_outputs(541)) and (layer3_outputs(5200));
    layer4_outputs(3879) <= not(layer3_outputs(6820)) or (layer3_outputs(4121));
    layer4_outputs(3880) <= layer3_outputs(5449);
    layer4_outputs(3881) <= layer3_outputs(7078);
    layer4_outputs(3882) <= (layer3_outputs(3704)) and not (layer3_outputs(5380));
    layer4_outputs(3883) <= layer3_outputs(1674);
    layer4_outputs(3884) <= not(layer3_outputs(1118)) or (layer3_outputs(5222));
    layer4_outputs(3885) <= layer3_outputs(246);
    layer4_outputs(3886) <= not(layer3_outputs(6545));
    layer4_outputs(3887) <= (layer3_outputs(198)) or (layer3_outputs(380));
    layer4_outputs(3888) <= not((layer3_outputs(4154)) xor (layer3_outputs(4378)));
    layer4_outputs(3889) <= layer3_outputs(5564);
    layer4_outputs(3890) <= not((layer3_outputs(4304)) or (layer3_outputs(1345)));
    layer4_outputs(3891) <= not(layer3_outputs(5707));
    layer4_outputs(3892) <= not((layer3_outputs(3137)) or (layer3_outputs(7590)));
    layer4_outputs(3893) <= layer3_outputs(2119);
    layer4_outputs(3894) <= not(layer3_outputs(7574));
    layer4_outputs(3895) <= layer3_outputs(6629);
    layer4_outputs(3896) <= layer3_outputs(1813);
    layer4_outputs(3897) <= not(layer3_outputs(363));
    layer4_outputs(3898) <= (layer3_outputs(6195)) xor (layer3_outputs(6698));
    layer4_outputs(3899) <= layer3_outputs(310);
    layer4_outputs(3900) <= not(layer3_outputs(7090)) or (layer3_outputs(6758));
    layer4_outputs(3901) <= (layer3_outputs(852)) xor (layer3_outputs(622));
    layer4_outputs(3902) <= (layer3_outputs(3118)) and not (layer3_outputs(2042));
    layer4_outputs(3903) <= not(layer3_outputs(497));
    layer4_outputs(3904) <= (layer3_outputs(6754)) and (layer3_outputs(1153));
    layer4_outputs(3905) <= layer3_outputs(263);
    layer4_outputs(3906) <= not(layer3_outputs(6956));
    layer4_outputs(3907) <= not((layer3_outputs(108)) and (layer3_outputs(2573)));
    layer4_outputs(3908) <= not(layer3_outputs(7293));
    layer4_outputs(3909) <= not(layer3_outputs(1056));
    layer4_outputs(3910) <= (layer3_outputs(4161)) and not (layer3_outputs(7390));
    layer4_outputs(3911) <= not(layer3_outputs(5913));
    layer4_outputs(3912) <= layer3_outputs(2202);
    layer4_outputs(3913) <= layer3_outputs(6444);
    layer4_outputs(3914) <= (layer3_outputs(5585)) and not (layer3_outputs(1666));
    layer4_outputs(3915) <= (layer3_outputs(5008)) xor (layer3_outputs(1332));
    layer4_outputs(3916) <= layer3_outputs(6300);
    layer4_outputs(3917) <= layer3_outputs(6630);
    layer4_outputs(3918) <= not((layer3_outputs(2491)) xor (layer3_outputs(5063)));
    layer4_outputs(3919) <= not(layer3_outputs(6377));
    layer4_outputs(3920) <= not(layer3_outputs(2917));
    layer4_outputs(3921) <= layer3_outputs(6279);
    layer4_outputs(3922) <= not(layer3_outputs(699)) or (layer3_outputs(3788));
    layer4_outputs(3923) <= not((layer3_outputs(5388)) xor (layer3_outputs(5478)));
    layer4_outputs(3924) <= not(layer3_outputs(973));
    layer4_outputs(3925) <= not(layer3_outputs(5229)) or (layer3_outputs(5792));
    layer4_outputs(3926) <= '0';
    layer4_outputs(3927) <= not(layer3_outputs(6538)) or (layer3_outputs(619));
    layer4_outputs(3928) <= not(layer3_outputs(4590));
    layer4_outputs(3929) <= layer3_outputs(5543);
    layer4_outputs(3930) <= (layer3_outputs(4010)) xor (layer3_outputs(2476));
    layer4_outputs(3931) <= (layer3_outputs(2587)) or (layer3_outputs(1147));
    layer4_outputs(3932) <= (layer3_outputs(1993)) or (layer3_outputs(4795));
    layer4_outputs(3933) <= (layer3_outputs(7552)) and (layer3_outputs(655));
    layer4_outputs(3934) <= not((layer3_outputs(3515)) or (layer3_outputs(5763)));
    layer4_outputs(3935) <= layer3_outputs(5207);
    layer4_outputs(3936) <= not(layer3_outputs(1326));
    layer4_outputs(3937) <= not((layer3_outputs(6521)) xor (layer3_outputs(1107)));
    layer4_outputs(3938) <= (layer3_outputs(540)) and not (layer3_outputs(6942));
    layer4_outputs(3939) <= '0';
    layer4_outputs(3940) <= (layer3_outputs(7005)) xor (layer3_outputs(4710));
    layer4_outputs(3941) <= not((layer3_outputs(6092)) xor (layer3_outputs(5854)));
    layer4_outputs(3942) <= layer3_outputs(4991);
    layer4_outputs(3943) <= layer3_outputs(3091);
    layer4_outputs(3944) <= not(layer3_outputs(2229));
    layer4_outputs(3945) <= not(layer3_outputs(1380)) or (layer3_outputs(4081));
    layer4_outputs(3946) <= not(layer3_outputs(4736));
    layer4_outputs(3947) <= (layer3_outputs(2407)) xor (layer3_outputs(2533));
    layer4_outputs(3948) <= not((layer3_outputs(2276)) xor (layer3_outputs(1877)));
    layer4_outputs(3949) <= not(layer3_outputs(176)) or (layer3_outputs(3562));
    layer4_outputs(3950) <= layer3_outputs(5320);
    layer4_outputs(3951) <= (layer3_outputs(556)) and not (layer3_outputs(221));
    layer4_outputs(3952) <= not(layer3_outputs(7351));
    layer4_outputs(3953) <= (layer3_outputs(6252)) or (layer3_outputs(1732));
    layer4_outputs(3954) <= not((layer3_outputs(3979)) or (layer3_outputs(7599)));
    layer4_outputs(3955) <= layer3_outputs(2217);
    layer4_outputs(3956) <= layer3_outputs(839);
    layer4_outputs(3957) <= layer3_outputs(6946);
    layer4_outputs(3958) <= (layer3_outputs(5055)) and (layer3_outputs(5468));
    layer4_outputs(3959) <= not((layer3_outputs(445)) and (layer3_outputs(1052)));
    layer4_outputs(3960) <= not(layer3_outputs(7522));
    layer4_outputs(3961) <= not(layer3_outputs(6058));
    layer4_outputs(3962) <= (layer3_outputs(3343)) xor (layer3_outputs(3190));
    layer4_outputs(3963) <= not(layer3_outputs(3581));
    layer4_outputs(3964) <= not(layer3_outputs(6992)) or (layer3_outputs(7283));
    layer4_outputs(3965) <= not(layer3_outputs(7374));
    layer4_outputs(3966) <= not(layer3_outputs(4334));
    layer4_outputs(3967) <= layer3_outputs(4374);
    layer4_outputs(3968) <= layer3_outputs(7668);
    layer4_outputs(3969) <= layer3_outputs(1750);
    layer4_outputs(3970) <= (layer3_outputs(236)) and (layer3_outputs(2909));
    layer4_outputs(3971) <= not(layer3_outputs(2086));
    layer4_outputs(3972) <= not(layer3_outputs(6513));
    layer4_outputs(3973) <= not(layer3_outputs(7606)) or (layer3_outputs(3530));
    layer4_outputs(3974) <= layer3_outputs(528);
    layer4_outputs(3975) <= layer3_outputs(1986);
    layer4_outputs(3976) <= '0';
    layer4_outputs(3977) <= layer3_outputs(6796);
    layer4_outputs(3978) <= (layer3_outputs(6457)) and not (layer3_outputs(1243));
    layer4_outputs(3979) <= not(layer3_outputs(7554));
    layer4_outputs(3980) <= layer3_outputs(5856);
    layer4_outputs(3981) <= not((layer3_outputs(2898)) xor (layer3_outputs(3385)));
    layer4_outputs(3982) <= (layer3_outputs(1867)) xor (layer3_outputs(1319));
    layer4_outputs(3983) <= not((layer3_outputs(6222)) xor (layer3_outputs(7636)));
    layer4_outputs(3984) <= not((layer3_outputs(2245)) xor (layer3_outputs(7121)));
    layer4_outputs(3985) <= not(layer3_outputs(3462));
    layer4_outputs(3986) <= not(layer3_outputs(2880));
    layer4_outputs(3987) <= layer3_outputs(121);
    layer4_outputs(3988) <= (layer3_outputs(4874)) xor (layer3_outputs(6299));
    layer4_outputs(3989) <= not(layer3_outputs(2781));
    layer4_outputs(3990) <= layer3_outputs(6397);
    layer4_outputs(3991) <= (layer3_outputs(2409)) and (layer3_outputs(5234));
    layer4_outputs(3992) <= not(layer3_outputs(4201));
    layer4_outputs(3993) <= not(layer3_outputs(4825));
    layer4_outputs(3994) <= not(layer3_outputs(5381)) or (layer3_outputs(1828));
    layer4_outputs(3995) <= (layer3_outputs(6064)) and not (layer3_outputs(983));
    layer4_outputs(3996) <= layer3_outputs(3600);
    layer4_outputs(3997) <= not(layer3_outputs(3033)) or (layer3_outputs(984));
    layer4_outputs(3998) <= not(layer3_outputs(4782));
    layer4_outputs(3999) <= not(layer3_outputs(7293));
    layer4_outputs(4000) <= not(layer3_outputs(6758)) or (layer3_outputs(4023));
    layer4_outputs(4001) <= (layer3_outputs(341)) xor (layer3_outputs(3006));
    layer4_outputs(4002) <= not(layer3_outputs(4075)) or (layer3_outputs(2664));
    layer4_outputs(4003) <= not(layer3_outputs(5894));
    layer4_outputs(4004) <= layer3_outputs(683);
    layer4_outputs(4005) <= layer3_outputs(4063);
    layer4_outputs(4006) <= layer3_outputs(3560);
    layer4_outputs(4007) <= (layer3_outputs(7585)) and not (layer3_outputs(5849));
    layer4_outputs(4008) <= not((layer3_outputs(5857)) and (layer3_outputs(614)));
    layer4_outputs(4009) <= not(layer3_outputs(1160));
    layer4_outputs(4010) <= (layer3_outputs(3581)) and (layer3_outputs(5689));
    layer4_outputs(4011) <= layer3_outputs(2039);
    layer4_outputs(4012) <= not(layer3_outputs(7224));
    layer4_outputs(4013) <= not(layer3_outputs(1003));
    layer4_outputs(4014) <= (layer3_outputs(7225)) xor (layer3_outputs(6646));
    layer4_outputs(4015) <= layer3_outputs(2443);
    layer4_outputs(4016) <= not(layer3_outputs(5649));
    layer4_outputs(4017) <= '0';
    layer4_outputs(4018) <= (layer3_outputs(4465)) xor (layer3_outputs(5911));
    layer4_outputs(4019) <= not((layer3_outputs(2500)) xor (layer3_outputs(3948)));
    layer4_outputs(4020) <= not((layer3_outputs(5932)) xor (layer3_outputs(4951)));
    layer4_outputs(4021) <= not(layer3_outputs(606));
    layer4_outputs(4022) <= layer3_outputs(1231);
    layer4_outputs(4023) <= not(layer3_outputs(3500)) or (layer3_outputs(2275));
    layer4_outputs(4024) <= layer3_outputs(3446);
    layer4_outputs(4025) <= layer3_outputs(5486);
    layer4_outputs(4026) <= not(layer3_outputs(4366)) or (layer3_outputs(5687));
    layer4_outputs(4027) <= (layer3_outputs(542)) xor (layer3_outputs(6202));
    layer4_outputs(4028) <= layer3_outputs(4863);
    layer4_outputs(4029) <= (layer3_outputs(7072)) or (layer3_outputs(1515));
    layer4_outputs(4030) <= not(layer3_outputs(296));
    layer4_outputs(4031) <= not(layer3_outputs(3164));
    layer4_outputs(4032) <= (layer3_outputs(4973)) xor (layer3_outputs(423));
    layer4_outputs(4033) <= not(layer3_outputs(7008));
    layer4_outputs(4034) <= layer3_outputs(3911);
    layer4_outputs(4035) <= not(layer3_outputs(1664)) or (layer3_outputs(2139));
    layer4_outputs(4036) <= (layer3_outputs(6746)) and (layer3_outputs(1190));
    layer4_outputs(4037) <= layer3_outputs(5080);
    layer4_outputs(4038) <= (layer3_outputs(6827)) and not (layer3_outputs(5483));
    layer4_outputs(4039) <= layer3_outputs(3089);
    layer4_outputs(4040) <= not(layer3_outputs(2056)) or (layer3_outputs(364));
    layer4_outputs(4041) <= (layer3_outputs(2906)) and not (layer3_outputs(746));
    layer4_outputs(4042) <= not((layer3_outputs(6631)) and (layer3_outputs(3611)));
    layer4_outputs(4043) <= layer3_outputs(488);
    layer4_outputs(4044) <= not(layer3_outputs(4054));
    layer4_outputs(4045) <= not(layer3_outputs(3162)) or (layer3_outputs(35));
    layer4_outputs(4046) <= layer3_outputs(5435);
    layer4_outputs(4047) <= not(layer3_outputs(2038));
    layer4_outputs(4048) <= layer3_outputs(6797);
    layer4_outputs(4049) <= not((layer3_outputs(536)) xor (layer3_outputs(2418)));
    layer4_outputs(4050) <= (layer3_outputs(263)) or (layer3_outputs(3195));
    layer4_outputs(4051) <= (layer3_outputs(2326)) and (layer3_outputs(5208));
    layer4_outputs(4052) <= (layer3_outputs(2881)) and (layer3_outputs(7401));
    layer4_outputs(4053) <= '1';
    layer4_outputs(4054) <= not(layer3_outputs(6795));
    layer4_outputs(4055) <= (layer3_outputs(6788)) or (layer3_outputs(2874));
    layer4_outputs(4056) <= not(layer3_outputs(4756));
    layer4_outputs(4057) <= not(layer3_outputs(89)) or (layer3_outputs(4242));
    layer4_outputs(4058) <= layer3_outputs(3791);
    layer4_outputs(4059) <= (layer3_outputs(2126)) and (layer3_outputs(3795));
    layer4_outputs(4060) <= not(layer3_outputs(5775));
    layer4_outputs(4061) <= layer3_outputs(6338);
    layer4_outputs(4062) <= layer3_outputs(1763);
    layer4_outputs(4063) <= layer3_outputs(5691);
    layer4_outputs(4064) <= (layer3_outputs(7504)) and not (layer3_outputs(922));
    layer4_outputs(4065) <= (layer3_outputs(5769)) and not (layer3_outputs(6158));
    layer4_outputs(4066) <= (layer3_outputs(559)) and (layer3_outputs(900));
    layer4_outputs(4067) <= not(layer3_outputs(158));
    layer4_outputs(4068) <= (layer3_outputs(6357)) and not (layer3_outputs(1000));
    layer4_outputs(4069) <= not(layer3_outputs(7356));
    layer4_outputs(4070) <= (layer3_outputs(3989)) or (layer3_outputs(4901));
    layer4_outputs(4071) <= layer3_outputs(6518);
    layer4_outputs(4072) <= not(layer3_outputs(7327));
    layer4_outputs(4073) <= layer3_outputs(2456);
    layer4_outputs(4074) <= layer3_outputs(7181);
    layer4_outputs(4075) <= (layer3_outputs(5997)) and (layer3_outputs(1903));
    layer4_outputs(4076) <= layer3_outputs(88);
    layer4_outputs(4077) <= layer3_outputs(455);
    layer4_outputs(4078) <= layer3_outputs(3870);
    layer4_outputs(4079) <= not(layer3_outputs(5566));
    layer4_outputs(4080) <= (layer3_outputs(5238)) and not (layer3_outputs(3577));
    layer4_outputs(4081) <= not(layer3_outputs(4344));
    layer4_outputs(4082) <= layer3_outputs(5561);
    layer4_outputs(4083) <= (layer3_outputs(2270)) or (layer3_outputs(5243));
    layer4_outputs(4084) <= not(layer3_outputs(6826));
    layer4_outputs(4085) <= not(layer3_outputs(2242)) or (layer3_outputs(1817));
    layer4_outputs(4086) <= not(layer3_outputs(5816));
    layer4_outputs(4087) <= not(layer3_outputs(3635));
    layer4_outputs(4088) <= layer3_outputs(2820);
    layer4_outputs(4089) <= layer3_outputs(6177);
    layer4_outputs(4090) <= not((layer3_outputs(3887)) xor (layer3_outputs(5010)));
    layer4_outputs(4091) <= layer3_outputs(7456);
    layer4_outputs(4092) <= not(layer3_outputs(3847));
    layer4_outputs(4093) <= not((layer3_outputs(3436)) or (layer3_outputs(1550)));
    layer4_outputs(4094) <= not(layer3_outputs(4744));
    layer4_outputs(4095) <= layer3_outputs(6872);
    layer4_outputs(4096) <= not((layer3_outputs(7126)) xor (layer3_outputs(2663)));
    layer4_outputs(4097) <= layer3_outputs(1852);
    layer4_outputs(4098) <= layer3_outputs(2213);
    layer4_outputs(4099) <= (layer3_outputs(5568)) and (layer3_outputs(1236));
    layer4_outputs(4100) <= layer3_outputs(1219);
    layer4_outputs(4101) <= not((layer3_outputs(1501)) xor (layer3_outputs(3471)));
    layer4_outputs(4102) <= layer3_outputs(7187);
    layer4_outputs(4103) <= (layer3_outputs(6702)) and not (layer3_outputs(4933));
    layer4_outputs(4104) <= not(layer3_outputs(7576)) or (layer3_outputs(6474));
    layer4_outputs(4105) <= not((layer3_outputs(5534)) and (layer3_outputs(2087)));
    layer4_outputs(4106) <= not((layer3_outputs(4904)) xor (layer3_outputs(2599)));
    layer4_outputs(4107) <= not((layer3_outputs(2343)) or (layer3_outputs(4164)));
    layer4_outputs(4108) <= layer3_outputs(4724);
    layer4_outputs(4109) <= not(layer3_outputs(4717)) or (layer3_outputs(3000));
    layer4_outputs(4110) <= not((layer3_outputs(2960)) or (layer3_outputs(6540)));
    layer4_outputs(4111) <= (layer3_outputs(4206)) and not (layer3_outputs(3882));
    layer4_outputs(4112) <= not(layer3_outputs(2127));
    layer4_outputs(4113) <= not(layer3_outputs(4777));
    layer4_outputs(4114) <= not(layer3_outputs(684));
    layer4_outputs(4115) <= not(layer3_outputs(4433));
    layer4_outputs(4116) <= not(layer3_outputs(949));
    layer4_outputs(4117) <= (layer3_outputs(3390)) and not (layer3_outputs(1786));
    layer4_outputs(4118) <= not(layer3_outputs(2130)) or (layer3_outputs(935));
    layer4_outputs(4119) <= (layer3_outputs(4036)) or (layer3_outputs(6582));
    layer4_outputs(4120) <= not(layer3_outputs(6647));
    layer4_outputs(4121) <= (layer3_outputs(4621)) and not (layer3_outputs(5265));
    layer4_outputs(4122) <= (layer3_outputs(3130)) or (layer3_outputs(3236));
    layer4_outputs(4123) <= '1';
    layer4_outputs(4124) <= (layer3_outputs(772)) xor (layer3_outputs(7383));
    layer4_outputs(4125) <= not(layer3_outputs(1979));
    layer4_outputs(4126) <= not(layer3_outputs(7376));
    layer4_outputs(4127) <= not(layer3_outputs(1016));
    layer4_outputs(4128) <= layer3_outputs(697);
    layer4_outputs(4129) <= not((layer3_outputs(1885)) xor (layer3_outputs(1678)));
    layer4_outputs(4130) <= not(layer3_outputs(381));
    layer4_outputs(4131) <= (layer3_outputs(2748)) xor (layer3_outputs(1995));
    layer4_outputs(4132) <= not((layer3_outputs(2145)) and (layer3_outputs(2639)));
    layer4_outputs(4133) <= (layer3_outputs(2173)) and not (layer3_outputs(7129));
    layer4_outputs(4134) <= layer3_outputs(4823);
    layer4_outputs(4135) <= (layer3_outputs(1982)) and not (layer3_outputs(1996));
    layer4_outputs(4136) <= (layer3_outputs(3752)) xor (layer3_outputs(7258));
    layer4_outputs(4137) <= layer3_outputs(336);
    layer4_outputs(4138) <= layer3_outputs(2897);
    layer4_outputs(4139) <= not((layer3_outputs(4941)) or (layer3_outputs(3792)));
    layer4_outputs(4140) <= layer3_outputs(6278);
    layer4_outputs(4141) <= layer3_outputs(6633);
    layer4_outputs(4142) <= layer3_outputs(2353);
    layer4_outputs(4143) <= not(layer3_outputs(7538));
    layer4_outputs(4144) <= not(layer3_outputs(7197)) or (layer3_outputs(1783));
    layer4_outputs(4145) <= layer3_outputs(2705);
    layer4_outputs(4146) <= not(layer3_outputs(107));
    layer4_outputs(4147) <= not(layer3_outputs(5627)) or (layer3_outputs(4353));
    layer4_outputs(4148) <= '1';
    layer4_outputs(4149) <= not((layer3_outputs(7318)) or (layer3_outputs(302)));
    layer4_outputs(4150) <= not(layer3_outputs(4616));
    layer4_outputs(4151) <= not(layer3_outputs(4155));
    layer4_outputs(4152) <= not(layer3_outputs(1331)) or (layer3_outputs(3275));
    layer4_outputs(4153) <= layer3_outputs(2273);
    layer4_outputs(4154) <= layer3_outputs(747);
    layer4_outputs(4155) <= (layer3_outputs(4090)) and (layer3_outputs(5707));
    layer4_outputs(4156) <= not(layer3_outputs(2259));
    layer4_outputs(4157) <= not((layer3_outputs(2060)) xor (layer3_outputs(6552)));
    layer4_outputs(4158) <= not(layer3_outputs(1883));
    layer4_outputs(4159) <= layer3_outputs(5896);
    layer4_outputs(4160) <= (layer3_outputs(2331)) or (layer3_outputs(5310));
    layer4_outputs(4161) <= layer3_outputs(3224);
    layer4_outputs(4162) <= not(layer3_outputs(7063));
    layer4_outputs(4163) <= (layer3_outputs(1100)) or (layer3_outputs(155));
    layer4_outputs(4164) <= not(layer3_outputs(2762));
    layer4_outputs(4165) <= not(layer3_outputs(6097)) or (layer3_outputs(6309));
    layer4_outputs(4166) <= layer3_outputs(4956);
    layer4_outputs(4167) <= not((layer3_outputs(5552)) xor (layer3_outputs(2330)));
    layer4_outputs(4168) <= '0';
    layer4_outputs(4169) <= not((layer3_outputs(4506)) xor (layer3_outputs(463)));
    layer4_outputs(4170) <= layer3_outputs(2808);
    layer4_outputs(4171) <= (layer3_outputs(2683)) and not (layer3_outputs(7645));
    layer4_outputs(4172) <= not(layer3_outputs(6406));
    layer4_outputs(4173) <= not(layer3_outputs(1119));
    layer4_outputs(4174) <= layer3_outputs(2577);
    layer4_outputs(4175) <= not(layer3_outputs(3330));
    layer4_outputs(4176) <= not(layer3_outputs(5642));
    layer4_outputs(4177) <= '0';
    layer4_outputs(4178) <= (layer3_outputs(6199)) and not (layer3_outputs(1238));
    layer4_outputs(4179) <= layer3_outputs(3766);
    layer4_outputs(4180) <= (layer3_outputs(5071)) xor (layer3_outputs(4891));
    layer4_outputs(4181) <= not(layer3_outputs(2365));
    layer4_outputs(4182) <= (layer3_outputs(3352)) and (layer3_outputs(376));
    layer4_outputs(4183) <= layer3_outputs(2233);
    layer4_outputs(4184) <= layer3_outputs(7105);
    layer4_outputs(4185) <= not(layer3_outputs(5216)) or (layer3_outputs(4813));
    layer4_outputs(4186) <= (layer3_outputs(778)) and not (layer3_outputs(3932));
    layer4_outputs(4187) <= not(layer3_outputs(345));
    layer4_outputs(4188) <= layer3_outputs(7153);
    layer4_outputs(4189) <= not((layer3_outputs(2319)) xor (layer3_outputs(2238)));
    layer4_outputs(4190) <= not(layer3_outputs(4808)) or (layer3_outputs(7375));
    layer4_outputs(4191) <= (layer3_outputs(418)) and not (layer3_outputs(1932));
    layer4_outputs(4192) <= not((layer3_outputs(828)) and (layer3_outputs(3299)));
    layer4_outputs(4193) <= not(layer3_outputs(4162));
    layer4_outputs(4194) <= not((layer3_outputs(6731)) or (layer3_outputs(6572)));
    layer4_outputs(4195) <= not(layer3_outputs(4432));
    layer4_outputs(4196) <= not(layer3_outputs(3233));
    layer4_outputs(4197) <= not(layer3_outputs(6905));
    layer4_outputs(4198) <= not(layer3_outputs(2831));
    layer4_outputs(4199) <= (layer3_outputs(2936)) and not (layer3_outputs(5767));
    layer4_outputs(4200) <= not(layer3_outputs(5990));
    layer4_outputs(4201) <= (layer3_outputs(6524)) and not (layer3_outputs(7484));
    layer4_outputs(4202) <= not(layer3_outputs(417)) or (layer3_outputs(2252));
    layer4_outputs(4203) <= (layer3_outputs(1104)) or (layer3_outputs(835));
    layer4_outputs(4204) <= layer3_outputs(3075);
    layer4_outputs(4205) <= (layer3_outputs(4654)) xor (layer3_outputs(7002));
    layer4_outputs(4206) <= not(layer3_outputs(4050)) or (layer3_outputs(3804));
    layer4_outputs(4207) <= not(layer3_outputs(3526)) or (layer3_outputs(4769));
    layer4_outputs(4208) <= (layer3_outputs(7080)) xor (layer3_outputs(7324));
    layer4_outputs(4209) <= (layer3_outputs(1563)) and (layer3_outputs(7362));
    layer4_outputs(4210) <= layer3_outputs(5204);
    layer4_outputs(4211) <= layer3_outputs(1792);
    layer4_outputs(4212) <= not((layer3_outputs(494)) or (layer3_outputs(5511)));
    layer4_outputs(4213) <= not(layer3_outputs(6355)) or (layer3_outputs(6671));
    layer4_outputs(4214) <= not(layer3_outputs(141));
    layer4_outputs(4215) <= not((layer3_outputs(5225)) or (layer3_outputs(5539)));
    layer4_outputs(4216) <= not(layer3_outputs(3391)) or (layer3_outputs(4648));
    layer4_outputs(4217) <= layer3_outputs(2948);
    layer4_outputs(4218) <= not(layer3_outputs(6544));
    layer4_outputs(4219) <= not(layer3_outputs(7189)) or (layer3_outputs(7429));
    layer4_outputs(4220) <= not((layer3_outputs(7022)) and (layer3_outputs(797)));
    layer4_outputs(4221) <= not(layer3_outputs(6272));
    layer4_outputs(4222) <= not(layer3_outputs(3703)) or (layer3_outputs(5674));
    layer4_outputs(4223) <= not(layer3_outputs(3223));
    layer4_outputs(4224) <= layer3_outputs(2509);
    layer4_outputs(4225) <= (layer3_outputs(4525)) and (layer3_outputs(981));
    layer4_outputs(4226) <= not(layer3_outputs(1323)) or (layer3_outputs(4722));
    layer4_outputs(4227) <= not(layer3_outputs(7638));
    layer4_outputs(4228) <= not((layer3_outputs(6982)) or (layer3_outputs(6065)));
    layer4_outputs(4229) <= (layer3_outputs(5576)) and not (layer3_outputs(7199));
    layer4_outputs(4230) <= not(layer3_outputs(3102));
    layer4_outputs(4231) <= not(layer3_outputs(7515));
    layer4_outputs(4232) <= layer3_outputs(6376);
    layer4_outputs(4233) <= (layer3_outputs(4567)) or (layer3_outputs(1167));
    layer4_outputs(4234) <= layer3_outputs(6775);
    layer4_outputs(4235) <= not((layer3_outputs(4167)) xor (layer3_outputs(6599)));
    layer4_outputs(4236) <= not(layer3_outputs(3521));
    layer4_outputs(4237) <= layer3_outputs(3701);
    layer4_outputs(4238) <= (layer3_outputs(3485)) or (layer3_outputs(6409));
    layer4_outputs(4239) <= (layer3_outputs(2976)) or (layer3_outputs(2521));
    layer4_outputs(4240) <= layer3_outputs(5488);
    layer4_outputs(4241) <= not((layer3_outputs(3813)) or (layer3_outputs(4873)));
    layer4_outputs(4242) <= layer3_outputs(6114);
    layer4_outputs(4243) <= not(layer3_outputs(201));
    layer4_outputs(4244) <= layer3_outputs(2283);
    layer4_outputs(4245) <= '0';
    layer4_outputs(4246) <= not((layer3_outputs(5450)) or (layer3_outputs(6850)));
    layer4_outputs(4247) <= layer3_outputs(5185);
    layer4_outputs(4248) <= not(layer3_outputs(5817)) or (layer3_outputs(6115));
    layer4_outputs(4249) <= (layer3_outputs(2383)) xor (layer3_outputs(6748));
    layer4_outputs(4250) <= (layer3_outputs(1029)) xor (layer3_outputs(6981));
    layer4_outputs(4251) <= (layer3_outputs(7217)) and not (layer3_outputs(2552));
    layer4_outputs(4252) <= (layer3_outputs(7159)) and not (layer3_outputs(7087));
    layer4_outputs(4253) <= not(layer3_outputs(6655)) or (layer3_outputs(3008));
    layer4_outputs(4254) <= layer3_outputs(4026);
    layer4_outputs(4255) <= not((layer3_outputs(603)) or (layer3_outputs(3517)));
    layer4_outputs(4256) <= (layer3_outputs(2824)) xor (layer3_outputs(5317));
    layer4_outputs(4257) <= layer3_outputs(7462);
    layer4_outputs(4258) <= not(layer3_outputs(7140)) or (layer3_outputs(2753));
    layer4_outputs(4259) <= (layer3_outputs(5219)) or (layer3_outputs(1094));
    layer4_outputs(4260) <= layer3_outputs(6712);
    layer4_outputs(4261) <= not(layer3_outputs(4462)) or (layer3_outputs(7614));
    layer4_outputs(4262) <= layer3_outputs(188);
    layer4_outputs(4263) <= layer3_outputs(1579);
    layer4_outputs(4264) <= layer3_outputs(2684);
    layer4_outputs(4265) <= (layer3_outputs(7655)) and (layer3_outputs(6253));
    layer4_outputs(4266) <= not((layer3_outputs(2080)) xor (layer3_outputs(3676)));
    layer4_outputs(4267) <= not(layer3_outputs(4676));
    layer4_outputs(4268) <= not(layer3_outputs(323)) or (layer3_outputs(7668));
    layer4_outputs(4269) <= not((layer3_outputs(419)) or (layer3_outputs(6260)));
    layer4_outputs(4270) <= layer3_outputs(4842);
    layer4_outputs(4271) <= not((layer3_outputs(2076)) xor (layer3_outputs(5850)));
    layer4_outputs(4272) <= not((layer3_outputs(3426)) xor (layer3_outputs(5651)));
    layer4_outputs(4273) <= not(layer3_outputs(2930));
    layer4_outputs(4274) <= not(layer3_outputs(6741)) or (layer3_outputs(7678));
    layer4_outputs(4275) <= layer3_outputs(5257);
    layer4_outputs(4276) <= (layer3_outputs(5606)) and (layer3_outputs(5098));
    layer4_outputs(4277) <= (layer3_outputs(308)) xor (layer3_outputs(3049));
    layer4_outputs(4278) <= not((layer3_outputs(3214)) xor (layer3_outputs(1488)));
    layer4_outputs(4279) <= not((layer3_outputs(5756)) xor (layer3_outputs(4185)));
    layer4_outputs(4280) <= layer3_outputs(299);
    layer4_outputs(4281) <= not(layer3_outputs(5378));
    layer4_outputs(4282) <= not(layer3_outputs(1378));
    layer4_outputs(4283) <= not(layer3_outputs(6823));
    layer4_outputs(4284) <= (layer3_outputs(6928)) xor (layer3_outputs(6690));
    layer4_outputs(4285) <= layer3_outputs(1536);
    layer4_outputs(4286) <= (layer3_outputs(1643)) and not (layer3_outputs(3376));
    layer4_outputs(4287) <= not(layer3_outputs(3765));
    layer4_outputs(4288) <= (layer3_outputs(574)) xor (layer3_outputs(6134));
    layer4_outputs(4289) <= not((layer3_outputs(986)) or (layer3_outputs(6770)));
    layer4_outputs(4290) <= not((layer3_outputs(6233)) xor (layer3_outputs(2772)));
    layer4_outputs(4291) <= layer3_outputs(6634);
    layer4_outputs(4292) <= layer3_outputs(1199);
    layer4_outputs(4293) <= layer3_outputs(7448);
    layer4_outputs(4294) <= (layer3_outputs(1531)) xor (layer3_outputs(1725));
    layer4_outputs(4295) <= not(layer3_outputs(7137));
    layer4_outputs(4296) <= not((layer3_outputs(2652)) xor (layer3_outputs(5574)));
    layer4_outputs(4297) <= layer3_outputs(6968);
    layer4_outputs(4298) <= layer3_outputs(1489);
    layer4_outputs(4299) <= layer3_outputs(5631);
    layer4_outputs(4300) <= not(layer3_outputs(3993)) or (layer3_outputs(5378));
    layer4_outputs(4301) <= not(layer3_outputs(2304));
    layer4_outputs(4302) <= layer3_outputs(7514);
    layer4_outputs(4303) <= not(layer3_outputs(2764)) or (layer3_outputs(5064));
    layer4_outputs(4304) <= not(layer3_outputs(2771));
    layer4_outputs(4305) <= (layer3_outputs(6746)) and (layer3_outputs(7587));
    layer4_outputs(4306) <= (layer3_outputs(547)) and not (layer3_outputs(9));
    layer4_outputs(4307) <= not(layer3_outputs(1666)) or (layer3_outputs(1746));
    layer4_outputs(4308) <= layer3_outputs(5837);
    layer4_outputs(4309) <= not(layer3_outputs(4963));
    layer4_outputs(4310) <= not((layer3_outputs(4818)) and (layer3_outputs(3715)));
    layer4_outputs(4311) <= layer3_outputs(3731);
    layer4_outputs(4312) <= '1';
    layer4_outputs(4313) <= not(layer3_outputs(5405));
    layer4_outputs(4314) <= layer3_outputs(25);
    layer4_outputs(4315) <= (layer3_outputs(677)) and not (layer3_outputs(962));
    layer4_outputs(4316) <= not(layer3_outputs(4759));
    layer4_outputs(4317) <= layer3_outputs(434);
    layer4_outputs(4318) <= not(layer3_outputs(966));
    layer4_outputs(4319) <= layer3_outputs(1679);
    layer4_outputs(4320) <= not((layer3_outputs(3699)) or (layer3_outputs(997)));
    layer4_outputs(4321) <= not(layer3_outputs(1381));
    layer4_outputs(4322) <= not(layer3_outputs(5749)) or (layer3_outputs(5751));
    layer4_outputs(4323) <= not(layer3_outputs(3861)) or (layer3_outputs(5521));
    layer4_outputs(4324) <= not(layer3_outputs(4798));
    layer4_outputs(4325) <= layer3_outputs(219);
    layer4_outputs(4326) <= (layer3_outputs(5510)) and not (layer3_outputs(3786));
    layer4_outputs(4327) <= (layer3_outputs(669)) and (layer3_outputs(2723));
    layer4_outputs(4328) <= not(layer3_outputs(6780));
    layer4_outputs(4329) <= not(layer3_outputs(5015)) or (layer3_outputs(7452));
    layer4_outputs(4330) <= not(layer3_outputs(4960)) or (layer3_outputs(485));
    layer4_outputs(4331) <= (layer3_outputs(2161)) and not (layer3_outputs(5383));
    layer4_outputs(4332) <= not((layer3_outputs(5072)) or (layer3_outputs(6729)));
    layer4_outputs(4333) <= not((layer3_outputs(7259)) and (layer3_outputs(663)));
    layer4_outputs(4334) <= not(layer3_outputs(4458));
    layer4_outputs(4335) <= layer3_outputs(5532);
    layer4_outputs(4336) <= (layer3_outputs(3524)) xor (layer3_outputs(3355));
    layer4_outputs(4337) <= (layer3_outputs(1975)) and not (layer3_outputs(5508));
    layer4_outputs(4338) <= layer3_outputs(4663);
    layer4_outputs(4339) <= layer3_outputs(6978);
    layer4_outputs(4340) <= not((layer3_outputs(2759)) xor (layer3_outputs(5340)));
    layer4_outputs(4341) <= (layer3_outputs(2070)) or (layer3_outputs(7124));
    layer4_outputs(4342) <= (layer3_outputs(5610)) xor (layer3_outputs(4342));
    layer4_outputs(4343) <= (layer3_outputs(159)) xor (layer3_outputs(2479));
    layer4_outputs(4344) <= (layer3_outputs(814)) and (layer3_outputs(6893));
    layer4_outputs(4345) <= layer3_outputs(2550);
    layer4_outputs(4346) <= not((layer3_outputs(6631)) xor (layer3_outputs(7188)));
    layer4_outputs(4347) <= layer3_outputs(6951);
    layer4_outputs(4348) <= layer3_outputs(3884);
    layer4_outputs(4349) <= (layer3_outputs(1486)) and not (layer3_outputs(3810));
    layer4_outputs(4350) <= not(layer3_outputs(424));
    layer4_outputs(4351) <= (layer3_outputs(7321)) or (layer3_outputs(206));
    layer4_outputs(4352) <= not(layer3_outputs(2253));
    layer4_outputs(4353) <= (layer3_outputs(6362)) xor (layer3_outputs(3024));
    layer4_outputs(4354) <= (layer3_outputs(514)) xor (layer3_outputs(2672));
    layer4_outputs(4355) <= layer3_outputs(3782);
    layer4_outputs(4356) <= layer3_outputs(4392);
    layer4_outputs(4357) <= not(layer3_outputs(5773)) or (layer3_outputs(7371));
    layer4_outputs(4358) <= (layer3_outputs(1741)) xor (layer3_outputs(806));
    layer4_outputs(4359) <= layer3_outputs(5311);
    layer4_outputs(4360) <= not(layer3_outputs(6143));
    layer4_outputs(4361) <= not(layer3_outputs(4932));
    layer4_outputs(4362) <= (layer3_outputs(2633)) xor (layer3_outputs(4709));
    layer4_outputs(4363) <= layer3_outputs(1848);
    layer4_outputs(4364) <= (layer3_outputs(3759)) and (layer3_outputs(5167));
    layer4_outputs(4365) <= (layer3_outputs(5681)) and not (layer3_outputs(3358));
    layer4_outputs(4366) <= (layer3_outputs(2408)) and not (layer3_outputs(3185));
    layer4_outputs(4367) <= not(layer3_outputs(358)) or (layer3_outputs(3731));
    layer4_outputs(4368) <= not(layer3_outputs(2856));
    layer4_outputs(4369) <= not(layer3_outputs(4141)) or (layer3_outputs(130));
    layer4_outputs(4370) <= (layer3_outputs(2878)) and (layer3_outputs(6595));
    layer4_outputs(4371) <= not(layer3_outputs(6323));
    layer4_outputs(4372) <= not((layer3_outputs(7223)) and (layer3_outputs(6865)));
    layer4_outputs(4373) <= not(layer3_outputs(727));
    layer4_outputs(4374) <= (layer3_outputs(1471)) xor (layer3_outputs(4629));
    layer4_outputs(4375) <= (layer3_outputs(5027)) or (layer3_outputs(6008));
    layer4_outputs(4376) <= not(layer3_outputs(2153)) or (layer3_outputs(500));
    layer4_outputs(4377) <= not((layer3_outputs(4136)) xor (layer3_outputs(5100)));
    layer4_outputs(4378) <= (layer3_outputs(559)) and (layer3_outputs(3672));
    layer4_outputs(4379) <= not((layer3_outputs(6265)) or (layer3_outputs(5411)));
    layer4_outputs(4380) <= (layer3_outputs(7395)) xor (layer3_outputs(4695));
    layer4_outputs(4381) <= (layer3_outputs(1440)) and not (layer3_outputs(5360));
    layer4_outputs(4382) <= layer3_outputs(2217);
    layer4_outputs(4383) <= not(layer3_outputs(7466));
    layer4_outputs(4384) <= not(layer3_outputs(2514));
    layer4_outputs(4385) <= not((layer3_outputs(4361)) or (layer3_outputs(6693)));
    layer4_outputs(4386) <= not(layer3_outputs(1196));
    layer4_outputs(4387) <= not((layer3_outputs(1425)) or (layer3_outputs(6487)));
    layer4_outputs(4388) <= (layer3_outputs(2763)) and (layer3_outputs(2586));
    layer4_outputs(4389) <= not(layer3_outputs(1466));
    layer4_outputs(4390) <= not(layer3_outputs(1448)) or (layer3_outputs(7621));
    layer4_outputs(4391) <= not((layer3_outputs(3973)) and (layer3_outputs(1901)));
    layer4_outputs(4392) <= layer3_outputs(7368);
    layer4_outputs(4393) <= not((layer3_outputs(3769)) xor (layer3_outputs(4831)));
    layer4_outputs(4394) <= (layer3_outputs(4495)) or (layer3_outputs(2338));
    layer4_outputs(4395) <= layer3_outputs(513);
    layer4_outputs(4396) <= not(layer3_outputs(5941)) or (layer3_outputs(1101));
    layer4_outputs(4397) <= layer3_outputs(5803);
    layer4_outputs(4398) <= layer3_outputs(2895);
    layer4_outputs(4399) <= not((layer3_outputs(6789)) xor (layer3_outputs(1867)));
    layer4_outputs(4400) <= not((layer3_outputs(5603)) or (layer3_outputs(2842)));
    layer4_outputs(4401) <= not(layer3_outputs(6056)) or (layer3_outputs(269));
    layer4_outputs(4402) <= layer3_outputs(7124);
    layer4_outputs(4403) <= not(layer3_outputs(4183)) or (layer3_outputs(3116));
    layer4_outputs(4404) <= layer3_outputs(1704);
    layer4_outputs(4405) <= not(layer3_outputs(1710)) or (layer3_outputs(1595));
    layer4_outputs(4406) <= not((layer3_outputs(3806)) or (layer3_outputs(327)));
    layer4_outputs(4407) <= not((layer3_outputs(229)) or (layer3_outputs(7392)));
    layer4_outputs(4408) <= layer3_outputs(4779);
    layer4_outputs(4409) <= layer3_outputs(936);
    layer4_outputs(4410) <= not((layer3_outputs(5781)) xor (layer3_outputs(1010)));
    layer4_outputs(4411) <= not(layer3_outputs(3429));
    layer4_outputs(4412) <= not((layer3_outputs(7491)) xor (layer3_outputs(5394)));
    layer4_outputs(4413) <= not(layer3_outputs(1788));
    layer4_outputs(4414) <= not(layer3_outputs(3060));
    layer4_outputs(4415) <= not((layer3_outputs(7328)) or (layer3_outputs(7316)));
    layer4_outputs(4416) <= (layer3_outputs(4801)) and (layer3_outputs(3329));
    layer4_outputs(4417) <= not(layer3_outputs(4601)) or (layer3_outputs(2822));
    layer4_outputs(4418) <= not(layer3_outputs(4423));
    layer4_outputs(4419) <= not((layer3_outputs(1150)) or (layer3_outputs(6526)));
    layer4_outputs(4420) <= not(layer3_outputs(4812));
    layer4_outputs(4421) <= layer3_outputs(2428);
    layer4_outputs(4422) <= (layer3_outputs(3338)) and (layer3_outputs(2065));
    layer4_outputs(4423) <= not(layer3_outputs(3048));
    layer4_outputs(4424) <= not(layer3_outputs(4749));
    layer4_outputs(4425) <= layer3_outputs(3902);
    layer4_outputs(4426) <= not(layer3_outputs(3315));
    layer4_outputs(4427) <= layer3_outputs(6934);
    layer4_outputs(4428) <= (layer3_outputs(7118)) and not (layer3_outputs(2079));
    layer4_outputs(4429) <= not((layer3_outputs(3611)) and (layer3_outputs(4025)));
    layer4_outputs(4430) <= not((layer3_outputs(4333)) xor (layer3_outputs(834)));
    layer4_outputs(4431) <= layer3_outputs(2241);
    layer4_outputs(4432) <= layer3_outputs(4665);
    layer4_outputs(4433) <= not(layer3_outputs(2264));
    layer4_outputs(4434) <= layer3_outputs(7300);
    layer4_outputs(4435) <= layer3_outputs(6243);
    layer4_outputs(4436) <= not((layer3_outputs(6980)) xor (layer3_outputs(64)));
    layer4_outputs(4437) <= not(layer3_outputs(157));
    layer4_outputs(4438) <= not(layer3_outputs(3180));
    layer4_outputs(4439) <= not(layer3_outputs(6353));
    layer4_outputs(4440) <= (layer3_outputs(6286)) or (layer3_outputs(2111));
    layer4_outputs(4441) <= layer3_outputs(2761);
    layer4_outputs(4442) <= (layer3_outputs(4715)) and not (layer3_outputs(388));
    layer4_outputs(4443) <= layer3_outputs(4119);
    layer4_outputs(4444) <= (layer3_outputs(7240)) and not (layer3_outputs(5117));
    layer4_outputs(4445) <= not(layer3_outputs(4199));
    layer4_outputs(4446) <= not((layer3_outputs(6511)) and (layer3_outputs(3074)));
    layer4_outputs(4447) <= not(layer3_outputs(6811)) or (layer3_outputs(1541));
    layer4_outputs(4448) <= not(layer3_outputs(2799)) or (layer3_outputs(3387));
    layer4_outputs(4449) <= (layer3_outputs(3106)) and not (layer3_outputs(3872));
    layer4_outputs(4450) <= (layer3_outputs(7219)) or (layer3_outputs(3577));
    layer4_outputs(4451) <= (layer3_outputs(6060)) or (layer3_outputs(7578));
    layer4_outputs(4452) <= (layer3_outputs(2657)) xor (layer3_outputs(4510));
    layer4_outputs(4453) <= not(layer3_outputs(1892));
    layer4_outputs(4454) <= layer3_outputs(6872);
    layer4_outputs(4455) <= layer3_outputs(4712);
    layer4_outputs(4456) <= not((layer3_outputs(1407)) or (layer3_outputs(5544)));
    layer4_outputs(4457) <= (layer3_outputs(87)) and (layer3_outputs(4857));
    layer4_outputs(4458) <= not((layer3_outputs(6320)) or (layer3_outputs(5030)));
    layer4_outputs(4459) <= not((layer3_outputs(3412)) and (layer3_outputs(4797)));
    layer4_outputs(4460) <= (layer3_outputs(2835)) or (layer3_outputs(330));
    layer4_outputs(4461) <= (layer3_outputs(7139)) or (layer3_outputs(3825));
    layer4_outputs(4462) <= not(layer3_outputs(4626));
    layer4_outputs(4463) <= not(layer3_outputs(3377));
    layer4_outputs(4464) <= not(layer3_outputs(600));
    layer4_outputs(4465) <= not((layer3_outputs(4032)) and (layer3_outputs(5190)));
    layer4_outputs(4466) <= not(layer3_outputs(4740));
    layer4_outputs(4467) <= not(layer3_outputs(3402));
    layer4_outputs(4468) <= not((layer3_outputs(2454)) or (layer3_outputs(1658)));
    layer4_outputs(4469) <= (layer3_outputs(4435)) and not (layer3_outputs(6779));
    layer4_outputs(4470) <= (layer3_outputs(295)) and (layer3_outputs(469));
    layer4_outputs(4471) <= not(layer3_outputs(7570));
    layer4_outputs(4472) <= layer3_outputs(7222);
    layer4_outputs(4473) <= not(layer3_outputs(4512));
    layer4_outputs(4474) <= (layer3_outputs(6083)) and (layer3_outputs(6264));
    layer4_outputs(4475) <= (layer3_outputs(3994)) xor (layer3_outputs(5121));
    layer4_outputs(4476) <= layer3_outputs(6184);
    layer4_outputs(4477) <= (layer3_outputs(843)) and not (layer3_outputs(2564));
    layer4_outputs(4478) <= (layer3_outputs(6958)) and (layer3_outputs(3007));
    layer4_outputs(4479) <= layer3_outputs(1492);
    layer4_outputs(4480) <= not(layer3_outputs(7132));
    layer4_outputs(4481) <= (layer3_outputs(4406)) xor (layer3_outputs(4034));
    layer4_outputs(4482) <= layer3_outputs(2189);
    layer4_outputs(4483) <= not((layer3_outputs(5229)) xor (layer3_outputs(436)));
    layer4_outputs(4484) <= not(layer3_outputs(6605));
    layer4_outputs(4485) <= layer3_outputs(3246);
    layer4_outputs(4486) <= not((layer3_outputs(964)) xor (layer3_outputs(3206)));
    layer4_outputs(4487) <= not(layer3_outputs(1015));
    layer4_outputs(4488) <= layer3_outputs(2098);
    layer4_outputs(4489) <= not((layer3_outputs(3962)) or (layer3_outputs(1089)));
    layer4_outputs(4490) <= not(layer3_outputs(2371));
    layer4_outputs(4491) <= not(layer3_outputs(4575));
    layer4_outputs(4492) <= not(layer3_outputs(6106)) or (layer3_outputs(3340));
    layer4_outputs(4493) <= not(layer3_outputs(5052));
    layer4_outputs(4494) <= (layer3_outputs(2964)) xor (layer3_outputs(7619));
    layer4_outputs(4495) <= not(layer3_outputs(5535));
    layer4_outputs(4496) <= not(layer3_outputs(6311)) or (layer3_outputs(3353));
    layer4_outputs(4497) <= not((layer3_outputs(5992)) and (layer3_outputs(1097)));
    layer4_outputs(4498) <= '0';
    layer4_outputs(4499) <= (layer3_outputs(1913)) and not (layer3_outputs(5882));
    layer4_outputs(4500) <= not(layer3_outputs(1372)) or (layer3_outputs(5836));
    layer4_outputs(4501) <= layer3_outputs(4838);
    layer4_outputs(4502) <= not(layer3_outputs(4943));
    layer4_outputs(4503) <= layer3_outputs(1105);
    layer4_outputs(4504) <= layer3_outputs(653);
    layer4_outputs(4505) <= not((layer3_outputs(7384)) xor (layer3_outputs(4917)));
    layer4_outputs(4506) <= not((layer3_outputs(4336)) or (layer3_outputs(5196)));
    layer4_outputs(4507) <= not((layer3_outputs(7305)) xor (layer3_outputs(3645)));
    layer4_outputs(4508) <= not((layer3_outputs(1289)) or (layer3_outputs(6753)));
    layer4_outputs(4509) <= (layer3_outputs(2104)) and not (layer3_outputs(602));
    layer4_outputs(4510) <= not((layer3_outputs(5063)) xor (layer3_outputs(5471)));
    layer4_outputs(4511) <= layer3_outputs(1700);
    layer4_outputs(4512) <= (layer3_outputs(6608)) and (layer3_outputs(4018));
    layer4_outputs(4513) <= not((layer3_outputs(5884)) xor (layer3_outputs(623)));
    layer4_outputs(4514) <= (layer3_outputs(2143)) and not (layer3_outputs(1371));
    layer4_outputs(4515) <= (layer3_outputs(3555)) and (layer3_outputs(4264));
    layer4_outputs(4516) <= (layer3_outputs(4597)) or (layer3_outputs(7103));
    layer4_outputs(4517) <= (layer3_outputs(6565)) xor (layer3_outputs(6099));
    layer4_outputs(4518) <= not(layer3_outputs(4294));
    layer4_outputs(4519) <= layer3_outputs(687);
    layer4_outputs(4520) <= not(layer3_outputs(7325)) or (layer3_outputs(145));
    layer4_outputs(4521) <= layer3_outputs(3638);
    layer4_outputs(4522) <= '0';
    layer4_outputs(4523) <= (layer3_outputs(2402)) and (layer3_outputs(5419));
    layer4_outputs(4524) <= (layer3_outputs(5815)) and not (layer3_outputs(3262));
    layer4_outputs(4525) <= layer3_outputs(23);
    layer4_outputs(4526) <= layer3_outputs(4508);
    layer4_outputs(4527) <= not((layer3_outputs(3111)) and (layer3_outputs(5943)));
    layer4_outputs(4528) <= not(layer3_outputs(5123));
    layer4_outputs(4529) <= not(layer3_outputs(1522));
    layer4_outputs(4530) <= layer3_outputs(1921);
    layer4_outputs(4531) <= not(layer3_outputs(3297));
    layer4_outputs(4532) <= layer3_outputs(447);
    layer4_outputs(4533) <= not(layer3_outputs(7679));
    layer4_outputs(4534) <= (layer3_outputs(4508)) and not (layer3_outputs(7559));
    layer4_outputs(4535) <= layer3_outputs(4120);
    layer4_outputs(4536) <= layer3_outputs(2399);
    layer4_outputs(4537) <= layer3_outputs(6096);
    layer4_outputs(4538) <= not(layer3_outputs(1686)) or (layer3_outputs(79));
    layer4_outputs(4539) <= not(layer3_outputs(2453));
    layer4_outputs(4540) <= layer3_outputs(440);
    layer4_outputs(4541) <= not(layer3_outputs(3929)) or (layer3_outputs(1402));
    layer4_outputs(4542) <= not(layer3_outputs(5742)) or (layer3_outputs(566));
    layer4_outputs(4543) <= '0';
    layer4_outputs(4544) <= not((layer3_outputs(2744)) xor (layer3_outputs(2366)));
    layer4_outputs(4545) <= not(layer3_outputs(5503));
    layer4_outputs(4546) <= not(layer3_outputs(1685)) or (layer3_outputs(7047));
    layer4_outputs(4547) <= layer3_outputs(1219);
    layer4_outputs(4548) <= not((layer3_outputs(7378)) or (layer3_outputs(1233)));
    layer4_outputs(4549) <= not((layer3_outputs(5607)) and (layer3_outputs(305)));
    layer4_outputs(4550) <= not(layer3_outputs(7370));
    layer4_outputs(4551) <= not(layer3_outputs(6548));
    layer4_outputs(4552) <= (layer3_outputs(1464)) and (layer3_outputs(6390));
    layer4_outputs(4553) <= layer3_outputs(147);
    layer4_outputs(4554) <= not(layer3_outputs(6381)) or (layer3_outputs(7451));
    layer4_outputs(4555) <= layer3_outputs(7142);
    layer4_outputs(4556) <= not((layer3_outputs(7344)) xor (layer3_outputs(6665)));
    layer4_outputs(4557) <= not(layer3_outputs(2871));
    layer4_outputs(4558) <= (layer3_outputs(5021)) xor (layer3_outputs(815));
    layer4_outputs(4559) <= layer3_outputs(7523);
    layer4_outputs(4560) <= not(layer3_outputs(3662));
    layer4_outputs(4561) <= layer3_outputs(2760);
    layer4_outputs(4562) <= not((layer3_outputs(3603)) or (layer3_outputs(2670)));
    layer4_outputs(4563) <= (layer3_outputs(3991)) and (layer3_outputs(6112));
    layer4_outputs(4564) <= not(layer3_outputs(4130));
    layer4_outputs(4565) <= layer3_outputs(2357);
    layer4_outputs(4566) <= not((layer3_outputs(2601)) and (layer3_outputs(1887)));
    layer4_outputs(4567) <= not(layer3_outputs(1646));
    layer4_outputs(4568) <= not(layer3_outputs(2079));
    layer4_outputs(4569) <= layer3_outputs(6998);
    layer4_outputs(4570) <= not(layer3_outputs(3248));
    layer4_outputs(4571) <= layer3_outputs(1129);
    layer4_outputs(4572) <= layer3_outputs(4523);
    layer4_outputs(4573) <= layer3_outputs(3801);
    layer4_outputs(4574) <= layer3_outputs(7673);
    layer4_outputs(4575) <= not(layer3_outputs(3043));
    layer4_outputs(4576) <= (layer3_outputs(7484)) and (layer3_outputs(502));
    layer4_outputs(4577) <= not(layer3_outputs(1227));
    layer4_outputs(4578) <= not((layer3_outputs(1876)) xor (layer3_outputs(4380)));
    layer4_outputs(4579) <= not(layer3_outputs(87));
    layer4_outputs(4580) <= not(layer3_outputs(5662));
    layer4_outputs(4581) <= (layer3_outputs(5245)) and (layer3_outputs(143));
    layer4_outputs(4582) <= layer3_outputs(4639);
    layer4_outputs(4583) <= not(layer3_outputs(6336));
    layer4_outputs(4584) <= not((layer3_outputs(6183)) xor (layer3_outputs(5685)));
    layer4_outputs(4585) <= (layer3_outputs(1900)) and not (layer3_outputs(4992));
    layer4_outputs(4586) <= not(layer3_outputs(7307)) or (layer3_outputs(3406));
    layer4_outputs(4587) <= layer3_outputs(1098);
    layer4_outputs(4588) <= layer3_outputs(81);
    layer4_outputs(4589) <= not(layer3_outputs(2303));
    layer4_outputs(4590) <= (layer3_outputs(4300)) and (layer3_outputs(26));
    layer4_outputs(4591) <= (layer3_outputs(701)) xor (layer3_outputs(7111));
    layer4_outputs(4592) <= (layer3_outputs(2733)) and (layer3_outputs(6855));
    layer4_outputs(4593) <= layer3_outputs(1787);
    layer4_outputs(4594) <= not((layer3_outputs(2442)) or (layer3_outputs(254)));
    layer4_outputs(4595) <= not(layer3_outputs(139)) or (layer3_outputs(5438));
    layer4_outputs(4596) <= '1';
    layer4_outputs(4597) <= not(layer3_outputs(3710));
    layer4_outputs(4598) <= not(layer3_outputs(2408));
    layer4_outputs(4599) <= layer3_outputs(3971);
    layer4_outputs(4600) <= layer3_outputs(5367);
    layer4_outputs(4601) <= not(layer3_outputs(7565));
    layer4_outputs(4602) <= not((layer3_outputs(3326)) or (layer3_outputs(6273)));
    layer4_outputs(4603) <= layer3_outputs(1598);
    layer4_outputs(4604) <= layer3_outputs(5765);
    layer4_outputs(4605) <= not(layer3_outputs(463)) or (layer3_outputs(2036));
    layer4_outputs(4606) <= not(layer3_outputs(7458)) or (layer3_outputs(7043));
    layer4_outputs(4607) <= layer3_outputs(524);
    layer4_outputs(4608) <= layer3_outputs(5119);
    layer4_outputs(4609) <= not((layer3_outputs(2269)) or (layer3_outputs(4016)));
    layer4_outputs(4610) <= not(layer3_outputs(6628));
    layer4_outputs(4611) <= not(layer3_outputs(2037)) or (layer3_outputs(403));
    layer4_outputs(4612) <= layer3_outputs(4225);
    layer4_outputs(4613) <= not(layer3_outputs(4908));
    layer4_outputs(4614) <= not(layer3_outputs(2872)) or (layer3_outputs(5347));
    layer4_outputs(4615) <= not(layer3_outputs(2868)) or (layer3_outputs(4279));
    layer4_outputs(4616) <= (layer3_outputs(3564)) or (layer3_outputs(3955));
    layer4_outputs(4617) <= (layer3_outputs(3131)) and not (layer3_outputs(3020));
    layer4_outputs(4618) <= not(layer3_outputs(6174));
    layer4_outputs(4619) <= layer3_outputs(2817);
    layer4_outputs(4620) <= not(layer3_outputs(6274));
    layer4_outputs(4621) <= not(layer3_outputs(5171));
    layer4_outputs(4622) <= not(layer3_outputs(5017));
    layer4_outputs(4623) <= (layer3_outputs(6957)) and not (layer3_outputs(3852));
    layer4_outputs(4624) <= (layer3_outputs(6331)) and not (layer3_outputs(6239));
    layer4_outputs(4625) <= not(layer3_outputs(928));
    layer4_outputs(4626) <= layer3_outputs(5429);
    layer4_outputs(4627) <= not(layer3_outputs(3086)) or (layer3_outputs(1185));
    layer4_outputs(4628) <= (layer3_outputs(4390)) xor (layer3_outputs(5825));
    layer4_outputs(4629) <= layer3_outputs(3682);
    layer4_outputs(4630) <= (layer3_outputs(6919)) and not (layer3_outputs(768));
    layer4_outputs(4631) <= not(layer3_outputs(2749)) or (layer3_outputs(4329));
    layer4_outputs(4632) <= not(layer3_outputs(6072));
    layer4_outputs(4633) <= not(layer3_outputs(4692));
    layer4_outputs(4634) <= not((layer3_outputs(7099)) or (layer3_outputs(5171)));
    layer4_outputs(4635) <= not(layer3_outputs(2946));
    layer4_outputs(4636) <= (layer3_outputs(4988)) xor (layer3_outputs(5703));
    layer4_outputs(4637) <= not(layer3_outputs(2118)) or (layer3_outputs(1820));
    layer4_outputs(4638) <= not(layer3_outputs(963));
    layer4_outputs(4639) <= layer3_outputs(7119);
    layer4_outputs(4640) <= (layer3_outputs(1845)) or (layer3_outputs(5843));
    layer4_outputs(4641) <= not(layer3_outputs(6200)) or (layer3_outputs(6127));
    layer4_outputs(4642) <= not((layer3_outputs(2099)) xor (layer3_outputs(4859)));
    layer4_outputs(4643) <= not(layer3_outputs(6063)) or (layer3_outputs(620));
    layer4_outputs(4644) <= not(layer3_outputs(3219));
    layer4_outputs(4645) <= layer3_outputs(4984);
    layer4_outputs(4646) <= layer3_outputs(4340);
    layer4_outputs(4647) <= not(layer3_outputs(1752)) or (layer3_outputs(2852));
    layer4_outputs(4648) <= not(layer3_outputs(7345));
    layer4_outputs(4649) <= '0';
    layer4_outputs(4650) <= not(layer3_outputs(6842)) or (layer3_outputs(520));
    layer4_outputs(4651) <= (layer3_outputs(4685)) or (layer3_outputs(6179));
    layer4_outputs(4652) <= layer3_outputs(7037);
    layer4_outputs(4653) <= layer3_outputs(2473);
    layer4_outputs(4654) <= layer3_outputs(5031);
    layer4_outputs(4655) <= not(layer3_outputs(1203));
    layer4_outputs(4656) <= not(layer3_outputs(2376)) or (layer3_outputs(5987));
    layer4_outputs(4657) <= (layer3_outputs(7519)) and (layer3_outputs(6904));
    layer4_outputs(4658) <= not(layer3_outputs(5305));
    layer4_outputs(4659) <= layer3_outputs(3979);
    layer4_outputs(4660) <= not(layer3_outputs(2328));
    layer4_outputs(4661) <= not(layer3_outputs(4788));
    layer4_outputs(4662) <= not(layer3_outputs(3627));
    layer4_outputs(4663) <= not(layer3_outputs(5567));
    layer4_outputs(4664) <= layer3_outputs(3380);
    layer4_outputs(4665) <= not(layer3_outputs(1396)) or (layer3_outputs(2113));
    layer4_outputs(4666) <= layer3_outputs(5592);
    layer4_outputs(4667) <= layer3_outputs(3790);
    layer4_outputs(4668) <= (layer3_outputs(7550)) and not (layer3_outputs(3177));
    layer4_outputs(4669) <= (layer3_outputs(4690)) xor (layer3_outputs(273));
    layer4_outputs(4670) <= (layer3_outputs(5122)) and not (layer3_outputs(4057));
    layer4_outputs(4671) <= not((layer3_outputs(1778)) or (layer3_outputs(6421)));
    layer4_outputs(4672) <= (layer3_outputs(1265)) xor (layer3_outputs(2254));
    layer4_outputs(4673) <= '1';
    layer4_outputs(4674) <= layer3_outputs(769);
    layer4_outputs(4675) <= layer3_outputs(5659);
    layer4_outputs(4676) <= not(layer3_outputs(2134));
    layer4_outputs(4677) <= not(layer3_outputs(6036)) or (layer3_outputs(5261));
    layer4_outputs(4678) <= (layer3_outputs(7517)) and (layer3_outputs(6672));
    layer4_outputs(4679) <= not(layer3_outputs(5735));
    layer4_outputs(4680) <= not(layer3_outputs(929)) or (layer3_outputs(3655));
    layer4_outputs(4681) <= layer3_outputs(1459);
    layer4_outputs(4682) <= (layer3_outputs(1450)) and not (layer3_outputs(6421));
    layer4_outputs(4683) <= layer3_outputs(6558);
    layer4_outputs(4684) <= not((layer3_outputs(1890)) xor (layer3_outputs(7510)));
    layer4_outputs(4685) <= (layer3_outputs(7594)) and not (layer3_outputs(996));
    layer4_outputs(4686) <= not((layer3_outputs(7156)) or (layer3_outputs(5284)));
    layer4_outputs(4687) <= not(layer3_outputs(3525));
    layer4_outputs(4688) <= not(layer3_outputs(6371)) or (layer3_outputs(3052));
    layer4_outputs(4689) <= (layer3_outputs(5430)) and (layer3_outputs(7278));
    layer4_outputs(4690) <= not(layer3_outputs(1384)) or (layer3_outputs(3548));
    layer4_outputs(4691) <= not(layer3_outputs(4385));
    layer4_outputs(4692) <= not(layer3_outputs(2553));
    layer4_outputs(4693) <= not(layer3_outputs(650));
    layer4_outputs(4694) <= (layer3_outputs(4335)) and (layer3_outputs(2089));
    layer4_outputs(4695) <= layer3_outputs(4644);
    layer4_outputs(4696) <= not((layer3_outputs(6277)) or (layer3_outputs(7461)));
    layer4_outputs(4697) <= not(layer3_outputs(697));
    layer4_outputs(4698) <= layer3_outputs(2664);
    layer4_outputs(4699) <= not(layer3_outputs(2801));
    layer4_outputs(4700) <= not(layer3_outputs(2424));
    layer4_outputs(4701) <= not(layer3_outputs(5806)) or (layer3_outputs(4279));
    layer4_outputs(4702) <= layer3_outputs(5441);
    layer4_outputs(4703) <= not(layer3_outputs(6654));
    layer4_outputs(4704) <= not(layer3_outputs(3401));
    layer4_outputs(4705) <= not(layer3_outputs(7078));
    layer4_outputs(4706) <= layer3_outputs(4994);
    layer4_outputs(4707) <= not((layer3_outputs(3177)) and (layer3_outputs(5694)));
    layer4_outputs(4708) <= (layer3_outputs(840)) and (layer3_outputs(5170));
    layer4_outputs(4709) <= layer3_outputs(2007);
    layer4_outputs(4710) <= not((layer3_outputs(4760)) and (layer3_outputs(2686)));
    layer4_outputs(4711) <= not(layer3_outputs(4173));
    layer4_outputs(4712) <= '1';
    layer4_outputs(4713) <= (layer3_outputs(2601)) or (layer3_outputs(7010));
    layer4_outputs(4714) <= not(layer3_outputs(6401));
    layer4_outputs(4715) <= (layer3_outputs(2097)) and not (layer3_outputs(1314));
    layer4_outputs(4716) <= (layer3_outputs(3998)) or (layer3_outputs(7282));
    layer4_outputs(4717) <= not(layer3_outputs(5739));
    layer4_outputs(4718) <= not(layer3_outputs(974)) or (layer3_outputs(555));
    layer4_outputs(4719) <= not(layer3_outputs(3899)) or (layer3_outputs(7370));
    layer4_outputs(4720) <= not(layer3_outputs(6371));
    layer4_outputs(4721) <= layer3_outputs(5737);
    layer4_outputs(4722) <= (layer3_outputs(6945)) or (layer3_outputs(4546));
    layer4_outputs(4723) <= (layer3_outputs(1188)) xor (layer3_outputs(1193));
    layer4_outputs(4724) <= not(layer3_outputs(7295));
    layer4_outputs(4725) <= layer3_outputs(6434);
    layer4_outputs(4726) <= not(layer3_outputs(4693));
    layer4_outputs(4727) <= not(layer3_outputs(3077)) or (layer3_outputs(531));
    layer4_outputs(4728) <= not(layer3_outputs(1729)) or (layer3_outputs(5470));
    layer4_outputs(4729) <= (layer3_outputs(2204)) xor (layer3_outputs(6595));
    layer4_outputs(4730) <= (layer3_outputs(1667)) and (layer3_outputs(4221));
    layer4_outputs(4731) <= not(layer3_outputs(4658)) or (layer3_outputs(5519));
    layer4_outputs(4732) <= not((layer3_outputs(1839)) xor (layer3_outputs(400)));
    layer4_outputs(4733) <= (layer3_outputs(1026)) and (layer3_outputs(5427));
    layer4_outputs(4734) <= not(layer3_outputs(5972));
    layer4_outputs(4735) <= not((layer3_outputs(3433)) xor (layer3_outputs(2123)));
    layer4_outputs(4736) <= (layer3_outputs(6410)) xor (layer3_outputs(4496));
    layer4_outputs(4737) <= layer3_outputs(2590);
    layer4_outputs(4738) <= not(layer3_outputs(3284));
    layer4_outputs(4739) <= not((layer3_outputs(7235)) or (layer3_outputs(1184)));
    layer4_outputs(4740) <= (layer3_outputs(959)) and not (layer3_outputs(784));
    layer4_outputs(4741) <= layer3_outputs(1937);
    layer4_outputs(4742) <= not(layer3_outputs(4897));
    layer4_outputs(4743) <= not((layer3_outputs(7491)) xor (layer3_outputs(4464)));
    layer4_outputs(4744) <= not(layer3_outputs(788));
    layer4_outputs(4745) <= layer3_outputs(5035);
    layer4_outputs(4746) <= not(layer3_outputs(1090));
    layer4_outputs(4747) <= not(layer3_outputs(5345));
    layer4_outputs(4748) <= layer3_outputs(6224);
    layer4_outputs(4749) <= not(layer3_outputs(68)) or (layer3_outputs(4595));
    layer4_outputs(4750) <= (layer3_outputs(7239)) xor (layer3_outputs(1860));
    layer4_outputs(4751) <= (layer3_outputs(3609)) or (layer3_outputs(4456));
    layer4_outputs(4752) <= not(layer3_outputs(2654));
    layer4_outputs(4753) <= not(layer3_outputs(579)) or (layer3_outputs(6034));
    layer4_outputs(4754) <= not(layer3_outputs(6804));
    layer4_outputs(4755) <= layer3_outputs(3601);
    layer4_outputs(4756) <= not(layer3_outputs(748));
    layer4_outputs(4757) <= not(layer3_outputs(6778));
    layer4_outputs(4758) <= layer3_outputs(6422);
    layer4_outputs(4759) <= (layer3_outputs(4290)) and not (layer3_outputs(1706));
    layer4_outputs(4760) <= not(layer3_outputs(6796));
    layer4_outputs(4761) <= not((layer3_outputs(3325)) xor (layer3_outputs(5166)));
    layer4_outputs(4762) <= (layer3_outputs(4442)) and not (layer3_outputs(1756));
    layer4_outputs(4763) <= not(layer3_outputs(2452)) or (layer3_outputs(4974));
    layer4_outputs(4764) <= not(layer3_outputs(4871));
    layer4_outputs(4765) <= not((layer3_outputs(128)) xor (layer3_outputs(53)));
    layer4_outputs(4766) <= not(layer3_outputs(1588));
    layer4_outputs(4767) <= not((layer3_outputs(6949)) or (layer3_outputs(3591)));
    layer4_outputs(4768) <= layer3_outputs(1545);
    layer4_outputs(4769) <= (layer3_outputs(3430)) and not (layer3_outputs(7019));
    layer4_outputs(4770) <= not(layer3_outputs(7389)) or (layer3_outputs(2162));
    layer4_outputs(4771) <= layer3_outputs(2635);
    layer4_outputs(4772) <= (layer3_outputs(6063)) and not (layer3_outputs(5252));
    layer4_outputs(4773) <= layer3_outputs(4516);
    layer4_outputs(4774) <= not(layer3_outputs(978)) or (layer3_outputs(2502));
    layer4_outputs(4775) <= not((layer3_outputs(195)) and (layer3_outputs(3543)));
    layer4_outputs(4776) <= (layer3_outputs(999)) or (layer3_outputs(6364));
    layer4_outputs(4777) <= (layer3_outputs(2400)) and (layer3_outputs(6734));
    layer4_outputs(4778) <= not(layer3_outputs(6811)) or (layer3_outputs(985));
    layer4_outputs(4779) <= layer3_outputs(3047);
    layer4_outputs(4780) <= not(layer3_outputs(866));
    layer4_outputs(4781) <= (layer3_outputs(4798)) and not (layer3_outputs(6642));
    layer4_outputs(4782) <= (layer3_outputs(7373)) and not (layer3_outputs(237));
    layer4_outputs(4783) <= not(layer3_outputs(387));
    layer4_outputs(4784) <= not(layer3_outputs(2740)) or (layer3_outputs(2203));
    layer4_outputs(4785) <= not(layer3_outputs(1581));
    layer4_outputs(4786) <= (layer3_outputs(6579)) or (layer3_outputs(2531));
    layer4_outputs(4787) <= layer3_outputs(5183);
    layer4_outputs(4788) <= not((layer3_outputs(3886)) xor (layer3_outputs(4451)));
    layer4_outputs(4789) <= (layer3_outputs(4703)) xor (layer3_outputs(297));
    layer4_outputs(4790) <= '0';
    layer4_outputs(4791) <= not(layer3_outputs(6146));
    layer4_outputs(4792) <= not(layer3_outputs(2791)) or (layer3_outputs(6));
    layer4_outputs(4793) <= '0';
    layer4_outputs(4794) <= not((layer3_outputs(384)) xor (layer3_outputs(3035)));
    layer4_outputs(4795) <= (layer3_outputs(4013)) or (layer3_outputs(2218));
    layer4_outputs(4796) <= layer3_outputs(1036);
    layer4_outputs(4797) <= (layer3_outputs(5594)) and not (layer3_outputs(7435));
    layer4_outputs(4798) <= layer3_outputs(7480);
    layer4_outputs(4799) <= not((layer3_outputs(3209)) xor (layer3_outputs(5874)));
    layer4_outputs(4800) <= (layer3_outputs(4959)) xor (layer3_outputs(1861));
    layer4_outputs(4801) <= not(layer3_outputs(4522));
    layer4_outputs(4802) <= (layer3_outputs(7437)) or (layer3_outputs(1062));
    layer4_outputs(4803) <= (layer3_outputs(181)) and (layer3_outputs(4862));
    layer4_outputs(4804) <= not((layer3_outputs(2242)) and (layer3_outputs(6238)));
    layer4_outputs(4805) <= not(layer3_outputs(1166));
    layer4_outputs(4806) <= not(layer3_outputs(7322));
    layer4_outputs(4807) <= layer3_outputs(2332);
    layer4_outputs(4808) <= not(layer3_outputs(676));
    layer4_outputs(4809) <= layer3_outputs(4707);
    layer4_outputs(4810) <= not(layer3_outputs(6213));
    layer4_outputs(4811) <= (layer3_outputs(7541)) or (layer3_outputs(91));
    layer4_outputs(4812) <= layer3_outputs(4810);
    layer4_outputs(4813) <= not(layer3_outputs(4674)) or (layer3_outputs(2617));
    layer4_outputs(4814) <= (layer3_outputs(3738)) xor (layer3_outputs(5403));
    layer4_outputs(4815) <= not((layer3_outputs(154)) and (layer3_outputs(2795)));
    layer4_outputs(4816) <= not((layer3_outputs(995)) or (layer3_outputs(1918)));
    layer4_outputs(4817) <= (layer3_outputs(2704)) and (layer3_outputs(736));
    layer4_outputs(4818) <= not(layer3_outputs(2177));
    layer4_outputs(4819) <= not(layer3_outputs(1976));
    layer4_outputs(4820) <= not(layer3_outputs(5738));
    layer4_outputs(4821) <= not(layer3_outputs(79));
    layer4_outputs(4822) <= not((layer3_outputs(5299)) and (layer3_outputs(6512)));
    layer4_outputs(4823) <= not((layer3_outputs(7422)) xor (layer3_outputs(4654)));
    layer4_outputs(4824) <= layer3_outputs(5179);
    layer4_outputs(4825) <= not(layer3_outputs(2190));
    layer4_outputs(4826) <= not(layer3_outputs(120)) or (layer3_outputs(4878));
    layer4_outputs(4827) <= not(layer3_outputs(5774));
    layer4_outputs(4828) <= not(layer3_outputs(2631));
    layer4_outputs(4829) <= not((layer3_outputs(1085)) or (layer3_outputs(5275)));
    layer4_outputs(4830) <= not(layer3_outputs(2937)) or (layer3_outputs(7291));
    layer4_outputs(4831) <= layer3_outputs(4813);
    layer4_outputs(4832) <= '1';
    layer4_outputs(4833) <= (layer3_outputs(473)) or (layer3_outputs(6109));
    layer4_outputs(4834) <= not(layer3_outputs(2650));
    layer4_outputs(4835) <= layer3_outputs(539);
    layer4_outputs(4836) <= not(layer3_outputs(538));
    layer4_outputs(4837) <= layer3_outputs(5159);
    layer4_outputs(4838) <= not(layer3_outputs(4198));
    layer4_outputs(4839) <= layer3_outputs(906);
    layer4_outputs(4840) <= layer3_outputs(3834);
    layer4_outputs(4841) <= not(layer3_outputs(4985)) or (layer3_outputs(1926));
    layer4_outputs(4842) <= layer3_outputs(220);
    layer4_outputs(4843) <= not(layer3_outputs(3496));
    layer4_outputs(4844) <= not(layer3_outputs(2539));
    layer4_outputs(4845) <= not(layer3_outputs(3437));
    layer4_outputs(4846) <= (layer3_outputs(6885)) xor (layer3_outputs(4043));
    layer4_outputs(4847) <= not(layer3_outputs(1015)) or (layer3_outputs(5333));
    layer4_outputs(4848) <= (layer3_outputs(3200)) xor (layer3_outputs(6410));
    layer4_outputs(4849) <= not((layer3_outputs(1309)) and (layer3_outputs(2409)));
    layer4_outputs(4850) <= (layer3_outputs(822)) xor (layer3_outputs(3158));
    layer4_outputs(4851) <= (layer3_outputs(567)) xor (layer3_outputs(6370));
    layer4_outputs(4852) <= not(layer3_outputs(47)) or (layer3_outputs(5293));
    layer4_outputs(4853) <= layer3_outputs(400);
    layer4_outputs(4854) <= '0';
    layer4_outputs(4855) <= not((layer3_outputs(1926)) xor (layer3_outputs(7464)));
    layer4_outputs(4856) <= layer3_outputs(2302);
    layer4_outputs(4857) <= layer3_outputs(2067);
    layer4_outputs(4858) <= (layer3_outputs(6658)) or (layer3_outputs(5295));
    layer4_outputs(4859) <= (layer3_outputs(5494)) or (layer3_outputs(6308));
    layer4_outputs(4860) <= not(layer3_outputs(5373)) or (layer3_outputs(3630));
    layer4_outputs(4861) <= layer3_outputs(6469);
    layer4_outputs(4862) <= layer3_outputs(4269);
    layer4_outputs(4863) <= not(layer3_outputs(7650)) or (layer3_outputs(1252));
    layer4_outputs(4864) <= not(layer3_outputs(6379));
    layer4_outputs(4865) <= not(layer3_outputs(1446));
    layer4_outputs(4866) <= not(layer3_outputs(2138));
    layer4_outputs(4867) <= not((layer3_outputs(4660)) and (layer3_outputs(7367)));
    layer4_outputs(4868) <= layer3_outputs(5014);
    layer4_outputs(4869) <= not(layer3_outputs(5092)) or (layer3_outputs(7130));
    layer4_outputs(4870) <= not(layer3_outputs(7500));
    layer4_outputs(4871) <= not(layer3_outputs(3779)) or (layer3_outputs(4289));
    layer4_outputs(4872) <= not((layer3_outputs(4688)) xor (layer3_outputs(4448)));
    layer4_outputs(4873) <= (layer3_outputs(6038)) and not (layer3_outputs(6515));
    layer4_outputs(4874) <= not(layer3_outputs(3545));
    layer4_outputs(4875) <= not(layer3_outputs(4237)) or (layer3_outputs(3907));
    layer4_outputs(4876) <= layer3_outputs(3608);
    layer4_outputs(4877) <= not((layer3_outputs(7405)) xor (layer3_outputs(4931)));
    layer4_outputs(4878) <= (layer3_outputs(1145)) and (layer3_outputs(7417));
    layer4_outputs(4879) <= not(layer3_outputs(329));
    layer4_outputs(4880) <= not((layer3_outputs(3854)) or (layer3_outputs(4618)));
    layer4_outputs(4881) <= not(layer3_outputs(5556));
    layer4_outputs(4882) <= not(layer3_outputs(4473));
    layer4_outputs(4883) <= not((layer3_outputs(1542)) and (layer3_outputs(4458)));
    layer4_outputs(4884) <= not(layer3_outputs(1120)) or (layer3_outputs(4364));
    layer4_outputs(4885) <= (layer3_outputs(2963)) xor (layer3_outputs(7535));
    layer4_outputs(4886) <= layer3_outputs(1157);
    layer4_outputs(4887) <= not(layer3_outputs(2589));
    layer4_outputs(4888) <= not(layer3_outputs(3620));
    layer4_outputs(4889) <= layer3_outputs(2787);
    layer4_outputs(4890) <= not(layer3_outputs(5715));
    layer4_outputs(4891) <= not((layer3_outputs(4200)) xor (layer3_outputs(5840)));
    layer4_outputs(4892) <= not(layer3_outputs(7046)) or (layer3_outputs(2012));
    layer4_outputs(4893) <= (layer3_outputs(4919)) and not (layer3_outputs(954));
    layer4_outputs(4894) <= not((layer3_outputs(4019)) or (layer3_outputs(5578)));
    layer4_outputs(4895) <= not(layer3_outputs(5291));
    layer4_outputs(4896) <= (layer3_outputs(4993)) or (layer3_outputs(7441));
    layer4_outputs(4897) <= not(layer3_outputs(4773));
    layer4_outputs(4898) <= not(layer3_outputs(2647));
    layer4_outputs(4899) <= not(layer3_outputs(2578));
    layer4_outputs(4900) <= layer3_outputs(4340);
    layer4_outputs(4901) <= not((layer3_outputs(2272)) or (layer3_outputs(3575)));
    layer4_outputs(4902) <= layer3_outputs(892);
    layer4_outputs(4903) <= layer3_outputs(6006);
    layer4_outputs(4904) <= (layer3_outputs(4576)) or (layer3_outputs(1516));
    layer4_outputs(4905) <= layer3_outputs(1945);
    layer4_outputs(4906) <= not((layer3_outputs(2769)) and (layer3_outputs(3708)));
    layer4_outputs(4907) <= layer3_outputs(3523);
    layer4_outputs(4908) <= not(layer3_outputs(711));
    layer4_outputs(4909) <= not((layer3_outputs(5893)) and (layer3_outputs(3062)));
    layer4_outputs(4910) <= not(layer3_outputs(3594)) or (layer3_outputs(4806));
    layer4_outputs(4911) <= not(layer3_outputs(1757));
    layer4_outputs(4912) <= (layer3_outputs(4628)) xor (layer3_outputs(7442));
    layer4_outputs(4913) <= layer3_outputs(1711);
    layer4_outputs(4914) <= not(layer3_outputs(6923));
    layer4_outputs(4915) <= layer3_outputs(6995);
    layer4_outputs(4916) <= not(layer3_outputs(5501));
    layer4_outputs(4917) <= not((layer3_outputs(5747)) or (layer3_outputs(3743)));
    layer4_outputs(4918) <= layer3_outputs(7467);
    layer4_outputs(4919) <= not(layer3_outputs(205));
    layer4_outputs(4920) <= layer3_outputs(4977);
    layer4_outputs(4921) <= layer3_outputs(1211);
    layer4_outputs(4922) <= '0';
    layer4_outputs(4923) <= not(layer3_outputs(20));
    layer4_outputs(4924) <= not((layer3_outputs(1162)) or (layer3_outputs(5109)));
    layer4_outputs(4925) <= not(layer3_outputs(5470));
    layer4_outputs(4926) <= layer3_outputs(815);
    layer4_outputs(4927) <= not(layer3_outputs(17));
    layer4_outputs(4928) <= not((layer3_outputs(6489)) xor (layer3_outputs(4282)));
    layer4_outputs(4929) <= not(layer3_outputs(1581));
    layer4_outputs(4930) <= not((layer3_outputs(3492)) xor (layer3_outputs(119)));
    layer4_outputs(4931) <= layer3_outputs(5887);
    layer4_outputs(4932) <= not(layer3_outputs(2019));
    layer4_outputs(4933) <= (layer3_outputs(4480)) and not (layer3_outputs(5512));
    layer4_outputs(4934) <= layer3_outputs(2824);
    layer4_outputs(4935) <= layer3_outputs(86);
    layer4_outputs(4936) <= not((layer3_outputs(2173)) or (layer3_outputs(2046)));
    layer4_outputs(4937) <= not(layer3_outputs(6549));
    layer4_outputs(4938) <= not(layer3_outputs(2444));
    layer4_outputs(4939) <= not(layer3_outputs(3231));
    layer4_outputs(4940) <= not((layer3_outputs(6394)) xor (layer3_outputs(7132)));
    layer4_outputs(4941) <= (layer3_outputs(4976)) and not (layer3_outputs(346));
    layer4_outputs(4942) <= (layer3_outputs(7047)) and (layer3_outputs(3242));
    layer4_outputs(4943) <= layer3_outputs(6786);
    layer4_outputs(4944) <= layer3_outputs(4267);
    layer4_outputs(4945) <= (layer3_outputs(7409)) and not (layer3_outputs(1866));
    layer4_outputs(4946) <= layer3_outputs(5593);
    layer4_outputs(4947) <= layer3_outputs(5921);
    layer4_outputs(4948) <= (layer3_outputs(5960)) and (layer3_outputs(611));
    layer4_outputs(4949) <= (layer3_outputs(3420)) and not (layer3_outputs(7243));
    layer4_outputs(4950) <= (layer3_outputs(4857)) or (layer3_outputs(3251));
    layer4_outputs(4951) <= layer3_outputs(4580);
    layer4_outputs(4952) <= not(layer3_outputs(36));
    layer4_outputs(4953) <= (layer3_outputs(2360)) and (layer3_outputs(2152));
    layer4_outputs(4954) <= not((layer3_outputs(2286)) xor (layer3_outputs(2875)));
    layer4_outputs(4955) <= layer3_outputs(2043);
    layer4_outputs(4956) <= not(layer3_outputs(1362));
    layer4_outputs(4957) <= layer3_outputs(6384);
    layer4_outputs(4958) <= (layer3_outputs(3807)) or (layer3_outputs(2914));
    layer4_outputs(4959) <= (layer3_outputs(3516)) and not (layer3_outputs(3786));
    layer4_outputs(4960) <= layer3_outputs(3264);
    layer4_outputs(4961) <= not(layer3_outputs(6189)) or (layer3_outputs(420));
    layer4_outputs(4962) <= not((layer3_outputs(1555)) xor (layer3_outputs(1113)));
    layer4_outputs(4963) <= layer3_outputs(4842);
    layer4_outputs(4964) <= not((layer3_outputs(4752)) xor (layer3_outputs(2907)));
    layer4_outputs(4965) <= not(layer3_outputs(2293));
    layer4_outputs(4966) <= layer3_outputs(2893);
    layer4_outputs(4967) <= (layer3_outputs(7175)) xor (layer3_outputs(4584));
    layer4_outputs(4968) <= not(layer3_outputs(4926));
    layer4_outputs(4969) <= layer3_outputs(963);
    layer4_outputs(4970) <= layer3_outputs(390);
    layer4_outputs(4971) <= layer3_outputs(7016);
    layer4_outputs(4972) <= (layer3_outputs(7231)) and not (layer3_outputs(3408));
    layer4_outputs(4973) <= layer3_outputs(305);
    layer4_outputs(4974) <= not(layer3_outputs(4774));
    layer4_outputs(4975) <= not(layer3_outputs(5614));
    layer4_outputs(4976) <= layer3_outputs(4165);
    layer4_outputs(4977) <= not(layer3_outputs(1953));
    layer4_outputs(4978) <= (layer3_outputs(2721)) and (layer3_outputs(560));
    layer4_outputs(4979) <= not(layer3_outputs(5975));
    layer4_outputs(4980) <= (layer3_outputs(4963)) xor (layer3_outputs(1109));
    layer4_outputs(4981) <= layer3_outputs(1733);
    layer4_outputs(4982) <= not(layer3_outputs(4276));
    layer4_outputs(4983) <= layer3_outputs(170);
    layer4_outputs(4984) <= (layer3_outputs(2827)) and not (layer3_outputs(258));
    layer4_outputs(4985) <= (layer3_outputs(5530)) or (layer3_outputs(5495));
    layer4_outputs(4986) <= (layer3_outputs(7416)) or (layer3_outputs(6125));
    layer4_outputs(4987) <= (layer3_outputs(5248)) or (layer3_outputs(1933));
    layer4_outputs(4988) <= not(layer3_outputs(462));
    layer4_outputs(4989) <= '0';
    layer4_outputs(4990) <= not(layer3_outputs(954));
    layer4_outputs(4991) <= not(layer3_outputs(2834));
    layer4_outputs(4992) <= layer3_outputs(2312);
    layer4_outputs(4993) <= not(layer3_outputs(4500));
    layer4_outputs(4994) <= not((layer3_outputs(1562)) xor (layer3_outputs(5980)));
    layer4_outputs(4995) <= not(layer3_outputs(5145)) or (layer3_outputs(6139));
    layer4_outputs(4996) <= (layer3_outputs(3204)) xor (layer3_outputs(7629));
    layer4_outputs(4997) <= not(layer3_outputs(5240));
    layer4_outputs(4998) <= not(layer3_outputs(2341));
    layer4_outputs(4999) <= not(layer3_outputs(1344));
    layer4_outputs(5000) <= layer3_outputs(1080);
    layer4_outputs(5001) <= not(layer3_outputs(3963));
    layer4_outputs(5002) <= (layer3_outputs(7581)) and not (layer3_outputs(5463));
    layer4_outputs(5003) <= (layer3_outputs(6591)) or (layer3_outputs(610));
    layer4_outputs(5004) <= not(layer3_outputs(3554));
    layer4_outputs(5005) <= layer3_outputs(4397);
    layer4_outputs(5006) <= layer3_outputs(1897);
    layer4_outputs(5007) <= not(layer3_outputs(2334)) or (layer3_outputs(694));
    layer4_outputs(5008) <= not(layer3_outputs(2235));
    layer4_outputs(5009) <= layer3_outputs(4786);
    layer4_outputs(5010) <= '1';
    layer4_outputs(5011) <= not(layer3_outputs(2522)) or (layer3_outputs(636));
    layer4_outputs(5012) <= not(layer3_outputs(585));
    layer4_outputs(5013) <= not((layer3_outputs(5272)) xor (layer3_outputs(7608)));
    layer4_outputs(5014) <= not((layer3_outputs(7558)) and (layer3_outputs(4235)));
    layer4_outputs(5015) <= not(layer3_outputs(6476)) or (layer3_outputs(4442));
    layer4_outputs(5016) <= not((layer3_outputs(4266)) or (layer3_outputs(1805)));
    layer4_outputs(5017) <= not(layer3_outputs(6126));
    layer4_outputs(5018) <= not(layer3_outputs(6521));
    layer4_outputs(5019) <= not((layer3_outputs(5228)) or (layer3_outputs(4197)));
    layer4_outputs(5020) <= not(layer3_outputs(7533));
    layer4_outputs(5021) <= (layer3_outputs(4615)) and not (layer3_outputs(7216));
    layer4_outputs(5022) <= layer3_outputs(3747);
    layer4_outputs(5023) <= (layer3_outputs(4150)) or (layer3_outputs(4999));
    layer4_outputs(5024) <= (layer3_outputs(7575)) xor (layer3_outputs(44));
    layer4_outputs(5025) <= not((layer3_outputs(6468)) xor (layer3_outputs(4076)));
    layer4_outputs(5026) <= not(layer3_outputs(2638));
    layer4_outputs(5027) <= layer3_outputs(7608);
    layer4_outputs(5028) <= not(layer3_outputs(5189));
    layer4_outputs(5029) <= not((layer3_outputs(782)) or (layer3_outputs(448)));
    layer4_outputs(5030) <= layer3_outputs(6941);
    layer4_outputs(5031) <= not(layer3_outputs(2828)) or (layer3_outputs(7525));
    layer4_outputs(5032) <= (layer3_outputs(6437)) xor (layer3_outputs(4760));
    layer4_outputs(5033) <= not((layer3_outputs(7425)) or (layer3_outputs(5685)));
    layer4_outputs(5034) <= not(layer3_outputs(6075));
    layer4_outputs(5035) <= not(layer3_outputs(5385)) or (layer3_outputs(5562));
    layer4_outputs(5036) <= layer3_outputs(5009);
    layer4_outputs(5037) <= layer3_outputs(5247);
    layer4_outputs(5038) <= not(layer3_outputs(192));
    layer4_outputs(5039) <= '1';
    layer4_outputs(5040) <= not(layer3_outputs(2619));
    layer4_outputs(5041) <= layer3_outputs(4293);
    layer4_outputs(5042) <= layer3_outputs(4957);
    layer4_outputs(5043) <= (layer3_outputs(7483)) or (layer3_outputs(4116));
    layer4_outputs(5044) <= (layer3_outputs(921)) and (layer3_outputs(4652));
    layer4_outputs(5045) <= not(layer3_outputs(3805));
    layer4_outputs(5046) <= not(layer3_outputs(3903));
    layer4_outputs(5047) <= not(layer3_outputs(1985));
    layer4_outputs(5048) <= (layer3_outputs(3411)) and not (layer3_outputs(108));
    layer4_outputs(5049) <= not((layer3_outputs(312)) and (layer3_outputs(464)));
    layer4_outputs(5050) <= (layer3_outputs(5227)) and (layer3_outputs(1631));
    layer4_outputs(5051) <= not(layer3_outputs(6660));
    layer4_outputs(5052) <= layer3_outputs(2137);
    layer4_outputs(5053) <= not(layer3_outputs(3922));
    layer4_outputs(5054) <= layer3_outputs(7551);
    layer4_outputs(5055) <= layer3_outputs(1994);
    layer4_outputs(5056) <= not(layer3_outputs(6253));
    layer4_outputs(5057) <= not((layer3_outputs(6879)) and (layer3_outputs(5794)));
    layer4_outputs(5058) <= layer3_outputs(4077);
    layer4_outputs(5059) <= not((layer3_outputs(3032)) or (layer3_outputs(3132)));
    layer4_outputs(5060) <= (layer3_outputs(5829)) xor (layer3_outputs(1230));
    layer4_outputs(5061) <= layer3_outputs(3123);
    layer4_outputs(5062) <= not(layer3_outputs(6079));
    layer4_outputs(5063) <= not(layer3_outputs(1584));
    layer4_outputs(5064) <= layer3_outputs(465);
    layer4_outputs(5065) <= (layer3_outputs(7376)) and (layer3_outputs(4666));
    layer4_outputs(5066) <= layer3_outputs(513);
    layer4_outputs(5067) <= layer3_outputs(3155);
    layer4_outputs(5068) <= layer3_outputs(4238);
    layer4_outputs(5069) <= not((layer3_outputs(2848)) xor (layer3_outputs(1850)));
    layer4_outputs(5070) <= not(layer3_outputs(136));
    layer4_outputs(5071) <= layer3_outputs(302);
    layer4_outputs(5072) <= not(layer3_outputs(7495));
    layer4_outputs(5073) <= layer3_outputs(2950);
    layer4_outputs(5074) <= layer3_outputs(2003);
    layer4_outputs(5075) <= (layer3_outputs(5108)) or (layer3_outputs(2646));
    layer4_outputs(5076) <= not(layer3_outputs(5473));
    layer4_outputs(5077) <= not(layer3_outputs(4805));
    layer4_outputs(5078) <= (layer3_outputs(2523)) xor (layer3_outputs(3748));
    layer4_outputs(5079) <= (layer3_outputs(7276)) or (layer3_outputs(7612));
    layer4_outputs(5080) <= not(layer3_outputs(2168));
    layer4_outputs(5081) <= layer3_outputs(2396);
    layer4_outputs(5082) <= not(layer3_outputs(2978)) or (layer3_outputs(6054));
    layer4_outputs(5083) <= not(layer3_outputs(5961));
    layer4_outputs(5084) <= (layer3_outputs(7648)) and not (layer3_outputs(7085));
    layer4_outputs(5085) <= not(layer3_outputs(3588)) or (layer3_outputs(7472));
    layer4_outputs(5086) <= not((layer3_outputs(4562)) and (layer3_outputs(3553)));
    layer4_outputs(5087) <= not((layer3_outputs(1221)) or (layer3_outputs(6915)));
    layer4_outputs(5088) <= not(layer3_outputs(5682));
    layer4_outputs(5089) <= not(layer3_outputs(7277));
    layer4_outputs(5090) <= (layer3_outputs(7126)) and not (layer3_outputs(2396));
    layer4_outputs(5091) <= not(layer3_outputs(7003));
    layer4_outputs(5092) <= layer3_outputs(4414);
    layer4_outputs(5093) <= (layer3_outputs(6808)) and not (layer3_outputs(5764));
    layer4_outputs(5094) <= not(layer3_outputs(6525));
    layer4_outputs(5095) <= layer3_outputs(1808);
    layer4_outputs(5096) <= layer3_outputs(1751);
    layer4_outputs(5097) <= (layer3_outputs(6026)) and not (layer3_outputs(4894));
    layer4_outputs(5098) <= layer3_outputs(5367);
    layer4_outputs(5099) <= '1';
    layer4_outputs(5100) <= layer3_outputs(4587);
    layer4_outputs(5101) <= not((layer3_outputs(1394)) and (layer3_outputs(3584)));
    layer4_outputs(5102) <= (layer3_outputs(3201)) and not (layer3_outputs(6166));
    layer4_outputs(5103) <= (layer3_outputs(1281)) and not (layer3_outputs(498));
    layer4_outputs(5104) <= not(layer3_outputs(6326));
    layer4_outputs(5105) <= layer3_outputs(3103);
    layer4_outputs(5106) <= layer3_outputs(2862);
    layer4_outputs(5107) <= not(layer3_outputs(5669));
    layer4_outputs(5108) <= (layer3_outputs(631)) and not (layer3_outputs(1693));
    layer4_outputs(5109) <= layer3_outputs(5114);
    layer4_outputs(5110) <= (layer3_outputs(4735)) and not (layer3_outputs(7357));
    layer4_outputs(5111) <= layer3_outputs(2527);
    layer4_outputs(5112) <= (layer3_outputs(7671)) xor (layer3_outputs(7336));
    layer4_outputs(5113) <= layer3_outputs(913);
    layer4_outputs(5114) <= not(layer3_outputs(4336)) or (layer3_outputs(6756));
    layer4_outputs(5115) <= not(layer3_outputs(5154)) or (layer3_outputs(2465));
    layer4_outputs(5116) <= layer3_outputs(5184);
    layer4_outputs(5117) <= not((layer3_outputs(124)) and (layer3_outputs(7401)));
    layer4_outputs(5118) <= layer3_outputs(5654);
    layer4_outputs(5119) <= not(layer3_outputs(3309));
    layer4_outputs(5120) <= (layer3_outputs(7576)) xor (layer3_outputs(7301));
    layer4_outputs(5121) <= not(layer3_outputs(1587));
    layer4_outputs(5122) <= not((layer3_outputs(3810)) xor (layer3_outputs(4083)));
    layer4_outputs(5123) <= layer3_outputs(2995);
    layer4_outputs(5124) <= not((layer3_outputs(5716)) and (layer3_outputs(2538)));
    layer4_outputs(5125) <= not((layer3_outputs(736)) xor (layer3_outputs(4940)));
    layer4_outputs(5126) <= not(layer3_outputs(4603));
    layer4_outputs(5127) <= (layer3_outputs(5033)) xor (layer3_outputs(3978));
    layer4_outputs(5128) <= (layer3_outputs(1672)) and not (layer3_outputs(2998));
    layer4_outputs(5129) <= not(layer3_outputs(2184));
    layer4_outputs(5130) <= layer3_outputs(4641);
    layer4_outputs(5131) <= (layer3_outputs(5731)) and (layer3_outputs(2533));
    layer4_outputs(5132) <= not(layer3_outputs(5753));
    layer4_outputs(5133) <= layer3_outputs(5424);
    layer4_outputs(5134) <= not((layer3_outputs(196)) and (layer3_outputs(540)));
    layer4_outputs(5135) <= (layer3_outputs(5223)) xor (layer3_outputs(260));
    layer4_outputs(5136) <= not((layer3_outputs(2547)) xor (layer3_outputs(6840)));
    layer4_outputs(5137) <= not(layer3_outputs(7182));
    layer4_outputs(5138) <= not((layer3_outputs(1606)) or (layer3_outputs(1249)));
    layer4_outputs(5139) <= not(layer3_outputs(5750));
    layer4_outputs(5140) <= not(layer3_outputs(3097));
    layer4_outputs(5141) <= layer3_outputs(4650);
    layer4_outputs(5142) <= layer3_outputs(6217);
    layer4_outputs(5143) <= not((layer3_outputs(3003)) or (layer3_outputs(1663)));
    layer4_outputs(5144) <= (layer3_outputs(2027)) and not (layer3_outputs(5418));
    layer4_outputs(5145) <= layer3_outputs(3015);
    layer4_outputs(5146) <= not(layer3_outputs(7319));
    layer4_outputs(5147) <= (layer3_outputs(1814)) and not (layer3_outputs(303));
    layer4_outputs(5148) <= not((layer3_outputs(1071)) or (layer3_outputs(2058)));
    layer4_outputs(5149) <= layer3_outputs(2868);
    layer4_outputs(5150) <= (layer3_outputs(5358)) or (layer3_outputs(4485));
    layer4_outputs(5151) <= (layer3_outputs(3726)) and not (layer3_outputs(7548));
    layer4_outputs(5152) <= layer3_outputs(4635);
    layer4_outputs(5153) <= layer3_outputs(2234);
    layer4_outputs(5154) <= (layer3_outputs(1068)) and (layer3_outputs(2974));
    layer4_outputs(5155) <= (layer3_outputs(6642)) and not (layer3_outputs(6615));
    layer4_outputs(5156) <= not(layer3_outputs(2482));
    layer4_outputs(5157) <= (layer3_outputs(1242)) and (layer3_outputs(6080));
    layer4_outputs(5158) <= not(layer3_outputs(7582));
    layer4_outputs(5159) <= (layer3_outputs(7622)) or (layer3_outputs(3547));
    layer4_outputs(5160) <= not((layer3_outputs(2158)) or (layer3_outputs(460)));
    layer4_outputs(5161) <= (layer3_outputs(543)) or (layer3_outputs(5201));
    layer4_outputs(5162) <= layer3_outputs(3403);
    layer4_outputs(5163) <= layer3_outputs(6856);
    layer4_outputs(5164) <= (layer3_outputs(2973)) and not (layer3_outputs(6331));
    layer4_outputs(5165) <= layer3_outputs(923);
    layer4_outputs(5166) <= layer3_outputs(1909);
    layer4_outputs(5167) <= not(layer3_outputs(5044)) or (layer3_outputs(3484));
    layer4_outputs(5168) <= layer3_outputs(4388);
    layer4_outputs(5169) <= layer3_outputs(1676);
    layer4_outputs(5170) <= not(layer3_outputs(1608));
    layer4_outputs(5171) <= not(layer3_outputs(5210));
    layer4_outputs(5172) <= not(layer3_outputs(2630));
    layer4_outputs(5173) <= layer3_outputs(2361);
    layer4_outputs(5174) <= (layer3_outputs(482)) and (layer3_outputs(5724));
    layer4_outputs(5175) <= not(layer3_outputs(4940)) or (layer3_outputs(7003));
    layer4_outputs(5176) <= layer3_outputs(1505);
    layer4_outputs(5177) <= not(layer3_outputs(1004));
    layer4_outputs(5178) <= (layer3_outputs(1331)) and not (layer3_outputs(775));
    layer4_outputs(5179) <= layer3_outputs(3265);
    layer4_outputs(5180) <= (layer3_outputs(5129)) or (layer3_outputs(6911));
    layer4_outputs(5181) <= layer3_outputs(7281);
    layer4_outputs(5182) <= not(layer3_outputs(7303)) or (layer3_outputs(6334));
    layer4_outputs(5183) <= (layer3_outputs(7146)) and (layer3_outputs(1972));
    layer4_outputs(5184) <= not(layer3_outputs(6977)) or (layer3_outputs(2602));
    layer4_outputs(5185) <= layer3_outputs(7153);
    layer4_outputs(5186) <= layer3_outputs(7407);
    layer4_outputs(5187) <= layer3_outputs(3725);
    layer4_outputs(5188) <= (layer3_outputs(7269)) and not (layer3_outputs(6047));
    layer4_outputs(5189) <= layer3_outputs(6015);
    layer4_outputs(5190) <= layer3_outputs(4525);
    layer4_outputs(5191) <= '0';
    layer4_outputs(5192) <= (layer3_outputs(3010)) xor (layer3_outputs(524));
    layer4_outputs(5193) <= (layer3_outputs(369)) or (layer3_outputs(5833));
    layer4_outputs(5194) <= not(layer3_outputs(6857));
    layer4_outputs(5195) <= not((layer3_outputs(4250)) or (layer3_outputs(644)));
    layer4_outputs(5196) <= not(layer3_outputs(6592)) or (layer3_outputs(3486));
    layer4_outputs(5197) <= layer3_outputs(5426);
    layer4_outputs(5198) <= layer3_outputs(992);
    layer4_outputs(5199) <= (layer3_outputs(2157)) or (layer3_outputs(501));
    layer4_outputs(5200) <= not(layer3_outputs(3935)) or (layer3_outputs(2466));
    layer4_outputs(5201) <= not(layer3_outputs(1498));
    layer4_outputs(5202) <= '0';
    layer4_outputs(5203) <= layer3_outputs(5762);
    layer4_outputs(5204) <= layer3_outputs(285);
    layer4_outputs(5205) <= not((layer3_outputs(5540)) xor (layer3_outputs(675)));
    layer4_outputs(5206) <= (layer3_outputs(1713)) and (layer3_outputs(2729));
    layer4_outputs(5207) <= not(layer3_outputs(5597));
    layer4_outputs(5208) <= not(layer3_outputs(5996)) or (layer3_outputs(1698));
    layer4_outputs(5209) <= not(layer3_outputs(6190));
    layer4_outputs(5210) <= not((layer3_outputs(4085)) and (layer3_outputs(5425)));
    layer4_outputs(5211) <= not((layer3_outputs(5869)) or (layer3_outputs(2183)));
    layer4_outputs(5212) <= (layer3_outputs(1878)) and (layer3_outputs(1942));
    layer4_outputs(5213) <= not(layer3_outputs(7421));
    layer4_outputs(5214) <= (layer3_outputs(1862)) and (layer3_outputs(2432));
    layer4_outputs(5215) <= (layer3_outputs(378)) xor (layer3_outputs(4124));
    layer4_outputs(5216) <= not((layer3_outputs(6848)) or (layer3_outputs(5888)));
    layer4_outputs(5217) <= layer3_outputs(6247);
    layer4_outputs(5218) <= layer3_outputs(7455);
    layer4_outputs(5219) <= not((layer3_outputs(6593)) xor (layer3_outputs(3540)));
    layer4_outputs(5220) <= layer3_outputs(3218);
    layer4_outputs(5221) <= not(layer3_outputs(5629));
    layer4_outputs(5222) <= '1';
    layer4_outputs(5223) <= (layer3_outputs(7120)) and not (layer3_outputs(3245));
    layer4_outputs(5224) <= not((layer3_outputs(3183)) or (layer3_outputs(1863)));
    layer4_outputs(5225) <= layer3_outputs(2364);
    layer4_outputs(5226) <= not(layer3_outputs(2820));
    layer4_outputs(5227) <= (layer3_outputs(5006)) xor (layer3_outputs(3085));
    layer4_outputs(5228) <= not(layer3_outputs(6030)) or (layer3_outputs(4771));
    layer4_outputs(5229) <= layer3_outputs(1284);
    layer4_outputs(5230) <= not(layer3_outputs(7079));
    layer4_outputs(5231) <= (layer3_outputs(5693)) xor (layer3_outputs(2256));
    layer4_outputs(5232) <= not(layer3_outputs(794));
    layer4_outputs(5233) <= layer3_outputs(4099);
    layer4_outputs(5234) <= not((layer3_outputs(1353)) xor (layer3_outputs(2593)));
    layer4_outputs(5235) <= layer3_outputs(4366);
    layer4_outputs(5236) <= layer3_outputs(404);
    layer4_outputs(5237) <= not((layer3_outputs(719)) xor (layer3_outputs(6264)));
    layer4_outputs(5238) <= (layer3_outputs(738)) xor (layer3_outputs(5398));
    layer4_outputs(5239) <= not(layer3_outputs(6842)) or (layer3_outputs(6181));
    layer4_outputs(5240) <= not(layer3_outputs(2772));
    layer4_outputs(5241) <= '0';
    layer4_outputs(5242) <= (layer3_outputs(5766)) and not (layer3_outputs(6059));
    layer4_outputs(5243) <= not(layer3_outputs(5384)) or (layer3_outputs(4566));
    layer4_outputs(5244) <= layer3_outputs(4387);
    layer4_outputs(5245) <= layer3_outputs(4866);
    layer4_outputs(5246) <= not(layer3_outputs(7194));
    layer4_outputs(5247) <= not(layer3_outputs(202));
    layer4_outputs(5248) <= not(layer3_outputs(5686));
    layer4_outputs(5249) <= layer3_outputs(4224);
    layer4_outputs(5250) <= not((layer3_outputs(3482)) or (layer3_outputs(1494)));
    layer4_outputs(5251) <= layer3_outputs(4345);
    layer4_outputs(5252) <= not((layer3_outputs(4078)) xor (layer3_outputs(1637)));
    layer4_outputs(5253) <= not(layer3_outputs(5993)) or (layer3_outputs(1197));
    layer4_outputs(5254) <= layer3_outputs(7632);
    layer4_outputs(5255) <= (layer3_outputs(6463)) and not (layer3_outputs(4181));
    layer4_outputs(5256) <= (layer3_outputs(2181)) and (layer3_outputs(2804));
    layer4_outputs(5257) <= not(layer3_outputs(1822)) or (layer3_outputs(2999));
    layer4_outputs(5258) <= layer3_outputs(3696);
    layer4_outputs(5259) <= layer3_outputs(5349);
    layer4_outputs(5260) <= layer3_outputs(6348);
    layer4_outputs(5261) <= not(layer3_outputs(1503));
    layer4_outputs(5262) <= not(layer3_outputs(4252)) or (layer3_outputs(6708));
    layer4_outputs(5263) <= layer3_outputs(3025);
    layer4_outputs(5264) <= not(layer3_outputs(6507));
    layer4_outputs(5265) <= (layer3_outputs(1697)) and not (layer3_outputs(7216));
    layer4_outputs(5266) <= layer3_outputs(335);
    layer4_outputs(5267) <= layer3_outputs(2921);
    layer4_outputs(5268) <= (layer3_outputs(2001)) or (layer3_outputs(6275));
    layer4_outputs(5269) <= (layer3_outputs(6674)) or (layer3_outputs(6005));
    layer4_outputs(5270) <= (layer3_outputs(6692)) and not (layer3_outputs(3095));
    layer4_outputs(5271) <= not(layer3_outputs(989));
    layer4_outputs(5272) <= (layer3_outputs(4445)) xor (layer3_outputs(6895));
    layer4_outputs(5273) <= not(layer3_outputs(3462));
    layer4_outputs(5274) <= layer3_outputs(2159);
    layer4_outputs(5275) <= (layer3_outputs(1081)) and (layer3_outputs(52));
    layer4_outputs(5276) <= layer3_outputs(4955);
    layer4_outputs(5277) <= layer3_outputs(4542);
    layer4_outputs(5278) <= '0';
    layer4_outputs(5279) <= not(layer3_outputs(5670));
    layer4_outputs(5280) <= (layer3_outputs(3239)) and not (layer3_outputs(1769));
    layer4_outputs(5281) <= not(layer3_outputs(2208));
    layer4_outputs(5282) <= (layer3_outputs(5191)) and (layer3_outputs(855));
    layer4_outputs(5283) <= (layer3_outputs(5061)) and (layer3_outputs(7490));
    layer4_outputs(5284) <= (layer3_outputs(3425)) xor (layer3_outputs(5193));
    layer4_outputs(5285) <= not(layer3_outputs(1849)) or (layer3_outputs(3412));
    layer4_outputs(5286) <= not(layer3_outputs(6898));
    layer4_outputs(5287) <= not((layer3_outputs(4142)) or (layer3_outputs(4789)));
    layer4_outputs(5288) <= layer3_outputs(4115);
    layer4_outputs(5289) <= not(layer3_outputs(5205));
    layer4_outputs(5290) <= layer3_outputs(7337);
    layer4_outputs(5291) <= (layer3_outputs(6742)) xor (layer3_outputs(238));
    layer4_outputs(5292) <= layer3_outputs(3078);
    layer4_outputs(5293) <= layer3_outputs(2594);
    layer4_outputs(5294) <= not((layer3_outputs(6193)) and (layer3_outputs(3303)));
    layer4_outputs(5295) <= not(layer3_outputs(5640));
    layer4_outputs(5296) <= (layer3_outputs(1197)) xor (layer3_outputs(2692));
    layer4_outputs(5297) <= layer3_outputs(474);
    layer4_outputs(5298) <= not(layer3_outputs(749));
    layer4_outputs(5299) <= not(layer3_outputs(6229));
    layer4_outputs(5300) <= (layer3_outputs(7475)) and (layer3_outputs(4728));
    layer4_outputs(5301) <= (layer3_outputs(3921)) or (layer3_outputs(4361));
    layer4_outputs(5302) <= not((layer3_outputs(2316)) xor (layer3_outputs(5235)));
    layer4_outputs(5303) <= not((layer3_outputs(3983)) or (layer3_outputs(6042)));
    layer4_outputs(5304) <= not(layer3_outputs(3223)) or (layer3_outputs(3769));
    layer4_outputs(5305) <= not(layer3_outputs(4843)) or (layer3_outputs(4988));
    layer4_outputs(5306) <= (layer3_outputs(1789)) and not (layer3_outputs(4570));
    layer4_outputs(5307) <= layer3_outputs(4515);
    layer4_outputs(5308) <= layer3_outputs(2492);
    layer4_outputs(5309) <= (layer3_outputs(4859)) and (layer3_outputs(2981));
    layer4_outputs(5310) <= (layer3_outputs(6078)) and not (layer3_outputs(5791));
    layer4_outputs(5311) <= not(layer3_outputs(5622)) or (layer3_outputs(582));
    layer4_outputs(5312) <= not(layer3_outputs(3023)) or (layer3_outputs(1225));
    layer4_outputs(5313) <= not(layer3_outputs(6498));
    layer4_outputs(5314) <= layer3_outputs(5913);
    layer4_outputs(5315) <= not(layer3_outputs(1641));
    layer4_outputs(5316) <= layer3_outputs(3020);
    layer4_outputs(5317) <= layer3_outputs(5170);
    layer4_outputs(5318) <= not(layer3_outputs(1517));
    layer4_outputs(5319) <= (layer3_outputs(184)) xor (layer3_outputs(2922));
    layer4_outputs(5320) <= not(layer3_outputs(1949));
    layer4_outputs(5321) <= layer3_outputs(3255);
    layer4_outputs(5322) <= not((layer3_outputs(1579)) xor (layer3_outputs(6531)));
    layer4_outputs(5323) <= (layer3_outputs(5697)) and not (layer3_outputs(1978));
    layer4_outputs(5324) <= not(layer3_outputs(1653));
    layer4_outputs(5325) <= (layer3_outputs(2773)) xor (layer3_outputs(6071));
    layer4_outputs(5326) <= layer3_outputs(7244);
    layer4_outputs(5327) <= not((layer3_outputs(2873)) and (layer3_outputs(7092)));
    layer4_outputs(5328) <= not((layer3_outputs(367)) and (layer3_outputs(5062)));
    layer4_outputs(5329) <= not(layer3_outputs(2955));
    layer4_outputs(5330) <= layer3_outputs(2385);
    layer4_outputs(5331) <= not(layer3_outputs(6927));
    layer4_outputs(5332) <= layer3_outputs(370);
    layer4_outputs(5333) <= not(layer3_outputs(5499)) or (layer3_outputs(163));
    layer4_outputs(5334) <= (layer3_outputs(3256)) and not (layer3_outputs(132));
    layer4_outputs(5335) <= not((layer3_outputs(7347)) or (layer3_outputs(3964)));
    layer4_outputs(5336) <= not(layer3_outputs(717));
    layer4_outputs(5337) <= not(layer3_outputs(5254)) or (layer3_outputs(3926));
    layer4_outputs(5338) <= layer3_outputs(1621);
    layer4_outputs(5339) <= (layer3_outputs(4295)) xor (layer3_outputs(3199));
    layer4_outputs(5340) <= layer3_outputs(2333);
    layer4_outputs(5341) <= not(layer3_outputs(3230));
    layer4_outputs(5342) <= not(layer3_outputs(4323));
    layer4_outputs(5343) <= not((layer3_outputs(6380)) xor (layer3_outputs(2869)));
    layer4_outputs(5344) <= not(layer3_outputs(1072));
    layer4_outputs(5345) <= layer3_outputs(4997);
    layer4_outputs(5346) <= layer3_outputs(2041);
    layer4_outputs(5347) <= not(layer3_outputs(4830));
    layer4_outputs(5348) <= layer3_outputs(6169);
    layer4_outputs(5349) <= not((layer3_outputs(2929)) or (layer3_outputs(2324)));
    layer4_outputs(5350) <= not((layer3_outputs(5782)) and (layer3_outputs(5602)));
    layer4_outputs(5351) <= not((layer3_outputs(5023)) and (layer3_outputs(6312)));
    layer4_outputs(5352) <= not((layer3_outputs(4254)) and (layer3_outputs(3650)));
    layer4_outputs(5353) <= layer3_outputs(3729);
    layer4_outputs(5354) <= layer3_outputs(990);
    layer4_outputs(5355) <= not((layer3_outputs(3740)) and (layer3_outputs(1964)));
    layer4_outputs(5356) <= layer3_outputs(2777);
    layer4_outputs(5357) <= not(layer3_outputs(3110));
    layer4_outputs(5358) <= layer3_outputs(6013);
    layer4_outputs(5359) <= layer3_outputs(1514);
    layer4_outputs(5360) <= not(layer3_outputs(2262)) or (layer3_outputs(1998));
    layer4_outputs(5361) <= not(layer3_outputs(5832));
    layer4_outputs(5362) <= not(layer3_outputs(2375)) or (layer3_outputs(5150));
    layer4_outputs(5363) <= not((layer3_outputs(163)) or (layer3_outputs(4153)));
    layer4_outputs(5364) <= layer3_outputs(2507);
    layer4_outputs(5365) <= not(layer3_outputs(96));
    layer4_outputs(5366) <= (layer3_outputs(5214)) and not (layer3_outputs(3034));
    layer4_outputs(5367) <= not(layer3_outputs(7235));
    layer4_outputs(5368) <= (layer3_outputs(1966)) and not (layer3_outputs(6386));
    layer4_outputs(5369) <= layer3_outputs(4322);
    layer4_outputs(5370) <= (layer3_outputs(2957)) and (layer3_outputs(1672));
    layer4_outputs(5371) <= not(layer3_outputs(3251));
    layer4_outputs(5372) <= not((layer3_outputs(4502)) or (layer3_outputs(3026)));
    layer4_outputs(5373) <= not(layer3_outputs(1734));
    layer4_outputs(5374) <= (layer3_outputs(4829)) xor (layer3_outputs(23));
    layer4_outputs(5375) <= layer3_outputs(1967);
    layer4_outputs(5376) <= not(layer3_outputs(1730));
    layer4_outputs(5377) <= not(layer3_outputs(281));
    layer4_outputs(5378) <= not(layer3_outputs(5790)) or (layer3_outputs(519));
    layer4_outputs(5379) <= layer3_outputs(7486);
    layer4_outputs(5380) <= not((layer3_outputs(3293)) or (layer3_outputs(5334)));
    layer4_outputs(5381) <= not(layer3_outputs(1933));
    layer4_outputs(5382) <= (layer3_outputs(2905)) xor (layer3_outputs(1104));
    layer4_outputs(5383) <= (layer3_outputs(1684)) or (layer3_outputs(3286));
    layer4_outputs(5384) <= (layer3_outputs(1776)) xor (layer3_outputs(7065));
    layer4_outputs(5385) <= (layer3_outputs(5688)) and (layer3_outputs(2813));
    layer4_outputs(5386) <= layer3_outputs(6885);
    layer4_outputs(5387) <= layer3_outputs(5539);
    layer4_outputs(5388) <= not(layer3_outputs(7080)) or (layer3_outputs(3641));
    layer4_outputs(5389) <= layer3_outputs(1275);
    layer4_outputs(5390) <= (layer3_outputs(1620)) or (layer3_outputs(5060));
    layer4_outputs(5391) <= not(layer3_outputs(2480));
    layer4_outputs(5392) <= (layer3_outputs(1897)) or (layer3_outputs(6851));
    layer4_outputs(5393) <= layer3_outputs(6918);
    layer4_outputs(5394) <= not((layer3_outputs(208)) and (layer3_outputs(3098)));
    layer4_outputs(5395) <= layer3_outputs(6445);
    layer4_outputs(5396) <= not(layer3_outputs(6844)) or (layer3_outputs(3074));
    layer4_outputs(5397) <= not((layer3_outputs(6271)) and (layer3_outputs(5089)));
    layer4_outputs(5398) <= not(layer3_outputs(2125));
    layer4_outputs(5399) <= layer3_outputs(2621);
    layer4_outputs(5400) <= (layer3_outputs(6462)) and (layer3_outputs(3563));
    layer4_outputs(5401) <= not(layer3_outputs(4968));
    layer4_outputs(5402) <= not(layer3_outputs(6341));
    layer4_outputs(5403) <= not(layer3_outputs(5154));
    layer4_outputs(5404) <= not(layer3_outputs(6077));
    layer4_outputs(5405) <= not(layer3_outputs(2759)) or (layer3_outputs(3597));
    layer4_outputs(5406) <= not((layer3_outputs(6067)) xor (layer3_outputs(1003)));
    layer4_outputs(5407) <= not(layer3_outputs(6159));
    layer4_outputs(5408) <= not(layer3_outputs(7198)) or (layer3_outputs(3165));
    layer4_outputs(5409) <= not((layer3_outputs(2821)) xor (layer3_outputs(3549)));
    layer4_outputs(5410) <= not(layer3_outputs(3651));
    layer4_outputs(5411) <= not((layer3_outputs(7071)) and (layer3_outputs(2672)));
    layer4_outputs(5412) <= (layer3_outputs(5581)) and not (layer3_outputs(1742));
    layer4_outputs(5413) <= not((layer3_outputs(153)) or (layer3_outputs(3970)));
    layer4_outputs(5414) <= not(layer3_outputs(427));
    layer4_outputs(5415) <= not(layer3_outputs(4829));
    layer4_outputs(5416) <= '0';
    layer4_outputs(5417) <= not((layer3_outputs(132)) xor (layer3_outputs(1313)));
    layer4_outputs(5418) <= not(layer3_outputs(6991));
    layer4_outputs(5419) <= (layer3_outputs(1501)) or (layer3_outputs(5684));
    layer4_outputs(5420) <= not(layer3_outputs(6951));
    layer4_outputs(5421) <= not(layer3_outputs(6483));
    layer4_outputs(5422) <= not(layer3_outputs(1649));
    layer4_outputs(5423) <= (layer3_outputs(4002)) and (layer3_outputs(3290));
    layer4_outputs(5424) <= (layer3_outputs(2117)) and not (layer3_outputs(261));
    layer4_outputs(5425) <= not(layer3_outputs(2716));
    layer4_outputs(5426) <= not(layer3_outputs(6698)) or (layer3_outputs(2629));
    layer4_outputs(5427) <= not(layer3_outputs(4875)) or (layer3_outputs(4133));
    layer4_outputs(5428) <= layer3_outputs(3013);
    layer4_outputs(5429) <= not((layer3_outputs(3763)) xor (layer3_outputs(184)));
    layer4_outputs(5430) <= not((layer3_outputs(3465)) or (layer3_outputs(6909)));
    layer4_outputs(5431) <= (layer3_outputs(3433)) or (layer3_outputs(4321));
    layer4_outputs(5432) <= not(layer3_outputs(5853));
    layer4_outputs(5433) <= '0';
    layer4_outputs(5434) <= not(layer3_outputs(6365));
    layer4_outputs(5435) <= not(layer3_outputs(3537));
    layer4_outputs(5436) <= layer3_outputs(4936);
    layer4_outputs(5437) <= not((layer3_outputs(3121)) and (layer3_outputs(868)));
    layer4_outputs(5438) <= (layer3_outputs(1250)) and not (layer3_outputs(6225));
    layer4_outputs(5439) <= not(layer3_outputs(5112));
    layer4_outputs(5440) <= not((layer3_outputs(6486)) or (layer3_outputs(7595)));
    layer4_outputs(5441) <= not(layer3_outputs(5133));
    layer4_outputs(5442) <= (layer3_outputs(3920)) and not (layer3_outputs(1293));
    layer4_outputs(5443) <= layer3_outputs(1018);
    layer4_outputs(5444) <= layer3_outputs(1456);
    layer4_outputs(5445) <= not((layer3_outputs(5801)) xor (layer3_outputs(5561)));
    layer4_outputs(5446) <= (layer3_outputs(4087)) and not (layer3_outputs(5250));
    layer4_outputs(5447) <= not(layer3_outputs(3687));
    layer4_outputs(5448) <= not(layer3_outputs(6418));
    layer4_outputs(5449) <= layer3_outputs(2975);
    layer4_outputs(5450) <= not((layer3_outputs(2092)) xor (layer3_outputs(5078)));
    layer4_outputs(5451) <= layer3_outputs(3148);
    layer4_outputs(5452) <= not((layer3_outputs(7048)) xor (layer3_outputs(5110)));
    layer4_outputs(5453) <= layer3_outputs(5212);
    layer4_outputs(5454) <= (layer3_outputs(6858)) and (layer3_outputs(7586));
    layer4_outputs(5455) <= (layer3_outputs(5618)) and not (layer3_outputs(7627));
    layer4_outputs(5456) <= not(layer3_outputs(7628)) or (layer3_outputs(2966));
    layer4_outputs(5457) <= not(layer3_outputs(3891));
    layer4_outputs(5458) <= (layer3_outputs(5861)) and (layer3_outputs(6170));
    layer4_outputs(5459) <= not((layer3_outputs(446)) xor (layer3_outputs(5941)));
    layer4_outputs(5460) <= (layer3_outputs(1220)) or (layer3_outputs(5983));
    layer4_outputs(5461) <= layer3_outputs(1346);
    layer4_outputs(5462) <= not(layer3_outputs(4520));
    layer4_outputs(5463) <= not(layer3_outputs(3864)) or (layer3_outputs(2212));
    layer4_outputs(5464) <= not(layer3_outputs(5276)) or (layer3_outputs(6818));
    layer4_outputs(5465) <= not(layer3_outputs(4624));
    layer4_outputs(5466) <= not(layer3_outputs(4726));
    layer4_outputs(5467) <= not(layer3_outputs(3961));
    layer4_outputs(5468) <= (layer3_outputs(3138)) xor (layer3_outputs(5818));
    layer4_outputs(5469) <= not(layer3_outputs(6579));
    layer4_outputs(5470) <= layer3_outputs(4930);
    layer4_outputs(5471) <= (layer3_outputs(5644)) or (layer3_outputs(5837));
    layer4_outputs(5472) <= '0';
    layer4_outputs(5473) <= not((layer3_outputs(1832)) and (layer3_outputs(3038)));
    layer4_outputs(5474) <= not((layer3_outputs(5669)) or (layer3_outputs(1523)));
    layer4_outputs(5475) <= not(layer3_outputs(2615));
    layer4_outputs(5476) <= not((layer3_outputs(1130)) or (layer3_outputs(5327)));
    layer4_outputs(5477) <= layer3_outputs(5314);
    layer4_outputs(5478) <= not(layer3_outputs(6342));
    layer4_outputs(5479) <= not(layer3_outputs(6964));
    layer4_outputs(5480) <= not(layer3_outputs(1722));
    layer4_outputs(5481) <= (layer3_outputs(1978)) or (layer3_outputs(5173));
    layer4_outputs(5482) <= (layer3_outputs(3342)) and (layer3_outputs(787));
    layer4_outputs(5483) <= not(layer3_outputs(4757)) or (layer3_outputs(3441));
    layer4_outputs(5484) <= not(layer3_outputs(6046)) or (layer3_outputs(670));
    layer4_outputs(5485) <= not(layer3_outputs(3617));
    layer4_outputs(5486) <= layer3_outputs(7329);
    layer4_outputs(5487) <= (layer3_outputs(1503)) and not (layer3_outputs(4359));
    layer4_outputs(5488) <= (layer3_outputs(3808)) and not (layer3_outputs(1228));
    layer4_outputs(5489) <= not((layer3_outputs(2416)) xor (layer3_outputs(1991)));
    layer4_outputs(5490) <= layer3_outputs(1428);
    layer4_outputs(5491) <= not(layer3_outputs(2100));
    layer4_outputs(5492) <= (layer3_outputs(5959)) and not (layer3_outputs(630));
    layer4_outputs(5493) <= not(layer3_outputs(4867)) or (layer3_outputs(4475));
    layer4_outputs(5494) <= (layer3_outputs(5797)) xor (layer3_outputs(6643));
    layer4_outputs(5495) <= layer3_outputs(1258);
    layer4_outputs(5496) <= layer3_outputs(6275);
    layer4_outputs(5497) <= layer3_outputs(7359);
    layer4_outputs(5498) <= not(layer3_outputs(2773)) or (layer3_outputs(7523));
    layer4_outputs(5499) <= layer3_outputs(2721);
    layer4_outputs(5500) <= layer3_outputs(4305);
    layer4_outputs(5501) <= (layer3_outputs(3027)) xor (layer3_outputs(5696));
    layer4_outputs(5502) <= (layer3_outputs(5749)) xor (layer3_outputs(6682));
    layer4_outputs(5503) <= layer3_outputs(1156);
    layer4_outputs(5504) <= not(layer3_outputs(4636));
    layer4_outputs(5505) <= (layer3_outputs(3505)) xor (layer3_outputs(2978));
    layer4_outputs(5506) <= not((layer3_outputs(486)) and (layer3_outputs(311)));
    layer4_outputs(5507) <= layer3_outputs(3631);
    layer4_outputs(5508) <= (layer3_outputs(4712)) or (layer3_outputs(140));
    layer4_outputs(5509) <= layer3_outputs(637);
    layer4_outputs(5510) <= (layer3_outputs(2543)) or (layer3_outputs(4925));
    layer4_outputs(5511) <= layer3_outputs(5828);
    layer4_outputs(5512) <= not(layer3_outputs(1474));
    layer4_outputs(5513) <= (layer3_outputs(1178)) and not (layer3_outputs(1509));
    layer4_outputs(5514) <= layer3_outputs(7397);
    layer4_outputs(5515) <= not(layer3_outputs(809));
    layer4_outputs(5516) <= (layer3_outputs(3322)) and not (layer3_outputs(290));
    layer4_outputs(5517) <= not(layer3_outputs(2221));
    layer4_outputs(5518) <= layer3_outputs(3239);
    layer4_outputs(5519) <= not(layer3_outputs(5569)) or (layer3_outputs(1654));
    layer4_outputs(5520) <= (layer3_outputs(6896)) or (layer3_outputs(4387));
    layer4_outputs(5521) <= (layer3_outputs(3167)) and (layer3_outputs(2213));
    layer4_outputs(5522) <= not((layer3_outputs(6600)) or (layer3_outputs(3864)));
    layer4_outputs(5523) <= layer3_outputs(4911);
    layer4_outputs(5524) <= layer3_outputs(5116);
    layer4_outputs(5525) <= (layer3_outputs(1573)) or (layer3_outputs(7603));
    layer4_outputs(5526) <= (layer3_outputs(124)) and (layer3_outputs(4861));
    layer4_outputs(5527) <= (layer3_outputs(3323)) and (layer3_outputs(2023));
    layer4_outputs(5528) <= not(layer3_outputs(2739));
    layer4_outputs(5529) <= layer3_outputs(1760);
    layer4_outputs(5530) <= (layer3_outputs(969)) and not (layer3_outputs(943));
    layer4_outputs(5531) <= (layer3_outputs(2732)) or (layer3_outputs(6360));
    layer4_outputs(5532) <= layer3_outputs(274);
    layer4_outputs(5533) <= not(layer3_outputs(1996));
    layer4_outputs(5534) <= not((layer3_outputs(5305)) and (layer3_outputs(2609)));
    layer4_outputs(5535) <= not(layer3_outputs(144));
    layer4_outputs(5536) <= not(layer3_outputs(32)) or (layer3_outputs(7456));
    layer4_outputs(5537) <= layer3_outputs(4345);
    layer4_outputs(5538) <= not((layer3_outputs(5723)) xor (layer3_outputs(2710)));
    layer4_outputs(5539) <= not((layer3_outputs(6290)) xor (layer3_outputs(1321)));
    layer4_outputs(5540) <= not((layer3_outputs(6748)) xor (layer3_outputs(4631)));
    layer4_outputs(5541) <= not(layer3_outputs(2934));
    layer4_outputs(5542) <= layer3_outputs(3259);
    layer4_outputs(5543) <= not(layer3_outputs(4204));
    layer4_outputs(5544) <= not(layer3_outputs(933));
    layer4_outputs(5545) <= not(layer3_outputs(1322)) or (layer3_outputs(6964));
    layer4_outputs(5546) <= not(layer3_outputs(3090));
    layer4_outputs(5547) <= layer3_outputs(1883);
    layer4_outputs(5548) <= layer3_outputs(3511);
    layer4_outputs(5549) <= not(layer3_outputs(2352));
    layer4_outputs(5550) <= (layer3_outputs(2520)) xor (layer3_outputs(1457));
    layer4_outputs(5551) <= not(layer3_outputs(2636));
    layer4_outputs(5552) <= not((layer3_outputs(2107)) or (layer3_outputs(3076)));
    layer4_outputs(5553) <= not(layer3_outputs(2103));
    layer4_outputs(5554) <= not(layer3_outputs(4320));
    layer4_outputs(5555) <= not(layer3_outputs(2741));
    layer4_outputs(5556) <= '1';
    layer4_outputs(5557) <= not(layer3_outputs(1215));
    layer4_outputs(5558) <= (layer3_outputs(7256)) xor (layer3_outputs(939));
    layer4_outputs(5559) <= (layer3_outputs(3543)) and (layer3_outputs(6369));
    layer4_outputs(5560) <= not(layer3_outputs(3028));
    layer4_outputs(5561) <= layer3_outputs(645);
    layer4_outputs(5562) <= not(layer3_outputs(2921));
    layer4_outputs(5563) <= layer3_outputs(1705);
    layer4_outputs(5564) <= not(layer3_outputs(7264));
    layer4_outputs(5565) <= layer3_outputs(5137);
    layer4_outputs(5566) <= layer3_outputs(1477);
    layer4_outputs(5567) <= not(layer3_outputs(6930)) or (layer3_outputs(4217));
    layer4_outputs(5568) <= not(layer3_outputs(1372)) or (layer3_outputs(901));
    layer4_outputs(5569) <= (layer3_outputs(7205)) and not (layer3_outputs(3793));
    layer4_outputs(5570) <= not(layer3_outputs(760));
    layer4_outputs(5571) <= not(layer3_outputs(5235));
    layer4_outputs(5572) <= (layer3_outputs(6352)) and (layer3_outputs(1354));
    layer4_outputs(5573) <= layer3_outputs(6110);
    layer4_outputs(5574) <= layer3_outputs(5979);
    layer4_outputs(5575) <= not((layer3_outputs(2210)) xor (layer3_outputs(1807)));
    layer4_outputs(5576) <= not(layer3_outputs(4914));
    layer4_outputs(5577) <= not((layer3_outputs(4561)) xor (layer3_outputs(5588)));
    layer4_outputs(5578) <= (layer3_outputs(5397)) or (layer3_outputs(5191));
    layer4_outputs(5579) <= layer3_outputs(1500);
    layer4_outputs(5580) <= not(layer3_outputs(6861));
    layer4_outputs(5581) <= not(layer3_outputs(2190));
    layer4_outputs(5582) <= not(layer3_outputs(1441));
    layer4_outputs(5583) <= not(layer3_outputs(6450)) or (layer3_outputs(4521));
    layer4_outputs(5584) <= not(layer3_outputs(2487));
    layer4_outputs(5585) <= layer3_outputs(5270);
    layer4_outputs(5586) <= not(layer3_outputs(1775));
    layer4_outputs(5587) <= not(layer3_outputs(5055));
    layer4_outputs(5588) <= (layer3_outputs(504)) and not (layer3_outputs(1183));
    layer4_outputs(5589) <= layer3_outputs(2073);
    layer4_outputs(5590) <= (layer3_outputs(6426)) or (layer3_outputs(3971));
    layer4_outputs(5591) <= layer3_outputs(3318);
    layer4_outputs(5592) <= (layer3_outputs(6073)) and not (layer3_outputs(3589));
    layer4_outputs(5593) <= (layer3_outputs(3476)) and not (layer3_outputs(1401));
    layer4_outputs(5594) <= not(layer3_outputs(3245));
    layer4_outputs(5595) <= not(layer3_outputs(4759)) or (layer3_outputs(2198));
    layer4_outputs(5596) <= layer3_outputs(6547);
    layer4_outputs(5597) <= not(layer3_outputs(4004)) or (layer3_outputs(4757));
    layer4_outputs(5598) <= layer3_outputs(2291);
    layer4_outputs(5599) <= (layer3_outputs(6718)) xor (layer3_outputs(3));
    layer4_outputs(5600) <= not(layer3_outputs(7131)) or (layer3_outputs(2182));
    layer4_outputs(5601) <= layer3_outputs(4546);
    layer4_outputs(5602) <= not(layer3_outputs(577));
    layer4_outputs(5603) <= layer3_outputs(2906);
    layer4_outputs(5604) <= not(layer3_outputs(5682));
    layer4_outputs(5605) <= not((layer3_outputs(3255)) xor (layer3_outputs(2857)));
    layer4_outputs(5606) <= layer3_outputs(3553);
    layer4_outputs(5607) <= layer3_outputs(290);
    layer4_outputs(5608) <= layer3_outputs(1863);
    layer4_outputs(5609) <= not(layer3_outputs(5522));
    layer4_outputs(5610) <= (layer3_outputs(4888)) xor (layer3_outputs(5126));
    layer4_outputs(5611) <= not(layer3_outputs(5476));
    layer4_outputs(5612) <= (layer3_outputs(1151)) xor (layer3_outputs(7271));
    layer4_outputs(5613) <= not(layer3_outputs(2178));
    layer4_outputs(5614) <= not(layer3_outputs(2101));
    layer4_outputs(5615) <= not(layer3_outputs(3281));
    layer4_outputs(5616) <= layer3_outputs(6946);
    layer4_outputs(5617) <= '1';
    layer4_outputs(5618) <= layer3_outputs(69);
    layer4_outputs(5619) <= not((layer3_outputs(5189)) and (layer3_outputs(6493)));
    layer4_outputs(5620) <= not(layer3_outputs(7539));
    layer4_outputs(5621) <= not((layer3_outputs(3651)) or (layer3_outputs(1054)));
    layer4_outputs(5622) <= (layer3_outputs(1339)) and not (layer3_outputs(284));
    layer4_outputs(5623) <= not(layer3_outputs(2747));
    layer4_outputs(5624) <= not(layer3_outputs(5303));
    layer4_outputs(5625) <= not(layer3_outputs(7206));
    layer4_outputs(5626) <= layer3_outputs(2740);
    layer4_outputs(5627) <= layer3_outputs(1422);
    layer4_outputs(5628) <= layer3_outputs(2900);
    layer4_outputs(5629) <= layer3_outputs(1459);
    layer4_outputs(5630) <= layer3_outputs(2775);
    layer4_outputs(5631) <= not(layer3_outputs(3043));
    layer4_outputs(5632) <= not(layer3_outputs(1636));
    layer4_outputs(5633) <= layer3_outputs(133);
    layer4_outputs(5634) <= not(layer3_outputs(6007)) or (layer3_outputs(1061));
    layer4_outputs(5635) <= (layer3_outputs(1642)) xor (layer3_outputs(4920));
    layer4_outputs(5636) <= (layer3_outputs(3796)) xor (layer3_outputs(1062));
    layer4_outputs(5637) <= not(layer3_outputs(7586));
    layer4_outputs(5638) <= (layer3_outputs(5145)) xor (layer3_outputs(6637));
    layer4_outputs(5639) <= layer3_outputs(4497);
    layer4_outputs(5640) <= layer3_outputs(5546);
    layer4_outputs(5641) <= not(layer3_outputs(4945));
    layer4_outputs(5642) <= layer3_outputs(5836);
    layer4_outputs(5643) <= not((layer3_outputs(2788)) and (layer3_outputs(7176)));
    layer4_outputs(5644) <= layer3_outputs(6638);
    layer4_outputs(5645) <= not(layer3_outputs(1444)) or (layer3_outputs(1862));
    layer4_outputs(5646) <= not((layer3_outputs(5475)) xor (layer3_outputs(4357)));
    layer4_outputs(5647) <= not(layer3_outputs(3830));
    layer4_outputs(5648) <= layer3_outputs(1597);
    layer4_outputs(5649) <= not((layer3_outputs(4804)) and (layer3_outputs(5852)));
    layer4_outputs(5650) <= not((layer3_outputs(6034)) or (layer3_outputs(2898)));
    layer4_outputs(5651) <= not(layer3_outputs(7512));
    layer4_outputs(5652) <= (layer3_outputs(4605)) and not (layer3_outputs(2635));
    layer4_outputs(5653) <= not(layer3_outputs(3816)) or (layer3_outputs(2136));
    layer4_outputs(5654) <= not(layer3_outputs(3767));
    layer4_outputs(5655) <= not(layer3_outputs(4157)) or (layer3_outputs(3836));
    layer4_outputs(5656) <= (layer3_outputs(3832)) and not (layer3_outputs(352));
    layer4_outputs(5657) <= not(layer3_outputs(5036)) or (layer3_outputs(5776));
    layer4_outputs(5658) <= not((layer3_outputs(5105)) or (layer3_outputs(4818)));
    layer4_outputs(5659) <= not(layer3_outputs(1404)) or (layer3_outputs(3333));
    layer4_outputs(5660) <= layer3_outputs(3781);
    layer4_outputs(5661) <= not(layer3_outputs(2992)) or (layer3_outputs(6569));
    layer4_outputs(5662) <= (layer3_outputs(4901)) xor (layer3_outputs(3099));
    layer4_outputs(5663) <= (layer3_outputs(4612)) xor (layer3_outputs(1254));
    layer4_outputs(5664) <= (layer3_outputs(3571)) and not (layer3_outputs(5714));
    layer4_outputs(5665) <= layer3_outputs(1827);
    layer4_outputs(5666) <= (layer3_outputs(2941)) xor (layer3_outputs(1770));
    layer4_outputs(5667) <= not(layer3_outputs(6196));
    layer4_outputs(5668) <= not((layer3_outputs(5246)) or (layer3_outputs(464)));
    layer4_outputs(5669) <= '0';
    layer4_outputs(5670) <= not(layer3_outputs(3688));
    layer4_outputs(5671) <= layer3_outputs(5111);
    layer4_outputs(5672) <= (layer3_outputs(5097)) xor (layer3_outputs(2972));
    layer4_outputs(5673) <= not(layer3_outputs(4275)) or (layer3_outputs(6917));
    layer4_outputs(5674) <= (layer3_outputs(1181)) and (layer3_outputs(4449));
    layer4_outputs(5675) <= (layer3_outputs(6715)) and not (layer3_outputs(3156));
    layer4_outputs(5676) <= layer3_outputs(7436);
    layer4_outputs(5677) <= not(layer3_outputs(5410));
    layer4_outputs(5678) <= layer3_outputs(3120);
    layer4_outputs(5679) <= not((layer3_outputs(3498)) and (layer3_outputs(3623)));
    layer4_outputs(5680) <= not(layer3_outputs(1141));
    layer4_outputs(5681) <= layer3_outputs(3893);
    layer4_outputs(5682) <= (layer3_outputs(2910)) xor (layer3_outputs(5389));
    layer4_outputs(5683) <= '1';
    layer4_outputs(5684) <= layer3_outputs(7394);
    layer4_outputs(5685) <= not(layer3_outputs(5458));
    layer4_outputs(5686) <= layer3_outputs(4917);
    layer4_outputs(5687) <= layer3_outputs(4405);
    layer4_outputs(5688) <= not(layer3_outputs(3105));
    layer4_outputs(5689) <= (layer3_outputs(3051)) and not (layer3_outputs(3690));
    layer4_outputs(5690) <= not(layer3_outputs(1124));
    layer4_outputs(5691) <= not(layer3_outputs(7604));
    layer4_outputs(5692) <= not(layer3_outputs(415));
    layer4_outputs(5693) <= layer3_outputs(6861);
    layer4_outputs(5694) <= not(layer3_outputs(6725));
    layer4_outputs(5695) <= (layer3_outputs(3232)) or (layer3_outputs(2837));
    layer4_outputs(5696) <= not(layer3_outputs(2891));
    layer4_outputs(5697) <= not(layer3_outputs(7027));
    layer4_outputs(5698) <= not(layer3_outputs(824)) or (layer3_outputs(1333));
    layer4_outputs(5699) <= not(layer3_outputs(4659));
    layer4_outputs(5700) <= not(layer3_outputs(2398));
    layer4_outputs(5701) <= not(layer3_outputs(4499)) or (layer3_outputs(1208));
    layer4_outputs(5702) <= not((layer3_outputs(3337)) or (layer3_outputs(4482)));
    layer4_outputs(5703) <= not(layer3_outputs(6997));
    layer4_outputs(5704) <= layer3_outputs(7479);
    layer4_outputs(5705) <= layer3_outputs(5715);
    layer4_outputs(5706) <= (layer3_outputs(2802)) and (layer3_outputs(2264));
    layer4_outputs(5707) <= (layer3_outputs(6511)) and not (layer3_outputs(5287));
    layer4_outputs(5708) <= (layer3_outputs(1773)) and (layer3_outputs(1045));
    layer4_outputs(5709) <= not((layer3_outputs(5680)) xor (layer3_outputs(3693)));
    layer4_outputs(5710) <= (layer3_outputs(3874)) or (layer3_outputs(4071));
    layer4_outputs(5711) <= not(layer3_outputs(2684));
    layer4_outputs(5712) <= layer3_outputs(2928);
    layer4_outputs(5713) <= not(layer3_outputs(5028));
    layer4_outputs(5714) <= (layer3_outputs(6747)) or (layer3_outputs(1050));
    layer4_outputs(5715) <= (layer3_outputs(5018)) and (layer3_outputs(7342));
    layer4_outputs(5716) <= not(layer3_outputs(4266));
    layer4_outputs(5717) <= layer3_outputs(7644);
    layer4_outputs(5718) <= not((layer3_outputs(6533)) xor (layer3_outputs(3925)));
    layer4_outputs(5719) <= (layer3_outputs(3970)) and (layer3_outputs(1871));
    layer4_outputs(5720) <= not(layer3_outputs(1117));
    layer4_outputs(5721) <= not(layer3_outputs(1705));
    layer4_outputs(5722) <= not((layer3_outputs(6346)) xor (layer3_outputs(7049)));
    layer4_outputs(5723) <= not(layer3_outputs(3841));
    layer4_outputs(5724) <= (layer3_outputs(5928)) and not (layer3_outputs(3031));
    layer4_outputs(5725) <= not(layer3_outputs(1));
    layer4_outputs(5726) <= not(layer3_outputs(3452));
    layer4_outputs(5727) <= (layer3_outputs(976)) and not (layer3_outputs(6220));
    layer4_outputs(5728) <= layer3_outputs(4711);
    layer4_outputs(5729) <= '0';
    layer4_outputs(5730) <= not(layer3_outputs(5847));
    layer4_outputs(5731) <= (layer3_outputs(4981)) and not (layer3_outputs(1791));
    layer4_outputs(5732) <= not((layer3_outputs(6603)) xor (layer3_outputs(2030)));
    layer4_outputs(5733) <= layer3_outputs(4799);
    layer4_outputs(5734) <= layer3_outputs(3829);
    layer4_outputs(5735) <= not(layer3_outputs(4495));
    layer4_outputs(5736) <= layer3_outputs(2966);
    layer4_outputs(5737) <= not(layer3_outputs(4664));
    layer4_outputs(5738) <= not(layer3_outputs(3528));
    layer4_outputs(5739) <= (layer3_outputs(2972)) and (layer3_outputs(1652));
    layer4_outputs(5740) <= (layer3_outputs(6886)) and not (layer3_outputs(3311));
    layer4_outputs(5741) <= not((layer3_outputs(2917)) or (layer3_outputs(6727)));
    layer4_outputs(5742) <= not(layer3_outputs(6634));
    layer4_outputs(5743) <= not(layer3_outputs(1635));
    layer4_outputs(5744) <= not(layer3_outputs(5230));
    layer4_outputs(5745) <= not(layer3_outputs(2654));
    layer4_outputs(5746) <= not(layer3_outputs(6293)) or (layer3_outputs(1483));
    layer4_outputs(5747) <= (layer3_outputs(5075)) xor (layer3_outputs(1574));
    layer4_outputs(5748) <= layer3_outputs(2419);
    layer4_outputs(5749) <= (layer3_outputs(825)) and not (layer3_outputs(1319));
    layer4_outputs(5750) <= not(layer3_outputs(3175));
    layer4_outputs(5751) <= (layer3_outputs(608)) xor (layer3_outputs(2899));
    layer4_outputs(5752) <= not(layer3_outputs(134));
    layer4_outputs(5753) <= not(layer3_outputs(2801));
    layer4_outputs(5754) <= layer3_outputs(7638);
    layer4_outputs(5755) <= layer3_outputs(1204);
    layer4_outputs(5756) <= not(layer3_outputs(4056));
    layer4_outputs(5757) <= (layer3_outputs(1442)) xor (layer3_outputs(1660));
    layer4_outputs(5758) <= (layer3_outputs(80)) and not (layer3_outputs(4592));
    layer4_outputs(5759) <= not(layer3_outputs(2312));
    layer4_outputs(5760) <= not(layer3_outputs(6723));
    layer4_outputs(5761) <= not((layer3_outputs(7117)) or (layer3_outputs(3745)));
    layer4_outputs(5762) <= not((layer3_outputs(4462)) or (layer3_outputs(7112)));
    layer4_outputs(5763) <= not(layer3_outputs(4006));
    layer4_outputs(5764) <= not(layer3_outputs(466)) or (layer3_outputs(6268));
    layer4_outputs(5765) <= (layer3_outputs(1369)) and not (layer3_outputs(4153));
    layer4_outputs(5766) <= (layer3_outputs(975)) and not (layer3_outputs(5975));
    layer4_outputs(5767) <= layer3_outputs(6227);
    layer4_outputs(5768) <= layer3_outputs(6232);
    layer4_outputs(5769) <= not((layer3_outputs(4489)) and (layer3_outputs(6302)));
    layer4_outputs(5770) <= layer3_outputs(4107);
    layer4_outputs(5771) <= layer3_outputs(4514);
    layer4_outputs(5772) <= (layer3_outputs(3779)) and (layer3_outputs(7492));
    layer4_outputs(5773) <= not(layer3_outputs(4930));
    layer4_outputs(5774) <= layer3_outputs(5909);
    layer4_outputs(5775) <= layer3_outputs(4727);
    layer4_outputs(5776) <= layer3_outputs(1625);
    layer4_outputs(5777) <= not(layer3_outputs(2486));
    layer4_outputs(5778) <= layer3_outputs(4529);
    layer4_outputs(5779) <= not(layer3_outputs(1620));
    layer4_outputs(5780) <= (layer3_outputs(1843)) and (layer3_outputs(6910));
    layer4_outputs(5781) <= not((layer3_outputs(7243)) or (layer3_outputs(5663)));
    layer4_outputs(5782) <= not((layer3_outputs(5386)) xor (layer3_outputs(7006)));
    layer4_outputs(5783) <= (layer3_outputs(7497)) and not (layer3_outputs(7196));
    layer4_outputs(5784) <= not(layer3_outputs(66));
    layer4_outputs(5785) <= not(layer3_outputs(823));
    layer4_outputs(5786) <= layer3_outputs(1123);
    layer4_outputs(5787) <= not(layer3_outputs(38));
    layer4_outputs(5788) <= (layer3_outputs(4891)) and not (layer3_outputs(187));
    layer4_outputs(5789) <= not((layer3_outputs(1590)) xor (layer3_outputs(2372)));
    layer4_outputs(5790) <= not(layer3_outputs(4089));
    layer4_outputs(5791) <= layer3_outputs(5702);
    layer4_outputs(5792) <= layer3_outputs(461);
    layer4_outputs(5793) <= not(layer3_outputs(2239));
    layer4_outputs(5794) <= not(layer3_outputs(1943));
    layer4_outputs(5795) <= not((layer3_outputs(3034)) xor (layer3_outputs(5032)));
    layer4_outputs(5796) <= layer3_outputs(5331);
    layer4_outputs(5797) <= (layer3_outputs(5449)) xor (layer3_outputs(3642));
    layer4_outputs(5798) <= not(layer3_outputs(6934));
    layer4_outputs(5799) <= not((layer3_outputs(5510)) xor (layer3_outputs(6006)));
    layer4_outputs(5800) <= layer3_outputs(321);
    layer4_outputs(5801) <= not((layer3_outputs(2713)) xor (layer3_outputs(1547)));
    layer4_outputs(5802) <= not(layer3_outputs(5881));
    layer4_outputs(5803) <= not(layer3_outputs(7607));
    layer4_outputs(5804) <= (layer3_outputs(1397)) and not (layer3_outputs(1387));
    layer4_outputs(5805) <= not(layer3_outputs(134));
    layer4_outputs(5806) <= not(layer3_outputs(4414));
    layer4_outputs(5807) <= (layer3_outputs(3247)) and not (layer3_outputs(6799));
    layer4_outputs(5808) <= not(layer3_outputs(4440));
    layer4_outputs(5809) <= not((layer3_outputs(6533)) or (layer3_outputs(4306)));
    layer4_outputs(5810) <= layer3_outputs(2681);
    layer4_outputs(5811) <= layer3_outputs(649);
    layer4_outputs(5812) <= not(layer3_outputs(7033));
    layer4_outputs(5813) <= not(layer3_outputs(1360));
    layer4_outputs(5814) <= '1';
    layer4_outputs(5815) <= (layer3_outputs(4231)) or (layer3_outputs(3877));
    layer4_outputs(5816) <= not(layer3_outputs(5932)) or (layer3_outputs(816));
    layer4_outputs(5817) <= (layer3_outputs(2378)) and not (layer3_outputs(1199));
    layer4_outputs(5818) <= (layer3_outputs(3578)) and not (layer3_outputs(2845));
    layer4_outputs(5819) <= layer3_outputs(1061);
    layer4_outputs(5820) <= (layer3_outputs(1396)) or (layer3_outputs(1899));
    layer4_outputs(5821) <= not(layer3_outputs(767));
    layer4_outputs(5822) <= layer3_outputs(6603);
    layer4_outputs(5823) <= layer3_outputs(309);
    layer4_outputs(5824) <= (layer3_outputs(2781)) and not (layer3_outputs(3206));
    layer4_outputs(5825) <= layer3_outputs(2793);
    layer4_outputs(5826) <= not(layer3_outputs(1060)) or (layer3_outputs(3294));
    layer4_outputs(5827) <= (layer3_outputs(1246)) and not (layer3_outputs(7241));
    layer4_outputs(5828) <= not(layer3_outputs(2313));
    layer4_outputs(5829) <= layer3_outputs(7150);
    layer4_outputs(5830) <= not(layer3_outputs(6150));
    layer4_outputs(5831) <= not(layer3_outputs(4847));
    layer4_outputs(5832) <= not(layer3_outputs(5268)) or (layer3_outputs(6086));
    layer4_outputs(5833) <= not((layer3_outputs(865)) and (layer3_outputs(6341)));
    layer4_outputs(5834) <= layer3_outputs(315);
    layer4_outputs(5835) <= not(layer3_outputs(477)) or (layer3_outputs(523));
    layer4_outputs(5836) <= not(layer3_outputs(6141));
    layer4_outputs(5837) <= not(layer3_outputs(6322));
    layer4_outputs(5838) <= not(layer3_outputs(3937));
    layer4_outputs(5839) <= not((layer3_outputs(4774)) or (layer3_outputs(3090)));
    layer4_outputs(5840) <= (layer3_outputs(3622)) xor (layer3_outputs(3055));
    layer4_outputs(5841) <= (layer3_outputs(2216)) and (layer3_outputs(4822));
    layer4_outputs(5842) <= (layer3_outputs(1748)) and (layer3_outputs(6604));
    layer4_outputs(5843) <= (layer3_outputs(5882)) or (layer3_outputs(3689));
    layer4_outputs(5844) <= layer3_outputs(138);
    layer4_outputs(5845) <= not(layer3_outputs(6494));
    layer4_outputs(5846) <= (layer3_outputs(6180)) and (layer3_outputs(6962));
    layer4_outputs(5847) <= layer3_outputs(6001);
    layer4_outputs(5848) <= layer3_outputs(5308);
    layer4_outputs(5849) <= not(layer3_outputs(3226));
    layer4_outputs(5850) <= layer3_outputs(7073);
    layer4_outputs(5851) <= (layer3_outputs(6198)) or (layer3_outputs(3018));
    layer4_outputs(5852) <= layer3_outputs(7095);
    layer4_outputs(5853) <= layer3_outputs(951);
    layer4_outputs(5854) <= layer3_outputs(1552);
    layer4_outputs(5855) <= layer3_outputs(1851);
    layer4_outputs(5856) <= layer3_outputs(4810);
    layer4_outputs(5857) <= layer3_outputs(435);
    layer4_outputs(5858) <= not((layer3_outputs(715)) and (layer3_outputs(1680)));
    layer4_outputs(5859) <= layer3_outputs(5096);
    layer4_outputs(5860) <= not(layer3_outputs(3140));
    layer4_outputs(5861) <= (layer3_outputs(5331)) and not (layer3_outputs(7270));
    layer4_outputs(5862) <= layer3_outputs(1605);
    layer4_outputs(5863) <= not(layer3_outputs(7554));
    layer4_outputs(5864) <= (layer3_outputs(4538)) xor (layer3_outputs(905));
    layer4_outputs(5865) <= not(layer3_outputs(5967));
    layer4_outputs(5866) <= not(layer3_outputs(3175));
    layer4_outputs(5867) <= not(layer3_outputs(5533));
    layer4_outputs(5868) <= (layer3_outputs(3306)) and not (layer3_outputs(216));
    layer4_outputs(5869) <= not((layer3_outputs(1527)) or (layer3_outputs(6980)));
    layer4_outputs(5870) <= layer3_outputs(455);
    layer4_outputs(5871) <= (layer3_outputs(5821)) and (layer3_outputs(916));
    layer4_outputs(5872) <= (layer3_outputs(1102)) and not (layer3_outputs(6283));
    layer4_outputs(5873) <= not(layer3_outputs(2271));
    layer4_outputs(5874) <= layer3_outputs(4352);
    layer4_outputs(5875) <= (layer3_outputs(1673)) xor (layer3_outputs(3743));
    layer4_outputs(5876) <= not(layer3_outputs(6787));
    layer4_outputs(5877) <= layer3_outputs(837);
    layer4_outputs(5878) <= not(layer3_outputs(839));
    layer4_outputs(5879) <= not(layer3_outputs(2427));
    layer4_outputs(5880) <= (layer3_outputs(2728)) and (layer3_outputs(5368));
    layer4_outputs(5881) <= (layer3_outputs(4807)) xor (layer3_outputs(3641));
    layer4_outputs(5882) <= not(layer3_outputs(3738)) or (layer3_outputs(1096));
    layer4_outputs(5883) <= not(layer3_outputs(2437));
    layer4_outputs(5884) <= not((layer3_outputs(7346)) xor (layer3_outputs(7531)));
    layer4_outputs(5885) <= not((layer3_outputs(6651)) xor (layer3_outputs(1476)));
    layer4_outputs(5886) <= (layer3_outputs(4560)) and not (layer3_outputs(5784));
    layer4_outputs(5887) <= not(layer3_outputs(1817));
    layer4_outputs(5888) <= not((layer3_outputs(6889)) and (layer3_outputs(2162)));
    layer4_outputs(5889) <= not(layer3_outputs(2805));
    layer4_outputs(5890) <= not(layer3_outputs(3257));
    layer4_outputs(5891) <= layer3_outputs(869);
    layer4_outputs(5892) <= (layer3_outputs(3072)) or (layer3_outputs(6817));
    layer4_outputs(5893) <= not((layer3_outputs(6673)) xor (layer3_outputs(4059)));
    layer4_outputs(5894) <= not(layer3_outputs(4625));
    layer4_outputs(5895) <= not(layer3_outputs(415)) or (layer3_outputs(4040));
    layer4_outputs(5896) <= (layer3_outputs(2485)) xor (layer3_outputs(7395));
    layer4_outputs(5897) <= '1';
    layer4_outputs(5898) <= not(layer3_outputs(5931));
    layer4_outputs(5899) <= not(layer3_outputs(825));
    layer4_outputs(5900) <= not((layer3_outputs(3740)) xor (layer3_outputs(4777)));
    layer4_outputs(5901) <= layer3_outputs(6812);
    layer4_outputs(5902) <= (layer3_outputs(6873)) and (layer3_outputs(4077));
    layer4_outputs(5903) <= (layer3_outputs(4477)) and not (layer3_outputs(551));
    layer4_outputs(5904) <= (layer3_outputs(5849)) and (layer3_outputs(4762));
    layer4_outputs(5905) <= layer3_outputs(1465);
    layer4_outputs(5906) <= not(layer3_outputs(1106));
    layer4_outputs(5907) <= not(layer3_outputs(6571)) or (layer3_outputs(3310));
    layer4_outputs(5908) <= '1';
    layer4_outputs(5909) <= not(layer3_outputs(4531));
    layer4_outputs(5910) <= (layer3_outputs(6454)) and not (layer3_outputs(3331));
    layer4_outputs(5911) <= not((layer3_outputs(5977)) xor (layer3_outputs(2953)));
    layer4_outputs(5912) <= layer3_outputs(6654);
    layer4_outputs(5913) <= not(layer3_outputs(6271)) or (layer3_outputs(1481));
    layer4_outputs(5914) <= not(layer3_outputs(2708)) or (layer3_outputs(6706));
    layer4_outputs(5915) <= layer3_outputs(2939);
    layer4_outputs(5916) <= layer3_outputs(2201);
    layer4_outputs(5917) <= not(layer3_outputs(1359)) or (layer3_outputs(7469));
    layer4_outputs(5918) <= layer3_outputs(1129);
    layer4_outputs(5919) <= not((layer3_outputs(2480)) and (layer3_outputs(2144)));
    layer4_outputs(5920) <= (layer3_outputs(6496)) and not (layer3_outputs(6858));
    layer4_outputs(5921) <= (layer3_outputs(1795)) and not (layer3_outputs(6907));
    layer4_outputs(5922) <= not(layer3_outputs(5784));
    layer4_outputs(5923) <= not(layer3_outputs(7338));
    layer4_outputs(5924) <= not(layer3_outputs(872)) or (layer3_outputs(2078));
    layer4_outputs(5925) <= (layer3_outputs(6989)) or (layer3_outputs(4673));
    layer4_outputs(5926) <= not(layer3_outputs(3322));
    layer4_outputs(5927) <= not(layer3_outputs(1024)) or (layer3_outputs(4492));
    layer4_outputs(5928) <= (layer3_outputs(2)) xor (layer3_outputs(4011));
    layer4_outputs(5929) <= (layer3_outputs(3954)) or (layer3_outputs(1256));
    layer4_outputs(5930) <= not(layer3_outputs(2504));
    layer4_outputs(5931) <= layer3_outputs(3968);
    layer4_outputs(5932) <= layer3_outputs(4075);
    layer4_outputs(5933) <= not(layer3_outputs(3467));
    layer4_outputs(5934) <= not(layer3_outputs(6270));
    layer4_outputs(5935) <= not((layer3_outputs(5144)) xor (layer3_outputs(7051)));
    layer4_outputs(5936) <= not(layer3_outputs(5159));
    layer4_outputs(5937) <= (layer3_outputs(5841)) or (layer3_outputs(3436));
    layer4_outputs(5938) <= layer3_outputs(7000);
    layer4_outputs(5939) <= not((layer3_outputs(7161)) and (layer3_outputs(4281)));
    layer4_outputs(5940) <= (layer3_outputs(4166)) xor (layer3_outputs(4851));
    layer4_outputs(5941) <= not(layer3_outputs(3458)) or (layer3_outputs(6008));
    layer4_outputs(5942) <= (layer3_outputs(6359)) and not (layer3_outputs(5590));
    layer4_outputs(5943) <= layer3_outputs(1216);
    layer4_outputs(5944) <= (layer3_outputs(7094)) and not (layer3_outputs(1687));
    layer4_outputs(5945) <= not((layer3_outputs(4828)) or (layer3_outputs(1048)));
    layer4_outputs(5946) <= not(layer3_outputs(5772));
    layer4_outputs(5947) <= not(layer3_outputs(2760));
    layer4_outputs(5948) <= layer3_outputs(6613);
    layer4_outputs(5949) <= (layer3_outputs(2444)) or (layer3_outputs(5726));
    layer4_outputs(5950) <= layer3_outputs(4370);
    layer4_outputs(5951) <= layer3_outputs(3595);
    layer4_outputs(5952) <= layer3_outputs(5518);
    layer4_outputs(5953) <= (layer3_outputs(7579)) and not (layer3_outputs(7028));
    layer4_outputs(5954) <= not(layer3_outputs(6909));
    layer4_outputs(5955) <= not(layer3_outputs(5024));
    layer4_outputs(5956) <= (layer3_outputs(4718)) xor (layer3_outputs(1544));
    layer4_outputs(5957) <= not((layer3_outputs(1794)) xor (layer3_outputs(878)));
    layer4_outputs(5958) <= '1';
    layer4_outputs(5959) <= not(layer3_outputs(634));
    layer4_outputs(5960) <= (layer3_outputs(4730)) and (layer3_outputs(2154));
    layer4_outputs(5961) <= (layer3_outputs(7408)) and (layer3_outputs(5314));
    layer4_outputs(5962) <= layer3_outputs(1225);
    layer4_outputs(5963) <= layer3_outputs(1407);
    layer4_outputs(5964) <= not(layer3_outputs(164));
    layer4_outputs(5965) <= not(layer3_outputs(4463)) or (layer3_outputs(1684));
    layer4_outputs(5966) <= (layer3_outputs(3356)) and not (layer3_outputs(3763));
    layer4_outputs(5967) <= not(layer3_outputs(6768)) or (layer3_outputs(863));
    layer4_outputs(5968) <= (layer3_outputs(3410)) xor (layer3_outputs(6775));
    layer4_outputs(5969) <= layer3_outputs(5451);
    layer4_outputs(5970) <= not(layer3_outputs(5679)) or (layer3_outputs(1879));
    layer4_outputs(5971) <= layer3_outputs(1837);
    layer4_outputs(5972) <= (layer3_outputs(1379)) xor (layer3_outputs(7663));
    layer4_outputs(5973) <= (layer3_outputs(6862)) and not (layer3_outputs(5271));
    layer4_outputs(5974) <= (layer3_outputs(2956)) and not (layer3_outputs(4020));
    layer4_outputs(5975) <= not((layer3_outputs(4285)) or (layer3_outputs(3513)));
    layer4_outputs(5976) <= layer3_outputs(4512);
    layer4_outputs(5977) <= not((layer3_outputs(3176)) or (layer3_outputs(1260)));
    layer4_outputs(5978) <= (layer3_outputs(2568)) or (layer3_outputs(1731));
    layer4_outputs(5979) <= not(layer3_outputs(1220));
    layer4_outputs(5980) <= (layer3_outputs(1202)) or (layer3_outputs(2844));
    layer4_outputs(5981) <= layer3_outputs(6037);
    layer4_outputs(5982) <= (layer3_outputs(493)) and not (layer3_outputs(3859));
    layer4_outputs(5983) <= layer3_outputs(848);
    layer4_outputs(5984) <= not(layer3_outputs(24)) or (layer3_outputs(3730));
    layer4_outputs(5985) <= not(layer3_outputs(3257)) or (layer3_outputs(2843));
    layer4_outputs(5986) <= (layer3_outputs(6242)) xor (layer3_outputs(4301));
    layer4_outputs(5987) <= not(layer3_outputs(3181)) or (layer3_outputs(4879));
    layer4_outputs(5988) <= not((layer3_outputs(1717)) and (layer3_outputs(4814)));
    layer4_outputs(5989) <= '0';
    layer4_outputs(5990) <= layer3_outputs(322);
    layer4_outputs(5991) <= (layer3_outputs(1401)) and (layer3_outputs(1553));
    layer4_outputs(5992) <= not(layer3_outputs(4318));
    layer4_outputs(5993) <= not(layer3_outputs(7040));
    layer4_outputs(5994) <= (layer3_outputs(98)) xor (layer3_outputs(2320));
    layer4_outputs(5995) <= not(layer3_outputs(7530));
    layer4_outputs(5996) <= (layer3_outputs(6225)) or (layer3_outputs(7278));
    layer4_outputs(5997) <= layer3_outputs(1934);
    layer4_outputs(5998) <= layer3_outputs(5499);
    layer4_outputs(5999) <= layer3_outputs(3432);
    layer4_outputs(6000) <= layer3_outputs(1168);
    layer4_outputs(6001) <= not(layer3_outputs(6783));
    layer4_outputs(6002) <= layer3_outputs(6645);
    layer4_outputs(6003) <= not(layer3_outputs(4297));
    layer4_outputs(6004) <= '1';
    layer4_outputs(6005) <= (layer3_outputs(6614)) and not (layer3_outputs(3837));
    layer4_outputs(6006) <= layer3_outputs(6072);
    layer4_outputs(6007) <= (layer3_outputs(1138)) xor (layer3_outputs(1625));
    layer4_outputs(6008) <= (layer3_outputs(3536)) and not (layer3_outputs(753));
    layer4_outputs(6009) <= not(layer3_outputs(2102));
    layer4_outputs(6010) <= layer3_outputs(6926);
    layer4_outputs(6011) <= layer3_outputs(2604);
    layer4_outputs(6012) <= (layer3_outputs(4883)) and not (layer3_outputs(678));
    layer4_outputs(6013) <= not(layer3_outputs(2103));
    layer4_outputs(6014) <= not(layer3_outputs(6826));
    layer4_outputs(6015) <= layer3_outputs(6868);
    layer4_outputs(6016) <= not((layer3_outputs(752)) xor (layer3_outputs(6130)));
    layer4_outputs(6017) <= not((layer3_outputs(1677)) xor (layer3_outputs(240)));
    layer4_outputs(6018) <= (layer3_outputs(6620)) and not (layer3_outputs(3789));
    layer4_outputs(6019) <= (layer3_outputs(1063)) or (layer3_outputs(418));
    layer4_outputs(6020) <= not(layer3_outputs(1305));
    layer4_outputs(6021) <= layer3_outputs(3334);
    layer4_outputs(6022) <= (layer3_outputs(2508)) and not (layer3_outputs(6993));
    layer4_outputs(6023) <= layer3_outputs(1251);
    layer4_outputs(6024) <= (layer3_outputs(4069)) and not (layer3_outputs(6393));
    layer4_outputs(6025) <= not((layer3_outputs(3261)) and (layer3_outputs(4771)));
    layer4_outputs(6026) <= (layer3_outputs(6349)) and not (layer3_outputs(1665));
    layer4_outputs(6027) <= (layer3_outputs(1410)) and not (layer3_outputs(4677));
    layer4_outputs(6028) <= not(layer3_outputs(6700));
    layer4_outputs(6029) <= not(layer3_outputs(4071)) or (layer3_outputs(4046));
    layer4_outputs(6030) <= not((layer3_outputs(4834)) and (layer3_outputs(6519)));
    layer4_outputs(6031) <= not((layer3_outputs(5927)) or (layer3_outputs(2596)));
    layer4_outputs(6032) <= layer3_outputs(877);
    layer4_outputs(6033) <= layer3_outputs(4278);
    layer4_outputs(6034) <= (layer3_outputs(2235)) and not (layer3_outputs(6643));
    layer4_outputs(6035) <= not(layer3_outputs(5937));
    layer4_outputs(6036) <= not(layer3_outputs(5411));
    layer4_outputs(6037) <= layer3_outputs(5005);
    layer4_outputs(6038) <= not(layer3_outputs(7186));
    layer4_outputs(6039) <= (layer3_outputs(2499)) or (layer3_outputs(755));
    layer4_outputs(6040) <= layer3_outputs(6549);
    layer4_outputs(6041) <= not(layer3_outputs(1576)) or (layer3_outputs(5813));
    layer4_outputs(6042) <= layer3_outputs(7295);
    layer4_outputs(6043) <= not(layer3_outputs(2630));
    layer4_outputs(6044) <= not(layer3_outputs(6437));
    layer4_outputs(6045) <= not((layer3_outputs(5438)) or (layer3_outputs(5066)));
    layer4_outputs(6046) <= not(layer3_outputs(4903));
    layer4_outputs(6047) <= not(layer3_outputs(4601));
    layer4_outputs(6048) <= layer3_outputs(3464);
    layer4_outputs(6049) <= (layer3_outputs(7141)) and (layer3_outputs(3446));
    layer4_outputs(6050) <= not(layer3_outputs(2367));
    layer4_outputs(6051) <= not((layer3_outputs(5737)) and (layer3_outputs(4062)));
    layer4_outputs(6052) <= not(layer3_outputs(3996)) or (layer3_outputs(1358));
    layer4_outputs(6053) <= not(layer3_outputs(915));
    layer4_outputs(6054) <= '0';
    layer4_outputs(6055) <= not(layer3_outputs(3014));
    layer4_outputs(6056) <= not(layer3_outputs(5549)) or (layer3_outputs(5354));
    layer4_outputs(6057) <= layer3_outputs(6953);
    layer4_outputs(6058) <= (layer3_outputs(3548)) and not (layer3_outputs(1159));
    layer4_outputs(6059) <= not(layer3_outputs(6162));
    layer4_outputs(6060) <= layer3_outputs(4883);
    layer4_outputs(6061) <= not(layer3_outputs(635));
    layer4_outputs(6062) <= (layer3_outputs(1948)) and not (layer3_outputs(7594));
    layer4_outputs(6063) <= (layer3_outputs(268)) xor (layer3_outputs(7355));
    layer4_outputs(6064) <= layer3_outputs(5996);
    layer4_outputs(6065) <= (layer3_outputs(2227)) and not (layer3_outputs(5264));
    layer4_outputs(6066) <= (layer3_outputs(7451)) and not (layer3_outputs(565));
    layer4_outputs(6067) <= not(layer3_outputs(123)) or (layer3_outputs(1273));
    layer4_outputs(6068) <= layer3_outputs(4262);
    layer4_outputs(6069) <= layer3_outputs(1662);
    layer4_outputs(6070) <= not((layer3_outputs(4806)) or (layer3_outputs(5531)));
    layer4_outputs(6071) <= (layer3_outputs(1694)) and (layer3_outputs(2816));
    layer4_outputs(6072) <= layer3_outputs(7180);
    layer4_outputs(6073) <= not(layer3_outputs(5855));
    layer4_outputs(6074) <= (layer3_outputs(4313)) and not (layer3_outputs(5454));
    layer4_outputs(6075) <= layer3_outputs(4965);
    layer4_outputs(6076) <= (layer3_outputs(3634)) or (layer3_outputs(2823));
    layer4_outputs(6077) <= layer3_outputs(503);
    layer4_outputs(6078) <= not(layer3_outputs(224)) or (layer3_outputs(6258));
    layer4_outputs(6079) <= not(layer3_outputs(6587)) or (layer3_outputs(2633));
    layer4_outputs(6080) <= '1';
    layer4_outputs(6081) <= (layer3_outputs(3989)) or (layer3_outputs(1576));
    layer4_outputs(6082) <= (layer3_outputs(5999)) or (layer3_outputs(889));
    layer4_outputs(6083) <= not(layer3_outputs(6912));
    layer4_outputs(6084) <= layer3_outputs(2478);
    layer4_outputs(6085) <= not((layer3_outputs(7465)) xor (layer3_outputs(6117)));
    layer4_outputs(6086) <= (layer3_outputs(2554)) and not (layer3_outputs(5404));
    layer4_outputs(6087) <= layer3_outputs(1531);
    layer4_outputs(6088) <= layer3_outputs(2289);
    layer4_outputs(6089) <= (layer3_outputs(5492)) and not (layer3_outputs(2474));
    layer4_outputs(6090) <= (layer3_outputs(3277)) and not (layer3_outputs(30));
    layer4_outputs(6091) <= layer3_outputs(2276);
    layer4_outputs(6092) <= not((layer3_outputs(2465)) and (layer3_outputs(924)));
    layer4_outputs(6093) <= layer3_outputs(1171);
    layer4_outputs(6094) <= layer3_outputs(3816);
    layer4_outputs(6095) <= layer3_outputs(1651);
    layer4_outputs(6096) <= not((layer3_outputs(1946)) and (layer3_outputs(5772)));
    layer4_outputs(6097) <= layer3_outputs(2897);
    layer4_outputs(6098) <= not((layer3_outputs(7352)) or (layer3_outputs(891)));
    layer4_outputs(6099) <= (layer3_outputs(5658)) and (layer3_outputs(7020));
    layer4_outputs(6100) <= not(layer3_outputs(3987));
    layer4_outputs(6101) <= not(layer3_outputs(6609));
    layer4_outputs(6102) <= (layer3_outputs(3985)) or (layer3_outputs(7352));
    layer4_outputs(6103) <= not(layer3_outputs(1701));
    layer4_outputs(6104) <= (layer3_outputs(1769)) and not (layer3_outputs(1855));
    layer4_outputs(6105) <= '1';
    layer4_outputs(6106) <= not(layer3_outputs(7039));
    layer4_outputs(6107) <= layer3_outputs(3592);
    layer4_outputs(6108) <= not(layer3_outputs(256));
    layer4_outputs(6109) <= (layer3_outputs(1152)) and not (layer3_outputs(3151));
    layer4_outputs(6110) <= (layer3_outputs(2693)) and (layer3_outputs(3879));
    layer4_outputs(6111) <= not(layer3_outputs(228)) or (layer3_outputs(5222));
    layer4_outputs(6112) <= not(layer3_outputs(5891)) or (layer3_outputs(5434));
    layer4_outputs(6113) <= layer3_outputs(1560);
    layer4_outputs(6114) <= not((layer3_outputs(3238)) xor (layer3_outputs(5166)));
    layer4_outputs(6115) <= (layer3_outputs(2488)) xor (layer3_outputs(2614));
    layer4_outputs(6116) <= (layer3_outputs(776)) and not (layer3_outputs(292));
    layer4_outputs(6117) <= layer3_outputs(5567);
    layer4_outputs(6118) <= not(layer3_outputs(3565));
    layer4_outputs(6119) <= (layer3_outputs(4232)) or (layer3_outputs(2032));
    layer4_outputs(6120) <= not((layer3_outputs(4599)) and (layer3_outputs(4348)));
    layer4_outputs(6121) <= not((layer3_outputs(2731)) and (layer3_outputs(5966)));
    layer4_outputs(6122) <= not(layer3_outputs(3867));
    layer4_outputs(6123) <= not(layer3_outputs(4532));
    layer4_outputs(6124) <= (layer3_outputs(6997)) and not (layer3_outputs(5559));
    layer4_outputs(6125) <= layer3_outputs(5288);
    layer4_outputs(6126) <= not((layer3_outputs(3984)) xor (layer3_outputs(5194)));
    layer4_outputs(6127) <= layer3_outputs(5086);
    layer4_outputs(6128) <= not(layer3_outputs(1566));
    layer4_outputs(6129) <= layer3_outputs(3599);
    layer4_outputs(6130) <= layer3_outputs(2134);
    layer4_outputs(6131) <= not((layer3_outputs(3507)) xor (layer3_outputs(5478)));
    layer4_outputs(6132) <= '0';
    layer4_outputs(6133) <= layer3_outputs(491);
    layer4_outputs(6134) <= not(layer3_outputs(2350));
    layer4_outputs(6135) <= layer3_outputs(6784);
    layer4_outputs(6136) <= not(layer3_outputs(280)) or (layer3_outputs(3616));
    layer4_outputs(6137) <= not(layer3_outputs(3904));
    layer4_outputs(6138) <= (layer3_outputs(3602)) and (layer3_outputs(1970));
    layer4_outputs(6139) <= (layer3_outputs(4014)) or (layer3_outputs(7559));
    layer4_outputs(6140) <= (layer3_outputs(1410)) or (layer3_outputs(2681));
    layer4_outputs(6141) <= layer3_outputs(1388);
    layer4_outputs(6142) <= not((layer3_outputs(5282)) xor (layer3_outputs(3430)));
    layer4_outputs(6143) <= not(layer3_outputs(402));
    layer4_outputs(6144) <= not(layer3_outputs(3894)) or (layer3_outputs(5731));
    layer4_outputs(6145) <= (layer3_outputs(123)) and not (layer3_outputs(4655));
    layer4_outputs(6146) <= layer3_outputs(429);
    layer4_outputs(6147) <= not(layer3_outputs(6395));
    layer4_outputs(6148) <= layer3_outputs(6515);
    layer4_outputs(6149) <= not(layer3_outputs(5007));
    layer4_outputs(6150) <= not(layer3_outputs(607)) or (layer3_outputs(343));
    layer4_outputs(6151) <= not(layer3_outputs(217));
    layer4_outputs(6152) <= not((layer3_outputs(450)) xor (layer3_outputs(6295)));
    layer4_outputs(6153) <= '0';
    layer4_outputs(6154) <= not((layer3_outputs(5824)) xor (layer3_outputs(1803)));
    layer4_outputs(6155) <= '0';
    layer4_outputs(6156) <= not(layer3_outputs(3824));
    layer4_outputs(6157) <= not((layer3_outputs(6004)) or (layer3_outputs(7314)));
    layer4_outputs(6158) <= layer3_outputs(41);
    layer4_outputs(6159) <= not((layer3_outputs(2348)) and (layer3_outputs(2814)));
    layer4_outputs(6160) <= layer3_outputs(1601);
    layer4_outputs(6161) <= layer3_outputs(5266);
    layer4_outputs(6162) <= (layer3_outputs(448)) and not (layer3_outputs(5969));
    layer4_outputs(6163) <= layer3_outputs(927);
    layer4_outputs(6164) <= (layer3_outputs(7151)) xor (layer3_outputs(3025));
    layer4_outputs(6165) <= not((layer3_outputs(2414)) or (layer3_outputs(2665)));
    layer4_outputs(6166) <= layer3_outputs(5379);
    layer4_outputs(6167) <= not(layer3_outputs(1027));
    layer4_outputs(6168) <= (layer3_outputs(1991)) xor (layer3_outputs(1735));
    layer4_outputs(6169) <= not(layer3_outputs(642));
    layer4_outputs(6170) <= not(layer3_outputs(7061)) or (layer3_outputs(1487));
    layer4_outputs(6171) <= not(layer3_outputs(2089));
    layer4_outputs(6172) <= (layer3_outputs(917)) and (layer3_outputs(549));
    layer4_outputs(6173) <= not(layer3_outputs(3755));
    layer4_outputs(6174) <= (layer3_outputs(3570)) and (layer3_outputs(5287));
    layer4_outputs(6175) <= not((layer3_outputs(6367)) xor (layer3_outputs(4009)));
    layer4_outputs(6176) <= not(layer3_outputs(1073)) or (layer3_outputs(3680));
    layer4_outputs(6177) <= (layer3_outputs(2563)) xor (layer3_outputs(7));
    layer4_outputs(6178) <= not(layer3_outputs(741));
    layer4_outputs(6179) <= (layer3_outputs(714)) xor (layer3_outputs(5579));
    layer4_outputs(6180) <= not(layer3_outputs(2797)) or (layer3_outputs(6776));
    layer4_outputs(6181) <= (layer3_outputs(5613)) and not (layer3_outputs(4927));
    layer4_outputs(6182) <= '1';
    layer4_outputs(6183) <= not((layer3_outputs(2459)) xor (layer3_outputs(6098)));
    layer4_outputs(6184) <= (layer3_outputs(2902)) or (layer3_outputs(6657));
    layer4_outputs(6185) <= not(layer3_outputs(4634));
    layer4_outputs(6186) <= layer3_outputs(1594);
    layer4_outputs(6187) <= not(layer3_outputs(2585));
    layer4_outputs(6188) <= layer3_outputs(2803);
    layer4_outputs(6189) <= (layer3_outputs(4551)) xor (layer3_outputs(6485));
    layer4_outputs(6190) <= layer3_outputs(5718);
    layer4_outputs(6191) <= (layer3_outputs(6257)) and (layer3_outputs(276));
    layer4_outputs(6192) <= not(layer3_outputs(4540));
    layer4_outputs(6193) <= layer3_outputs(1669);
    layer4_outputs(6194) <= layer3_outputs(2329);
    layer4_outputs(6195) <= (layer3_outputs(6551)) xor (layer3_outputs(6610));
    layer4_outputs(6196) <= layer3_outputs(6220);
    layer4_outputs(6197) <= (layer3_outputs(5352)) or (layer3_outputs(467));
    layer4_outputs(6198) <= (layer3_outputs(2936)) or (layer3_outputs(5590));
    layer4_outputs(6199) <= layer3_outputs(6370);
    layer4_outputs(6200) <= layer3_outputs(4881);
    layer4_outputs(6201) <= layer3_outputs(5172);
    layer4_outputs(6202) <= (layer3_outputs(709)) and not (layer3_outputs(5364));
    layer4_outputs(6203) <= not(layer3_outputs(7168));
    layer4_outputs(6204) <= layer3_outputs(3552);
    layer4_outputs(6205) <= layer3_outputs(227);
    layer4_outputs(6206) <= not(layer3_outputs(1369));
    layer4_outputs(6207) <= not(layer3_outputs(5944));
    layer4_outputs(6208) <= not(layer3_outputs(6245));
    layer4_outputs(6209) <= not((layer3_outputs(6357)) and (layer3_outputs(1917)));
    layer4_outputs(6210) <= (layer3_outputs(190)) and not (layer3_outputs(1736));
    layer4_outputs(6211) <= not(layer3_outputs(546)) or (layer3_outputs(2359));
    layer4_outputs(6212) <= not(layer3_outputs(5865));
    layer4_outputs(6213) <= (layer3_outputs(4178)) or (layer3_outputs(808));
    layer4_outputs(6214) <= not(layer3_outputs(6830));
    layer4_outputs(6215) <= (layer3_outputs(3749)) and (layer3_outputs(4102));
    layer4_outputs(6216) <= (layer3_outputs(2943)) or (layer3_outputs(2015));
    layer4_outputs(6217) <= not(layer3_outputs(5653));
    layer4_outputs(6218) <= layer3_outputs(5359);
    layer4_outputs(6219) <= layer3_outputs(121);
    layer4_outputs(6220) <= layer3_outputs(5178);
    layer4_outputs(6221) <= layer3_outputs(2561);
    layer4_outputs(6222) <= (layer3_outputs(5333)) xor (layer3_outputs(6152));
    layer4_outputs(6223) <= not(layer3_outputs(4902));
    layer4_outputs(6224) <= not(layer3_outputs(5146)) or (layer3_outputs(2737));
    layer4_outputs(6225) <= layer3_outputs(4530);
    layer4_outputs(6226) <= (layer3_outputs(5971)) xor (layer3_outputs(6093));
    layer4_outputs(6227) <= not(layer3_outputs(1468)) or (layer3_outputs(1955));
    layer4_outputs(6228) <= not(layer3_outputs(3231));
    layer4_outputs(6229) <= not(layer3_outputs(1263));
    layer4_outputs(6230) <= not((layer3_outputs(732)) and (layer3_outputs(7534)));
    layer4_outputs(6231) <= layer3_outputs(114);
    layer4_outputs(6232) <= (layer3_outputs(730)) and (layer3_outputs(433));
    layer4_outputs(6233) <= not(layer3_outputs(325));
    layer4_outputs(6234) <= layer3_outputs(1506);
    layer4_outputs(6235) <= layer3_outputs(333);
    layer4_outputs(6236) <= not(layer3_outputs(2920));
    layer4_outputs(6237) <= layer3_outputs(437);
    layer4_outputs(6238) <= not((layer3_outputs(5349)) xor (layer3_outputs(5971)));
    layer4_outputs(6239) <= layer3_outputs(5769);
    layer4_outputs(6240) <= not(layer3_outputs(4326)) or (layer3_outputs(677));
    layer4_outputs(6241) <= not(layer3_outputs(2494));
    layer4_outputs(6242) <= layer3_outputs(215);
    layer4_outputs(6243) <= not(layer3_outputs(4816));
    layer4_outputs(6244) <= (layer3_outputs(3977)) xor (layer3_outputs(6867));
    layer4_outputs(6245) <= not(layer3_outputs(2350)) or (layer3_outputs(3621));
    layer4_outputs(6246) <= not(layer3_outputs(3876));
    layer4_outputs(6247) <= not(layer3_outputs(854));
    layer4_outputs(6248) <= not(layer3_outputs(1965));
    layer4_outputs(6249) <= '1';
    layer4_outputs(6250) <= (layer3_outputs(2256)) or (layer3_outputs(2572));
    layer4_outputs(6251) <= not(layer3_outputs(320));
    layer4_outputs(6252) <= layer3_outputs(6188);
    layer4_outputs(6253) <= (layer3_outputs(6610)) and not (layer3_outputs(5584));
    layer4_outputs(6254) <= not((layer3_outputs(2124)) or (layer3_outputs(4205)));
    layer4_outputs(6255) <= not((layer3_outputs(2224)) and (layer3_outputs(4952)));
    layer4_outputs(6256) <= layer3_outputs(4257);
    layer4_outputs(6257) <= not(layer3_outputs(2561));
    layer4_outputs(6258) <= not(layer3_outputs(6888)) or (layer3_outputs(2018));
    layer4_outputs(6259) <= (layer3_outputs(2371)) or (layer3_outputs(5095));
    layer4_outputs(6260) <= not(layer3_outputs(2643));
    layer4_outputs(6261) <= (layer3_outputs(3546)) xor (layer3_outputs(5622));
    layer4_outputs(6262) <= (layer3_outputs(890)) and not (layer3_outputs(7));
    layer4_outputs(6263) <= not(layer3_outputs(7187));
    layer4_outputs(6264) <= (layer3_outputs(3148)) and (layer3_outputs(1707));
    layer4_outputs(6265) <= layer3_outputs(2395);
    layer4_outputs(6266) <= layer3_outputs(7463);
    layer4_outputs(6267) <= '1';
    layer4_outputs(6268) <= (layer3_outputs(6839)) and not (layer3_outputs(871));
    layer4_outputs(6269) <= (layer3_outputs(1818)) xor (layer3_outputs(5756));
    layer4_outputs(6270) <= not((layer3_outputs(6691)) and (layer3_outputs(3672)));
    layer4_outputs(6271) <= not(layer3_outputs(6910));
    layer4_outputs(6272) <= not((layer3_outputs(5559)) and (layer3_outputs(6391)));
    layer4_outputs(6273) <= (layer3_outputs(2406)) or (layer3_outputs(5514));
    layer4_outputs(6274) <= not(layer3_outputs(6877));
    layer4_outputs(6275) <= (layer3_outputs(3311)) xor (layer3_outputs(126));
    layer4_outputs(6276) <= (layer3_outputs(3663)) and not (layer3_outputs(5374));
    layer4_outputs(6277) <= layer3_outputs(885);
    layer4_outputs(6278) <= (layer3_outputs(3598)) or (layer3_outputs(3774));
    layer4_outputs(6279) <= not((layer3_outputs(2420)) and (layer3_outputs(201)));
    layer4_outputs(6280) <= (layer3_outputs(7281)) or (layer3_outputs(1507));
    layer4_outputs(6281) <= not((layer3_outputs(6123)) and (layer3_outputs(1147)));
    layer4_outputs(6282) <= not((layer3_outputs(5891)) or (layer3_outputs(4234)));
    layer4_outputs(6283) <= layer3_outputs(7090);
    layer4_outputs(6284) <= layer3_outputs(2518);
    layer4_outputs(6285) <= layer3_outputs(6620);
    layer4_outputs(6286) <= not(layer3_outputs(6368));
    layer4_outputs(6287) <= layer3_outputs(4471);
    layer4_outputs(6288) <= not((layer3_outputs(5516)) xor (layer3_outputs(5023)));
    layer4_outputs(6289) <= not(layer3_outputs(7155)) or (layer3_outputs(3195));
    layer4_outputs(6290) <= layer3_outputs(5968);
    layer4_outputs(6291) <= not(layer3_outputs(1009)) or (layer3_outputs(7326));
    layer4_outputs(6292) <= layer3_outputs(5504);
    layer4_outputs(6293) <= not(layer3_outputs(1411));
    layer4_outputs(6294) <= (layer3_outputs(6680)) xor (layer3_outputs(2588));
    layer4_outputs(6295) <= not(layer3_outputs(7309));
    layer4_outputs(6296) <= layer3_outputs(6382);
    layer4_outputs(6297) <= layer3_outputs(6292);
    layer4_outputs(6298) <= not(layer3_outputs(38)) or (layer3_outputs(3170));
    layer4_outputs(6299) <= not(layer3_outputs(4136));
    layer4_outputs(6300) <= layer3_outputs(2792);
    layer4_outputs(6301) <= (layer3_outputs(6714)) xor (layer3_outputs(5294));
    layer4_outputs(6302) <= not(layer3_outputs(7158));
    layer4_outputs(6303) <= not(layer3_outputs(2171));
    layer4_outputs(6304) <= not(layer3_outputs(1229)) or (layer3_outputs(3712));
    layer4_outputs(6305) <= layer3_outputs(859);
    layer4_outputs(6306) <= layer3_outputs(4613);
    layer4_outputs(6307) <= layer3_outputs(3815);
    layer4_outputs(6308) <= (layer3_outputs(3341)) or (layer3_outputs(1340));
    layer4_outputs(6309) <= layer3_outputs(416);
    layer4_outputs(6310) <= not((layer3_outputs(3282)) xor (layer3_outputs(3630)));
    layer4_outputs(6311) <= layer3_outputs(3101);
    layer4_outputs(6312) <= layer3_outputs(4243);
    layer4_outputs(6313) <= not((layer3_outputs(4886)) or (layer3_outputs(2749)));
    layer4_outputs(6314) <= not(layer3_outputs(3114)) or (layer3_outputs(3226));
    layer4_outputs(6315) <= (layer3_outputs(6655)) or (layer3_outputs(7483));
    layer4_outputs(6316) <= layer3_outputs(6586);
    layer4_outputs(6317) <= not(layer3_outputs(7583));
    layer4_outputs(6318) <= (layer3_outputs(4406)) and not (layer3_outputs(3847));
    layer4_outputs(6319) <= not(layer3_outputs(5892));
    layer4_outputs(6320) <= not((layer3_outputs(3111)) and (layer3_outputs(1509)));
    layer4_outputs(6321) <= layer3_outputs(4415);
    layer4_outputs(6322) <= not(layer3_outputs(1974));
    layer4_outputs(6323) <= layer3_outputs(5295);
    layer4_outputs(6324) <= (layer3_outputs(3386)) and not (layer3_outputs(1599));
    layer4_outputs(6325) <= not((layer3_outputs(717)) or (layer3_outputs(5206)));
    layer4_outputs(6326) <= (layer3_outputs(3263)) and not (layer3_outputs(7021));
    layer4_outputs(6327) <= layer3_outputs(3778);
    layer4_outputs(6328) <= layer3_outputs(5090);
    layer4_outputs(6329) <= layer3_outputs(6843);
    layer4_outputs(6330) <= not(layer3_outputs(3259));
    layer4_outputs(6331) <= layer3_outputs(7221);
    layer4_outputs(6332) <= layer3_outputs(2284);
    layer4_outputs(6333) <= (layer3_outputs(4390)) and not (layer3_outputs(4773));
    layer4_outputs(6334) <= not(layer3_outputs(6591));
    layer4_outputs(6335) <= not(layer3_outputs(1557));
    layer4_outputs(6336) <= not((layer3_outputs(4904)) xor (layer3_outputs(2751)));
    layer4_outputs(6337) <= not(layer3_outputs(78));
    layer4_outputs(6338) <= not(layer3_outputs(484));
    layer4_outputs(6339) <= layer3_outputs(911);
    layer4_outputs(6340) <= layer3_outputs(4241);
    layer4_outputs(6341) <= (layer3_outputs(3976)) or (layer3_outputs(4642));
    layer4_outputs(6342) <= not((layer3_outputs(2181)) or (layer3_outputs(3519)));
    layer4_outputs(6343) <= (layer3_outputs(1566)) or (layer3_outputs(3924));
    layer4_outputs(6344) <= not(layer3_outputs(1327)) or (layer3_outputs(2623));
    layer4_outputs(6345) <= (layer3_outputs(5187)) xor (layer3_outputs(4989));
    layer4_outputs(6346) <= not(layer3_outputs(3488));
    layer4_outputs(6347) <= not(layer3_outputs(6392));
    layer4_outputs(6348) <= not(layer3_outputs(3782));
    layer4_outputs(6349) <= (layer3_outputs(1875)) or (layer3_outputs(4750));
    layer4_outputs(6350) <= not(layer3_outputs(2345));
    layer4_outputs(6351) <= not((layer3_outputs(1703)) and (layer3_outputs(3648)));
    layer4_outputs(6352) <= layer3_outputs(6113);
    layer4_outputs(6353) <= layer3_outputs(3360);
    layer4_outputs(6354) <= (layer3_outputs(6452)) and not (layer3_outputs(6554));
    layer4_outputs(6355) <= not(layer3_outputs(5148));
    layer4_outputs(6356) <= not((layer3_outputs(6396)) and (layer3_outputs(6899)));
    layer4_outputs(6357) <= (layer3_outputs(1398)) or (layer3_outputs(3383));
    layer4_outputs(6358) <= not(layer3_outputs(498)) or (layer3_outputs(1636));
    layer4_outputs(6359) <= layer3_outputs(6733);
    layer4_outputs(6360) <= not(layer3_outputs(4587));
    layer4_outputs(6361) <= not(layer3_outputs(5297)) or (layer3_outputs(6261));
    layer4_outputs(6362) <= not((layer3_outputs(4010)) or (layer3_outputs(271)));
    layer4_outputs(6363) <= (layer3_outputs(6695)) and not (layer3_outputs(7177));
    layer4_outputs(6364) <= layer3_outputs(6813);
    layer4_outputs(6365) <= not(layer3_outputs(6272));
    layer4_outputs(6366) <= not(layer3_outputs(478));
    layer4_outputs(6367) <= '0';
    layer4_outputs(6368) <= (layer3_outputs(4682)) or (layer3_outputs(259));
    layer4_outputs(6369) <= not((layer3_outputs(4835)) xor (layer3_outputs(6974)));
    layer4_outputs(6370) <= (layer3_outputs(6705)) and not (layer3_outputs(348));
    layer4_outputs(6371) <= not(layer3_outputs(3573));
    layer4_outputs(6372) <= not((layer3_outputs(650)) xor (layer3_outputs(5664)));
    layer4_outputs(6373) <= not((layer3_outputs(6638)) and (layer3_outputs(1804)));
    layer4_outputs(6374) <= layer3_outputs(1151);
    layer4_outputs(6375) <= not(layer3_outputs(2927));
    layer4_outputs(6376) <= (layer3_outputs(5489)) xor (layer3_outputs(7412));
    layer4_outputs(6377) <= layer3_outputs(6819);
    layer4_outputs(6378) <= not((layer3_outputs(5321)) or (layer3_outputs(1592)));
    layer4_outputs(6379) <= not((layer3_outputs(7100)) or (layer3_outputs(4978)));
    layer4_outputs(6380) <= not(layer3_outputs(1298)) or (layer3_outputs(5312));
    layer4_outputs(6381) <= not(layer3_outputs(4739));
    layer4_outputs(6382) <= layer3_outputs(6142);
    layer4_outputs(6383) <= layer3_outputs(6839);
    layer4_outputs(6384) <= not((layer3_outputs(4606)) and (layer3_outputs(1074)));
    layer4_outputs(6385) <= not(layer3_outputs(4051));
    layer4_outputs(6386) <= not(layer3_outputs(1905)) or (layer3_outputs(3575));
    layer4_outputs(6387) <= not(layer3_outputs(7393));
    layer4_outputs(6388) <= layer3_outputs(7339);
    layer4_outputs(6389) <= (layer3_outputs(6614)) and (layer3_outputs(1582));
    layer4_outputs(6390) <= (layer3_outputs(6372)) or (layer3_outputs(4466));
    layer4_outputs(6391) <= not(layer3_outputs(4219));
    layer4_outputs(6392) <= not(layer3_outputs(5169));
    layer4_outputs(6393) <= (layer3_outputs(1880)) and not (layer3_outputs(1475));
    layer4_outputs(6394) <= layer3_outputs(7166);
    layer4_outputs(6395) <= not((layer3_outputs(6983)) and (layer3_outputs(6849)));
    layer4_outputs(6396) <= (layer3_outputs(6990)) xor (layer3_outputs(6348));
    layer4_outputs(6397) <= not(layer3_outputs(3442));
    layer4_outputs(6398) <= not(layer3_outputs(5730)) or (layer3_outputs(1850));
    layer4_outputs(6399) <= layer3_outputs(6876);
    layer4_outputs(6400) <= not(layer3_outputs(4447));
    layer4_outputs(6401) <= (layer3_outputs(1821)) and (layer3_outputs(2567));
    layer4_outputs(6402) <= (layer3_outputs(6976)) and not (layer3_outputs(5421));
    layer4_outputs(6403) <= not(layer3_outputs(4738));
    layer4_outputs(6404) <= layer3_outputs(3367);
    layer4_outputs(6405) <= not(layer3_outputs(177));
    layer4_outputs(6406) <= not(layer3_outputs(4834));
    layer4_outputs(6407) <= layer3_outputs(3931);
    layer4_outputs(6408) <= (layer3_outputs(2642)) and not (layer3_outputs(7537));
    layer4_outputs(6409) <= (layer3_outputs(2316)) and not (layer3_outputs(6841));
    layer4_outputs(6410) <= layer3_outputs(7521);
    layer4_outputs(6411) <= layer3_outputs(4225);
    layer4_outputs(6412) <= (layer3_outputs(762)) and (layer3_outputs(2775));
    layer4_outputs(6413) <= not(layer3_outputs(1234));
    layer4_outputs(6414) <= not((layer3_outputs(1304)) and (layer3_outputs(385)));
    layer4_outputs(6415) <= not(layer3_outputs(2931)) or (layer3_outputs(1346));
    layer4_outputs(6416) <= (layer3_outputs(2336)) and not (layer3_outputs(6878));
    layer4_outputs(6417) <= layer3_outputs(781);
    layer4_outputs(6418) <= not((layer3_outputs(7163)) xor (layer3_outputs(6913)));
    layer4_outputs(6419) <= layer3_outputs(2339);
    layer4_outputs(6420) <= (layer3_outputs(5178)) and not (layer3_outputs(73));
    layer4_outputs(6421) <= not(layer3_outputs(2423));
    layer4_outputs(6422) <= not(layer3_outputs(638)) or (layer3_outputs(426));
    layer4_outputs(6423) <= not(layer3_outputs(1530)) or (layer3_outputs(1608));
    layer4_outputs(6424) <= layer3_outputs(4262);
    layer4_outputs(6425) <= not(layer3_outputs(2081)) or (layer3_outputs(7524));
    layer4_outputs(6426) <= layer3_outputs(6589);
    layer4_outputs(6427) <= (layer3_outputs(1523)) or (layer3_outputs(2069));
    layer4_outputs(6428) <= layer3_outputs(1686);
    layer4_outputs(6429) <= not(layer3_outputs(866)) or (layer3_outputs(1037));
    layer4_outputs(6430) <= not((layer3_outputs(2827)) xor (layer3_outputs(4024)));
    layer4_outputs(6431) <= not(layer3_outputs(5326));
    layer4_outputs(6432) <= layer3_outputs(3712);
    layer4_outputs(6433) <= layer3_outputs(1325);
    layer4_outputs(6434) <= not(layer3_outputs(2282));
    layer4_outputs(6435) <= not(layer3_outputs(1462));
    layer4_outputs(6436) <= not(layer3_outputs(5966));
    layer4_outputs(6437) <= (layer3_outputs(7341)) and not (layer3_outputs(190));
    layer4_outputs(6438) <= not((layer3_outputs(3753)) or (layer3_outputs(4646)));
    layer4_outputs(6439) <= layer3_outputs(2262);
    layer4_outputs(6440) <= not((layer3_outputs(2514)) or (layer3_outputs(3306)));
    layer4_outputs(6441) <= (layer3_outputs(2095)) and (layer3_outputs(193));
    layer4_outputs(6442) <= '0';
    layer4_outputs(6443) <= not(layer3_outputs(6954));
    layer4_outputs(6444) <= (layer3_outputs(3654)) or (layer3_outputs(4201));
    layer4_outputs(6445) <= layer3_outputs(4195);
    layer4_outputs(6446) <= not((layer3_outputs(558)) or (layer3_outputs(6505)));
    layer4_outputs(6447) <= not((layer3_outputs(4999)) or (layer3_outputs(1412)));
    layer4_outputs(6448) <= layer3_outputs(2057);
    layer4_outputs(6449) <= not(layer3_outputs(2585));
    layer4_outputs(6450) <= not(layer3_outputs(7282));
    layer4_outputs(6451) <= layer3_outputs(5347);
    layer4_outputs(6452) <= not(layer3_outputs(3050));
    layer4_outputs(6453) <= (layer3_outputs(4892)) and (layer3_outputs(1308));
    layer4_outputs(6454) <= not((layer3_outputs(2020)) and (layer3_outputs(2807)));
    layer4_outputs(6455) <= not(layer3_outputs(6590));
    layer4_outputs(6456) <= layer3_outputs(2010);
    layer4_outputs(6457) <= not(layer3_outputs(5642));
    layer4_outputs(6458) <= not(layer3_outputs(1437));
    layer4_outputs(6459) <= not(layer3_outputs(7423));
    layer4_outputs(6460) <= layer3_outputs(5467);
    layer4_outputs(6461) <= (layer3_outputs(2687)) and (layer3_outputs(754));
    layer4_outputs(6462) <= (layer3_outputs(1155)) and not (layer3_outputs(3296));
    layer4_outputs(6463) <= layer3_outputs(5515);
    layer4_outputs(6464) <= not((layer3_outputs(991)) or (layer3_outputs(2713)));
    layer4_outputs(6465) <= (layer3_outputs(1454)) or (layer3_outputs(1846));
    layer4_outputs(6466) <= not(layer3_outputs(2719)) or (layer3_outputs(4755));
    layer4_outputs(6467) <= not((layer3_outputs(1680)) or (layer3_outputs(482)));
    layer4_outputs(6468) <= (layer3_outputs(4568)) and not (layer3_outputs(7360));
    layer4_outputs(6469) <= not(layer3_outputs(58));
    layer4_outputs(6470) <= not(layer3_outputs(6470));
    layer4_outputs(6471) <= not((layer3_outputs(3096)) and (layer3_outputs(3817)));
    layer4_outputs(6472) <= layer3_outputs(370);
    layer4_outputs(6473) <= (layer3_outputs(6337)) or (layer3_outputs(7183));
    layer4_outputs(6474) <= (layer3_outputs(1750)) and not (layer3_outputs(2322));
    layer4_outputs(6475) <= layer3_outputs(194);
    layer4_outputs(6476) <= not(layer3_outputs(1367));
    layer4_outputs(6477) <= not(layer3_outputs(5372));
    layer4_outputs(6478) <= not((layer3_outputs(5221)) or (layer3_outputs(654)));
    layer4_outputs(6479) <= (layer3_outputs(1021)) xor (layer3_outputs(682));
    layer4_outputs(6480) <= layer3_outputs(4378);
    layer4_outputs(6481) <= layer3_outputs(4892);
    layer4_outputs(6482) <= layer3_outputs(5948);
    layer4_outputs(6483) <= not(layer3_outputs(2914)) or (layer3_outputs(5393));
    layer4_outputs(6484) <= layer3_outputs(1905);
    layer4_outputs(6485) <= layer3_outputs(3529);
    layer4_outputs(6486) <= (layer3_outputs(4271)) and (layer3_outputs(1537));
    layer4_outputs(6487) <= not(layer3_outputs(5620)) or (layer3_outputs(711));
    layer4_outputs(6488) <= not(layer3_outputs(7677));
    layer4_outputs(6489) <= not((layer3_outputs(6403)) and (layer3_outputs(5068)));
    layer4_outputs(6490) <= not(layer3_outputs(4889)) or (layer3_outputs(4171));
    layer4_outputs(6491) <= layer3_outputs(3440);
    layer4_outputs(6492) <= not(layer3_outputs(1743)) or (layer3_outputs(3618));
    layer4_outputs(6493) <= not((layer3_outputs(1970)) and (layer3_outputs(6724)));
    layer4_outputs(6494) <= (layer3_outputs(5899)) and not (layer3_outputs(6960));
    layer4_outputs(6495) <= not((layer3_outputs(5113)) xor (layer3_outputs(2144)));
    layer4_outputs(6496) <= not(layer3_outputs(6501)) or (layer3_outputs(6350));
    layer4_outputs(6497) <= not((layer3_outputs(802)) xor (layer3_outputs(97)));
    layer4_outputs(6498) <= layer3_outputs(7605);
    layer4_outputs(6499) <= (layer3_outputs(664)) and not (layer3_outputs(1091));
    layer4_outputs(6500) <= (layer3_outputs(6906)) and (layer3_outputs(4551));
    layer4_outputs(6501) <= not(layer3_outputs(106));
    layer4_outputs(6502) <= layer3_outputs(695);
    layer4_outputs(6503) <= layer3_outputs(1604);
    layer4_outputs(6504) <= (layer3_outputs(351)) and not (layer3_outputs(7660));
    layer4_outputs(6505) <= layer3_outputs(5486);
    layer4_outputs(6506) <= not(layer3_outputs(6848));
    layer4_outputs(6507) <= not(layer3_outputs(2826));
    layer4_outputs(6508) <= not(layer3_outputs(2369));
    layer4_outputs(6509) <= layer3_outputs(6481);
    layer4_outputs(6510) <= not(layer3_outputs(4707));
    layer4_outputs(6511) <= not(layer3_outputs(5131));
    layer4_outputs(6512) <= not((layer3_outputs(6241)) or (layer3_outputs(6837)));
    layer4_outputs(6513) <= layer3_outputs(6606);
    layer4_outputs(6514) <= (layer3_outputs(2596)) xor (layer3_outputs(353));
    layer4_outputs(6515) <= (layer3_outputs(4346)) xor (layer3_outputs(2540));
    layer4_outputs(6516) <= not(layer3_outputs(2671)) or (layer3_outputs(4639));
    layer4_outputs(6517) <= (layer3_outputs(4352)) xor (layer3_outputs(6047));
    layer4_outputs(6518) <= layer3_outputs(197);
    layer4_outputs(6519) <= not(layer3_outputs(2149));
    layer4_outputs(6520) <= (layer3_outputs(4112)) and (layer3_outputs(4569));
    layer4_outputs(6521) <= (layer3_outputs(948)) xor (layer3_outputs(3975));
    layer4_outputs(6522) <= not(layer3_outputs(5199));
    layer4_outputs(6523) <= not((layer3_outputs(5742)) xor (layer3_outputs(1662)));
    layer4_outputs(6524) <= not((layer3_outputs(7669)) and (layer3_outputs(6580)));
    layer4_outputs(6525) <= (layer3_outputs(1520)) and not (layer3_outputs(2835));
    layer4_outputs(6526) <= not(layer3_outputs(3)) or (layer3_outputs(5935));
    layer4_outputs(6527) <= layer3_outputs(1416);
    layer4_outputs(6528) <= layer3_outputs(5989);
    layer4_outputs(6529) <= not(layer3_outputs(7570));
    layer4_outputs(6530) <= layer3_outputs(5047);
    layer4_outputs(6531) <= not(layer3_outputs(3964)) or (layer3_outputs(2742));
    layer4_outputs(6532) <= layer3_outputs(3540);
    layer4_outputs(6533) <= not((layer3_outputs(1977)) xor (layer3_outputs(182)));
    layer4_outputs(6534) <= layer3_outputs(6307);
    layer4_outputs(6535) <= layer3_outputs(2174);
    layer4_outputs(6536) <= '0';
    layer4_outputs(6537) <= (layer3_outputs(6492)) and not (layer3_outputs(6234));
    layer4_outputs(6538) <= (layer3_outputs(1187)) and (layer3_outputs(772));
    layer4_outputs(6539) <= layer3_outputs(6375);
    layer4_outputs(6540) <= (layer3_outputs(224)) and (layer3_outputs(6145));
    layer4_outputs(6541) <= layer3_outputs(1957);
    layer4_outputs(6542) <= not(layer3_outputs(5130));
    layer4_outputs(6543) <= not((layer3_outputs(5116)) xor (layer3_outputs(1782)));
    layer4_outputs(6544) <= not(layer3_outputs(5469));
    layer4_outputs(6545) <= not(layer3_outputs(6516));
    layer4_outputs(6546) <= not((layer3_outputs(7500)) xor (layer3_outputs(5537)));
    layer4_outputs(6547) <= layer3_outputs(2388);
    layer4_outputs(6548) <= (layer3_outputs(3775)) and not (layer3_outputs(988));
    layer4_outputs(6549) <= not(layer3_outputs(140));
    layer4_outputs(6550) <= (layer3_outputs(5080)) and (layer3_outputs(2315));
    layer4_outputs(6551) <= not((layer3_outputs(1067)) or (layer3_outputs(6354)));
    layer4_outputs(6552) <= (layer3_outputs(1643)) and not (layer3_outputs(1458));
    layer4_outputs(6553) <= not((layer3_outputs(358)) and (layer3_outputs(5266)));
    layer4_outputs(6554) <= layer3_outputs(3943);
    layer4_outputs(6555) <= not(layer3_outputs(7667));
    layer4_outputs(6556) <= layer3_outputs(6983);
    layer4_outputs(6557) <= not(layer3_outputs(3798));
    layer4_outputs(6558) <= (layer3_outputs(746)) and not (layer3_outputs(7624));
    layer4_outputs(6559) <= not(layer3_outputs(5609)) or (layer3_outputs(366));
    layer4_outputs(6560) <= (layer3_outputs(6340)) xor (layer3_outputs(7366));
    layer4_outputs(6561) <= (layer3_outputs(5703)) or (layer3_outputs(5797));
    layer4_outputs(6562) <= not((layer3_outputs(7115)) or (layer3_outputs(4115)));
    layer4_outputs(6563) <= layer3_outputs(4566);
    layer4_outputs(6564) <= (layer3_outputs(6212)) and not (layer3_outputs(3660));
    layer4_outputs(6565) <= (layer3_outputs(1288)) xor (layer3_outputs(7297));
    layer4_outputs(6566) <= (layer3_outputs(598)) xor (layer3_outputs(6218));
    layer4_outputs(6567) <= (layer3_outputs(4554)) or (layer3_outputs(1870));
    layer4_outputs(6568) <= (layer3_outputs(4619)) and not (layer3_outputs(3844));
    layer4_outputs(6569) <= not(layer3_outputs(7481));
    layer4_outputs(6570) <= layer3_outputs(5881);
    layer4_outputs(6571) <= (layer3_outputs(5334)) xor (layer3_outputs(6730));
    layer4_outputs(6572) <= not((layer3_outputs(1477)) and (layer3_outputs(7527)));
    layer4_outputs(6573) <= '1';
    layer4_outputs(6574) <= layer3_outputs(7086);
    layer4_outputs(6575) <= '0';
    layer4_outputs(6576) <= not(layer3_outputs(3968));
    layer4_outputs(6577) <= layer3_outputs(3590);
    layer4_outputs(6578) <= layer3_outputs(2608);
    layer4_outputs(6579) <= layer3_outputs(7131);
    layer4_outputs(6580) <= (layer3_outputs(2041)) xor (layer3_outputs(2261));
    layer4_outputs(6581) <= layer3_outputs(7607);
    layer4_outputs(6582) <= not(layer3_outputs(429));
    layer4_outputs(6583) <= layer3_outputs(2521);
    layer4_outputs(6584) <= not(layer3_outputs(4149));
    layer4_outputs(6585) <= layer3_outputs(111);
    layer4_outputs(6586) <= (layer3_outputs(3064)) and not (layer3_outputs(5236));
    layer4_outputs(6587) <= (layer3_outputs(639)) xor (layer3_outputs(5147));
    layer4_outputs(6588) <= not(layer3_outputs(735));
    layer4_outputs(6589) <= (layer3_outputs(7230)) or (layer3_outputs(7511));
    layer4_outputs(6590) <= layer3_outputs(6480);
    layer4_outputs(6591) <= not(layer3_outputs(7545));
    layer4_outputs(6592) <= not((layer3_outputs(4865)) or (layer3_outputs(6860)));
    layer4_outputs(6593) <= layer3_outputs(2977);
    layer4_outputs(6594) <= (layer3_outputs(6818)) xor (layer3_outputs(289));
    layer4_outputs(6595) <= layer3_outputs(1164);
    layer4_outputs(6596) <= not((layer3_outputs(908)) or (layer3_outputs(6896)));
    layer4_outputs(6597) <= (layer3_outputs(6458)) and not (layer3_outputs(1930));
    layer4_outputs(6598) <= layer3_outputs(3210);
    layer4_outputs(6599) <= not(layer3_outputs(7569));
    layer4_outputs(6600) <= layer3_outputs(5474);
    layer4_outputs(6601) <= (layer3_outputs(6891)) xor (layer3_outputs(1158));
    layer4_outputs(6602) <= '0';
    layer4_outputs(6603) <= not((layer3_outputs(5406)) or (layer3_outputs(4105)));
    layer4_outputs(6604) <= not(layer3_outputs(5485));
    layer4_outputs(6605) <= not((layer3_outputs(7058)) or (layer3_outputs(3250)));
    layer4_outputs(6606) <= not(layer3_outputs(7095));
    layer4_outputs(6607) <= not((layer3_outputs(6645)) or (layer3_outputs(2137)));
    layer4_outputs(6608) <= not(layer3_outputs(5951)) or (layer3_outputs(1521));
    layer4_outputs(6609) <= layer3_outputs(1800);
    layer4_outputs(6610) <= not(layer3_outputs(5019)) or (layer3_outputs(6196));
    layer4_outputs(6611) <= layer3_outputs(6567);
    layer4_outputs(6612) <= layer3_outputs(4723);
    layer4_outputs(6613) <= (layer3_outputs(6837)) or (layer3_outputs(930));
    layer4_outputs(6614) <= not(layer3_outputs(6541));
    layer4_outputs(6615) <= layer3_outputs(4900);
    layer4_outputs(6616) <= layer3_outputs(1899);
    layer4_outputs(6617) <= '1';
    layer4_outputs(6618) <= (layer3_outputs(6899)) xor (layer3_outputs(1593));
    layer4_outputs(6619) <= (layer3_outputs(6018)) and (layer3_outputs(2202));
    layer4_outputs(6620) <= not(layer3_outputs(6077));
    layer4_outputs(6621) <= (layer3_outputs(4939)) xor (layer3_outputs(7466));
    layer4_outputs(6622) <= not(layer3_outputs(1602));
    layer4_outputs(6623) <= layer3_outputs(5127);
    layer4_outputs(6624) <= layer3_outputs(981);
    layer4_outputs(6625) <= layer3_outputs(6617);
    layer4_outputs(6626) <= (layer3_outputs(6440)) and (layer3_outputs(707));
    layer4_outputs(6627) <= not((layer3_outputs(5135)) or (layer3_outputs(5285)));
    layer4_outputs(6628) <= (layer3_outputs(6648)) and (layer3_outputs(1702));
    layer4_outputs(6629) <= layer3_outputs(9);
    layer4_outputs(6630) <= layer3_outputs(3272);
    layer4_outputs(6631) <= layer3_outputs(6329);
    layer4_outputs(6632) <= not(layer3_outputs(5236));
    layer4_outputs(6633) <= not(layer3_outputs(5434));
    layer4_outputs(6634) <= not(layer3_outputs(7477));
    layer4_outputs(6635) <= (layer3_outputs(207)) xor (layer3_outputs(2471));
    layer4_outputs(6636) <= layer3_outputs(2400);
    layer4_outputs(6637) <= not(layer3_outputs(4590));
    layer4_outputs(6638) <= not(layer3_outputs(7089));
    layer4_outputs(6639) <= layer3_outputs(6557);
    layer4_outputs(6640) <= not((layer3_outputs(3063)) and (layer3_outputs(3799)));
    layer4_outputs(6641) <= '1';
    layer4_outputs(6642) <= (layer3_outputs(2669)) or (layer3_outputs(5027));
    layer4_outputs(6643) <= not(layer3_outputs(4699)) or (layer3_outputs(1927));
    layer4_outputs(6644) <= (layer3_outputs(2484)) and not (layer3_outputs(5260));
    layer4_outputs(6645) <= (layer3_outputs(5949)) and not (layer3_outputs(6704));
    layer4_outputs(6646) <= not(layer3_outputs(6749));
    layer4_outputs(6647) <= not((layer3_outputs(266)) and (layer3_outputs(2117)));
    layer4_outputs(6648) <= layer3_outputs(412);
    layer4_outputs(6649) <= (layer3_outputs(279)) or (layer3_outputs(6933));
    layer4_outputs(6650) <= not((layer3_outputs(4042)) and (layer3_outputs(2767)));
    layer4_outputs(6651) <= not((layer3_outputs(4013)) and (layer3_outputs(6487)));
    layer4_outputs(6652) <= (layer3_outputs(4431)) and not (layer3_outputs(2385));
    layer4_outputs(6653) <= (layer3_outputs(4155)) xor (layer3_outputs(6325));
    layer4_outputs(6654) <= layer3_outputs(6726);
    layer4_outputs(6655) <= not(layer3_outputs(4282)) or (layer3_outputs(2776));
    layer4_outputs(6656) <= not(layer3_outputs(2819));
    layer4_outputs(6657) <= not(layer3_outputs(2431));
    layer4_outputs(6658) <= (layer3_outputs(5708)) or (layer3_outputs(5679));
    layer4_outputs(6659) <= layer3_outputs(4571);
    layer4_outputs(6660) <= layer3_outputs(3609);
    layer4_outputs(6661) <= not((layer3_outputs(3466)) xor (layer3_outputs(1572)));
    layer4_outputs(6662) <= not((layer3_outputs(3541)) xor (layer3_outputs(2702)));
    layer4_outputs(6663) <= layer3_outputs(2250);
    layer4_outputs(6664) <= not(layer3_outputs(5953));
    layer4_outputs(6665) <= not(layer3_outputs(6701));
    layer4_outputs(6666) <= not(layer3_outputs(2003));
    layer4_outputs(6667) <= not((layer3_outputs(5057)) xor (layer3_outputs(4790)));
    layer4_outputs(6668) <= '1';
    layer4_outputs(6669) <= (layer3_outputs(7614)) and not (layer3_outputs(6076));
    layer4_outputs(6670) <= layer3_outputs(3490);
    layer4_outputs(6671) <= not(layer3_outputs(242)) or (layer3_outputs(2656));
    layer4_outputs(6672) <= layer3_outputs(3842);
    layer4_outputs(6673) <= layer3_outputs(1518);
    layer4_outputs(6674) <= not(layer3_outputs(651));
    layer4_outputs(6675) <= not(layer3_outputs(4408)) or (layer3_outputs(3357));
    layer4_outputs(6676) <= not(layer3_outputs(1255));
    layer4_outputs(6677) <= layer3_outputs(3827);
    layer4_outputs(6678) <= layer3_outputs(4425);
    layer4_outputs(6679) <= layer3_outputs(4277);
    layer4_outputs(6680) <= layer3_outputs(531);
    layer4_outputs(6681) <= layer3_outputs(6553);
    layer4_outputs(6682) <= (layer3_outputs(2246)) and not (layer3_outputs(7579));
    layer4_outputs(6683) <= (layer3_outputs(4198)) and not (layer3_outputs(4324));
    layer4_outputs(6684) <= not(layer3_outputs(1591));
    layer4_outputs(6685) <= layer3_outputs(1393);
    layer4_outputs(6686) <= layer3_outputs(1285);
    layer4_outputs(6687) <= not(layer3_outputs(326)) or (layer3_outputs(3343));
    layer4_outputs(6688) <= not(layer3_outputs(5408));
    layer4_outputs(6689) <= layer3_outputs(4365);
    layer4_outputs(6690) <= (layer3_outputs(6586)) and not (layer3_outputs(269));
    layer4_outputs(6691) <= not((layer3_outputs(4127)) or (layer3_outputs(3388)));
    layer4_outputs(6692) <= not(layer3_outputs(7247));
    layer4_outputs(6693) <= (layer3_outputs(6446)) xor (layer3_outputs(5076));
    layer4_outputs(6694) <= not(layer3_outputs(4962)) or (layer3_outputs(2427));
    layer4_outputs(6695) <= not((layer3_outputs(5822)) and (layer3_outputs(2075)));
    layer4_outputs(6696) <= layer3_outputs(2659);
    layer4_outputs(6697) <= layer3_outputs(4951);
    layer4_outputs(6698) <= layer3_outputs(3889);
    layer4_outputs(6699) <= layer3_outputs(4430);
    layer4_outputs(6700) <= not((layer3_outputs(6999)) and (layer3_outputs(3846)));
    layer4_outputs(6701) <= (layer3_outputs(5163)) and not (layer3_outputs(406));
    layer4_outputs(6702) <= not((layer3_outputs(5132)) xor (layer3_outputs(4468)));
    layer4_outputs(6703) <= (layer3_outputs(1755)) and not (layer3_outputs(3697));
    layer4_outputs(6704) <= not(layer3_outputs(2260));
    layer4_outputs(6705) <= not(layer3_outputs(7115));
    layer4_outputs(6706) <= layer3_outputs(2226);
    layer4_outputs(6707) <= layer3_outputs(4218);
    layer4_outputs(6708) <= not(layer3_outputs(7037));
    layer4_outputs(6709) <= not(layer3_outputs(185));
    layer4_outputs(6710) <= (layer3_outputs(5589)) and not (layer3_outputs(6575));
    layer4_outputs(6711) <= (layer3_outputs(6744)) xor (layer3_outputs(695));
    layer4_outputs(6712) <= '0';
    layer4_outputs(6713) <= (layer3_outputs(6833)) and (layer3_outputs(2198));
    layer4_outputs(6714) <= layer3_outputs(7616);
    layer4_outputs(6715) <= not((layer3_outputs(1045)) and (layer3_outputs(48)));
    layer4_outputs(6716) <= layer3_outputs(4395);
    layer4_outputs(6717) <= not((layer3_outputs(2391)) and (layer3_outputs(5793)));
    layer4_outputs(6718) <= layer3_outputs(309);
    layer4_outputs(6719) <= layer3_outputs(802);
    layer4_outputs(6720) <= (layer3_outputs(2809)) and not (layer3_outputs(1440));
    layer4_outputs(6721) <= not(layer3_outputs(4899));
    layer4_outputs(6722) <= not(layer3_outputs(5034));
    layer4_outputs(6723) <= layer3_outputs(4932);
    layer4_outputs(6724) <= (layer3_outputs(6026)) and not (layer3_outputs(6215));
    layer4_outputs(6725) <= not(layer3_outputs(2368));
    layer4_outputs(6726) <= not(layer3_outputs(3787));
    layer4_outputs(6727) <= (layer3_outputs(1235)) or (layer3_outputs(3680));
    layer4_outputs(6728) <= layer3_outputs(2231);
    layer4_outputs(6729) <= not(layer3_outputs(342)) or (layer3_outputs(2621));
    layer4_outputs(6730) <= not(layer3_outputs(2169));
    layer4_outputs(6731) <= (layer3_outputs(3631)) or (layer3_outputs(2131));
    layer4_outputs(6732) <= (layer3_outputs(3729)) or (layer3_outputs(33));
    layer4_outputs(6733) <= layer3_outputs(4124);
    layer4_outputs(6734) <= layer3_outputs(4751);
    layer4_outputs(6735) <= (layer3_outputs(2671)) and (layer3_outputs(6057));
    layer4_outputs(6736) <= not(layer3_outputs(2167)) or (layer3_outputs(2429));
    layer4_outputs(6737) <= not(layer3_outputs(4260));
    layer4_outputs(6738) <= layer3_outputs(3988);
    layer4_outputs(6739) <= (layer3_outputs(2331)) and (layer3_outputs(3285));
    layer4_outputs(6740) <= not(layer3_outputs(1816));
    layer4_outputs(6741) <= not(layer3_outputs(4086));
    layer4_outputs(6742) <= (layer3_outputs(6939)) and not (layer3_outputs(755));
    layer4_outputs(6743) <= not(layer3_outputs(6671));
    layer4_outputs(6744) <= (layer3_outputs(4500)) and not (layer3_outputs(1616));
    layer4_outputs(6745) <= not((layer3_outputs(4755)) xor (layer3_outputs(6897)));
    layer4_outputs(6746) <= layer3_outputs(4494);
    layer4_outputs(6747) <= not(layer3_outputs(5733)) or (layer3_outputs(6041));
    layer4_outputs(6748) <= (layer3_outputs(2148)) or (layer3_outputs(6583));
    layer4_outputs(6749) <= not(layer3_outputs(2532));
    layer4_outputs(6750) <= not((layer3_outputs(1753)) or (layer3_outputs(250)));
    layer4_outputs(6751) <= not((layer3_outputs(365)) xor (layer3_outputs(226)));
    layer4_outputs(6752) <= not(layer3_outputs(6297));
    layer4_outputs(6753) <= (layer3_outputs(7495)) and not (layer3_outputs(7039));
    layer4_outputs(6754) <= layer3_outputs(6919);
    layer4_outputs(6755) <= layer3_outputs(3887);
    layer4_outputs(6756) <= not(layer3_outputs(4125));
    layer4_outputs(6757) <= (layer3_outputs(1484)) or (layer3_outputs(2389));
    layer4_outputs(6758) <= (layer3_outputs(1738)) and not (layer3_outputs(5391));
    layer4_outputs(6759) <= layer3_outputs(454);
    layer4_outputs(6760) <= (layer3_outputs(6293)) and (layer3_outputs(758));
    layer4_outputs(6761) <= layer3_outputs(7546);
    layer4_outputs(6762) <= layer3_outputs(934);
    layer4_outputs(6763) <= layer3_outputs(4325);
    layer4_outputs(6764) <= (layer3_outputs(372)) and not (layer3_outputs(5173));
    layer4_outputs(6765) <= layer3_outputs(3422);
    layer4_outputs(6766) <= layer3_outputs(2183);
    layer4_outputs(6767) <= layer3_outputs(3289);
    layer4_outputs(6768) <= (layer3_outputs(6881)) xor (layer3_outputs(932));
    layer4_outputs(6769) <= (layer3_outputs(4617)) and (layer3_outputs(6033));
    layer4_outputs(6770) <= (layer3_outputs(5057)) xor (layer3_outputs(245));
    layer4_outputs(6771) <= layer3_outputs(7418);
    layer4_outputs(6772) <= (layer3_outputs(2954)) xor (layer3_outputs(3387));
    layer4_outputs(6773) <= (layer3_outputs(2967)) or (layer3_outputs(7011));
    layer4_outputs(6774) <= layer3_outputs(2247);
    layer4_outputs(6775) <= (layer3_outputs(910)) and not (layer3_outputs(228));
    layer4_outputs(6776) <= layer3_outputs(476);
    layer4_outputs(6777) <= not(layer3_outputs(6277)) or (layer3_outputs(330));
    layer4_outputs(6778) <= not(layer3_outputs(936));
    layer4_outputs(6779) <= not(layer3_outputs(2387));
    layer4_outputs(6780) <= layer3_outputs(4716);
    layer4_outputs(6781) <= not(layer3_outputs(865));
    layer4_outputs(6782) <= not(layer3_outputs(3038));
    layer4_outputs(6783) <= layer3_outputs(3350);
    layer4_outputs(6784) <= (layer3_outputs(676)) and (layer3_outputs(318));
    layer4_outputs(6785) <= not(layer3_outputs(4158));
    layer4_outputs(6786) <= layer3_outputs(3661);
    layer4_outputs(6787) <= not(layer3_outputs(4096));
    layer4_outputs(6788) <= not(layer3_outputs(5711)) or (layer3_outputs(6791));
    layer4_outputs(6789) <= not((layer3_outputs(5993)) xor (layer3_outputs(480)));
    layer4_outputs(6790) <= not((layer3_outputs(6014)) or (layer3_outputs(114)));
    layer4_outputs(6791) <= layer3_outputs(1193);
    layer4_outputs(6792) <= layer3_outputs(4853);
    layer4_outputs(6793) <= layer3_outputs(2478);
    layer4_outputs(6794) <= not(layer3_outputs(2244));
    layer4_outputs(6795) <= layer3_outputs(2833);
    layer4_outputs(6796) <= not(layer3_outputs(3775));
    layer4_outputs(6797) <= layer3_outputs(6217);
    layer4_outputs(6798) <= (layer3_outputs(4841)) and (layer3_outputs(4470));
    layer4_outputs(6799) <= not(layer3_outputs(2623)) or (layer3_outputs(7443));
    layer4_outputs(6800) <= not(layer3_outputs(384));
    layer4_outputs(6801) <= (layer3_outputs(5369)) and not (layer3_outputs(3941));
    layer4_outputs(6802) <= layer3_outputs(1656);
    layer4_outputs(6803) <= '1';
    layer4_outputs(6804) <= '1';
    layer4_outputs(6805) <= not((layer3_outputs(1746)) xor (layer3_outputs(658)));
    layer4_outputs(6806) <= (layer3_outputs(5210)) and (layer3_outputs(7075));
    layer4_outputs(6807) <= (layer3_outputs(6895)) xor (layer3_outputs(3323));
    layer4_outputs(6808) <= not(layer3_outputs(6030));
    layer4_outputs(6809) <= (layer3_outputs(3735)) and (layer3_outputs(4432));
    layer4_outputs(6810) <= not(layer3_outputs(3254)) or (layer3_outputs(6657));
    layer4_outputs(6811) <= layer3_outputs(1655);
    layer4_outputs(6812) <= not(layer3_outputs(798)) or (layer3_outputs(4644));
    layer4_outputs(6813) <= layer3_outputs(5500);
    layer4_outputs(6814) <= not(layer3_outputs(1727));
    layer4_outputs(6815) <= (layer3_outputs(1928)) and not (layer3_outputs(80));
    layer4_outputs(6816) <= not(layer3_outputs(5106));
    layer4_outputs(6817) <= not(layer3_outputs(1886));
    layer4_outputs(6818) <= not(layer3_outputs(7167));
    layer4_outputs(6819) <= not((layer3_outputs(3279)) and (layer3_outputs(8)));
    layer4_outputs(6820) <= layer3_outputs(6032);
    layer4_outputs(6821) <= layer3_outputs(2344);
    layer4_outputs(6822) <= not((layer3_outputs(164)) or (layer3_outputs(3039)));
    layer4_outputs(6823) <= not(layer3_outputs(3744)) or (layer3_outputs(2028));
    layer4_outputs(6824) <= not((layer3_outputs(7634)) or (layer3_outputs(1946)));
    layer4_outputs(6825) <= not((layer3_outputs(1204)) or (layer3_outputs(3559)));
    layer4_outputs(6826) <= not(layer3_outputs(3028)) or (layer3_outputs(6836));
    layer4_outputs(6827) <= (layer3_outputs(1960)) xor (layer3_outputs(7185));
    layer4_outputs(6828) <= not(layer3_outputs(6767));
    layer4_outputs(6829) <= not((layer3_outputs(467)) or (layer3_outputs(7589)));
    layer4_outputs(6830) <= not((layer3_outputs(4118)) xor (layer3_outputs(3415)));
    layer4_outputs(6831) <= (layer3_outputs(3572)) xor (layer3_outputs(6322));
    layer4_outputs(6832) <= not((layer3_outputs(5394)) xor (layer3_outputs(1300)));
    layer4_outputs(6833) <= (layer3_outputs(399)) and not (layer3_outputs(5130));
    layer4_outputs(6834) <= not(layer3_outputs(4429));
    layer4_outputs(6835) <= not((layer3_outputs(5534)) or (layer3_outputs(3234)));
    layer4_outputs(6836) <= not((layer3_outputs(6100)) xor (layer3_outputs(4213)));
    layer4_outputs(6837) <= not(layer3_outputs(6984));
    layer4_outputs(6838) <= layer3_outputs(5265);
    layer4_outputs(6839) <= (layer3_outputs(7649)) xor (layer3_outputs(445));
    layer4_outputs(6840) <= not((layer3_outputs(324)) xor (layer3_outputs(775)));
    layer4_outputs(6841) <= (layer3_outputs(3527)) and (layer3_outputs(4470));
    layer4_outputs(6842) <= layer3_outputs(2940);
    layer4_outputs(6843) <= not(layer3_outputs(2010));
    layer4_outputs(6844) <= not((layer3_outputs(1719)) xor (layer3_outputs(1888)));
    layer4_outputs(6845) <= not(layer3_outputs(1350));
    layer4_outputs(6846) <= not((layer3_outputs(1341)) or (layer3_outputs(5147)));
    layer4_outputs(6847) <= layer3_outputs(1840);
    layer4_outputs(6848) <= (layer3_outputs(7647)) and not (layer3_outputs(7053));
    layer4_outputs(6849) <= not((layer3_outputs(3448)) xor (layer3_outputs(2738)));
    layer4_outputs(6850) <= not(layer3_outputs(477));
    layer4_outputs(6851) <= (layer3_outputs(1127)) or (layer3_outputs(5125));
    layer4_outputs(6852) <= not((layer3_outputs(2611)) or (layer3_outputs(5190)));
    layer4_outputs(6853) <= not(layer3_outputs(7006)) or (layer3_outputs(461));
    layer4_outputs(6854) <= layer3_outputs(3494);
    layer4_outputs(6855) <= layer3_outputs(6575);
    layer4_outputs(6856) <= layer3_outputs(6650);
    layer4_outputs(6857) <= layer3_outputs(4856);
    layer4_outputs(6858) <= not((layer3_outputs(784)) or (layer3_outputs(4362)));
    layer4_outputs(6859) <= layer3_outputs(6012);
    layer4_outputs(6860) <= not(layer3_outputs(2167)) or (layer3_outputs(5388));
    layer4_outputs(6861) <= layer3_outputs(3023);
    layer4_outputs(6862) <= not(layer3_outputs(487));
    layer4_outputs(6863) <= layer3_outputs(1277);
    layer4_outputs(6864) <= not((layer3_outputs(7584)) or (layer3_outputs(4742)));
    layer4_outputs(6865) <= not(layer3_outputs(1241));
    layer4_outputs(6866) <= not(layer3_outputs(6184));
    layer4_outputs(6867) <= layer3_outputs(2540);
    layer4_outputs(6868) <= not(layer3_outputs(3287));
    layer4_outputs(6869) <= (layer3_outputs(4486)) or (layer3_outputs(6544));
    layer4_outputs(6870) <= not((layer3_outputs(5672)) xor (layer3_outputs(1857)));
    layer4_outputs(6871) <= (layer3_outputs(6238)) and not (layer3_outputs(5969));
    layer4_outputs(6872) <= (layer3_outputs(5919)) and (layer3_outputs(849));
    layer4_outputs(6873) <= (layer3_outputs(118)) and not (layer3_outputs(6959));
    layer4_outputs(6874) <= not(layer3_outputs(238)) or (layer3_outputs(6079));
    layer4_outputs(6875) <= layer3_outputs(1228);
    layer4_outputs(6876) <= not((layer3_outputs(7299)) and (layer3_outputs(3194)));
    layer4_outputs(6877) <= layer3_outputs(39);
    layer4_outputs(6878) <= (layer3_outputs(6686)) or (layer3_outputs(1409));
    layer4_outputs(6879) <= not(layer3_outputs(5329));
    layer4_outputs(6880) <= '1';
    layer4_outputs(6881) <= layer3_outputs(686);
    layer4_outputs(6882) <= not(layer3_outputs(956));
    layer4_outputs(6883) <= (layer3_outputs(6123)) and not (layer3_outputs(5513));
    layer4_outputs(6884) <= (layer3_outputs(271)) and not (layer3_outputs(970));
    layer4_outputs(6885) <= not(layer3_outputs(6161)) or (layer3_outputs(6528));
    layer4_outputs(6886) <= layer3_outputs(2985);
    layer4_outputs(6887) <= layer3_outputs(2947);
    layer4_outputs(6888) <= layer3_outputs(2145);
    layer4_outputs(6889) <= (layer3_outputs(4821)) xor (layer3_outputs(398));
    layer4_outputs(6890) <= (layer3_outputs(2096)) and not (layer3_outputs(629));
    layer4_outputs(6891) <= (layer3_outputs(3046)) and not (layer3_outputs(5764));
    layer4_outputs(6892) <= layer3_outputs(3633);
    layer4_outputs(6893) <= not(layer3_outputs(4023));
    layer4_outputs(6894) <= (layer3_outputs(2607)) and (layer3_outputs(6989));
    layer4_outputs(6895) <= (layer3_outputs(2968)) and not (layer3_outputs(5608));
    layer4_outputs(6896) <= not(layer3_outputs(4450)) or (layer3_outputs(885));
    layer4_outputs(6897) <= layer3_outputs(1264);
    layer4_outputs(6898) <= not(layer3_outputs(5139));
    layer4_outputs(6899) <= layer3_outputs(4216);
    layer4_outputs(6900) <= (layer3_outputs(2915)) and not (layer3_outputs(4375));
    layer4_outputs(6901) <= layer3_outputs(7174);
    layer4_outputs(6902) <= not(layer3_outputs(3109)) or (layer3_outputs(5605));
    layer4_outputs(6903) <= not(layer3_outputs(5879));
    layer4_outputs(6904) <= not(layer3_outputs(5935)) or (layer3_outputs(3632));
    layer4_outputs(6905) <= not(layer3_outputs(1145));
    layer4_outputs(6906) <= not(layer3_outputs(782));
    layer4_outputs(6907) <= not(layer3_outputs(4718));
    layer4_outputs(6908) <= not((layer3_outputs(824)) and (layer3_outputs(6529)));
    layer4_outputs(6909) <= (layer3_outputs(1198)) or (layer3_outputs(4977));
    layer4_outputs(6910) <= (layer3_outputs(733)) and not (layer3_outputs(2470));
    layer4_outputs(6911) <= layer3_outputs(5205);
    layer4_outputs(6912) <= not(layer3_outputs(7154)) or (layer3_outputs(4217));
    layer4_outputs(6913) <= (layer3_outputs(938)) or (layer3_outputs(5366));
    layer4_outputs(6914) <= not((layer3_outputs(1017)) xor (layer3_outputs(7056)));
    layer4_outputs(6915) <= not(layer3_outputs(2980));
    layer4_outputs(6916) <= not(layer3_outputs(1317)) or (layer3_outputs(7267));
    layer4_outputs(6917) <= not(layer3_outputs(4948));
    layer4_outputs(6918) <= (layer3_outputs(1824)) and not (layer3_outputs(4108));
    layer4_outputs(6919) <= layer3_outputs(609);
    layer4_outputs(6920) <= (layer3_outputs(2332)) xor (layer3_outputs(2715));
    layer4_outputs(6921) <= not(layer3_outputs(2576)) or (layer3_outputs(3819));
    layer4_outputs(6922) <= not(layer3_outputs(5280));
    layer4_outputs(6923) <= (layer3_outputs(1048)) and not (layer3_outputs(5001));
    layer4_outputs(6924) <= layer3_outputs(3184);
    layer4_outputs(6925) <= (layer3_outputs(4241)) and (layer3_outputs(5012));
    layer4_outputs(6926) <= (layer3_outputs(2325)) and (layer3_outputs(2057));
    layer4_outputs(6927) <= (layer3_outputs(1218)) and not (layer3_outputs(316));
    layer4_outputs(6928) <= not(layer3_outputs(6484));
    layer4_outputs(6929) <= not(layer3_outputs(4122));
    layer4_outputs(6930) <= not(layer3_outputs(4541));
    layer4_outputs(6931) <= not(layer3_outputs(4138)) or (layer3_outputs(6499));
    layer4_outputs(6932) <= not(layer3_outputs(243));
    layer4_outputs(6933) <= layer3_outputs(749);
    layer4_outputs(6934) <= not(layer3_outputs(948));
    layer4_outputs(6935) <= not(layer3_outputs(1761));
    layer4_outputs(6936) <= layer3_outputs(71);
    layer4_outputs(6937) <= (layer3_outputs(291)) and not (layer3_outputs(3005));
    layer4_outputs(6938) <= layer3_outputs(1725);
    layer4_outputs(6939) <= (layer3_outputs(5758)) and (layer3_outputs(7520));
    layer4_outputs(6940) <= not(layer3_outputs(1334));
    layer4_outputs(6941) <= layer3_outputs(3469);
    layer4_outputs(6942) <= not((layer3_outputs(2662)) and (layer3_outputs(7232)));
    layer4_outputs(6943) <= layer3_outputs(6593);
    layer4_outputs(6944) <= (layer3_outputs(4617)) or (layer3_outputs(4046));
    layer4_outputs(6945) <= not(layer3_outputs(225));
    layer4_outputs(6946) <= (layer3_outputs(7532)) and not (layer3_outputs(2209));
    layer4_outputs(6947) <= layer3_outputs(3019);
    layer4_outputs(6948) <= not((layer3_outputs(909)) or (layer3_outputs(6479)));
    layer4_outputs(6949) <= (layer3_outputs(7462)) or (layer3_outputs(7099));
    layer4_outputs(6950) <= (layer3_outputs(908)) or (layer3_outputs(1414));
    layer4_outputs(6951) <= (layer3_outputs(2486)) xor (layer3_outputs(3995));
    layer4_outputs(6952) <= not(layer3_outputs(5153)) or (layer3_outputs(2206));
    layer4_outputs(6953) <= layer3_outputs(1046);
    layer4_outputs(6954) <= not(layer3_outputs(1508));
    layer4_outputs(6955) <= layer3_outputs(5864);
    layer4_outputs(6956) <= not(layer3_outputs(1205)) or (layer3_outputs(649));
    layer4_outputs(6957) <= layer3_outputs(1259);
    layer4_outputs(6958) <= layer3_outputs(4646);
    layer4_outputs(6959) <= layer3_outputs(5518);
    layer4_outputs(6960) <= layer3_outputs(368);
    layer4_outputs(6961) <= (layer3_outputs(6916)) xor (layer3_outputs(7459));
    layer4_outputs(6962) <= layer3_outputs(4591);
    layer4_outputs(6963) <= not((layer3_outputs(633)) and (layer3_outputs(700)));
    layer4_outputs(6964) <= layer3_outputs(7565);
    layer4_outputs(6965) <= layer3_outputs(1689);
    layer4_outputs(6966) <= not(layer3_outputs(7013));
    layer4_outputs(6967) <= not((layer3_outputs(6085)) xor (layer3_outputs(1055)));
    layer4_outputs(6968) <= layer3_outputs(5826);
    layer4_outputs(6969) <= not(layer3_outputs(1519));
    layer4_outputs(6970) <= not(layer3_outputs(4895)) or (layer3_outputs(1674));
    layer4_outputs(6971) <= not((layer3_outputs(1675)) xor (layer3_outputs(2370)));
    layer4_outputs(6972) <= not((layer3_outputs(5641)) xor (layer3_outputs(5880)));
    layer4_outputs(6973) <= layer3_outputs(4638);
    layer4_outputs(6974) <= not(layer3_outputs(4313));
    layer4_outputs(6975) <= not((layer3_outputs(6025)) and (layer3_outputs(6314)));
    layer4_outputs(6976) <= not((layer3_outputs(2393)) and (layer3_outputs(842)));
    layer4_outputs(6977) <= not(layer3_outputs(1413)) or (layer3_outputs(3030));
    layer4_outputs(6978) <= not((layer3_outputs(969)) and (layer3_outputs(6806)));
    layer4_outputs(6979) <= layer3_outputs(7441);
    layer4_outputs(6980) <= not((layer3_outputs(6361)) xor (layer3_outputs(7599)));
    layer4_outputs(6981) <= not((layer3_outputs(1395)) or (layer3_outputs(938)));
    layer4_outputs(6982) <= layer3_outputs(7255);
    layer4_outputs(6983) <= layer3_outputs(1378);
    layer4_outputs(6984) <= not(layer3_outputs(6734));
    layer4_outputs(6985) <= layer3_outputs(3213);
    layer4_outputs(6986) <= not(layer3_outputs(2300)) or (layer3_outputs(443));
    layer4_outputs(6987) <= (layer3_outputs(3249)) xor (layer3_outputs(5362));
    layer4_outputs(6988) <= layer3_outputs(5883);
    layer4_outputs(6989) <= layer3_outputs(2517);
    layer4_outputs(6990) <= not((layer3_outputs(6397)) or (layer3_outputs(2132)));
    layer4_outputs(6991) <= not(layer3_outputs(6003));
    layer4_outputs(6992) <= not((layer3_outputs(1163)) and (layer3_outputs(3840)));
    layer4_outputs(6993) <= (layer3_outputs(598)) or (layer3_outputs(3813));
    layer4_outputs(6994) <= (layer3_outputs(925)) and not (layer3_outputs(1476));
    layer4_outputs(6995) <= (layer3_outputs(2367)) or (layer3_outputs(4258));
    layer4_outputs(6996) <= layer3_outputs(5905);
    layer4_outputs(6997) <= not(layer3_outputs(3865));
    layer4_outputs(6998) <= not(layer3_outputs(282));
    layer4_outputs(6999) <= (layer3_outputs(5292)) and not (layer3_outputs(5563));
    layer4_outputs(7000) <= not(layer3_outputs(2895));
    layer4_outputs(7001) <= (layer3_outputs(6711)) or (layer3_outputs(7135));
    layer4_outputs(7002) <= (layer3_outputs(2095)) or (layer3_outputs(1785));
    layer4_outputs(7003) <= not((layer3_outputs(5505)) or (layer3_outputs(3184)));
    layer4_outputs(7004) <= layer3_outputs(5912);
    layer4_outputs(7005) <= (layer3_outputs(5180)) or (layer3_outputs(5601));
    layer4_outputs(7006) <= not(layer3_outputs(4837));
    layer4_outputs(7007) <= not(layer3_outputs(1508));
    layer4_outputs(7008) <= layer3_outputs(3379);
    layer4_outputs(7009) <= not(layer3_outputs(4711));
    layer4_outputs(7010) <= not(layer3_outputs(7528));
    layer4_outputs(7011) <= not(layer3_outputs(389)) or (layer3_outputs(127));
    layer4_outputs(7012) <= not((layer3_outputs(4869)) or (layer3_outputs(918)));
    layer4_outputs(7013) <= not((layer3_outputs(7041)) xor (layer3_outputs(2825)));
    layer4_outputs(7014) <= (layer3_outputs(2494)) and (layer3_outputs(3270));
    layer4_outputs(7015) <= not(layer3_outputs(3396)) or (layer3_outputs(5026));
    layer4_outputs(7016) <= (layer3_outputs(7351)) or (layer3_outputs(1766));
    layer4_outputs(7017) <= '0';
    layer4_outputs(7018) <= not((layer3_outputs(4855)) or (layer3_outputs(4866)));
    layer4_outputs(7019) <= not(layer3_outputs(6294)) or (layer3_outputs(5424));
    layer4_outputs(7020) <= (layer3_outputs(5420)) and not (layer3_outputs(3009));
    layer4_outputs(7021) <= not(layer3_outputs(6845));
    layer4_outputs(7022) <= not((layer3_outputs(3057)) xor (layer3_outputs(572)));
    layer4_outputs(7023) <= not(layer3_outputs(2248));
    layer4_outputs(7024) <= layer3_outputs(4764);
    layer4_outputs(7025) <= layer3_outputs(4066);
    layer4_outputs(7026) <= not(layer3_outputs(7381));
    layer4_outputs(7027) <= (layer3_outputs(7144)) xor (layer3_outputs(4177));
    layer4_outputs(7028) <= layer3_outputs(5563);
    layer4_outputs(7029) <= layer3_outputs(6009);
    layer4_outputs(7030) <= (layer3_outputs(6689)) xor (layer3_outputs(2146));
    layer4_outputs(7031) <= not((layer3_outputs(357)) or (layer3_outputs(2839)));
    layer4_outputs(7032) <= (layer3_outputs(1308)) and not (layer3_outputs(2129));
    layer4_outputs(7033) <= layer3_outputs(1690);
    layer4_outputs(7034) <= not(layer3_outputs(1901)) or (layer3_outputs(7169));
    layer4_outputs(7035) <= layer3_outputs(6396);
    layer4_outputs(7036) <= (layer3_outputs(3773)) and not (layer3_outputs(1804));
    layer4_outputs(7037) <= (layer3_outputs(5099)) and not (layer3_outputs(6289));
    layer4_outputs(7038) <= (layer3_outputs(4197)) xor (layer3_outputs(3219));
    layer4_outputs(7039) <= not(layer3_outputs(3533));
    layer4_outputs(7040) <= (layer3_outputs(2774)) and (layer3_outputs(7174));
    layer4_outputs(7041) <= not((layer3_outputs(4128)) xor (layer3_outputs(5550)));
    layer4_outputs(7042) <= layer3_outputs(4396);
    layer4_outputs(7043) <= not((layer3_outputs(131)) and (layer3_outputs(7403)));
    layer4_outputs(7044) <= layer3_outputs(6959);
    layer4_outputs(7045) <= layer3_outputs(6635);
    layer4_outputs(7046) <= not(layer3_outputs(5754)) or (layer3_outputs(6236));
    layer4_outputs(7047) <= layer3_outputs(4585);
    layer4_outputs(7048) <= (layer3_outputs(5324)) and (layer3_outputs(5665));
    layer4_outputs(7049) <= layer3_outputs(4138);
    layer4_outputs(7050) <= not(layer3_outputs(2659));
    layer4_outputs(7051) <= not(layer3_outputs(6104));
    layer4_outputs(7052) <= not(layer3_outputs(291)) or (layer3_outputs(3135));
    layer4_outputs(7053) <= not(layer3_outputs(7482));
    layer4_outputs(7054) <= not(layer3_outputs(6363)) or (layer3_outputs(533));
    layer4_outputs(7055) <= not(layer3_outputs(5677));
    layer4_outputs(7056) <= (layer3_outputs(6943)) and not (layer3_outputs(1239));
    layer4_outputs(7057) <= not(layer3_outputs(1513)) or (layer3_outputs(5588));
    layer4_outputs(7058) <= layer3_outputs(5958);
    layer4_outputs(7059) <= not((layer3_outputs(7673)) or (layer3_outputs(4727)));
    layer4_outputs(7060) <= layer3_outputs(5249);
    layer4_outputs(7061) <= layer3_outputs(7563);
    layer4_outputs(7062) <= layer3_outputs(4949);
    layer4_outputs(7063) <= not(layer3_outputs(4518)) or (layer3_outputs(5093));
    layer4_outputs(7064) <= layer3_outputs(3274);
    layer4_outputs(7065) <= (layer3_outputs(5944)) and not (layer3_outputs(1838));
    layer4_outputs(7066) <= (layer3_outputs(1182)) and not (layer3_outputs(3181));
    layer4_outputs(7067) <= not((layer3_outputs(4007)) or (layer3_outputs(2347)));
    layer4_outputs(7068) <= not((layer3_outputs(1026)) xor (layer3_outputs(6717)));
    layer4_outputs(7069) <= layer3_outputs(1276);
    layer4_outputs(7070) <= layer3_outputs(3319);
    layer4_outputs(7071) <= layer3_outputs(4182);
    layer4_outputs(7072) <= not(layer3_outputs(1837));
    layer4_outputs(7073) <= (layer3_outputs(5820)) and (layer3_outputs(7648));
    layer4_outputs(7074) <= '1';
    layer4_outputs(7075) <= (layer3_outputs(371)) or (layer3_outputs(7287));
    layer4_outputs(7076) <= not(layer3_outputs(7476));
    layer4_outputs(7077) <= not(layer3_outputs(437)) or (layer3_outputs(1645));
    layer4_outputs(7078) <= not((layer3_outputs(1240)) xor (layer3_outputs(7322)));
    layer4_outputs(7079) <= not((layer3_outputs(6167)) xor (layer3_outputs(5889)));
    layer4_outputs(7080) <= (layer3_outputs(4776)) and not (layer3_outputs(7494));
    layer4_outputs(7081) <= not((layer3_outputs(6659)) and (layer3_outputs(4254)));
    layer4_outputs(7082) <= (layer3_outputs(7547)) or (layer3_outputs(2072));
    layer4_outputs(7083) <= (layer3_outputs(2901)) and not (layer3_outputs(951));
    layer4_outputs(7084) <= layer3_outputs(5699);
    layer4_outputs(7085) <= (layer3_outputs(5356)) and not (layer3_outputs(2902));
    layer4_outputs(7086) <= (layer3_outputs(3722)) and (layer3_outputs(7639));
    layer4_outputs(7087) <= not((layer3_outputs(2290)) xor (layer3_outputs(7238)));
    layer4_outputs(7088) <= not(layer3_outputs(1914));
    layer4_outputs(7089) <= (layer3_outputs(2765)) and not (layer3_outputs(42));
    layer4_outputs(7090) <= not(layer3_outputs(3674)) or (layer3_outputs(2507));
    layer4_outputs(7091) <= not((layer3_outputs(5596)) xor (layer3_outputs(1409)));
    layer4_outputs(7092) <= (layer3_outputs(1925)) xor (layer3_outputs(5104));
    layer4_outputs(7093) <= layer3_outputs(1389);
    layer4_outputs(7094) <= (layer3_outputs(721)) and (layer3_outputs(3283));
    layer4_outputs(7095) <= not(layer3_outputs(6254));
    layer4_outputs(7096) <= not(layer3_outputs(771));
    layer4_outputs(7097) <= not(layer3_outputs(1868));
    layer4_outputs(7098) <= layer3_outputs(5084);
    layer4_outputs(7099) <= (layer3_outputs(3926)) or (layer3_outputs(5167));
    layer4_outputs(7100) <= not((layer3_outputs(6166)) xor (layer3_outputs(570)));
    layer4_outputs(7101) <= not(layer3_outputs(6967)) or (layer3_outputs(6670));
    layer4_outputs(7102) <= (layer3_outputs(5514)) and not (layer3_outputs(1257));
    layer4_outputs(7103) <= layer3_outputs(3045);
    layer4_outputs(7104) <= not(layer3_outputs(2053)) or (layer3_outputs(7133));
    layer4_outputs(7105) <= (layer3_outputs(1835)) or (layer3_outputs(2779));
    layer4_outputs(7106) <= not(layer3_outputs(7066)) or (layer3_outputs(4381));
    layer4_outputs(7107) <= (layer3_outputs(3399)) and not (layer3_outputs(267));
    layer4_outputs(7108) <= (layer3_outputs(5710)) and not (layer3_outputs(6841));
    layer4_outputs(7109) <= (layer3_outputs(3295)) and not (layer3_outputs(6351));
    layer4_outputs(7110) <= (layer3_outputs(355)) and (layer3_outputs(1420));
    layer4_outputs(7111) <= not((layer3_outputs(2812)) xor (layer3_outputs(6559)));
    layer4_outputs(7112) <= layer3_outputs(5237);
    layer4_outputs(7113) <= not(layer3_outputs(2757)) or (layer3_outputs(5354));
    layer4_outputs(7114) <= (layer3_outputs(5775)) or (layer3_outputs(125));
    layer4_outputs(7115) <= (layer3_outputs(3870)) and not (layer3_outputs(167));
    layer4_outputs(7116) <= layer3_outputs(3456);
    layer4_outputs(7117) <= not((layer3_outputs(2428)) xor (layer3_outputs(2281)));
    layer4_outputs(7118) <= (layer3_outputs(3615)) and not (layer3_outputs(3228));
    layer4_outputs(7119) <= not(layer3_outputs(6335));
    layer4_outputs(7120) <= layer3_outputs(3924);
    layer4_outputs(7121) <= (layer3_outputs(211)) xor (layer3_outputs(2251));
    layer4_outputs(7122) <= not(layer3_outputs(2565));
    layer4_outputs(7123) <= not(layer3_outputs(4721));
    layer4_outputs(7124) <= layer3_outputs(5056);
    layer4_outputs(7125) <= layer3_outputs(7038);
    layer4_outputs(7126) <= not((layer3_outputs(1421)) xor (layer3_outputs(6136)));
    layer4_outputs(7127) <= layer3_outputs(753);
    layer4_outputs(7128) <= not(layer3_outputs(5795));
    layer4_outputs(7129) <= not(layer3_outputs(851));
    layer4_outputs(7130) <= (layer3_outputs(5158)) or (layer3_outputs(710));
    layer4_outputs(7131) <= layer3_outputs(7348);
    layer4_outputs(7132) <= (layer3_outputs(6122)) and not (layer3_outputs(6866));
    layer4_outputs(7133) <= (layer3_outputs(3371)) or (layer3_outputs(6378));
    layer4_outputs(7134) <= layer3_outputs(4517);
    layer4_outputs(7135) <= layer3_outputs(2718);
    layer4_outputs(7136) <= (layer3_outputs(6801)) and not (layer3_outputs(1430));
    layer4_outputs(7137) <= not(layer3_outputs(4922));
    layer4_outputs(7138) <= layer3_outputs(3510);
    layer4_outputs(7139) <= (layer3_outputs(518)) xor (layer3_outputs(1001));
    layer4_outputs(7140) <= not(layer3_outputs(5570));
    layer4_outputs(7141) <= layer3_outputs(5024);
    layer4_outputs(7142) <= layer3_outputs(3522);
    layer4_outputs(7143) <= layer3_outputs(2011);
    layer4_outputs(7144) <= not(layer3_outputs(3865));
    layer4_outputs(7145) <= layer3_outputs(1538);
    layer4_outputs(7146) <= not(layer3_outputs(3098));
    layer4_outputs(7147) <= not(layer3_outputs(4699)) or (layer3_outputs(4530));
    layer4_outputs(7148) <= layer3_outputs(5004);
    layer4_outputs(7149) <= not((layer3_outputs(5867)) xor (layer3_outputs(6230)));
    layer4_outputs(7150) <= not(layer3_outputs(952)) or (layer3_outputs(897));
    layer4_outputs(7151) <= not((layer3_outputs(7353)) and (layer3_outputs(1226)));
    layer4_outputs(7152) <= not(layer3_outputs(4893));
    layer4_outputs(7153) <= layer3_outputs(1427);
    layer4_outputs(7154) <= (layer3_outputs(1312)) xor (layer3_outputs(2243));
    layer4_outputs(7155) <= not((layer3_outputs(2927)) and (layer3_outputs(6908)));
    layer4_outputs(7156) <= (layer3_outputs(3629)) or (layer3_outputs(7386));
    layer4_outputs(7157) <= (layer3_outputs(5051)) xor (layer3_outputs(1590));
    layer4_outputs(7158) <= not(layer3_outputs(1342));
    layer4_outputs(7159) <= not(layer3_outputs(7225));
    layer4_outputs(7160) <= not(layer3_outputs(5800));
    layer4_outputs(7161) <= layer3_outputs(3938);
    layer4_outputs(7162) <= not(layer3_outputs(3805));
    layer4_outputs(7163) <= layer3_outputs(6099);
    layer4_outputs(7164) <= not(layer3_outputs(4483));
    layer4_outputs(7165) <= not((layer3_outputs(2531)) xor (layer3_outputs(6759)));
    layer4_outputs(7166) <= (layer3_outputs(2706)) xor (layer3_outputs(4678));
    layer4_outputs(7167) <= layer3_outputs(767);
    layer4_outputs(7168) <= not((layer3_outputs(2526)) xor (layer3_outputs(4176)));
    layer4_outputs(7169) <= (layer3_outputs(5735)) xor (layer3_outputs(1739));
    layer4_outputs(7170) <= layer3_outputs(4326);
    layer4_outputs(7171) <= layer3_outputs(1215);
    layer4_outputs(7172) <= '0';
    layer4_outputs(7173) <= (layer3_outputs(7212)) and not (layer3_outputs(3344));
    layer4_outputs(7174) <= not((layer3_outputs(1488)) or (layer3_outputs(1630)));
    layer4_outputs(7175) <= not(layer3_outputs(7640));
    layer4_outputs(7176) <= layer3_outputs(770);
    layer4_outputs(7177) <= not((layer3_outputs(6373)) xor (layer3_outputs(1597)));
    layer4_outputs(7178) <= (layer3_outputs(422)) xor (layer3_outputs(813));
    layer4_outputs(7179) <= (layer3_outputs(3244)) xor (layer3_outputs(1846));
    layer4_outputs(7180) <= not(layer3_outputs(5453));
    layer4_outputs(7181) <= layer3_outputs(4680);
    layer4_outputs(7182) <= not(layer3_outputs(7068));
    layer4_outputs(7183) <= (layer3_outputs(4790)) xor (layer3_outputs(4565));
    layer4_outputs(7184) <= layer3_outputs(4319);
    layer4_outputs(7185) <= not(layer3_outputs(993)) or (layer3_outputs(6160));
    layer4_outputs(7186) <= not(layer3_outputs(1993));
    layer4_outputs(7187) <= not((layer3_outputs(116)) or (layer3_outputs(3097)));
    layer4_outputs(7188) <= not(layer3_outputs(2059));
    layer4_outputs(7189) <= not(layer3_outputs(3011));
    layer4_outputs(7190) <= not(layer3_outputs(177)) or (layer3_outputs(1634));
    layer4_outputs(7191) <= not(layer3_outputs(762));
    layer4_outputs(7192) <= not(layer3_outputs(2816)) or (layer3_outputs(1363));
    layer4_outputs(7193) <= (layer3_outputs(5390)) xor (layer3_outputs(1412));
    layer4_outputs(7194) <= not(layer3_outputs(5226));
    layer4_outputs(7195) <= (layer3_outputs(5162)) and not (layer3_outputs(1950));
    layer4_outputs(7196) <= not((layer3_outputs(2258)) xor (layer3_outputs(1137)));
    layer4_outputs(7197) <= not(layer3_outputs(6713));
    layer4_outputs(7198) <= layer3_outputs(7308);
    layer4_outputs(7199) <= not(layer3_outputs(1678));
    layer4_outputs(7200) <= (layer3_outputs(2268)) xor (layer3_outputs(6816));
    layer4_outputs(7201) <= not((layer3_outputs(438)) or (layer3_outputs(6707)));
    layer4_outputs(7202) <= not((layer3_outputs(7052)) or (layer3_outputs(5811)));
    layer4_outputs(7203) <= layer3_outputs(7092);
    layer4_outputs(7204) <= layer3_outputs(4802);
    layer4_outputs(7205) <= not(layer3_outputs(834));
    layer4_outputs(7206) <= not(layer3_outputs(5180)) or (layer3_outputs(199));
    layer4_outputs(7207) <= not(layer3_outputs(913));
    layer4_outputs(7208) <= (layer3_outputs(1606)) or (layer3_outputs(7168));
    layer4_outputs(7209) <= not(layer3_outputs(5719));
    layer4_outputs(7210) <= not((layer3_outputs(2996)) xor (layer3_outputs(5487)));
    layer4_outputs(7211) <= not((layer3_outputs(6505)) or (layer3_outputs(401)));
    layer4_outputs(7212) <= not(layer3_outputs(6140));
    layer4_outputs(7213) <= (layer3_outputs(1514)) and not (layer3_outputs(506));
    layer4_outputs(7214) <= (layer3_outputs(7555)) and not (layer3_outputs(2811));
    layer4_outputs(7215) <= (layer3_outputs(7009)) and not (layer3_outputs(7285));
    layer4_outputs(7216) <= not((layer3_outputs(1203)) and (layer3_outputs(6334)));
    layer4_outputs(7217) <= (layer3_outputs(1210)) and not (layer3_outputs(3205));
    layer4_outputs(7218) <= (layer3_outputs(60)) or (layer3_outputs(5363));
    layer4_outputs(7219) <= not(layer3_outputs(4402));
    layer4_outputs(7220) <= not(layer3_outputs(5785));
    layer4_outputs(7221) <= (layer3_outputs(3853)) or (layer3_outputs(2108));
    layer4_outputs(7222) <= not((layer3_outputs(220)) and (layer3_outputs(6188)));
    layer4_outputs(7223) <= '0';
    layer4_outputs(7224) <= not((layer3_outputs(4838)) or (layer3_outputs(3629)));
    layer4_outputs(7225) <= (layer3_outputs(6777)) and not (layer3_outputs(5060));
    layer4_outputs(7226) <= not(layer3_outputs(4295)) or (layer3_outputs(160));
    layer4_outputs(7227) <= (layer3_outputs(6059)) and not (layer3_outputs(3069));
    layer4_outputs(7228) <= layer3_outputs(2127);
    layer4_outputs(7229) <= not(layer3_outputs(791)) or (layer3_outputs(1271));
    layer4_outputs(7230) <= not((layer3_outputs(3080)) and (layer3_outputs(1383)));
    layer4_outputs(7231) <= layer3_outputs(5464);
    layer4_outputs(7232) <= (layer3_outputs(6752)) or (layer3_outputs(4961));
    layer4_outputs(7233) <= not(layer3_outputs(5441));
    layer4_outputs(7234) <= (layer3_outputs(7191)) xor (layer3_outputs(1935));
    layer4_outputs(7235) <= layer3_outputs(6576);
    layer4_outputs(7236) <= not(layer3_outputs(7224)) or (layer3_outputs(6817));
    layer4_outputs(7237) <= layer3_outputs(5152);
    layer4_outputs(7238) <= layer3_outputs(780);
    layer4_outputs(7239) <= not((layer3_outputs(812)) or (layer3_outputs(1499)));
    layer4_outputs(7240) <= layer3_outputs(2994);
    layer4_outputs(7241) <= (layer3_outputs(4334)) or (layer3_outputs(6523));
    layer4_outputs(7242) <= not((layer3_outputs(6807)) or (layer3_outputs(5161)));
    layer4_outputs(7243) <= not(layer3_outputs(4240)) or (layer3_outputs(113));
    layer4_outputs(7244) <= not(layer3_outputs(2390));
    layer4_outputs(7245) <= '1';
    layer4_outputs(7246) <= not((layer3_outputs(1822)) and (layer3_outputs(3432)));
    layer4_outputs(7247) <= not((layer3_outputs(5808)) and (layer3_outputs(7057)));
    layer4_outputs(7248) <= not((layer3_outputs(1302)) xor (layer3_outputs(2326)));
    layer4_outputs(7249) <= not((layer3_outputs(3967)) or (layer3_outputs(3736)));
    layer4_outputs(7250) <= not((layer3_outputs(127)) or (layer3_outputs(7185)));
    layer4_outputs(7251) <= (layer3_outputs(5506)) and not (layer3_outputs(2032));
    layer4_outputs(7252) <= not(layer3_outputs(4038)) or (layer3_outputs(7355));
    layer4_outputs(7253) <= not((layer3_outputs(3914)) xor (layer3_outputs(573)));
    layer4_outputs(7254) <= not(layer3_outputs(1967));
    layer4_outputs(7255) <= not((layer3_outputs(4021)) or (layer3_outputs(1186)));
    layer4_outputs(7256) <= not(layer3_outputs(931));
    layer4_outputs(7257) <= not(layer3_outputs(1005)) or (layer3_outputs(6674));
    layer4_outputs(7258) <= (layer3_outputs(4788)) xor (layer3_outputs(4428));
    layer4_outputs(7259) <= not(layer3_outputs(1570));
    layer4_outputs(7260) <= not(layer3_outputs(3506));
    layer4_outputs(7261) <= not(layer3_outputs(2002));
    layer4_outputs(7262) <= layer3_outputs(62);
    layer4_outputs(7263) <= (layer3_outputs(7195)) and not (layer3_outputs(6832));
    layer4_outputs(7264) <= not(layer3_outputs(2398)) or (layer3_outputs(2151));
    layer4_outputs(7265) <= (layer3_outputs(5743)) or (layer3_outputs(423));
    layer4_outputs(7266) <= (layer3_outputs(4186)) xor (layer3_outputs(7212));
    layer4_outputs(7267) <= (layer3_outputs(2440)) and (layer3_outputs(2500));
    layer4_outputs(7268) <= (layer3_outputs(6991)) and not (layer3_outputs(7498));
    layer4_outputs(7269) <= (layer3_outputs(5404)) xor (layer3_outputs(922));
    layer4_outputs(7270) <= (layer3_outputs(4417)) or (layer3_outputs(78));
    layer4_outputs(7271) <= not((layer3_outputs(5090)) and (layer3_outputs(4645)));
    layer4_outputs(7272) <= not(layer3_outputs(3491));
    layer4_outputs(7273) <= layer3_outputs(7064);
    layer4_outputs(7274) <= not(layer3_outputs(1639));
    layer4_outputs(7275) <= (layer3_outputs(5967)) and not (layer3_outputs(2291));
    layer4_outputs(7276) <= not(layer3_outputs(2656));
    layer4_outputs(7277) <= not((layer3_outputs(6797)) and (layer3_outputs(247)));
    layer4_outputs(7278) <= (layer3_outputs(5048)) or (layer3_outputs(5481));
    layer4_outputs(7279) <= not(layer3_outputs(253));
    layer4_outputs(7280) <= not(layer3_outputs(265));
    layer4_outputs(7281) <= layer3_outputs(5871);
    layer4_outputs(7282) <= layer3_outputs(2598);
    layer4_outputs(7283) <= not((layer3_outputs(275)) and (layer3_outputs(3237)));
    layer4_outputs(7284) <= not(layer3_outputs(6489)) or (layer3_outputs(5177));
    layer4_outputs(7285) <= layer3_outputs(1030);
    layer4_outputs(7286) <= not((layer3_outputs(4816)) or (layer3_outputs(5548)));
    layer4_outputs(7287) <= not(layer3_outputs(1452));
    layer4_outputs(7288) <= not(layer3_outputs(5071));
    layer4_outputs(7289) <= not(layer3_outputs(5705)) or (layer3_outputs(1908));
    layer4_outputs(7290) <= not(layer3_outputs(3669));
    layer4_outputs(7291) <= (layer3_outputs(4000)) xor (layer3_outputs(4996));
    layer4_outputs(7292) <= not(layer3_outputs(7273)) or (layer3_outputs(3875));
    layer4_outputs(7293) <= (layer3_outputs(5091)) and not (layer3_outputs(4002));
    layer4_outputs(7294) <= not(layer3_outputs(5447)) or (layer3_outputs(1733));
    layer4_outputs(7295) <= '0';
    layer4_outputs(7296) <= not(layer3_outputs(2245));
    layer4_outputs(7297) <= not((layer3_outputs(3647)) or (layer3_outputs(4613)));
    layer4_outputs(7298) <= layer3_outputs(3136);
    layer4_outputs(7299) <= not(layer3_outputs(636)) or (layer3_outputs(4109));
    layer4_outputs(7300) <= not((layer3_outputs(4715)) and (layer3_outputs(1610)));
    layer4_outputs(7301) <= (layer3_outputs(4435)) or (layer3_outputs(6761));
    layer4_outputs(7302) <= (layer3_outputs(4259)) and (layer3_outputs(7299));
    layer4_outputs(7303) <= not(layer3_outputs(3593)) or (layer3_outputs(5700));
    layer4_outputs(7304) <= layer3_outputs(5666);
    layer4_outputs(7305) <= (layer3_outputs(2315)) and (layer3_outputs(3113));
    layer4_outputs(7306) <= (layer3_outputs(4535)) or (layer3_outputs(6214));
    layer4_outputs(7307) <= layer3_outputs(1940);
    layer4_outputs(7308) <= not(layer3_outputs(3487));
    layer4_outputs(7309) <= layer3_outputs(6219);
    layer4_outputs(7310) <= layer3_outputs(3104);
    layer4_outputs(7311) <= not((layer3_outputs(1374)) or (layer3_outputs(618)));
    layer4_outputs(7312) <= (layer3_outputs(4004)) and (layer3_outputs(1432));
    layer4_outputs(7313) <= layer3_outputs(3490);
    layer4_outputs(7314) <= (layer3_outputs(6552)) and not (layer3_outputs(1815));
    layer4_outputs(7315) <= not(layer3_outputs(6369));
    layer4_outputs(7316) <= layer3_outputs(5274);
    layer4_outputs(7317) <= (layer3_outputs(943)) xor (layer3_outputs(6441));
    layer4_outputs(7318) <= layer3_outputs(4291);
    layer4_outputs(7319) <= (layer3_outputs(907)) or (layer3_outputs(4169));
    layer4_outputs(7320) <= not(layer3_outputs(1139));
    layer4_outputs(7321) <= not(layer3_outputs(4659)) or (layer3_outputs(622));
    layer4_outputs(7322) <= not((layer3_outputs(2879)) and (layer3_outputs(4600)));
    layer4_outputs(7323) <= (layer3_outputs(6279)) and not (layer3_outputs(2456));
    layer4_outputs(7324) <= not(layer3_outputs(6809));
    layer4_outputs(7325) <= layer3_outputs(7049);
    layer4_outputs(7326) <= not((layer3_outputs(2423)) xor (layer3_outputs(701)));
    layer4_outputs(7327) <= not(layer3_outputs(1035));
    layer4_outputs(7328) <= (layer3_outputs(374)) xor (layer3_outputs(2450));
    layer4_outputs(7329) <= not((layer3_outputs(4585)) and (layer3_outputs(7375)));
    layer4_outputs(7330) <= not((layer3_outputs(7136)) xor (layer3_outputs(810)));
    layer4_outputs(7331) <= layer3_outputs(1528);
    layer4_outputs(7332) <= layer3_outputs(5681);
    layer4_outputs(7333) <= (layer3_outputs(2417)) and not (layer3_outputs(2434));
    layer4_outputs(7334) <= not(layer3_outputs(5289));
    layer4_outputs(7335) <= not(layer3_outputs(5939)) or (layer3_outputs(6107));
    layer4_outputs(7336) <= layer3_outputs(3463);
    layer4_outputs(7337) <= layer3_outputs(6920);
    layer4_outputs(7338) <= not(layer3_outputs(7465));
    layer4_outputs(7339) <= layer3_outputs(4616);
    layer4_outputs(7340) <= not((layer3_outputs(5929)) xor (layer3_outputs(7661)));
    layer4_outputs(7341) <= layer3_outputs(2083);
    layer4_outputs(7342) <= not(layer3_outputs(3400)) or (layer3_outputs(3671));
    layer4_outputs(7343) <= not((layer3_outputs(5974)) xor (layer3_outputs(7391)));
    layer4_outputs(7344) <= not((layer3_outputs(2576)) or (layer3_outputs(1848)));
    layer4_outputs(7345) <= layer3_outputs(6175);
    layer4_outputs(7346) <= (layer3_outputs(2872)) or (layer3_outputs(6966));
    layer4_outputs(7347) <= (layer3_outputs(7440)) and (layer3_outputs(7399));
    layer4_outputs(7348) <= layer3_outputs(2043);
    layer4_outputs(7349) <= not(layer3_outputs(4576));
    layer4_outputs(7350) <= (layer3_outputs(4083)) and (layer3_outputs(920));
    layer4_outputs(7351) <= not(layer3_outputs(4765));
    layer4_outputs(7352) <= not(layer3_outputs(6283)) or (layer3_outputs(1510));
    layer4_outputs(7353) <= not((layer3_outputs(3196)) or (layer3_outputs(777)));
    layer4_outputs(7354) <= (layer3_outputs(6321)) and (layer3_outputs(3732));
    layer4_outputs(7355) <= layer3_outputs(381);
    layer4_outputs(7356) <= not(layer3_outputs(6870));
    layer4_outputs(7357) <= not(layer3_outputs(5667));
    layer4_outputs(7358) <= not(layer3_outputs(3288)) or (layer3_outputs(165));
    layer4_outputs(7359) <= not(layer3_outputs(6440));
    layer4_outputs(7360) <= (layer3_outputs(2156)) or (layer3_outputs(5855));
    layer4_outputs(7361) <= layer3_outputs(3905);
    layer4_outputs(7362) <= layer3_outputs(3843);
    layer4_outputs(7363) <= layer3_outputs(2838);
    layer4_outputs(7364) <= not(layer3_outputs(7053));
    layer4_outputs(7365) <= layer3_outputs(1772);
    layer4_outputs(7366) <= not(layer3_outputs(6045));
    layer4_outputs(7367) <= not(layer3_outputs(411));
    layer4_outputs(7368) <= layer3_outputs(3501);
    layer4_outputs(7369) <= not((layer3_outputs(2040)) and (layer3_outputs(4125)));
    layer4_outputs(7370) <= not((layer3_outputs(2701)) xor (layer3_outputs(2763)));
    layer4_outputs(7371) <= not(layer3_outputs(6430)) or (layer3_outputs(1166));
    layer4_outputs(7372) <= not((layer3_outputs(6665)) xor (layer3_outputs(188)));
    layer4_outputs(7373) <= not((layer3_outputs(1734)) xor (layer3_outputs(1695)));
    layer4_outputs(7374) <= not(layer3_outputs(4434));
    layer4_outputs(7375) <= not(layer3_outputs(2420));
    layer4_outputs(7376) <= layer3_outputs(7571);
    layer4_outputs(7377) <= (layer3_outputs(333)) or (layer3_outputs(1240));
    layer4_outputs(7378) <= not(layer3_outputs(5711));
    layer4_outputs(7379) <= (layer3_outputs(1433)) and not (layer3_outputs(3550));
    layer4_outputs(7380) <= not(layer3_outputs(511));
    layer4_outputs(7381) <= (layer3_outputs(522)) or (layer3_outputs(6178));
    layer4_outputs(7382) <= not((layer3_outputs(5301)) or (layer3_outputs(7658)));
    layer4_outputs(7383) <= not((layer3_outputs(7138)) xor (layer3_outputs(7447)));
    layer4_outputs(7384) <= not(layer3_outputs(751));
    layer4_outputs(7385) <= not(layer3_outputs(5006));
    layer4_outputs(7386) <= not(layer3_outputs(2748));
    layer4_outputs(7387) <= (layer3_outputs(1297)) or (layer3_outputs(2298));
    layer4_outputs(7388) <= layer3_outputs(7359);
    layer4_outputs(7389) <= layer3_outputs(3457);
    layer4_outputs(7390) <= not(layer3_outputs(4962)) or (layer3_outputs(75));
    layer4_outputs(7391) <= not(layer3_outputs(671)) or (layer3_outputs(670));
    layer4_outputs(7392) <= (layer3_outputs(4935)) and (layer3_outputs(3320));
    layer4_outputs(7393) <= layer3_outputs(2006);
    layer4_outputs(7394) <= not((layer3_outputs(3517)) and (layer3_outputs(3381)));
    layer4_outputs(7395) <= (layer3_outputs(3302)) or (layer3_outputs(5650));
    layer4_outputs(7396) <= layer3_outputs(5838);
    layer4_outputs(7397) <= (layer3_outputs(1093)) and not (layer3_outputs(5637));
    layer4_outputs(7398) <= not(layer3_outputs(4006));
    layer4_outputs(7399) <= (layer3_outputs(107)) and (layer3_outputs(2752));
    layer4_outputs(7400) <= not((layer3_outputs(2413)) or (layer3_outputs(803)));
    layer4_outputs(7401) <= '1';
    layer4_outputs(7402) <= (layer3_outputs(5307)) and not (layer3_outputs(1754));
    layer4_outputs(7403) <= (layer3_outputs(2935)) and (layer3_outputs(4974));
    layer4_outputs(7404) <= not((layer3_outputs(5342)) and (layer3_outputs(4256)));
    layer4_outputs(7405) <= not((layer3_outputs(5979)) or (layer3_outputs(2542)));
    layer4_outputs(7406) <= not(layer3_outputs(6725));
    layer4_outputs(7407) <= not(layer3_outputs(712));
    layer4_outputs(7408) <= (layer3_outputs(6854)) or (layer3_outputs(1535));
    layer4_outputs(7409) <= layer3_outputs(5785);
    layer4_outputs(7410) <= not((layer3_outputs(1053)) or (layer3_outputs(5937)));
    layer4_outputs(7411) <= not((layer3_outputs(5878)) or (layer3_outputs(5726)));
    layer4_outputs(7412) <= (layer3_outputs(681)) and (layer3_outputs(3675));
    layer4_outputs(7413) <= not(layer3_outputs(4087));
    layer4_outputs(7414) <= (layer3_outputs(1480)) and not (layer3_outputs(2174));
    layer4_outputs(7415) <= not(layer3_outputs(1105));
    layer4_outputs(7416) <= not((layer3_outputs(2629)) or (layer3_outputs(3854)));
    layer4_outputs(7417) <= not(layer3_outputs(770));
    layer4_outputs(7418) <= layer3_outputs(3243);
    layer4_outputs(7419) <= not(layer3_outputs(6102));
    layer4_outputs(7420) <= (layer3_outputs(640)) or (layer3_outputs(6772));
    layer4_outputs(7421) <= not(layer3_outputs(1941)) or (layer3_outputs(360));
    layer4_outputs(7422) <= not((layer3_outputs(2729)) or (layer3_outputs(5921)));
    layer4_outputs(7423) <= (layer3_outputs(4008)) xor (layer3_outputs(5997));
    layer4_outputs(7424) <= not(layer3_outputs(1548));
    layer4_outputs(7425) <= (layer3_outputs(2511)) and not (layer3_outputs(6866));
    layer4_outputs(7426) <= (layer3_outputs(2750)) and not (layer3_outputs(2247));
    layer4_outputs(7427) <= layer3_outputs(647);
    layer4_outputs(7428) <= layer3_outputs(4478);
    layer4_outputs(7429) <= not(layer3_outputs(7403));
    layer4_outputs(7430) <= not(layer3_outputs(2223)) or (layer3_outputs(1696));
    layer4_outputs(7431) <= not((layer3_outputs(2510)) or (layer3_outputs(2407)));
    layer4_outputs(7432) <= (layer3_outputs(2536)) xor (layer3_outputs(2237));
    layer4_outputs(7433) <= (layer3_outputs(4202)) and (layer3_outputs(2121));
    layer4_outputs(7434) <= (layer3_outputs(3720)) xor (layer3_outputs(7252));
    layer4_outputs(7435) <= not((layer3_outputs(5489)) or (layer3_outputs(2829)));
    layer4_outputs(7436) <= (layer3_outputs(2301)) and not (layer3_outputs(6925));
    layer4_outputs(7437) <= not(layer3_outputs(5417));
    layer4_outputs(7438) <= not(layer3_outputs(3863));
    layer4_outputs(7439) <= layer3_outputs(142);
    layer4_outputs(7440) <= not(layer3_outputs(5321)) or (layer3_outputs(2618));
    layer4_outputs(7441) <= not(layer3_outputs(3042));
    layer4_outputs(7442) <= not((layer3_outputs(4412)) and (layer3_outputs(169)));
    layer4_outputs(7443) <= (layer3_outputs(2717)) xor (layer3_outputs(4277));
    layer4_outputs(7444) <= layer3_outputs(894);
    layer4_outputs(7445) <= (layer3_outputs(7379)) or (layer3_outputs(7471));
    layer4_outputs(7446) <= (layer3_outputs(3103)) or (layer3_outputs(5819));
    layer4_outputs(7447) <= not(layer3_outputs(4449));
    layer4_outputs(7448) <= (layer3_outputs(2240)) or (layer3_outputs(4558));
    layer4_outputs(7449) <= not(layer3_outputs(6137)) or (layer3_outputs(5626));
    layer4_outputs(7450) <= layer3_outputs(4174);
    layer4_outputs(7451) <= layer3_outputs(2216);
    layer4_outputs(7452) <= (layer3_outputs(5583)) xor (layer3_outputs(6435));
    layer4_outputs(7453) <= (layer3_outputs(7051)) and not (layer3_outputs(3602));
    layer4_outputs(7454) <= (layer3_outputs(5315)) xor (layer3_outputs(63));
    layer4_outputs(7455) <= not(layer3_outputs(751)) or (layer3_outputs(454));
    layer4_outputs(7456) <= not(layer3_outputs(6768));
    layer4_outputs(7457) <= not(layer3_outputs(3044));
    layer4_outputs(7458) <= layer3_outputs(2734);
    layer4_outputs(7459) <= layer3_outputs(3974);
    layer4_outputs(7460) <= not((layer3_outputs(3362)) or (layer3_outputs(5814)));
    layer4_outputs(7461) <= not((layer3_outputs(6472)) and (layer3_outputs(4553)));
    layer4_outputs(7462) <= layer3_outputs(6994);
    layer4_outputs(7463) <= (layer3_outputs(141)) and not (layer3_outputs(7428));
    layer4_outputs(7464) <= not(layer3_outputs(3726));
    layer4_outputs(7465) <= not(layer3_outputs(3445)) or (layer3_outputs(640));
    layer4_outputs(7466) <= (layer3_outputs(653)) xor (layer3_outputs(6532));
    layer4_outputs(7467) <= (layer3_outputs(7302)) xor (layer3_outputs(1671));
    layer4_outputs(7468) <= (layer3_outputs(6176)) and not (layer3_outputs(1072));
    layer4_outputs(7469) <= layer3_outputs(3561);
    layer4_outputs(7470) <= not(layer3_outputs(912));
    layer4_outputs(7471) <= (layer3_outputs(6391)) xor (layer3_outputs(95));
    layer4_outputs(7472) <= (layer3_outputs(7536)) and not (layer3_outputs(2851));
    layer4_outputs(7473) <= layer3_outputs(4299);
    layer4_outputs(7474) <= (layer3_outputs(3154)) and not (layer3_outputs(5069));
    layer4_outputs(7475) <= (layer3_outputs(2323)) xor (layer3_outputs(7318));
    layer4_outputs(7476) <= (layer3_outputs(6965)) and (layer3_outputs(4570));
    layer4_outputs(7477) <= not(layer3_outputs(6427));
    layer4_outputs(7478) <= not(layer3_outputs(1274));
    layer4_outputs(7479) <= not(layer3_outputs(6539)) or (layer3_outputs(1972));
    layer4_outputs(7480) <= not(layer3_outputs(2200));
    layer4_outputs(7481) <= (layer3_outputs(2997)) or (layer3_outputs(3794));
    layer4_outputs(7482) <= not(layer3_outputs(6132));
    layer4_outputs(7483) <= '1';
    layer4_outputs(7484) <= not(layer3_outputs(5777));
    layer4_outputs(7485) <= not(layer3_outputs(7031)) or (layer3_outputs(233));
    layer4_outputs(7486) <= (layer3_outputs(4086)) and not (layer3_outputs(2771));
    layer4_outputs(7487) <= not((layer3_outputs(5186)) and (layer3_outputs(7567)));
    layer4_outputs(7488) <= not((layer3_outputs(6939)) xor (layer3_outputs(5475)));
    layer4_outputs(7489) <= (layer3_outputs(4248)) and not (layer3_outputs(4127));
    layer4_outputs(7490) <= not(layer3_outputs(1415));
    layer4_outputs(7491) <= not(layer3_outputs(3624));
    layer4_outputs(7492) <= not((layer3_outputs(578)) and (layer3_outputs(4984)));
    layer4_outputs(7493) <= not(layer3_outputs(1889)) or (layer3_outputs(891));
    layer4_outputs(7494) <= not(layer3_outputs(8));
    layer4_outputs(7495) <= (layer3_outputs(3512)) and not (layer3_outputs(1763));
    layer4_outputs(7496) <= not(layer3_outputs(4147));
    layer4_outputs(7497) <= not(layer3_outputs(6802));
    layer4_outputs(7498) <= layer3_outputs(5897);
    layer4_outputs(7499) <= not((layer3_outputs(5016)) and (layer3_outputs(7631)));
    layer4_outputs(7500) <= layer3_outputs(3736);
    layer4_outputs(7501) <= (layer3_outputs(5165)) and not (layer3_outputs(4612));
    layer4_outputs(7502) <= (layer3_outputs(2784)) and (layer3_outputs(3076));
    layer4_outputs(7503) <= not((layer3_outputs(729)) or (layer3_outputs(72)));
    layer4_outputs(7504) <= layer3_outputs(1917);
    layer4_outputs(7505) <= not(layer3_outputs(5293));
    layer4_outputs(7506) <= (layer3_outputs(2295)) or (layer3_outputs(3265));
    layer4_outputs(7507) <= layer3_outputs(1801);
    layer4_outputs(7508) <= (layer3_outputs(5101)) or (layer3_outputs(5779));
    layer4_outputs(7509) <= layer3_outputs(4876);
    layer4_outputs(7510) <= (layer3_outputs(5972)) and (layer3_outputs(1688));
    layer4_outputs(7511) <= not(layer3_outputs(4273));
    layer4_outputs(7512) <= not(layer3_outputs(5375)) or (layer3_outputs(1366));
    layer4_outputs(7513) <= not((layer3_outputs(3297)) and (layer3_outputs(84)));
    layer4_outputs(7514) <= layer3_outputs(3502);
    layer4_outputs(7515) <= not((layer3_outputs(3426)) xor (layer3_outputs(5244)));
    layer4_outputs(7516) <= layer3_outputs(425);
    layer4_outputs(7517) <= not(layer3_outputs(950));
    layer4_outputs(7518) <= not(layer3_outputs(745)) or (layer3_outputs(6069));
    layer4_outputs(7519) <= not(layer3_outputs(1543)) or (layer3_outputs(1506));
    layer4_outputs(7520) <= not(layer3_outputs(869));
    layer4_outputs(7521) <= not((layer3_outputs(532)) xor (layer3_outputs(6304)));
    layer4_outputs(7522) <= not(layer3_outputs(49));
    layer4_outputs(7523) <= (layer3_outputs(4794)) and (layer3_outputs(6232));
    layer4_outputs(7524) <= (layer3_outputs(7573)) and (layer3_outputs(6736));
    layer4_outputs(7525) <= '0';
    layer4_outputs(7526) <= not((layer3_outputs(6715)) and (layer3_outputs(6660)));
    layer4_outputs(7527) <= layer3_outputs(4723);
    layer4_outputs(7528) <= layer3_outputs(2800);
    layer4_outputs(7529) <= not(layer3_outputs(5525));
    layer4_outputs(7530) <= layer3_outputs(2930);
    layer4_outputs(7531) <= not(layer3_outputs(2105));
    layer4_outputs(7532) <= layer3_outputs(5462);
    layer4_outputs(7533) <= not(layer3_outputs(5495));
    layer4_outputs(7534) <= not(layer3_outputs(2462)) or (layer3_outputs(3187));
    layer4_outputs(7535) <= layer3_outputs(6119);
    layer4_outputs(7536) <= layer3_outputs(1875);
    layer4_outputs(7537) <= layer3_outputs(1961);
    layer4_outputs(7538) <= not(layer3_outputs(7070));
    layer4_outputs(7539) <= layer3_outputs(4268);
    layer4_outputs(7540) <= (layer3_outputs(4852)) and not (layer3_outputs(2666));
    layer4_outputs(7541) <= not((layer3_outputs(4683)) and (layer3_outputs(70)));
    layer4_outputs(7542) <= not(layer3_outputs(1286));
    layer4_outputs(7543) <= not(layer3_outputs(499));
    layer4_outputs(7544) <= not((layer3_outputs(4752)) and (layer3_outputs(1841)));
    layer4_outputs(7545) <= '1';
    layer4_outputs(7546) <= not((layer3_outputs(7423)) xor (layer3_outputs(5315)));
    layer4_outputs(7547) <= not(layer3_outputs(2035));
    layer4_outputs(7548) <= not(layer3_outputs(840)) or (layer3_outputs(4515));
    layer4_outputs(7549) <= not(layer3_outputs(4897));
    layer4_outputs(7550) <= layer3_outputs(6509);
    layer4_outputs(7551) <= not(layer3_outputs(800));
    layer4_outputs(7552) <= (layer3_outputs(5417)) or (layer3_outputs(7106));
    layer4_outputs(7553) <= layer3_outputs(2769);
    layer4_outputs(7554) <= not(layer3_outputs(3860));
    layer4_outputs(7555) <= not((layer3_outputs(6204)) and (layer3_outputs(7190)));
    layer4_outputs(7556) <= layer3_outputs(1557);
    layer4_outputs(7557) <= (layer3_outputs(5579)) xor (layer3_outputs(5850));
    layer4_outputs(7558) <= layer3_outputs(7457);
    layer4_outputs(7559) <= layer3_outputs(911);
    layer4_outputs(7560) <= not((layer3_outputs(3364)) xor (layer3_outputs(4251)));
    layer4_outputs(7561) <= not(layer3_outputs(5285));
    layer4_outputs(7562) <= not(layer3_outputs(7100)) or (layer3_outputs(3748));
    layer4_outputs(7563) <= not(layer3_outputs(6669));
    layer4_outputs(7564) <= layer3_outputs(5525);
    layer4_outputs(7565) <= layer3_outputs(2742);
    layer4_outputs(7566) <= (layer3_outputs(530)) and not (layer3_outputs(2756));
    layer4_outputs(7567) <= layer3_outputs(635);
    layer4_outputs(7568) <= not((layer3_outputs(3376)) and (layer3_outputs(7109)));
    layer4_outputs(7569) <= not(layer3_outputs(1594));
    layer4_outputs(7570) <= not(layer3_outputs(3652)) or (layer3_outputs(3546));
    layer4_outputs(7571) <= (layer3_outputs(1063)) or (layer3_outputs(3659));
    layer4_outputs(7572) <= layer3_outputs(470);
    layer4_outputs(7573) <= (layer3_outputs(2958)) or (layer3_outputs(329));
    layer4_outputs(7574) <= not(layer3_outputs(1919));
    layer4_outputs(7575) <= not(layer3_outputs(7082));
    layer4_outputs(7576) <= not(layer3_outputs(3152));
    layer4_outputs(7577) <= not(layer3_outputs(3407));
    layer4_outputs(7578) <= not(layer3_outputs(292));
    layer4_outputs(7579) <= (layer3_outputs(4937)) or (layer3_outputs(1807));
    layer4_outputs(7580) <= (layer3_outputs(4373)) or (layer3_outputs(2669));
    layer4_outputs(7581) <= not((layer3_outputs(6690)) or (layer3_outputs(3519)));
    layer4_outputs(7582) <= (layer3_outputs(3855)) and not (layer3_outputs(3987));
    layer4_outputs(7583) <= layer3_outputs(6473);
    layer4_outputs(7584) <= (layer3_outputs(152)) and (layer3_outputs(1462));
    layer4_outputs(7585) <= layer3_outputs(3590);
    layer4_outputs(7586) <= layer3_outputs(3751);
    layer4_outputs(7587) <= (layer3_outputs(2691)) and (layer3_outputs(170));
    layer4_outputs(7588) <= not(layer3_outputs(2847));
    layer4_outputs(7589) <= not(layer3_outputs(6795));
    layer4_outputs(7590) <= not(layer3_outputs(6407));
    layer4_outputs(7591) <= not(layer3_outputs(1913));
    layer4_outputs(7592) <= not((layer3_outputs(2551)) xor (layer3_outputs(2382)));
    layer4_outputs(7593) <= (layer3_outputs(512)) or (layer3_outputs(2751));
    layer4_outputs(7594) <= layer3_outputs(2815);
    layer4_outputs(7595) <= (layer3_outputs(702)) or (layer3_outputs(5472));
    layer4_outputs(7596) <= layer3_outputs(1512);
    layer4_outputs(7597) <= (layer3_outputs(301)) or (layer3_outputs(288));
    layer4_outputs(7598) <= (layer3_outputs(5526)) and not (layer3_outputs(3448));
    layer4_outputs(7599) <= not(layer3_outputs(3143)) or (layer3_outputs(3271));
    layer4_outputs(7600) <= not(layer3_outputs(1377)) or (layer3_outputs(4341));
    layer4_outputs(7601) <= (layer3_outputs(166)) xor (layer3_outputs(2509));
    layer4_outputs(7602) <= (layer3_outputs(5739)) and not (layer3_outputs(3906));
    layer4_outputs(7603) <= layer3_outputs(4661);
    layer4_outputs(7604) <= (layer3_outputs(4941)) xor (layer3_outputs(5962));
    layer4_outputs(7605) <= (layer3_outputs(2844)) and not (layer3_outputs(1525));
    layer4_outputs(7606) <= not((layer3_outputs(904)) xor (layer3_outputs(1894)));
    layer4_outputs(7607) <= layer3_outputs(5124);
    layer4_outputs(7608) <= not((layer3_outputs(2849)) or (layer3_outputs(5786)));
    layer4_outputs(7609) <= layer3_outputs(2743);
    layer4_outputs(7610) <= not((layer3_outputs(5720)) or (layer3_outputs(204)));
    layer4_outputs(7611) <= (layer3_outputs(4382)) and not (layer3_outputs(4610));
    layer4_outputs(7612) <= (layer3_outputs(1638)) and (layer3_outputs(6556));
    layer4_outputs(7613) <= not(layer3_outputs(6530));
    layer4_outputs(7614) <= layer3_outputs(288);
    layer4_outputs(7615) <= (layer3_outputs(5273)) xor (layer3_outputs(1221));
    layer4_outputs(7616) <= (layer3_outputs(3382)) xor (layer3_outputs(7385));
    layer4_outputs(7617) <= (layer3_outputs(1836)) and not (layer3_outputs(4362));
    layer4_outputs(7618) <= not((layer3_outputs(1411)) and (layer3_outputs(3654)));
    layer4_outputs(7619) <= (layer3_outputs(1891)) and (layer3_outputs(5118));
    layer4_outputs(7620) <= (layer3_outputs(5713)) xor (layer3_outputs(2727));
    layer4_outputs(7621) <= not((layer3_outputs(3145)) and (layer3_outputs(4145)));
    layer4_outputs(7622) <= (layer3_outputs(4072)) and (layer3_outputs(5022));
    layer4_outputs(7623) <= layer3_outputs(1691);
    layer4_outputs(7624) <= (layer3_outputs(1420)) and not (layer3_outputs(5237));
    layer4_outputs(7625) <= not((layer3_outputs(7298)) xor (layer3_outputs(1131)));
    layer4_outputs(7626) <= not(layer3_outputs(7657)) or (layer3_outputs(6904));
    layer4_outputs(7627) <= (layer3_outputs(3686)) or (layer3_outputs(6721));
    layer4_outputs(7628) <= not((layer3_outputs(6605)) or (layer3_outputs(818)));
    layer4_outputs(7629) <= (layer3_outputs(5484)) and not (layer3_outputs(2524));
    layer4_outputs(7630) <= layer3_outputs(3152);
    layer4_outputs(7631) <= not(layer3_outputs(5037));
    layer4_outputs(7632) <= layer3_outputs(6636);
    layer4_outputs(7633) <= layer3_outputs(6419);
    layer4_outputs(7634) <= not(layer3_outputs(1133));
    layer4_outputs(7635) <= layer3_outputs(4766);
    layer4_outputs(7636) <= (layer3_outputs(5744)) xor (layer3_outputs(6705));
    layer4_outputs(7637) <= layer3_outputs(1939);
    layer4_outputs(7638) <= not(layer3_outputs(2197)) or (layer3_outputs(3962));
    layer4_outputs(7639) <= (layer3_outputs(4596)) and not (layer3_outputs(3607));
    layer4_outputs(7640) <= not(layer3_outputs(6193)) or (layer3_outputs(4210));
    layer4_outputs(7641) <= not(layer3_outputs(4296));
    layer4_outputs(7642) <= (layer3_outputs(5613)) and not (layer3_outputs(7022));
    layer4_outputs(7643) <= not(layer3_outputs(5084));
    layer4_outputs(7644) <= not((layer3_outputs(4486)) or (layer3_outputs(6223)));
    layer4_outputs(7645) <= layer3_outputs(3122);
    layer4_outputs(7646) <= not(layer3_outputs(4745)) or (layer3_outputs(4895));
    layer4_outputs(7647) <= layer3_outputs(4650);
    layer4_outputs(7648) <= (layer3_outputs(742)) and not (layer3_outputs(3120));
    layer4_outputs(7649) <= layer3_outputs(3495);
    layer4_outputs(7650) <= not(layer3_outputs(7402));
    layer4_outputs(7651) <= (layer3_outputs(3157)) or (layer3_outputs(4986));
    layer4_outputs(7652) <= not(layer3_outputs(1891));
    layer4_outputs(7653) <= not(layer3_outputs(5401));
    layer4_outputs(7654) <= not(layer3_outputs(4864));
    layer4_outputs(7655) <= (layer3_outputs(1405)) or (layer3_outputs(6056));
    layer4_outputs(7656) <= (layer3_outputs(486)) and (layer3_outputs(2785));
    layer4_outputs(7657) <= layer3_outputs(2073);
    layer4_outputs(7658) <= not(layer3_outputs(3898)) or (layer3_outputs(5547));
    layer4_outputs(7659) <= not(layer3_outputs(18));
    layer4_outputs(7660) <= not(layer3_outputs(5234));
    layer4_outputs(7661) <= layer3_outputs(7504);
    layer4_outputs(7662) <= not(layer3_outputs(2254)) or (layer3_outputs(2782));
    layer4_outputs(7663) <= layer3_outputs(3055);
    layer4_outputs(7664) <= not(layer3_outputs(1644));
    layer4_outputs(7665) <= not((layer3_outputs(835)) xor (layer3_outputs(1556)));
    layer4_outputs(7666) <= layer3_outputs(1661);
    layer4_outputs(7667) <= layer3_outputs(6147);
    layer4_outputs(7668) <= not(layer3_outputs(6473));
    layer4_outputs(7669) <= not(layer3_outputs(1096)) or (layer3_outputs(3503));
    layer4_outputs(7670) <= not(layer3_outputs(4330)) or (layer3_outputs(2436));
    layer4_outputs(7671) <= not((layer3_outputs(894)) or (layer3_outputs(7526)));
    layer4_outputs(7672) <= layer3_outputs(6136);
    layer4_outputs(7673) <= layer3_outputs(895);
    layer4_outputs(7674) <= layer3_outputs(1894);
    layer4_outputs(7675) <= not(layer3_outputs(1895)) or (layer3_outputs(6151));
    layer4_outputs(7676) <= not(layer3_outputs(1583));
    layer4_outputs(7677) <= not(layer3_outputs(5805));
    layer4_outputs(7678) <= (layer3_outputs(5156)) or (layer3_outputs(7529));
    layer4_outputs(7679) <= layer3_outputs(5787);
    outputs(0) <= not(layer4_outputs(2377));
    outputs(1) <= not(layer4_outputs(60));
    outputs(2) <= layer4_outputs(581);
    outputs(3) <= (layer4_outputs(2053)) xor (layer4_outputs(6358));
    outputs(4) <= not((layer4_outputs(7405)) or (layer4_outputs(7149)));
    outputs(5) <= not(layer4_outputs(469));
    outputs(6) <= (layer4_outputs(6594)) xor (layer4_outputs(6418));
    outputs(7) <= not(layer4_outputs(3985));
    outputs(8) <= not((layer4_outputs(4044)) xor (layer4_outputs(5058)));
    outputs(9) <= not((layer4_outputs(5273)) or (layer4_outputs(4837)));
    outputs(10) <= (layer4_outputs(2835)) and (layer4_outputs(3487));
    outputs(11) <= not(layer4_outputs(5918));
    outputs(12) <= (layer4_outputs(1214)) and (layer4_outputs(6821));
    outputs(13) <= not(layer4_outputs(1012));
    outputs(14) <= (layer4_outputs(1463)) xor (layer4_outputs(1591));
    outputs(15) <= layer4_outputs(2052);
    outputs(16) <= not((layer4_outputs(2967)) xor (layer4_outputs(6557)));
    outputs(17) <= not(layer4_outputs(66));
    outputs(18) <= (layer4_outputs(2669)) and not (layer4_outputs(1055));
    outputs(19) <= layer4_outputs(6009);
    outputs(20) <= not(layer4_outputs(5670));
    outputs(21) <= layer4_outputs(6040);
    outputs(22) <= layer4_outputs(7157);
    outputs(23) <= (layer4_outputs(261)) and not (layer4_outputs(7521));
    outputs(24) <= layer4_outputs(1096);
    outputs(25) <= layer4_outputs(6892);
    outputs(26) <= not(layer4_outputs(7314));
    outputs(27) <= not(layer4_outputs(5096));
    outputs(28) <= layer4_outputs(7663);
    outputs(29) <= not((layer4_outputs(5079)) xor (layer4_outputs(3660)));
    outputs(30) <= layer4_outputs(2797);
    outputs(31) <= not((layer4_outputs(7620)) and (layer4_outputs(5833)));
    outputs(32) <= not(layer4_outputs(6662));
    outputs(33) <= not(layer4_outputs(4163)) or (layer4_outputs(891));
    outputs(34) <= (layer4_outputs(135)) and (layer4_outputs(5525));
    outputs(35) <= layer4_outputs(1117);
    outputs(36) <= not(layer4_outputs(5766));
    outputs(37) <= layer4_outputs(2497);
    outputs(38) <= layer4_outputs(817);
    outputs(39) <= not((layer4_outputs(360)) xor (layer4_outputs(5101)));
    outputs(40) <= not(layer4_outputs(4055));
    outputs(41) <= not(layer4_outputs(6095));
    outputs(42) <= not(layer4_outputs(3325));
    outputs(43) <= (layer4_outputs(6075)) xor (layer4_outputs(1749));
    outputs(44) <= layer4_outputs(7176);
    outputs(45) <= not(layer4_outputs(2242));
    outputs(46) <= layer4_outputs(4754);
    outputs(47) <= not((layer4_outputs(5510)) xor (layer4_outputs(1070)));
    outputs(48) <= not(layer4_outputs(6843));
    outputs(49) <= not(layer4_outputs(886));
    outputs(50) <= not(layer4_outputs(4153));
    outputs(51) <= not(layer4_outputs(3650)) or (layer4_outputs(1833));
    outputs(52) <= (layer4_outputs(2749)) or (layer4_outputs(5169));
    outputs(53) <= layer4_outputs(1260);
    outputs(54) <= layer4_outputs(2323);
    outputs(55) <= (layer4_outputs(7481)) xor (layer4_outputs(1097));
    outputs(56) <= not((layer4_outputs(5679)) or (layer4_outputs(2090)));
    outputs(57) <= (layer4_outputs(4593)) and not (layer4_outputs(2188));
    outputs(58) <= not(layer4_outputs(1777));
    outputs(59) <= layer4_outputs(7632);
    outputs(60) <= layer4_outputs(7530);
    outputs(61) <= layer4_outputs(5860);
    outputs(62) <= (layer4_outputs(3703)) xor (layer4_outputs(2045));
    outputs(63) <= (layer4_outputs(450)) and not (layer4_outputs(2509));
    outputs(64) <= layer4_outputs(1322);
    outputs(65) <= not((layer4_outputs(3180)) xor (layer4_outputs(6248)));
    outputs(66) <= (layer4_outputs(1649)) and (layer4_outputs(3396));
    outputs(67) <= not(layer4_outputs(2321));
    outputs(68) <= layer4_outputs(3107);
    outputs(69) <= layer4_outputs(5334);
    outputs(70) <= not((layer4_outputs(5694)) xor (layer4_outputs(5667)));
    outputs(71) <= (layer4_outputs(5361)) xor (layer4_outputs(1498));
    outputs(72) <= not(layer4_outputs(7370));
    outputs(73) <= layer4_outputs(2172);
    outputs(74) <= (layer4_outputs(6048)) and not (layer4_outputs(548));
    outputs(75) <= layer4_outputs(5523);
    outputs(76) <= layer4_outputs(5954);
    outputs(77) <= layer4_outputs(1130);
    outputs(78) <= not(layer4_outputs(2043)) or (layer4_outputs(2489));
    outputs(79) <= not((layer4_outputs(249)) and (layer4_outputs(2118)));
    outputs(80) <= (layer4_outputs(3607)) xor (layer4_outputs(4501));
    outputs(81) <= not((layer4_outputs(6507)) xor (layer4_outputs(1174)));
    outputs(82) <= (layer4_outputs(6545)) xor (layer4_outputs(2764));
    outputs(83) <= layer4_outputs(934);
    outputs(84) <= layer4_outputs(4254);
    outputs(85) <= not(layer4_outputs(7320));
    outputs(86) <= (layer4_outputs(2229)) xor (layer4_outputs(3546));
    outputs(87) <= layer4_outputs(6375);
    outputs(88) <= not((layer4_outputs(872)) or (layer4_outputs(3654)));
    outputs(89) <= layer4_outputs(854);
    outputs(90) <= layer4_outputs(5465);
    outputs(91) <= not(layer4_outputs(2429));
    outputs(92) <= not(layer4_outputs(6725));
    outputs(93) <= not(layer4_outputs(1764));
    outputs(94) <= not(layer4_outputs(6578));
    outputs(95) <= layer4_outputs(419);
    outputs(96) <= not(layer4_outputs(2237));
    outputs(97) <= not(layer4_outputs(5888));
    outputs(98) <= layer4_outputs(4097);
    outputs(99) <= (layer4_outputs(3341)) xor (layer4_outputs(2058));
    outputs(100) <= layer4_outputs(4325);
    outputs(101) <= not(layer4_outputs(3154));
    outputs(102) <= not(layer4_outputs(1855));
    outputs(103) <= not(layer4_outputs(2753));
    outputs(104) <= not(layer4_outputs(1032));
    outputs(105) <= (layer4_outputs(5830)) xor (layer4_outputs(2580));
    outputs(106) <= not(layer4_outputs(5452));
    outputs(107) <= layer4_outputs(3965);
    outputs(108) <= not(layer4_outputs(6713));
    outputs(109) <= layer4_outputs(5507);
    outputs(110) <= layer4_outputs(1454);
    outputs(111) <= not((layer4_outputs(6804)) xor (layer4_outputs(6379)));
    outputs(112) <= not(layer4_outputs(3945));
    outputs(113) <= layer4_outputs(857);
    outputs(114) <= layer4_outputs(1163);
    outputs(115) <= not(layer4_outputs(6871));
    outputs(116) <= not((layer4_outputs(6230)) xor (layer4_outputs(7588)));
    outputs(117) <= layer4_outputs(4433);
    outputs(118) <= not((layer4_outputs(5579)) xor (layer4_outputs(72)));
    outputs(119) <= not((layer4_outputs(5510)) xor (layer4_outputs(191)));
    outputs(120) <= layer4_outputs(277);
    outputs(121) <= not(layer4_outputs(7473));
    outputs(122) <= (layer4_outputs(6655)) or (layer4_outputs(1849));
    outputs(123) <= layer4_outputs(7475);
    outputs(124) <= layer4_outputs(1923);
    outputs(125) <= not(layer4_outputs(5756));
    outputs(126) <= (layer4_outputs(6361)) and (layer4_outputs(488));
    outputs(127) <= (layer4_outputs(2336)) and not (layer4_outputs(3713));
    outputs(128) <= not(layer4_outputs(6254)) or (layer4_outputs(6541));
    outputs(129) <= layer4_outputs(7180);
    outputs(130) <= not(layer4_outputs(1550));
    outputs(131) <= (layer4_outputs(811)) and not (layer4_outputs(4221));
    outputs(132) <= not((layer4_outputs(3526)) xor (layer4_outputs(1948)));
    outputs(133) <= not(layer4_outputs(3582));
    outputs(134) <= layer4_outputs(2563);
    outputs(135) <= layer4_outputs(6252);
    outputs(136) <= layer4_outputs(7233);
    outputs(137) <= layer4_outputs(4788);
    outputs(138) <= not((layer4_outputs(7231)) or (layer4_outputs(3072)));
    outputs(139) <= layer4_outputs(2350);
    outputs(140) <= not(layer4_outputs(5855));
    outputs(141) <= (layer4_outputs(5401)) and not (layer4_outputs(3145));
    outputs(142) <= layer4_outputs(4756);
    outputs(143) <= layer4_outputs(5450);
    outputs(144) <= not(layer4_outputs(4648));
    outputs(145) <= layer4_outputs(7056);
    outputs(146) <= layer4_outputs(7497);
    outputs(147) <= not((layer4_outputs(2431)) or (layer4_outputs(1253)));
    outputs(148) <= (layer4_outputs(6745)) xor (layer4_outputs(1533));
    outputs(149) <= not((layer4_outputs(4760)) xor (layer4_outputs(6090)));
    outputs(150) <= layer4_outputs(3050);
    outputs(151) <= not((layer4_outputs(120)) xor (layer4_outputs(4311)));
    outputs(152) <= layer4_outputs(6320);
    outputs(153) <= not((layer4_outputs(4843)) and (layer4_outputs(5907)));
    outputs(154) <= layer4_outputs(2919);
    outputs(155) <= not((layer4_outputs(3642)) xor (layer4_outputs(6894)));
    outputs(156) <= not(layer4_outputs(2969));
    outputs(157) <= not(layer4_outputs(667));
    outputs(158) <= layer4_outputs(3600);
    outputs(159) <= layer4_outputs(5812);
    outputs(160) <= not(layer4_outputs(1572));
    outputs(161) <= not(layer4_outputs(2047));
    outputs(162) <= (layer4_outputs(3732)) and (layer4_outputs(1787));
    outputs(163) <= not(layer4_outputs(5183));
    outputs(164) <= not(layer4_outputs(7564));
    outputs(165) <= layer4_outputs(6570);
    outputs(166) <= (layer4_outputs(2662)) and (layer4_outputs(3156));
    outputs(167) <= not(layer4_outputs(5215));
    outputs(168) <= not(layer4_outputs(5622));
    outputs(169) <= (layer4_outputs(415)) xor (layer4_outputs(3061));
    outputs(170) <= not(layer4_outputs(6522));
    outputs(171) <= not((layer4_outputs(5367)) or (layer4_outputs(5108)));
    outputs(172) <= not((layer4_outputs(2511)) xor (layer4_outputs(466)));
    outputs(173) <= layer4_outputs(5838);
    outputs(174) <= layer4_outputs(3134);
    outputs(175) <= layer4_outputs(1150);
    outputs(176) <= not((layer4_outputs(5814)) and (layer4_outputs(657)));
    outputs(177) <= not(layer4_outputs(361));
    outputs(178) <= not(layer4_outputs(4827));
    outputs(179) <= layer4_outputs(6794);
    outputs(180) <= (layer4_outputs(3987)) xor (layer4_outputs(7397));
    outputs(181) <= not((layer4_outputs(456)) xor (layer4_outputs(4563)));
    outputs(182) <= not((layer4_outputs(4003)) xor (layer4_outputs(3875)));
    outputs(183) <= (layer4_outputs(7676)) and (layer4_outputs(6759));
    outputs(184) <= layer4_outputs(5370);
    outputs(185) <= not((layer4_outputs(2955)) and (layer4_outputs(290)));
    outputs(186) <= layer4_outputs(6081);
    outputs(187) <= (layer4_outputs(3211)) or (layer4_outputs(1332));
    outputs(188) <= layer4_outputs(4772);
    outputs(189) <= not(layer4_outputs(2710));
    outputs(190) <= not(layer4_outputs(3267));
    outputs(191) <= not(layer4_outputs(6038));
    outputs(192) <= layer4_outputs(2);
    outputs(193) <= (layer4_outputs(438)) and not (layer4_outputs(4410));
    outputs(194) <= not(layer4_outputs(1481));
    outputs(195) <= not((layer4_outputs(3947)) xor (layer4_outputs(4408)));
    outputs(196) <= layer4_outputs(2170);
    outputs(197) <= not((layer4_outputs(3584)) xor (layer4_outputs(4281)));
    outputs(198) <= layer4_outputs(7050);
    outputs(199) <= (layer4_outputs(2238)) and not (layer4_outputs(2842));
    outputs(200) <= not((layer4_outputs(4550)) or (layer4_outputs(2761)));
    outputs(201) <= layer4_outputs(2025);
    outputs(202) <= (layer4_outputs(474)) and not (layer4_outputs(5723));
    outputs(203) <= layer4_outputs(4341);
    outputs(204) <= layer4_outputs(143);
    outputs(205) <= layer4_outputs(4584);
    outputs(206) <= (layer4_outputs(5160)) xor (layer4_outputs(5377));
    outputs(207) <= (layer4_outputs(5536)) xor (layer4_outputs(5980));
    outputs(208) <= (layer4_outputs(1471)) and not (layer4_outputs(5651));
    outputs(209) <= layer4_outputs(2760);
    outputs(210) <= not(layer4_outputs(2826));
    outputs(211) <= not((layer4_outputs(2204)) xor (layer4_outputs(955)));
    outputs(212) <= not(layer4_outputs(7515));
    outputs(213) <= not(layer4_outputs(4553));
    outputs(214) <= not(layer4_outputs(4167));
    outputs(215) <= layer4_outputs(5761);
    outputs(216) <= layer4_outputs(1245);
    outputs(217) <= not(layer4_outputs(5895)) or (layer4_outputs(5719));
    outputs(218) <= (layer4_outputs(1052)) xor (layer4_outputs(7429));
    outputs(219) <= layer4_outputs(1664);
    outputs(220) <= not(layer4_outputs(1497));
    outputs(221) <= not(layer4_outputs(7469));
    outputs(222) <= (layer4_outputs(3651)) and (layer4_outputs(2128));
    outputs(223) <= (layer4_outputs(7448)) xor (layer4_outputs(5742));
    outputs(224) <= not(layer4_outputs(5786));
    outputs(225) <= layer4_outputs(3864);
    outputs(226) <= layer4_outputs(5112);
    outputs(227) <= layer4_outputs(5135);
    outputs(228) <= (layer4_outputs(1536)) xor (layer4_outputs(5082));
    outputs(229) <= (layer4_outputs(453)) and not (layer4_outputs(540));
    outputs(230) <= layer4_outputs(1500);
    outputs(231) <= not(layer4_outputs(2178));
    outputs(232) <= layer4_outputs(3967);
    outputs(233) <= (layer4_outputs(635)) xor (layer4_outputs(1589));
    outputs(234) <= (layer4_outputs(2692)) and not (layer4_outputs(5664));
    outputs(235) <= layer4_outputs(5444);
    outputs(236) <= not(layer4_outputs(2603));
    outputs(237) <= not(layer4_outputs(5720));
    outputs(238) <= (layer4_outputs(297)) xor (layer4_outputs(1324));
    outputs(239) <= (layer4_outputs(5908)) xor (layer4_outputs(1807));
    outputs(240) <= not(layer4_outputs(5914));
    outputs(241) <= layer4_outputs(643);
    outputs(242) <= not(layer4_outputs(753));
    outputs(243) <= (layer4_outputs(5245)) xor (layer4_outputs(3927));
    outputs(244) <= not(layer4_outputs(2904));
    outputs(245) <= not(layer4_outputs(2268)) or (layer4_outputs(4382));
    outputs(246) <= layer4_outputs(3635);
    outputs(247) <= layer4_outputs(930);
    outputs(248) <= layer4_outputs(3192);
    outputs(249) <= not(layer4_outputs(2778));
    outputs(250) <= not(layer4_outputs(464));
    outputs(251) <= not(layer4_outputs(7462));
    outputs(252) <= (layer4_outputs(4181)) xor (layer4_outputs(7417));
    outputs(253) <= not(layer4_outputs(6489));
    outputs(254) <= not(layer4_outputs(4620));
    outputs(255) <= (layer4_outputs(240)) xor (layer4_outputs(2408));
    outputs(256) <= not((layer4_outputs(2788)) xor (layer4_outputs(7590)));
    outputs(257) <= not(layer4_outputs(6441));
    outputs(258) <= not(layer4_outputs(3019));
    outputs(259) <= not(layer4_outputs(3855));
    outputs(260) <= not(layer4_outputs(3101));
    outputs(261) <= layer4_outputs(1980);
    outputs(262) <= not(layer4_outputs(5257)) or (layer4_outputs(2815));
    outputs(263) <= not(layer4_outputs(3196));
    outputs(264) <= (layer4_outputs(3300)) and not (layer4_outputs(74));
    outputs(265) <= (layer4_outputs(6006)) and not (layer4_outputs(1185));
    outputs(266) <= layer4_outputs(7677);
    outputs(267) <= not(layer4_outputs(1518));
    outputs(268) <= not((layer4_outputs(1910)) xor (layer4_outputs(2242)));
    outputs(269) <= layer4_outputs(7094);
    outputs(270) <= (layer4_outputs(7580)) and (layer4_outputs(3016));
    outputs(271) <= not(layer4_outputs(5583));
    outputs(272) <= layer4_outputs(3409);
    outputs(273) <= not(layer4_outputs(463));
    outputs(274) <= layer4_outputs(1542);
    outputs(275) <= not(layer4_outputs(5868));
    outputs(276) <= layer4_outputs(1235);
    outputs(277) <= layer4_outputs(6911);
    outputs(278) <= not((layer4_outputs(1772)) xor (layer4_outputs(3463)));
    outputs(279) <= not(layer4_outputs(1608));
    outputs(280) <= layer4_outputs(7378);
    outputs(281) <= layer4_outputs(2383);
    outputs(282) <= layer4_outputs(4860);
    outputs(283) <= not(layer4_outputs(5733));
    outputs(284) <= not((layer4_outputs(3508)) or (layer4_outputs(5741)));
    outputs(285) <= not(layer4_outputs(7540));
    outputs(286) <= not(layer4_outputs(4684));
    outputs(287) <= not((layer4_outputs(1446)) xor (layer4_outputs(3062)));
    outputs(288) <= not((layer4_outputs(4067)) xor (layer4_outputs(6382)));
    outputs(289) <= not(layer4_outputs(815));
    outputs(290) <= layer4_outputs(6558);
    outputs(291) <= layer4_outputs(3868);
    outputs(292) <= not(layer4_outputs(7326));
    outputs(293) <= not(layer4_outputs(5570));
    outputs(294) <= not((layer4_outputs(2087)) xor (layer4_outputs(418)));
    outputs(295) <= not(layer4_outputs(6657));
    outputs(296) <= not((layer4_outputs(3741)) xor (layer4_outputs(792)));
    outputs(297) <= not((layer4_outputs(4280)) xor (layer4_outputs(4039)));
    outputs(298) <= not(layer4_outputs(6656));
    outputs(299) <= (layer4_outputs(1318)) and not (layer4_outputs(3979));
    outputs(300) <= layer4_outputs(6088);
    outputs(301) <= (layer4_outputs(4770)) xor (layer4_outputs(5759));
    outputs(302) <= not((layer4_outputs(960)) xor (layer4_outputs(3316)));
    outputs(303) <= (layer4_outputs(2844)) xor (layer4_outputs(4099));
    outputs(304) <= layer4_outputs(148);
    outputs(305) <= not(layer4_outputs(721));
    outputs(306) <= layer4_outputs(7677);
    outputs(307) <= not((layer4_outputs(4920)) or (layer4_outputs(3081)));
    outputs(308) <= not(layer4_outputs(6930));
    outputs(309) <= layer4_outputs(1344);
    outputs(310) <= not(layer4_outputs(2717));
    outputs(311) <= (layer4_outputs(2161)) or (layer4_outputs(1161));
    outputs(312) <= (layer4_outputs(5373)) and not (layer4_outputs(4187));
    outputs(313) <= layer4_outputs(2568);
    outputs(314) <= layer4_outputs(4365);
    outputs(315) <= not(layer4_outputs(4218));
    outputs(316) <= layer4_outputs(5579);
    outputs(317) <= layer4_outputs(3293);
    outputs(318) <= not(layer4_outputs(6930));
    outputs(319) <= not(layer4_outputs(1962)) or (layer4_outputs(2279));
    outputs(320) <= layer4_outputs(7567);
    outputs(321) <= not(layer4_outputs(3285));
    outputs(322) <= layer4_outputs(3222);
    outputs(323) <= layer4_outputs(3551);
    outputs(324) <= not(layer4_outputs(5802));
    outputs(325) <= not((layer4_outputs(2164)) xor (layer4_outputs(80)));
    outputs(326) <= layer4_outputs(7199);
    outputs(327) <= layer4_outputs(1952);
    outputs(328) <= layer4_outputs(5342);
    outputs(329) <= not(layer4_outputs(6717));
    outputs(330) <= not((layer4_outputs(1548)) xor (layer4_outputs(2173)));
    outputs(331) <= layer4_outputs(3542);
    outputs(332) <= not((layer4_outputs(614)) and (layer4_outputs(326)));
    outputs(333) <= layer4_outputs(1248);
    outputs(334) <= (layer4_outputs(6456)) and not (layer4_outputs(7311));
    outputs(335) <= (layer4_outputs(139)) xor (layer4_outputs(440));
    outputs(336) <= (layer4_outputs(3724)) or (layer4_outputs(4347));
    outputs(337) <= not(layer4_outputs(6041));
    outputs(338) <= not(layer4_outputs(1492));
    outputs(339) <= not(layer4_outputs(473));
    outputs(340) <= not(layer4_outputs(2382));
    outputs(341) <= not((layer4_outputs(594)) and (layer4_outputs(4362)));
    outputs(342) <= layer4_outputs(3415);
    outputs(343) <= not((layer4_outputs(1546)) xor (layer4_outputs(7043)));
    outputs(344) <= (layer4_outputs(0)) xor (layer4_outputs(2151));
    outputs(345) <= (layer4_outputs(2090)) xor (layer4_outputs(4507));
    outputs(346) <= layer4_outputs(3522);
    outputs(347) <= (layer4_outputs(265)) xor (layer4_outputs(6131));
    outputs(348) <= not(layer4_outputs(290));
    outputs(349) <= layer4_outputs(3787);
    outputs(350) <= layer4_outputs(5154);
    outputs(351) <= (layer4_outputs(3452)) and (layer4_outputs(6731));
    outputs(352) <= not(layer4_outputs(4808));
    outputs(353) <= layer4_outputs(954);
    outputs(354) <= not((layer4_outputs(142)) or (layer4_outputs(6326)));
    outputs(355) <= layer4_outputs(6791);
    outputs(356) <= layer4_outputs(5836);
    outputs(357) <= not((layer4_outputs(1519)) xor (layer4_outputs(6997)));
    outputs(358) <= not(layer4_outputs(4985));
    outputs(359) <= layer4_outputs(2749);
    outputs(360) <= not(layer4_outputs(6908));
    outputs(361) <= (layer4_outputs(6828)) and (layer4_outputs(5264));
    outputs(362) <= layer4_outputs(7284);
    outputs(363) <= layer4_outputs(1795);
    outputs(364) <= not(layer4_outputs(6998));
    outputs(365) <= (layer4_outputs(2713)) or (layer4_outputs(1884));
    outputs(366) <= layer4_outputs(2299);
    outputs(367) <= not(layer4_outputs(5923)) or (layer4_outputs(2869));
    outputs(368) <= not(layer4_outputs(1078));
    outputs(369) <= (layer4_outputs(382)) and not (layer4_outputs(3665));
    outputs(370) <= not(layer4_outputs(5948));
    outputs(371) <= (layer4_outputs(7470)) and (layer4_outputs(6990));
    outputs(372) <= not((layer4_outputs(7426)) or (layer4_outputs(2887)));
    outputs(373) <= (layer4_outputs(1470)) and not (layer4_outputs(7263));
    outputs(374) <= (layer4_outputs(6231)) xor (layer4_outputs(2074));
    outputs(375) <= layer4_outputs(3954);
    outputs(376) <= not(layer4_outputs(2138));
    outputs(377) <= layer4_outputs(5826);
    outputs(378) <= not(layer4_outputs(6387));
    outputs(379) <= layer4_outputs(5170);
    outputs(380) <= not(layer4_outputs(7420));
    outputs(381) <= layer4_outputs(7663);
    outputs(382) <= not(layer4_outputs(6630)) or (layer4_outputs(1233));
    outputs(383) <= (layer4_outputs(5612)) xor (layer4_outputs(5638));
    outputs(384) <= (layer4_outputs(6418)) xor (layer4_outputs(2343));
    outputs(385) <= not((layer4_outputs(4234)) xor (layer4_outputs(5854)));
    outputs(386) <= layer4_outputs(2534);
    outputs(387) <= not(layer4_outputs(2320));
    outputs(388) <= not(layer4_outputs(3121));
    outputs(389) <= not((layer4_outputs(7552)) xor (layer4_outputs(2059)));
    outputs(390) <= layer4_outputs(77);
    outputs(391) <= layer4_outputs(7629);
    outputs(392) <= not(layer4_outputs(3294));
    outputs(393) <= layer4_outputs(2126);
    outputs(394) <= layer4_outputs(2469);
    outputs(395) <= (layer4_outputs(3197)) xor (layer4_outputs(1132));
    outputs(396) <= not(layer4_outputs(6611));
    outputs(397) <= not(layer4_outputs(6491));
    outputs(398) <= (layer4_outputs(1373)) xor (layer4_outputs(2207));
    outputs(399) <= layer4_outputs(2355);
    outputs(400) <= (layer4_outputs(3380)) or (layer4_outputs(314));
    outputs(401) <= (layer4_outputs(7349)) and not (layer4_outputs(971));
    outputs(402) <= not((layer4_outputs(4175)) or (layer4_outputs(1203)));
    outputs(403) <= layer4_outputs(847);
    outputs(404) <= (layer4_outputs(1561)) xor (layer4_outputs(4331));
    outputs(405) <= not((layer4_outputs(7382)) or (layer4_outputs(4223)));
    outputs(406) <= not(layer4_outputs(3243));
    outputs(407) <= layer4_outputs(3208);
    outputs(408) <= not(layer4_outputs(1726));
    outputs(409) <= not(layer4_outputs(5626));
    outputs(410) <= not((layer4_outputs(713)) xor (layer4_outputs(6823)));
    outputs(411) <= not(layer4_outputs(5967));
    outputs(412) <= not(layer4_outputs(1284));
    outputs(413) <= layer4_outputs(3227);
    outputs(414) <= (layer4_outputs(1818)) and not (layer4_outputs(324));
    outputs(415) <= not((layer4_outputs(7369)) xor (layer4_outputs(6593)));
    outputs(416) <= (layer4_outputs(5187)) or (layer4_outputs(3174));
    outputs(417) <= (layer4_outputs(1116)) xor (layer4_outputs(5031));
    outputs(418) <= not(layer4_outputs(2460));
    outputs(419) <= not(layer4_outputs(4562));
    outputs(420) <= (layer4_outputs(4526)) xor (layer4_outputs(5213));
    outputs(421) <= layer4_outputs(4356);
    outputs(422) <= layer4_outputs(4593);
    outputs(423) <= layer4_outputs(173);
    outputs(424) <= (layer4_outputs(5689)) and not (layer4_outputs(1380));
    outputs(425) <= not((layer4_outputs(4037)) xor (layer4_outputs(914)));
    outputs(426) <= (layer4_outputs(169)) and not (layer4_outputs(2545));
    outputs(427) <= (layer4_outputs(2615)) xor (layer4_outputs(6741));
    outputs(428) <= not(layer4_outputs(4892));
    outputs(429) <= not((layer4_outputs(3485)) or (layer4_outputs(5923)));
    outputs(430) <= not(layer4_outputs(2471));
    outputs(431) <= layer4_outputs(2667);
    outputs(432) <= layer4_outputs(928);
    outputs(433) <= not((layer4_outputs(1715)) xor (layer4_outputs(4522)));
    outputs(434) <= not((layer4_outputs(7215)) or (layer4_outputs(7314)));
    outputs(435) <= (layer4_outputs(6024)) and not (layer4_outputs(2553));
    outputs(436) <= not(layer4_outputs(6503));
    outputs(437) <= not(layer4_outputs(456));
    outputs(438) <= not((layer4_outputs(6299)) or (layer4_outputs(556)));
    outputs(439) <= not(layer4_outputs(3562));
    outputs(440) <= not((layer4_outputs(2156)) xor (layer4_outputs(5055)));
    outputs(441) <= not((layer4_outputs(3922)) xor (layer4_outputs(1372)));
    outputs(442) <= not((layer4_outputs(3131)) and (layer4_outputs(6409)));
    outputs(443) <= (layer4_outputs(3539)) xor (layer4_outputs(5750));
    outputs(444) <= not(layer4_outputs(6598));
    outputs(445) <= (layer4_outputs(1843)) or (layer4_outputs(6815));
    outputs(446) <= layer4_outputs(3049);
    outputs(447) <= not(layer4_outputs(1346));
    outputs(448) <= not(layer4_outputs(6702));
    outputs(449) <= not(layer4_outputs(944));
    outputs(450) <= not(layer4_outputs(1097));
    outputs(451) <= not(layer4_outputs(7064));
    outputs(452) <= layer4_outputs(1403);
    outputs(453) <= layer4_outputs(5773);
    outputs(454) <= not(layer4_outputs(6492));
    outputs(455) <= (layer4_outputs(2594)) xor (layer4_outputs(4257));
    outputs(456) <= (layer4_outputs(4674)) and not (layer4_outputs(461));
    outputs(457) <= layer4_outputs(5363);
    outputs(458) <= not(layer4_outputs(4029));
    outputs(459) <= not((layer4_outputs(781)) xor (layer4_outputs(6987)));
    outputs(460) <= not((layer4_outputs(5007)) and (layer4_outputs(2979)));
    outputs(461) <= layer4_outputs(1509);
    outputs(462) <= layer4_outputs(1585);
    outputs(463) <= layer4_outputs(7301);
    outputs(464) <= not(layer4_outputs(7354)) or (layer4_outputs(7472));
    outputs(465) <= not(layer4_outputs(6122));
    outputs(466) <= (layer4_outputs(437)) and not (layer4_outputs(5236));
    outputs(467) <= not(layer4_outputs(157));
    outputs(468) <= not(layer4_outputs(3462));
    outputs(469) <= not(layer4_outputs(4216));
    outputs(470) <= not(layer4_outputs(856));
    outputs(471) <= layer4_outputs(3238);
    outputs(472) <= not(layer4_outputs(1476));
    outputs(473) <= not(layer4_outputs(6254));
    outputs(474) <= layer4_outputs(2577);
    outputs(475) <= not(layer4_outputs(4027));
    outputs(476) <= (layer4_outputs(2482)) or (layer4_outputs(7295));
    outputs(477) <= not(layer4_outputs(1960));
    outputs(478) <= not(layer4_outputs(6030));
    outputs(479) <= not((layer4_outputs(5698)) and (layer4_outputs(1962)));
    outputs(480) <= (layer4_outputs(1585)) and (layer4_outputs(1458));
    outputs(481) <= not((layer4_outputs(4692)) xor (layer4_outputs(2902)));
    outputs(482) <= not((layer4_outputs(5901)) or (layer4_outputs(4929)));
    outputs(483) <= not(layer4_outputs(7276));
    outputs(484) <= not(layer4_outputs(5415));
    outputs(485) <= not((layer4_outputs(1975)) xor (layer4_outputs(4023)));
    outputs(486) <= (layer4_outputs(3733)) and not (layer4_outputs(5571));
    outputs(487) <= not(layer4_outputs(1202));
    outputs(488) <= (layer4_outputs(4086)) xor (layer4_outputs(2070));
    outputs(489) <= not((layer4_outputs(4703)) xor (layer4_outputs(2514)));
    outputs(490) <= not(layer4_outputs(5183));
    outputs(491) <= not(layer4_outputs(1234));
    outputs(492) <= layer4_outputs(6012);
    outputs(493) <= not(layer4_outputs(1681));
    outputs(494) <= not(layer4_outputs(6));
    outputs(495) <= layer4_outputs(5071);
    outputs(496) <= not((layer4_outputs(347)) xor (layer4_outputs(6201)));
    outputs(497) <= layer4_outputs(6417);
    outputs(498) <= layer4_outputs(308);
    outputs(499) <= not(layer4_outputs(4448));
    outputs(500) <= layer4_outputs(5942);
    outputs(501) <= not(layer4_outputs(7032));
    outputs(502) <= not(layer4_outputs(2640));
    outputs(503) <= not((layer4_outputs(3578)) or (layer4_outputs(327)));
    outputs(504) <= not((layer4_outputs(3632)) xor (layer4_outputs(153)));
    outputs(505) <= not((layer4_outputs(3348)) xor (layer4_outputs(819)));
    outputs(506) <= layer4_outputs(767);
    outputs(507) <= layer4_outputs(6044);
    outputs(508) <= not(layer4_outputs(4374));
    outputs(509) <= not((layer4_outputs(3429)) or (layer4_outputs(681)));
    outputs(510) <= layer4_outputs(5461);
    outputs(511) <= not((layer4_outputs(5944)) xor (layer4_outputs(3283)));
    outputs(512) <= not(layer4_outputs(1448)) or (layer4_outputs(7143));
    outputs(513) <= not(layer4_outputs(1119));
    outputs(514) <= not((layer4_outputs(662)) or (layer4_outputs(6859)));
    outputs(515) <= (layer4_outputs(2389)) and not (layer4_outputs(3242));
    outputs(516) <= layer4_outputs(6119);
    outputs(517) <= not((layer4_outputs(1623)) or (layer4_outputs(2404)));
    outputs(518) <= (layer4_outputs(2402)) and not (layer4_outputs(565));
    outputs(519) <= not(layer4_outputs(1050)) or (layer4_outputs(6416));
    outputs(520) <= layer4_outputs(6646);
    outputs(521) <= not(layer4_outputs(3774));
    outputs(522) <= not(layer4_outputs(685));
    outputs(523) <= (layer4_outputs(1458)) and (layer4_outputs(216));
    outputs(524) <= not((layer4_outputs(1347)) or (layer4_outputs(7628)));
    outputs(525) <= (layer4_outputs(5293)) and not (layer4_outputs(6517));
    outputs(526) <= not(layer4_outputs(184));
    outputs(527) <= not((layer4_outputs(1321)) or (layer4_outputs(5592)));
    outputs(528) <= not(layer4_outputs(3340));
    outputs(529) <= (layer4_outputs(526)) xor (layer4_outputs(4121));
    outputs(530) <= layer4_outputs(2466);
    outputs(531) <= layer4_outputs(4618);
    outputs(532) <= (layer4_outputs(1453)) xor (layer4_outputs(6644));
    outputs(533) <= (layer4_outputs(1098)) xor (layer4_outputs(3535));
    outputs(534) <= not(layer4_outputs(446));
    outputs(535) <= not(layer4_outputs(7222));
    outputs(536) <= layer4_outputs(3317);
    outputs(537) <= not(layer4_outputs(4146));
    outputs(538) <= layer4_outputs(7559);
    outputs(539) <= not((layer4_outputs(3507)) and (layer4_outputs(4351)));
    outputs(540) <= (layer4_outputs(6563)) xor (layer4_outputs(4107));
    outputs(541) <= layer4_outputs(4947);
    outputs(542) <= not((layer4_outputs(112)) or (layer4_outputs(3781)));
    outputs(543) <= layer4_outputs(4769);
    outputs(544) <= (layer4_outputs(1108)) or (layer4_outputs(3066));
    outputs(545) <= not(layer4_outputs(1705));
    outputs(546) <= not(layer4_outputs(4281));
    outputs(547) <= not(layer4_outputs(2640));
    outputs(548) <= not(layer4_outputs(6704));
    outputs(549) <= (layer4_outputs(1196)) and not (layer4_outputs(6926));
    outputs(550) <= not(layer4_outputs(5303));
    outputs(551) <= not(layer4_outputs(6397));
    outputs(552) <= (layer4_outputs(2167)) and (layer4_outputs(6288));
    outputs(553) <= not(layer4_outputs(852));
    outputs(554) <= (layer4_outputs(3706)) xor (layer4_outputs(1861));
    outputs(555) <= (layer4_outputs(6462)) and (layer4_outputs(4873));
    outputs(556) <= (layer4_outputs(1051)) or (layer4_outputs(5674));
    outputs(557) <= layer4_outputs(7356);
    outputs(558) <= layer4_outputs(5511);
    outputs(559) <= not(layer4_outputs(4990));
    outputs(560) <= layer4_outputs(232);
    outputs(561) <= not(layer4_outputs(5030));
    outputs(562) <= not((layer4_outputs(5320)) xor (layer4_outputs(6676)));
    outputs(563) <= not((layer4_outputs(1059)) xor (layer4_outputs(6380)));
    outputs(564) <= not(layer4_outputs(5303));
    outputs(565) <= not(layer4_outputs(3219));
    outputs(566) <= layer4_outputs(6971);
    outputs(567) <= not(layer4_outputs(7442));
    outputs(568) <= layer4_outputs(1802);
    outputs(569) <= (layer4_outputs(1927)) and not (layer4_outputs(7051));
    outputs(570) <= layer4_outputs(2950);
    outputs(571) <= not(layer4_outputs(4551));
    outputs(572) <= (layer4_outputs(2257)) xor (layer4_outputs(5411));
    outputs(573) <= not(layer4_outputs(4160));
    outputs(574) <= (layer4_outputs(3618)) and (layer4_outputs(5590));
    outputs(575) <= layer4_outputs(3587);
    outputs(576) <= not((layer4_outputs(2588)) xor (layer4_outputs(6127)));
    outputs(577) <= not(layer4_outputs(17));
    outputs(578) <= not(layer4_outputs(2337));
    outputs(579) <= layer4_outputs(3970);
    outputs(580) <= layer4_outputs(3434);
    outputs(581) <= not(layer4_outputs(3158));
    outputs(582) <= (layer4_outputs(2641)) xor (layer4_outputs(5885));
    outputs(583) <= layer4_outputs(5468);
    outputs(584) <= layer4_outputs(7636);
    outputs(585) <= layer4_outputs(2910);
    outputs(586) <= (layer4_outputs(1376)) xor (layer4_outputs(646));
    outputs(587) <= not(layer4_outputs(6226));
    outputs(588) <= layer4_outputs(3293);
    outputs(589) <= layer4_outputs(5936);
    outputs(590) <= layer4_outputs(5135);
    outputs(591) <= layer4_outputs(353);
    outputs(592) <= not((layer4_outputs(6129)) xor (layer4_outputs(3338)));
    outputs(593) <= (layer4_outputs(5756)) xor (layer4_outputs(966));
    outputs(594) <= (layer4_outputs(383)) and not (layer4_outputs(4301));
    outputs(595) <= not((layer4_outputs(4107)) or (layer4_outputs(1628)));
    outputs(596) <= not(layer4_outputs(4851)) or (layer4_outputs(2143));
    outputs(597) <= not(layer4_outputs(5575));
    outputs(598) <= not((layer4_outputs(5805)) xor (layer4_outputs(6167)));
    outputs(599) <= not(layer4_outputs(6503));
    outputs(600) <= not(layer4_outputs(162));
    outputs(601) <= layer4_outputs(4070);
    outputs(602) <= not(layer4_outputs(7482));
    outputs(603) <= layer4_outputs(6992);
    outputs(604) <= layer4_outputs(6027);
    outputs(605) <= (layer4_outputs(3105)) and (layer4_outputs(2755));
    outputs(606) <= layer4_outputs(4971);
    outputs(607) <= (layer4_outputs(7408)) xor (layer4_outputs(1990));
    outputs(608) <= layer4_outputs(722);
    outputs(609) <= (layer4_outputs(790)) and not (layer4_outputs(1169));
    outputs(610) <= (layer4_outputs(1895)) xor (layer4_outputs(5536));
    outputs(611) <= not((layer4_outputs(6106)) xor (layer4_outputs(1822)));
    outputs(612) <= not((layer4_outputs(6801)) xor (layer4_outputs(3684)));
    outputs(613) <= not(layer4_outputs(5322));
    outputs(614) <= not((layer4_outputs(1077)) xor (layer4_outputs(803)));
    outputs(615) <= layer4_outputs(922);
    outputs(616) <= (layer4_outputs(6849)) xor (layer4_outputs(1410));
    outputs(617) <= (layer4_outputs(3923)) xor (layer4_outputs(5024));
    outputs(618) <= not((layer4_outputs(1260)) xor (layer4_outputs(5104)));
    outputs(619) <= not((layer4_outputs(5027)) and (layer4_outputs(2093)));
    outputs(620) <= not(layer4_outputs(5987));
    outputs(621) <= layer4_outputs(740);
    outputs(622) <= layer4_outputs(2121);
    outputs(623) <= layer4_outputs(3134);
    outputs(624) <= (layer4_outputs(7233)) and (layer4_outputs(1637));
    outputs(625) <= layer4_outputs(220);
    outputs(626) <= (layer4_outputs(4017)) xor (layer4_outputs(3995));
    outputs(627) <= not((layer4_outputs(5416)) or (layer4_outputs(1418)));
    outputs(628) <= not((layer4_outputs(4950)) and (layer4_outputs(4538)));
    outputs(629) <= not((layer4_outputs(4894)) xor (layer4_outputs(6537)));
    outputs(630) <= layer4_outputs(2563);
    outputs(631) <= (layer4_outputs(3192)) and not (layer4_outputs(4082));
    outputs(632) <= (layer4_outputs(6290)) and not (layer4_outputs(3579));
    outputs(633) <= layer4_outputs(7197);
    outputs(634) <= not(layer4_outputs(5332)) or (layer4_outputs(1076));
    outputs(635) <= not(layer4_outputs(586));
    outputs(636) <= (layer4_outputs(1910)) xor (layer4_outputs(4263));
    outputs(637) <= layer4_outputs(2397);
    outputs(638) <= not(layer4_outputs(1198));
    outputs(639) <= not(layer4_outputs(2329));
    outputs(640) <= not((layer4_outputs(552)) xor (layer4_outputs(6870)));
    outputs(641) <= not(layer4_outputs(1807));
    outputs(642) <= not(layer4_outputs(7042));
    outputs(643) <= layer4_outputs(1827);
    outputs(644) <= layer4_outputs(2891);
    outputs(645) <= not(layer4_outputs(7053));
    outputs(646) <= layer4_outputs(15);
    outputs(647) <= not((layer4_outputs(6355)) xor (layer4_outputs(7000)));
    outputs(648) <= (layer4_outputs(1808)) xor (layer4_outputs(3993));
    outputs(649) <= (layer4_outputs(3522)) and not (layer4_outputs(4604));
    outputs(650) <= not((layer4_outputs(6890)) xor (layer4_outputs(3937)));
    outputs(651) <= layer4_outputs(7485);
    outputs(652) <= not((layer4_outputs(1875)) or (layer4_outputs(2619)));
    outputs(653) <= layer4_outputs(7171);
    outputs(654) <= layer4_outputs(3107);
    outputs(655) <= not(layer4_outputs(5849));
    outputs(656) <= (layer4_outputs(4319)) and not (layer4_outputs(7123));
    outputs(657) <= layer4_outputs(3635);
    outputs(658) <= (layer4_outputs(7409)) and not (layer4_outputs(1949));
    outputs(659) <= not((layer4_outputs(5055)) xor (layer4_outputs(1279)));
    outputs(660) <= (layer4_outputs(5110)) and not (layer4_outputs(6032));
    outputs(661) <= (layer4_outputs(6112)) xor (layer4_outputs(5641));
    outputs(662) <= not(layer4_outputs(770));
    outputs(663) <= (layer4_outputs(6543)) and (layer4_outputs(3313));
    outputs(664) <= not((layer4_outputs(5941)) or (layer4_outputs(367)));
    outputs(665) <= layer4_outputs(7666);
    outputs(666) <= layer4_outputs(3040);
    outputs(667) <= (layer4_outputs(2163)) and (layer4_outputs(4004));
    outputs(668) <= (layer4_outputs(1693)) and not (layer4_outputs(3267));
    outputs(669) <= not((layer4_outputs(1153)) xor (layer4_outputs(7561)));
    outputs(670) <= not(layer4_outputs(4184));
    outputs(671) <= (layer4_outputs(4429)) and (layer4_outputs(6918));
    outputs(672) <= not(layer4_outputs(6277)) or (layer4_outputs(5486));
    outputs(673) <= not(layer4_outputs(1863));
    outputs(674) <= not(layer4_outputs(3492)) or (layer4_outputs(1136));
    outputs(675) <= (layer4_outputs(2025)) and not (layer4_outputs(4895));
    outputs(676) <= not(layer4_outputs(754)) or (layer4_outputs(6012));
    outputs(677) <= not(layer4_outputs(5733));
    outputs(678) <= (layer4_outputs(2617)) and (layer4_outputs(21));
    outputs(679) <= layer4_outputs(7061);
    outputs(680) <= not(layer4_outputs(7509));
    outputs(681) <= not((layer4_outputs(6491)) or (layer4_outputs(918)));
    outputs(682) <= (layer4_outputs(5866)) xor (layer4_outputs(231));
    outputs(683) <= not(layer4_outputs(5440));
    outputs(684) <= (layer4_outputs(1232)) and not (layer4_outputs(1003));
    outputs(685) <= layer4_outputs(6282);
    outputs(686) <= not((layer4_outputs(1395)) or (layer4_outputs(7309)));
    outputs(687) <= not(layer4_outputs(7298)) or (layer4_outputs(5487));
    outputs(688) <= layer4_outputs(7111);
    outputs(689) <= layer4_outputs(166);
    outputs(690) <= (layer4_outputs(5529)) xor (layer4_outputs(385));
    outputs(691) <= layer4_outputs(4999);
    outputs(692) <= layer4_outputs(414);
    outputs(693) <= not((layer4_outputs(5796)) xor (layer4_outputs(892)));
    outputs(694) <= (layer4_outputs(3312)) xor (layer4_outputs(1201));
    outputs(695) <= (layer4_outputs(2116)) and not (layer4_outputs(4729));
    outputs(696) <= not(layer4_outputs(3768)) or (layer4_outputs(2172));
    outputs(697) <= (layer4_outputs(6098)) and not (layer4_outputs(2405));
    outputs(698) <= not(layer4_outputs(4837));
    outputs(699) <= layer4_outputs(164);
    outputs(700) <= not(layer4_outputs(4598));
    outputs(701) <= layer4_outputs(4079);
    outputs(702) <= not(layer4_outputs(3309));
    outputs(703) <= not(layer4_outputs(5645));
    outputs(704) <= layer4_outputs(5625);
    outputs(705) <= not((layer4_outputs(1060)) xor (layer4_outputs(1779)));
    outputs(706) <= not((layer4_outputs(7396)) xor (layer4_outputs(3397)));
    outputs(707) <= not(layer4_outputs(6076));
    outputs(708) <= (layer4_outputs(1554)) and (layer4_outputs(2417));
    outputs(709) <= layer4_outputs(4024);
    outputs(710) <= layer4_outputs(1542);
    outputs(711) <= not(layer4_outputs(4632));
    outputs(712) <= layer4_outputs(3633);
    outputs(713) <= not((layer4_outputs(3690)) or (layer4_outputs(2616)));
    outputs(714) <= not(layer4_outputs(1058));
    outputs(715) <= layer4_outputs(2530);
    outputs(716) <= not(layer4_outputs(3990));
    outputs(717) <= not(layer4_outputs(4749));
    outputs(718) <= not(layer4_outputs(7660));
    outputs(719) <= layer4_outputs(2538);
    outputs(720) <= layer4_outputs(3837);
    outputs(721) <= not(layer4_outputs(5759));
    outputs(722) <= (layer4_outputs(7257)) xor (layer4_outputs(5917));
    outputs(723) <= not(layer4_outputs(1495));
    outputs(724) <= layer4_outputs(2020);
    outputs(725) <= (layer4_outputs(7235)) xor (layer4_outputs(4519));
    outputs(726) <= not((layer4_outputs(4564)) or (layer4_outputs(3933)));
    outputs(727) <= not(layer4_outputs(3838));
    outputs(728) <= not(layer4_outputs(1966));
    outputs(729) <= not(layer4_outputs(938));
    outputs(730) <= layer4_outputs(1638);
    outputs(731) <= layer4_outputs(3087);
    outputs(732) <= (layer4_outputs(5485)) xor (layer4_outputs(3431));
    outputs(733) <= layer4_outputs(6894);
    outputs(734) <= not(layer4_outputs(3155));
    outputs(735) <= layer4_outputs(7195);
    outputs(736) <= layer4_outputs(4966);
    outputs(737) <= layer4_outputs(88);
    outputs(738) <= not((layer4_outputs(1900)) or (layer4_outputs(1102)));
    outputs(739) <= not(layer4_outputs(6725));
    outputs(740) <= not((layer4_outputs(3271)) xor (layer4_outputs(5005)));
    outputs(741) <= not(layer4_outputs(1319));
    outputs(742) <= not(layer4_outputs(1168));
    outputs(743) <= not((layer4_outputs(3006)) xor (layer4_outputs(7609)));
    outputs(744) <= not(layer4_outputs(6700));
    outputs(745) <= not(layer4_outputs(1185));
    outputs(746) <= not(layer4_outputs(7420));
    outputs(747) <= layer4_outputs(6126);
    outputs(748) <= (layer4_outputs(6243)) and not (layer4_outputs(5460));
    outputs(749) <= layer4_outputs(5362);
    outputs(750) <= layer4_outputs(6846);
    outputs(751) <= not(layer4_outputs(1750));
    outputs(752) <= (layer4_outputs(5893)) xor (layer4_outputs(5961));
    outputs(753) <= (layer4_outputs(7675)) xor (layer4_outputs(1851));
    outputs(754) <= not(layer4_outputs(1576));
    outputs(755) <= layer4_outputs(203);
    outputs(756) <= not((layer4_outputs(3614)) or (layer4_outputs(3858)));
    outputs(757) <= not(layer4_outputs(6273));
    outputs(758) <= not((layer4_outputs(2179)) xor (layer4_outputs(4387)));
    outputs(759) <= layer4_outputs(525);
    outputs(760) <= layer4_outputs(4943);
    outputs(761) <= not((layer4_outputs(4818)) xor (layer4_outputs(1243)));
    outputs(762) <= (layer4_outputs(5177)) and not (layer4_outputs(2655));
    outputs(763) <= (layer4_outputs(3557)) or (layer4_outputs(1229));
    outputs(764) <= layer4_outputs(9);
    outputs(765) <= not(layer4_outputs(5221));
    outputs(766) <= not((layer4_outputs(4381)) or (layer4_outputs(5024)));
    outputs(767) <= not(layer4_outputs(3232));
    outputs(768) <= '0';
    outputs(769) <= not((layer4_outputs(5003)) or (layer4_outputs(1574)));
    outputs(770) <= (layer4_outputs(1685)) and not (layer4_outputs(1707));
    outputs(771) <= (layer4_outputs(4111)) and (layer4_outputs(6737));
    outputs(772) <= not(layer4_outputs(7169));
    outputs(773) <= layer4_outputs(5216);
    outputs(774) <= not((layer4_outputs(5449)) xor (layer4_outputs(6607)));
    outputs(775) <= layer4_outputs(6266);
    outputs(776) <= layer4_outputs(3155);
    outputs(777) <= layer4_outputs(6437);
    outputs(778) <= layer4_outputs(5931);
    outputs(779) <= (layer4_outputs(1522)) xor (layer4_outputs(7386));
    outputs(780) <= not(layer4_outputs(434)) or (layer4_outputs(740));
    outputs(781) <= layer4_outputs(902);
    outputs(782) <= (layer4_outputs(6863)) and not (layer4_outputs(306));
    outputs(783) <= layer4_outputs(5800);
    outputs(784) <= layer4_outputs(6773);
    outputs(785) <= not((layer4_outputs(1584)) xor (layer4_outputs(5450)));
    outputs(786) <= (layer4_outputs(1397)) and not (layer4_outputs(5378));
    outputs(787) <= (layer4_outputs(336)) and not (layer4_outputs(4124));
    outputs(788) <= layer4_outputs(4465);
    outputs(789) <= layer4_outputs(3901);
    outputs(790) <= not(layer4_outputs(2730));
    outputs(791) <= not(layer4_outputs(3281));
    outputs(792) <= (layer4_outputs(993)) xor (layer4_outputs(6184));
    outputs(793) <= (layer4_outputs(1157)) xor (layer4_outputs(3984));
    outputs(794) <= layer4_outputs(1255);
    outputs(795) <= layer4_outputs(6520);
    outputs(796) <= not((layer4_outputs(1053)) xor (layer4_outputs(2106)));
    outputs(797) <= not(layer4_outputs(2768));
    outputs(798) <= (layer4_outputs(7495)) xor (layer4_outputs(2844));
    outputs(799) <= (layer4_outputs(5772)) xor (layer4_outputs(1081));
    outputs(800) <= (layer4_outputs(53)) and (layer4_outputs(1285));
    outputs(801) <= layer4_outputs(3500);
    outputs(802) <= not(layer4_outputs(6868));
    outputs(803) <= layer4_outputs(389);
    outputs(804) <= (layer4_outputs(204)) and not (layer4_outputs(73));
    outputs(805) <= not(layer4_outputs(4899));
    outputs(806) <= not(layer4_outputs(6014));
    outputs(807) <= not((layer4_outputs(1250)) or (layer4_outputs(2291)));
    outputs(808) <= layer4_outputs(4087);
    outputs(809) <= layer4_outputs(855);
    outputs(810) <= not((layer4_outputs(686)) or (layer4_outputs(2174)));
    outputs(811) <= (layer4_outputs(1033)) and not (layer4_outputs(7418));
    outputs(812) <= (layer4_outputs(6614)) and (layer4_outputs(2886));
    outputs(813) <= (layer4_outputs(2549)) and (layer4_outputs(6755));
    outputs(814) <= not((layer4_outputs(6786)) or (layer4_outputs(7438)));
    outputs(815) <= layer4_outputs(1044);
    outputs(816) <= not(layer4_outputs(1366));
    outputs(817) <= (layer4_outputs(5691)) and (layer4_outputs(1965));
    outputs(818) <= (layer4_outputs(1159)) and (layer4_outputs(954));
    outputs(819) <= (layer4_outputs(5932)) and (layer4_outputs(4644));
    outputs(820) <= not(layer4_outputs(1099));
    outputs(821) <= layer4_outputs(7132);
    outputs(822) <= layer4_outputs(2145);
    outputs(823) <= layer4_outputs(6237);
    outputs(824) <= not(layer4_outputs(6185));
    outputs(825) <= (layer4_outputs(5167)) and not (layer4_outputs(5364));
    outputs(826) <= not(layer4_outputs(5457));
    outputs(827) <= layer4_outputs(3593);
    outputs(828) <= (layer4_outputs(3882)) xor (layer4_outputs(7052));
    outputs(829) <= layer4_outputs(7266);
    outputs(830) <= (layer4_outputs(873)) and not (layer4_outputs(822));
    outputs(831) <= (layer4_outputs(3121)) xor (layer4_outputs(6512));
    outputs(832) <= not(layer4_outputs(4446));
    outputs(833) <= (layer4_outputs(5850)) and not (layer4_outputs(4178));
    outputs(834) <= not((layer4_outputs(5901)) xor (layer4_outputs(86)));
    outputs(835) <= layer4_outputs(7200);
    outputs(836) <= not((layer4_outputs(7394)) xor (layer4_outputs(1840)));
    outputs(837) <= not(layer4_outputs(4792));
    outputs(838) <= layer4_outputs(5948);
    outputs(839) <= layer4_outputs(4470);
    outputs(840) <= not((layer4_outputs(2789)) xor (layer4_outputs(4888)));
    outputs(841) <= (layer4_outputs(656)) and not (layer4_outputs(5347));
    outputs(842) <= not(layer4_outputs(4446));
    outputs(843) <= (layer4_outputs(3556)) and not (layer4_outputs(1972));
    outputs(844) <= (layer4_outputs(3027)) xor (layer4_outputs(7184));
    outputs(845) <= (layer4_outputs(3418)) and (layer4_outputs(5164));
    outputs(846) <= (layer4_outputs(3977)) and not (layer4_outputs(3148));
    outputs(847) <= layer4_outputs(6007);
    outputs(848) <= (layer4_outputs(4208)) and not (layer4_outputs(2898));
    outputs(849) <= (layer4_outputs(7241)) and not (layer4_outputs(6228));
    outputs(850) <= (layer4_outputs(4878)) and not (layer4_outputs(2486));
    outputs(851) <= layer4_outputs(6619);
    outputs(852) <= layer4_outputs(4382);
    outputs(853) <= (layer4_outputs(4796)) and not (layer4_outputs(3936));
    outputs(854) <= not((layer4_outputs(5734)) and (layer4_outputs(910)));
    outputs(855) <= (layer4_outputs(7440)) and not (layer4_outputs(7642));
    outputs(856) <= not(layer4_outputs(5775));
    outputs(857) <= not(layer4_outputs(1353)) or (layer4_outputs(3563));
    outputs(858) <= not(layer4_outputs(3237));
    outputs(859) <= not((layer4_outputs(6445)) or (layer4_outputs(7073)));
    outputs(860) <= not((layer4_outputs(2222)) and (layer4_outputs(6466)));
    outputs(861) <= (layer4_outputs(4637)) and not (layer4_outputs(678));
    outputs(862) <= (layer4_outputs(6633)) and not (layer4_outputs(4783));
    outputs(863) <= not((layer4_outputs(545)) xor (layer4_outputs(769)));
    outputs(864) <= not(layer4_outputs(6289));
    outputs(865) <= not((layer4_outputs(1363)) or (layer4_outputs(108)));
    outputs(866) <= layer4_outputs(5048);
    outputs(867) <= not((layer4_outputs(4335)) xor (layer4_outputs(5176)));
    outputs(868) <= layer4_outputs(7089);
    outputs(869) <= layer4_outputs(7384);
    outputs(870) <= not(layer4_outputs(2554));
    outputs(871) <= not((layer4_outputs(3865)) xor (layer4_outputs(6816)));
    outputs(872) <= (layer4_outputs(1372)) and not (layer4_outputs(3073));
    outputs(873) <= (layer4_outputs(5194)) and (layer4_outputs(5451));
    outputs(874) <= not((layer4_outputs(3159)) or (layer4_outputs(4358)));
    outputs(875) <= (layer4_outputs(7161)) and not (layer4_outputs(69));
    outputs(876) <= layer4_outputs(2201);
    outputs(877) <= (layer4_outputs(1439)) xor (layer4_outputs(6291));
    outputs(878) <= layer4_outputs(7014);
    outputs(879) <= (layer4_outputs(1581)) and (layer4_outputs(1868));
    outputs(880) <= not((layer4_outputs(3755)) or (layer4_outputs(2261)));
    outputs(881) <= layer4_outputs(3649);
    outputs(882) <= layer4_outputs(547);
    outputs(883) <= layer4_outputs(4251);
    outputs(884) <= (layer4_outputs(1789)) and (layer4_outputs(3351));
    outputs(885) <= layer4_outputs(4937);
    outputs(886) <= not(layer4_outputs(7422));
    outputs(887) <= layer4_outputs(3490);
    outputs(888) <= (layer4_outputs(4616)) and not (layer4_outputs(3519));
    outputs(889) <= not(layer4_outputs(2040));
    outputs(890) <= (layer4_outputs(2805)) or (layer4_outputs(6597));
    outputs(891) <= (layer4_outputs(4573)) xor (layer4_outputs(4777));
    outputs(892) <= layer4_outputs(1476);
    outputs(893) <= not((layer4_outputs(2890)) or (layer4_outputs(5414)));
    outputs(894) <= layer4_outputs(1708);
    outputs(895) <= (layer4_outputs(1565)) xor (layer4_outputs(4513));
    outputs(896) <= not(layer4_outputs(542));
    outputs(897) <= layer4_outputs(1904);
    outputs(898) <= layer4_outputs(4291);
    outputs(899) <= layer4_outputs(710);
    outputs(900) <= (layer4_outputs(5615)) and not (layer4_outputs(28));
    outputs(901) <= not((layer4_outputs(7270)) or (layer4_outputs(3660)));
    outputs(902) <= (layer4_outputs(4333)) and not (layer4_outputs(7096));
    outputs(903) <= not((layer4_outputs(7627)) xor (layer4_outputs(6952)));
    outputs(904) <= not((layer4_outputs(1577)) xor (layer4_outputs(2348)));
    outputs(905) <= layer4_outputs(3366);
    outputs(906) <= layer4_outputs(3862);
    outputs(907) <= (layer4_outputs(3581)) xor (layer4_outputs(5969));
    outputs(908) <= not((layer4_outputs(5929)) xor (layer4_outputs(6071)));
    outputs(909) <= (layer4_outputs(1212)) xor (layer4_outputs(4731));
    outputs(910) <= not(layer4_outputs(5337));
    outputs(911) <= not(layer4_outputs(6642));
    outputs(912) <= (layer4_outputs(6900)) and not (layer4_outputs(1444));
    outputs(913) <= (layer4_outputs(539)) and not (layer4_outputs(3564));
    outputs(914) <= not((layer4_outputs(3321)) or (layer4_outputs(1434)));
    outputs(915) <= not((layer4_outputs(6337)) xor (layer4_outputs(839)));
    outputs(916) <= not((layer4_outputs(7370)) xor (layer4_outputs(4270)));
    outputs(917) <= not((layer4_outputs(6457)) xor (layer4_outputs(5488)));
    outputs(918) <= (layer4_outputs(5629)) and not (layer4_outputs(4732));
    outputs(919) <= not((layer4_outputs(2400)) xor (layer4_outputs(2478)));
    outputs(920) <= not((layer4_outputs(4660)) xor (layer4_outputs(1680)));
    outputs(921) <= (layer4_outputs(3333)) or (layer4_outputs(2671));
    outputs(922) <= (layer4_outputs(1328)) and (layer4_outputs(639));
    outputs(923) <= (layer4_outputs(2474)) and not (layer4_outputs(5792));
    outputs(924) <= not(layer4_outputs(3488));
    outputs(925) <= not((layer4_outputs(4512)) or (layer4_outputs(5584)));
    outputs(926) <= (layer4_outputs(882)) xor (layer4_outputs(2667));
    outputs(927) <= not((layer4_outputs(716)) and (layer4_outputs(3742)));
    outputs(928) <= (layer4_outputs(6248)) and not (layer4_outputs(1049));
    outputs(929) <= not(layer4_outputs(3792));
    outputs(930) <= not((layer4_outputs(86)) xor (layer4_outputs(5398)));
    outputs(931) <= (layer4_outputs(1061)) and (layer4_outputs(4566));
    outputs(932) <= not((layer4_outputs(3488)) or (layer4_outputs(3540)));
    outputs(933) <= (layer4_outputs(1345)) xor (layer4_outputs(7306));
    outputs(934) <= layer4_outputs(577);
    outputs(935) <= layer4_outputs(3648);
    outputs(936) <= not(layer4_outputs(6368));
    outputs(937) <= not(layer4_outputs(3545));
    outputs(938) <= not((layer4_outputs(6140)) xor (layer4_outputs(2270)));
    outputs(939) <= not((layer4_outputs(3499)) xor (layer4_outputs(3881)));
    outputs(940) <= (layer4_outputs(2170)) xor (layer4_outputs(7539));
    outputs(941) <= not(layer4_outputs(4689));
    outputs(942) <= not((layer4_outputs(624)) xor (layer4_outputs(2651)));
    outputs(943) <= layer4_outputs(3557);
    outputs(944) <= not((layer4_outputs(1945)) xor (layer4_outputs(3841)));
    outputs(945) <= layer4_outputs(4846);
    outputs(946) <= (layer4_outputs(55)) xor (layer4_outputs(1773));
    outputs(947) <= not(layer4_outputs(5841));
    outputs(948) <= not((layer4_outputs(4539)) or (layer4_outputs(323)));
    outputs(949) <= (layer4_outputs(5943)) xor (layer4_outputs(4285));
    outputs(950) <= layer4_outputs(6434);
    outputs(951) <= not(layer4_outputs(261));
    outputs(952) <= (layer4_outputs(3753)) or (layer4_outputs(4545));
    outputs(953) <= (layer4_outputs(2953)) xor (layer4_outputs(1441));
    outputs(954) <= (layer4_outputs(1571)) xor (layer4_outputs(3422));
    outputs(955) <= not(layer4_outputs(1999));
    outputs(956) <= not(layer4_outputs(1951));
    outputs(957) <= not((layer4_outputs(4355)) xor (layer4_outputs(6615)));
    outputs(958) <= layer4_outputs(2235);
    outputs(959) <= layer4_outputs(2913);
    outputs(960) <= not((layer4_outputs(6004)) and (layer4_outputs(3574)));
    outputs(961) <= (layer4_outputs(6692)) and (layer4_outputs(3616));
    outputs(962) <= layer4_outputs(3647);
    outputs(963) <= layer4_outputs(4945);
    outputs(964) <= not((layer4_outputs(4549)) or (layer4_outputs(2546)));
    outputs(965) <= not(layer4_outputs(3301));
    outputs(966) <= (layer4_outputs(2689)) and not (layer4_outputs(3640));
    outputs(967) <= layer4_outputs(6901);
    outputs(968) <= layer4_outputs(703);
    outputs(969) <= layer4_outputs(2726);
    outputs(970) <= not(layer4_outputs(100));
    outputs(971) <= not(layer4_outputs(7070));
    outputs(972) <= (layer4_outputs(3799)) and not (layer4_outputs(2659));
    outputs(973) <= not(layer4_outputs(965));
    outputs(974) <= layer4_outputs(3586);
    outputs(975) <= not((layer4_outputs(5188)) xor (layer4_outputs(41)));
    outputs(976) <= not((layer4_outputs(3136)) or (layer4_outputs(5622)));
    outputs(977) <= layer4_outputs(4350);
    outputs(978) <= not((layer4_outputs(2206)) or (layer4_outputs(3444)));
    outputs(979) <= (layer4_outputs(1312)) xor (layer4_outputs(5982));
    outputs(980) <= layer4_outputs(7495);
    outputs(981) <= (layer4_outputs(1653)) and not (layer4_outputs(6594));
    outputs(982) <= not(layer4_outputs(4537));
    outputs(983) <= (layer4_outputs(3470)) xor (layer4_outputs(6948));
    outputs(984) <= (layer4_outputs(1176)) and not (layer4_outputs(1616));
    outputs(985) <= not(layer4_outputs(5248));
    outputs(986) <= (layer4_outputs(4140)) and not (layer4_outputs(931));
    outputs(987) <= not(layer4_outputs(7618));
    outputs(988) <= not(layer4_outputs(7652));
    outputs(989) <= not(layer4_outputs(308)) or (layer4_outputs(1721));
    outputs(990) <= not((layer4_outputs(7109)) or (layer4_outputs(2426)));
    outputs(991) <= not(layer4_outputs(938));
    outputs(992) <= not(layer4_outputs(7553));
    outputs(993) <= not(layer4_outputs(5690));
    outputs(994) <= not(layer4_outputs(3424));
    outputs(995) <= layer4_outputs(2648);
    outputs(996) <= not(layer4_outputs(5470));
    outputs(997) <= (layer4_outputs(3427)) and not (layer4_outputs(3804));
    outputs(998) <= (layer4_outputs(5214)) and not (layer4_outputs(7041));
    outputs(999) <= not((layer4_outputs(2185)) xor (layer4_outputs(6460)));
    outputs(1000) <= not(layer4_outputs(968)) or (layer4_outputs(4256));
    outputs(1001) <= not(layer4_outputs(5424));
    outputs(1002) <= not((layer4_outputs(3752)) xor (layer4_outputs(1204)));
    outputs(1003) <= layer4_outputs(4953);
    outputs(1004) <= layer4_outputs(3502);
    outputs(1005) <= not(layer4_outputs(4539));
    outputs(1006) <= layer4_outputs(1497);
    outputs(1007) <= not(layer4_outputs(3135)) or (layer4_outputs(5252));
    outputs(1008) <= not(layer4_outputs(5114));
    outputs(1009) <= layer4_outputs(2816);
    outputs(1010) <= (layer4_outputs(7220)) and not (layer4_outputs(2536));
    outputs(1011) <= not((layer4_outputs(3758)) or (layer4_outputs(5574)));
    outputs(1012) <= not(layer4_outputs(6659));
    outputs(1013) <= not(layer4_outputs(1874));
    outputs(1014) <= (layer4_outputs(6763)) xor (layer4_outputs(1537));
    outputs(1015) <= not(layer4_outputs(1653));
    outputs(1016) <= not((layer4_outputs(6647)) or (layer4_outputs(4695)));
    outputs(1017) <= not((layer4_outputs(6515)) and (layer4_outputs(7403)));
    outputs(1018) <= not(layer4_outputs(814));
    outputs(1019) <= not((layer4_outputs(871)) xor (layer4_outputs(3645)));
    outputs(1020) <= layer4_outputs(2542);
    outputs(1021) <= layer4_outputs(5788);
    outputs(1022) <= not((layer4_outputs(1816)) xor (layer4_outputs(610)));
    outputs(1023) <= (layer4_outputs(5073)) and not (layer4_outputs(2280));
    outputs(1024) <= (layer4_outputs(4800)) and not (layer4_outputs(5521));
    outputs(1025) <= not(layer4_outputs(5376));
    outputs(1026) <= not(layer4_outputs(2357));
    outputs(1027) <= (layer4_outputs(5924)) xor (layer4_outputs(1614));
    outputs(1028) <= (layer4_outputs(5400)) and not (layer4_outputs(7474));
    outputs(1029) <= (layer4_outputs(7489)) and not (layer4_outputs(3543));
    outputs(1030) <= not(layer4_outputs(1270));
    outputs(1031) <= (layer4_outputs(6744)) and (layer4_outputs(2637));
    outputs(1032) <= layer4_outputs(1275);
    outputs(1033) <= (layer4_outputs(6644)) or (layer4_outputs(68));
    outputs(1034) <= (layer4_outputs(2018)) and not (layer4_outputs(7002));
    outputs(1035) <= not((layer4_outputs(3709)) xor (layer4_outputs(6848)));
    outputs(1036) <= not(layer4_outputs(4242));
    outputs(1037) <= not(layer4_outputs(4621));
    outputs(1038) <= (layer4_outputs(559)) xor (layer4_outputs(4957));
    outputs(1039) <= not(layer4_outputs(5062));
    outputs(1040) <= not(layer4_outputs(2939));
    outputs(1041) <= layer4_outputs(3474);
    outputs(1042) <= not((layer4_outputs(7444)) xor (layer4_outputs(4098)));
    outputs(1043) <= (layer4_outputs(4547)) and not (layer4_outputs(7008));
    outputs(1044) <= (layer4_outputs(6128)) and (layer4_outputs(4459));
    outputs(1045) <= (layer4_outputs(700)) xor (layer4_outputs(4030));
    outputs(1046) <= (layer4_outputs(1840)) or (layer4_outputs(3665));
    outputs(1047) <= (layer4_outputs(3615)) and not (layer4_outputs(6797));
    outputs(1048) <= layer4_outputs(7313);
    outputs(1049) <= (layer4_outputs(7637)) xor (layer4_outputs(2359));
    outputs(1050) <= not((layer4_outputs(1363)) or (layer4_outputs(5719)));
    outputs(1051) <= (layer4_outputs(1879)) xor (layer4_outputs(2284));
    outputs(1052) <= not(layer4_outputs(3043));
    outputs(1053) <= not((layer4_outputs(4206)) xor (layer4_outputs(6463)));
    outputs(1054) <= (layer4_outputs(7067)) xor (layer4_outputs(2279));
    outputs(1055) <= not(layer4_outputs(4430));
    outputs(1056) <= (layer4_outputs(4544)) and not (layer4_outputs(1009));
    outputs(1057) <= not(layer4_outputs(5599));
    outputs(1058) <= (layer4_outputs(855)) xor (layer4_outputs(6951));
    outputs(1059) <= layer4_outputs(7653);
    outputs(1060) <= not((layer4_outputs(7333)) or (layer4_outputs(6862)));
    outputs(1061) <= (layer4_outputs(3275)) and not (layer4_outputs(3161));
    outputs(1062) <= not(layer4_outputs(5548));
    outputs(1063) <= (layer4_outputs(2225)) and not (layer4_outputs(6241));
    outputs(1064) <= not(layer4_outputs(2340));
    outputs(1065) <= (layer4_outputs(5912)) and (layer4_outputs(6006));
    outputs(1066) <= (layer4_outputs(6857)) and not (layer4_outputs(3199));
    outputs(1067) <= (layer4_outputs(2178)) and not (layer4_outputs(2198));
    outputs(1068) <= not((layer4_outputs(256)) xor (layer4_outputs(4708)));
    outputs(1069) <= (layer4_outputs(2678)) xor (layer4_outputs(3672));
    outputs(1070) <= not((layer4_outputs(2855)) xor (layer4_outputs(7057)));
    outputs(1071) <= (layer4_outputs(5960)) xor (layer4_outputs(5033));
    outputs(1072) <= (layer4_outputs(7248)) xor (layer4_outputs(6734));
    outputs(1073) <= not(layer4_outputs(3783));
    outputs(1074) <= (layer4_outputs(2318)) and not (layer4_outputs(5816));
    outputs(1075) <= layer4_outputs(3912);
    outputs(1076) <= (layer4_outputs(211)) xor (layer4_outputs(747));
    outputs(1077) <= not(layer4_outputs(6496));
    outputs(1078) <= (layer4_outputs(6154)) xor (layer4_outputs(1823));
    outputs(1079) <= not((layer4_outputs(2672)) or (layer4_outputs(1568)));
    outputs(1080) <= layer4_outputs(3032);
    outputs(1081) <= layer4_outputs(5357);
    outputs(1082) <= not(layer4_outputs(111));
    outputs(1083) <= not((layer4_outputs(6068)) or (layer4_outputs(6174)));
    outputs(1084) <= layer4_outputs(4730);
    outputs(1085) <= (layer4_outputs(5896)) xor (layer4_outputs(4894));
    outputs(1086) <= layer4_outputs(1423);
    outputs(1087) <= not(layer4_outputs(2332));
    outputs(1088) <= (layer4_outputs(6569)) and (layer4_outputs(5962));
    outputs(1089) <= not(layer4_outputs(5908));
    outputs(1090) <= not(layer4_outputs(5827));
    outputs(1091) <= (layer4_outputs(5035)) xor (layer4_outputs(4071));
    outputs(1092) <= (layer4_outputs(3543)) xor (layer4_outputs(579));
    outputs(1093) <= (layer4_outputs(3493)) and not (layer4_outputs(6139));
    outputs(1094) <= not((layer4_outputs(3541)) xor (layer4_outputs(2234)));
    outputs(1095) <= not(layer4_outputs(3765));
    outputs(1096) <= (layer4_outputs(1157)) and not (layer4_outputs(224));
    outputs(1097) <= not(layer4_outputs(5567));
    outputs(1098) <= layer4_outputs(4276);
    outputs(1099) <= layer4_outputs(5157);
    outputs(1100) <= not(layer4_outputs(6357));
    outputs(1101) <= (layer4_outputs(4698)) xor (layer4_outputs(4106));
    outputs(1102) <= not((layer4_outputs(3934)) xor (layer4_outputs(3275)));
    outputs(1103) <= not(layer4_outputs(5403));
    outputs(1104) <= layer4_outputs(4444);
    outputs(1105) <= not(layer4_outputs(1905)) or (layer4_outputs(4265));
    outputs(1106) <= (layer4_outputs(4897)) xor (layer4_outputs(2454));
    outputs(1107) <= layer4_outputs(658);
    outputs(1108) <= not(layer4_outputs(4792));
    outputs(1109) <= not(layer4_outputs(4841));
    outputs(1110) <= not(layer4_outputs(3986));
    outputs(1111) <= (layer4_outputs(2485)) xor (layer4_outputs(1177));
    outputs(1112) <= not(layer4_outputs(6428));
    outputs(1113) <= (layer4_outputs(6580)) and not (layer4_outputs(4124));
    outputs(1114) <= not(layer4_outputs(2310));
    outputs(1115) <= not((layer4_outputs(1590)) xor (layer4_outputs(2686)));
    outputs(1116) <= not(layer4_outputs(728));
    outputs(1117) <= not(layer4_outputs(4247));
    outputs(1118) <= not(layer4_outputs(3959));
    outputs(1119) <= layer4_outputs(2619);
    outputs(1120) <= layer4_outputs(2912);
    outputs(1121) <= not((layer4_outputs(2796)) xor (layer4_outputs(3751)));
    outputs(1122) <= (layer4_outputs(532)) xor (layer4_outputs(1709));
    outputs(1123) <= (layer4_outputs(5718)) and (layer4_outputs(5281));
    outputs(1124) <= not(layer4_outputs(5464));
    outputs(1125) <= layer4_outputs(5301);
    outputs(1126) <= (layer4_outputs(7398)) and (layer4_outputs(5884));
    outputs(1127) <= (layer4_outputs(1600)) xor (layer4_outputs(5133));
    outputs(1128) <= not((layer4_outputs(5765)) or (layer4_outputs(3118)));
    outputs(1129) <= layer4_outputs(544);
    outputs(1130) <= (layer4_outputs(6124)) or (layer4_outputs(5926));
    outputs(1131) <= (layer4_outputs(3679)) xor (layer4_outputs(6011));
    outputs(1132) <= not((layer4_outputs(4219)) or (layer4_outputs(2901)));
    outputs(1133) <= not(layer4_outputs(2885));
    outputs(1134) <= not(layer4_outputs(2851));
    outputs(1135) <= not((layer4_outputs(1041)) xor (layer4_outputs(998)));
    outputs(1136) <= (layer4_outputs(3807)) and not (layer4_outputs(5434));
    outputs(1137) <= (layer4_outputs(5949)) and not (layer4_outputs(3066));
    outputs(1138) <= layer4_outputs(7184);
    outputs(1139) <= layer4_outputs(1774);
    outputs(1140) <= layer4_outputs(4231);
    outputs(1141) <= layer4_outputs(7341);
    outputs(1142) <= layer4_outputs(1612);
    outputs(1143) <= not(layer4_outputs(2339));
    outputs(1144) <= not(layer4_outputs(2708));
    outputs(1145) <= not((layer4_outputs(4911)) xor (layer4_outputs(4147)));
    outputs(1146) <= (layer4_outputs(5414)) xor (layer4_outputs(6538));
    outputs(1147) <= not(layer4_outputs(320));
    outputs(1148) <= (layer4_outputs(6344)) and not (layer4_outputs(2771));
    outputs(1149) <= layer4_outputs(6164);
    outputs(1150) <= not(layer4_outputs(5834));
    outputs(1151) <= layer4_outputs(4735);
    outputs(1152) <= layer4_outputs(6736);
    outputs(1153) <= not((layer4_outputs(2739)) xor (layer4_outputs(2699)));
    outputs(1154) <= (layer4_outputs(616)) and not (layer4_outputs(5894));
    outputs(1155) <= (layer4_outputs(2428)) xor (layer4_outputs(3074));
    outputs(1156) <= not((layer4_outputs(2523)) or (layer4_outputs(3336)));
    outputs(1157) <= layer4_outputs(424);
    outputs(1158) <= layer4_outputs(3280);
    outputs(1159) <= layer4_outputs(3773);
    outputs(1160) <= not((layer4_outputs(6425)) and (layer4_outputs(4596)));
    outputs(1161) <= (layer4_outputs(6972)) and (layer4_outputs(2879));
    outputs(1162) <= not((layer4_outputs(5633)) xor (layer4_outputs(6665)));
    outputs(1163) <= (layer4_outputs(5201)) and not (layer4_outputs(1043));
    outputs(1164) <= not((layer4_outputs(1671)) xor (layer4_outputs(5489)));
    outputs(1165) <= layer4_outputs(1620);
    outputs(1166) <= not(layer4_outputs(3373));
    outputs(1167) <= not(layer4_outputs(6727));
    outputs(1168) <= not((layer4_outputs(132)) xor (layer4_outputs(6470)));
    outputs(1169) <= (layer4_outputs(2545)) and not (layer4_outputs(2734));
    outputs(1170) <= (layer4_outputs(1778)) and not (layer4_outputs(6539));
    outputs(1171) <= not(layer4_outputs(1863));
    outputs(1172) <= (layer4_outputs(5249)) and not (layer4_outputs(5573));
    outputs(1173) <= not(layer4_outputs(2953));
    outputs(1174) <= layer4_outputs(4208);
    outputs(1175) <= not(layer4_outputs(3019));
    outputs(1176) <= not(layer4_outputs(1584));
    outputs(1177) <= not((layer4_outputs(4088)) or (layer4_outputs(7101)));
    outputs(1178) <= layer4_outputs(2406);
    outputs(1179) <= (layer4_outputs(2973)) and (layer4_outputs(1612));
    outputs(1180) <= not(layer4_outputs(1375));
    outputs(1181) <= not(layer4_outputs(3297));
    outputs(1182) <= not((layer4_outputs(2451)) xor (layer4_outputs(2566)));
    outputs(1183) <= not((layer4_outputs(915)) xor (layer4_outputs(7550)));
    outputs(1184) <= not((layer4_outputs(1250)) or (layer4_outputs(6960)));
    outputs(1185) <= layer4_outputs(1016);
    outputs(1186) <= not(layer4_outputs(2171));
    outputs(1187) <= not(layer4_outputs(5848)) or (layer4_outputs(3333));
    outputs(1188) <= layer4_outputs(7384);
    outputs(1189) <= layer4_outputs(7110);
    outputs(1190) <= (layer4_outputs(457)) and (layer4_outputs(47));
    outputs(1191) <= layer4_outputs(4809);
    outputs(1192) <= not((layer4_outputs(7650)) or (layer4_outputs(258)));
    outputs(1193) <= layer4_outputs(7132);
    outputs(1194) <= not((layer4_outputs(6136)) xor (layer4_outputs(1249)));
    outputs(1195) <= not(layer4_outputs(5881));
    outputs(1196) <= layer4_outputs(7148);
    outputs(1197) <= not((layer4_outputs(4158)) xor (layer4_outputs(7517)));
    outputs(1198) <= layer4_outputs(32);
    outputs(1199) <= (layer4_outputs(2092)) xor (layer4_outputs(948));
    outputs(1200) <= not(layer4_outputs(965));
    outputs(1201) <= not((layer4_outputs(1561)) or (layer4_outputs(3630)));
    outputs(1202) <= not((layer4_outputs(6185)) or (layer4_outputs(1926)));
    outputs(1203) <= not(layer4_outputs(2935));
    outputs(1204) <= (layer4_outputs(7009)) xor (layer4_outputs(198));
    outputs(1205) <= (layer4_outputs(4694)) xor (layer4_outputs(4308));
    outputs(1206) <= not((layer4_outputs(6646)) xor (layer4_outputs(567)));
    outputs(1207) <= not((layer4_outputs(3219)) xor (layer4_outputs(2730)));
    outputs(1208) <= layer4_outputs(3871);
    outputs(1209) <= not(layer4_outputs(6443));
    outputs(1210) <= not(layer4_outputs(6170));
    outputs(1211) <= not(layer4_outputs(4558));
    outputs(1212) <= layer4_outputs(7347);
    outputs(1213) <= not(layer4_outputs(3795));
    outputs(1214) <= not((layer4_outputs(7188)) xor (layer4_outputs(4775)));
    outputs(1215) <= (layer4_outputs(7367)) or (layer4_outputs(3010));
    outputs(1216) <= not(layer4_outputs(5161));
    outputs(1217) <= layer4_outputs(2524);
    outputs(1218) <= (layer4_outputs(4909)) xor (layer4_outputs(627));
    outputs(1219) <= layer4_outputs(2517);
    outputs(1220) <= layer4_outputs(944);
    outputs(1221) <= layer4_outputs(4984);
    outputs(1222) <= layer4_outputs(2944);
    outputs(1223) <= not(layer4_outputs(2681));
    outputs(1224) <= (layer4_outputs(6950)) xor (layer4_outputs(5580));
    outputs(1225) <= (layer4_outputs(5219)) xor (layer4_outputs(7018));
    outputs(1226) <= layer4_outputs(5977);
    outputs(1227) <= (layer4_outputs(4736)) and not (layer4_outputs(3707));
    outputs(1228) <= (layer4_outputs(7106)) xor (layer4_outputs(474));
    outputs(1229) <= not((layer4_outputs(5795)) or (layer4_outputs(1232)));
    outputs(1230) <= layer4_outputs(3667);
    outputs(1231) <= not(layer4_outputs(2068));
    outputs(1232) <= (layer4_outputs(6302)) and not (layer4_outputs(7193));
    outputs(1233) <= not(layer4_outputs(860)) or (layer4_outputs(2811));
    outputs(1234) <= layer4_outputs(6157);
    outputs(1235) <= layer4_outputs(3123);
    outputs(1236) <= (layer4_outputs(2377)) and (layer4_outputs(1000));
    outputs(1237) <= not((layer4_outputs(2093)) xor (layer4_outputs(7007)));
    outputs(1238) <= not(layer4_outputs(2614));
    outputs(1239) <= not(layer4_outputs(7506));
    outputs(1240) <= not((layer4_outputs(6329)) or (layer4_outputs(4762)));
    outputs(1241) <= not((layer4_outputs(5453)) and (layer4_outputs(4789)));
    outputs(1242) <= not((layer4_outputs(1695)) or (layer4_outputs(4243)));
    outputs(1243) <= (layer4_outputs(984)) and not (layer4_outputs(6785));
    outputs(1244) <= not(layer4_outputs(1693));
    outputs(1245) <= not(layer4_outputs(5777));
    outputs(1246) <= layer4_outputs(3690);
    outputs(1247) <= (layer4_outputs(3597)) and not (layer4_outputs(5245));
    outputs(1248) <= (layer4_outputs(2335)) and (layer4_outputs(5809));
    outputs(1249) <= (layer4_outputs(3178)) and not (layer4_outputs(133));
    outputs(1250) <= (layer4_outputs(3958)) and not (layer4_outputs(3230));
    outputs(1251) <= not((layer4_outputs(524)) xor (layer4_outputs(7673)));
    outputs(1252) <= (layer4_outputs(6300)) xor (layer4_outputs(4251));
    outputs(1253) <= not((layer4_outputs(6183)) or (layer4_outputs(2236)));
    outputs(1254) <= not(layer4_outputs(6062));
    outputs(1255) <= not((layer4_outputs(2218)) or (layer4_outputs(7358)));
    outputs(1256) <= not(layer4_outputs(6289));
    outputs(1257) <= not((layer4_outputs(4443)) or (layer4_outputs(246)));
    outputs(1258) <= (layer4_outputs(3361)) and not (layer4_outputs(2783));
    outputs(1259) <= not(layer4_outputs(5594));
    outputs(1260) <= layer4_outputs(5042);
    outputs(1261) <= not((layer4_outputs(4613)) and (layer4_outputs(4561)));
    outputs(1262) <= layer4_outputs(4875);
    outputs(1263) <= (layer4_outputs(2972)) and not (layer4_outputs(7247));
    outputs(1264) <= (layer4_outputs(3255)) and not (layer4_outputs(4810));
    outputs(1265) <= layer4_outputs(6588);
    outputs(1266) <= (layer4_outputs(5768)) and not (layer4_outputs(146));
    outputs(1267) <= not(layer4_outputs(6255));
    outputs(1268) <= (layer4_outputs(5957)) and not (layer4_outputs(3755));
    outputs(1269) <= not(layer4_outputs(2897));
    outputs(1270) <= layer4_outputs(6354);
    outputs(1271) <= (layer4_outputs(7591)) xor (layer4_outputs(7351));
    outputs(1272) <= layer4_outputs(1920);
    outputs(1273) <= layer4_outputs(4420);
    outputs(1274) <= not(layer4_outputs(3846));
    outputs(1275) <= (layer4_outputs(2196)) and (layer4_outputs(4829));
    outputs(1276) <= not(layer4_outputs(6983));
    outputs(1277) <= not((layer4_outputs(4390)) and (layer4_outputs(7343)));
    outputs(1278) <= not((layer4_outputs(6476)) xor (layer4_outputs(681)));
    outputs(1279) <= layer4_outputs(7059);
    outputs(1280) <= not(layer4_outputs(328));
    outputs(1281) <= not(layer4_outputs(6807));
    outputs(1282) <= not((layer4_outputs(2852)) or (layer4_outputs(5544)));
    outputs(1283) <= (layer4_outputs(4870)) and (layer4_outputs(878));
    outputs(1284) <= layer4_outputs(5034);
    outputs(1285) <= not(layer4_outputs(5384));
    outputs(1286) <= (layer4_outputs(1789)) and (layer4_outputs(1485));
    outputs(1287) <= not((layer4_outputs(421)) xor (layer4_outputs(403)));
    outputs(1288) <= (layer4_outputs(1227)) and not (layer4_outputs(3888));
    outputs(1289) <= (layer4_outputs(4788)) and (layer4_outputs(7213));
    outputs(1290) <= layer4_outputs(2487);
    outputs(1291) <= (layer4_outputs(1)) and not (layer4_outputs(5823));
    outputs(1292) <= not(layer4_outputs(7125));
    outputs(1293) <= layer4_outputs(3060);
    outputs(1294) <= layer4_outputs(483);
    outputs(1295) <= (layer4_outputs(3170)) and (layer4_outputs(7664));
    outputs(1296) <= layer4_outputs(4455);
    outputs(1297) <= (layer4_outputs(7678)) and not (layer4_outputs(6741));
    outputs(1298) <= not((layer4_outputs(2980)) xor (layer4_outputs(3807)));
    outputs(1299) <= (layer4_outputs(3501)) xor (layer4_outputs(6060));
    outputs(1300) <= not(layer4_outputs(6777));
    outputs(1301) <= layer4_outputs(2751);
    outputs(1302) <= layer4_outputs(1991);
    outputs(1303) <= layer4_outputs(5829);
    outputs(1304) <= layer4_outputs(5045);
    outputs(1305) <= not((layer4_outputs(5728)) or (layer4_outputs(5789)));
    outputs(1306) <= layer4_outputs(6586);
    outputs(1307) <= layer4_outputs(6200);
    outputs(1308) <= layer4_outputs(7355);
    outputs(1309) <= (layer4_outputs(1356)) and not (layer4_outputs(1059));
    outputs(1310) <= layer4_outputs(6591);
    outputs(1311) <= layer4_outputs(1617);
    outputs(1312) <= layer4_outputs(1656);
    outputs(1313) <= (layer4_outputs(7004)) xor (layer4_outputs(6855));
    outputs(1314) <= (layer4_outputs(2530)) xor (layer4_outputs(4267));
    outputs(1315) <= layer4_outputs(4467);
    outputs(1316) <= not((layer4_outputs(3251)) xor (layer4_outputs(848)));
    outputs(1317) <= not(layer4_outputs(6885));
    outputs(1318) <= layer4_outputs(2326);
    outputs(1319) <= (layer4_outputs(3075)) and not (layer4_outputs(38));
    outputs(1320) <= not(layer4_outputs(482));
    outputs(1321) <= (layer4_outputs(5482)) and (layer4_outputs(6449));
    outputs(1322) <= not(layer4_outputs(986));
    outputs(1323) <= layer4_outputs(942);
    outputs(1324) <= not(layer4_outputs(2755));
    outputs(1325) <= layer4_outputs(1997);
    outputs(1326) <= (layer4_outputs(1942)) and not (layer4_outputs(1195));
    outputs(1327) <= not(layer4_outputs(3704));
    outputs(1328) <= not(layer4_outputs(1147));
    outputs(1329) <= (layer4_outputs(2621)) xor (layer4_outputs(87));
    outputs(1330) <= (layer4_outputs(5472)) or (layer4_outputs(4725));
    outputs(1331) <= (layer4_outputs(7536)) xor (layer4_outputs(83));
    outputs(1332) <= not((layer4_outputs(5383)) and (layer4_outputs(3782)));
    outputs(1333) <= (layer4_outputs(2862)) and not (layer4_outputs(2257));
    outputs(1334) <= not((layer4_outputs(311)) xor (layer4_outputs(6568)));
    outputs(1335) <= not((layer4_outputs(1635)) xor (layer4_outputs(3429)));
    outputs(1336) <= (layer4_outputs(4217)) and (layer4_outputs(5404));
    outputs(1337) <= (layer4_outputs(3109)) and not (layer4_outputs(5553));
    outputs(1338) <= layer4_outputs(1204);
    outputs(1339) <= not(layer4_outputs(1252));
    outputs(1340) <= (layer4_outputs(1273)) and (layer4_outputs(4380));
    outputs(1341) <= layer4_outputs(4277);
    outputs(1342) <= not(layer4_outputs(7226));
    outputs(1343) <= not(layer4_outputs(1515)) or (layer4_outputs(123));
    outputs(1344) <= (layer4_outputs(500)) and not (layer4_outputs(2786));
    outputs(1345) <= not(layer4_outputs(3220));
    outputs(1346) <= (layer4_outputs(3917)) xor (layer4_outputs(870));
    outputs(1347) <= not(layer4_outputs(6066));
    outputs(1348) <= not(layer4_outputs(3887));
    outputs(1349) <= layer4_outputs(6340);
    outputs(1350) <= not(layer4_outputs(429));
    outputs(1351) <= layer4_outputs(3026);
    outputs(1352) <= not((layer4_outputs(7669)) or (layer4_outputs(6797)));
    outputs(1353) <= not(layer4_outputs(4453));
    outputs(1354) <= not(layer4_outputs(5402));
    outputs(1355) <= layer4_outputs(5148);
    outputs(1356) <= layer4_outputs(4203);
    outputs(1357) <= not(layer4_outputs(3850));
    outputs(1358) <= layer4_outputs(3705);
    outputs(1359) <= layer4_outputs(3812);
    outputs(1360) <= not((layer4_outputs(5527)) xor (layer4_outputs(7002)));
    outputs(1361) <= layer4_outputs(2256);
    outputs(1362) <= not((layer4_outputs(3609)) xor (layer4_outputs(2846)));
    outputs(1363) <= not(layer4_outputs(2905));
    outputs(1364) <= not(layer4_outputs(2958));
    outputs(1365) <= not(layer4_outputs(7655));
    outputs(1366) <= not(layer4_outputs(2724)) or (layer4_outputs(3869));
    outputs(1367) <= layer4_outputs(1467);
    outputs(1368) <= (layer4_outputs(6903)) xor (layer4_outputs(5189));
    outputs(1369) <= layer4_outputs(2569);
    outputs(1370) <= layer4_outputs(5314);
    outputs(1371) <= not(layer4_outputs(6524));
    outputs(1372) <= layer4_outputs(912);
    outputs(1373) <= layer4_outputs(5437);
    outputs(1374) <= not(layer4_outputs(3686));
    outputs(1375) <= not((layer4_outputs(7230)) xor (layer4_outputs(762)));
    outputs(1376) <= (layer4_outputs(6872)) and (layer4_outputs(5381));
    outputs(1377) <= not(layer4_outputs(7146));
    outputs(1378) <= (layer4_outputs(4853)) and not (layer4_outputs(2291));
    outputs(1379) <= not(layer4_outputs(2558)) or (layer4_outputs(4295));
    outputs(1380) <= not(layer4_outputs(3858));
    outputs(1381) <= layer4_outputs(5575);
    outputs(1382) <= (layer4_outputs(7014)) and not (layer4_outputs(1494));
    outputs(1383) <= not(layer4_outputs(3023));
    outputs(1384) <= layer4_outputs(5475);
    outputs(1385) <= (layer4_outputs(3706)) xor (layer4_outputs(2970));
    outputs(1386) <= not(layer4_outputs(3312));
    outputs(1387) <= not(layer4_outputs(3195));
    outputs(1388) <= (layer4_outputs(1409)) xor (layer4_outputs(3999));
    outputs(1389) <= not((layer4_outputs(2379)) xor (layer4_outputs(887)));
    outputs(1390) <= not((layer4_outputs(6709)) or (layer4_outputs(2692)));
    outputs(1391) <= (layer4_outputs(6935)) and not (layer4_outputs(4899));
    outputs(1392) <= not(layer4_outputs(301));
    outputs(1393) <= not((layer4_outputs(5547)) xor (layer4_outputs(6301)));
    outputs(1394) <= (layer4_outputs(3113)) and not (layer4_outputs(102));
    outputs(1395) <= layer4_outputs(5647);
    outputs(1396) <= not((layer4_outputs(2731)) xor (layer4_outputs(5227)));
    outputs(1397) <= layer4_outputs(3132);
    outputs(1398) <= (layer4_outputs(4893)) and not (layer4_outputs(5115));
    outputs(1399) <= (layer4_outputs(3383)) xor (layer4_outputs(6722));
    outputs(1400) <= not(layer4_outputs(6590));
    outputs(1401) <= layer4_outputs(5532);
    outputs(1402) <= not(layer4_outputs(6152));
    outputs(1403) <= layer4_outputs(3384);
    outputs(1404) <= (layer4_outputs(3240)) and (layer4_outputs(5238));
    outputs(1405) <= not((layer4_outputs(6045)) xor (layer4_outputs(678)));
    outputs(1406) <= layer4_outputs(4212);
    outputs(1407) <= (layer4_outputs(3406)) xor (layer4_outputs(5133));
    outputs(1408) <= not(layer4_outputs(2722));
    outputs(1409) <= layer4_outputs(5585);
    outputs(1410) <= not(layer4_outputs(1651));
    outputs(1411) <= layer4_outputs(5275);
    outputs(1412) <= layer4_outputs(5040);
    outputs(1413) <= (layer4_outputs(978)) and (layer4_outputs(3916));
    outputs(1414) <= layer4_outputs(1122);
    outputs(1415) <= layer4_outputs(5138);
    outputs(1416) <= (layer4_outputs(2560)) xor (layer4_outputs(4782));
    outputs(1417) <= layer4_outputs(1984);
    outputs(1418) <= not((layer4_outputs(7497)) xor (layer4_outputs(1796)));
    outputs(1419) <= not(layer4_outputs(5657));
    outputs(1420) <= layer4_outputs(2272);
    outputs(1421) <= (layer4_outputs(2652)) and not (layer4_outputs(2684));
    outputs(1422) <= (layer4_outputs(3224)) and not (layer4_outputs(252));
    outputs(1423) <= not((layer4_outputs(1080)) or (layer4_outputs(6701)));
    outputs(1424) <= not((layer4_outputs(6436)) xor (layer4_outputs(5304)));
    outputs(1425) <= layer4_outputs(6822);
    outputs(1426) <= layer4_outputs(6439);
    outputs(1427) <= (layer4_outputs(6563)) xor (layer4_outputs(5886));
    outputs(1428) <= not(layer4_outputs(7169));
    outputs(1429) <= layer4_outputs(4001);
    outputs(1430) <= layer4_outputs(4870);
    outputs(1431) <= (layer4_outputs(4417)) and (layer4_outputs(3451));
    outputs(1432) <= not(layer4_outputs(6120));
    outputs(1433) <= not((layer4_outputs(4723)) or (layer4_outputs(7025)));
    outputs(1434) <= layer4_outputs(4275);
    outputs(1435) <= (layer4_outputs(7162)) and not (layer4_outputs(3969));
    outputs(1436) <= (layer4_outputs(1732)) xor (layer4_outputs(2458));
    outputs(1437) <= not((layer4_outputs(1615)) xor (layer4_outputs(1508)));
    outputs(1438) <= not((layer4_outputs(3337)) or (layer4_outputs(5170)));
    outputs(1439) <= layer4_outputs(5629);
    outputs(1440) <= not(layer4_outputs(3296));
    outputs(1441) <= (layer4_outputs(152)) and not (layer4_outputs(4926));
    outputs(1442) <= '0';
    outputs(1443) <= not((layer4_outputs(5107)) xor (layer4_outputs(2331)));
    outputs(1444) <= (layer4_outputs(7365)) and not (layer4_outputs(7369));
    outputs(1445) <= layer4_outputs(2076);
    outputs(1446) <= layer4_outputs(1724);
    outputs(1447) <= layer4_outputs(1329);
    outputs(1448) <= (layer4_outputs(3323)) xor (layer4_outputs(2650));
    outputs(1449) <= not(layer4_outputs(2426));
    outputs(1450) <= (layer4_outputs(1400)) and not (layer4_outputs(6350));
    outputs(1451) <= not((layer4_outputs(6057)) xor (layer4_outputs(1607)));
    outputs(1452) <= layer4_outputs(4726);
    outputs(1453) <= not((layer4_outputs(2608)) xor (layer4_outputs(1624)));
    outputs(1454) <= not(layer4_outputs(7047)) or (layer4_outputs(3592));
    outputs(1455) <= not((layer4_outputs(7032)) xor (layer4_outputs(4526)));
    outputs(1456) <= layer4_outputs(5224);
    outputs(1457) <= not((layer4_outputs(6796)) and (layer4_outputs(1408)));
    outputs(1458) <= (layer4_outputs(5665)) and not (layer4_outputs(3937));
    outputs(1459) <= not((layer4_outputs(3269)) or (layer4_outputs(6608)));
    outputs(1460) <= not(layer4_outputs(2010));
    outputs(1461) <= not(layer4_outputs(1126));
    outputs(1462) <= (layer4_outputs(839)) xor (layer4_outputs(1632));
    outputs(1463) <= not((layer4_outputs(2785)) xor (layer4_outputs(7023)));
    outputs(1464) <= not(layer4_outputs(7034));
    outputs(1465) <= layer4_outputs(1725);
    outputs(1466) <= not(layer4_outputs(7274));
    outputs(1467) <= not(layer4_outputs(1479));
    outputs(1468) <= layer4_outputs(5139);
    outputs(1469) <= not(layer4_outputs(2415));
    outputs(1470) <= not((layer4_outputs(430)) or (layer4_outputs(4242)));
    outputs(1471) <= not((layer4_outputs(7055)) xor (layer4_outputs(5516)));
    outputs(1472) <= not(layer4_outputs(1297));
    outputs(1473) <= not(layer4_outputs(3249));
    outputs(1474) <= (layer4_outputs(2440)) xor (layer4_outputs(642));
    outputs(1475) <= not(layer4_outputs(2502));
    outputs(1476) <= not(layer4_outputs(5360));
    outputs(1477) <= layer4_outputs(1131);
    outputs(1478) <= (layer4_outputs(5398)) and (layer4_outputs(5981));
    outputs(1479) <= not((layer4_outputs(1008)) xor (layer4_outputs(3141)));
    outputs(1480) <= layer4_outputs(1083);
    outputs(1481) <= (layer4_outputs(5725)) xor (layer4_outputs(1305));
    outputs(1482) <= not((layer4_outputs(4916)) xor (layer4_outputs(6721)));
    outputs(1483) <= not(layer4_outputs(4207));
    outputs(1484) <= (layer4_outputs(6814)) xor (layer4_outputs(6634));
    outputs(1485) <= not(layer4_outputs(5031)) or (layer4_outputs(2719));
    outputs(1486) <= (layer4_outputs(601)) xor (layer4_outputs(4986));
    outputs(1487) <= not(layer4_outputs(6518));
    outputs(1488) <= layer4_outputs(773);
    outputs(1489) <= not(layer4_outputs(6196));
    outputs(1490) <= not(layer4_outputs(1267));
    outputs(1491) <= not((layer4_outputs(4471)) or (layer4_outputs(6788)));
    outputs(1492) <= not(layer4_outputs(2774)) or (layer4_outputs(5458));
    outputs(1493) <= (layer4_outputs(3928)) and not (layer4_outputs(3931));
    outputs(1494) <= not(layer4_outputs(4731));
    outputs(1495) <= not(layer4_outputs(494)) or (layer4_outputs(339));
    outputs(1496) <= (layer4_outputs(4104)) and not (layer4_outputs(7353));
    outputs(1497) <= not((layer4_outputs(360)) or (layer4_outputs(4739)));
    outputs(1498) <= not((layer4_outputs(907)) or (layer4_outputs(4715)));
    outputs(1499) <= (layer4_outputs(5167)) and not (layer4_outputs(2655));
    outputs(1500) <= (layer4_outputs(5423)) xor (layer4_outputs(11));
    outputs(1501) <= (layer4_outputs(354)) and not (layer4_outputs(4391));
    outputs(1502) <= not(layer4_outputs(4739)) or (layer4_outputs(2926));
    outputs(1503) <= (layer4_outputs(6030)) xor (layer4_outputs(67));
    outputs(1504) <= (layer4_outputs(1094)) and not (layer4_outputs(2967));
    outputs(1505) <= (layer4_outputs(6826)) and (layer4_outputs(5067));
    outputs(1506) <= layer4_outputs(2811);
    outputs(1507) <= not(layer4_outputs(7011));
    outputs(1508) <= layer4_outputs(915);
    outputs(1509) <= layer4_outputs(1563);
    outputs(1510) <= not((layer4_outputs(2846)) xor (layer4_outputs(4058)));
    outputs(1511) <= (layer4_outputs(5517)) xor (layer4_outputs(836));
    outputs(1512) <= not(layer4_outputs(6105));
    outputs(1513) <= (layer4_outputs(1723)) xor (layer4_outputs(2595));
    outputs(1514) <= not(layer4_outputs(4713));
    outputs(1515) <= (layer4_outputs(3498)) xor (layer4_outputs(6853));
    outputs(1516) <= not(layer4_outputs(3220));
    outputs(1517) <= (layer4_outputs(7010)) xor (layer4_outputs(3767));
    outputs(1518) <= (layer4_outputs(1772)) and not (layer4_outputs(1613));
    outputs(1519) <= not(layer4_outputs(2189));
    outputs(1520) <= layer4_outputs(2414);
    outputs(1521) <= (layer4_outputs(4211)) and not (layer4_outputs(5296));
    outputs(1522) <= (layer4_outputs(4826)) xor (layer4_outputs(6970));
    outputs(1523) <= (layer4_outputs(4360)) xor (layer4_outputs(6470));
    outputs(1524) <= (layer4_outputs(370)) and not (layer4_outputs(2666));
    outputs(1525) <= not((layer4_outputs(3471)) or (layer4_outputs(366)));
    outputs(1526) <= not((layer4_outputs(2265)) xor (layer4_outputs(3467)));
    outputs(1527) <= (layer4_outputs(5065)) and not (layer4_outputs(2119));
    outputs(1528) <= not(layer4_outputs(3994));
    outputs(1529) <= layer4_outputs(4781);
    outputs(1530) <= (layer4_outputs(2748)) and not (layer4_outputs(7669));
    outputs(1531) <= (layer4_outputs(4645)) and (layer4_outputs(6178));
    outputs(1532) <= (layer4_outputs(1950)) and (layer4_outputs(1365));
    outputs(1533) <= layer4_outputs(610);
    outputs(1534) <= layer4_outputs(5652);
    outputs(1535) <= not((layer4_outputs(4166)) or (layer4_outputs(3421)));
    outputs(1536) <= not(layer4_outputs(5684));
    outputs(1537) <= not(layer4_outputs(783));
    outputs(1538) <= not(layer4_outputs(2976));
    outputs(1539) <= layer4_outputs(4105);
    outputs(1540) <= not(layer4_outputs(3257));
    outputs(1541) <= (layer4_outputs(5331)) and not (layer4_outputs(6050));
    outputs(1542) <= not(layer4_outputs(6635));
    outputs(1543) <= not(layer4_outputs(7071));
    outputs(1544) <= not(layer4_outputs(4668));
    outputs(1545) <= not(layer4_outputs(3898));
    outputs(1546) <= layer4_outputs(2154);
    outputs(1547) <= not(layer4_outputs(5290));
    outputs(1548) <= layer4_outputs(6951);
    outputs(1549) <= (layer4_outputs(2435)) and not (layer4_outputs(3077));
    outputs(1550) <= not((layer4_outputs(4790)) xor (layer4_outputs(6428)));
    outputs(1551) <= not(layer4_outputs(7578));
    outputs(1552) <= not((layer4_outputs(627)) xor (layer4_outputs(7189)));
    outputs(1553) <= not(layer4_outputs(5760));
    outputs(1554) <= layer4_outputs(7643);
    outputs(1555) <= not(layer4_outputs(4997));
    outputs(1556) <= layer4_outputs(4022);
    outputs(1557) <= not(layer4_outputs(1684));
    outputs(1558) <= not((layer4_outputs(7093)) xor (layer4_outputs(6508)));
    outputs(1559) <= (layer4_outputs(4414)) xor (layer4_outputs(1535));
    outputs(1560) <= layer4_outputs(4612);
    outputs(1561) <= layer4_outputs(4132);
    outputs(1562) <= not(layer4_outputs(439));
    outputs(1563) <= layer4_outputs(243);
    outputs(1564) <= layer4_outputs(7120);
    outputs(1565) <= (layer4_outputs(1545)) and (layer4_outputs(5357));
    outputs(1566) <= layer4_outputs(6687);
    outputs(1567) <= (layer4_outputs(4266)) xor (layer4_outputs(1325));
    outputs(1568) <= layer4_outputs(3303);
    outputs(1569) <= (layer4_outputs(3902)) or (layer4_outputs(3485));
    outputs(1570) <= not(layer4_outputs(6738));
    outputs(1571) <= not((layer4_outputs(7329)) xor (layer4_outputs(5600)));
    outputs(1572) <= (layer4_outputs(5551)) and not (layer4_outputs(6148));
    outputs(1573) <= (layer4_outputs(3128)) and not (layer4_outputs(6070));
    outputs(1574) <= not((layer4_outputs(6656)) xor (layer4_outputs(7630)));
    outputs(1575) <= not(layer4_outputs(3775));
    outputs(1576) <= layer4_outputs(5352);
    outputs(1577) <= layer4_outputs(3167);
    outputs(1578) <= layer4_outputs(6645);
    outputs(1579) <= layer4_outputs(461);
    outputs(1580) <= layer4_outputs(7421);
    outputs(1581) <= not(layer4_outputs(3043));
    outputs(1582) <= layer4_outputs(6485);
    outputs(1583) <= not(layer4_outputs(5000));
    outputs(1584) <= not(layer4_outputs(5188));
    outputs(1585) <= not((layer4_outputs(7142)) xor (layer4_outputs(6276)));
    outputs(1586) <= not(layer4_outputs(3623));
    outputs(1587) <= layer4_outputs(4346);
    outputs(1588) <= (layer4_outputs(4650)) xor (layer4_outputs(1213));
    outputs(1589) <= layer4_outputs(4275);
    outputs(1590) <= not((layer4_outputs(6000)) xor (layer4_outputs(6352)));
    outputs(1591) <= layer4_outputs(5933);
    outputs(1592) <= layer4_outputs(2721);
    outputs(1593) <= not(layer4_outputs(957));
    outputs(1594) <= layer4_outputs(630);
    outputs(1595) <= (layer4_outputs(2873)) xor (layer4_outputs(6352));
    outputs(1596) <= not(layer4_outputs(3572));
    outputs(1597) <= not(layer4_outputs(4761));
    outputs(1598) <= layer4_outputs(3554);
    outputs(1599) <= not(layer4_outputs(2319));
    outputs(1600) <= not(layer4_outputs(5891));
    outputs(1601) <= not((layer4_outputs(4110)) xor (layer4_outputs(6748)));
    outputs(1602) <= (layer4_outputs(2633)) and not (layer4_outputs(2157));
    outputs(1603) <= layer4_outputs(2943);
    outputs(1604) <= not(layer4_outputs(785));
    outputs(1605) <= (layer4_outputs(2276)) xor (layer4_outputs(4295));
    outputs(1606) <= not(layer4_outputs(1278));
    outputs(1607) <= not((layer4_outputs(3812)) or (layer4_outputs(4473)));
    outputs(1608) <= not(layer4_outputs(2097));
    outputs(1609) <= layer4_outputs(1275);
    outputs(1610) <= layer4_outputs(773);
    outputs(1611) <= not(layer4_outputs(6022));
    outputs(1612) <= (layer4_outputs(3961)) xor (layer4_outputs(3114));
    outputs(1613) <= layer4_outputs(2515);
    outputs(1614) <= not(layer4_outputs(995));
    outputs(1615) <= not(layer4_outputs(1864)) or (layer4_outputs(2175));
    outputs(1616) <= layer4_outputs(6659);
    outputs(1617) <= layer4_outputs(362);
    outputs(1618) <= (layer4_outputs(4496)) and (layer4_outputs(1225));
    outputs(1619) <= layer4_outputs(5745);
    outputs(1620) <= not(layer4_outputs(973));
    outputs(1621) <= (layer4_outputs(6382)) xor (layer4_outputs(4099));
    outputs(1622) <= not(layer4_outputs(2968));
    outputs(1623) <= layer4_outputs(1893);
    outputs(1624) <= layer4_outputs(2054);
    outputs(1625) <= layer4_outputs(4820);
    outputs(1626) <= layer4_outputs(3646);
    outputs(1627) <= not(layer4_outputs(6984));
    outputs(1628) <= layer4_outputs(2106);
    outputs(1629) <= not(layer4_outputs(966));
    outputs(1630) <= not(layer4_outputs(3848));
    outputs(1631) <= not(layer4_outputs(1657)) or (layer4_outputs(3363));
    outputs(1632) <= not(layer4_outputs(4163));
    outputs(1633) <= layer4_outputs(3371);
    outputs(1634) <= not(layer4_outputs(7247));
    outputs(1635) <= (layer4_outputs(5262)) xor (layer4_outputs(2860));
    outputs(1636) <= layer4_outputs(5582);
    outputs(1637) <= layer4_outputs(3560);
    outputs(1638) <= layer4_outputs(1105);
    outputs(1639) <= not((layer4_outputs(5568)) and (layer4_outputs(4043)));
    outputs(1640) <= not(layer4_outputs(3264));
    outputs(1641) <= not(layer4_outputs(900)) or (layer4_outputs(7641));
    outputs(1642) <= layer4_outputs(6728);
    outputs(1643) <= (layer4_outputs(2537)) and not (layer4_outputs(3402));
    outputs(1644) <= (layer4_outputs(1570)) or (layer4_outputs(6210));
    outputs(1645) <= layer4_outputs(4423);
    outputs(1646) <= not(layer4_outputs(841));
    outputs(1647) <= not(layer4_outputs(6743));
    outputs(1648) <= (layer4_outputs(7046)) and not (layer4_outputs(3252));
    outputs(1649) <= layer4_outputs(4324);
    outputs(1650) <= not(layer4_outputs(1241));
    outputs(1651) <= not((layer4_outputs(7087)) and (layer4_outputs(2433)));
    outputs(1652) <= layer4_outputs(680);
    outputs(1653) <= not((layer4_outputs(786)) and (layer4_outputs(4668)));
    outputs(1654) <= not(layer4_outputs(5763));
    outputs(1655) <= not((layer4_outputs(7039)) and (layer4_outputs(5006)));
    outputs(1656) <= not(layer4_outputs(4912));
    outputs(1657) <= (layer4_outputs(3457)) and not (layer4_outputs(22));
    outputs(1658) <= not(layer4_outputs(100));
    outputs(1659) <= (layer4_outputs(4369)) and not (layer4_outputs(7187));
    outputs(1660) <= (layer4_outputs(6247)) and not (layer4_outputs(5598));
    outputs(1661) <= layer4_outputs(6513);
    outputs(1662) <= layer4_outputs(789);
    outputs(1663) <= layer4_outputs(4859);
    outputs(1664) <= not(layer4_outputs(5892));
    outputs(1665) <= not(layer4_outputs(2109));
    outputs(1666) <= (layer4_outputs(6325)) and not (layer4_outputs(5875));
    outputs(1667) <= not(layer4_outputs(5771));
    outputs(1668) <= not(layer4_outputs(7173));
    outputs(1669) <= not(layer4_outputs(5784));
    outputs(1670) <= not(layer4_outputs(3524));
    outputs(1671) <= layer4_outputs(6752);
    outputs(1672) <= not(layer4_outputs(3266));
    outputs(1673) <= not(layer4_outputs(6748)) or (layer4_outputs(193));
    outputs(1674) <= not(layer4_outputs(2404));
    outputs(1675) <= not(layer4_outputs(7550));
    outputs(1676) <= (layer4_outputs(364)) and not (layer4_outputs(3514));
    outputs(1677) <= not(layer4_outputs(148));
    outputs(1678) <= layer4_outputs(1688);
    outputs(1679) <= (layer4_outputs(2772)) xor (layer4_outputs(5726));
    outputs(1680) <= not((layer4_outputs(6358)) xor (layer4_outputs(511)));
    outputs(1681) <= layer4_outputs(1815);
    outputs(1682) <= layer4_outputs(119);
    outputs(1683) <= layer4_outputs(2645);
    outputs(1684) <= layer4_outputs(4967);
    outputs(1685) <= layer4_outputs(3003);
    outputs(1686) <= (layer4_outputs(1633)) and not (layer4_outputs(7049));
    outputs(1687) <= not((layer4_outputs(7594)) xor (layer4_outputs(6162)));
    outputs(1688) <= layer4_outputs(6678);
    outputs(1689) <= layer4_outputs(3468);
    outputs(1690) <= layer4_outputs(6724);
    outputs(1691) <= not(layer4_outputs(793));
    outputs(1692) <= not(layer4_outputs(3296)) or (layer4_outputs(6915));
    outputs(1693) <= not(layer4_outputs(5865));
    outputs(1694) <= not(layer4_outputs(5569));
    outputs(1695) <= (layer4_outputs(5219)) or (layer4_outputs(5041));
    outputs(1696) <= layer4_outputs(2704);
    outputs(1697) <= (layer4_outputs(6163)) and (layer4_outputs(563));
    outputs(1698) <= not(layer4_outputs(2894));
    outputs(1699) <= not((layer4_outputs(115)) and (layer4_outputs(575)));
    outputs(1700) <= layer4_outputs(3614);
    outputs(1701) <= layer4_outputs(2164);
    outputs(1702) <= layer4_outputs(7290);
    outputs(1703) <= not(layer4_outputs(752)) or (layer4_outputs(5390));
    outputs(1704) <= layer4_outputs(7424);
    outputs(1705) <= layer4_outputs(2500);
    outputs(1706) <= layer4_outputs(5834);
    outputs(1707) <= not(layer4_outputs(7475)) or (layer4_outputs(2387));
    outputs(1708) <= layer4_outputs(7493);
    outputs(1709) <= layer4_outputs(516);
    outputs(1710) <= not(layer4_outputs(7114));
    outputs(1711) <= not((layer4_outputs(2609)) xor (layer4_outputs(7063)));
    outputs(1712) <= not((layer4_outputs(5869)) and (layer4_outputs(7524)));
    outputs(1713) <= not(layer4_outputs(1901));
    outputs(1714) <= layer4_outputs(4112);
    outputs(1715) <= (layer4_outputs(1456)) xor (layer4_outputs(6413));
    outputs(1716) <= (layer4_outputs(1207)) xor (layer4_outputs(776));
    outputs(1717) <= not((layer4_outputs(6738)) xor (layer4_outputs(3210)));
    outputs(1718) <= not((layer4_outputs(3090)) and (layer4_outputs(3757)));
    outputs(1719) <= not(layer4_outputs(4157));
    outputs(1720) <= layer4_outputs(477);
    outputs(1721) <= (layer4_outputs(619)) and not (layer4_outputs(2845));
    outputs(1722) <= not(layer4_outputs(6871));
    outputs(1723) <= (layer4_outputs(4130)) and not (layer4_outputs(7598));
    outputs(1724) <= not(layer4_outputs(5233));
    outputs(1725) <= not(layer4_outputs(3176));
    outputs(1726) <= (layer4_outputs(6554)) xor (layer4_outputs(821));
    outputs(1727) <= (layer4_outputs(2422)) xor (layer4_outputs(827));
    outputs(1728) <= not((layer4_outputs(4103)) or (layer4_outputs(967)));
    outputs(1729) <= not((layer4_outputs(1511)) xor (layer4_outputs(6825)));
    outputs(1730) <= not(layer4_outputs(6226));
    outputs(1731) <= (layer4_outputs(4654)) xor (layer4_outputs(6239));
    outputs(1732) <= not((layer4_outputs(6046)) and (layer4_outputs(343)));
    outputs(1733) <= layer4_outputs(1970);
    outputs(1734) <= not(layer4_outputs(6190));
    outputs(1735) <= layer4_outputs(1638);
    outputs(1736) <= not(layer4_outputs(4065));
    outputs(1737) <= not(layer4_outputs(2345));
    outputs(1738) <= not(layer4_outputs(1983)) or (layer4_outputs(272));
    outputs(1739) <= (layer4_outputs(2247)) or (layer4_outputs(6784));
    outputs(1740) <= (layer4_outputs(2359)) xor (layer4_outputs(5345));
    outputs(1741) <= layer4_outputs(5542);
    outputs(1742) <= not(layer4_outputs(3358));
    outputs(1743) <= not(layer4_outputs(4222)) or (layer4_outputs(5557));
    outputs(1744) <= layer4_outputs(2490);
    outputs(1745) <= (layer4_outputs(1031)) xor (layer4_outputs(294));
    outputs(1746) <= not(layer4_outputs(5140));
    outputs(1747) <= not((layer4_outputs(704)) or (layer4_outputs(4063)));
    outputs(1748) <= not((layer4_outputs(1932)) or (layer4_outputs(1944)));
    outputs(1749) <= not(layer4_outputs(7126));
    outputs(1750) <= layer4_outputs(4943);
    outputs(1751) <= not(layer4_outputs(2544));
    outputs(1752) <= not((layer4_outputs(4274)) xor (layer4_outputs(535)));
    outputs(1753) <= layer4_outputs(7510);
    outputs(1754) <= (layer4_outputs(85)) xor (layer4_outputs(7223));
    outputs(1755) <= layer4_outputs(818);
    outputs(1756) <= not(layer4_outputs(6113)) or (layer4_outputs(3610));
    outputs(1757) <= layer4_outputs(6565);
    outputs(1758) <= layer4_outputs(4602);
    outputs(1759) <= (layer4_outputs(1411)) and not (layer4_outputs(1418));
    outputs(1760) <= layer4_outputs(4646);
    outputs(1761) <= (layer4_outputs(1723)) xor (layer4_outputs(7242));
    outputs(1762) <= not(layer4_outputs(6688));
    outputs(1763) <= (layer4_outputs(850)) and (layer4_outputs(7334));
    outputs(1764) <= (layer4_outputs(3529)) and not (layer4_outputs(3700));
    outputs(1765) <= not(layer4_outputs(3535));
    outputs(1766) <= not(layer4_outputs(359));
    outputs(1767) <= (layer4_outputs(5111)) and not (layer4_outputs(5454));
    outputs(1768) <= not(layer4_outputs(5934));
    outputs(1769) <= not(layer4_outputs(3752));
    outputs(1770) <= layer4_outputs(4956);
    outputs(1771) <= layer4_outputs(2638);
    outputs(1772) <= not((layer4_outputs(3288)) xor (layer4_outputs(7293)));
    outputs(1773) <= (layer4_outputs(333)) and not (layer4_outputs(734));
    outputs(1774) <= layer4_outputs(6632);
    outputs(1775) <= not(layer4_outputs(5606));
    outputs(1776) <= (layer4_outputs(542)) and not (layer4_outputs(1792));
    outputs(1777) <= not(layer4_outputs(2724));
    outputs(1778) <= layer4_outputs(3138);
    outputs(1779) <= layer4_outputs(668);
    outputs(1780) <= not((layer4_outputs(1362)) xor (layer4_outputs(7576)));
    outputs(1781) <= not(layer4_outputs(1482));
    outputs(1782) <= not(layer4_outputs(3735));
    outputs(1783) <= not((layer4_outputs(4363)) or (layer4_outputs(4458)));
    outputs(1784) <= (layer4_outputs(7040)) and not (layer4_outputs(133));
    outputs(1785) <= layer4_outputs(3253);
    outputs(1786) <= layer4_outputs(1255);
    outputs(1787) <= not(layer4_outputs(3123));
    outputs(1788) <= not((layer4_outputs(5714)) and (layer4_outputs(91)));
    outputs(1789) <= (layer4_outputs(6619)) xor (layer4_outputs(4710));
    outputs(1790) <= not((layer4_outputs(4230)) or (layer4_outputs(1333)));
    outputs(1791) <= not(layer4_outputs(392));
    outputs(1792) <= not((layer4_outputs(6638)) and (layer4_outputs(3701)));
    outputs(1793) <= not(layer4_outputs(1831)) or (layer4_outputs(5230));
    outputs(1794) <= not((layer4_outputs(4972)) or (layer4_outputs(349)));
    outputs(1795) <= layer4_outputs(2014);
    outputs(1796) <= layer4_outputs(6343);
    outputs(1797) <= layer4_outputs(3989);
    outputs(1798) <= (layer4_outputs(2531)) and (layer4_outputs(7060));
    outputs(1799) <= not(layer4_outputs(4778)) or (layer4_outputs(1134));
    outputs(1800) <= not(layer4_outputs(7419));
    outputs(1801) <= not(layer4_outputs(3830));
    outputs(1802) <= layer4_outputs(6632);
    outputs(1803) <= layer4_outputs(6327);
    outputs(1804) <= (layer4_outputs(7517)) and not (layer4_outputs(7613));
    outputs(1805) <= layer4_outputs(7162);
    outputs(1806) <= not(layer4_outputs(4588));
    outputs(1807) <= (layer4_outputs(2284)) and (layer4_outputs(1900));
    outputs(1808) <= layer4_outputs(835);
    outputs(1809) <= not((layer4_outputs(5864)) xor (layer4_outputs(5268)));
    outputs(1810) <= (layer4_outputs(7070)) and (layer4_outputs(5076));
    outputs(1811) <= layer4_outputs(2716);
    outputs(1812) <= not((layer4_outputs(2391)) xor (layer4_outputs(6278)));
    outputs(1813) <= layer4_outputs(5199);
    outputs(1814) <= not(layer4_outputs(1045));
    outputs(1815) <= layer4_outputs(1882);
    outputs(1816) <= (layer4_outputs(4927)) xor (layer4_outputs(3171));
    outputs(1817) <= not(layer4_outputs(6111));
    outputs(1818) <= layer4_outputs(1283);
    outputs(1819) <= (layer4_outputs(2139)) xor (layer4_outputs(1701));
    outputs(1820) <= (layer4_outputs(823)) xor (layer4_outputs(4439));
    outputs(1821) <= not((layer4_outputs(759)) or (layer4_outputs(5023)));
    outputs(1822) <= (layer4_outputs(2531)) and not (layer4_outputs(2147));
    outputs(1823) <= not(layer4_outputs(1195));
    outputs(1824) <= (layer4_outputs(5276)) and (layer4_outputs(2547));
    outputs(1825) <= (layer4_outputs(5604)) and not (layer4_outputs(5212));
    outputs(1826) <= not(layer4_outputs(6341));
    outputs(1827) <= layer4_outputs(645);
    outputs(1828) <= not(layer4_outputs(4278));
    outputs(1829) <= layer4_outputs(732);
    outputs(1830) <= not(layer4_outputs(5195));
    outputs(1831) <= not(layer4_outputs(4977));
    outputs(1832) <= layer4_outputs(655);
    outputs(1833) <= not(layer4_outputs(3338));
    outputs(1834) <= not((layer4_outputs(5973)) xor (layer4_outputs(7113)));
    outputs(1835) <= not(layer4_outputs(5803));
    outputs(1836) <= (layer4_outputs(2190)) xor (layer4_outputs(6196));
    outputs(1837) <= not(layer4_outputs(6592));
    outputs(1838) <= not((layer4_outputs(4950)) xor (layer4_outputs(4361)));
    outputs(1839) <= not(layer4_outputs(1192));
    outputs(1840) <= not((layer4_outputs(6640)) or (layer4_outputs(4933)));
    outputs(1841) <= not(layer4_outputs(4255));
    outputs(1842) <= layer4_outputs(2997);
    outputs(1843) <= not(layer4_outputs(7087)) or (layer4_outputs(293));
    outputs(1844) <= not(layer4_outputs(3825));
    outputs(1845) <= layer4_outputs(6567);
    outputs(1846) <= layer4_outputs(5086);
    outputs(1847) <= not(layer4_outputs(3273));
    outputs(1848) <= not(layer4_outputs(3567));
    outputs(1849) <= not(layer4_outputs(2297));
    outputs(1850) <= layer4_outputs(4082);
    outputs(1851) <= layer4_outputs(2589);
    outputs(1852) <= (layer4_outputs(4224)) xor (layer4_outputs(535));
    outputs(1853) <= (layer4_outputs(2075)) and (layer4_outputs(5297));
    outputs(1854) <= (layer4_outputs(506)) and not (layer4_outputs(4194));
    outputs(1855) <= not(layer4_outputs(2103));
    outputs(1856) <= not((layer4_outputs(5607)) xor (layer4_outputs(3692)));
    outputs(1857) <= layer4_outputs(6280);
    outputs(1858) <= not(layer4_outputs(2288));
    outputs(1859) <= (layer4_outputs(7445)) and not (layer4_outputs(2976));
    outputs(1860) <= layer4_outputs(1394);
    outputs(1861) <= not(layer4_outputs(7506));
    outputs(1862) <= layer4_outputs(2230);
    outputs(1863) <= (layer4_outputs(6469)) and not (layer4_outputs(6540));
    outputs(1864) <= not(layer4_outputs(1141));
    outputs(1865) <= not(layer4_outputs(25));
    outputs(1866) <= (layer4_outputs(969)) and not (layer4_outputs(4145));
    outputs(1867) <= (layer4_outputs(4459)) and (layer4_outputs(5289));
    outputs(1868) <= layer4_outputs(5659);
    outputs(1869) <= layer4_outputs(2386);
    outputs(1870) <= not((layer4_outputs(969)) xor (layer4_outputs(5045)));
    outputs(1871) <= layer4_outputs(3413);
    outputs(1872) <= (layer4_outputs(443)) and (layer4_outputs(5358));
    outputs(1873) <= layer4_outputs(5173);
    outputs(1874) <= not(layer4_outputs(6634));
    outputs(1875) <= (layer4_outputs(1558)) and (layer4_outputs(3570));
    outputs(1876) <= not((layer4_outputs(1630)) and (layer4_outputs(6189)));
    outputs(1877) <= not(layer4_outputs(2));
    outputs(1878) <= not(layer4_outputs(3953));
    outputs(1879) <= layer4_outputs(7647);
    outputs(1880) <= (layer4_outputs(3335)) and not (layer4_outputs(7516));
    outputs(1881) <= not((layer4_outputs(4260)) and (layer4_outputs(3708)));
    outputs(1882) <= not((layer4_outputs(1452)) xor (layer4_outputs(533)));
    outputs(1883) <= (layer4_outputs(1047)) and not (layer4_outputs(2005));
    outputs(1884) <= layer4_outputs(5442);
    outputs(1885) <= (layer4_outputs(4252)) xor (layer4_outputs(6603));
    outputs(1886) <= not(layer4_outputs(5270));
    outputs(1887) <= (layer4_outputs(6714)) and (layer4_outputs(1543));
    outputs(1888) <= (layer4_outputs(1452)) and not (layer4_outputs(817));
    outputs(1889) <= (layer4_outputs(4644)) xor (layer4_outputs(4085));
    outputs(1890) <= layer4_outputs(1125);
    outputs(1891) <= not(layer4_outputs(3620));
    outputs(1892) <= (layer4_outputs(4762)) xor (layer4_outputs(5783));
    outputs(1893) <= not(layer4_outputs(1430)) or (layer4_outputs(2636));
    outputs(1894) <= layer4_outputs(4080);
    outputs(1895) <= not(layer4_outputs(3355));
    outputs(1896) <= layer4_outputs(2900);
    outputs(1897) <= not(layer4_outputs(4904));
    outputs(1898) <= not(layer4_outputs(377));
    outputs(1899) <= (layer4_outputs(32)) xor (layer4_outputs(6274));
    outputs(1900) <= (layer4_outputs(4938)) xor (layer4_outputs(7594));
    outputs(1901) <= not(layer4_outputs(504));
    outputs(1902) <= not((layer4_outputs(6265)) xor (layer4_outputs(5120)));
    outputs(1903) <= not(layer4_outputs(1527));
    outputs(1904) <= layer4_outputs(3938);
    outputs(1905) <= not(layer4_outputs(3785));
    outputs(1906) <= layer4_outputs(2227);
    outputs(1907) <= not((layer4_outputs(5255)) xor (layer4_outputs(5100)));
    outputs(1908) <= not(layer4_outputs(4734));
    outputs(1909) <= layer4_outputs(378);
    outputs(1910) <= not(layer4_outputs(5617)) or (layer4_outputs(4819));
    outputs(1911) <= layer4_outputs(7159);
    outputs(1912) <= not(layer4_outputs(614));
    outputs(1913) <= (layer4_outputs(287)) xor (layer4_outputs(2380));
    outputs(1914) <= (layer4_outputs(3039)) and (layer4_outputs(686));
    outputs(1915) <= layer4_outputs(4913);
    outputs(1916) <= layer4_outputs(1004);
    outputs(1917) <= not(layer4_outputs(2390));
    outputs(1918) <= not(layer4_outputs(7581));
    outputs(1919) <= not((layer4_outputs(7393)) xor (layer4_outputs(4578)));
    outputs(1920) <= layer4_outputs(2597);
    outputs(1921) <= not(layer4_outputs(3933));
    outputs(1922) <= (layer4_outputs(5600)) and not (layer4_outputs(3823));
    outputs(1923) <= layer4_outputs(7673);
    outputs(1924) <= not(layer4_outputs(5619));
    outputs(1925) <= not((layer4_outputs(5946)) or (layer4_outputs(4273)));
    outputs(1926) <= layer4_outputs(1468);
    outputs(1927) <= layer4_outputs(1677);
    outputs(1928) <= (layer4_outputs(7197)) or (layer4_outputs(988));
    outputs(1929) <= not(layer4_outputs(407));
    outputs(1930) <= layer4_outputs(5997);
    outputs(1931) <= (layer4_outputs(5530)) xor (layer4_outputs(1237));
    outputs(1932) <= (layer4_outputs(3802)) xor (layer4_outputs(16));
    outputs(1933) <= not(layer4_outputs(4785));
    outputs(1934) <= (layer4_outputs(6016)) and (layer4_outputs(4776));
    outputs(1935) <= not(layer4_outputs(2038));
    outputs(1936) <= layer4_outputs(333);
    outputs(1937) <= not(layer4_outputs(5686));
    outputs(1938) <= not(layer4_outputs(640)) or (layer4_outputs(182));
    outputs(1939) <= layer4_outputs(1311);
    outputs(1940) <= (layer4_outputs(358)) and (layer4_outputs(7631));
    outputs(1941) <= layer4_outputs(1985);
    outputs(1942) <= not(layer4_outputs(2906));
    outputs(1943) <= layer4_outputs(200);
    outputs(1944) <= (layer4_outputs(7188)) and not (layer4_outputs(4879));
    outputs(1945) <= not(layer4_outputs(3734));
    outputs(1946) <= not(layer4_outputs(6264));
    outputs(1947) <= (layer4_outputs(6296)) xor (layer4_outputs(1449));
    outputs(1948) <= not((layer4_outputs(218)) and (layer4_outputs(3604)));
    outputs(1949) <= not(layer4_outputs(2840));
    outputs(1950) <= not(layer4_outputs(5859));
    outputs(1951) <= not(layer4_outputs(48));
    outputs(1952) <= (layer4_outputs(1049)) xor (layer4_outputs(4136));
    outputs(1953) <= layer4_outputs(6925);
    outputs(1954) <= not(layer4_outputs(2557));
    outputs(1955) <= (layer4_outputs(3823)) xor (layer4_outputs(2959));
    outputs(1956) <= layer4_outputs(2704);
    outputs(1957) <= layer4_outputs(3729);
    outputs(1958) <= layer4_outputs(7275);
    outputs(1959) <= not(layer4_outputs(1505)) or (layer4_outputs(925));
    outputs(1960) <= not(layer4_outputs(2693));
    outputs(1961) <= not(layer4_outputs(6100));
    outputs(1962) <= layer4_outputs(5783);
    outputs(1963) <= layer4_outputs(7624);
    outputs(1964) <= not(layer4_outputs(1381));
    outputs(1965) <= not(layer4_outputs(4940));
    outputs(1966) <= not(layer4_outputs(2992));
    outputs(1967) <= not(layer4_outputs(991));
    outputs(1968) <= not(layer4_outputs(2585));
    outputs(1969) <= (layer4_outputs(212)) and not (layer4_outputs(6680));
    outputs(1970) <= (layer4_outputs(1722)) or (layer4_outputs(2155));
    outputs(1971) <= layer4_outputs(6595);
    outputs(1972) <= not(layer4_outputs(2146));
    outputs(1973) <= layer4_outputs(1326);
    outputs(1974) <= not(layer4_outputs(2146));
    outputs(1975) <= layer4_outputs(2813);
    outputs(1976) <= not(layer4_outputs(3165));
    outputs(1977) <= layer4_outputs(7454);
    outputs(1978) <= layer4_outputs(34);
    outputs(1979) <= (layer4_outputs(2898)) xor (layer4_outputs(6020));
    outputs(1980) <= layer4_outputs(7000);
    outputs(1981) <= not(layer4_outputs(602)) or (layer4_outputs(3935));
    outputs(1982) <= not(layer4_outputs(5952));
    outputs(1983) <= (layer4_outputs(296)) xor (layer4_outputs(4095));
    outputs(1984) <= not(layer4_outputs(5010)) or (layer4_outputs(6401));
    outputs(1985) <= layer4_outputs(2399);
    outputs(1986) <= layer4_outputs(1890);
    outputs(1987) <= layer4_outputs(2399);
    outputs(1988) <= not((layer4_outputs(127)) and (layer4_outputs(6104)));
    outputs(1989) <= not(layer4_outputs(3257));
    outputs(1990) <= (layer4_outputs(6720)) xor (layer4_outputs(3777));
    outputs(1991) <= not((layer4_outputs(5708)) or (layer4_outputs(4565)));
    outputs(1992) <= not(layer4_outputs(2046));
    outputs(1993) <= not(layer4_outputs(2879));
    outputs(1994) <= layer4_outputs(7457);
    outputs(1995) <= not(layer4_outputs(635));
    outputs(1996) <= not(layer4_outputs(7240)) or (layer4_outputs(6272));
    outputs(1997) <= not((layer4_outputs(4868)) and (layer4_outputs(221)));
    outputs(1998) <= (layer4_outputs(5779)) xor (layer4_outputs(4721));
    outputs(1999) <= not(layer4_outputs(3034));
    outputs(2000) <= layer4_outputs(2801);
    outputs(2001) <= layer4_outputs(4094);
    outputs(2002) <= (layer4_outputs(3382)) and not (layer4_outputs(1923));
    outputs(2003) <= layer4_outputs(5387);
    outputs(2004) <= not(layer4_outputs(1907));
    outputs(2005) <= not(layer4_outputs(6236)) or (layer4_outputs(1188));
    outputs(2006) <= layer4_outputs(916);
    outputs(2007) <= not(layer4_outputs(217));
    outputs(2008) <= (layer4_outputs(1462)) xor (layer4_outputs(1222));
    outputs(2009) <= not(layer4_outputs(3872));
    outputs(2010) <= (layer4_outputs(5628)) xor (layer4_outputs(3336));
    outputs(2011) <= layer4_outputs(5835);
    outputs(2012) <= not(layer4_outputs(4741));
    outputs(2013) <= not(layer4_outputs(3433));
    outputs(2014) <= layer4_outputs(4385);
    outputs(2015) <= layer4_outputs(2295);
    outputs(2016) <= layer4_outputs(118);
    outputs(2017) <= layer4_outputs(1160);
    outputs(2018) <= (layer4_outputs(6939)) xor (layer4_outputs(61));
    outputs(2019) <= layer4_outputs(3099);
    outputs(2020) <= layer4_outputs(1724);
    outputs(2021) <= not(layer4_outputs(4940));
    outputs(2022) <= not(layer4_outputs(7149));
    outputs(2023) <= not((layer4_outputs(5630)) or (layer4_outputs(4536)));
    outputs(2024) <= not((layer4_outputs(6581)) xor (layer4_outputs(6545)));
    outputs(2025) <= (layer4_outputs(1504)) xor (layer4_outputs(2905));
    outputs(2026) <= not(layer4_outputs(1197));
    outputs(2027) <= layer4_outputs(7116);
    outputs(2028) <= not(layer4_outputs(3578));
    outputs(2029) <= not(layer4_outputs(5497));
    outputs(2030) <= (layer4_outputs(6385)) and (layer4_outputs(4285));
    outputs(2031) <= layer4_outputs(2694);
    outputs(2032) <= layer4_outputs(1427);
    outputs(2033) <= not(layer4_outputs(4487));
    outputs(2034) <= (layer4_outputs(7568)) xor (layer4_outputs(1760));
    outputs(2035) <= not((layer4_outputs(2995)) or (layer4_outputs(772)));
    outputs(2036) <= (layer4_outputs(7416)) or (layer4_outputs(4763));
    outputs(2037) <= layer4_outputs(3037);
    outputs(2038) <= not(layer4_outputs(3584));
    outputs(2039) <= (layer4_outputs(7313)) xor (layer4_outputs(6146));
    outputs(2040) <= not((layer4_outputs(1793)) and (layer4_outputs(292)));
    outputs(2041) <= not(layer4_outputs(525));
    outputs(2042) <= not((layer4_outputs(4134)) or (layer4_outputs(4457)));
    outputs(2043) <= layer4_outputs(1685);
    outputs(2044) <= not(layer4_outputs(7593)) or (layer4_outputs(2187));
    outputs(2045) <= not(layer4_outputs(2071));
    outputs(2046) <= layer4_outputs(1280);
    outputs(2047) <= not(layer4_outputs(6746));
    outputs(2048) <= layer4_outputs(949);
    outputs(2049) <= not((layer4_outputs(319)) xor (layer4_outputs(195)));
    outputs(2050) <= not((layer4_outputs(1695)) xor (layer4_outputs(5662)));
    outputs(2051) <= not(layer4_outputs(4699));
    outputs(2052) <= not(layer4_outputs(7171));
    outputs(2053) <= layer4_outputs(4999);
    outputs(2054) <= (layer4_outputs(3285)) and not (layer4_outputs(2254));
    outputs(2055) <= not(layer4_outputs(2499)) or (layer4_outputs(898));
    outputs(2056) <= not(layer4_outputs(7062));
    outputs(2057) <= (layer4_outputs(5710)) xor (layer4_outputs(3254));
    outputs(2058) <= layer4_outputs(7521);
    outputs(2059) <= layer4_outputs(3445);
    outputs(2060) <= layer4_outputs(3126);
    outputs(2061) <= layer4_outputs(2525);
    outputs(2062) <= not(layer4_outputs(4364));
    outputs(2063) <= layer4_outputs(75);
    outputs(2064) <= layer4_outputs(2903);
    outputs(2065) <= layer4_outputs(6287);
    outputs(2066) <= not(layer4_outputs(711));
    outputs(2067) <= layer4_outputs(3445);
    outputs(2068) <= (layer4_outputs(5289)) and not (layer4_outputs(2878));
    outputs(2069) <= (layer4_outputs(2452)) xor (layer4_outputs(4709));
    outputs(2070) <= not(layer4_outputs(3574));
    outputs(2071) <= not(layer4_outputs(3455));
    outputs(2072) <= layer4_outputs(4406);
    outputs(2073) <= (layer4_outputs(1276)) or (layer4_outputs(2823));
    outputs(2074) <= (layer4_outputs(620)) xor (layer4_outputs(7334));
    outputs(2075) <= (layer4_outputs(6339)) and not (layer4_outputs(2364));
    outputs(2076) <= (layer4_outputs(2634)) xor (layer4_outputs(4491));
    outputs(2077) <= not((layer4_outputs(7209)) and (layer4_outputs(4621)));
    outputs(2078) <= not(layer4_outputs(3228));
    outputs(2079) <= (layer4_outputs(4597)) and not (layer4_outputs(3012));
    outputs(2080) <= not((layer4_outputs(4248)) xor (layer4_outputs(2793)));
    outputs(2081) <= layer4_outputs(7457);
    outputs(2082) <= not(layer4_outputs(5679)) or (layer4_outputs(737));
    outputs(2083) <= not(layer4_outputs(5254));
    outputs(2084) <= layer4_outputs(274);
    outputs(2085) <= (layer4_outputs(398)) or (layer4_outputs(1072));
    outputs(2086) <= layer4_outputs(5710);
    outputs(2087) <= layer4_outputs(2638);
    outputs(2088) <= not(layer4_outputs(1625));
    outputs(2089) <= not(layer4_outputs(5392));
    outputs(2090) <= (layer4_outputs(2650)) and not (layer4_outputs(137));
    outputs(2091) <= not(layer4_outputs(4364));
    outputs(2092) <= not(layer4_outputs(5515));
    outputs(2093) <= (layer4_outputs(3600)) xor (layer4_outputs(6102));
    outputs(2094) <= not(layer4_outputs(3547));
    outputs(2095) <= not((layer4_outputs(2973)) xor (layer4_outputs(4170)));
    outputs(2096) <= not(layer4_outputs(2503));
    outputs(2097) <= layer4_outputs(1709);
    outputs(2098) <= not(layer4_outputs(3636));
    outputs(2099) <= (layer4_outputs(1174)) xor (layer4_outputs(3353));
    outputs(2100) <= not(layer4_outputs(2981));
    outputs(2101) <= layer4_outputs(455);
    outputs(2102) <= not((layer4_outputs(698)) xor (layer4_outputs(6963)));
    outputs(2103) <= not(layer4_outputs(3359));
    outputs(2104) <= layer4_outputs(3638);
    outputs(2105) <= (layer4_outputs(5404)) xor (layer4_outputs(3368));
    outputs(2106) <= not(layer4_outputs(4867));
    outputs(2107) <= not(layer4_outputs(1897)) or (layer4_outputs(601));
    outputs(2108) <= not(layer4_outputs(2046));
    outputs(2109) <= (layer4_outputs(6431)) xor (layer4_outputs(6673));
    outputs(2110) <= layer4_outputs(2862);
    outputs(2111) <= (layer4_outputs(5634)) and (layer4_outputs(4857));
    outputs(2112) <= not(layer4_outputs(4103));
    outputs(2113) <= not(layer4_outputs(4973));
    outputs(2114) <= layer4_outputs(6931);
    outputs(2115) <= not(layer4_outputs(6834));
    outputs(2116) <= not(layer4_outputs(3370));
    outputs(2117) <= not(layer4_outputs(2338));
    outputs(2118) <= not(layer4_outputs(5323));
    outputs(2119) <= not(layer4_outputs(6390));
    outputs(2120) <= layer4_outputs(1763);
    outputs(2121) <= layer4_outputs(3745);
    outputs(2122) <= not(layer4_outputs(3323));
    outputs(2123) <= layer4_outputs(2745);
    outputs(2124) <= layer4_outputs(3072);
    outputs(2125) <= not(layer4_outputs(2626));
    outputs(2126) <= not((layer4_outputs(4653)) and (layer4_outputs(2554)));
    outputs(2127) <= not(layer4_outputs(5078));
    outputs(2128) <= not(layer4_outputs(1221));
    outputs(2129) <= not(layer4_outputs(6812));
    outputs(2130) <= (layer4_outputs(6845)) and not (layer4_outputs(7501));
    outputs(2131) <= layer4_outputs(2203);
    outputs(2132) <= layer4_outputs(3895);
    outputs(2133) <= layer4_outputs(5786);
    outputs(2134) <= (layer4_outputs(2186)) or (layer4_outputs(3248));
    outputs(2135) <= layer4_outputs(2219);
    outputs(2136) <= layer4_outputs(1688);
    outputs(2137) <= (layer4_outputs(20)) and not (layer4_outputs(4247));
    outputs(2138) <= not((layer4_outputs(2720)) and (layer4_outputs(6610)));
    outputs(2139) <= (layer4_outputs(509)) xor (layer4_outputs(7119));
    outputs(2140) <= layer4_outputs(2078);
    outputs(2141) <= not((layer4_outputs(5975)) xor (layer4_outputs(7531)));
    outputs(2142) <= not((layer4_outputs(5546)) xor (layer4_outputs(3438)));
    outputs(2143) <= not(layer4_outputs(3461)) or (layer4_outputs(5989));
    outputs(2144) <= not(layer4_outputs(5146));
    outputs(2145) <= layer4_outputs(1677);
    outputs(2146) <= layer4_outputs(2154);
    outputs(2147) <= layer4_outputs(1601);
    outputs(2148) <= (layer4_outputs(5123)) xor (layer4_outputs(6031));
    outputs(2149) <= layer4_outputs(1024);
    outputs(2150) <= not(layer4_outputs(7453));
    outputs(2151) <= not(layer4_outputs(1784));
    outputs(2152) <= (layer4_outputs(331)) or (layer4_outputs(2769));
    outputs(2153) <= not(layer4_outputs(1067)) or (layer4_outputs(5156));
    outputs(2154) <= not(layer4_outputs(3246));
    outputs(2155) <= (layer4_outputs(7062)) xor (layer4_outputs(4236));
    outputs(2156) <= not(layer4_outputs(7505));
    outputs(2157) <= layer4_outputs(2743);
    outputs(2158) <= layer4_outputs(4517);
    outputs(2159) <= not(layer4_outputs(1368));
    outputs(2160) <= not((layer4_outputs(380)) or (layer4_outputs(2024)));
    outputs(2161) <= not((layer4_outputs(2302)) xor (layer4_outputs(3712)));
    outputs(2162) <= layer4_outputs(1292);
    outputs(2163) <= layer4_outputs(434);
    outputs(2164) <= not((layer4_outputs(307)) xor (layer4_outputs(1517)));
    outputs(2165) <= not(layer4_outputs(1070));
    outputs(2166) <= not(layer4_outputs(7134));
    outputs(2167) <= (layer4_outputs(2181)) and not (layer4_outputs(481));
    outputs(2168) <= not((layer4_outputs(6058)) xor (layer4_outputs(6393)));
    outputs(2169) <= layer4_outputs(7185);
    outputs(2170) <= layer4_outputs(1525);
    outputs(2171) <= layer4_outputs(238);
    outputs(2172) <= not(layer4_outputs(2032));
    outputs(2173) <= not(layer4_outputs(3034));
    outputs(2174) <= not(layer4_outputs(3502)) or (layer4_outputs(5983));
    outputs(2175) <= layer4_outputs(35);
    outputs(2176) <= not(layer4_outputs(6855)) or (layer4_outputs(3182));
    outputs(2177) <= (layer4_outputs(2073)) or (layer4_outputs(2911));
    outputs(2178) <= not(layer4_outputs(6023)) or (layer4_outputs(3662));
    outputs(2179) <= layer4_outputs(3537);
    outputs(2180) <= (layer4_outputs(6356)) xor (layer4_outputs(706));
    outputs(2181) <= (layer4_outputs(6513)) and (layer4_outputs(3811));
    outputs(2182) <= not(layer4_outputs(3909));
    outputs(2183) <= not(layer4_outputs(7623));
    outputs(2184) <= not(layer4_outputs(1241));
    outputs(2185) <= not(layer4_outputs(3352));
    outputs(2186) <= not((layer4_outputs(7318)) and (layer4_outputs(5493)));
    outputs(2187) <= not(layer4_outputs(2055));
    outputs(2188) <= layer4_outputs(2123);
    outputs(2189) <= (layer4_outputs(7273)) xor (layer4_outputs(2689));
    outputs(2190) <= layer4_outputs(2470);
    outputs(2191) <= layer4_outputs(5358);
    outputs(2192) <= layer4_outputs(4821);
    outputs(2193) <= layer4_outputs(6837);
    outputs(2194) <= (layer4_outputs(1140)) and not (layer4_outputs(2206));
    outputs(2195) <= layer4_outputs(2280);
    outputs(2196) <= (layer4_outputs(3465)) and not (layer4_outputs(772));
    outputs(2197) <= not(layer4_outputs(1975));
    outputs(2198) <= layer4_outputs(1112);
    outputs(2199) <= (layer4_outputs(4211)) and (layer4_outputs(4921));
    outputs(2200) <= not(layer4_outputs(7124));
    outputs(2201) <= layer4_outputs(1140);
    outputs(2202) <= not(layer4_outputs(3048));
    outputs(2203) <= not(layer4_outputs(233));
    outputs(2204) <= layer4_outputs(4905);
    outputs(2205) <= not(layer4_outputs(5736));
    outputs(2206) <= layer4_outputs(4890);
    outputs(2207) <= not(layer4_outputs(5247));
    outputs(2208) <= layer4_outputs(543);
    outputs(2209) <= not(layer4_outputs(3069));
    outputs(2210) <= layer4_outputs(248);
    outputs(2211) <= not(layer4_outputs(3454));
    outputs(2212) <= layer4_outputs(3305);
    outputs(2213) <= (layer4_outputs(4546)) and not (layer4_outputs(302));
    outputs(2214) <= not((layer4_outputs(5374)) xor (layer4_outputs(1431)));
    outputs(2215) <= layer4_outputs(1491);
    outputs(2216) <= layer4_outputs(7288);
    outputs(2217) <= (layer4_outputs(5264)) and (layer4_outputs(2333));
    outputs(2218) <= (layer4_outputs(5535)) xor (layer4_outputs(5177));
    outputs(2219) <= not(layer4_outputs(5285));
    outputs(2220) <= not((layer4_outputs(7193)) xor (layer4_outputs(747)));
    outputs(2221) <= not(layer4_outputs(578)) or (layer4_outputs(700));
    outputs(2222) <= not(layer4_outputs(5818));
    outputs(2223) <= layer4_outputs(357);
    outputs(2224) <= not((layer4_outputs(702)) or (layer4_outputs(2847)));
    outputs(2225) <= not(layer4_outputs(2757));
    outputs(2226) <= (layer4_outputs(4477)) xor (layer4_outputs(4881));
    outputs(2227) <= not(layer4_outputs(7362));
    outputs(2228) <= layer4_outputs(2385);
    outputs(2229) <= not(layer4_outputs(3996)) or (layer4_outputs(5271));
    outputs(2230) <= not(layer4_outputs(4929));
    outputs(2231) <= layer4_outputs(5369);
    outputs(2232) <= layer4_outputs(3748);
    outputs(2233) <= (layer4_outputs(6988)) xor (layer4_outputs(3988));
    outputs(2234) <= not(layer4_outputs(207));
    outputs(2235) <= (layer4_outputs(353)) or (layer4_outputs(3216));
    outputs(2236) <= not((layer4_outputs(7293)) xor (layer4_outputs(6261)));
    outputs(2237) <= not(layer4_outputs(6762));
    outputs(2238) <= not(layer4_outputs(3898));
    outputs(2239) <= not(layer4_outputs(4240));
    outputs(2240) <= layer4_outputs(3646);
    outputs(2241) <= layer4_outputs(2227);
    outputs(2242) <= (layer4_outputs(415)) xor (layer4_outputs(6059));
    outputs(2243) <= (layer4_outputs(4423)) and (layer4_outputs(4343));
    outputs(2244) <= (layer4_outputs(3803)) and not (layer4_outputs(5769));
    outputs(2245) <= (layer4_outputs(3110)) xor (layer4_outputs(4445));
    outputs(2246) <= (layer4_outputs(7262)) and (layer4_outputs(409));
    outputs(2247) <= not(layer4_outputs(49));
    outputs(2248) <= (layer4_outputs(1839)) and not (layer4_outputs(4014));
    outputs(2249) <= layer4_outputs(727);
    outputs(2250) <= layer4_outputs(6408);
    outputs(2251) <= (layer4_outputs(900)) xor (layer4_outputs(1913));
    outputs(2252) <= not(layer4_outputs(6947));
    outputs(2253) <= layer4_outputs(7565);
    outputs(2254) <= layer4_outputs(4553);
    outputs(2255) <= not(layer4_outputs(3701));
    outputs(2256) <= not(layer4_outputs(6223));
    outputs(2257) <= not(layer4_outputs(5823));
    outputs(2258) <= layer4_outputs(438);
    outputs(2259) <= not(layer4_outputs(1644));
    outputs(2260) <= not((layer4_outputs(6716)) xor (layer4_outputs(5052)));
    outputs(2261) <= not(layer4_outputs(2999));
    outputs(2262) <= not(layer4_outputs(5586));
    outputs(2263) <= not(layer4_outputs(3410)) or (layer4_outputs(6678));
    outputs(2264) <= (layer4_outputs(6176)) and not (layer4_outputs(3903));
    outputs(2265) <= (layer4_outputs(7552)) and not (layer4_outputs(6346));
    outputs(2266) <= layer4_outputs(7590);
    outputs(2267) <= not(layer4_outputs(6754)) or (layer4_outputs(3177));
    outputs(2268) <= (layer4_outputs(4034)) or (layer4_outputs(3726));
    outputs(2269) <= not(layer4_outputs(1756));
    outputs(2270) <= not(layer4_outputs(4570));
    outputs(2271) <= (layer4_outputs(7648)) xor (layer4_outputs(6706));
    outputs(2272) <= layer4_outputs(2541);
    outputs(2273) <= layer4_outputs(7026);
    outputs(2274) <= not(layer4_outputs(3668)) or (layer4_outputs(1982));
    outputs(2275) <= (layer4_outputs(351)) and (layer4_outputs(5360));
    outputs(2276) <= not(layer4_outputs(7455));
    outputs(2277) <= not(layer4_outputs(7304));
    outputs(2278) <= not(layer4_outputs(6023)) or (layer4_outputs(6138));
    outputs(2279) <= (layer4_outputs(6241)) or (layer4_outputs(4186));
    outputs(2280) <= layer4_outputs(6473);
    outputs(2281) <= not((layer4_outputs(97)) xor (layer4_outputs(4571)));
    outputs(2282) <= not(layer4_outputs(2259));
    outputs(2283) <= (layer4_outputs(6247)) xor (layer4_outputs(2179));
    outputs(2284) <= not((layer4_outputs(2094)) xor (layer4_outputs(2447)));
    outputs(2285) <= layer4_outputs(1557);
    outputs(2286) <= layer4_outputs(6515);
    outputs(2287) <= layer4_outputs(316);
    outputs(2288) <= not(layer4_outputs(1482));
    outputs(2289) <= not(layer4_outputs(3652));
    outputs(2290) <= layer4_outputs(6078);
    outputs(2291) <= (layer4_outputs(7661)) and (layer4_outputs(84));
    outputs(2292) <= not(layer4_outputs(73));
    outputs(2293) <= not(layer4_outputs(5140));
    outputs(2294) <= layer4_outputs(7141);
    outputs(2295) <= layer4_outputs(1662);
    outputs(2296) <= layer4_outputs(6480);
    outputs(2297) <= not(layer4_outputs(4634)) or (layer4_outputs(5092));
    outputs(2298) <= not(layer4_outputs(6326));
    outputs(2299) <= layer4_outputs(4180);
    outputs(2300) <= layer4_outputs(5944);
    outputs(2301) <= layer4_outputs(387);
    outputs(2302) <= layer4_outputs(2594);
    outputs(2303) <= layer4_outputs(7349);
    outputs(2304) <= layer4_outputs(2980);
    outputs(2305) <= layer4_outputs(2055);
    outputs(2306) <= layer4_outputs(4293);
    outputs(2307) <= not((layer4_outputs(4856)) and (layer4_outputs(1228)));
    outputs(2308) <= not(layer4_outputs(1291));
    outputs(2309) <= layer4_outputs(4620);
    outputs(2310) <= not(layer4_outputs(3133));
    outputs(2311) <= (layer4_outputs(6281)) and not (layer4_outputs(550));
    outputs(2312) <= not(layer4_outputs(7155)) or (layer4_outputs(6054));
    outputs(2313) <= (layer4_outputs(282)) xor (layer4_outputs(7512));
    outputs(2314) <= layer4_outputs(6609);
    outputs(2315) <= layer4_outputs(6);
    outputs(2316) <= (layer4_outputs(2853)) or (layer4_outputs(5336));
    outputs(2317) <= not((layer4_outputs(1402)) or (layer4_outputs(5126)));
    outputs(2318) <= layer4_outputs(4404);
    outputs(2319) <= layer4_outputs(3816);
    outputs(2320) <= not(layer4_outputs(7389));
    outputs(2321) <= not(layer4_outputs(2148));
    outputs(2322) <= not(layer4_outputs(7428));
    outputs(2323) <= layer4_outputs(3978);
    outputs(2324) <= (layer4_outputs(6211)) and not (layer4_outputs(4977));
    outputs(2325) <= not(layer4_outputs(4897));
    outputs(2326) <= (layer4_outputs(2403)) and not (layer4_outputs(3781));
    outputs(2327) <= (layer4_outputs(3070)) xor (layer4_outputs(832));
    outputs(2328) <= not(layer4_outputs(2444));
    outputs(2329) <= (layer4_outputs(4914)) xor (layer4_outputs(1826));
    outputs(2330) <= not((layer4_outputs(782)) xor (layer4_outputs(6165)));
    outputs(2331) <= (layer4_outputs(1014)) xor (layer4_outputs(6879));
    outputs(2332) <= not(layer4_outputs(1295));
    outputs(2333) <= not(layer4_outputs(5552));
    outputs(2334) <= (layer4_outputs(6526)) xor (layer4_outputs(6736));
    outputs(2335) <= (layer4_outputs(4961)) and not (layer4_outputs(111));
    outputs(2336) <= not(layer4_outputs(7084));
    outputs(2337) <= (layer4_outputs(172)) and (layer4_outputs(4826));
    outputs(2338) <= not((layer4_outputs(3151)) xor (layer4_outputs(1887)));
    outputs(2339) <= not(layer4_outputs(3657));
    outputs(2340) <= not(layer4_outputs(5439));
    outputs(2341) <= not(layer4_outputs(5153));
    outputs(2342) <= layer4_outputs(3576);
    outputs(2343) <= (layer4_outputs(1974)) and (layer4_outputs(2021));
    outputs(2344) <= layer4_outputs(1159);
    outputs(2345) <= not(layer4_outputs(4979));
    outputs(2346) <= layer4_outputs(3596);
    outputs(2347) <= layer4_outputs(4598);
    outputs(2348) <= not((layer4_outputs(5831)) or (layer4_outputs(3441)));
    outputs(2349) <= layer4_outputs(5844);
    outputs(2350) <= not(layer4_outputs(5302));
    outputs(2351) <= (layer4_outputs(7179)) and not (layer4_outputs(1273));
    outputs(2352) <= layer4_outputs(1990);
    outputs(2353) <= layer4_outputs(6766);
    outputs(2354) <= not(layer4_outputs(291));
    outputs(2355) <= not((layer4_outputs(6672)) xor (layer4_outputs(1496)));
    outputs(2356) <= not((layer4_outputs(2700)) xor (layer4_outputs(6526)));
    outputs(2357) <= (layer4_outputs(2616)) and not (layer4_outputs(6810));
    outputs(2358) <= (layer4_outputs(288)) or (layer4_outputs(7031));
    outputs(2359) <= not(layer4_outputs(7029));
    outputs(2360) <= layer4_outputs(5870);
    outputs(2361) <= (layer4_outputs(1124)) and (layer4_outputs(7036));
    outputs(2362) <= (layer4_outputs(1242)) xor (layer4_outputs(4952));
    outputs(2363) <= not(layer4_outputs(286));
    outputs(2364) <= not(layer4_outputs(7099)) or (layer4_outputs(2768));
    outputs(2365) <= not(layer4_outputs(5555));
    outputs(2366) <= (layer4_outputs(398)) xor (layer4_outputs(2472));
    outputs(2367) <= not((layer4_outputs(3376)) or (layer4_outputs(3450)));
    outputs(2368) <= not((layer4_outputs(5033)) or (layer4_outputs(7137)));
    outputs(2369) <= not(layer4_outputs(1930));
    outputs(2370) <= not((layer4_outputs(1588)) xor (layer4_outputs(4170)));
    outputs(2371) <= layer4_outputs(7071);
    outputs(2372) <= layer4_outputs(5315);
    outputs(2373) <= not(layer4_outputs(2604));
    outputs(2374) <= layer4_outputs(6688);
    outputs(2375) <= (layer4_outputs(6455)) xor (layer4_outputs(977));
    outputs(2376) <= (layer4_outputs(2587)) and (layer4_outputs(404));
    outputs(2377) <= not(layer4_outputs(1784));
    outputs(2378) <= not(layer4_outputs(5332)) or (layer4_outputs(1419));
    outputs(2379) <= not(layer4_outputs(6570));
    outputs(2380) <= not((layer4_outputs(4327)) or (layer4_outputs(4567)));
    outputs(2381) <= layer4_outputs(3120);
    outputs(2382) <= (layer4_outputs(5850)) xor (layer4_outputs(2714));
    outputs(2383) <= (layer4_outputs(3643)) and (layer4_outputs(1582));
    outputs(2384) <= not(layer4_outputs(880));
    outputs(2385) <= (layer4_outputs(7412)) xor (layer4_outputs(5571));
    outputs(2386) <= layer4_outputs(2860);
    outputs(2387) <= not(layer4_outputs(6956));
    outputs(2388) <= not(layer4_outputs(3420));
    outputs(2389) <= not(layer4_outputs(2340));
    outputs(2390) <= not(layer4_outputs(7364));
    outputs(2391) <= not((layer4_outputs(5762)) or (layer4_outputs(3930)));
    outputs(2392) <= layer4_outputs(6181);
    outputs(2393) <= layer4_outputs(6212);
    outputs(2394) <= not(layer4_outputs(7428));
    outputs(2395) <= (layer4_outputs(1075)) and (layer4_outputs(3041));
    outputs(2396) <= not(layer4_outputs(4244));
    outputs(2397) <= not(layer4_outputs(5764));
    outputs(2398) <= not(layer4_outputs(3411));
    outputs(2399) <= layer4_outputs(10);
    outputs(2400) <= not((layer4_outputs(235)) or (layer4_outputs(127)));
    outputs(2401) <= not(layer4_outputs(6846));
    outputs(2402) <= not(layer4_outputs(2684));
    outputs(2403) <= not(layer4_outputs(6891));
    outputs(2404) <= not(layer4_outputs(6422));
    outputs(2405) <= not((layer4_outputs(1213)) xor (layer4_outputs(4797)));
    outputs(2406) <= layer4_outputs(7671);
    outputs(2407) <= not(layer4_outputs(7508));
    outputs(2408) <= not(layer4_outputs(6156));
    outputs(2409) <= layer4_outputs(2368);
    outputs(2410) <= not((layer4_outputs(7361)) xor (layer4_outputs(991)));
    outputs(2411) <= not(layer4_outputs(6715));
    outputs(2412) <= layer4_outputs(6611);
    outputs(2413) <= not((layer4_outputs(1694)) xor (layer4_outputs(1395)));
    outputs(2414) <= not(layer4_outputs(5845)) or (layer4_outputs(1085));
    outputs(2415) <= not((layer4_outputs(5528)) and (layer4_outputs(52)));
    outputs(2416) <= not(layer4_outputs(5430));
    outputs(2417) <= not(layer4_outputs(5905)) or (layer4_outputs(7642));
    outputs(2418) <= not(layer4_outputs(2479));
    outputs(2419) <= layer4_outputs(6459);
    outputs(2420) <= layer4_outputs(974);
    outputs(2421) <= layer4_outputs(5593);
    outputs(2422) <= not((layer4_outputs(4262)) and (layer4_outputs(7161)));
    outputs(2423) <= not(layer4_outputs(1815));
    outputs(2424) <= not(layer4_outputs(6666));
    outputs(2425) <= not((layer4_outputs(7153)) xor (layer4_outputs(5642)));
    outputs(2426) <= (layer4_outputs(4370)) and not (layer4_outputs(5451));
    outputs(2427) <= layer4_outputs(7224);
    outputs(2428) <= not(layer4_outputs(1928));
    outputs(2429) <= layer4_outputs(3870);
    outputs(2430) <= (layer4_outputs(5656)) or (layer4_outputs(4665));
    outputs(2431) <= layer4_outputs(2896);
    outputs(2432) <= not(layer4_outputs(3760));
    outputs(2433) <= layer4_outputs(1674);
    outputs(2434) <= not(layer4_outputs(2210));
    outputs(2435) <= (layer4_outputs(3096)) and not (layer4_outputs(5877));
    outputs(2436) <= layer4_outputs(863);
    outputs(2437) <= (layer4_outputs(199)) or (layer4_outputs(5586));
    outputs(2438) <= not(layer4_outputs(1872));
    outputs(2439) <= not(layer4_outputs(4088));
    outputs(2440) <= not(layer4_outputs(7168));
    outputs(2441) <= (layer4_outputs(6957)) and (layer4_outputs(2335));
    outputs(2442) <= not(layer4_outputs(947));
    outputs(2443) <= not(layer4_outputs(4716));
    outputs(2444) <= layer4_outputs(4930);
    outputs(2445) <= layer4_outputs(4886);
    outputs(2446) <= layer4_outputs(6501);
    outputs(2447) <= not(layer4_outputs(1732));
    outputs(2448) <= (layer4_outputs(4651)) and not (layer4_outputs(4269));
    outputs(2449) <= not((layer4_outputs(7045)) or (layer4_outputs(6209)));
    outputs(2450) <= not(layer4_outputs(1247)) or (layer4_outputs(5044));
    outputs(2451) <= not(layer4_outputs(3185)) or (layer4_outputs(6293));
    outputs(2452) <= (layer4_outputs(5568)) and (layer4_outputs(937));
    outputs(2453) <= not(layer4_outputs(3324));
    outputs(2454) <= layer4_outputs(4494);
    outputs(2455) <= layer4_outputs(150);
    outputs(2456) <= layer4_outputs(6882);
    outputs(2457) <= layer4_outputs(5868);
    outputs(2458) <= layer4_outputs(422);
    outputs(2459) <= not((layer4_outputs(7526)) xor (layer4_outputs(589)));
    outputs(2460) <= layer4_outputs(105);
    outputs(2461) <= not((layer4_outputs(1332)) xor (layer4_outputs(1150)));
    outputs(2462) <= layer4_outputs(1091);
    outputs(2463) <= not(layer4_outputs(4808));
    outputs(2464) <= layer4_outputs(2966);
    outputs(2465) <= (layer4_outputs(3372)) xor (layer4_outputs(4270));
    outputs(2466) <= layer4_outputs(604);
    outputs(2467) <= not(layer4_outputs(1871));
    outputs(2468) <= not((layer4_outputs(4557)) xor (layer4_outputs(487)));
    outputs(2469) <= layer4_outputs(5708);
    outputs(2470) <= (layer4_outputs(7635)) and not (layer4_outputs(70));
    outputs(2471) <= layer4_outputs(2345);
    outputs(2472) <= not(layer4_outputs(5613)) or (layer4_outputs(411));
    outputs(2473) <= (layer4_outputs(4764)) and (layer4_outputs(1797));
    outputs(2474) <= not((layer4_outputs(6991)) xor (layer4_outputs(6046)));
    outputs(2475) <= not((layer4_outputs(7591)) xor (layer4_outputs(858)));
    outputs(2476) <= (layer4_outputs(4139)) and (layer4_outputs(4705));
    outputs(2477) <= layer4_outputs(6710);
    outputs(2478) <= layer4_outputs(1968);
    outputs(2479) <= not((layer4_outputs(7501)) xor (layer4_outputs(842)));
    outputs(2480) <= (layer4_outputs(3810)) xor (layer4_outputs(7079));
    outputs(2481) <= not(layer4_outputs(465));
    outputs(2482) <= layer4_outputs(2237);
    outputs(2483) <= not(layer4_outputs(5302));
    outputs(2484) <= not((layer4_outputs(1149)) or (layer4_outputs(2527)));
    outputs(2485) <= not(layer4_outputs(4022));
    outputs(2486) <= not(layer4_outputs(1781));
    outputs(2487) <= not(layer4_outputs(6506));
    outputs(2488) <= layer4_outputs(329);
    outputs(2489) <= not(layer4_outputs(7407));
    outputs(2490) <= not(layer4_outputs(4784));
    outputs(2491) <= (layer4_outputs(1348)) and not (layer4_outputs(4755));
    outputs(2492) <= not(layer4_outputs(6719));
    outputs(2493) <= layer4_outputs(537);
    outputs(2494) <= layer4_outputs(2613);
    outputs(2495) <= not((layer4_outputs(7411)) or (layer4_outputs(5283)));
    outputs(2496) <= layer4_outputs(1884);
    outputs(2497) <= layer4_outputs(4193);
    outputs(2498) <= not(layer4_outputs(4884));
    outputs(2499) <= (layer4_outputs(1127)) and not (layer4_outputs(4315));
    outputs(2500) <= not((layer4_outputs(6242)) xor (layer4_outputs(5127)));
    outputs(2501) <= layer4_outputs(4891);
    outputs(2502) <= not(layer4_outputs(6561));
    outputs(2503) <= layer4_outputs(644);
    outputs(2504) <= (layer4_outputs(714)) xor (layer4_outputs(1545));
    outputs(2505) <= not(layer4_outputs(2049)) or (layer4_outputs(2642));
    outputs(2506) <= not(layer4_outputs(4065));
    outputs(2507) <= (layer4_outputs(7674)) xor (layer4_outputs(5354));
    outputs(2508) <= not(layer4_outputs(690));
    outputs(2509) <= layer4_outputs(2294);
    outputs(2510) <= layer4_outputs(6983);
    outputs(2511) <= not(layer4_outputs(6322));
    outputs(2512) <= not(layer4_outputs(1262));
    outputs(2513) <= (layer4_outputs(5589)) xor (layer4_outputs(5012));
    outputs(2514) <= not(layer4_outputs(6391));
    outputs(2515) <= not(layer4_outputs(448));
    outputs(2516) <= not(layer4_outputs(5920));
    outputs(2517) <= (layer4_outputs(3179)) or (layer4_outputs(7492));
    outputs(2518) <= not(layer4_outputs(3067));
    outputs(2519) <= not((layer4_outputs(1433)) xor (layer4_outputs(5562)));
    outputs(2520) <= layer4_outputs(6405);
    outputs(2521) <= layer4_outputs(6308);
    outputs(2522) <= layer4_outputs(621);
    outputs(2523) <= not(layer4_outputs(7561));
    outputs(2524) <= (layer4_outputs(2894)) and (layer4_outputs(6177));
    outputs(2525) <= layer4_outputs(2099);
    outputs(2526) <= not(layer4_outputs(633)) or (layer4_outputs(3661));
    outputs(2527) <= (layer4_outputs(1226)) and (layer4_outputs(7485));
    outputs(2528) <= layer4_outputs(107);
    outputs(2529) <= layer4_outputs(3115);
    outputs(2530) <= not((layer4_outputs(6256)) xor (layer4_outputs(4015)));
    outputs(2531) <= not(layer4_outputs(573));
    outputs(2532) <= layer4_outputs(4442);
    outputs(2533) <= layer4_outputs(5840);
    outputs(2534) <= (layer4_outputs(3127)) xor (layer4_outputs(3147));
    outputs(2535) <= not(layer4_outputs(6271));
    outputs(2536) <= not((layer4_outputs(4397)) xor (layer4_outputs(642)));
    outputs(2537) <= not(layer4_outputs(3236)) or (layer4_outputs(6065));
    outputs(2538) <= not(layer4_outputs(5673)) or (layer4_outputs(4723));
    outputs(2539) <= not(layer4_outputs(1115));
    outputs(2540) <= not(layer4_outputs(5205));
    outputs(2541) <= layer4_outputs(3129);
    outputs(2542) <= not(layer4_outputs(241));
    outputs(2543) <= (layer4_outputs(6454)) xor (layer4_outputs(281));
    outputs(2544) <= not(layer4_outputs(1741));
    outputs(2545) <= layer4_outputs(6968);
    outputs(2546) <= (layer4_outputs(3762)) and not (layer4_outputs(4696));
    outputs(2547) <= layer4_outputs(6628);
    outputs(2548) <= not(layer4_outputs(5990));
    outputs(2549) <= layer4_outputs(7210);
    outputs(2550) <= layer4_outputs(5266);
    outputs(2551) <= not(layer4_outputs(6502));
    outputs(2552) <= (layer4_outputs(7423)) xor (layer4_outputs(1971));
    outputs(2553) <= not(layer4_outputs(3325));
    outputs(2554) <= (layer4_outputs(3306)) and not (layer4_outputs(1134));
    outputs(2555) <= not(layer4_outputs(598));
    outputs(2556) <= layer4_outputs(5554);
    outputs(2557) <= not(layer4_outputs(2675));
    outputs(2558) <= layer4_outputs(3968);
    outputs(2559) <= not(layer4_outputs(2221));
    outputs(2560) <= not((layer4_outputs(1056)) xor (layer4_outputs(1916)));
    outputs(2561) <= layer4_outputs(1512);
    outputs(2562) <= layer4_outputs(7316);
    outputs(2563) <= layer4_outputs(63);
    outputs(2564) <= not(layer4_outputs(5159));
    outputs(2565) <= layer4_outputs(3347);
    outputs(2566) <= layer4_outputs(1977);
    outputs(2567) <= (layer4_outputs(4485)) and (layer4_outputs(576));
    outputs(2568) <= (layer4_outputs(2308)) and not (layer4_outputs(1427));
    outputs(2569) <= layer4_outputs(3260);
    outputs(2570) <= not(layer4_outputs(4018));
    outputs(2571) <= layer4_outputs(4479);
    outputs(2572) <= not(layer4_outputs(477));
    outputs(2573) <= not(layer4_outputs(4399));
    outputs(2574) <= layer4_outputs(2486);
    outputs(2575) <= not((layer4_outputs(1804)) xor (layer4_outputs(6943)));
    outputs(2576) <= (layer4_outputs(2807)) and (layer4_outputs(5244));
    outputs(2577) <= layer4_outputs(5109);
    outputs(2578) <= not(layer4_outputs(327));
    outputs(2579) <= not((layer4_outputs(7374)) xor (layer4_outputs(4499)));
    outputs(2580) <= layer4_outputs(1968);
    outputs(2581) <= not((layer4_outputs(1075)) xor (layer4_outputs(3391)));
    outputs(2582) <= not(layer4_outputs(7236));
    outputs(2583) <= not(layer4_outputs(4716));
    outputs(2584) <= not(layer4_outputs(1698));
    outputs(2585) <= not((layer4_outputs(3112)) or (layer4_outputs(7112)));
    outputs(2586) <= layer4_outputs(6450);
    outputs(2587) <= not(layer4_outputs(489));
    outputs(2588) <= not(layer4_outputs(6471));
    outputs(2589) <= (layer4_outputs(4309)) and not (layer4_outputs(5056));
    outputs(2590) <= (layer4_outputs(3208)) xor (layer4_outputs(1343));
    outputs(2591) <= layer4_outputs(802);
    outputs(2592) <= not(layer4_outputs(7639));
    outputs(2593) <= layer4_outputs(6872);
    outputs(2594) <= not((layer4_outputs(3033)) and (layer4_outputs(5736)));
    outputs(2595) <= not((layer4_outputs(830)) xor (layer4_outputs(3401)));
    outputs(2596) <= layer4_outputs(5089);
    outputs(2597) <= not(layer4_outputs(7260));
    outputs(2598) <= layer4_outputs(4814);
    outputs(2599) <= not(layer4_outputs(5634));
    outputs(2600) <= (layer4_outputs(5713)) xor (layer4_outputs(5662));
    outputs(2601) <= (layer4_outputs(3307)) xor (layer4_outputs(1510));
    outputs(2602) <= layer4_outputs(7608);
    outputs(2603) <= not(layer4_outputs(4437));
    outputs(2604) <= (layer4_outputs(5680)) and not (layer4_outputs(2697));
    outputs(2605) <= not(layer4_outputs(1352));
    outputs(2606) <= not((layer4_outputs(6589)) or (layer4_outputs(5300)));
    outputs(2607) <= not(layer4_outputs(466)) or (layer4_outputs(1876));
    outputs(2608) <= (layer4_outputs(6728)) and not (layer4_outputs(1759));
    outputs(2609) <= not(layer4_outputs(3236));
    outputs(2610) <= layer4_outputs(2653);
    outputs(2611) <= (layer4_outputs(3169)) and (layer4_outputs(607));
    outputs(2612) <= (layer4_outputs(5637)) and (layer4_outputs(6237));
    outputs(2613) <= not(layer4_outputs(153));
    outputs(2614) <= not(layer4_outputs(1087));
    outputs(2615) <= layer4_outputs(6495);
    outputs(2616) <= not(layer4_outputs(5075)) or (layer4_outputs(4400));
    outputs(2617) <= layer4_outputs(2732);
    outputs(2618) <= (layer4_outputs(3496)) and not (layer4_outputs(669));
    outputs(2619) <= layer4_outputs(6363);
    outputs(2620) <= not(layer4_outputs(3881));
    outputs(2621) <= layer4_outputs(7190);
    outputs(2622) <= not(layer4_outputs(4092));
    outputs(2623) <= not(layer4_outputs(1892));
    outputs(2624) <= (layer4_outputs(6369)) xor (layer4_outputs(3625));
    outputs(2625) <= not((layer4_outputs(1467)) xor (layer4_outputs(7287)));
    outputs(2626) <= not(layer4_outputs(3925)) or (layer4_outputs(3093));
    outputs(2627) <= (layer4_outputs(5053)) and not (layer4_outputs(5574));
    outputs(2628) <= not(layer4_outputs(1279));
    outputs(2629) <= layer4_outputs(6541);
    outputs(2630) <= not(layer4_outputs(1142));
    outputs(2631) <= not(layer4_outputs(5673));
    outputs(2632) <= not(layer4_outputs(4636));
    outputs(2633) <= (layer4_outputs(3308)) and not (layer4_outputs(1158));
    outputs(2634) <= not(layer4_outputs(3945));
    outputs(2635) <= not(layer4_outputs(7278)) or (layer4_outputs(2010));
    outputs(2636) <= (layer4_outputs(5963)) and not (layer4_outputs(2434));
    outputs(2637) <= layer4_outputs(2629);
    outputs(2638) <= (layer4_outputs(1552)) xor (layer4_outputs(826));
    outputs(2639) <= layer4_outputs(5428);
    outputs(2640) <= not(layer4_outputs(2098));
    outputs(2641) <= layer4_outputs(5496);
    outputs(2642) <= not((layer4_outputs(5715)) xor (layer4_outputs(3526)));
    outputs(2643) <= not(layer4_outputs(4815));
    outputs(2644) <= layer4_outputs(4975);
    outputs(2645) <= layer4_outputs(3203);
    outputs(2646) <= not(layer4_outputs(5304));
    outputs(2647) <= not(layer4_outputs(5200));
    outputs(2648) <= not(layer4_outputs(4420));
    outputs(2649) <= not((layer4_outputs(7303)) xor (layer4_outputs(4869)));
    outputs(2650) <= not((layer4_outputs(1039)) xor (layer4_outputs(5364)));
    outputs(2651) <= (layer4_outputs(5436)) xor (layer4_outputs(4409));
    outputs(2652) <= not(layer4_outputs(4670));
    outputs(2653) <= not(layer4_outputs(1827));
    outputs(2654) <= (layer4_outputs(4111)) xor (layer4_outputs(2385));
    outputs(2655) <= not((layer4_outputs(3754)) and (layer4_outputs(486)));
    outputs(2656) <= layer4_outputs(2308);
    outputs(2657) <= layer4_outputs(4430);
    outputs(2658) <= not((layer4_outputs(5061)) or (layer4_outputs(6745)));
    outputs(2659) <= not(layer4_outputs(6757)) or (layer4_outputs(1586));
    outputs(2660) <= not((layer4_outputs(7127)) or (layer4_outputs(3270)));
    outputs(2661) <= layer4_outputs(2812);
    outputs(2662) <= not(layer4_outputs(3124));
    outputs(2663) <= not(layer4_outputs(6414)) or (layer4_outputs(5648));
    outputs(2664) <= layer4_outputs(5117);
    outputs(2665) <= layer4_outputs(4798);
    outputs(2666) <= (layer4_outputs(1376)) and not (layer4_outputs(2050));
    outputs(2667) <= not(layer4_outputs(448));
    outputs(2668) <= (layer4_outputs(4035)) and (layer4_outputs(820));
    outputs(2669) <= (layer4_outputs(2610)) and (layer4_outputs(7300));
    outputs(2670) <= not((layer4_outputs(4846)) xor (layer4_outputs(5738)));
    outputs(2671) <= not((layer4_outputs(5136)) or (layer4_outputs(1660)));
    outputs(2672) <= (layer4_outputs(6635)) xor (layer4_outputs(6249));
    outputs(2673) <= not(layer4_outputs(6831));
    outputs(2674) <= not((layer4_outputs(7644)) or (layer4_outputs(7582)));
    outputs(2675) <= layer4_outputs(718);
    outputs(2676) <= not(layer4_outputs(2617));
    outputs(2677) <= not(layer4_outputs(4491));
    outputs(2678) <= layer4_outputs(5486);
    outputs(2679) <= not((layer4_outputs(6449)) xor (layer4_outputs(2419)));
    outputs(2680) <= (layer4_outputs(2160)) xor (layer4_outputs(1499));
    outputs(2681) <= not(layer4_outputs(4774));
    outputs(2682) <= not(layer4_outputs(5820));
    outputs(2683) <= layer4_outputs(3627);
    outputs(2684) <= not(layer4_outputs(4538));
    outputs(2685) <= not(layer4_outputs(5342));
    outputs(2686) <= layer4_outputs(5974);
    outputs(2687) <= not(layer4_outputs(3466));
    outputs(2688) <= not(layer4_outputs(2228));
    outputs(2689) <= not(layer4_outputs(2327));
    outputs(2690) <= (layer4_outputs(5341)) and not (layer4_outputs(7221));
    outputs(2691) <= not(layer4_outputs(3052));
    outputs(2692) <= layer4_outputs(7355);
    outputs(2693) <= layer4_outputs(7214);
    outputs(2694) <= not((layer4_outputs(2656)) xor (layer4_outputs(924)));
    outputs(2695) <= not(layer4_outputs(2942));
    outputs(2696) <= not(layer4_outputs(5225));
    outputs(2697) <= not(layer4_outputs(7309));
    outputs(2698) <= not(layer4_outputs(503));
    outputs(2699) <= not((layer4_outputs(4049)) xor (layer4_outputs(4261)));
    outputs(2700) <= layer4_outputs(785);
    outputs(2701) <= not(layer4_outputs(504)) or (layer4_outputs(4161));
    outputs(2702) <= (layer4_outputs(1820)) xor (layer4_outputs(101));
    outputs(2703) <= not((layer4_outputs(1040)) and (layer4_outputs(1710)));
    outputs(2704) <= not(layer4_outputs(2027)) or (layer4_outputs(7477));
    outputs(2705) <= not((layer4_outputs(4955)) and (layer4_outputs(4320)));
    outputs(2706) <= not(layer4_outputs(1006));
    outputs(2707) <= layer4_outputs(6161);
    outputs(2708) <= not((layer4_outputs(5609)) or (layer4_outputs(5513)));
    outputs(2709) <= (layer4_outputs(421)) and (layer4_outputs(2293));
    outputs(2710) <= not(layer4_outputs(254));
    outputs(2711) <= layer4_outputs(1914);
    outputs(2712) <= layer4_outputs(958);
    outputs(2713) <= layer4_outputs(183);
    outputs(2714) <= not((layer4_outputs(7668)) xor (layer4_outputs(6806)));
    outputs(2715) <= not((layer4_outputs(1765)) and (layer4_outputs(6942)));
    outputs(2716) <= not(layer4_outputs(6756)) or (layer4_outputs(939));
    outputs(2717) <= not(layer4_outputs(4100));
    outputs(2718) <= not((layer4_outputs(871)) or (layer4_outputs(192)));
    outputs(2719) <= not((layer4_outputs(6493)) xor (layer4_outputs(853)));
    outputs(2720) <= not(layer4_outputs(7363));
    outputs(2721) <= (layer4_outputs(3454)) xor (layer4_outputs(3497));
    outputs(2722) <= layer4_outputs(2642);
    outputs(2723) <= (layer4_outputs(5941)) and not (layer4_outputs(3353));
    outputs(2724) <= not(layer4_outputs(7281));
    outputs(2725) <= (layer4_outputs(1425)) and not (layer4_outputs(6452));
    outputs(2726) <= not(layer4_outputs(5953));
    outputs(2727) <= (layer4_outputs(5128)) xor (layer4_outputs(2392));
    outputs(2728) <= (layer4_outputs(6091)) and not (layer4_outputs(104));
    outputs(2729) <= (layer4_outputs(2446)) and (layer4_outputs(4359));
    outputs(2730) <= not(layer4_outputs(6844));
    outputs(2731) <= (layer4_outputs(196)) and (layer4_outputs(6103));
    outputs(2732) <= layer4_outputs(7570);
    outputs(2733) <= (layer4_outputs(2386)) xor (layer4_outputs(3307));
    outputs(2734) <= (layer4_outputs(3670)) xor (layer4_outputs(4416));
    outputs(2735) <= not(layer4_outputs(385));
    outputs(2736) <= (layer4_outputs(3054)) xor (layer4_outputs(7140));
    outputs(2737) <= layer4_outputs(3313);
    outputs(2738) <= not(layer4_outputs(410)) or (layer4_outputs(5542));
    outputs(2739) <= not((layer4_outputs(6347)) xor (layer4_outputs(945)));
    outputs(2740) <= not(layer4_outputs(3736));
    outputs(2741) <= layer4_outputs(3631);
    outputs(2742) <= (layer4_outputs(136)) and not (layer4_outputs(5505));
    outputs(2743) <= (layer4_outputs(6680)) xor (layer4_outputs(4600));
    outputs(2744) <= layer4_outputs(2311);
    outputs(2745) <= not((layer4_outputs(2353)) or (layer4_outputs(1420)));
    outputs(2746) <= not(layer4_outputs(4566));
    outputs(2747) <= layer4_outputs(6427);
    outputs(2748) <= not((layer4_outputs(2633)) xor (layer4_outputs(3960)));
    outputs(2749) <= layer4_outputs(3104);
    outputs(2750) <= (layer4_outputs(6117)) and (layer4_outputs(7426));
    outputs(2751) <= (layer4_outputs(6606)) and not (layer4_outputs(7109));
    outputs(2752) <= layer4_outputs(3306);
    outputs(2753) <= layer4_outputs(2294);
    outputs(2754) <= not((layer4_outputs(1528)) or (layer4_outputs(4237)));
    outputs(2755) <= layer4_outputs(2581);
    outputs(2756) <= layer4_outputs(6525);
    outputs(2757) <= not((layer4_outputs(5762)) or (layer4_outputs(1899)));
    outputs(2758) <= not(layer4_outputs(3053));
    outputs(2759) <= layer4_outputs(3884);
    outputs(2760) <= (layer4_outputs(7496)) and (layer4_outputs(2998));
    outputs(2761) <= not(layer4_outputs(1100));
    outputs(2762) <= layer4_outputs(6037);
    outputs(2763) <= layer4_outputs(4562);
    outputs(2764) <= layer4_outputs(1341);
    outputs(2765) <= not((layer4_outputs(7554)) or (layer4_outputs(4689)));
    outputs(2766) <= (layer4_outputs(3695)) xor (layer4_outputs(4266));
    outputs(2767) <= layer4_outputs(7209);
    outputs(2768) <= not((layer4_outputs(6922)) xor (layer4_outputs(5703)));
    outputs(2769) <= not(layer4_outputs(5655));
    outputs(2770) <= not(layer4_outputs(6527));
    outputs(2771) <= not((layer4_outputs(1436)) xor (layer4_outputs(2788)));
    outputs(2772) <= layer4_outputs(1564);
    outputs(2773) <= not(layer4_outputs(1133)) or (layer4_outputs(3707));
    outputs(2774) <= layer4_outputs(515);
    outputs(2775) <= not((layer4_outputs(5086)) and (layer4_outputs(6371)));
    outputs(2776) <= layer4_outputs(278);
    outputs(2777) <= (layer4_outputs(4527)) and not (layer4_outputs(1848));
    outputs(2778) <= not(layer4_outputs(2890));
    outputs(2779) <= not((layer4_outputs(269)) or (layer4_outputs(3144)));
    outputs(2780) <= layer4_outputs(904);
    outputs(2781) <= not((layer4_outputs(5383)) and (layer4_outputs(7170)));
    outputs(2782) <= (layer4_outputs(6856)) and not (layer4_outputs(5509));
    outputs(2783) <= not((layer4_outputs(4820)) or (layer4_outputs(5399)));
    outputs(2784) <= layer4_outputs(6849);
    outputs(2785) <= layer4_outputs(1549);
    outputs(2786) <= layer4_outputs(4313);
    outputs(2787) <= not((layer4_outputs(1291)) xor (layer4_outputs(4498)));
    outputs(2788) <= not((layer4_outputs(5661)) xor (layer4_outputs(1604)));
    outputs(2789) <= not(layer4_outputs(6695)) or (layer4_outputs(5797));
    outputs(2790) <= (layer4_outputs(5408)) xor (layer4_outputs(5179));
    outputs(2791) <= not(layer4_outputs(7592));
    outputs(2792) <= layer4_outputs(5244);
    outputs(2793) <= not(layer4_outputs(2889)) or (layer4_outputs(7413));
    outputs(2794) <= not((layer4_outputs(1463)) or (layer4_outputs(6776)));
    outputs(2795) <= layer4_outputs(2473);
    outputs(2796) <= layer4_outputs(5928);
    outputs(2797) <= not(layer4_outputs(3480));
    outputs(2798) <= not(layer4_outputs(1163));
    outputs(2799) <= not(layer4_outputs(206));
    outputs(2800) <= not((layer4_outputs(3097)) and (layer4_outputs(2549)));
    outputs(2801) <= not((layer4_outputs(275)) xor (layer4_outputs(3269)));
    outputs(2802) <= not(layer4_outputs(7509));
    outputs(2803) <= (layer4_outputs(503)) xor (layer4_outputs(1176));
    outputs(2804) <= not(layer4_outputs(342));
    outputs(2805) <= (layer4_outputs(1541)) or (layer4_outputs(3862));
    outputs(2806) <= not((layer4_outputs(3188)) xor (layer4_outputs(541)));
    outputs(2807) <= (layer4_outputs(4152)) xor (layer4_outputs(3477));
    outputs(2808) <= layer4_outputs(1605);
    outputs(2809) <= not(layer4_outputs(6889)) or (layer4_outputs(2371));
    outputs(2810) <= not(layer4_outputs(5299));
    outputs(2811) <= layer4_outputs(6829);
    outputs(2812) <= not(layer4_outputs(6664));
    outputs(2813) <= not(layer4_outputs(7640)) or (layer4_outputs(6596));
    outputs(2814) <= (layer4_outputs(5014)) and (layer4_outputs(2026));
    outputs(2815) <= layer4_outputs(23);
    outputs(2816) <= (layer4_outputs(3853)) and (layer4_outputs(445));
    outputs(2817) <= (layer4_outputs(2861)) and not (layer4_outputs(3512));
    outputs(2818) <= layer4_outputs(956);
    outputs(2819) <= layer4_outputs(3402);
    outputs(2820) <= not(layer4_outputs(7450));
    outputs(2821) <= layer4_outputs(5806);
    outputs(2822) <= (layer4_outputs(5098)) and not (layer4_outputs(620));
    outputs(2823) <= (layer4_outputs(1615)) or (layer4_outputs(2492));
    outputs(2824) <= not(layer4_outputs(4157)) or (layer4_outputs(6523));
    outputs(2825) <= (layer4_outputs(3083)) and (layer4_outputs(1498));
    outputs(2826) <= not((layer4_outputs(4767)) xor (layer4_outputs(4725)));
    outputs(2827) <= not(layer4_outputs(1838));
    outputs(2828) <= (layer4_outputs(3341)) and not (layer4_outputs(5020));
    outputs(2829) <= (layer4_outputs(3149)) xor (layer4_outputs(6172));
    outputs(2830) <= not(layer4_outputs(7667));
    outputs(2831) <= not(layer4_outputs(1761));
    outputs(2832) <= not(layer4_outputs(1667));
    outputs(2833) <= layer4_outputs(498);
    outputs(2834) <= not(layer4_outputs(2552));
    outputs(2835) <= not(layer4_outputs(6074));
    outputs(2836) <= layer4_outputs(6531);
    outputs(2837) <= layer4_outputs(6084);
    outputs(2838) <= layer4_outputs(4432);
    outputs(2839) <= (layer4_outputs(5172)) and (layer4_outputs(1335));
    outputs(2840) <= (layer4_outputs(6053)) and not (layer4_outputs(6287));
    outputs(2841) <= layer4_outputs(4972);
    outputs(2842) <= not(layer4_outputs(3146));
    outputs(2843) <= not(layer4_outputs(5232));
    outputs(2844) <= not(layer4_outputs(3474)) or (layer4_outputs(1318));
    outputs(2845) <= layer4_outputs(6964);
    outputs(2846) <= not((layer4_outputs(4756)) or (layer4_outputs(2736)));
    outputs(2847) <= not(layer4_outputs(4835));
    outputs(2848) <= layer4_outputs(1019);
    outputs(2849) <= (layer4_outputs(1785)) xor (layer4_outputs(530));
    outputs(2850) <= not(layer4_outputs(1636));
    outputs(2851) <= layer4_outputs(1882);
    outputs(2852) <= not((layer4_outputs(6262)) xor (layer4_outputs(7632)));
    outputs(2853) <= layer4_outputs(1164);
    outputs(2854) <= not(layer4_outputs(877));
    outputs(2855) <= layer4_outputs(56);
    outputs(2856) <= (layer4_outputs(6785)) or (layer4_outputs(6968));
    outputs(2857) <= not(layer4_outputs(1956));
    outputs(2858) <= not(layer4_outputs(4559));
    outputs(2859) <= not(layer4_outputs(2866));
    outputs(2860) <= layer4_outputs(814);
    outputs(2861) <= not(layer4_outputs(2715));
    outputs(2862) <= layer4_outputs(4707);
    outputs(2863) <= (layer4_outputs(3775)) and (layer4_outputs(7210));
    outputs(2864) <= not((layer4_outputs(6260)) or (layer4_outputs(3173)));
    outputs(2865) <= (layer4_outputs(5929)) and not (layer4_outputs(1745));
    outputs(2866) <= not(layer4_outputs(3122));
    outputs(2867) <= (layer4_outputs(3792)) xor (layer4_outputs(3537));
    outputs(2868) <= not(layer4_outputs(3628));
    outputs(2869) <= (layer4_outputs(3280)) xor (layer4_outputs(1824));
    outputs(2870) <= layer4_outputs(1551);
    outputs(2871) <= layer4_outputs(6592);
    outputs(2872) <= (layer4_outputs(847)) and not (layer4_outputs(2958));
    outputs(2873) <= not(layer4_outputs(5541));
    outputs(2874) <= not(layer4_outputs(5116));
    outputs(2875) <= layer4_outputs(6089);
    outputs(2876) <= layer4_outputs(145);
    outputs(2877) <= not(layer4_outputs(3745)) or (layer4_outputs(177));
    outputs(2878) <= not(layer4_outputs(3962));
    outputs(2879) <= not((layer4_outputs(1760)) or (layer4_outputs(3211)));
    outputs(2880) <= (layer4_outputs(7156)) xor (layer4_outputs(6904));
    outputs(2881) <= layer4_outputs(2798);
    outputs(2882) <= layer4_outputs(2562);
    outputs(2883) <= (layer4_outputs(5539)) xor (layer4_outputs(1323));
    outputs(2884) <= not(layer4_outputs(580));
    outputs(2885) <= layer4_outputs(6610);
    outputs(2886) <= not((layer4_outputs(4815)) and (layer4_outputs(6633)));
    outputs(2887) <= (layer4_outputs(1081)) and not (layer4_outputs(3268));
    outputs(2888) <= layer4_outputs(6426);
    outputs(2889) <= not(layer4_outputs(1004)) or (layer4_outputs(4076));
    outputs(2890) <= not(layer4_outputs(1469));
    outputs(2891) <= not((layer4_outputs(4606)) xor (layer4_outputs(2417)));
    outputs(2892) <= layer4_outputs(4264);
    outputs(2893) <= (layer4_outputs(5895)) and not (layer4_outputs(2491));
    outputs(2894) <= layer4_outputs(1716);
    outputs(2895) <= not(layer4_outputs(3786));
    outputs(2896) <= layer4_outputs(3159);
    outputs(2897) <= not((layer4_outputs(3856)) or (layer4_outputs(5275)));
    outputs(2898) <= layer4_outputs(2512);
    outputs(2899) <= layer4_outputs(2984);
    outputs(2900) <= layer4_outputs(3978);
    outputs(2901) <= not(layer4_outputs(2201)) or (layer4_outputs(6313));
    outputs(2902) <= layer4_outputs(3221);
    outputs(2903) <= not((layer4_outputs(6916)) xor (layer4_outputs(2243)));
    outputs(2904) <= layer4_outputs(5226);
    outputs(2905) <= (layer4_outputs(7337)) xor (layer4_outputs(1118));
    outputs(2906) <= not(layer4_outputs(3163));
    outputs(2907) <= not(layer4_outputs(6895));
    outputs(2908) <= not(layer4_outputs(408));
    outputs(2909) <= (layer4_outputs(4535)) and not (layer4_outputs(2384));
    outputs(2910) <= layer4_outputs(6913);
    outputs(2911) <= not(layer4_outputs(5283));
    outputs(2912) <= layer4_outputs(5419);
    outputs(2913) <= not(layer4_outputs(6636));
    outputs(2914) <= not((layer4_outputs(5217)) xor (layer4_outputs(1074)));
    outputs(2915) <= layer4_outputs(1334);
    outputs(2916) <= not(layer4_outputs(372));
    outputs(2917) <= layer4_outputs(886);
    outputs(2918) <= not((layer4_outputs(6602)) xor (layer4_outputs(7508)));
    outputs(2919) <= layer4_outputs(903);
    outputs(2920) <= (layer4_outputs(6373)) and not (layer4_outputs(4865));
    outputs(2921) <= (layer4_outputs(19)) and not (layer4_outputs(1986));
    outputs(2922) <= (layer4_outputs(4048)) and not (layer4_outputs(4493));
    outputs(2923) <= (layer4_outputs(3151)) xor (layer4_outputs(7679));
    outputs(2924) <= (layer4_outputs(1282)) and not (layer4_outputs(2204));
    outputs(2925) <= (layer4_outputs(2313)) and not (layer4_outputs(2434));
    outputs(2926) <= layer4_outputs(5240);
    outputs(2927) <= layer4_outputs(2906);
    outputs(2928) <= (layer4_outputs(4750)) and not (layer4_outputs(1239));
    outputs(2929) <= (layer4_outputs(6466)) and (layer4_outputs(3119));
    outputs(2930) <= layer4_outputs(399);
    outputs(2931) <= layer4_outputs(724);
    outputs(2932) <= not(layer4_outputs(6795));
    outputs(2933) <= (layer4_outputs(611)) and not (layer4_outputs(7097));
    outputs(2934) <= layer4_outputs(3426);
    outputs(2935) <= (layer4_outputs(5899)) xor (layer4_outputs(6623));
    outputs(2936) <= (layer4_outputs(7404)) xor (layer4_outputs(655));
    outputs(2937) <= not(layer4_outputs(3146));
    outputs(2938) <= layer4_outputs(3559);
    outputs(2939) <= not(layer4_outputs(5992));
    outputs(2940) <= not(layer4_outputs(643)) or (layer4_outputs(2107));
    outputs(2941) <= layer4_outputs(1580);
    outputs(2942) <= (layer4_outputs(3638)) and (layer4_outputs(1270));
    outputs(2943) <= not(layer4_outputs(2929)) or (layer4_outputs(1091));
    outputs(2944) <= not((layer4_outputs(1269)) xor (layer4_outputs(4317)));
    outputs(2945) <= layer4_outputs(7542);
    outputs(2946) <= (layer4_outputs(982)) and not (layer4_outputs(5395));
    outputs(2947) <= layer4_outputs(1905);
    outputs(2948) <= not(layer4_outputs(1133));
    outputs(2949) <= not(layer4_outputs(3060));
    outputs(2950) <= not(layer4_outputs(345));
    outputs(2951) <= layer4_outputs(5376);
    outputs(2952) <= layer4_outputs(6143);
    outputs(2953) <= not(layer4_outputs(4863));
    outputs(2954) <= not((layer4_outputs(1658)) xor (layer4_outputs(3562)));
    outputs(2955) <= not(layer4_outputs(5187));
    outputs(2956) <= not(layer4_outputs(3322));
    outputs(2957) <= (layer4_outputs(2410)) and (layer4_outputs(7387));
    outputs(2958) <= not((layer4_outputs(1184)) xor (layer4_outputs(6468)));
    outputs(2959) <= layer4_outputs(3196);
    outputs(2960) <= layer4_outputs(236);
    outputs(2961) <= not(layer4_outputs(2606));
    outputs(2962) <= layer4_outputs(5934);
    outputs(2963) <= not(layer4_outputs(779));
    outputs(2964) <= layer4_outputs(6544);
    outputs(2965) <= layer4_outputs(3873);
    outputs(2966) <= not(layer4_outputs(879));
    outputs(2967) <= layer4_outputs(2477);
    outputs(2968) <= not(layer4_outputs(6460));
    outputs(2969) <= (layer4_outputs(5599)) and (layer4_outputs(558));
    outputs(2970) <= not(layer4_outputs(6199));
    outputs(2971) <= layer4_outputs(6722);
    outputs(2972) <= not((layer4_outputs(7130)) xor (layer4_outputs(4917)));
    outputs(2973) <= not((layer4_outputs(6828)) xor (layer4_outputs(6682)));
    outputs(2974) <= layer4_outputs(6781);
    outputs(2975) <= not(layer4_outputs(368));
    outputs(2976) <= not((layer4_outputs(3142)) xor (layer4_outputs(5203)));
    outputs(2977) <= not(layer4_outputs(4799));
    outputs(2978) <= (layer4_outputs(1969)) and not (layer4_outputs(4185));
    outputs(2979) <= not(layer4_outputs(2356));
    outputs(2980) <= layer4_outputs(341);
    outputs(2981) <= not(layer4_outputs(4855));
    outputs(2982) <= layer4_outputs(6495);
    outputs(2983) <= layer4_outputs(2388);
    outputs(2984) <= (layer4_outputs(1183)) xor (layer4_outputs(4460));
    outputs(2985) <= not((layer4_outputs(5933)) xor (layer4_outputs(44)));
    outputs(2986) <= layer4_outputs(3299);
    outputs(2987) <= (layer4_outputs(749)) and not (layer4_outputs(2644));
    outputs(2988) <= not(layer4_outputs(7567));
    outputs(2989) <= not(layer4_outputs(652));
    outputs(2990) <= not(layer4_outputs(5159));
    outputs(2991) <= (layer4_outputs(6048)) xor (layer4_outputs(4342));
    outputs(2992) <= not(layer4_outputs(2743));
    outputs(2993) <= not(layer4_outputs(4269));
    outputs(2994) <= (layer4_outputs(7265)) xor (layer4_outputs(713));
    outputs(2995) <= (layer4_outputs(6842)) and not (layer4_outputs(331));
    outputs(2996) <= layer4_outputs(2341);
    outputs(2997) <= not(layer4_outputs(6751)) or (layer4_outputs(3398));
    outputs(2998) <= not(layer4_outputs(496));
    outputs(2999) <= not(layer4_outputs(4928));
    outputs(3000) <= not(layer4_outputs(6075));
    outputs(3001) <= layer4_outputs(7572);
    outputs(3002) <= layer4_outputs(4874);
    outputs(3003) <= (layer4_outputs(2706)) or (layer4_outputs(4838));
    outputs(3004) <= not(layer4_outputs(1846));
    outputs(3005) <= not((layer4_outputs(529)) xor (layer4_outputs(7437)));
    outputs(3006) <= not(layer4_outputs(4018));
    outputs(3007) <= (layer4_outputs(3931)) xor (layer4_outputs(5300));
    outputs(3008) <= layer4_outputs(3375);
    outputs(3009) <= layer4_outputs(1513);
    outputs(3010) <= not(layer4_outputs(3906));
    outputs(3011) <= not(layer4_outputs(4802));
    outputs(3012) <= (layer4_outputs(1106)) xor (layer4_outputs(4025));
    outputs(3013) <= (layer4_outputs(5021)) and (layer4_outputs(3922));
    outputs(3014) <= (layer4_outputs(4263)) or (layer4_outputs(3282));
    outputs(3015) <= not(layer4_outputs(4197));
    outputs(3016) <= not((layer4_outputs(3997)) xor (layer4_outputs(337)));
    outputs(3017) <= not(layer4_outputs(6304));
    outputs(3018) <= not(layer4_outputs(2407));
    outputs(3019) <= not((layer4_outputs(1717)) xor (layer4_outputs(3179)));
    outputs(3020) <= (layer4_outputs(6182)) and not (layer4_outputs(3218));
    outputs(3021) <= layer4_outputs(5339);
    outputs(3022) <= not((layer4_outputs(1367)) or (layer4_outputs(6768)));
    outputs(3023) <= not(layer4_outputs(2946));
    outputs(3024) <= layer4_outputs(3718);
    outputs(3025) <= not(layer4_outputs(2766));
    outputs(3026) <= layer4_outputs(6444);
    outputs(3027) <= layer4_outputs(377);
    outputs(3028) <= layer4_outputs(2823);
    outputs(3029) <= layer4_outputs(4877);
    outputs(3030) <= not(layer4_outputs(50));
    outputs(3031) <= not(layer4_outputs(264));
    outputs(3032) <= layer4_outputs(347);
    outputs(3033) <= not(layer4_outputs(6812));
    outputs(3034) <= (layer4_outputs(7191)) or (layer4_outputs(4793));
    outputs(3035) <= layer4_outputs(2225);
    outputs(3036) <= not(layer4_outputs(6187));
    outputs(3037) <= (layer4_outputs(5986)) and (layer4_outputs(7538));
    outputs(3038) <= (layer4_outputs(2896)) and not (layer4_outputs(207));
    outputs(3039) <= layer4_outputs(2094);
    outputs(3040) <= layer4_outputs(7107);
    outputs(3041) <= not((layer4_outputs(3847)) and (layer4_outputs(1999)));
    outputs(3042) <= layer4_outputs(5);
    outputs(3043) <= not(layer4_outputs(1879));
    outputs(3044) <= not(layer4_outputs(2921));
    outputs(3045) <= layer4_outputs(3455);
    outputs(3046) <= not(layer4_outputs(5076));
    outputs(3047) <= not(layer4_outputs(7498)) or (layer4_outputs(6974));
    outputs(3048) <= layer4_outputs(5017);
    outputs(3049) <= layer4_outputs(6396);
    outputs(3050) <= not(layer4_outputs(7304));
    outputs(3051) <= layer4_outputs(2410);
    outputs(3052) <= not((layer4_outputs(5752)) xor (layer4_outputs(7040)));
    outputs(3053) <= not(layer4_outputs(4447));
    outputs(3054) <= not(layer4_outputs(6600));
    outputs(3055) <= (layer4_outputs(4056)) xor (layer4_outputs(2753));
    outputs(3056) <= not((layer4_outputs(890)) xor (layer4_outputs(5911)));
    outputs(3057) <= layer4_outputs(3287);
    outputs(3058) <= layer4_outputs(626);
    outputs(3059) <= layer4_outputs(2198);
    outputs(3060) <= layer4_outputs(5226);
    outputs(3061) <= (layer4_outputs(7645)) and not (layer4_outputs(1566));
    outputs(3062) <= (layer4_outputs(5864)) or (layer4_outputs(1645));
    outputs(3063) <= not((layer4_outputs(551)) xor (layer4_outputs(4399)));
    outputs(3064) <= (layer4_outputs(3528)) and (layer4_outputs(4556));
    outputs(3065) <= layer4_outputs(1852);
    outputs(3066) <= not(layer4_outputs(6277));
    outputs(3067) <= not(layer4_outputs(7322));
    outputs(3068) <= layer4_outputs(458);
    outputs(3069) <= layer4_outputs(6236);
    outputs(3070) <= (layer4_outputs(4214)) and (layer4_outputs(55));
    outputs(3071) <= layer4_outputs(1382);
    outputs(3072) <= (layer4_outputs(1403)) xor (layer4_outputs(2250));
    outputs(3073) <= layer4_outputs(5476);
    outputs(3074) <= not(layer4_outputs(5924));
    outputs(3075) <= layer4_outputs(5964);
    outputs(3076) <= layer4_outputs(3818);
    outputs(3077) <= layer4_outputs(1082);
    outputs(3078) <= layer4_outputs(7360);
    outputs(3079) <= (layer4_outputs(3122)) and (layer4_outputs(1850));
    outputs(3080) <= layer4_outputs(13);
    outputs(3081) <= (layer4_outputs(5447)) and (layer4_outputs(3038));
    outputs(3082) <= not(layer4_outputs(7424));
    outputs(3083) <= (layer4_outputs(1908)) xor (layer4_outputs(7036));
    outputs(3084) <= (layer4_outputs(2983)) and not (layer4_outputs(5975));
    outputs(3085) <= layer4_outputs(7085);
    outputs(3086) <= (layer4_outputs(6397)) and not (layer4_outputs(3479));
    outputs(3087) <= (layer4_outputs(784)) and not (layer4_outputs(1998));
    outputs(3088) <= (layer4_outputs(2414)) and not (layer4_outputs(5844));
    outputs(3089) <= (layer4_outputs(6991)) xor (layer4_outputs(2945));
    outputs(3090) <= not((layer4_outputs(185)) xor (layer4_outputs(3022)));
    outputs(3091) <= not(layer4_outputs(4795));
    outputs(3092) <= (layer4_outputs(7010)) xor (layer4_outputs(1673));
    outputs(3093) <= (layer4_outputs(5955)) and not (layer4_outputs(4246));
    outputs(3094) <= not(layer4_outputs(1955));
    outputs(3095) <= not((layer4_outputs(3688)) and (layer4_outputs(109)));
    outputs(3096) <= not((layer4_outputs(6499)) or (layer4_outputs(6343)));
    outputs(3097) <= (layer4_outputs(305)) xor (layer4_outputs(6965));
    outputs(3098) <= (layer4_outputs(3809)) xor (layer4_outputs(692));
    outputs(3099) <= layer4_outputs(4227);
    outputs(3100) <= (layer4_outputs(2711)) and not (layer4_outputs(5406));
    outputs(3101) <= layer4_outputs(1759);
    outputs(3102) <= (layer4_outputs(7053)) xor (layer4_outputs(6320));
    outputs(3103) <= not(layer4_outputs(3563));
    outputs(3104) <= not(layer4_outputs(3183));
    outputs(3105) <= (layer4_outputs(6216)) and (layer4_outputs(2759));
    outputs(3106) <= layer4_outputs(5984);
    outputs(3107) <= not((layer4_outputs(5147)) xor (layer4_outputs(4743)));
    outputs(3108) <= (layer4_outputs(6311)) and (layer4_outputs(1993));
    outputs(3109) <= not(layer4_outputs(7449));
    outputs(3110) <= not(layer4_outputs(1666)) or (layer4_outputs(2382));
    outputs(3111) <= layer4_outputs(6924);
    outputs(3112) <= layer4_outputs(1912);
    outputs(3113) <= layer4_outputs(6925);
    outputs(3114) <= not(layer4_outputs(2330));
    outputs(3115) <= (layer4_outputs(223)) xor (layer4_outputs(3001));
    outputs(3116) <= layer4_outputs(1391);
    outputs(3117) <= layer4_outputs(7186);
    outputs(3118) <= not(layer4_outputs(5581));
    outputs(3119) <= not((layer4_outputs(851)) or (layer4_outputs(693)));
    outputs(3120) <= layer4_outputs(1393);
    outputs(3121) <= (layer4_outputs(1586)) xor (layer4_outputs(870));
    outputs(3122) <= layer4_outputs(3176);
    outputs(3123) <= not(layer4_outputs(6339));
    outputs(3124) <= not(layer4_outputs(4970)) or (layer4_outputs(4288));
    outputs(3125) <= layer4_outputs(5540);
    outputs(3126) <= not((layer4_outputs(7466)) xor (layer4_outputs(677)));
    outputs(3127) <= layer4_outputs(1787);
    outputs(3128) <= not((layer4_outputs(3249)) xor (layer4_outputs(3948)));
    outputs(3129) <= not((layer4_outputs(451)) or (layer4_outputs(1106)));
    outputs(3130) <= not(layer4_outputs(5081)) or (layer4_outputs(4696));
    outputs(3131) <= not(layer4_outputs(4876));
    outputs(3132) <= (layer4_outputs(6186)) xor (layer4_outputs(6551));
    outputs(3133) <= not(layer4_outputs(6016));
    outputs(3134) <= layer4_outputs(7468);
    outputs(3135) <= not(layer4_outputs(3952));
    outputs(3136) <= layer4_outputs(2797);
    outputs(3137) <= not(layer4_outputs(893));
    outputs(3138) <= layer4_outputs(1993);
    outputs(3139) <= layer4_outputs(7112);
    outputs(3140) <= (layer4_outputs(1650)) xor (layer4_outputs(7276));
    outputs(3141) <= (layer4_outputs(5987)) and (layer4_outputs(2292));
    outputs(3142) <= not(layer4_outputs(6365)) or (layer4_outputs(5587));
    outputs(3143) <= not((layer4_outputs(5276)) xor (layer4_outputs(7060)));
    outputs(3144) <= not((layer4_outputs(247)) xor (layer4_outputs(1399)));
    outputs(3145) <= not((layer4_outputs(7376)) xor (layer4_outputs(1700)));
    outputs(3146) <= not(layer4_outputs(7597));
    outputs(3147) <= not(layer4_outputs(7259));
    outputs(3148) <= layer4_outputs(2874);
    outputs(3149) <= not(layer4_outputs(1915));
    outputs(3150) <= layer4_outputs(4434);
    outputs(3151) <= (layer4_outputs(3855)) and not (layer4_outputs(5718));
    outputs(3152) <= layer4_outputs(1190);
    outputs(3153) <= (layer4_outputs(4813)) and not (layer4_outputs(848));
    outputs(3154) <= layer4_outputs(180);
    outputs(3155) <= layer4_outputs(1532);
    outputs(3156) <= layer4_outputs(5842);
    outputs(3157) <= layer4_outputs(5653);
    outputs(3158) <= layer4_outputs(3730);
    outputs(3159) <= (layer4_outputs(6092)) and not (layer4_outputs(7324));
    outputs(3160) <= not(layer4_outputs(2756)) or (layer4_outputs(6747));
    outputs(3161) <= layer4_outputs(7649);
    outputs(3162) <= layer4_outputs(2006);
    outputs(3163) <= (layer4_outputs(1872)) or (layer4_outputs(2609));
    outputs(3164) <= not((layer4_outputs(4697)) xor (layer4_outputs(4641)));
    outputs(3165) <= (layer4_outputs(2994)) xor (layer4_outputs(6572));
    outputs(3166) <= not(layer4_outputs(3676));
    outputs(3167) <= not(layer4_outputs(7575));
    outputs(3168) <= (layer4_outputs(3068)) or (layer4_outputs(2644));
    outputs(3169) <= (layer4_outputs(7031)) xor (layer4_outputs(5880));
    outputs(3170) <= not(layer4_outputs(3058));
    outputs(3171) <= (layer4_outputs(534)) and (layer4_outputs(2100));
    outputs(3172) <= layer4_outputs(6605);
    outputs(3173) <= layer4_outputs(4229);
    outputs(3174) <= (layer4_outputs(5146)) and not (layer4_outputs(7100));
    outputs(3175) <= not(layer4_outputs(5549));
    outputs(3176) <= not((layer4_outputs(829)) or (layer4_outputs(4010)));
    outputs(3177) <= (layer4_outputs(7198)) and not (layer4_outputs(662));
    outputs(3178) <= not((layer4_outputs(731)) and (layer4_outputs(3624)));
    outputs(3179) <= layer4_outputs(945);
    outputs(3180) <= not(layer4_outputs(6888));
    outputs(3181) <= layer4_outputs(3636);
    outputs(3182) <= (layer4_outputs(254)) and (layer4_outputs(4583));
    outputs(3183) <= not(layer4_outputs(2260));
    outputs(3184) <= not((layer4_outputs(4889)) or (layer4_outputs(2857)));
    outputs(3185) <= not(layer4_outputs(3089));
    outputs(3186) <= (layer4_outputs(4884)) and not (layer4_outputs(5618));
    outputs(3187) <= not(layer4_outputs(775));
    outputs(3188) <= layer4_outputs(1455);
    outputs(3189) <= not((layer4_outputs(1128)) xor (layer4_outputs(2274)));
    outputs(3190) <= (layer4_outputs(6639)) and not (layer4_outputs(563));
    outputs(3191) <= layer4_outputs(4957);
    outputs(3192) <= not((layer4_outputs(5545)) or (layer4_outputs(6488)));
    outputs(3193) <= not(layer4_outputs(3388)) or (layer4_outputs(3711));
    outputs(3194) <= not(layer4_outputs(5268));
    outputs(3195) <= not(layer4_outputs(1405));
    outputs(3196) <= (layer4_outputs(5396)) xor (layer4_outputs(3089));
    outputs(3197) <= layer4_outputs(936);
    outputs(3198) <= layer4_outputs(1539);
    outputs(3199) <= not(layer4_outputs(3231));
    outputs(3200) <= not(layer4_outputs(2275));
    outputs(3201) <= not((layer4_outputs(134)) xor (layer4_outputs(5429)));
    outputs(3202) <= not(layer4_outputs(4651));
    outputs(3203) <= layer4_outputs(4147);
    outputs(3204) <= layer4_outputs(1216);
    outputs(3205) <= (layer4_outputs(1484)) and not (layer4_outputs(2087));
    outputs(3206) <= not((layer4_outputs(699)) xor (layer4_outputs(5810)));
    outputs(3207) <= (layer4_outputs(166)) xor (layer4_outputs(5950));
    outputs(3208) <= layer4_outputs(2166);
    outputs(3209) <= not(layer4_outputs(1599));
    outputs(3210) <= not((layer4_outputs(7539)) xor (layer4_outputs(708)));
    outputs(3211) <= layer4_outputs(2977);
    outputs(3212) <= not((layer4_outputs(5932)) xor (layer4_outputs(5305)));
    outputs(3213) <= (layer4_outputs(6313)) xor (layer4_outputs(7299));
    outputs(3214) <= (layer4_outputs(4230)) xor (layer4_outputs(1307));
    outputs(3215) <= not((layer4_outputs(5748)) xor (layer4_outputs(530)));
    outputs(3216) <= not((layer4_outputs(4174)) xor (layer4_outputs(3022)));
    outputs(3217) <= layer4_outputs(3278);
    outputs(3218) <= layer4_outputs(6474);
    outputs(3219) <= not(layer4_outputs(4403));
    outputs(3220) <= layer4_outputs(99);
    outputs(3221) <= (layer4_outputs(1753)) and (layer4_outputs(6681));
    outputs(3222) <= layer4_outputs(7077);
    outputs(3223) <= not(layer4_outputs(3587));
    outputs(3224) <= (layer4_outputs(2316)) xor (layer4_outputs(2520));
    outputs(3225) <= not((layer4_outputs(2143)) or (layer4_outputs(3911)));
    outputs(3226) <= not(layer4_outputs(741));
    outputs(3227) <= not(layer4_outputs(4486)) or (layer4_outputs(6753));
    outputs(3228) <= (layer4_outputs(4704)) and not (layer4_outputs(6376));
    outputs(3229) <= layer4_outputs(1139);
    outputs(3230) <= not(layer4_outputs(4619));
    outputs(3231) <= not(layer4_outputs(1529));
    outputs(3232) <= not(layer4_outputs(1166));
    outputs(3233) <= layer4_outputs(2149);
    outputs(3234) <= not(layer4_outputs(7037));
    outputs(3235) <= not((layer4_outputs(7487)) or (layer4_outputs(6364)));
    outputs(3236) <= not(layer4_outputs(158));
    outputs(3237) <= (layer4_outputs(4590)) xor (layer4_outputs(4407));
    outputs(3238) <= not(layer4_outputs(6270));
    outputs(3239) <= layer4_outputs(5591);
    outputs(3240) <= (layer4_outputs(6389)) or (layer4_outputs(2500));
    outputs(3241) <= not(layer4_outputs(4852));
    outputs(3242) <= not(layer4_outputs(3200));
    outputs(3243) <= not(layer4_outputs(5371));
    outputs(3244) <= layer4_outputs(2824);
    outputs(3245) <= not(layer4_outputs(3472));
    outputs(3246) <= not((layer4_outputs(1101)) or (layer4_outputs(898)));
    outputs(3247) <= (layer4_outputs(3719)) and (layer4_outputs(1880));
    outputs(3248) <= (layer4_outputs(1477)) and (layer4_outputs(5447));
    outputs(3249) <= not((layer4_outputs(1079)) xor (layer4_outputs(1191)));
    outputs(3250) <= layer4_outputs(2038);
    outputs(3251) <= not(layer4_outputs(5251)) or (layer4_outputs(1055));
    outputs(3252) <= (layer4_outputs(5996)) and not (layer4_outputs(5704));
    outputs(3253) <= layer4_outputs(638);
    outputs(3254) <= (layer4_outputs(7412)) or (layer4_outputs(3626));
    outputs(3255) <= layer4_outputs(6934);
    outputs(3256) <= (layer4_outputs(6677)) xor (layer4_outputs(6750));
    outputs(3257) <= not((layer4_outputs(2176)) xor (layer4_outputs(7484)));
    outputs(3258) <= layer4_outputs(2923);
    outputs(3259) <= not((layer4_outputs(2238)) xor (layer4_outputs(6028)));
    outputs(3260) <= not(layer4_outputs(7056));
    outputs(3261) <= layer4_outputs(1357);
    outputs(3262) <= layer4_outputs(1794);
    outputs(3263) <= layer4_outputs(3362);
    outputs(3264) <= (layer4_outputs(1751)) and not (layer4_outputs(1845));
    outputs(3265) <= layer4_outputs(4277);
    outputs(3266) <= not(layer4_outputs(202)) or (layer4_outputs(5036));
    outputs(3267) <= not(layer4_outputs(1609));
    outputs(3268) <= (layer4_outputs(1206)) and (layer4_outputs(6719));
    outputs(3269) <= (layer4_outputs(1607)) and not (layer4_outputs(7427));
    outputs(3270) <= not(layer4_outputs(2623));
    outputs(3271) <= (layer4_outputs(4454)) and (layer4_outputs(918));
    outputs(3272) <= not((layer4_outputs(4492)) and (layer4_outputs(4535)));
    outputs(3273) <= (layer4_outputs(325)) and (layer4_outputs(3673));
    outputs(3274) <= not(layer4_outputs(2925));
    outputs(3275) <= not((layer4_outputs(4403)) xor (layer4_outputs(2186)));
    outputs(3276) <= not(layer4_outputs(2661));
    outputs(3277) <= (layer4_outputs(1029)) and not (layer4_outputs(1862));
    outputs(3278) <= not(layer4_outputs(5841));
    outputs(3279) <= not((layer4_outputs(5501)) and (layer4_outputs(1306)));
    outputs(3280) <= not(layer4_outputs(6218)) or (layer4_outputs(2507));
    outputs(3281) <= layer4_outputs(7460);
    outputs(3282) <= not(layer4_outputs(775));
    outputs(3283) <= (layer4_outputs(370)) and (layer4_outputs(417));
    outputs(3284) <= not((layer4_outputs(1669)) or (layer4_outputs(6761)));
    outputs(3285) <= layer4_outputs(6566);
    outputs(3286) <= (layer4_outputs(2519)) or (layer4_outputs(3585));
    outputs(3287) <= layer4_outputs(5319);
    outputs(3288) <= layer4_outputs(912);
    outputs(3289) <= not(layer4_outputs(1328));
    outputs(3290) <= not(layer4_outputs(3786));
    outputs(3291) <= layer4_outputs(7616);
    outputs(3292) <= not(layer4_outputs(1507));
    outputs(3293) <= not(layer4_outputs(6603));
    outputs(3294) <= not(layer4_outputs(2096));
    outputs(3295) <= (layer4_outputs(4463)) or (layer4_outputs(6861));
    outputs(3296) <= not(layer4_outputs(6373));
    outputs(3297) <= not((layer4_outputs(1806)) xor (layer4_outputs(3495)));
    outputs(3298) <= layer4_outputs(3712);
    outputs(3299) <= not(layer4_outputs(2551));
    outputs(3300) <= not((layer4_outputs(2372)) and (layer4_outputs(2700)));
    outputs(3301) <= layer4_outputs(761);
    outputs(3302) <= layer4_outputs(7203);
    outputs(3303) <= (layer4_outputs(5405)) xor (layer4_outputs(257));
    outputs(3304) <= not((layer4_outputs(4300)) xor (layer4_outputs(7086)));
    outputs(3305) <= not(layer4_outputs(6462));
    outputs(3306) <= not(layer4_outputs(3439)) or (layer4_outputs(5791));
    outputs(3307) <= layer4_outputs(1109);
    outputs(3308) <= layer4_outputs(4278);
    outputs(3309) <= not((layer4_outputs(1158)) xor (layer4_outputs(5473)));
    outputs(3310) <= layer4_outputs(4424);
    outputs(3311) <= layer4_outputs(3673);
    outputs(3312) <= layer4_outputs(1678);
    outputs(3313) <= not(layer4_outputs(6376));
    outputs(3314) <= not(layer4_outputs(7317));
    outputs(3315) <= not((layer4_outputs(117)) xor (layer4_outputs(2015)));
    outputs(3316) <= layer4_outputs(6453);
    outputs(3317) <= (layer4_outputs(271)) xor (layer4_outputs(2870));
    outputs(3318) <= layer4_outputs(2012);
    outputs(3319) <= layer4_outputs(4073);
    outputs(3320) <= not(layer4_outputs(831));
    outputs(3321) <= (layer4_outputs(4647)) and not (layer4_outputs(6394));
    outputs(3322) <= not(layer4_outputs(6995));
    outputs(3323) <= layer4_outputs(692);
    outputs(3324) <= layer4_outputs(2977);
    outputs(3325) <= not(layer4_outputs(711));
    outputs(3326) <= not(layer4_outputs(431));
    outputs(3327) <= (layer4_outputs(4720)) and not (layer4_outputs(3728));
    outputs(3328) <= layer4_outputs(1623);
    outputs(3329) <= (layer4_outputs(5836)) and not (layer4_outputs(2600));
    outputs(3330) <= layer4_outputs(4282);
    outputs(3331) <= layer4_outputs(4503);
    outputs(3332) <= (layer4_outputs(3939)) xor (layer4_outputs(6695));
    outputs(3333) <= layer4_outputs(879);
    outputs(3334) <= not(layer4_outputs(5107));
    outputs(3335) <= not((layer4_outputs(6578)) or (layer4_outputs(7398)));
    outputs(3336) <= layer4_outputs(7167);
    outputs(3337) <= layer4_outputs(155);
    outputs(3338) <= not(layer4_outputs(4582));
    outputs(3339) <= layer4_outputs(7623);
    outputs(3340) <= layer4_outputs(1721);
    outputs(3341) <= not(layer4_outputs(2081));
    outputs(3342) <= not(layer4_outputs(1828));
    outputs(3343) <= not(layer4_outputs(5100));
    outputs(3344) <= not((layer4_outputs(3539)) xor (layer4_outputs(5988)));
    outputs(3345) <= not(layer4_outputs(6415));
    outputs(3346) <= not(layer4_outputs(7237));
    outputs(3347) <= (layer4_outputs(5899)) xor (layer4_outputs(6573));
    outputs(3348) <= (layer4_outputs(707)) and (layer4_outputs(633));
    outputs(3349) <= not(layer4_outputs(4326));
    outputs(3350) <= layer4_outputs(1360);
    outputs(3351) <= not(layer4_outputs(1439));
    outputs(3352) <= not(layer4_outputs(4845));
    outputs(3353) <= layer4_outputs(994);
    outputs(3354) <= (layer4_outputs(6566)) xor (layer4_outputs(7503));
    outputs(3355) <= not(layer4_outputs(1080));
    outputs(3356) <= layer4_outputs(4629);
    outputs(3357) <= (layer4_outputs(6585)) or (layer4_outputs(488));
    outputs(3358) <= not((layer4_outputs(7607)) xor (layer4_outputs(1942)));
    outputs(3359) <= not((layer4_outputs(562)) xor (layer4_outputs(6232)));
    outputs(3360) <= (layer4_outputs(4476)) or (layer4_outputs(3201));
    outputs(3361) <= (layer4_outputs(517)) and not (layer4_outputs(2535));
    outputs(3362) <= layer4_outputs(5479);
    outputs(3363) <= not(layer4_outputs(4319)) or (layer4_outputs(7402));
    outputs(3364) <= layer4_outputs(971);
    outputs(3365) <= not(layer4_outputs(5437));
    outputs(3366) <= layer4_outputs(7158);
    outputs(3367) <= not(layer4_outputs(3739));
    outputs(3368) <= (layer4_outputs(5142)) and not (layer4_outputs(2218));
    outputs(3369) <= not(layer4_outputs(7415));
    outputs(3370) <= (layer4_outputs(4858)) and not (layer4_outputs(6837));
    outputs(3371) <= layer4_outputs(2292);
    outputs(3372) <= layer4_outputs(1061);
    outputs(3373) <= not(layer4_outputs(1609));
    outputs(3374) <= (layer4_outputs(2124)) and (layer4_outputs(6546));
    outputs(3375) <= not(layer4_outputs(4418));
    outputs(3376) <= layer4_outputs(3255);
    outputs(3377) <= not((layer4_outputs(4271)) xor (layer4_outputs(3017)));
    outputs(3378) <= not(layer4_outputs(4691)) or (layer4_outputs(7604));
    outputs(3379) <= (layer4_outputs(1830)) and not (layer4_outputs(2091));
    outputs(3380) <= not(layer4_outputs(3932)) or (layer4_outputs(1104));
    outputs(3381) <= not(layer4_outputs(451));
    outputs(3382) <= not((layer4_outputs(4396)) xor (layer4_outputs(3430)));
    outputs(3383) <= not(layer4_outputs(2251)) or (layer4_outputs(7297));
    outputs(3384) <= (layer4_outputs(3395)) and (layer4_outputs(7528));
    outputs(3385) <= layer4_outputs(6437);
    outputs(3386) <= layer4_outputs(7243);
    outputs(3387) <= layer4_outputs(108);
    outputs(3388) <= not(layer4_outputs(5430));
    outputs(3389) <= (layer4_outputs(529)) and not (layer4_outputs(2248));
    outputs(3390) <= not(layer4_outputs(3548));
    outputs(3391) <= not((layer4_outputs(1166)) xor (layer4_outputs(7282)));
    outputs(3392) <= not((layer4_outputs(1399)) and (layer4_outputs(1809)));
    outputs(3393) <= layer4_outputs(6193);
    outputs(3394) <= (layer4_outputs(4771)) and (layer4_outputs(376));
    outputs(3395) <= not(layer4_outputs(2982));
    outputs(3396) <= not(layer4_outputs(1429));
    outputs(3397) <= not(layer4_outputs(2897));
    outputs(3398) <= not(layer4_outputs(7064));
    outputs(3399) <= layer4_outputs(4166);
    outputs(3400) <= not(layer4_outputs(6451));
    outputs(3401) <= (layer4_outputs(3149)) and (layer4_outputs(890));
    outputs(3402) <= not(layer4_outputs(6708));
    outputs(3403) <= (layer4_outputs(1167)) xor (layer4_outputs(684));
    outputs(3404) <= not(layer4_outputs(7523));
    outputs(3405) <= (layer4_outputs(1634)) or (layer4_outputs(7368));
    outputs(3406) <= layer4_outputs(5427);
    outputs(3407) <= (layer4_outputs(2974)) xor (layer4_outputs(5280));
    outputs(3408) <= not(layer4_outputs(4857));
    outputs(3409) <= not((layer4_outputs(2471)) xor (layer4_outputs(4312)));
    outputs(3410) <= (layer4_outputs(637)) and not (layer4_outputs(2871));
    outputs(3411) <= (layer4_outputs(337)) and (layer4_outputs(1289));
    outputs(3412) <= not(layer4_outputs(5122));
    outputs(3413) <= layer4_outputs(4398);
    outputs(3414) <= layer4_outputs(5921);
    outputs(3415) <= layer4_outputs(6604);
    outputs(3416) <= not(layer4_outputs(737));
    outputs(3417) <= layer4_outputs(5805);
    outputs(3418) <= not((layer4_outputs(5441)) or (layer4_outputs(7337)));
    outputs(3419) <= layer4_outputs(3204);
    outputs(3420) <= not((layer4_outputs(3467)) xor (layer4_outputs(4948)));
    outputs(3421) <= not(layer4_outputs(4732));
    outputs(3422) <= not((layer4_outputs(6595)) xor (layer4_outputs(4138)));
    outputs(3423) <= layer4_outputs(345);
    outputs(3424) <= not(layer4_outputs(1551));
    outputs(3425) <= layer4_outputs(2951);
    outputs(3426) <= not(layer4_outputs(7310));
    outputs(3427) <= (layer4_outputs(4091)) and (layer4_outputs(2302));
    outputs(3428) <= layer4_outputs(4241);
    outputs(3429) <= not(layer4_outputs(5514));
    outputs(3430) <= layer4_outputs(6740);
    outputs(3431) <= not(layer4_outputs(549));
    outputs(3432) <= not(layer4_outputs(7666));
    outputs(3433) <= layer4_outputs(302);
    outputs(3434) <= not(layer4_outputs(1137));
    outputs(3435) <= layer4_outputs(40);
    outputs(3436) <= not(layer4_outputs(3253));
    outputs(3437) <= not(layer4_outputs(4654));
    outputs(3438) <= not((layer4_outputs(356)) and (layer4_outputs(1489)));
    outputs(3439) <= not((layer4_outputs(4182)) xor (layer4_outputs(3473)));
    outputs(3440) <= not((layer4_outputs(1690)) xor (layer4_outputs(4669)));
    outputs(3441) <= layer4_outputs(4704);
    outputs(3442) <= not(layer4_outputs(5088));
    outputs(3443) <= layer4_outputs(7516);
    outputs(3444) <= layer4_outputs(2991);
    outputs(3445) <= not(layer4_outputs(4850));
    outputs(3446) <= not(layer4_outputs(5813));
    outputs(3447) <= (layer4_outputs(2322)) or (layer4_outputs(594));
    outputs(3448) <= (layer4_outputs(1808)) and not (layer4_outputs(6225));
    outputs(3449) <= not((layer4_outputs(2153)) xor (layer4_outputs(3139)));
    outputs(3450) <= not((layer4_outputs(5311)) or (layer4_outputs(2957)));
    outputs(3451) <= not((layer4_outputs(2880)) xor (layer4_outputs(1160)));
    outputs(3452) <= layer4_outputs(4927);
    outputs(3453) <= layer4_outputs(5764);
    outputs(3454) <= not((layer4_outputs(4089)) xor (layer4_outputs(1371)));
    outputs(3455) <= (layer4_outputs(3966)) xor (layer4_outputs(1263));
    outputs(3456) <= layer4_outputs(2727);
    outputs(3457) <= (layer4_outputs(7078)) and (layer4_outputs(6276));
    outputs(3458) <= not(layer4_outputs(1588));
    outputs(3459) <= (layer4_outputs(4338)) and (layer4_outputs(6330));
    outputs(3460) <= not(layer4_outputs(595));
    outputs(3461) <= not((layer4_outputs(1812)) xor (layer4_outputs(2043)));
    outputs(3462) <= not(layer4_outputs(1697));
    outputs(3463) <= layer4_outputs(4273);
    outputs(3464) <= not((layer4_outputs(6521)) xor (layer4_outputs(6851)));
    outputs(3465) <= (layer4_outputs(3075)) and not (layer4_outputs(1552));
    outputs(3466) <= not((layer4_outputs(1803)) xor (layer4_outputs(1108)));
    outputs(3467) <= (layer4_outputs(4554)) and (layer4_outputs(6476));
    outputs(3468) <= not((layer4_outputs(4575)) and (layer4_outputs(1916)));
    outputs(3469) <= (layer4_outputs(222)) and not (layer4_outputs(5037));
    outputs(3470) <= layer4_outputs(3909);
    outputs(3471) <= not(layer4_outputs(5003));
    outputs(3472) <= layer4_outputs(4238);
    outputs(3473) <= not(layer4_outputs(7647)) or (layer4_outputs(4854));
    outputs(3474) <= (layer4_outputs(4508)) and (layer4_outputs(1918));
    outputs(3475) <= layer4_outputs(923);
    outputs(3476) <= not(layer4_outputs(2537));
    outputs(3477) <= not(layer4_outputs(1873)) or (layer4_outputs(368));
    outputs(3478) <= layer4_outputs(7221);
    outputs(3479) <= not(layer4_outputs(5194));
    outputs(3480) <= (layer4_outputs(6311)) xor (layer4_outputs(1857));
    outputs(3481) <= not((layer4_outputs(2528)) xor (layer4_outputs(4104)));
    outputs(3482) <= (layer4_outputs(2828)) and not (layer4_outputs(190));
    outputs(3483) <= layer4_outputs(801);
    outputs(3484) <= not(layer4_outputs(6314)) or (layer4_outputs(3374));
    outputs(3485) <= not(layer4_outputs(1111));
    outputs(3486) <= layer4_outputs(6699);
    outputs(3487) <= (layer4_outputs(3613)) and not (layer4_outputs(1103));
    outputs(3488) <= not((layer4_outputs(195)) xor (layer4_outputs(6684)));
    outputs(3489) <= not((layer4_outputs(546)) xor (layer4_outputs(289)));
    outputs(3490) <= not(layer4_outputs(1243));
    outputs(3491) <= (layer4_outputs(67)) and (layer4_outputs(6405));
    outputs(3492) <= layer4_outputs(3901);
    outputs(3493) <= (layer4_outputs(204)) xor (layer4_outputs(4590));
    outputs(3494) <= not(layer4_outputs(6268));
    outputs(3495) <= layer4_outputs(827);
    outputs(3496) <= layer4_outputs(305);
    outputs(3497) <= not(layer4_outputs(3627));
    outputs(3498) <= not((layer4_outputs(2347)) xor (layer4_outputs(4677)));
    outputs(3499) <= not((layer4_outputs(1857)) or (layer4_outputs(4900)));
    outputs(3500) <= layer4_outputs(22);
    outputs(3501) <= layer4_outputs(1443);
    outputs(3502) <= not(layer4_outputs(1632));
    outputs(3503) <= layer4_outputs(3928);
    outputs(3504) <= not(layer4_outputs(260));
    outputs(3505) <= (layer4_outputs(4473)) and (layer4_outputs(3508));
    outputs(3506) <= not(layer4_outputs(3074));
    outputs(3507) <= not(layer4_outputs(6560)) or (layer4_outputs(2329));
    outputs(3508) <= not((layer4_outputs(899)) or (layer4_outputs(7065)));
    outputs(3509) <= layer4_outputs(340);
    outputs(3510) <= layer4_outputs(5760);
    outputs(3511) <= not((layer4_outputs(4607)) or (layer4_outputs(6525)));
    outputs(3512) <= layer4_outputs(1171);
    outputs(3513) <= layer4_outputs(2149);
    outputs(3514) <= (layer4_outputs(57)) and (layer4_outputs(3000));
    outputs(3515) <= not(layer4_outputs(3118));
    outputs(3516) <= layer4_outputs(40);
    outputs(3517) <= (layer4_outputs(7515)) and not (layer4_outputs(6109));
    outputs(3518) <= (layer4_outputs(4356)) and (layer4_outputs(6847));
    outputs(3519) <= not(layer4_outputs(5172));
    outputs(3520) <= not((layer4_outputs(3450)) xor (layer4_outputs(1123)));
    outputs(3521) <= layer4_outputs(6818);
    outputs(3522) <= not((layer4_outputs(7446)) and (layer4_outputs(3505)));
    outputs(3523) <= not(layer4_outputs(478));
    outputs(3524) <= not(layer4_outputs(590));
    outputs(3525) <= (layer4_outputs(5735)) and not (layer4_outputs(164));
    outputs(3526) <= not(layer4_outputs(289));
    outputs(3527) <= not(layer4_outputs(6353));
    outputs(3528) <= layer4_outputs(872);
    outputs(3529) <= layer4_outputs(6858);
    outputs(3530) <= not(layer4_outputs(6967));
    outputs(3531) <= (layer4_outputs(5499)) and not (layer4_outputs(1024));
    outputs(3532) <= layer4_outputs(5261);
    outputs(3533) <= not(layer4_outputs(2744));
    outputs(3534) <= not(layer4_outputs(7565));
    outputs(3535) <= (layer4_outputs(5333)) and (layer4_outputs(2990));
    outputs(3536) <= layer4_outputs(4530);
    outputs(3537) <= layer4_outputs(125);
    outputs(3538) <= layer4_outputs(4591);
    outputs(3539) <= layer4_outputs(3808);
    outputs(3540) <= layer4_outputs(1209);
    outputs(3541) <= not(layer4_outputs(5210)) or (layer4_outputs(149));
    outputs(3542) <= layer4_outputs(4779);
    outputs(3543) <= layer4_outputs(756);
    outputs(3544) <= not(layer4_outputs(4753));
    outputs(3545) <= not(layer4_outputs(3297));
    outputs(3546) <= not((layer4_outputs(7095)) xor (layer4_outputs(4171)));
    outputs(3547) <= not(layer4_outputs(23));
    outputs(3548) <= (layer4_outputs(3988)) and not (layer4_outputs(1891));
    outputs(3549) <= not(layer4_outputs(5638));
    outputs(3550) <= not(layer4_outputs(7639));
    outputs(3551) <= not((layer4_outputs(1961)) or (layer4_outputs(5095)));
    outputs(3552) <= layer4_outputs(4084);
    outputs(3553) <= layer4_outputs(317);
    outputs(3554) <= not(layer4_outputs(693));
    outputs(3555) <= (layer4_outputs(1156)) xor (layer4_outputs(4797));
    outputs(3556) <= (layer4_outputs(7124)) xor (layer4_outputs(2162));
    outputs(3557) <= not((layer4_outputs(6365)) or (layer4_outputs(3991)));
    outputs(3558) <= (layer4_outputs(2397)) or (layer4_outputs(3320));
    outputs(3559) <= layer4_outputs(3890);
    outputs(3560) <= layer4_outputs(6638);
    outputs(3561) <= (layer4_outputs(407)) and not (layer4_outputs(763));
    outputs(3562) <= layer4_outputs(2834);
    outputs(3563) <= (layer4_outputs(7245)) and not (layer4_outputs(6782));
    outputs(3564) <= not(layer4_outputs(1017));
    outputs(3565) <= not(layer4_outputs(3571));
    outputs(3566) <= not(layer4_outputs(5474));
    outputs(3567) <= not(layer4_outputs(3550));
    outputs(3568) <= (layer4_outputs(6014)) and not (layer4_outputs(7316));
    outputs(3569) <= not(layer4_outputs(4795));
    outputs(3570) <= not((layer4_outputs(952)) xor (layer4_outputs(3554)));
    outputs(3571) <= not(layer4_outputs(18));
    outputs(3572) <= (layer4_outputs(5969)) and (layer4_outputs(1068));
    outputs(3573) <= (layer4_outputs(6420)) or (layer4_outputs(7266));
    outputs(3574) <= not((layer4_outputs(6180)) xor (layer4_outputs(1971)));
    outputs(3575) <= not(layer4_outputs(2416));
    outputs(3576) <= not(layer4_outputs(6469)) or (layer4_outputs(6152));
    outputs(3577) <= layer4_outputs(6074);
    outputs(3578) <= not(layer4_outputs(3879));
    outputs(3579) <= not(layer4_outputs(1601));
    outputs(3580) <= not(layer4_outputs(6430)) or (layer4_outputs(5721));
    outputs(3581) <= layer4_outputs(3591);
    outputs(3582) <= not(layer4_outputs(3143));
    outputs(3583) <= layer4_outputs(4765);
    outputs(3584) <= (layer4_outputs(4109)) and (layer4_outputs(5318));
    outputs(3585) <= not(layer4_outputs(1881));
    outputs(3586) <= not(layer4_outputs(3231));
    outputs(3587) <= not(layer4_outputs(6055));
    outputs(3588) <= (layer4_outputs(6880)) xor (layer4_outputs(216));
    outputs(3589) <= layer4_outputs(3172);
    outputs(3590) <= (layer4_outputs(1954)) and (layer4_outputs(7534));
    outputs(3591) <= (layer4_outputs(5573)) or (layer4_outputs(3890));
    outputs(3592) <= not(layer4_outputs(3824));
    outputs(3593) <= layer4_outputs(973);
    outputs(3594) <= not(layer4_outputs(6564));
    outputs(3595) <= not(layer4_outputs(837));
    outputs(3596) <= layer4_outputs(1495);
    outputs(3597) <= layer4_outputs(5380);
    outputs(3598) <= (layer4_outputs(502)) and not (layer4_outputs(1364));
    outputs(3599) <= not(layer4_outputs(5616));
    outputs(3600) <= (layer4_outputs(2665)) xor (layer4_outputs(3305));
    outputs(3601) <= layer4_outputs(6224);
    outputs(3602) <= not(layer4_outputs(2108));
    outputs(3603) <= not(layer4_outputs(5627));
    outputs(3604) <= not(layer4_outputs(1342));
    outputs(3605) <= layer4_outputs(697);
    outputs(3606) <= layer4_outputs(2552);
    outputs(3607) <= layer4_outputs(866);
    outputs(3608) <= layer4_outputs(4586);
    outputs(3609) <= (layer4_outputs(865)) and (layer4_outputs(221));
    outputs(3610) <= not((layer4_outputs(7249)) or (layer4_outputs(3311)));
    outputs(3611) <= not((layer4_outputs(1935)) or (layer4_outputs(1330)));
    outputs(3612) <= (layer4_outputs(3591)) and not (layer4_outputs(3598));
    outputs(3613) <= (layer4_outputs(2465)) xor (layer4_outputs(6946));
    outputs(3614) <= layer4_outputs(5991);
    outputs(3615) <= not(layer4_outputs(1829));
    outputs(3616) <= not((layer4_outputs(1066)) xor (layer4_outputs(1814)));
    outputs(3617) <= layer4_outputs(3417);
    outputs(3618) <= not(layer4_outputs(4150));
    outputs(3619) <= not(layer4_outputs(5115));
    outputs(3620) <= (layer4_outputs(480)) and not (layer4_outputs(6620));
    outputs(3621) <= not(layer4_outputs(5577));
    outputs(3622) <= not(layer4_outputs(4394));
    outputs(3623) <= (layer4_outputs(4603)) and (layer4_outputs(1475));
    outputs(3624) <= layer4_outputs(6965);
    outputs(3625) <= not((layer4_outputs(4151)) xor (layer4_outputs(3608)));
    outputs(3626) <= layer4_outputs(4063);
    outputs(3627) <= (layer4_outputs(2759)) and (layer4_outputs(3024));
    outputs(3628) <= layer4_outputs(4258);
    outputs(3629) <= (layer4_outputs(3356)) xor (layer4_outputs(1210));
    outputs(3630) <= layer4_outputs(7468);
    outputs(3631) <= not(layer4_outputs(7242));
    outputs(3632) <= (layer4_outputs(5281)) xor (layer4_outputs(3209));
    outputs(3633) <= layer4_outputs(7114);
    outputs(3634) <= (layer4_outputs(5018)) and not (layer4_outputs(6052));
    outputs(3635) <= layer4_outputs(3573);
    outputs(3636) <= layer4_outputs(5603);
    outputs(3637) <= (layer4_outputs(4775)) xor (layer4_outputs(4287));
    outputs(3638) <= layer4_outputs(6533);
    outputs(3639) <= not((layer4_outputs(2458)) xor (layer4_outputs(167)));
    outputs(3640) <= not(layer4_outputs(1972));
    outputs(3641) <= not((layer4_outputs(1371)) xor (layer4_outputs(3730)));
    outputs(3642) <= not(layer4_outputs(5347));
    outputs(3643) <= layer4_outputs(3845);
    outputs(3644) <= not((layer4_outputs(2293)) or (layer4_outputs(1027)));
    outputs(3645) <= not(layer4_outputs(5768));
    outputs(3646) <= layer4_outputs(6559);
    outputs(3647) <= (layer4_outputs(5142)) and not (layer4_outputs(6378));
    outputs(3648) <= layer4_outputs(5886);
    outputs(3649) <= layer4_outputs(3758);
    outputs(3650) <= not(layer4_outputs(4921));
    outputs(3651) <= (layer4_outputs(6059)) xor (layer4_outputs(1796));
    outputs(3652) <= not(layer4_outputs(7408));
    outputs(3653) <= (layer4_outputs(5758)) xor (layer4_outputs(1752));
    outputs(3654) <= not(layer4_outputs(2629));
    outputs(3655) <= not(layer4_outputs(5640));
    outputs(3656) <= layer4_outputs(980);
    outputs(3657) <= (layer4_outputs(5119)) and (layer4_outputs(1035));
    outputs(3658) <= (layer4_outputs(7321)) and not (layer4_outputs(6835));
    outputs(3659) <= (layer4_outputs(911)) xor (layer4_outputs(3384));
    outputs(3660) <= not(layer4_outputs(6548));
    outputs(3661) <= not((layer4_outputs(1377)) or (layer4_outputs(5320)));
    outputs(3662) <= (layer4_outputs(6973)) xor (layer4_outputs(6224));
    outputs(3663) <= not(layer4_outputs(885));
    outputs(3664) <= not(layer4_outputs(7028)) or (layer4_outputs(6441));
    outputs(3665) <= layer4_outputs(3079);
    outputs(3666) <= (layer4_outputs(607)) and (layer4_outputs(7098));
    outputs(3667) <= (layer4_outputs(2115)) and not (layer4_outputs(6399));
    outputs(3668) <= layer4_outputs(4201);
    outputs(3669) <= (layer4_outputs(6229)) and (layer4_outputs(5653));
    outputs(3670) <= not((layer4_outputs(134)) or (layer4_outputs(5277)));
    outputs(3671) <= layer4_outputs(7302);
    outputs(3672) <= not(layer4_outputs(5166));
    outputs(3673) <= (layer4_outputs(2605)) xor (layer4_outputs(6398));
    outputs(3674) <= layer4_outputs(3595);
    outputs(3675) <= layer4_outputs(4945);
    outputs(3676) <= layer4_outputs(2686);
    outputs(3677) <= not(layer4_outputs(1404));
    outputs(3678) <= (layer4_outputs(6309)) and (layer4_outputs(2212));
    outputs(3679) <= layer4_outputs(285);
    outputs(3680) <= layer4_outputs(6148);
    outputs(3681) <= not(layer4_outputs(541));
    outputs(3682) <= layer4_outputs(250);
    outputs(3683) <= not(layer4_outputs(596));
    outputs(3684) <= not(layer4_outputs(2361));
    outputs(3685) <= (layer4_outputs(4714)) and (layer4_outputs(676));
    outputs(3686) <= not(layer4_outputs(5665));
    outputs(3687) <= not((layer4_outputs(5062)) xor (layer4_outputs(1988)));
    outputs(3688) <= not(layer4_outputs(4627));
    outputs(3689) <= (layer4_outputs(4222)) xor (layer4_outputs(2241));
    outputs(3690) <= not((layer4_outputs(1286)) xor (layer4_outputs(2076)));
    outputs(3691) <= layer4_outputs(1116);
    outputs(3692) <= not((layer4_outputs(5051)) xor (layer4_outputs(1521)));
    outputs(3693) <= not(layer4_outputs(1670));
    outputs(3694) <= not(layer4_outputs(3262));
    outputs(3695) <= layer4_outputs(3835);
    outputs(3696) <= layer4_outputs(4578);
    outputs(3697) <= layer4_outputs(4534);
    outputs(3698) <= (layer4_outputs(7535)) and (layer4_outputs(1743));
    outputs(3699) <= layer4_outputs(4066);
    outputs(3700) <= (layer4_outputs(1901)) and (layer4_outputs(2258));
    outputs(3701) <= not(layer4_outputs(6621));
    outputs(3702) <= (layer4_outputs(3057)) and not (layer4_outputs(5130));
    outputs(3703) <= (layer4_outputs(371)) xor (layer4_outputs(170));
    outputs(3704) <= not(layer4_outputs(4608));
    outputs(3705) <= (layer4_outputs(3693)) and not (layer4_outputs(1529));
    outputs(3706) <= not((layer4_outputs(2587)) or (layer4_outputs(2694)));
    outputs(3707) <= (layer4_outputs(2688)) and (layer4_outputs(2349));
    outputs(3708) <= not(layer4_outputs(24)) or (layer4_outputs(3814));
    outputs(3709) <= not(layer4_outputs(7385));
    outputs(3710) <= (layer4_outputs(1352)) and not (layer4_outputs(293));
    outputs(3711) <= layer4_outputs(1407);
    outputs(3712) <= not(layer4_outputs(1952));
    outputs(3713) <= (layer4_outputs(5152)) and not (layer4_outputs(7122));
    outputs(3714) <= layer4_outputs(4805);
    outputs(3715) <= not(layer4_outputs(4626));
    outputs(3716) <= layer4_outputs(878);
    outputs(3717) <= not(layer4_outputs(5643));
    outputs(3718) <= not(layer4_outputs(3016));
    outputs(3719) <= layer4_outputs(3643);
    outputs(3720) <= layer4_outputs(2249);
    outputs(3721) <= not(layer4_outputs(5555)) or (layer4_outputs(4225));
    outputs(3722) <= not((layer4_outputs(688)) or (layer4_outputs(6499)));
    outputs(3723) <= layer4_outputs(3719);
    outputs(3724) <= layer4_outputs(4041);
    outputs(3725) <= layer4_outputs(1587);
    outputs(3726) <= layer4_outputs(1859);
    outputs(3727) <= layer4_outputs(5699);
    outputs(3728) <= layer4_outputs(4840);
    outputs(3729) <= not(layer4_outputs(4801)) or (layer4_outputs(7491));
    outputs(3730) <= layer4_outputs(6479);
    outputs(3731) <= layer4_outputs(7610);
    outputs(3732) <= not((layer4_outputs(6903)) xor (layer4_outputs(1568)));
    outputs(3733) <= layer4_outputs(609);
    outputs(3734) <= (layer4_outputs(6253)) or (layer4_outputs(6190));
    outputs(3735) <= layer4_outputs(490);
    outputs(3736) <= (layer4_outputs(7157)) and not (layer4_outputs(6910));
    outputs(3737) <= not(layer4_outputs(588));
    outputs(3738) <= (layer4_outputs(1780)) or (layer4_outputs(1720));
    outputs(3739) <= layer4_outputs(7431);
    outputs(3740) <= (layer4_outputs(5909)) and (layer4_outputs(628));
    outputs(3741) <= layer4_outputs(7382);
    outputs(3742) <= not(layer4_outputs(2132)) or (layer4_outputs(1978));
    outputs(3743) <= layer4_outputs(5084);
    outputs(3744) <= (layer4_outputs(4436)) and not (layer4_outputs(4752));
    outputs(3745) <= (layer4_outputs(2456)) xor (layer4_outputs(7505));
    outputs(3746) <= not(layer4_outputs(3164));
    outputs(3747) <= not(layer4_outputs(4450));
    outputs(3748) <= (layer4_outputs(6304)) and not (layer4_outputs(2016));
    outputs(3749) <= not(layer4_outputs(2612));
    outputs(3750) <= not(layer4_outputs(3150));
    outputs(3751) <= (layer4_outputs(4190)) and not (layer4_outputs(7441));
    outputs(3752) <= layer4_outputs(1628);
    outputs(3753) <= layer4_outputs(4830);
    outputs(3754) <= layer4_outputs(53);
    outputs(3755) <= not(layer4_outputs(1933));
    outputs(3756) <= (layer4_outputs(1841)) xor (layer4_outputs(1747));
    outputs(3757) <= (layer4_outputs(3168)) and (layer4_outputs(5484));
    outputs(3758) <= not((layer4_outputs(5681)) xor (layer4_outputs(63)));
    outputs(3759) <= (layer4_outputs(6553)) xor (layer4_outputs(65));
    outputs(3760) <= not(layer4_outputs(526));
    outputs(3761) <= layer4_outputs(4932);
    outputs(3762) <= (layer4_outputs(7105)) and (layer4_outputs(3982));
    outputs(3763) <= (layer4_outputs(4091)) and not (layer4_outputs(4900));
    outputs(3764) <= not((layer4_outputs(4877)) or (layer4_outputs(6923)));
    outputs(3765) <= layer4_outputs(3442);
    outputs(3766) <= not(layer4_outputs(4925)) or (layer4_outputs(2570));
    outputs(3767) <= layer4_outputs(228);
    outputs(3768) <= not((layer4_outputs(629)) xor (layer4_outputs(4243)));
    outputs(3769) <= (layer4_outputs(4574)) xor (layer4_outputs(3896));
    outputs(3770) <= not((layer4_outputs(6689)) xor (layer4_outputs(7308)));
    outputs(3771) <= not(layer4_outputs(5784));
    outputs(3772) <= not(layer4_outputs(156));
    outputs(3773) <= not((layer4_outputs(4552)) xor (layer4_outputs(5331)));
    outputs(3774) <= (layer4_outputs(766)) and (layer4_outputs(3489));
    outputs(3775) <= layer4_outputs(2285);
    outputs(3776) <= (layer4_outputs(4462)) and (layer4_outputs(7058));
    outputs(3777) <= layer4_outputs(638);
    outputs(3778) <= not(layer4_outputs(566));
    outputs(3779) <= (layer4_outputs(3498)) xor (layer4_outputs(2063));
    outputs(3780) <= layer4_outputs(828);
    outputs(3781) <= layer4_outputs(2727);
    outputs(3782) <= not((layer4_outputs(522)) xor (layer4_outputs(500)));
    outputs(3783) <= (layer4_outputs(6976)) xor (layer4_outputs(7069));
    outputs(3784) <= not(layer4_outputs(5072)) or (layer4_outputs(2963));
    outputs(3785) <= layer4_outputs(697);
    outputs(3786) <= layer4_outputs(5921);
    outputs(3787) <= not(layer4_outputs(2674));
    outputs(3788) <= layer4_outputs(2601);
    outputs(3789) <= layer4_outputs(1190);
    outputs(3790) <= not((layer4_outputs(1950)) and (layer4_outputs(3029)));
    outputs(3791) <= layer4_outputs(3011);
    outputs(3792) <= layer4_outputs(1001);
    outputs(3793) <= (layer4_outputs(6676)) xor (layer4_outputs(430));
    outputs(3794) <= layer4_outputs(4898);
    outputs(3795) <= not(layer4_outputs(5080));
    outputs(3796) <= not(layer4_outputs(45));
    outputs(3797) <= not((layer4_outputs(1729)) or (layer4_outputs(4498)));
    outputs(3798) <= layer4_outputs(2036);
    outputs(3799) <= not((layer4_outputs(4874)) xor (layer4_outputs(1406)));
    outputs(3800) <= layer4_outputs(5075);
    outputs(3801) <= not(layer4_outputs(3274));
    outputs(3802) <= layer4_outputs(5314);
    outputs(3803) <= not(layer4_outputs(1238));
    outputs(3804) <= not(layer4_outputs(4068));
    outputs(3805) <= not(layer4_outputs(147));
    outputs(3806) <= layer4_outputs(5985);
    outputs(3807) <= not(layer4_outputs(509));
    outputs(3808) <= layer4_outputs(3344);
    outputs(3809) <= layer4_outputs(4581);
    outputs(3810) <= not(layer4_outputs(2760));
    outputs(3811) <= not((layer4_outputs(3051)) or (layer4_outputs(6679)));
    outputs(3812) <= not((layer4_outputs(5915)) xor (layer4_outputs(2737)));
    outputs(3813) <= (layer4_outputs(5508)) and not (layer4_outputs(5712));
    outputs(3814) <= (layer4_outputs(929)) and (layer4_outputs(766));
    outputs(3815) <= (layer4_outputs(5480)) xor (layer4_outputs(5175));
    outputs(3816) <= (layer4_outputs(1621)) xor (layer4_outputs(1366));
    outputs(3817) <= not(layer4_outputs(1530));
    outputs(3818) <= not(layer4_outputs(5209));
    outputs(3819) <= not(layer4_outputs(3108));
    outputs(3820) <= layer4_outputs(2803);
    outputs(3821) <= layer4_outputs(1156);
    outputs(3822) <= not(layer4_outputs(3824));
    outputs(3823) <= not((layer4_outputs(3331)) or (layer4_outputs(7500)));
    outputs(3824) <= not((layer4_outputs(2578)) and (layer4_outputs(6488)));
    outputs(3825) <= not(layer4_outputs(3131));
    outputs(3826) <= layer4_outputs(1813);
    outputs(3827) <= (layer4_outputs(6093)) and not (layer4_outputs(5966));
    outputs(3828) <= not(layer4_outputs(1762));
    outputs(3829) <= not((layer4_outputs(6121)) or (layer4_outputs(4228)));
    outputs(3830) <= not(layer4_outputs(2565));
    outputs(3831) <= layer4_outputs(7469);
    outputs(3832) <= not(layer4_outputs(3286));
    outputs(3833) <= not(layer4_outputs(3424));
    outputs(3834) <= layer4_outputs(4662);
    outputs(3835) <= (layer4_outputs(2277)) and not (layer4_outputs(6616));
    outputs(3836) <= layer4_outputs(2023);
    outputs(3837) <= not((layer4_outputs(6679)) or (layer4_outputs(6350)));
    outputs(3838) <= (layer4_outputs(1456)) and not (layer4_outputs(1729));
    outputs(3839) <= layer4_outputs(1527);
    outputs(3840) <= (layer4_outputs(1434)) and not (layer4_outputs(2355));
    outputs(3841) <= not(layer4_outputs(6345));
    outputs(3842) <= (layer4_outputs(5370)) xor (layer4_outputs(2376));
    outputs(3843) <= not(layer4_outputs(6626));
    outputs(3844) <= not(layer4_outputs(7096));
    outputs(3845) <= not(layer4_outputs(4054));
    outputs(3846) <= not(layer4_outputs(4990));
    outputs(3847) <= layer4_outputs(5013);
    outputs(3848) <= not(layer4_outputs(6858));
    outputs(3849) <= not((layer4_outputs(4759)) xor (layer4_outputs(5034)));
    outputs(3850) <= not(layer4_outputs(5192)) or (layer4_outputs(277));
    outputs(3851) <= not(layer4_outputs(3509)) or (layer4_outputs(7080));
    outputs(3852) <= (layer4_outputs(3137)) xor (layer4_outputs(5711));
    outputs(3853) <= layer4_outputs(6197);
    outputs(3854) <= not(layer4_outputs(6840));
    outputs(3855) <= not((layer4_outputs(4472)) xor (layer4_outputs(2993)));
    outputs(3856) <= not((layer4_outputs(5615)) xor (layer4_outputs(3139)));
    outputs(3857) <= not((layer4_outputs(6083)) xor (layer4_outputs(1603)));
    outputs(3858) <= (layer4_outputs(5524)) and not (layer4_outputs(6107));
    outputs(3859) <= not((layer4_outputs(4078)) or (layer4_outputs(4529)));
    outputs(3860) <= not(layer4_outputs(3128));
    outputs(3861) <= (layer4_outputs(1062)) xor (layer4_outputs(329));
    outputs(3862) <= not(layer4_outputs(6175));
    outputs(3863) <= not((layer4_outputs(7445)) and (layer4_outputs(6230)));
    outputs(3864) <= layer4_outputs(6832);
    outputs(3865) <= not(layer4_outputs(2192)) or (layer4_outputs(4618));
    outputs(3866) <= not(layer4_outputs(4887)) or (layer4_outputs(5502));
    outputs(3867) <= not((layer4_outputs(7088)) xor (layer4_outputs(7589)));
    outputs(3868) <= not(layer4_outputs(2136));
    outputs(3869) <= (layer4_outputs(2512)) and not (layer4_outputs(2576));
    outputs(3870) <= not(layer4_outputs(2431));
    outputs(3871) <= layer4_outputs(7144);
    outputs(3872) <= not(layer4_outputs(3995));
    outputs(3873) <= layer4_outputs(4512);
    outputs(3874) <= not((layer4_outputs(6417)) xor (layer4_outputs(4783)));
    outputs(3875) <= (layer4_outputs(5198)) and (layer4_outputs(6480));
    outputs(3876) <= (layer4_outputs(2140)) xor (layer4_outputs(1425));
    outputs(3877) <= (layer4_outputs(5422)) and not (layer4_outputs(30));
    outputs(3878) <= layer4_outputs(1896);
    outputs(3879) <= (layer4_outputs(4959)) and not (layer4_outputs(1547));
    outputs(3880) <= layer4_outputs(6842);
    outputs(3881) <= not(layer4_outputs(246));
    outputs(3882) <= not(layer4_outputs(2614));
    outputs(3883) <= layer4_outputs(6964);
    outputs(3884) <= (layer4_outputs(439)) and not (layer4_outputs(1219));
    outputs(3885) <= not(layer4_outputs(3697));
    outputs(3886) <= not(layer4_outputs(5237)) or (layer4_outputs(6101));
    outputs(3887) <= not(layer4_outputs(7357));
    outputs(3888) <= layer4_outputs(2925);
    outputs(3889) <= not((layer4_outputs(6876)) xor (layer4_outputs(7091)));
    outputs(3890) <= not(layer4_outputs(168));
    outputs(3891) <= (layer4_outputs(3947)) and not (layer4_outputs(5940));
    outputs(3892) <= (layer4_outputs(6497)) and not (layer4_outputs(5288));
    outputs(3893) <= (layer4_outputs(2835)) xor (layer4_outputs(3580));
    outputs(3894) <= layer4_outputs(6306);
    outputs(3895) <= (layer4_outputs(4184)) xor (layer4_outputs(2882));
    outputs(3896) <= layer4_outputs(7486);
    outputs(3897) <= layer4_outputs(5330);
    outputs(3898) <= (layer4_outputs(3612)) xor (layer4_outputs(1121));
    outputs(3899) <= (layer4_outputs(3654)) and not (layer4_outputs(1937));
    outputs(3900) <= not(layer4_outputs(2442));
    outputs(3901) <= layer4_outputs(972);
    outputs(3902) <= (layer4_outputs(7327)) and not (layer4_outputs(869));
    outputs(3903) <= not(layer4_outputs(6227));
    outputs(3904) <= not(layer4_outputs(538));
    outputs(3905) <= layer4_outputs(200);
    outputs(3906) <= not(layer4_outputs(1825));
    outputs(3907) <= (layer4_outputs(5379)) and (layer4_outputs(576));
    outputs(3908) <= (layer4_outputs(6231)) xor (layer4_outputs(5019));
    outputs(3909) <= not((layer4_outputs(7430)) xor (layer4_outputs(3766)));
    outputs(3910) <= (layer4_outputs(3992)) xor (layer4_outputs(5624));
    outputs(3911) <= not(layer4_outputs(5227));
    outputs(3912) <= not(layer4_outputs(7461));
    outputs(3913) <= layer4_outputs(4182);
    outputs(3914) <= not(layer4_outputs(6325));
    outputs(3915) <= layer4_outputs(1769);
    outputs(3916) <= (layer4_outputs(1022)) xor (layer4_outputs(7425));
    outputs(3917) <= layer4_outputs(5263);
    outputs(3918) <= (layer4_outputs(4483)) and not (layer4_outputs(7052));
    outputs(3919) <= not((layer4_outputs(6928)) xor (layer4_outputs(1797)));
    outputs(3920) <= layer4_outputs(2845);
    outputs(3921) <= not((layer4_outputs(3787)) or (layer4_outputs(589)));
    outputs(3922) <= layer4_outputs(2070);
    outputs(3923) <= layer4_outputs(1792);
    outputs(3924) <= (layer4_outputs(6007)) and not (layer4_outputs(2120));
    outputs(3925) <= (layer4_outputs(6145)) xor (layer4_outputs(4342));
    outputs(3926) <= not(layer4_outputs(5402));
    outputs(3927) <= layer4_outputs(3459);
    outputs(3928) <= not(layer4_outputs(5498));
    outputs(3929) <= not(layer4_outputs(6643));
    outputs(3930) <= (layer4_outputs(7467)) xor (layer4_outputs(3815));
    outputs(3931) <= (layer4_outputs(484)) xor (layer4_outputs(3515));
    outputs(3932) <= (layer4_outputs(6137)) and not (layer4_outputs(3443));
    outputs(3933) <= layer4_outputs(2425);
    outputs(3934) <= not((layer4_outputs(2806)) and (layer4_outputs(953)));
    outputs(3935) <= layer4_outputs(5631);
    outputs(3936) <= layer4_outputs(1361);
    outputs(3937) <= not((layer4_outputs(1268)) xor (layer4_outputs(2442)));
    outputs(3938) <= layer4_outputs(4387);
    outputs(3939) <= (layer4_outputs(1151)) xor (layer4_outputs(1924));
    outputs(3940) <= (layer4_outputs(6085)) or (layer4_outputs(4935));
    outputs(3941) <= not((layer4_outputs(6582)) xor (layer4_outputs(3242)));
    outputs(3942) <= not((layer4_outputs(7055)) xor (layer4_outputs(6590)));
    outputs(3943) <= layer4_outputs(6865);
    outputs(3944) <= (layer4_outputs(2048)) xor (layer4_outputs(3618));
    outputs(3945) <= not((layer4_outputs(1992)) and (layer4_outputs(6434)));
    outputs(3946) <= not(layer4_outputs(5610));
    outputs(3947) <= layer4_outputs(2513);
    outputs(3948) <= not((layer4_outputs(4378)) or (layer4_outputs(4075)));
    outputs(3949) <= layer4_outputs(6935);
    outputs(3950) <= layer4_outputs(1113);
    outputs(3951) <= not(layer4_outputs(6841));
    outputs(3952) <= not(layer4_outputs(2424));
    outputs(3953) <= layer4_outputs(1941);
    outputs(3954) <= not(layer4_outputs(5894));
    outputs(3955) <= layer4_outputs(2654);
    outputs(3956) <= not((layer4_outputs(1143)) xor (layer4_outputs(4172)));
    outputs(3957) <= not(layer4_outputs(2215));
    outputs(3958) <= (layer4_outputs(2464)) xor (layer4_outputs(6726));
    outputs(3959) <= not(layer4_outputs(2994));
    outputs(3960) <= (layer4_outputs(521)) and not (layer4_outputs(6214));
    outputs(3961) <= not((layer4_outputs(1560)) xor (layer4_outputs(3892)));
    outputs(3962) <= layer4_outputs(210);
    outputs(3963) <= layer4_outputs(381);
    outputs(3964) <= not((layer4_outputs(4322)) and (layer4_outputs(600)));
    outputs(3965) <= layer4_outputs(1340);
    outputs(3966) <= not(layer4_outputs(3222));
    outputs(3967) <= layer4_outputs(1518);
    outputs(3968) <= layer4_outputs(1915);
    outputs(3969) <= layer4_outputs(1873);
    outputs(3970) <= not(layer4_outputs(7487));
    outputs(3971) <= not((layer4_outputs(2216)) xor (layer4_outputs(1404)));
    outputs(3972) <= not((layer4_outputs(7325)) xor (layer4_outputs(1401)));
    outputs(3973) <= not((layer4_outputs(6990)) xor (layer4_outputs(2842)));
    outputs(3974) <= layer4_outputs(6669);
    outputs(3975) <= not((layer4_outputs(5472)) xor (layer4_outputs(4223)));
    outputs(3976) <= not((layer4_outputs(3678)) xor (layer4_outputs(1618)));
    outputs(3977) <= not(layer4_outputs(2445));
    outputs(3978) <= not(layer4_outputs(4676));
    outputs(3979) <= layer4_outputs(4131);
    outputs(3980) <= layer4_outputs(2457);
    outputs(3981) <= (layer4_outputs(371)) or (layer4_outputs(3017));
    outputs(3982) <= layer4_outputs(836);
    outputs(3983) <= layer4_outputs(5025);
    outputs(3984) <= not((layer4_outputs(739)) xor (layer4_outputs(3668)));
    outputs(3985) <= (layer4_outputs(3891)) and (layer4_outputs(4432));
    outputs(3986) <= (layer4_outputs(6535)) xor (layer4_outputs(5529));
    outputs(3987) <= (layer4_outputs(4951)) xor (layer4_outputs(568));
    outputs(3988) <= not(layer4_outputs(3027));
    outputs(3989) <= (layer4_outputs(121)) xor (layer4_outputs(6140));
    outputs(3990) <= not((layer4_outputs(5500)) xor (layer4_outputs(6081)));
    outputs(3991) <= not(layer4_outputs(6790));
    outputs(3992) <= (layer4_outputs(441)) xor (layer4_outputs(512));
    outputs(3993) <= not(layer4_outputs(3814));
    outputs(3994) <= (layer4_outputs(1503)) xor (layer4_outputs(6168));
    outputs(3995) <= (layer4_outputs(3797)) and (layer4_outputs(5305));
    outputs(3996) <= layer4_outputs(2600);
    outputs(3997) <= layer4_outputs(4746);
    outputs(3998) <= not(layer4_outputs(7585));
    outputs(3999) <= not((layer4_outputs(2033)) or (layer4_outputs(4334)));
    outputs(4000) <= layer4_outputs(6100);
    outputs(4001) <= not(layer4_outputs(3458));
    outputs(4002) <= not((layer4_outputs(1320)) xor (layer4_outputs(2121)));
    outputs(4003) <= not(layer4_outputs(1492));
    outputs(4004) <= not(layer4_outputs(3921));
    outputs(4005) <= not((layer4_outputs(3904)) xor (layer4_outputs(608)));
    outputs(4006) <= layer4_outputs(6085);
    outputs(4007) <= not((layer4_outputs(5365)) and (layer4_outputs(3440)));
    outputs(4008) <= not((layer4_outputs(159)) and (layer4_outputs(795)));
    outputs(4009) <= (layer4_outputs(4196)) xor (layer4_outputs(5032));
    outputs(4010) <= layer4_outputs(5454);
    outputs(4011) <= (layer4_outputs(4213)) xor (layer4_outputs(6897));
    outputs(4012) <= (layer4_outputs(708)) xor (layer4_outputs(5819));
    outputs(4013) <= layer4_outputs(771);
    outputs(4014) <= (layer4_outputs(330)) xor (layer4_outputs(2347));
    outputs(4015) <= not(layer4_outputs(7657));
    outputs(4016) <= layer4_outputs(2881);
    outputs(4017) <= not(layer4_outputs(2439));
    outputs(4018) <= layer4_outputs(4437);
    outputs(4019) <= not(layer4_outputs(7012));
    outputs(4020) <= layer4_outputs(1929);
    outputs(4021) <= (layer4_outputs(6873)) xor (layer4_outputs(1432));
    outputs(4022) <= not(layer4_outputs(4428));
    outputs(4023) <= not((layer4_outputs(3985)) xor (layer4_outputs(2098)));
    outputs(4024) <= layer4_outputs(1844);
    outputs(4025) <= not(layer4_outputs(2698));
    outputs(4026) <= not(layer4_outputs(6380));
    outputs(4027) <= (layer4_outputs(440)) or (layer4_outputs(5705));
    outputs(4028) <= not((layer4_outputs(4819)) xor (layer4_outputs(5220)));
    outputs(4029) <= not(layer4_outputs(5));
    outputs(4030) <= not((layer4_outputs(3817)) xor (layer4_outputs(593)));
    outputs(4031) <= not((layer4_outputs(5646)) xor (layer4_outputs(3749)));
    outputs(4032) <= not((layer4_outputs(4866)) and (layer4_outputs(5035)));
    outputs(4033) <= layer4_outputs(6850);
    outputs(4034) <= not((layer4_outputs(3565)) or (layer4_outputs(3592)));
    outputs(4035) <= (layer4_outputs(4628)) xor (layer4_outputs(6718));
    outputs(4036) <= layer4_outputs(3461);
    outputs(4037) <= not((layer4_outputs(5717)) or (layer4_outputs(2516)));
    outputs(4038) <= not((layer4_outputs(7034)) xor (layer4_outputs(5094)));
    outputs(4039) <= not(layer4_outputs(993));
    outputs(4040) <= layer4_outputs(2580);
    outputs(4041) <= (layer4_outputs(5090)) or (layer4_outputs(4569));
    outputs(4042) <= (layer4_outputs(4804)) xor (layer4_outputs(274));
    outputs(4043) <= not(layer4_outputs(6915));
    outputs(4044) <= (layer4_outputs(2696)) xor (layer4_outputs(5499));
    outputs(4045) <= not((layer4_outputs(5767)) xor (layer4_outputs(6820)));
    outputs(4046) <= not(layer4_outputs(1619));
    outputs(4047) <= not(layer4_outputs(3084)) or (layer4_outputs(7366));
    outputs(4048) <= not(layer4_outputs(7217)) or (layer4_outputs(2572));
    outputs(4049) <= (layer4_outputs(3760)) xor (layer4_outputs(3702));
    outputs(4050) <= layer4_outputs(5001);
    outputs(4051) <= layer4_outputs(6613);
    outputs(4052) <= layer4_outputs(6415);
    outputs(4053) <= not((layer4_outputs(6274)) xor (layer4_outputs(6501)));
    outputs(4054) <= layer4_outputs(6217);
    outputs(4055) <= not(layer4_outputs(3357)) or (layer4_outputs(5749));
    outputs(4056) <= layer4_outputs(1217);
    outputs(4057) <= not(layer4_outputs(401));
    outputs(4058) <= not((layer4_outputs(718)) or (layer4_outputs(7199)));
    outputs(4059) <= not(layer4_outputs(6017)) or (layer4_outputs(717));
    outputs(4060) <= layer4_outputs(380);
    outputs(4061) <= not((layer4_outputs(2669)) xor (layer4_outputs(6689)));
    outputs(4062) <= not(layer4_outputs(3163));
    outputs(4063) <= not(layer4_outputs(2239)) or (layer4_outputs(1057));
    outputs(4064) <= not((layer4_outputs(6291)) xor (layer4_outputs(910)));
    outputs(4065) <= not(layer4_outputs(2989));
    outputs(4066) <= (layer4_outputs(1230)) and not (layer4_outputs(7122));
    outputs(4067) <= layer4_outputs(3873);
    outputs(4068) <= not(layer4_outputs(7603));
    outputs(4069) <= not(layer4_outputs(1308));
    outputs(4070) <= (layer4_outputs(6836)) or (layer4_outputs(5433));
    outputs(4071) <= (layer4_outputs(7492)) and not (layer4_outputs(3393));
    outputs(4072) <= not((layer4_outputs(7664)) xor (layer4_outputs(5930)));
    outputs(4073) <= layer4_outputs(7108);
    outputs(4074) <= not((layer4_outputs(1836)) and (layer4_outputs(6360)));
    outputs(4075) <= (layer4_outputs(4332)) xor (layer4_outputs(5830));
    outputs(4076) <= not(layer4_outputs(126));
    outputs(4077) <= layer4_outputs(1047);
    outputs(4078) <= not(layer4_outputs(5589));
    outputs(4079) <= not((layer4_outputs(3832)) and (layer4_outputs(3157)));
    outputs(4080) <= not(layer4_outputs(527));
    outputs(4081) <= (layer4_outputs(5959)) xor (layer4_outputs(6636));
    outputs(4082) <= layer4_outputs(6616);
    outputs(4083) <= (layer4_outputs(2520)) xor (layer4_outputs(1128));
    outputs(4084) <= not((layer4_outputs(4323)) xor (layer4_outputs(1981)));
    outputs(4085) <= (layer4_outputs(1834)) xor (layer4_outputs(1457));
    outputs(4086) <= (layer4_outputs(3198)) xor (layer4_outputs(3682));
    outputs(4087) <= not(layer4_outputs(4456));
    outputs(4088) <= not((layer4_outputs(2130)) or (layer4_outputs(940)));
    outputs(4089) <= not((layer4_outputs(5560)) xor (layer4_outputs(4013)));
    outputs(4090) <= not(layer4_outputs(5083));
    outputs(4091) <= not(layer4_outputs(7476));
    outputs(4092) <= not((layer4_outputs(6338)) xor (layer4_outputs(3637)));
    outputs(4093) <= (layer4_outputs(6094)) and (layer4_outputs(3279));
    outputs(4094) <= not((layer4_outputs(3727)) xor (layer4_outputs(6869)));
    outputs(4095) <= not((layer4_outputs(5060)) xor (layer4_outputs(2991)));
    outputs(4096) <= layer4_outputs(2221);
    outputs(4097) <= not(layer4_outputs(7030));
    outputs(4098) <= layer4_outputs(7526);
    outputs(4099) <= not(layer4_outputs(5505));
    outputs(4100) <= not(layer4_outputs(4648));
    outputs(4101) <= (layer4_outputs(2022)) xor (layer4_outputs(6383));
    outputs(4102) <= (layer4_outputs(291)) xor (layer4_outputs(4631));
    outputs(4103) <= not((layer4_outputs(6640)) xor (layer4_outputs(68)));
    outputs(4104) <= not(layer4_outputs(7271)) or (layer4_outputs(3071));
    outputs(4105) <= not(layer4_outputs(2665)) or (layer4_outputs(5643));
    outputs(4106) <= layer4_outputs(6562);
    outputs(4107) <= layer4_outputs(2936);
    outputs(4108) <= not((layer4_outputs(757)) xor (layer4_outputs(1878)));
    outputs(4109) <= not(layer4_outputs(4579));
    outputs(4110) <= not(layer4_outputs(2941)) or (layer4_outputs(6225));
    outputs(4111) <= not((layer4_outputs(6263)) xor (layer4_outputs(4609)));
    outputs(4112) <= (layer4_outputs(2607)) xor (layer4_outputs(5148));
    outputs(4113) <= not(layer4_outputs(2158));
    outputs(4114) <= (layer4_outputs(4059)) or (layer4_outputs(3150));
    outputs(4115) <= layer4_outputs(5480);
    outputs(4116) <= not(layer4_outputs(338));
    outputs(4117) <= not(layer4_outputs(37));
    outputs(4118) <= not(layer4_outputs(99));
    outputs(4119) <= not(layer4_outputs(2857));
    outputs(4120) <= layer4_outputs(1007);
    outputs(4121) <= layer4_outputs(838);
    outputs(4122) <= (layer4_outputs(1650)) and not (layer4_outputs(5808));
    outputs(4123) <= not(layer4_outputs(2883));
    outputs(4124) <= not(layer4_outputs(7145));
    outputs(4125) <= layer4_outputs(4406);
    outputs(4126) <= (layer4_outputs(889)) xor (layer4_outputs(4069));
    outputs(4127) <= not((layer4_outputs(3165)) and (layer4_outputs(5232)));
    outputs(4128) <= not(layer4_outputs(1913)) or (layer4_outputs(2591));
    outputs(4129) <= not(layer4_outputs(1069));
    outputs(4130) <= (layer4_outputs(5692)) xor (layer4_outputs(205));
    outputs(4131) <= not((layer4_outputs(3198)) xor (layer4_outputs(5731)));
    outputs(4132) <= layer4_outputs(4585);
    outputs(4133) <= not(layer4_outputs(2962));
    outputs(4134) <= not(layer4_outputs(7338));
    outputs(4135) <= not(layer4_outputs(3886));
    outputs(4136) <= not(layer4_outputs(2833));
    outputs(4137) <= not(layer4_outputs(4443));
    outputs(4138) <= not(layer4_outputs(4393));
    outputs(4139) <= not(layer4_outputs(3854));
    outputs(4140) <= not(layer4_outputs(6568));
    outputs(4141) <= layer4_outputs(1342);
    outputs(4142) <= not(layer4_outputs(587));
    outputs(4143) <= not((layer4_outputs(7286)) xor (layer4_outputs(2158)));
    outputs(4144) <= layer4_outputs(514);
    outputs(4145) <= not(layer4_outputs(5940));
    outputs(4146) <= layer4_outputs(2321);
    outputs(4147) <= layer4_outputs(2241);
    outputs(4148) <= (layer4_outputs(1659)) xor (layer4_outputs(2838));
    outputs(4149) <= not(layer4_outputs(3709));
    outputs(4150) <= layer4_outputs(6239);
    outputs(4151) <= not(layer4_outputs(3509));
    outputs(4152) <= not((layer4_outputs(7482)) xor (layer4_outputs(6159)));
    outputs(4153) <= not(layer4_outputs(7129)) or (layer4_outputs(2865));
    outputs(4154) <= layer4_outputs(3967);
    outputs(4155) <= not(layer4_outputs(94)) or (layer4_outputs(2378));
    outputs(4156) <= (layer4_outputs(4528)) and not (layer4_outputs(4917));
    outputs(4157) <= layer4_outputs(613);
    outputs(4158) <= not((layer4_outputs(117)) xor (layer4_outputs(4919)));
    outputs(4159) <= not(layer4_outputs(1408));
    outputs(4160) <= (layer4_outputs(4156)) xor (layer4_outputs(6045));
    outputs(4161) <= (layer4_outputs(4062)) xor (layer4_outputs(3446));
    outputs(4162) <= layer4_outputs(6770);
    outputs(4163) <= not((layer4_outputs(2495)) xor (layer4_outputs(6591)));
    outputs(4164) <= layer4_outputs(1378);
    outputs(4165) <= layer4_outputs(7350);
    outputs(4166) <= not(layer4_outputs(7342));
    outputs(4167) <= not(layer4_outputs(5284));
    outputs(4168) <= (layer4_outputs(6524)) xor (layer4_outputs(3542));
    outputs(4169) <= (layer4_outputs(428)) xor (layer4_outputs(1594));
    outputs(4170) <= (layer4_outputs(3763)) and (layer4_outputs(309));
    outputs(4171) <= (layer4_outputs(5749)) or (layer4_outputs(4139));
    outputs(4172) <= not((layer4_outputs(3784)) and (layer4_outputs(1240)));
    outputs(4173) <= not(layer4_outputs(2014));
    outputs(4174) <= not(layer4_outputs(3953));
    outputs(4175) <= not(layer4_outputs(7340));
    outputs(4176) <= (layer4_outputs(6207)) and not (layer4_outputs(4617));
    outputs(4177) <= (layer4_outputs(2252)) xor (layer4_outputs(6465));
    outputs(4178) <= not(layer4_outputs(1052));
    outputs(4179) <= not((layer4_outputs(6744)) or (layer4_outputs(911)));
    outputs(4180) <= not(layer4_outputs(3610));
    outputs(4181) <= (layer4_outputs(7377)) and not (layer4_outputs(2166));
    outputs(4182) <= not(layer4_outputs(4909));
    outputs(4183) <= (layer4_outputs(1964)) and not (layer4_outputs(323));
    outputs(4184) <= (layer4_outputs(2817)) xor (layer4_outputs(5713));
    outputs(4185) <= layer4_outputs(7462);
    outputs(4186) <= not((layer4_outputs(7277)) or (layer4_outputs(4774)));
    outputs(4187) <= not((layer4_outputs(7443)) xor (layer4_outputs(2815)));
    outputs(4188) <= layer4_outputs(3506);
    outputs(4189) <= not((layer4_outputs(3913)) xor (layer4_outputs(984)));
    outputs(4190) <= not(layer4_outputs(2144));
    outputs(4191) <= not(layer4_outputs(4719));
    outputs(4192) <= layer4_outputs(3207);
    outputs(4193) <= (layer4_outputs(2264)) or (layer4_outputs(1037));
    outputs(4194) <= not((layer4_outputs(5696)) xor (layer4_outputs(3833)));
    outputs(4195) <= not(layer4_outputs(4847));
    outputs(4196) <= layer4_outputs(6694);
    outputs(4197) <= not((layer4_outputs(1050)) xor (layer4_outputs(4391)));
    outputs(4198) <= layer4_outputs(5776);
    outputs(4199) <= not((layer4_outputs(7246)) or (layer4_outputs(6639)));
    outputs(4200) <= layer4_outputs(266);
    outputs(4201) <= not(layer4_outputs(6483));
    outputs(4202) <= layer4_outputs(7134);
    outputs(4203) <= not(layer4_outputs(1485));
    outputs(4204) <= not(layer4_outputs(1619));
    outputs(4205) <= not(layer4_outputs(4442));
    outputs(4206) <= not(layer4_outputs(2895));
    outputs(4207) <= not(layer4_outputs(146));
    outputs(4208) <= not((layer4_outputs(5748)) xor (layer4_outputs(801)));
    outputs(4209) <= not(layer4_outputs(7541));
    outputs(4210) <= (layer4_outputs(5274)) and not (layer4_outputs(1737));
    outputs(4211) <= layer4_outputs(1032);
    outputs(4212) <= not(layer4_outputs(2441));
    outputs(4213) <= not(layer4_outputs(2040));
    outputs(4214) <= not(layer4_outputs(2439));
    outputs(4215) <= not((layer4_outputs(1060)) xor (layer4_outputs(1013)));
    outputs(4216) <= not(layer4_outputs(1909));
    outputs(4217) <= not(layer4_outputs(2137));
    outputs(4218) <= (layer4_outputs(1654)) xor (layer4_outputs(4360));
    outputs(4219) <= (layer4_outputs(5961)) xor (layer4_outputs(2954));
    outputs(4220) <= not((layer4_outputs(6942)) and (layer4_outputs(3925)));
    outputs(4221) <= (layer4_outputs(4318)) xor (layer4_outputs(6815));
    outputs(4222) <= not(layer4_outputs(2037));
    outputs(4223) <= not(layer4_outputs(3008));
    outputs(4224) <= not(layer4_outputs(6555));
    outputs(4225) <= not(layer4_outputs(7020));
    outputs(4226) <= (layer4_outputs(2691)) xor (layer4_outputs(1906));
    outputs(4227) <= not((layer4_outputs(6516)) xor (layer4_outputs(1330)));
    outputs(4228) <= (layer4_outputs(932)) and not (layer4_outputs(3136));
    outputs(4229) <= not(layer4_outputs(1894));
    outputs(4230) <= layer4_outputs(4643);
    outputs(4231) <= (layer4_outputs(1821)) xor (layer4_outputs(7208));
    outputs(4232) <= (layer4_outputs(7121)) and (layer4_outputs(4068));
    outputs(4233) <= not(layer4_outputs(868));
    outputs(4234) <= not(layer4_outputs(2766));
    outputs(4235) <= not(layer4_outputs(782));
    outputs(4236) <= (layer4_outputs(776)) xor (layer4_outputs(2039));
    outputs(4237) <= (layer4_outputs(1312)) xor (layer4_outputs(6886));
    outputs(4238) <= not(layer4_outputs(6521));
    outputs(4239) <= (layer4_outputs(926)) xor (layer4_outputs(7670));
    outputs(4240) <= layer4_outputs(4548);
    outputs(4241) <= layer4_outputs(1555);
    outputs(4242) <= not(layer4_outputs(3385));
    outputs(4243) <= layer4_outputs(602);
    outputs(4244) <= not(layer4_outputs(3476));
    outputs(4245) <= not(layer4_outputs(2466));
    outputs(4246) <= layer4_outputs(1447);
    outputs(4247) <= not(layer4_outputs(899)) or (layer4_outputs(1540));
    outputs(4248) <= layer4_outputs(2927);
    outputs(4249) <= layer4_outputs(3400);
    outputs(4250) <= (layer4_outputs(5000)) xor (layer4_outputs(4807));
    outputs(4251) <= not((layer4_outputs(6348)) xor (layer4_outputs(2001)));
    outputs(4252) <= layer4_outputs(1384);
    outputs(4253) <= layer4_outputs(3698);
    outputs(4254) <= not((layer4_outputs(6647)) and (layer4_outputs(5284)));
    outputs(4255) <= not(layer4_outputs(1358));
    outputs(4256) <= layer4_outputs(5705);
    outputs(4257) <= not((layer4_outputs(1886)) and (layer4_outputs(7269)));
    outputs(4258) <= layer4_outputs(1521);
    outputs(4259) <= not(layer4_outputs(44));
    outputs(4260) <= not(layer4_outputs(6312));
    outputs(4261) <= layer4_outputs(3459);
    outputs(4262) <= (layer4_outputs(7466)) and not (layer4_outputs(4126));
    outputs(4263) <= not(layer4_outputs(7335));
    outputs(4264) <= not(layer4_outputs(849));
    outputs(4265) <= layer4_outputs(2159);
    outputs(4266) <= (layer4_outputs(4146)) and not (layer4_outputs(3443));
    outputs(4267) <= not(layer4_outputs(2589));
    outputs(4268) <= layer4_outputs(1768);
    outputs(4269) <= (layer4_outputs(6989)) and not (layer4_outputs(2395));
    outputs(4270) <= layer4_outputs(3463);
    outputs(4271) <= not((layer4_outputs(4555)) xor (layer4_outputs(7104)));
    outputs(4272) <= layer4_outputs(6305);
    outputs(4273) <= not(layer4_outputs(1368));
    outputs(4274) <= layer4_outputs(230);
    outputs(4275) <= layer4_outputs(7163);
    outputs(4276) <= layer4_outputs(1339);
    outputs(4277) <= (layer4_outputs(2372)) and (layer4_outputs(6705));
    outputs(4278) <= not(layer4_outputs(7631));
    outputs(4279) <= not(layer4_outputs(6954));
    outputs(4280) <= layer4_outputs(875);
    outputs(4281) <= not(layer4_outputs(81));
    outputs(4282) <= layer4_outputs(1428);
    outputs(4283) <= not(layer4_outputs(742));
    outputs(4284) <= (layer4_outputs(4479)) xor (layer4_outputs(5639));
    outputs(4285) <= not(layer4_outputs(3974));
    outputs(4286) <= not(layer4_outputs(6345));
    outputs(4287) <= layer4_outputs(7529);
    outputs(4288) <= not((layer4_outputs(5513)) xor (layer4_outputs(978)));
    outputs(4289) <= not((layer4_outputs(5857)) xor (layer4_outputs(2380)));
    outputs(4290) <= not((layer4_outputs(5978)) and (layer4_outputs(7019)));
    outputs(4291) <= not(layer4_outputs(2817));
    outputs(4292) <= layer4_outputs(6083);
    outputs(4293) <= not(layer4_outputs(6672));
    outputs(4294) <= not(layer4_outputs(3503));
    outputs(4295) <= (layer4_outputs(386)) xor (layer4_outputs(3753));
    outputs(4296) <= layer4_outputs(5900);
    outputs(4297) <= not((layer4_outputs(1028)) xor (layer4_outputs(268)));
    outputs(4298) <= not((layer4_outputs(5249)) and (layer4_outputs(3031)));
    outputs(4299) <= not((layer4_outputs(2436)) xor (layer4_outputs(2928)));
    outputs(4300) <= layer4_outputs(5092);
    outputs(4301) <= layer4_outputs(469);
    outputs(4302) <= not((layer4_outputs(3421)) or (layer4_outputs(6895)));
    outputs(4303) <= not((layer4_outputs(3416)) and (layer4_outputs(2030)));
    outputs(4304) <= not(layer4_outputs(4414));
    outputs(4305) <= (layer4_outputs(641)) and (layer4_outputs(6881));
    outputs(4306) <= layer4_outputs(1338);
    outputs(4307) <= not(layer4_outputs(2649)) or (layer4_outputs(2419));
    outputs(4308) <= layer4_outputs(2193);
    outputs(4309) <= not(layer4_outputs(6198)) or (layer4_outputs(2150));
    outputs(4310) <= (layer4_outputs(1991)) and not (layer4_outputs(3435));
    outputs(4311) <= layer4_outputs(1397);
    outputs(4312) <= layer4_outputs(3261);
    outputs(4313) <= (layer4_outputs(1769)) xor (layer4_outputs(3848));
    outputs(4314) <= not((layer4_outputs(6768)) xor (layer4_outputs(1390)));
    outputs(4315) <= (layer4_outputs(887)) xor (layer4_outputs(5479));
    outputs(4316) <= not(layer4_outputs(1926)) or (layer4_outputs(7154));
    outputs(4317) <= (layer4_outputs(1536)) or (layer4_outputs(7137));
    outputs(4318) <= not(layer4_outputs(3308));
    outputs(4319) <= not(layer4_outputs(3354));
    outputs(4320) <= layer4_outputs(2646);
    outputs(4321) <= not(layer4_outputs(3168));
    outputs(4322) <= (layer4_outputs(7575)) xor (layer4_outputs(927));
    outputs(4323) <= not((layer4_outputs(4426)) xor (layer4_outputs(3314)));
    outputs(4324) <= not(layer4_outputs(2675));
    outputs(4325) <= layer4_outputs(1598);
    outputs(4326) <= (layer4_outputs(2528)) xor (layer4_outputs(2295));
    outputs(4327) <= not(layer4_outputs(396)) or (layer4_outputs(2861));
    outputs(4328) <= (layer4_outputs(2162)) xor (layer4_outputs(6874));
    outputs(4329) <= not((layer4_outputs(513)) xor (layer4_outputs(7042)));
    outputs(4330) <= not(layer4_outputs(4294));
    outputs(4331) <= (layer4_outputs(355)) xor (layer4_outputs(4599));
    outputs(4332) <= layer4_outputs(6116);
    outputs(4333) <= layer4_outputs(4896);
    outputs(4334) <= layer4_outputs(6472);
    outputs(4335) <= (layer4_outputs(3514)) and (layer4_outputs(6684));
    outputs(4336) <= (layer4_outputs(4523)) xor (layer4_outputs(4381));
    outputs(4337) <= layer4_outputs(6362);
    outputs(4338) <= (layer4_outputs(5979)) xor (layer4_outputs(3153));
    outputs(4339) <= not(layer4_outputs(3662));
    outputs(4340) <= not(layer4_outputs(3903));
    outputs(4341) <= not((layer4_outputs(522)) or (layer4_outputs(506)));
    outputs(4342) <= (layer4_outputs(2247)) and not (layer4_outputs(581));
    outputs(4343) <= (layer4_outputs(7496)) and (layer4_outputs(2950));
    outputs(4344) <= not(layer4_outputs(6208));
    outputs(4345) <= layer4_outputs(7094);
    outputs(4346) <= not((layer4_outputs(3658)) xor (layer4_outputs(1936)));
    outputs(4347) <= not(layer4_outputs(970));
    outputs(4348) <= not(layer4_outputs(6971));
    outputs(4349) <= layer4_outputs(7105);
    outputs(4350) <= not(layer4_outputs(2468));
    outputs(4351) <= layer4_outputs(2940);
    outputs(4352) <= (layer4_outputs(6761)) or (layer4_outputs(6066));
    outputs(4353) <= layer4_outputs(6510);
    outputs(4354) <= layer4_outputs(251);
    outputs(4355) <= (layer4_outputs(480)) xor (layer4_outputs(3529));
    outputs(4356) <= not((layer4_outputs(4289)) and (layer4_outputs(729)));
    outputs(4357) <= (layer4_outputs(3013)) xor (layer4_outputs(1744));
    outputs(4358) <= not(layer4_outputs(1271));
    outputs(4359) <= not(layer4_outputs(4770)) or (layer4_outputs(4625));
    outputs(4360) <= not(layer4_outputs(1465));
    outputs(4361) <= not(layer4_outputs(3295));
    outputs(4362) <= layer4_outputs(7500);
    outputs(4363) <= not((layer4_outputs(176)) or (layer4_outputs(6317)));
    outputs(4364) <= layer4_outputs(5741);
    outputs(4365) <= not(layer4_outputs(1583));
    outputs(4366) <= layer4_outputs(5535);
    outputs(4367) <= (layer4_outputs(2610)) xor (layer4_outputs(3908));
    outputs(4368) <= not(layer4_outputs(6961));
    outputs(4369) <= layer4_outputs(7041);
    outputs(4370) <= layer4_outputs(5001);
    outputs(4371) <= layer4_outputs(6172);
    outputs(4372) <= not(layer4_outputs(5340));
    outputs(4373) <= layer4_outputs(2786);
    outputs(4374) <= layer4_outputs(493);
    outputs(4375) <= layer4_outputs(4296);
    outputs(4376) <= (layer4_outputs(6764)) xor (layer4_outputs(295));
    outputs(4377) <= layer4_outputs(7381);
    outputs(4378) <= not((layer4_outputs(6433)) xor (layer4_outputs(3164)));
    outputs(4379) <= not(layer4_outputs(6009));
    outputs(4380) <= (layer4_outputs(7100)) and not (layer4_outputs(1983));
    outputs(4381) <= layer4_outputs(2946);
    outputs(4382) <= not((layer4_outputs(4073)) xor (layer4_outputs(983)));
    outputs(4383) <= layer4_outputs(3162);
    outputs(4384) <= layer4_outputs(6500);
    outputs(4385) <= not((layer4_outputs(5567)) or (layer4_outputs(7066)));
    outputs(4386) <= not((layer4_outputs(4395)) xor (layer4_outputs(2333)));
    outputs(4387) <= (layer4_outputs(5083)) xor (layer4_outputs(52));
    outputs(4388) <= not(layer4_outputs(1947));
    outputs(4389) <= not((layer4_outputs(2509)) xor (layer4_outputs(1117)));
    outputs(4390) <= not((layer4_outputs(5504)) xor (layer4_outputs(1136)));
    outputs(4391) <= layer4_outputs(968);
    outputs(4392) <= layer4_outputs(1957);
    outputs(4393) <= layer4_outputs(3189);
    outputs(4394) <= layer4_outputs(612);
    outputs(4395) <= (layer4_outputs(1236)) and not (layer4_outputs(4431));
    outputs(4396) <= not((layer4_outputs(4738)) xor (layer4_outputs(6912)));
    outputs(4397) <= (layer4_outputs(6118)) and not (layer4_outputs(4155));
    outputs(4398) <= not(layer4_outputs(7430));
    outputs(4399) <= not(layer4_outputs(6798));
    outputs(4400) <= layer4_outputs(2363);
    outputs(4401) <= not(layer4_outputs(6144));
    outputs(4402) <= (layer4_outputs(1386)) xor (layer4_outputs(4476));
    outputs(4403) <= not(layer4_outputs(225));
    outputs(4404) <= not(layer4_outputs(2042));
    outputs(4405) <= layer4_outputs(5152);
    outputs(4406) <= (layer4_outputs(1407)) xor (layer4_outputs(7196));
    outputs(4407) <= (layer4_outputs(3746)) and (layer4_outputs(7601));
    outputs(4408) <= not(layer4_outputs(4640));
    outputs(4409) <= not(layer4_outputs(1283));
    outputs(4410) <= layer4_outputs(5213);
    outputs(4411) <= layer4_outputs(5986);
    outputs(4412) <= layer4_outputs(5516);
    outputs(4413) <= not((layer4_outputs(1054)) xor (layer4_outputs(4836)));
    outputs(4414) <= (layer4_outputs(6099)) or (layer4_outputs(6691));
    outputs(4415) <= layer4_outputs(6260);
    outputs(4416) <= not(layer4_outputs(1349)) or (layer4_outputs(283));
    outputs(4417) <= not(layer4_outputs(7464));
    outputs(4418) <= layer4_outputs(7560);
    outputs(4419) <= not(layer4_outputs(4705));
    outputs(4420) <= not(layer4_outputs(4075));
    outputs(4421) <= not(layer4_outputs(462));
    outputs(4422) <= not(layer4_outputs(1484));
    outputs(4423) <= not((layer4_outputs(4256)) xor (layer4_outputs(2944)));
    outputs(4424) <= not((layer4_outputs(2011)) xor (layer4_outputs(1954)));
    outputs(4425) <= not((layer4_outputs(6597)) xor (layer4_outputs(5259)));
    outputs(4426) <= layer4_outputs(1172);
    outputs(4427) <= not((layer4_outputs(7248)) xor (layer4_outputs(4504)));
    outputs(4428) <= not((layer4_outputs(5178)) xor (layer4_outputs(1569)));
    outputs(4429) <= (layer4_outputs(5701)) xor (layer4_outputs(6175));
    outputs(4430) <= layer4_outputs(1727);
    outputs(4431) <= layer4_outputs(1817);
    outputs(4432) <= not(layer4_outputs(4619));
    outputs(4433) <= (layer4_outputs(1501)) xor (layer4_outputs(4573));
    outputs(4434) <= not(layer4_outputs(5726));
    outputs(4435) <= layer4_outputs(4297);
    outputs(4436) <= (layer4_outputs(2363)) xor (layer4_outputs(5050));
    outputs(4437) <= not(layer4_outputs(6505));
    outputs(4438) <= not(layer4_outputs(636)) or (layer4_outputs(2028));
    outputs(4439) <= layer4_outputs(7651);
    outputs(4440) <= layer4_outputs(3555);
    outputs(4441) <= not((layer4_outputs(6733)) xor (layer4_outputs(2066)));
    outputs(4442) <= not((layer4_outputs(4916)) xor (layer4_outputs(5660)));
    outputs(4443) <= (layer4_outputs(2396)) xor (layer4_outputs(1606));
    outputs(4444) <= not(layer4_outputs(7528));
    outputs(4445) <= not(layer4_outputs(2117));
    outputs(4446) <= (layer4_outputs(1310)) xor (layer4_outputs(3617));
    outputs(4447) <= layer4_outputs(2327);
    outputs(4448) <= layer4_outputs(2573);
    outputs(4449) <= not(layer4_outputs(357));
    outputs(4450) <= not(layer4_outputs(5254));
    outputs(4451) <= (layer4_outputs(476)) and (layer4_outputs(5942));
    outputs(4452) <= (layer4_outputs(771)) xor (layer4_outputs(2101));
    outputs(4453) <= (layer4_outputs(7113)) and not (layer4_outputs(1696));
    outputs(4454) <= (layer4_outputs(6714)) or (layer4_outputs(2375));
    outputs(4455) <= layer4_outputs(442);
    outputs(4456) <= not((layer4_outputs(420)) xor (layer4_outputs(7059)));
    outputs(4457) <= (layer4_outputs(4303)) and not (layer4_outputs(2904));
    outputs(4458) <= not(layer4_outputs(1788));
    outputs(4459) <= layer4_outputs(4660);
    outputs(4460) <= layer4_outputs(788);
    outputs(4461) <= layer4_outputs(6746);
    outputs(4462) <= (layer4_outputs(3860)) and not (layer4_outputs(3435));
    outputs(4463) <= layer4_outputs(62);
    outputs(4464) <= (layer4_outputs(5971)) xor (layer4_outputs(4439));
    outputs(4465) <= layer4_outputs(2880);
    outputs(4466) <= layer4_outputs(796);
    outputs(4467) <= layer4_outputs(3959);
    outputs(4468) <= not((layer4_outputs(4094)) xor (layer4_outputs(6061)));
    outputs(4469) <= not(layer4_outputs(4683));
    outputs(4470) <= layer4_outputs(5185);
    outputs(4471) <= not(layer4_outputs(6486));
    outputs(4472) <= not((layer4_outputs(7419)) xor (layer4_outputs(1364)));
    outputs(4473) <= not(layer4_outputs(2929));
    outputs(4474) <= (layer4_outputs(3880)) or (layer4_outputs(381));
    outputs(4475) <= not(layer4_outputs(1919));
    outputs(4476) <= not(layer4_outputs(600));
    outputs(4477) <= not(layer4_outputs(1357));
    outputs(4478) <= layer4_outputs(5544);
    outputs(4479) <= not(layer4_outputs(5564));
    outputs(4480) <= not((layer4_outputs(4096)) or (layer4_outputs(2522)));
    outputs(4481) <= layer4_outputs(7228);
    outputs(4482) <= layer4_outputs(279);
    outputs(4483) <= layer4_outputs(4865);
    outputs(4484) <= not(layer4_outputs(4673)) or (layer4_outputs(3860));
    outputs(4485) <= not(layer4_outputs(3581));
    outputs(4486) <= layer4_outputs(3904);
    outputs(4487) <= (layer4_outputs(964)) xor (layer4_outputs(1246));
    outputs(4488) <= (layer4_outputs(7346)) xor (layer4_outputs(1953));
    outputs(4489) <= layer4_outputs(3482);
    outputs(4490) <= (layer4_outputs(1525)) xor (layer4_outputs(6867));
    outputs(4491) <= layer4_outputs(1340);
    outputs(4492) <= not(layer4_outputs(6781));
    outputs(4493) <= not(layer4_outputs(4782));
    outputs(4494) <= layer4_outputs(5608);
    outputs(4495) <= not((layer4_outputs(524)) xor (layer4_outputs(1960)));
    outputs(4496) <= not(layer4_outputs(4686));
    outputs(4497) <= layer4_outputs(6713);
    outputs(4498) <= layer4_outputs(4215);
    outputs(4499) <= (layer4_outputs(7251)) or (layer4_outputs(3386));
    outputs(4500) <= layer4_outputs(6412);
    outputs(4501) <= not((layer4_outputs(4721)) xor (layer4_outputs(5019)));
    outputs(4502) <= not(layer4_outputs(6348));
    outputs(4503) <= not(layer4_outputs(2267));
    outputs(4504) <= layer4_outputs(5330);
    outputs(4505) <= not(layer4_outputs(482));
    outputs(4506) <= (layer4_outputs(6929)) and not (layer4_outputs(6234));
    outputs(4507) <= not(layer4_outputs(6917)) or (layer4_outputs(3871));
    outputs(4508) <= layer4_outputs(2623);
    outputs(4509) <= not(layer4_outputs(6447));
    outputs(4510) <= not((layer4_outputs(2546)) xor (layer4_outputs(3172)));
    outputs(4511) <= not((layer4_outputs(3996)) and (layer4_outputs(3362)));
    outputs(4512) <= layer4_outputs(2318);
    outputs(4513) <= not(layer4_outputs(2506));
    outputs(4514) <= not(layer4_outputs(3414));
    outputs(4515) <= (layer4_outputs(5199)) and (layer4_outputs(5263));
    outputs(4516) <= not(layer4_outputs(5668));
    outputs(4517) <= not(layer4_outputs(4183));
    outputs(4518) <= not(layer4_outputs(2195));
    outputs(4519) <= layer4_outputs(3291);
    outputs(4520) <= layer4_outputs(3942);
    outputs(4521) <= not((layer4_outputs(7653)) xor (layer4_outputs(3669)));
    outputs(4522) <= layer4_outputs(5418);
    outputs(4523) <= layer4_outputs(5979);
    outputs(4524) <= layer4_outputs(6178);
    outputs(4525) <= (layer4_outputs(5690)) and not (layer4_outputs(5902));
    outputs(4526) <= not(layer4_outputs(2834));
    outputs(4527) <= (layer4_outputs(4674)) xor (layer4_outputs(1263));
    outputs(4528) <= not(layer4_outputs(3517));
    outputs(4529) <= not(layer4_outputs(6218));
    outputs(4530) <= not(layer4_outputs(864));
    outputs(4531) <= not(layer4_outputs(7133));
    outputs(4532) <= not(layer4_outputs(1524));
    outputs(4533) <= (layer4_outputs(3006)) and (layer4_outputs(6125));
    outputs(4534) <= not((layer4_outputs(2202)) xor (layer4_outputs(1596)));
    outputs(4535) <= not(layer4_outputs(4072));
    outputs(4536) <= layer4_outputs(3425);
    outputs(4537) <= not((layer4_outputs(4083)) and (layer4_outputs(6127)));
    outputs(4538) <= not(layer4_outputs(5832));
    outputs(4539) <= not(layer4_outputs(2448));
    outputs(4540) <= not(layer4_outputs(864));
    outputs(4541) <= not((layer4_outputs(648)) xor (layer4_outputs(4371)));
    outputs(4542) <= (layer4_outputs(4470)) xor (layer4_outputs(2657));
    outputs(4543) <= not(layer4_outputs(5845));
    outputs(4544) <= layer4_outputs(3619);
    outputs(4545) <= layer4_outputs(4198);
    outputs(4546) <= not(layer4_outputs(3024));
    outputs(4547) <= layer4_outputs(5884);
    outputs(4548) <= not(layer4_outputs(3170));
    outputs(4549) <= layer4_outputs(4842);
    outputs(4550) <= layer4_outputs(5898);
    outputs(4551) <= not(layer4_outputs(648)) or (layer4_outputs(1203));
    outputs(4552) <= not(layer4_outputs(6531));
    outputs(4553) <= not(layer4_outputs(1583));
    outputs(4554) <= layer4_outputs(3345);
    outputs(4555) <= (layer4_outputs(6042)) xor (layer4_outputs(7240));
    outputs(4556) <= not((layer4_outputs(7583)) xor (layer4_outputs(6752)));
    outputs(4557) <= not((layer4_outputs(4614)) and (layer4_outputs(4466)));
    outputs(4558) <= (layer4_outputs(110)) xor (layer4_outputs(3078));
    outputs(4559) <= not((layer4_outputs(6133)) xor (layer4_outputs(6026)));
    outputs(4560) <= (layer4_outputs(437)) xor (layer4_outputs(4589));
    outputs(4561) <= not((layer4_outputs(7252)) xor (layer4_outputs(6760)));
    outputs(4562) <= not(layer4_outputs(1181));
    outputs(4563) <= not(layer4_outputs(7360));
    outputs(4564) <= layer4_outputs(7359);
    outputs(4565) <= not(layer4_outputs(6184));
    outputs(4566) <= not(layer4_outputs(3041));
    outputs(4567) <= (layer4_outputs(126)) xor (layer4_outputs(1823));
    outputs(4568) <= not(layer4_outputs(7305));
    outputs(4569) <= not(layer4_outputs(7191));
    outputs(4570) <= (layer4_outputs(1411)) and not (layer4_outputs(1173));
    outputs(4571) <= (layer4_outputs(6844)) xor (layer4_outputs(4096));
    outputs(4572) <= not(layer4_outputs(3403));
    outputs(4573) <= not((layer4_outputs(2301)) xor (layer4_outputs(5798)));
    outputs(4574) <= not((layer4_outputs(1973)) or (layer4_outputs(2208)));
    outputs(4575) <= not((layer4_outputs(4632)) xor (layer4_outputs(4133)));
    outputs(4576) <= not((layer4_outputs(2416)) xor (layer4_outputs(1835)));
    outputs(4577) <= not((layer4_outputs(5674)) or (layer4_outputs(4678)));
    outputs(4578) <= not(layer4_outputs(7206)) or (layer4_outputs(3732));
    outputs(4579) <= not(layer4_outputs(3571));
    outputs(4580) <= not((layer4_outputs(7617)) xor (layer4_outputs(6478)));
    outputs(4581) <= layer4_outputs(5066);
    outputs(4582) <= (layer4_outputs(4796)) xor (layer4_outputs(5518));
    outputs(4583) <= layer4_outputs(2296);
    outputs(4584) <= (layer4_outputs(2240)) and not (layer4_outputs(423));
    outputs(4585) <= not(layer4_outputs(3852)) or (layer4_outputs(3018));
    outputs(4586) <= not(layer4_outputs(2645));
    outputs(4587) <= not((layer4_outputs(3116)) xor (layer4_outputs(4440)));
    outputs(4588) <= layer4_outputs(1520);
    outputs(4589) <= not(layer4_outputs(7670));
    outputs(4590) <= not(layer4_outputs(3768)) or (layer4_outputs(5151));
    outputs(4591) <= not(layer4_outputs(2411));
    outputs(4592) <= (layer4_outputs(4044)) xor (layer4_outputs(2373));
    outputs(4593) <= (layer4_outputs(1302)) and not (layer4_outputs(1071));
    outputs(4594) <= not((layer4_outputs(492)) or (layer4_outputs(5699)));
    outputs(4595) <= not((layer4_outputs(404)) xor (layer4_outputs(7125)));
    outputs(4596) <= not(layer4_outputs(3648)) or (layer4_outputs(5113));
    outputs(4597) <= not(layer4_outputs(3030));
    outputs(4598) <= not((layer4_outputs(2022)) or (layer4_outputs(1978)));
    outputs(4599) <= layer4_outputs(2281);
    outputs(4600) <= (layer4_outputs(7464)) xor (layer4_outputs(5907));
    outputs(4601) <= (layer4_outputs(2524)) xor (layer4_outputs(1114));
    outputs(4602) <= not(layer4_outputs(4630)) or (layer4_outputs(6823));
    outputs(4603) <= layer4_outputs(1938);
    outputs(4604) <= (layer4_outputs(4772)) xor (layer4_outputs(4179));
    outputs(4605) <= not(layer4_outputs(7455)) or (layer4_outputs(6089));
    outputs(4606) <= layer4_outputs(7121);
    outputs(4607) <= not(layer4_outputs(3697));
    outputs(4608) <= layer4_outputs(7323);
    outputs(4609) <= layer4_outputs(5947);
    outputs(4610) <= not(layer4_outputs(1265));
    outputs(4611) <= not(layer4_outputs(2683));
    outputs(4612) <= not(layer4_outputs(3568));
    outputs(4613) <= not(layer4_outputs(4314));
    outputs(4614) <= not((layer4_outputs(3014)) or (layer4_outputs(2504)));
    outputs(4615) <= not((layer4_outputs(1057)) or (layer4_outputs(1643)));
    outputs(4616) <= layer4_outputs(4036);
    outputs(4617) <= not(layer4_outputs(7257));
    outputs(4618) <= layer4_outputs(4064);
    outputs(4619) <= (layer4_outputs(3009)) and not (layer4_outputs(4125));
    outputs(4620) <= not((layer4_outputs(4143)) and (layer4_outputs(5927)));
    outputs(4621) <= not(layer4_outputs(5432));
    outputs(4622) <= (layer4_outputs(6072)) and not (layer4_outputs(5015));
    outputs(4623) <= not((layer4_outputs(5617)) xor (layer4_outputs(5093)));
    outputs(4624) <= not(layer4_outputs(869));
    outputs(4625) <= not(layer4_outputs(3252));
    outputs(4626) <= layer4_outputs(6709);
    outputs(4627) <= (layer4_outputs(6696)) xor (layer4_outputs(3800));
    outputs(4628) <= not((layer4_outputs(2519)) xor (layer4_outputs(1686)));
    outputs(4629) <= not(layer4_outputs(5288));
    outputs(4630) <= (layer4_outputs(4641)) and not (layer4_outputs(4070));
    outputs(4631) <= not((layer4_outputs(1295)) xor (layer4_outputs(7095)));
    outputs(4632) <= not(layer4_outputs(6791)) or (layer4_outputs(6317));
    outputs(4633) <= layer4_outputs(6742);
    outputs(4634) <= not(layer4_outputs(4635));
    outputs(4635) <= layer4_outputs(4497);
    outputs(4636) <= not((layer4_outputs(6653)) or (layer4_outputs(1180)));
    outputs(4637) <= not(layer4_outputs(3079));
    outputs(4638) <= not(layer4_outputs(2019));
    outputs(4639) <= not(layer4_outputs(2529));
    outputs(4640) <= layer4_outputs(7488);
    outputs(4641) <= not(layer4_outputs(1731));
    outputs(4642) <= (layer4_outputs(4518)) xor (layer4_outputs(4388));
    outputs(4643) <= not(layer4_outputs(7543));
    outputs(4644) <= layer4_outputs(5455);
    outputs(4645) <= layer4_outputs(5776);
    outputs(4646) <= layer4_outputs(5876);
    outputs(4647) <= layer4_outputs(6221);
    outputs(4648) <= layer4_outputs(2807);
    outputs(4649) <= (layer4_outputs(4100)) and not (layer4_outputs(7341));
    outputs(4650) <= not((layer4_outputs(6703)) or (layer4_outputs(6202)));
    outputs(4651) <= layer4_outputs(1344);
    outputs(4652) <= (layer4_outputs(4745)) and not (layer4_outputs(4918));
    outputs(4653) <= not((layer4_outputs(3103)) and (layer4_outputs(3642)));
    outputs(4654) <= layer4_outputs(498);
    outputs(4655) <= (layer4_outputs(739)) and (layer4_outputs(1294));
    outputs(4656) <= layer4_outputs(6943);
    outputs(4657) <= not(layer4_outputs(1597));
    outputs(4658) <= not(layer4_outputs(1989));
    outputs(4659) <= not((layer4_outputs(6852)) xor (layer4_outputs(4971)));
    outputs(4660) <= layer4_outputs(3778);
    outputs(4661) <= not(layer4_outputs(50));
    outputs(4662) <= not((layer4_outputs(2120)) or (layer4_outputs(4164)));
    outputs(4663) <= not(layer4_outputs(97)) or (layer4_outputs(1446));
    outputs(4664) <= layer4_outputs(6335);
    outputs(4665) <= (layer4_outputs(2841)) and not (layer4_outputs(4880));
    outputs(4666) <= layer4_outputs(4031);
    outputs(4667) <= not((layer4_outputs(242)) or (layer4_outputs(6549)));
    outputs(4668) <= not((layer4_outputs(7172)) xor (layer4_outputs(4402)));
    outputs(4669) <= not(layer4_outputs(4035));
    outputs(4670) <= not(layer4_outputs(7638));
    outputs(4671) <= (layer4_outputs(2298)) xor (layer4_outputs(2402));
    outputs(4672) <= layer4_outputs(3209);
    outputs(4673) <= not((layer4_outputs(1849)) or (layer4_outputs(6144)));
    outputs(4674) <= (layer4_outputs(4246)) xor (layer4_outputs(349));
    outputs(4675) <= not((layer4_outputs(507)) and (layer4_outputs(341)));
    outputs(4676) <= not(layer4_outputs(4733));
    outputs(4677) <= not(layer4_outputs(1980)) or (layer4_outputs(3437));
    outputs(4678) <= not(layer4_outputs(3186));
    outputs(4679) <= layer4_outputs(2362);
    outputs(4680) <= (layer4_outputs(3896)) or (layer4_outputs(5902));
    outputs(4681) <= layer4_outputs(1258);
    outputs(4682) <= layer4_outputs(4176);
    outputs(4683) <= not(layer4_outputs(3935));
    outputs(4684) <= (layer4_outputs(2059)) and not (layer4_outputs(3794));
    outputs(4685) <= layer4_outputs(2859);
    outputs(4686) <= layer4_outputs(5858);
    outputs(4687) <= not((layer4_outputs(4000)) or (layer4_outputs(4367)));
    outputs(4688) <= (layer4_outputs(6484)) and not (layer4_outputs(6370));
    outputs(4689) <= layer4_outputs(5231);
    outputs(4690) <= (layer4_outputs(5677)) xor (layer4_outputs(5774));
    outputs(4691) <= not(layer4_outputs(7016));
    outputs(4692) <= layer4_outputs(6371);
    outputs(4693) <= (layer4_outputs(5671)) and (layer4_outputs(0));
    outputs(4694) <= layer4_outputs(4532);
    outputs(4695) <= layer4_outputs(1130);
    outputs(4696) <= not(layer4_outputs(4736));
    outputs(4697) <= layer4_outputs(5781);
    outputs(4698) <= (layer4_outputs(7033)) and (layer4_outputs(650));
    outputs(4699) <= (layer4_outputs(726)) and not (layer4_outputs(1287));
    outputs(4700) <= not(layer4_outputs(6519));
    outputs(4701) <= not(layer4_outputs(2161));
    outputs(4702) <= not(layer4_outputs(6845));
    outputs(4703) <= layer4_outputs(3025);
    outputs(4704) <= layer4_outputs(1761);
    outputs(4705) <= not(layer4_outputs(3677));
    outputs(4706) <= layer4_outputs(265);
    outputs(4707) <= layer4_outputs(7);
    outputs(4708) <= layer4_outputs(1556);
    outputs(4709) <= layer4_outputs(4371);
    outputs(4710) <= layer4_outputs(1578);
    outputs(4711) <= layer4_outputs(5722);
    outputs(4712) <= not((layer4_outputs(6229)) and (layer4_outputs(4404)));
    outputs(4713) <= not((layer4_outputs(1595)) xor (layer4_outputs(1665)));
    outputs(4714) <= (layer4_outputs(4086)) and not (layer4_outputs(3251));
    outputs(4715) <= not(layer4_outputs(1063)) or (layer4_outputs(2871));
    outputs(4716) <= layer4_outputs(3243);
    outputs(4717) <= not((layer4_outputs(5258)) and (layer4_outputs(5794)));
    outputs(4718) <= layer4_outputs(5286);
    outputs(4719) <= not((layer4_outputs(4931)) and (layer4_outputs(1086)));
    outputs(4720) <= layer4_outputs(4537);
    outputs(4721) <= not(layer4_outputs(2799));
    outputs(4722) <= (layer4_outputs(5375)) and not (layer4_outputs(5057));
    outputs(4723) <= layer4_outputs(6756);
    outputs(4724) <= not(layer4_outputs(1733));
    outputs(4725) <= layer4_outputs(5518);
    outputs(4726) <= not(layer4_outputs(6767));
    outputs(4727) <= not((layer4_outputs(5229)) or (layer4_outputs(4728)));
    outputs(4728) <= not(layer4_outputs(1362));
    outputs(4729) <= not(layer4_outputs(5301));
    outputs(4730) <= not(layer4_outputs(1805));
    outputs(4731) <= (layer4_outputs(1310)) and not (layer4_outputs(2282));
    outputs(4732) <= not(layer4_outputs(6257));
    outputs(4733) <= layer4_outputs(414);
    outputs(4734) <= layer4_outputs(5316);
    outputs(4735) <= (layer4_outputs(4744)) and (layer4_outputs(2909));
    outputs(4736) <= layer4_outputs(2026);
    outputs(4737) <= not((layer4_outputs(6547)) xor (layer4_outputs(6406)));
    outputs(4738) <= layer4_outputs(6674);
    outputs(4739) <= not(layer4_outputs(6922));
    outputs(4740) <= not(layer4_outputs(3847));
    outputs(4741) <= (layer4_outputs(5493)) and (layer4_outputs(1871));
    outputs(4742) <= not(layer4_outputs(7645));
    outputs(4743) <= (layer4_outputs(999)) and not (layer4_outputs(7490));
    outputs(4744) <= (layer4_outputs(4393)) and not (layer4_outputs(197));
    outputs(4745) <= not(layer4_outputs(116));
    outputs(4746) <= not(layer4_outputs(3883));
    outputs(4747) <= (layer4_outputs(4724)) and (layer4_outputs(6199));
    outputs(4748) <= not(layer4_outputs(1689));
    outputs(4749) <= not(layer4_outputs(5367));
    outputs(4750) <= not(layer4_outputs(1035));
    outputs(4751) <= not(layer4_outputs(1088)) or (layer4_outputs(6452));
    outputs(4752) <= not(layer4_outputs(5463));
    outputs(4753) <= (layer4_outputs(147)) and not (layer4_outputs(2674));
    outputs(4754) <= not((layer4_outputs(3769)) xor (layer4_outputs(3974)));
    outputs(4755) <= layer4_outputs(5602);
    outputs(4756) <= layer4_outputs(3549);
    outputs(4757) <= not(layer4_outputs(6952));
    outputs(4758) <= (layer4_outputs(3)) and not (layer4_outputs(1420));
    outputs(4759) <= (layer4_outputs(1565)) xor (layer4_outputs(7004));
    outputs(4760) <= (layer4_outputs(3738)) xor (layer4_outputs(4685));
    outputs(4761) <= not(layer4_outputs(5815));
    outputs(4762) <= layer4_outputs(796);
    outputs(4763) <= not(layer4_outputs(334));
    outputs(4764) <= not(layer4_outputs(623));
    outputs(4765) <= not(layer4_outputs(6879));
    outputs(4766) <= layer4_outputs(4200);
    outputs(4767) <= layer4_outputs(1680);
    outputs(4768) <= layer4_outputs(3315);
    outputs(4769) <= layer4_outputs(3971);
    outputs(4770) <= not(layer4_outputs(2782));
    outputs(4771) <= (layer4_outputs(3779)) and not (layer4_outputs(4878));
    outputs(4772) <= (layer4_outputs(3214)) and (layer4_outputs(7085));
    outputs(4773) <= (layer4_outputs(71)) and (layer4_outputs(6853));
    outputs(4774) <= not(layer4_outputs(3408));
    outputs(4775) <= not(layer4_outputs(1862));
    outputs(4776) <= not(layer4_outputs(3655));
    outputs(4777) <= (layer4_outputs(272)) and (layer4_outputs(6909));
    outputs(4778) <= not(layer4_outputs(1611));
    outputs(4779) <= (layer4_outputs(1211)) xor (layer4_outputs(4502));
    outputs(4780) <= layer4_outputs(139);
    outputs(4781) <= not(layer4_outputs(5228));
    outputs(4782) <= not(layer4_outputs(3414));
    outputs(4783) <= layer4_outputs(3100);
    outputs(4784) <= (layer4_outputs(5114)) and (layer4_outputs(4896));
    outputs(4785) <= (layer4_outputs(5596)) xor (layer4_outputs(3742));
    outputs(4786) <= layer4_outputs(5700);
    outputs(4787) <= not(layer4_outputs(6019));
    outputs(4788) <= not(layer4_outputs(3096)) or (layer4_outputs(717));
    outputs(4789) <= layer4_outputs(3982);
    outputs(4790) <= (layer4_outputs(6810)) and not (layer4_outputs(3801));
    outputs(4791) <= not(layer4_outputs(987));
    outputs(4792) <= layer4_outputs(2080);
    outputs(4793) <= layer4_outputs(803);
    outputs(4794) <= layer4_outputs(6440);
    outputs(4795) <= not(layer4_outputs(7220)) or (layer4_outputs(192));
    outputs(4796) <= layer4_outputs(1381);
    outputs(4797) <= not(layer4_outputs(2547));
    outputs(4798) <= not(layer4_outputs(4154));
    outputs(4799) <= not((layer4_outputs(4575)) xor (layer4_outputs(6486)));
    outputs(4800) <= not(layer4_outputs(2591));
    outputs(4801) <= not((layer4_outputs(5477)) and (layer4_outputs(6549)));
    outputs(4802) <= (layer4_outputs(1603)) and not (layer4_outputs(4149));
    outputs(4803) <= layer4_outputs(4419);
    outputs(4804) <= not((layer4_outputs(4388)) xor (layer4_outputs(2332)));
    outputs(4805) <= layer4_outputs(473);
    outputs(4806) <= not(layer4_outputs(6483));
    outputs(4807) <= layer4_outputs(6988);
    outputs(4808) <= (layer4_outputs(6802)) xor (layer4_outputs(5139));
    outputs(4809) <= layer4_outputs(2346);
    outputs(4810) <= layer4_outputs(2800);
    outputs(4811) <= not(layer4_outputs(4710));
    outputs(4812) <= (layer4_outputs(1591)) xor (layer4_outputs(1388));
    outputs(4813) <= layer4_outputs(2220);
    outputs(4814) <= (layer4_outputs(3339)) and (layer4_outputs(1717));
    outputs(4815) <= layer4_outputs(7557);
    outputs(4816) <= (layer4_outputs(286)) xor (layer4_outputs(4348));
    outputs(4817) <= (layer4_outputs(4976)) and not (layer4_outputs(2951));
    outputs(4818) <= layer4_outputs(3882);
    outputs(4819) <= layer4_outputs(4700);
    outputs(4820) <= not(layer4_outputs(3501));
    outputs(4821) <= not(layer4_outputs(15));
    outputs(4822) <= not(layer4_outputs(278));
    outputs(4823) <= (layer4_outputs(7308)) and not (layer4_outputs(4804));
    outputs(4824) <= not((layer4_outputs(5121)) xor (layer4_outputs(4675)));
    outputs(4825) <= layer4_outputs(4949);
    outputs(4826) <= not((layer4_outputs(4464)) xor (layer4_outputs(6482)));
    outputs(4827) <= layer4_outputs(6584);
    outputs(4828) <= layer4_outputs(5028);
    outputs(4829) <= not(layer4_outputs(5503));
    outputs(4830) <= not(layer4_outputs(6770));
    outputs(4831) <= layer4_outputs(3015);
    outputs(4832) <= (layer4_outputs(491)) or (layer4_outputs(1664));
    outputs(4833) <= not(layer4_outputs(791));
    outputs(4834) <= (layer4_outputs(4824)) and not (layer4_outputs(7476));
    outputs(4835) <= (layer4_outputs(861)) and not (layer4_outputs(2576));
    outputs(4836) <= not(layer4_outputs(3504));
    outputs(4837) <= (layer4_outputs(4455)) and not (layer4_outputs(743));
    outputs(4838) <= not(layer4_outputs(33));
    outputs(4839) <= (layer4_outputs(5520)) and not (layer4_outputs(338));
    outputs(4840) <= not(layer4_outputs(975));
    outputs(4841) <= (layer4_outputs(7201)) xor (layer4_outputs(4959));
    outputs(4842) <= not(layer4_outputs(1224));
    outputs(4843) <= (layer4_outputs(7285)) and not (layer4_outputs(5909));
    outputs(4844) <= layer4_outputs(553);
    outputs(4845) <= not(layer4_outputs(4487));
    outputs(4846) <= not(layer4_outputs(426));
    outputs(4847) <= not(layer4_outputs(2559));
    outputs(4848) <= layer4_outputs(1336);
    outputs(4849) <= layer4_outputs(7194);
    outputs(4850) <= (layer4_outputs(2888)) xor (layer4_outputs(4210));
    outputs(4851) <= layer4_outputs(1090);
    outputs(4852) <= (layer4_outputs(4426)) and (layer4_outputs(670));
    outputs(4853) <= not(layer4_outputs(6530));
    outputs(4854) <= layer4_outputs(7285);
    outputs(4855) <= not((layer4_outputs(683)) or (layer4_outputs(2444)));
    outputs(4856) <= layer4_outputs(49);
    outputs(4857) <= (layer4_outputs(3346)) and not (layer4_outputs(6005));
    outputs(4858) <= not((layer4_outputs(561)) or (layer4_outputs(5971)));
    outputs(4859) <= not(layer4_outputs(7269));
    outputs(4860) <= not((layer4_outputs(1299)) or (layer4_outputs(2713)));
    outputs(4861) <= not(layer4_outputs(4280)) or (layer4_outputs(6809));
    outputs(4862) <= not(layer4_outputs(1145));
    outputs(4863) <= not((layer4_outputs(3258)) or (layer4_outputs(2969)));
    outputs(4864) <= (layer4_outputs(698)) and not (layer4_outputs(2338));
    outputs(4865) <= (layer4_outputs(6280)) xor (layer4_outputs(4834));
    outputs(4866) <= layer4_outputs(1021);
    outputs(4867) <= not(layer4_outputs(1272));
    outputs(4868) <= not(layer4_outputs(6269));
    outputs(4869) <= layer4_outputs(1634);
    outputs(4870) <= not(layer4_outputs(6933));
    outputs(4871) <= layer4_outputs(2663);
    outputs(4872) <= not((layer4_outputs(2808)) and (layer4_outputs(3763)));
    outputs(4873) <= layer4_outputs(3106);
    outputs(4874) <= not(layer4_outputs(6448));
    outputs(4875) <= (layer4_outputs(1294)) xor (layer4_outputs(6841));
    outputs(4876) <= (layer4_outputs(2927)) xor (layer4_outputs(4257));
    outputs(4877) <= (layer4_outputs(113)) and not (layer4_outputs(5279));
    outputs(4878) <= not(layer4_outputs(4584));
    outputs(4879) <= not((layer4_outputs(423)) xor (layer4_outputs(298)));
    outputs(4880) <= not((layer4_outputs(209)) or (layer4_outputs(5640)));
    outputs(4881) <= not((layer4_outputs(2030)) and (layer4_outputs(2051)));
    outputs(4882) <= layer4_outputs(5036);
    outputs(4883) <= layer4_outputs(2533);
    outputs(4884) <= not(layer4_outputs(948));
    outputs(4885) <= layer4_outputs(6305);
    outputs(4886) <= (layer4_outputs(6160)) and (layer4_outputs(4585));
    outputs(4887) <= layer4_outputs(765);
    outputs(4888) <= not(layer4_outputs(2367));
    outputs(4889) <= layer4_outputs(2194);
    outputs(4890) <= not(layer4_outputs(4052));
    outputs(4891) <= (layer4_outputs(3309)) and (layer4_outputs(605));
    outputs(4892) <= (layer4_outputs(6084)) and not (layer4_outputs(1490));
    outputs(4893) <= not(layer4_outputs(2770));
    outputs(4894) <= layer4_outputs(6157);
    outputs(4895) <= layer4_outputs(6290);
    outputs(4896) <= not((layer4_outputs(4936)) and (layer4_outputs(6213)));
    outputs(4897) <= (layer4_outputs(4220)) and not (layer4_outputs(3840));
    outputs(4898) <= not(layer4_outputs(499));
    outputs(4899) <= not((layer4_outputs(379)) xor (layer4_outputs(3290)));
    outputs(4900) <= not(layer4_outputs(5123));
    outputs(4901) <= layer4_outputs(1277);
    outputs(4902) <= layer4_outputs(979);
    outputs(4903) <= not(layer4_outputs(754));
    outputs(4904) <= layer4_outputs(5888);
    outputs(4905) <= layer4_outputs(7322);
    outputs(4906) <= layer4_outputs(5922);
    outputs(4907) <= layer4_outputs(996);
    outputs(4908) <= not(layer4_outputs(1669));
    outputs(4909) <= not(layer4_outputs(6982));
    outputs(4910) <= (layer4_outputs(6118)) and not (layer4_outputs(1054));
    outputs(4911) <= not((layer4_outputs(5313)) and (layer4_outputs(5456)));
    outputs(4912) <= (layer4_outputs(2776)) and not (layer4_outputs(3152));
    outputs(4913) <= not((layer4_outputs(7553)) or (layer4_outputs(2173)));
    outputs(4914) <= layer4_outputs(7619);
    outputs(4915) <= not((layer4_outputs(2491)) or (layer4_outputs(1767)));
    outputs(4916) <= not(layer4_outputs(7207));
    outputs(4917) <= not(layer4_outputs(721));
    outputs(4918) <= not(layer4_outputs(1373));
    outputs(4919) <= not((layer4_outputs(4151)) xor (layer4_outputs(1374)));
    outputs(4920) <= not(layer4_outputs(6034));
    outputs(4921) <= layer4_outputs(1672);
    outputs(4922) <= not(layer4_outputs(972));
    outputs(4923) <= (layer4_outputs(4854)) xor (layer4_outputs(5427));
    outputs(4924) <= not(layer4_outputs(6095));
    outputs(4925) <= (layer4_outputs(1687)) and (layer4_outputs(5422));
    outputs(4926) <= layer4_outputs(212);
    outputs(4927) <= not(layer4_outputs(2687));
    outputs(4928) <= layer4_outputs(1818);
    outputs(4929) <= not((layer4_outputs(3457)) xor (layer4_outputs(4914)));
    outputs(4930) <= not(layer4_outputs(5269));
    outputs(4931) <= not((layer4_outputs(4998)) xor (layer4_outputs(3647)));
    outputs(4932) <= layer4_outputs(2709);
    outputs(4933) <= layer4_outputs(629);
    outputs(4934) <= not((layer4_outputs(237)) xor (layer4_outputs(5951)));
    outputs(4935) <= layer4_outputs(1865);
    outputs(4936) <= (layer4_outputs(7278)) and not (layer4_outputs(6529));
    outputs(4937) <= not(layer4_outputs(1725));
    outputs(4938) <= layer4_outputs(3448);
    outputs(4939) <= not((layer4_outputs(402)) and (layer4_outputs(6729)));
    outputs(4940) <= layer4_outputs(2122);
    outputs(4941) <= not(layer4_outputs(6458));
    outputs(4942) <= not((layer4_outputs(6342)) or (layer4_outputs(4315)));
    outputs(4943) <= not(layer4_outputs(1718));
    outputs(4944) <= not(layer4_outputs(2799));
    outputs(4945) <= (layer4_outputs(2829)) and not (layer4_outputs(4161));
    outputs(4946) <= not((layer4_outputs(468)) xor (layer4_outputs(7312)));
    outputs(4947) <= not((layer4_outputs(3950)) and (layer4_outputs(6888)));
    outputs(4948) <= not(layer4_outputs(5426));
    outputs(4949) <= layer4_outputs(1309);
    outputs(4950) <= layer4_outputs(1300);
    outputs(4951) <= layer4_outputs(2535);
    outputs(4952) <= (layer4_outputs(3083)) and not (layer4_outputs(7338));
    outputs(4953) <= layer4_outputs(5843);
    outputs(4954) <= (layer4_outputs(1925)) xor (layer4_outputs(4253));
    outputs(4955) <= not(layer4_outputs(793));
    outputs(4956) <= layer4_outputs(3328);
    outputs(4957) <= layer4_outputs(557);
    outputs(4958) <= not(layer4_outputs(1129));
    outputs(4959) <= (layer4_outputs(7030)) and not (layer4_outputs(4638));
    outputs(4960) <= not(layer4_outputs(3844));
    outputs(4961) <= (layer4_outputs(569)) or (layer4_outputs(4384));
    outputs(4962) <= layer4_outputs(6805);
    outputs(4963) <= not((layer4_outputs(3536)) xor (layer4_outputs(3815)));
    outputs(4964) <= layer4_outputs(3941);
    outputs(4965) <= not(layer4_outputs(1526));
    outputs(4966) <= layer4_outputs(6979);
    outputs(4967) <= (layer4_outputs(2690)) xor (layer4_outputs(2115));
    outputs(4968) <= not(layer4_outputs(1331));
    outputs(4969) <= (layer4_outputs(3918)) xor (layer4_outputs(6571));
    outputs(4970) <= not((layer4_outputs(7435)) xor (layer4_outputs(2133)));
    outputs(4971) <= (layer4_outputs(1891)) and not (layer4_outputs(6204));
    outputs(4972) <= layer4_outputs(7072);
    outputs(4973) <= not((layer4_outputs(631)) or (layer4_outputs(4093)));
    outputs(4974) <= not(layer4_outputs(791));
    outputs(4975) <= layer4_outputs(3090);
    outputs(4976) <= layer4_outputs(2810);
    outputs(4977) <= not(layer4_outputs(5609));
    outputs(4978) <= layer4_outputs(3390);
    outputs(4979) <= not(layer4_outputs(3283));
    outputs(4980) <= not((layer4_outputs(2208)) or (layer4_outputs(3681)));
    outputs(4981) <= not((layer4_outputs(6615)) xor (layer4_outputs(4608)));
    outputs(4982) <= not(layer4_outputs(1821));
    outputs(4983) <= (layer4_outputs(7045)) and not (layer4_outputs(3580));
    outputs(4984) <= (layer4_outputs(2013)) and (layer4_outputs(5827));
    outputs(4985) <= layer4_outputs(3225);
    outputs(4986) <= not(layer4_outputs(5554));
    outputs(4987) <= layer4_outputs(5847);
    outputs(4988) <= not(layer4_outputs(1885));
    outputs(4989) <= not(layer4_outputs(2627));
    outputs(4990) <= layer4_outputs(852);
    outputs(4991) <= (layer4_outputs(4129)) and (layer4_outputs(7454));
    outputs(4992) <= not((layer4_outputs(2191)) or (layer4_outputs(5676)));
    outputs(4993) <= not((layer4_outputs(2750)) and (layer4_outputs(2525)));
    outputs(4994) <= not((layer4_outputs(2066)) xor (layer4_outputs(6344)));
    outputs(4995) <= not(layer4_outputs(958));
    outputs(4996) <= not((layer4_outputs(5049)) xor (layer4_outputs(1774)));
    outputs(4997) <= layer4_outputs(5286);
    outputs(4998) <= (layer4_outputs(214)) xor (layer4_outputs(787));
    outputs(4999) <= (layer4_outputs(4738)) xor (layer4_outputs(444));
    outputs(5000) <= (layer4_outputs(428)) xor (layer4_outputs(7533));
    outputs(5001) <= not(layer4_outputs(121));
    outputs(5002) <= not((layer4_outputs(5501)) xor (layer4_outputs(5163)));
    outputs(5003) <= not(layer4_outputs(1380));
    outputs(5004) <= layer4_outputs(4408);
    outputs(5005) <= not(layer4_outputs(5900));
    outputs(5006) <= layer4_outputs(4882);
    outputs(5007) <= not(layer4_outputs(3575));
    outputs(5008) <= (layer4_outputs(4798)) xor (layer4_outputs(3086));
    outputs(5009) <= not(layer4_outputs(6996));
    outputs(5010) <= layer4_outputs(4290);
    outputs(5011) <= (layer4_outputs(5312)) xor (layer4_outputs(5939));
    outputs(5012) <= not(layer4_outputs(6427));
    outputs(5013) <= layer4_outputs(5743);
    outputs(5014) <= not(layer4_outputs(957));
    outputs(5015) <= not(layer4_outputs(6039));
    outputs(5016) <= not(layer4_outputs(4309));
    outputs(5017) <= not(layer4_outputs(7556));
    outputs(5018) <= not(layer4_outputs(1356));
    outputs(5019) <= layer4_outputs(6008);
    outputs(5020) <= layer4_outputs(4681);
    outputs(5021) <= (layer4_outputs(3878)) xor (layer4_outputs(1798));
    outputs(5022) <= (layer4_outputs(3683)) xor (layer4_outputs(4920));
    outputs(5023) <= not(layer4_outputs(2289));
    outputs(5024) <= (layer4_outputs(2794)) xor (layer4_outputs(3153));
    outputs(5025) <= layer4_outputs(963);
    outputs(5026) <= not(layer4_outputs(7504));
    outputs(5027) <= not(layer4_outputs(584));
    outputs(5028) <= layer4_outputs(1478);
    outputs(5029) <= (layer4_outputs(7657)) xor (layer4_outputs(6333));
    outputs(5030) <= (layer4_outputs(4144)) and not (layer4_outputs(4855));
    outputs(5031) <= layer4_outputs(3478);
    outputs(5032) <= layer4_outputs(3734);
    outputs(5033) <= layer4_outputs(2532);
    outputs(5034) <= (layer4_outputs(1995)) and not (layer4_outputs(6402));
    outputs(5035) <= not(layer4_outputs(7234));
    outputs(5036) <= layer4_outputs(4419);
    outputs(5037) <= not(layer4_outputs(2501));
    outputs(5038) <= (layer4_outputs(4397)) and (layer4_outputs(3987));
    outputs(5039) <= layer4_outputs(4290);
    outputs(5040) <= not(layer4_outputs(6212));
    outputs(5041) <= (layer4_outputs(6493)) and (layer4_outputs(4980));
    outputs(5042) <= not((layer4_outputs(29)) or (layer4_outputs(1111)));
    outputs(5043) <= layer4_outputs(2819);
    outputs(5044) <= layer4_outputs(1870);
    outputs(5045) <= layer4_outputs(2468);
    outputs(5046) <= not(layer4_outputs(5794));
    outputs(5047) <= layer4_outputs(228);
    outputs(5048) <= not(layer4_outputs(4125));
    outputs(5049) <= not(layer4_outputs(592));
    outputs(5050) <= (layer4_outputs(3692)) xor (layer4_outputs(3544));
    outputs(5051) <= not(layer4_outputs(1939));
    outputs(5052) <= layer4_outputs(76);
    outputs(5053) <= layer4_outputs(3599);
    outputs(5054) <= layer4_outputs(2856);
    outputs(5055) <= not(layer4_outputs(4000));
    outputs(5056) <= not((layer4_outputs(3951)) or (layer4_outputs(1350)));
    outputs(5057) <= (layer4_outputs(5467)) and not (layer4_outputs(5569));
    outputs(5058) <= (layer4_outputs(4586)) and not (layer4_outputs(6899));
    outputs(5059) <= not((layer4_outputs(7388)) xor (layer4_outputs(1847)));
    outputs(5060) <= layer4_outputs(2831);
    outputs(5061) <= not(layer4_outputs(1678));
    outputs(5062) <= not((layer4_outputs(3237)) xor (layer4_outputs(1154)));
    outputs(5063) <= not(layer4_outputs(2908));
    outputs(5064) <= layer4_outputs(5702);
    outputs(5065) <= not(layer4_outputs(2188));
    outputs(5066) <= not((layer4_outputs(6978)) xor (layer4_outputs(2148)));
    outputs(5067) <= layer4_outputs(5316);
    outputs(5068) <= not((layer4_outputs(7597)) or (layer4_outputs(184)));
    outputs(5069) <= layer4_outputs(154);
    outputs(5070) <= layer4_outputs(1464);
    outputs(5071) <= (layer4_outputs(6022)) xor (layer4_outputs(3920));
    outputs(5072) <= layer4_outputs(2676);
    outputs(5073) <= not((layer4_outputs(2858)) xor (layer4_outputs(4229)));
    outputs(5074) <= (layer4_outputs(2175)) and not (layer4_outputs(4286));
    outputs(5075) <= not((layer4_outputs(227)) xor (layer4_outputs(2134)));
    outputs(5076) <= layer4_outputs(6050);
    outputs(5077) <= (layer4_outputs(815)) xor (layer4_outputs(7183));
    outputs(5078) <= layer4_outputs(919);
    outputs(5079) <= layer4_outputs(6674);
    outputs(5080) <= layer4_outputs(5696);
    outputs(5081) <= layer4_outputs(5171);
    outputs(5082) <= layer4_outputs(4901);
    outputs(5083) <= not(layer4_outputs(422));
    outputs(5084) <= not(layer4_outputs(5998));
    outputs(5085) <= layer4_outputs(4347);
    outputs(5086) <= not((layer4_outputs(1733)) and (layer4_outputs(2394)));
    outputs(5087) <= not(layer4_outputs(1855));
    outputs(5088) <= not(layer4_outputs(4264));
    outputs(5089) <= layer4_outputs(4306);
    outputs(5090) <= not(layer4_outputs(5420));
    outputs(5091) <= not(layer4_outputs(2543)) or (layer4_outputs(1170));
    outputs(5092) <= layer4_outputs(2936);
    outputs(5093) <= layer4_outputs(7253);
    outputs(5094) <= not((layer4_outputs(6372)) xor (layer4_outputs(7545)));
    outputs(5095) <= not(layer4_outputs(294));
    outputs(5096) <= layer4_outputs(6539);
    outputs(5097) <= layer4_outputs(6893);
    outputs(5098) <= not(layer4_outputs(1883));
    outputs(5099) <= layer4_outputs(7080);
    outputs(5100) <= not((layer4_outputs(1510)) xor (layer4_outputs(2725)));
    outputs(5101) <= not(layer4_outputs(4372));
    outputs(5102) <= layer4_outputs(1267);
    outputs(5103) <= (layer4_outputs(5382)) or (layer4_outputs(3919));
    outputs(5104) <= not(layer4_outputs(5091));
    outputs(5105) <= not(layer4_outputs(3834));
    outputs(5106) <= layer4_outputs(2287);
    outputs(5107) <= layer4_outputs(4167);
    outputs(5108) <= layer4_outputs(3358);
    outputs(5109) <= layer4_outputs(7181);
    outputs(5110) <= layer4_outputs(4969);
    outputs(5111) <= (layer4_outputs(6648)) and not (layer4_outputs(7556));
    outputs(5112) <= not(layer4_outputs(1806));
    outputs(5113) <= layer4_outputs(7212);
    outputs(5114) <= not(layer4_outputs(2830));
    outputs(5115) <= not((layer4_outputs(4214)) xor (layer4_outputs(2440)));
    outputs(5116) <= not((layer4_outputs(628)) and (layer4_outputs(2989)));
    outputs(5117) <= not(layer4_outputs(5434));
    outputs(5118) <= layer4_outputs(4737);
    outputs(5119) <= not(layer4_outputs(3930));
    outputs(5120) <= layer4_outputs(2757);
    outputs(5121) <= not(layer4_outputs(2677));
    outputs(5122) <= layer4_outputs(5448);
    outputs(5123) <= layer4_outputs(6479);
    outputs(5124) <= not(layer4_outputs(6970));
    outputs(5125) <= not(layer4_outputs(3471));
    outputs(5126) <= (layer4_outputs(5028)) xor (layer4_outputs(5214));
    outputs(5127) <= (layer4_outputs(5614)) and not (layer4_outputs(7287));
    outputs(5128) <= layer4_outputs(4828);
    outputs(5129) <= not(layer4_outputs(1864));
    outputs(5130) <= (layer4_outputs(6279)) xor (layer4_outputs(7009));
    outputs(5131) <= layer4_outputs(7118);
    outputs(5132) <= layer4_outputs(6431);
    outputs(5133) <= layer4_outputs(2102);
    outputs(5134) <= layer4_outputs(3020);
    outputs(5135) <= not(layer4_outputs(6377)) or (layer4_outputs(6934));
    outputs(5136) <= not((layer4_outputs(2601)) xor (layer4_outputs(5965)));
    outputs(5137) <= not((layer4_outputs(6388)) xor (layer4_outputs(7172)));
    outputs(5138) <= not(layer4_outputs(1987));
    outputs(5139) <= not(layer4_outputs(508));
    outputs(5140) <= (layer4_outputs(2965)) xor (layer4_outputs(6097));
    outputs(5141) <= not(layer4_outputs(6261));
    outputs(5142) <= layer4_outputs(1758);
    outputs(5143) <= not((layer4_outputs(400)) xor (layer4_outputs(6160)));
    outputs(5144) <= layer4_outputs(5598);
    outputs(5145) <= layer4_outputs(397);
    outputs(5146) <= not((layer4_outputs(6817)) and (layer4_outputs(5688)));
    outputs(5147) <= not(layer4_outputs(5246));
    outputs(5148) <= (layer4_outputs(5004)) and not (layer4_outputs(5022));
    outputs(5149) <= layer4_outputs(5375);
    outputs(5150) <= not(layer4_outputs(846));
    outputs(5151) <= (layer4_outputs(132)) xor (layer4_outputs(6102));
    outputs(5152) <= not(layer4_outputs(5419));
    outputs(5153) <= layer4_outputs(5602);
    outputs(5154) <= (layer4_outputs(6487)) xor (layer4_outputs(1488));
    outputs(5155) <= (layer4_outputs(4964)) and not (layer4_outputs(1992));
    outputs(5156) <= (layer4_outputs(6509)) and not (layer4_outputs(3093));
    outputs(5157) <= not(layer4_outputs(671));
    outputs(5158) <= layer4_outputs(5132);
    outputs(5159) <= layer4_outputs(2461);
    outputs(5160) <= not(layer4_outputs(3782));
    outputs(5161) <= not(layer4_outputs(6522));
    outputs(5162) <= not((layer4_outputs(2182)) and (layer4_outputs(3138)));
    outputs(5163) <= (layer4_outputs(6589)) xor (layer4_outputs(6577));
    outputs(5164) <= layer4_outputs(6205);
    outputs(5165) <= layer4_outputs(4203);
    outputs(5166) <= not(layer4_outputs(6031));
    outputs(5167) <= layer4_outputs(4495);
    outputs(5168) <= not((layer4_outputs(2041)) and (layer4_outputs(5481)));
    outputs(5169) <= (layer4_outputs(5457)) or (layer4_outputs(3117));
    outputs(5170) <= layer4_outputs(3640);
    outputs(5171) <= layer4_outputs(3395);
    outputs(5172) <= not(layer4_outputs(1125));
    outputs(5173) <= (layer4_outputs(5790)) and not (layer4_outputs(335));
    outputs(5174) <= (layer4_outputs(113)) and not (layer4_outputs(6134));
    outputs(5175) <= (layer4_outputs(7143)) xor (layer4_outputs(4813));
    outputs(5176) <= not(layer4_outputs(3169));
    outputs(5177) <= layer4_outputs(2582);
    outputs(5178) <= not(layer4_outputs(2877));
    outputs(5179) <= layer4_outputs(2322);
    outputs(5180) <= layer4_outputs(5271);
    outputs(5181) <= not((layer4_outputs(1183)) xor (layer4_outputs(7510)));
    outputs(5182) <= (layer4_outputs(7447)) and (layer4_outputs(4137));
    outputs(5183) <= not(layer4_outputs(3777));
    outputs(5184) <= not(layer4_outputs(2624));
    outputs(5185) <= not(layer4_outputs(4849)) or (layer4_outputs(5395));
    outputs(5186) <= not(layer4_outputs(6396));
    outputs(5187) <= not((layer4_outputs(5730)) and (layer4_outputs(259)));
    outputs(5188) <= layer4_outputs(1833);
    outputs(5189) <= layer4_outputs(2082);
    outputs(5190) <= not(layer4_outputs(6323));
    outputs(5191) <= not(layer4_outputs(2245));
    outputs(5192) <= not(layer4_outputs(3204));
    outputs(5193) <= not(layer4_outputs(2737));
    outputs(5194) <= (layer4_outputs(3102)) and not (layer4_outputs(5087));
    outputs(5195) <= not(layer4_outputs(7478));
    outputs(5196) <= (layer4_outputs(2729)) and (layer4_outputs(5197));
    outputs(5197) <= (layer4_outputs(5578)) and (layer4_outputs(4842));
    outputs(5198) <= not(layer4_outputs(468));
    outputs(5199) <= not(layer4_outputs(6819));
    outputs(5200) <= not(layer4_outputs(6128));
    outputs(5201) <= layer4_outputs(1315);
    outputs(5202) <= layer4_outputs(1172);
    outputs(5203) <= layer4_outputs(6825);
    outputs(5204) <= layer4_outputs(5113);
    outputs(5205) <= not(layer4_outputs(3964));
    outputs(5206) <= not(layer4_outputs(4944));
    outputs(5207) <= (layer4_outputs(3827)) and (layer4_outputs(5359));
    outputs(5208) <= not(layer4_outputs(5871));
    outputs(5209) <= (layer4_outputs(1259)) xor (layer4_outputs(1480));
    outputs(5210) <= not(layer4_outputs(6625));
    outputs(5211) <= not(layer4_outputs(6859)) or (layer4_outputs(1076));
    outputs(5212) <= (layer4_outputs(2697)) and not (layer4_outputs(2473));
    outputs(5213) <= not((layer4_outputs(845)) xor (layer4_outputs(3714)));
    outputs(5214) <= not(layer4_outputs(5732));
    outputs(5215) <= layer4_outputs(553);
    outputs(5216) <= not((layer4_outputs(2957)) xor (layer4_outputs(2105)));
    outputs(5217) <= not(layer4_outputs(2351));
    outputs(5218) <= (layer4_outputs(3328)) and not (layer4_outputs(1167));
    outputs(5219) <= (layer4_outputs(6534)) and (layer4_outputs(4206));
    outputs(5220) <= layer4_outputs(3516);
    outputs(5221) <= not((layer4_outputs(5874)) xor (layer4_outputs(5775)));
    outputs(5222) <= not(layer4_outputs(7473));
    outputs(5223) <= (layer4_outputs(6877)) xor (layer4_outputs(4697));
    outputs(5224) <= (layer4_outputs(3078)) xor (layer4_outputs(6816));
    outputs(5225) <= not(layer4_outputs(7465)) or (layer4_outputs(1676));
    outputs(5226) <= layer4_outputs(7146);
    outputs(5227) <= not(layer4_outputs(7394)) or (layer4_outputs(3820));
    outputs(5228) <= not(layer4_outputs(5709));
    outputs(5229) <= not(layer4_outputs(7005)) or (layer4_outputs(3972));
    outputs(5230) <= not(layer4_outputs(1795));
    outputs(5231) <= not(layer4_outputs(2301));
    outputs(5232) <= (layer4_outputs(2863)) xor (layer4_outputs(6088));
    outputs(5233) <= layer4_outputs(4472);
    outputs(5234) <= layer4_outputs(4571);
    outputs(5235) <= not(layer4_outputs(2006));
    outputs(5236) <= not(layer4_outputs(4042));
    outputs(5237) <= layer4_outputs(7225);
    outputs(5238) <= not(layer4_outputs(6981));
    outputs(5239) <= (layer4_outputs(4817)) xor (layer4_outputs(3811));
    outputs(5240) <= not(layer4_outputs(1713));
    outputs(5241) <= layer4_outputs(5580);
    outputs(5242) <= not((layer4_outputs(4265)) or (layer4_outputs(1847)));
    outputs(5243) <= layer4_outputs(996);
    outputs(5244) <= not(layer4_outputs(5390));
    outputs(5245) <= layer4_outputs(3292);
    outputs(5246) <= not(layer4_outputs(4702)) or (layer4_outputs(3689));
    outputs(5247) <= layer4_outputs(7470);
    outputs(5248) <= layer4_outputs(4633);
    outputs(5249) <= (layer4_outputs(986)) and not (layer4_outputs(4812));
    outputs(5250) <= not(layer4_outputs(3950));
    outputs(5251) <= not(layer4_outputs(2393));
    outputs(5252) <= layer4_outputs(1877);
    outputs(5253) <= not((layer4_outputs(4155)) xor (layer4_outputs(3809)));
    outputs(5254) <= layer4_outputs(3691);
    outputs(5255) <= not(layer4_outputs(2270)) or (layer4_outputs(2960));
    outputs(5256) <= (layer4_outputs(1392)) and (layer4_outputs(7177));
    outputs(5257) <= not((layer4_outputs(2437)) xor (layer4_outputs(6994)));
    outputs(5258) <= (layer4_outputs(7668)) and not (layer4_outputs(1412));
    outputs(5259) <= not(layer4_outputs(137)) or (layer4_outputs(5779));
    outputs(5260) <= layer4_outputs(275);
    outputs(5261) <= layer4_outputs(4633);
    outputs(5262) <= layer4_outputs(2453);
    outputs(5263) <= (layer4_outputs(317)) xor (layer4_outputs(5326));
    outputs(5264) <= layer4_outputs(7288);
    outputs(5265) <= not((layer4_outputs(4047)) or (layer4_outputs(4536)));
    outputs(5266) <= layer4_outputs(5995);
    outputs(5267) <= not((layer4_outputs(4413)) xor (layer4_outputs(1958)));
    outputs(5268) <= not(layer4_outputs(2775));
    outputs(5269) <= not(layer4_outputs(1037));
    outputs(5270) <= layer4_outputs(6161);
    outputs(5271) <= not(layer4_outputs(7571));
    outputs(5272) <= not(layer4_outputs(5495));
    outputs(5273) <= layer4_outputs(1618);
    outputs(5274) <= (layer4_outputs(825)) and (layer4_outputs(3790));
    outputs(5275) <= layer4_outputs(3850);
    outputs(5276) <= layer4_outputs(5110);
    outputs(5277) <= not(layer4_outputs(3656));
    outputs(5278) <= not(layer4_outputs(6490));
    outputs(5279) <= not((layer4_outputs(3229)) xor (layer4_outputs(6885)));
    outputs(5280) <= (layer4_outputs(3046)) and not (layer4_outputs(3908));
    outputs(5281) <= not((layer4_outputs(2853)) or (layer4_outputs(6356)));
    outputs(5282) <= layer4_outputs(7135);
    outputs(5283) <= not((layer4_outputs(6416)) xor (layer4_outputs(7292)));
    outputs(5284) <= not(layer4_outputs(6749));
    outputs(5285) <= layer4_outputs(7678);
    outputs(5286) <= layer4_outputs(5777);
    outputs(5287) <= (layer4_outputs(7099)) and (layer4_outputs(1077));
    outputs(5288) <= not(layer4_outputs(4645)) or (layer4_outputs(4489));
    outputs(5289) <= not(layer4_outputs(6458));
    outputs(5290) <= not((layer4_outputs(2818)) or (layer4_outputs(3872)));
    outputs(5291) <= not((layer4_outputs(5230)) xor (layer4_outputs(3035)));
    outputs(5292) <= (layer4_outputs(5876)) and not (layer4_outputs(4207));
    outputs(5293) <= not((layer4_outputs(1974)) or (layer4_outputs(2207)));
    outputs(5294) <= not(layer4_outputs(2403));
    outputs(5295) <= (layer4_outputs(5785)) and not (layer4_outputs(7277));
    outputs(5296) <= (layer4_outputs(714)) or (layer4_outputs(6740));
    outputs(5297) <= (layer4_outputs(1592)) xor (layer4_outputs(5186));
    outputs(5298) <= not(layer4_outputs(6388));
    outputs(5299) <= layer4_outputs(1325);
    outputs(5300) <= layer4_outputs(4057);
    outputs(5301) <= (layer4_outputs(1240)) and (layer4_outputs(2876));
    outputs(5302) <= not(layer4_outputs(2314));
    outputs(5303) <= layer4_outputs(3376);
    outputs(5304) <= not(layer4_outputs(6508));
    outputs(5305) <= not(layer4_outputs(1196));
    outputs(5306) <= not(layer4_outputs(6808));
    outputs(5307) <= (layer4_outputs(4693)) or (layer4_outputs(6848));
    outputs(5308) <= (layer4_outputs(4140)) and (layer4_outputs(4296));
    outputs(5309) <= not(layer4_outputs(2518));
    outputs(5310) <= layer4_outputs(2891);
    outputs(5311) <= not(layer4_outputs(4567));
    outputs(5312) <= (layer4_outputs(6650)) xor (layer4_outputs(48));
    outputs(5313) <= (layer4_outputs(5366)) xor (layer4_outputs(5224));
    outputs(5314) <= (layer4_outputs(4949)) and not (layer4_outputs(5522));
    outputs(5315) <= layer4_outputs(3842);
    outputs(5316) <= not((layer4_outputs(6087)) xor (layer4_outputs(3652)));
    outputs(5317) <= layer4_outputs(6693);
    outputs(5318) <= layer4_outputs(351);
    outputs(5319) <= not(layer4_outputs(6459));
    outputs(5320) <= not(layer4_outputs(4711));
    outputs(5321) <= (layer4_outputs(3373)) and not (layer4_outputs(4028));
    outputs(5322) <= not((layer4_outputs(96)) xor (layer4_outputs(3304)));
    outputs(5323) <= (layer4_outputs(4986)) xor (layer4_outputs(2997));
    outputs(5324) <= layer4_outputs(6681);
    outputs(5325) <= layer4_outputs(4131);
    outputs(5326) <= not(layer4_outputs(2067));
    outputs(5327) <= layer4_outputs(2209);
    outputs(5328) <= not(layer4_outputs(6577));
    outputs(5329) <= layer4_outputs(5298);
    outputs(5330) <= layer4_outputs(2312);
    outputs(5331) <= (layer4_outputs(5537)) and not (layer4_outputs(5211));
    outputs(5332) <= (layer4_outputs(2465)) or (layer4_outputs(4366));
    outputs(5333) <= (layer4_outputs(5938)) and (layer4_outputs(1017));
    outputs(5334) <= layer4_outputs(2104);
    outputs(5335) <= layer4_outputs(4718);
    outputs(5336) <= not(layer4_outputs(1193));
    outputs(5337) <= (layer4_outputs(3968)) xor (layer4_outputs(2567));
    outputs(5338) <= (layer4_outputs(2455)) xor (layer4_outputs(3290));
    outputs(5339) <= layer4_outputs(4110);
    outputs(5340) <= not(layer4_outputs(2205));
    outputs(5341) <= not(layer4_outputs(2130));
    outputs(5342) <= layer4_outputs(2498);
    outputs(5343) <= layer4_outputs(2312);
    outputs(5344) <= layer4_outputs(6278);
    outputs(5345) <= (layer4_outputs(4361)) and not (layer4_outputs(5607));
    outputs(5346) <= not(layer4_outputs(554));
    outputs(5347) <= not(layer4_outputs(616)) or (layer4_outputs(644));
    outputs(5348) <= not(layer4_outputs(2056));
    outputs(5349) <= layer4_outputs(3863);
    outputs(5350) <= (layer4_outputs(1819)) xor (layer4_outputs(1914));
    outputs(5351) <= not((layer4_outputs(1595)) xor (layer4_outputs(352)));
    outputs(5352) <= not(layer4_outputs(3391));
    outputs(5353) <= (layer4_outputs(6911)) or (layer4_outputs(3530));
    outputs(5354) <= not(layer4_outputs(4963));
    outputs(5355) <= not(layer4_outputs(4871));
    outputs(5356) <= (layer4_outputs(2230)) and (layer4_outputs(1633));
    outputs(5357) <= not(layer4_outputs(1710)) or (layer4_outputs(4428));
    outputs(5358) <= layer4_outputs(3992);
    outputs(5359) <= layer4_outputs(5158);
    outputs(5360) <= not(layer4_outputs(2008));
    outputs(5361) <= layer4_outputs(4722);
    outputs(5362) <= layer4_outputs(4901);
    outputs(5363) <= not(layer4_outputs(1223));
    outputs(5364) <= layer4_outputs(7655);
    outputs(5365) <= not((layer4_outputs(2078)) xor (layer4_outputs(287)));
    outputs(5366) <= not((layer4_outputs(4960)) or (layer4_outputs(7563)));
    outputs(5367) <= layer4_outputs(6098);
    outputs(5368) <= not((layer4_outputs(5697)) xor (layer4_outputs(6330)));
    outputs(5369) <= not((layer4_outputs(271)) xor (layer4_outputs(5922)));
    outputs(5370) <= not((layer4_outputs(5121)) xor (layer4_outputs(6627)));
    outputs(5371) <= layer4_outputs(4254);
    outputs(5372) <= layer4_outputs(2415);
    outputs(5373) <= (layer4_outputs(420)) and (layer4_outputs(492));
    outputs(5374) <= not(layer4_outputs(5747)) or (layer4_outputs(3810));
    outputs(5375) <= not((layer4_outputs(2226)) or (layer4_outputs(6877)));
    outputs(5376) <= (layer4_outputs(6617)) xor (layer4_outputs(5553));
    outputs(5377) <= layer4_outputs(1095);
    outputs(5378) <= not(layer4_outputs(5171)) or (layer4_outputs(1671));
    outputs(5379) <= layer4_outputs(3980);
    outputs(5380) <= not(layer4_outputs(1402));
    outputs(5381) <= layer4_outputs(3617);
    outputs(5382) <= not((layer4_outputs(1333)) and (layer4_outputs(2728)));
    outputs(5383) <= not(layer4_outputs(2917));
    outputs(5384) <= (layer4_outputs(4204)) xor (layer4_outputs(4505));
    outputs(5385) <= not(layer4_outputs(2698));
    outputs(5386) <= not((layer4_outputs(2007)) and (layer4_outputs(941)));
    outputs(5387) <= (layer4_outputs(4656)) xor (layer4_outputs(1702));
    outputs(5388) <= (layer4_outputs(4974)) and not (layer4_outputs(1027));
    outputs(5389) <= (layer4_outputs(2748)) xor (layer4_outputs(1320));
    outputs(5390) <= layer4_outputs(1179);
    outputs(5391) <= layer4_outputs(1358);
    outputs(5392) <= layer4_outputs(7254);
    outputs(5393) <= (layer4_outputs(2805)) and (layer4_outputs(3884));
    outputs(5394) <= not(layer4_outputs(3339));
    outputs(5395) <= not(layer4_outputs(6599));
    outputs(5396) <= (layer4_outputs(6375)) xor (layer4_outputs(1197));
    outputs(5397) <= (layer4_outputs(1778)) xor (layer4_outputs(4976));
    outputs(5398) <= (layer4_outputs(5164)) and not (layer4_outputs(2747));
    outputs(5399) <= not(layer4_outputs(4253));
    outputs(5400) <= not(layer4_outputs(6932));
    outputs(5401) <= not(layer4_outputs(6651));
    outputs(5402) <= layer4_outputs(4564);
    outputs(5403) <= not(layer4_outputs(5485));
    outputs(5404) <= layer4_outputs(6316);
    outputs(5405) <= layer4_outputs(4066);
    outputs(5406) <= not(layer4_outputs(6324)) or (layer4_outputs(788));
    outputs(5407) <= not((layer4_outputs(3757)) or (layer4_outputs(262)));
    outputs(5408) <= not(layer4_outputs(93));
    outputs(5409) <= layer4_outputs(94);
    outputs(5410) <= not(layer4_outputs(4898));
    outputs(5411) <= layer4_outputs(5423);
    outputs(5412) <= not(layer4_outputs(7203));
    outputs(5413) <= layer4_outputs(188);
    outputs(5414) <= not(layer4_outputs(5917));
    outputs(5415) <= layer4_outputs(5136);
    outputs(5416) <= not(layer4_outputs(4486));
    outputs(5417) <= layer4_outputs(1738);
    outputs(5418) <= not(layer4_outputs(2032));
    outputs(5419) <= layer4_outputs(5488);
    outputs(5420) <= layer4_outputs(4126);
    outputs(5421) <= (layer4_outputs(3200)) xor (layer4_outputs(6637));
    outputs(5422) <= not(layer4_outputs(7331));
    outputs(5423) <= layer4_outputs(4415);
    outputs(5424) <= not((layer4_outputs(2726)) xor (layer4_outputs(4469)));
    outputs(5425) <= (layer4_outputs(1451)) and (layer4_outputs(6444));
    outputs(5426) <= layer4_outputs(5540);
    outputs(5427) <= (layer4_outputs(1006)) and (layer4_outputs(3805));
    outputs(5428) <= (layer4_outputs(2343)) and not (layer4_outputs(6498));
    outputs(5429) <= not(layer4_outputs(3948));
    outputs(5430) <= (layer4_outputs(2492)) or (layer4_outputs(2636));
    outputs(5431) <= not((layer4_outputs(4993)) xor (layer4_outputs(3738)));
    outputs(5432) <= not(layer4_outputs(1907));
    outputs(5433) <= (layer4_outputs(1487)) and (layer4_outputs(276));
    outputs(5434) <= not((layer4_outputs(5561)) and (layer4_outputs(1414)));
    outputs(5435) <= layer4_outputs(1820);
    outputs(5436) <= not(layer4_outputs(6916));
    outputs(5437) <= (layer4_outputs(2510)) xor (layer4_outputs(571));
    outputs(5438) <= not(layer4_outputs(3042));
    outputs(5439) <= (layer4_outputs(4191)) xor (layer4_outputs(7564));
    outputs(5440) <= not(layer4_outputs(1970));
    outputs(5441) <= layer4_outputs(3520);
    outputs(5442) <= (layer4_outputs(7566)) or (layer4_outputs(5559));
    outputs(5443) <= not(layer4_outputs(1758));
    outputs(5444) <= not(layer4_outputs(2276));
    outputs(5445) <= not(layer4_outputs(6250));
    outputs(5446) <= layer4_outputs(4425);
    outputs(5447) <= layer4_outputs(3575);
    outputs(5448) <= layer4_outputs(5040);
    outputs(5449) <= not(layer4_outputs(4262));
    outputs(5450) <= not(layer4_outputs(5978)) or (layer4_outputs(7656));
    outputs(5451) <= (layer4_outputs(3054)) xor (layer4_outputs(306));
    outputs(5452) <= not((layer4_outputs(1947)) xor (layer4_outputs(5350)));
    outputs(5453) <= not(layer4_outputs(4679));
    outputs(5454) <= layer4_outputs(2579);
    outputs(5455) <= not(layer4_outputs(4867)) or (layer4_outputs(797));
    outputs(5456) <= not(layer4_outputs(2199));
    outputs(5457) <= not(layer4_outputs(497));
    outputs(5458) <= not(layer4_outputs(6474)) or (layer4_outputs(5215));
    outputs(5459) <= (layer4_outputs(6033)) xor (layer4_outputs(3345));
    outputs(5460) <= not((layer4_outputs(3608)) or (layer4_outputs(6391)));
    outputs(5461) <= not(layer4_outputs(3076));
    outputs(5462) <= layer4_outputs(1317);
    outputs(5463) <= layer4_outputs(5236);
    outputs(5464) <= layer4_outputs(2409);
    outputs(5465) <= (layer4_outputs(6926)) and not (layer4_outputs(1575));
    outputs(5466) <= not(layer4_outputs(3063));
    outputs(5467) <= not((layer4_outputs(5047)) or (layer4_outputs(5173)));
    outputs(5468) <= (layer4_outputs(5103)) xor (layer4_outputs(6771));
    outputs(5469) <= (layer4_outputs(6867)) and not (layer4_outputs(244));
    outputs(5470) <= (layer4_outputs(4611)) and (layer4_outputs(5677));
    outputs(5471) <= (layer4_outputs(4128)) xor (layer4_outputs(3716));
    outputs(5472) <= not(layer4_outputs(3759));
    outputs(5473) <= not(layer4_outputs(5494));
    outputs(5474) <= not((layer4_outputs(4709)) or (layer4_outputs(444)));
    outputs(5475) <= not(layer4_outputs(1949));
    outputs(5476) <= layer4_outputs(6408);
    outputs(5477) <= not(layer4_outputs(6015));
    outputs(5478) <= not(layer4_outputs(6547));
    outputs(5479) <= not(layer4_outputs(7335));
    outputs(5480) <= layer4_outputs(4087);
    outputs(5481) <= (layer4_outputs(868)) and not (layer4_outputs(2516));
    outputs(5482) <= not(layer4_outputs(4903));
    outputs(5483) <= not(layer4_outputs(6518));
    outputs(5484) <= layer4_outputs(2018);
    outputs(5485) <= layer4_outputs(597);
    outputs(5486) <= not(layer4_outputs(4358));
    outputs(5487) <= not(layer4_outputs(3565));
    outputs(5488) <= not((layer4_outputs(2702)) or (layer4_outputs(4325)));
    outputs(5489) <= (layer4_outputs(2233)) and (layer4_outputs(5663));
    outputs(5490) <= (layer4_outputs(570)) and not (layer4_outputs(4449));
    outputs(5491) <= not(layer4_outputs(7533)) or (layer4_outputs(4520));
    outputs(5492) <= not(layer4_outputs(3012));
    outputs(5493) <= not(layer4_outputs(3246));
    outputs(5494) <= not(layer4_outputs(556));
    outputs(5495) <= (layer4_outputs(1480)) and not (layer4_outputs(6228));
    outputs(5496) <= (layer4_outputs(7662)) and not (layer4_outputs(3813));
    outputs(5497) <= layer4_outputs(6034);
    outputs(5498) <= layer4_outputs(2413);
    outputs(5499) <= (layer4_outputs(4527)) and not (layer4_outputs(2317));
    outputs(5500) <= (layer4_outputs(579)) xor (layer4_outputs(6569));
    outputs(5501) <= not(layer4_outputs(43));
    outputs(5502) <= not(layer4_outputs(4933));
    outputs(5503) <= not(layer4_outputs(2499));
    outputs(5504) <= not(layer4_outputs(2663));
    outputs(5505) <= not((layer4_outputs(5206)) xor (layer4_outputs(3951)));
    outputs(5506) <= not(layer4_outputs(7020));
    outputs(5507) <= layer4_outputs(980);
    outputs(5508) <= (layer4_outputs(1005)) and (layer4_outputs(5196));
    outputs(5509) <= not((layer4_outputs(4452)) xor (layer4_outputs(1573)));
    outputs(5510) <= not(layer4_outputs(2092));
    outputs(5511) <= not(layer4_outputs(4892)) or (layer4_outputs(1339));
    outputs(5512) <= layer4_outputs(1466);
    outputs(5513) <= not(layer4_outputs(4982));
    outputs(5514) <= (layer4_outputs(821)) and (layer4_outputs(2943));
    outputs(5515) <= not(layer4_outputs(1483));
    outputs(5516) <= layer4_outputs(6883);
    outputs(5517) <= (layer4_outputs(2940)) and not (layer4_outputs(7202));
    outputs(5518) <= layer4_outputs(2787);
    outputs(5519) <= layer4_outputs(2314);
    outputs(5520) <= (layer4_outputs(177)) xor (layer4_outputs(1637));
    outputs(5521) <= (layer4_outputs(5104)) xor (layer4_outputs(6130));
    outputs(5522) <= not(layer4_outputs(519));
    outputs(5523) <= not((layer4_outputs(1660)) xor (layer4_outputs(4002)));
    outputs(5524) <= (layer4_outputs(1254)) and not (layer4_outputs(6574));
    outputs(5525) <= not(layer4_outputs(4232));
    outputs(5526) <= not(layer4_outputs(7091));
    outputs(5527) <= not((layer4_outputs(3891)) or (layer4_outputs(2131)));
    outputs(5528) <= (layer4_outputs(927)) and (layer4_outputs(382));
    outputs(5529) <= not((layer4_outputs(3223)) xor (layer4_outputs(5099)));
    outputs(5530) <= (layer4_outputs(4072)) and not (layer4_outputs(2324));
    outputs(5531) <= layer4_outputs(2624);
    outputs(5532) <= layer4_outputs(3556);
    outputs(5533) <= not(layer4_outputs(1835));
    outputs(5534) <= layer4_outputs(7596);
    outputs(5535) <= not((layer4_outputs(3468)) xor (layer4_outputs(3331)));
    outputs(5536) <= not(layer4_outputs(4482));
    outputs(5537) <= (layer4_outputs(5724)) or (layer4_outputs(1931));
    outputs(5538) <= not((layer4_outputs(5919)) and (layer4_outputs(4303)));
    outputs(5539) <= not((layer4_outputs(6307)) or (layer4_outputs(3687)));
    outputs(5540) <= layer4_outputs(5860);
    outputs(5541) <= (layer4_outputs(6298)) xor (layer4_outputs(6051));
    outputs(5542) <= not(layer4_outputs(3061));
    outputs(5543) <= not(layer4_outputs(5633));
    outputs(5544) <= layer4_outputs(2918);
    outputs(5545) <= not((layer4_outputs(6251)) or (layer4_outputs(613)));
    outputs(5546) <= layer4_outputs(7178);
    outputs(5547) <= layer4_outputs(1620);
    outputs(5548) <= not((layer4_outputs(3779)) or (layer4_outputs(1374)));
    outputs(5549) <= (layer4_outputs(4978)) and (layer4_outputs(4215));
    outputs(5550) <= layer4_outputs(3521);
    outputs(5551) <= not((layer4_outputs(5372)) or (layer4_outputs(7397)));
    outputs(5552) <= not((layer4_outputs(59)) or (layer4_outputs(4836)));
    outputs(5553) <= layer4_outputs(1665);
    outputs(5554) <= (layer4_outputs(2782)) and (layer4_outputs(3403));
    outputs(5555) <= layer4_outputs(3051);
    outputs(5556) <= not(layer4_outputs(5687));
    outputs(5557) <= (layer4_outputs(391)) xor (layer4_outputs(7027));
    outputs(5558) <= not(layer4_outputs(3879));
    outputs(5559) <= (layer4_outputs(849)) and (layer4_outputs(5258));
    outputs(5560) <= (layer4_outputs(3234)) xor (layer4_outputs(6977));
    outputs(5561) <= not(layer4_outputs(6786));
    outputs(5562) <= (layer4_outputs(196)) and not (layer4_outputs(6235));
    outputs(5563) <= not((layer4_outputs(5534)) xor (layer4_outputs(4902)));
    outputs(5564) <= (layer4_outputs(7540)) xor (layer4_outputs(6054));
    outputs(5565) <= not(layer4_outputs(3185));
    outputs(5566) <= not((layer4_outputs(5262)) xor (layer4_outputs(7659)));
    outputs(5567) <= layer4_outputs(2824);
    outputs(5568) <= not(layer4_outputs(3382));
    outputs(5569) <= (layer4_outputs(1313)) xor (layer4_outputs(970));
    outputs(5570) <= (layer4_outputs(2036)) and not (layer4_outputs(427));
    outputs(5571) <= not((layer4_outputs(7626)) or (layer4_outputs(875)));
    outputs(5572) <= not(layer4_outputs(1676));
    outputs(5573) <= (layer4_outputs(6309)) and (layer4_outputs(5630));
    outputs(5574) <= (layer4_outputs(5435)) and not (layer4_outputs(3553));
    outputs(5575) <= not(layer4_outputs(3386));
    outputs(5576) <= layer4_outputs(4367);
    outputs(5577) <= (layer4_outputs(543)) and not (layer4_outputs(4405));
    outputs(5578) <= layer4_outputs(185);
    outputs(5579) <= not(layer4_outputs(5995));
    outputs(5580) <= not(layer4_outputs(2974));
    outputs(5581) <= layer4_outputs(5385);
    outputs(5582) <= layer4_outputs(846);
    outputs(5583) <= (layer4_outputs(2816)) and (layer4_outputs(588));
    outputs(5584) <= layer4_outputs(6189);
    outputs(5585) <= (layer4_outputs(1413)) and not (layer4_outputs(4495));
    outputs(5586) <= layer4_outputs(1102);
    outputs(5587) <= not(layer4_outputs(2679));
    outputs(5588) <= not((layer4_outputs(3696)) or (layer4_outputs(1365)));
    outputs(5589) <= not(layer4_outputs(1672));
    outputs(5590) <= not((layer4_outputs(615)) or (layer4_outputs(5658)));
    outputs(5591) <= (layer4_outputs(7481)) and (layer4_outputs(660));
    outputs(5592) <= not(layer4_outputs(1483));
    outputs(5593) <= (layer4_outputs(3659)) and not (layer4_outputs(2606));
    outputs(5594) <= (layer4_outputs(4662)) and not (layer4_outputs(5964));
    outputs(5595) <= layer4_outputs(3295);
    outputs(5596) <= (layer4_outputs(4952)) and not (layer4_outputs(515));
    outputs(5597) <= not(layer4_outputs(977));
    outputs(5598) <= not((layer4_outputs(2574)) or (layer4_outputs(3381)));
    outputs(5599) <= not(layer4_outputs(1090));
    outputs(5600) <= (layer4_outputs(4613)) xor (layer4_outputs(2000));
    outputs(5601) <= layer4_outputs(5068);
    outputs(5602) <= layer4_outputs(3205);
    outputs(5603) <= not(layer4_outputs(6747));
    outputs(5604) <= layer4_outputs(7048);
    outputs(5605) <= (layer4_outputs(6906)) and (layer4_outputs(1553));
    outputs(5606) <= layer4_outputs(5310);
    outputs(5607) <= layer4_outputs(413);
    outputs(5608) <= not(layer4_outputs(5324));
    outputs(5609) <= layer4_outputs(4915);
    outputs(5610) <= not(layer4_outputs(4427));
    outputs(5611) <= not(layer4_outputs(2543));
    outputs(5612) <= (layer4_outputs(5670)) and not (layer4_outputs(2348));
    outputs(5613) <= not(layer4_outputs(7131));
    outputs(5614) <= (layer4_outputs(1022)) and (layer4_outputs(6413));
    outputs(5615) <= not(layer4_outputs(2255)) or (layer4_outputs(3705));
    outputs(5616) <= not(layer4_outputs(3664));
    outputs(5617) <= (layer4_outputs(5982)) or (layer4_outputs(2389));
    outputs(5618) <= layer4_outputs(3147);
    outputs(5619) <= not(layer4_outputs(7204));
    outputs(5620) <= (layer4_outputs(7524)) xor (layer4_outputs(5557));
    outputs(5621) <= not((layer4_outputs(5411)) xor (layer4_outputs(7139)));
    outputs(5622) <= not(layer4_outputs(1168));
    outputs(5623) <= (layer4_outputs(3659)) and (layer4_outputs(1071));
    outputs(5624) <= layer4_outputs(4516);
    outputs(5625) <= not((layer4_outputs(5626)) or (layer4_outputs(312)));
    outputs(5626) <= not(layer4_outputs(7409));
    outputs(5627) <= (layer4_outputs(3470)) and (layer4_outputs(2019));
    outputs(5628) <= not((layer4_outputs(7451)) xor (layer4_outputs(3375)));
    outputs(5629) <= (layer4_outputs(310)) and (layer4_outputs(5064));
    outputs(5630) <= not((layer4_outputs(6917)) xor (layer4_outputs(122)));
    outputs(5631) <= not((layer4_outputs(5348)) or (layer4_outputs(6043)));
    outputs(5632) <= not(layer4_outputs(172));
    outputs(5633) <= layer4_outputs(6268);
    outputs(5634) <= not((layer4_outputs(6481)) or (layer4_outputs(3319)));
    outputs(5635) <= (layer4_outputs(6013)) xor (layer4_outputs(7395));
    outputs(5636) <= layer4_outputs(3595);
    outputs(5637) <= (layer4_outputs(65)) and (layer4_outputs(5999));
    outputs(5638) <= layer4_outputs(4559);
    outputs(5639) <= (layer4_outputs(6188)) and (layer4_outputs(1902));
    outputs(5640) <= (layer4_outputs(6113)) and not (layer4_outputs(1225));
    outputs(5641) <= (layer4_outputs(5432)) and not (layer4_outputs(4714));
    outputs(5642) <= (layer4_outputs(1324)) and not (layer4_outputs(2975));
    outputs(5643) <= (layer4_outputs(1224)) and (layer4_outputs(3036));
    outputs(5644) <= not(layer4_outputs(266));
    outputs(5645) <= layer4_outputs(5461);
    outputs(5646) <= layer4_outputs(4042);
    outputs(5647) <= not(layer4_outputs(7038));
    outputs(5648) <= layer4_outputs(845);
    outputs(5649) <= layer4_outputs(3374);
    outputs(5650) <= not(layer4_outputs(7165));
    outputs(5651) <= (layer4_outputs(4778)) and not (layer4_outputs(1460));
    outputs(5652) <= layer4_outputs(2776);
    outputs(5653) <= not(layer4_outputs(736));
    outputs(5654) <= not(layer4_outputs(3381));
    outputs(5655) <= (layer4_outputs(4444)) and (layer4_outputs(6394));
    outputs(5656) <= layer4_outputs(5548);
    outputs(5657) <= not(layer4_outputs(2611));
    outputs(5658) <= layer4_outputs(6263);
    outputs(5659) <= not(layer4_outputs(774)) or (layer4_outputs(4805));
    outputs(5660) <= not(layer4_outputs(5771));
    outputs(5661) <= not(layer4_outputs(2483));
    outputs(5662) <= layer4_outputs(4600);
    outputs(5663) <= layer4_outputs(2407);
    outputs(5664) <= not(layer4_outputs(3106));
    outputs(5665) <= (layer4_outputs(174)) and not (layer4_outputs(893));
    outputs(5666) <= layer4_outputs(2913);
    outputs(5667) <= layer4_outputs(1095);
    outputs(5668) <= (layer4_outputs(4451)) xor (layer4_outputs(5059));
    outputs(5669) <= not((layer4_outputs(330)) or (layer4_outputs(994)));
    outputs(5670) <= not(layer4_outputs(804));
    outputs(5671) <= layer4_outputs(2564);
    outputs(5672) <= not((layer4_outputs(5127)) xor (layer4_outputs(2758)));
    outputs(5673) <= not(layer4_outputs(5508));
    outputs(5674) <= layer4_outputs(1415);
    outputs(5675) <= (layer4_outputs(4016)) and not (layer4_outputs(6135));
    outputs(5676) <= (layer4_outputs(6729)) and not (layer4_outputs(4034));
    outputs(5677) <= not(layer4_outputs(2831));
    outputs(5678) <= not(layer4_outputs(5270));
    outputs(5679) <= layer4_outputs(896);
    outputs(5680) <= not(layer4_outputs(4998));
    outputs(5681) <= (layer4_outputs(3615)) and (layer4_outputs(6064));
    outputs(5682) <= layer4_outputs(7574);
    outputs(5683) <= layer4_outputs(7018);
    outputs(5684) <= layer4_outputs(4713);
    outputs(5685) <= not(layer4_outputs(7518));
    outputs(5686) <= not((layer4_outputs(2893)) or (layer4_outputs(3480)));
    outputs(5687) <= not(layer4_outputs(3588));
    outputs(5688) <= (layer4_outputs(4610)) xor (layer4_outputs(3091));
    outputs(5689) <= layer4_outputs(5523);
    outputs(5690) <= layer4_outputs(6053);
    outputs(5691) <= not((layer4_outputs(1744)) xor (layer4_outputs(7453)));
    outputs(5692) <= not(layer4_outputs(5817));
    outputs(5693) <= layer4_outputs(4236);
    outputs(5694) <= layer4_outputs(6884);
    outputs(5695) <= layer4_outputs(961);
    outputs(5696) <= not(layer4_outputs(6167));
    outputs(5697) <= not(layer4_outputs(7375));
    outputs(5698) <= not(layer4_outputs(3346)) or (layer4_outputs(4357));
    outputs(5699) <= not(layer4_outputs(3971));
    outputs(5700) <= not(layer4_outputs(6003));
    outputs(5701) <= (layer4_outputs(6948)) and (layer4_outputs(6080));
    outputs(5702) <= (layer4_outputs(4020)) or (layer4_outputs(4509));
    outputs(5703) <= layer4_outputs(1893);
    outputs(5704) <= not((layer4_outputs(7083)) xor (layer4_outputs(6565)));
    outputs(5705) <= (layer4_outputs(6671)) and not (layer4_outputs(7163));
    outputs(5706) <= not((layer4_outputs(5467)) xor (layer4_outputs(2719)));
    outputs(5707) <= not(layer4_outputs(6882));
    outputs(5708) <= not(layer4_outputs(2142));
    outputs(5709) <= layer4_outputs(7602);
    outputs(5710) <= layer4_outputs(665);
    outputs(5711) <= not(layer4_outputs(4791));
    outputs(5712) <= (layer4_outputs(1231)) and not (layer4_outputs(4226));
    outputs(5713) <= not(layer4_outputs(936));
    outputs(5714) <= layer4_outputs(3979);
    outputs(5715) <= layer4_outputs(3907);
    outputs(5716) <= not(layer4_outputs(1461));
    outputs(5717) <= not((layer4_outputs(217)) xor (layer4_outputs(3497)));
    outputs(5718) <= (layer4_outputs(7057)) and not (layer4_outputs(6114));
    outputs(5719) <= layer4_outputs(5021);
    outputs(5720) <= (layer4_outputs(2920)) and (layer4_outputs(5945));
    outputs(5721) <= not(layer4_outputs(6324));
    outputs(5722) <= not((layer4_outputs(5587)) xor (layer4_outputs(745)));
    outputs(5723) <= not(layer4_outputs(4923));
    outputs(5724) <= not((layer4_outputs(3456)) or (layer4_outputs(1499)));
    outputs(5725) <= (layer4_outputs(4271)) and (layer4_outputs(833));
    outputs(5726) <= (layer4_outputs(2075)) and not (layer4_outputs(5727));
    outputs(5727) <= not(layer4_outputs(4961)) or (layer4_outputs(78));
    outputs(5728) <= not(layer4_outputs(7518)) or (layer4_outputs(6422));
    outputs(5729) <= layer4_outputs(5216);
    outputs(5730) <= layer4_outputs(7023);
    outputs(5731) <= not(layer4_outputs(7331));
    outputs(5732) <= (layer4_outputs(1343)) and (layer4_outputs(2311));
    outputs(5733) <= layer4_outputs(3111);
    outputs(5734) <= (layer4_outputs(7051)) and not (layer4_outputs(1171));
    outputs(5735) <= not(layer4_outputs(3802));
    outputs(5736) <= layer4_outputs(1388);
    outputs(5737) <= layer4_outputs(2081);
    outputs(5738) <= not((layer4_outputs(3015)) or (layer4_outputs(5413)));
    outputs(5739) <= (layer4_outputs(4209)) and (layer4_outputs(7559));
    outputs(5740) <= (layer4_outputs(3423)) and not (layer4_outputs(5880));
    outputs(5741) <= not(layer4_outputs(7439));
    outputs(5742) <= (layer4_outputs(7217)) and not (layer4_outputs(7537));
    outputs(5743) <= layer4_outputs(2701);
    outputs(5744) <= not(layer4_outputs(1031));
    outputs(5745) <= (layer4_outputs(5956)) and (layer4_outputs(5565));
    outputs(5746) <= not(layer4_outputs(4806));
    outputs(5747) <= (layer4_outputs(5453)) xor (layer4_outputs(142));
    outputs(5748) <= not(layer4_outputs(3064));
    outputs(5749) <= not(layer4_outputs(4165));
    outputs(5750) <= layer4_outputs(5220);
    outputs(5751) <= not((layer4_outputs(4885)) or (layer4_outputs(4463)));
    outputs(5752) <= layer4_outputs(7324);
    outputs(5753) <= not((layer4_outputs(3300)) or (layer4_outputs(5793)));
    outputs(5754) <= not((layer4_outputs(3762)) or (layer4_outputs(2152)));
    outputs(5755) <= (layer4_outputs(219)) and (layer4_outputs(2156));
    outputs(5756) <= layer4_outputs(7511);
    outputs(5757) <= not(layer4_outputs(4304));
    outputs(5758) <= not((layer4_outputs(1123)) xor (layer4_outputs(4199)));
    outputs(5759) <= layer4_outputs(1562);
    outputs(5760) <= not((layer4_outputs(5209)) or (layer4_outputs(3322)));
    outputs(5761) <= not(layer4_outputs(1739));
    outputs(5762) <= not(layer4_outputs(2934));
    outputs(5763) <= not(layer4_outputs(4435));
    outputs(5764) <= (layer4_outputs(7448)) and not (layer4_outputs(6432));
    outputs(5765) <= not(layer4_outputs(6497));
    outputs(5766) <= not((layer4_outputs(2262)) or (layer4_outputs(1892)));
    outputs(5767) <= not(layer4_outputs(2277));
    outputs(5768) <= (layer4_outputs(4626)) and (layer4_outputs(5205));
    outputs(5769) <= not((layer4_outputs(6227)) xor (layer4_outputs(5168)));
    outputs(5770) <= layer4_outputs(7164);
    outputs(5771) <= layer4_outputs(2883);
    outputs(5772) <= (layer4_outputs(4190)) and not (layer4_outputs(7224));
    outputs(5773) <= not(layer4_outputs(5359));
    outputs(5774) <= not(layer4_outputs(3104));
    outputs(5775) <= not((layer4_outputs(2028)) or (layer4_outputs(7459)));
    outputs(5776) <= (layer4_outputs(4363)) and not (layer4_outputs(1382));
    outputs(5777) <= not(layer4_outputs(1500));
    outputs(5778) <= layer4_outputs(6393);
    outputs(5779) <= (layer4_outputs(891)) or (layer4_outputs(25));
    outputs(5780) <= layer4_outputs(1790);
    outputs(5781) <= not(layer4_outputs(5925));
    outputs(5782) <= layer4_outputs(4895);
    outputs(5783) <= (layer4_outputs(1396)) and not (layer4_outputs(7286));
    outputs(5784) <= not((layer4_outputs(7289)) xor (layer4_outputs(4582)));
    outputs(5785) <= not(layer4_outputs(6258));
    outputs(5786) <= layer4_outputs(5207);
    outputs(5787) <= not((layer4_outputs(411)) and (layer4_outputs(4673)));
    outputs(5788) <= (layer4_outputs(12)) xor (layer4_outputs(2921));
    outputs(5789) <= (layer4_outputs(394)) and (layer4_outputs(3800));
    outputs(5790) <= layer4_outputs(4661);
    outputs(5791) <= layer4_outputs(6091);
    outputs(5792) <= (layer4_outputs(3367)) and not (layer4_outputs(3115));
    outputs(5793) <= not(layer4_outputs(6205));
    outputs(5794) <= (layer4_outputs(2830)) and not (layer4_outputs(5865));
    outputs(5795) <= (layer4_outputs(5235)) and not (layer4_outputs(3851));
    outputs(5796) <= not((layer4_outputs(1034)) xor (layer4_outputs(3258)));
    outputs(5797) <= layer4_outputs(768);
    outputs(5798) <= (layer4_outputs(7090)) xor (layer4_outputs(1771));
    outputs(5799) <= not(layer4_outputs(1494));
    outputs(5800) <= not(layer4_outputs(612));
    outputs(5801) <= not(layer4_outputs(5208));
    outputs(5802) <= not(layer4_outputs(3098));
    outputs(5803) <= not(layer4_outputs(6219));
    outputs(5804) <= layer4_outputs(5837);
    outputs(5805) <= layer4_outputs(6809);
    outputs(5806) <= not(layer4_outputs(2224));
    outputs(5807) <= not((layer4_outputs(6912)) xor (layer4_outputs(1092)));
    outputs(5808) <= not((layer4_outputs(1934)) xor (layer4_outputs(4322)));
    outputs(5809) <= layer4_outputs(37);
    outputs(5810) <= not(layer4_outputs(6864));
    outputs(5811) <= layer4_outputs(1474);
    outputs(5812) <= layer4_outputs(4594);
    outputs(5813) <= (layer4_outputs(6737)) and (layer4_outputs(3399));
    outputs(5814) <= layer4_outputs(2986);
    outputs(5815) <= (layer4_outputs(7644)) and not (layer4_outputs(3018));
    outputs(5816) <= not(layer4_outputs(2378));
    outputs(5817) <= (layer4_outputs(1856)) and not (layer4_outputs(2765));
    outputs(5818) <= (layer4_outputs(654)) xor (layer4_outputs(3418));
    outputs(5819) <= layer4_outputs(6609);
    outputs(5820) <= layer4_outputs(7484);
    outputs(5821) <= layer4_outputs(5803);
    outputs(5822) <= (layer4_outputs(1249)) and (layer4_outputs(1600));
    outputs(5823) <= not(layer4_outputs(1048));
    outputs(5824) <= (layer4_outputs(1996)) and not (layer4_outputs(1315));
    outputs(5825) <= not(layer4_outputs(2910));
    outputs(5826) <= layer4_outputs(7065);
    outputs(5827) <= layer4_outputs(6419);
    outputs(5828) <= layer4_outputs(4944);
    outputs(5829) <= not(layer4_outputs(6384));
    outputs(5830) <= not(layer4_outputs(156));
    outputs(5831) <= not(layer4_outputs(2810));
    outputs(5832) <= not(layer4_outputs(1311));
    outputs(5833) <= (layer4_outputs(6192)) or (layer4_outputs(2920));
    outputs(5834) <= not(layer4_outputs(4217));
    outputs(5835) <= not(layer4_outputs(1598));
    outputs(5836) <= layer4_outputs(7624);
    outputs(5837) <= not(layer4_outputs(964));
    outputs(5838) <= (layer4_outputs(4558)) and not (layer4_outputs(5561));
    outputs(5839) <= (layer4_outputs(2632)) xor (layer4_outputs(3003));
    outputs(5840) <= layer4_outputs(7170);
    outputs(5841) <= layer4_outputs(5097);
    outputs(5842) <= (layer4_outputs(7090)) and not (layer4_outputs(923));
    outputs(5843) <= (layer4_outputs(5321)) and not (layer4_outputs(2841));
    outputs(5844) <= not(layer4_outputs(2887));
    outputs(5845) <= not(layer4_outputs(3678));
    outputs(5846) <= (layer4_outputs(215)) xor (layer4_outputs(4666));
    outputs(5847) <= layer4_outputs(454);
    outputs(5848) <= (layer4_outputs(7039)) and (layer4_outputs(1459));
    outputs(5849) <= layer4_outputs(4946);
    outputs(5850) <= layer4_outputs(372);
    outputs(5851) <= layer4_outputs(2787);
    outputs(5852) <= layer4_outputs(6021);
    outputs(5853) <= not(layer4_outputs(4102)) or (layer4_outputs(6359));
    outputs(5854) <= layer4_outputs(1268);
    outputs(5855) <= not((layer4_outputs(5373)) or (layer4_outputs(4666)));
    outputs(5856) <= (layer4_outputs(4015)) xor (layer4_outputs(4185));
    outputs(5857) <= layer4_outputs(7102);
    outputs(5858) <= (layer4_outputs(6040)) and (layer4_outputs(1377));
    outputs(5859) <= not(layer4_outputs(4910));
    outputs(5860) <= layer4_outputs(659);
    outputs(5861) <= not(layer4_outputs(5197));
    outputs(5862) <= layer4_outputs(499);
    outputs(5863) <= layer4_outputs(5581);
    outputs(5864) <= layer4_outputs(5976);
    outputs(5865) <= layer4_outputs(4844);
    outputs(5866) <= not((layer4_outputs(3493)) or (layer4_outputs(4011)));
    outputs(5867) <= (layer4_outputs(1173)) and not (layer4_outputs(4232));
    outputs(5868) <= layer4_outputs(3400);
    outputs(5869) <= layer4_outputs(6883);
    outputs(5870) <= not(layer4_outputs(7033));
    outputs(5871) <= not((layer4_outputs(634)) xor (layer4_outputs(7403)));
    outputs(5872) <= (layer4_outputs(1179)) xor (layer4_outputs(161));
    outputs(5873) <= (layer4_outputs(6981)) and (layer4_outputs(720));
    outputs(5874) <= not(layer4_outputs(4205));
    outputs(5875) <= (layer4_outputs(4465)) and not (layer4_outputs(5539));
    outputs(5876) <= layer4_outputs(4767);
    outputs(5877) <= layer4_outputs(3993);
    outputs(5878) <= not((layer4_outputs(6209)) xor (layer4_outputs(3052)));
    outputs(5879) <= layer4_outputs(4519);
    outputs(5880) <= not(layer4_outputs(5362));
    outputs(5881) <= layer4_outputs(465);
    outputs(5882) <= (layer4_outputs(2877)) and (layer4_outputs(2484));
    outputs(5883) <= layer4_outputs(1937);
    outputs(5884) <= not((layer4_outputs(58)) or (layer4_outputs(7579)));
    outputs(5885) <= layer4_outputs(7244);
    outputs(5886) <= not(layer4_outputs(6897));
    outputs(5887) <= not(layer4_outputs(5811));
    outputs(5888) <= layer4_outputs(7641);
    outputs(5889) <= (layer4_outputs(5343)) and (layer4_outputs(1486));
    outputs(5890) <= not(layer4_outputs(3496));
    outputs(5891) <= (layer4_outputs(1018)) and (layer4_outputs(5839));
    outputs(5892) <= not((layer4_outputs(378)) xor (layer4_outputs(5903)));
    outputs(5893) <= (layer4_outputs(4301)) and (layer4_outputs(5145));
    outputs(5894) <= layer4_outputs(6295);
    outputs(5895) <= not(layer4_outputs(2224));
    outputs(5896) <= not(layer4_outputs(7443)) or (layer4_outputs(5273));
    outputs(5897) <= (layer4_outputs(6149)) xor (layer4_outputs(5804));
    outputs(5898) <= (layer4_outputs(2596)) and not (layer4_outputs(4975));
    outputs(5899) <= not(layer4_outputs(4272));
    outputs(5900) <= (layer4_outputs(4663)) xor (layer4_outputs(6306));
    outputs(5901) <= not(layer4_outputs(6130));
    outputs(5902) <= layer4_outputs(1899);
    outputs(5903) <= layer4_outputs(5243);
    outputs(5904) <= layer4_outputs(2517);
    outputs(5905) <= not(layer4_outputs(722)) or (layer4_outputs(1313));
    outputs(5906) <= layer4_outputs(6703);
    outputs(5907) <= (layer4_outputs(807)) and not (layer4_outputs(6587));
    outputs(5908) <= not(layer4_outputs(2709));
    outputs(5909) <= not(layer4_outputs(4786));
    outputs(5910) <= layer4_outputs(828);
    outputs(5911) <= (layer4_outputs(3399)) xor (layer4_outputs(565));
    outputs(5912) <= not((layer4_outputs(5890)) or (layer4_outputs(5025)));
    outputs(5913) <= not((layer4_outputs(1662)) xor (layer4_outputs(705)));
    outputs(5914) <= not(layer4_outputs(5635));
    outputs(5915) <= layer4_outputs(1110);
    outputs(5916) <= (layer4_outputs(352)) and not (layer4_outputs(4831));
    outputs(5917) <= layer4_outputs(5863);
    outputs(5918) <= not(layer4_outputs(1355));
    outputs(5919) <= not(layer4_outputs(6631));
    outputs(5920) <= not(layer4_outputs(6984));
    outputs(5921) <= (layer4_outputs(5439)) and (layer4_outputs(1051));
    outputs(5922) <= (layer4_outputs(4974)) and (layer4_outputs(2168));
    outputs(5923) <= layer4_outputs(4706);
    outputs(5924) <= layer4_outputs(656);
    outputs(5925) <= not(layer4_outputs(4494));
    outputs(5926) <= (layer4_outputs(6941)) and not (layer4_outputs(4934));
    outputs(5927) <= not((layer4_outputs(3740)) xor (layer4_outputs(2555)));
    outputs(5928) <= layer4_outputs(5815);
    outputs(5929) <= layer4_outputs(3748);
    outputs(5930) <= layer4_outputs(3801);
    outputs(5931) <= layer4_outputs(10);
    outputs(5932) <= not(layer4_outputs(3187));
    outputs(5933) <= not(layer4_outputs(6099));
    outputs(5934) <= layer4_outputs(5105);
    outputs(5935) <= not(layer4_outputs(1631));
    outputs(5936) <= layer4_outputs(2266);
    outputs(5937) <= not(layer4_outputs(4904));
    outputs(5938) <= (layer4_outputs(920)) and (layer4_outputs(1629));
    outputs(5939) <= (layer4_outputs(7386)) and not (layer4_outputs(1148));
    outputs(5940) <= layer4_outputs(2548);
    outputs(5941) <= layer4_outputs(3841);
    outputs(5942) <= not((layer4_outputs(5534)) and (layer4_outputs(2960)));
    outputs(5943) <= not(layer4_outputs(1008));
    outputs(5944) <= not(layer4_outputs(1271)) or (layer4_outputs(5327));
    outputs(5945) <= not(layer4_outputs(840));
    outputs(5946) <= not(layer4_outputs(2213));
    outputs(5947) <= not(layer4_outputs(5122));
    outputs(5948) <= not(layer4_outputs(3187)) or (layer4_outputs(5016));
    outputs(5949) <= not((layer4_outputs(1570)) xor (layer4_outputs(59)));
    outputs(5950) <= not(layer4_outputs(5174));
    outputs(5951) <= not(layer4_outputs(5644));
    outputs(5952) <= layer4_outputs(4154);
    outputs(5953) <= not(layer4_outputs(3944));
    outputs(5954) <= not((layer4_outputs(5444)) xor (layer4_outputs(447)));
    outputs(5955) <= not(layer4_outputs(2453));
    outputs(5956) <= (layer4_outputs(4433)) and (layer4_outputs(5565));
    outputs(5957) <= layer4_outputs(57);
    outputs(5958) <= not(layer4_outputs(6043));
    outputs(5959) <= not(layer4_outputs(6826));
    outputs(5960) <= not(layer4_outputs(211));
    outputs(5961) <= not(layer4_outputs(6004)) or (layer4_outputs(2051));
    outputs(5962) <= not(layer4_outputs(4329));
    outputs(5963) <= layer4_outputs(6654);
    outputs(5964) <= (layer4_outputs(6778)) xor (layer4_outputs(7108));
    outputs(5965) <= layer4_outputs(5769);
    outputs(5966) <= layer4_outputs(4509);
    outputs(5967) <= layer4_outputs(1413);
    outputs(5968) <= not(layer4_outputs(6556));
    outputs(5969) <= not(layer4_outputs(6246));
    outputs(5970) <= layer4_outputs(834);
    outputs(5971) <= layer4_outputs(1848);
    outputs(5972) <= not(layer4_outputs(1690));
    outputs(5973) <= layer4_outputs(1526);
    outputs(5974) <= not(layer4_outputs(755));
    outputs(5975) <= not(layer4_outputs(5381));
    outputs(5976) <= (layer4_outputs(1063)) and not (layer4_outputs(4503));
    outputs(5977) <= (layer4_outputs(3934)) or (layer4_outputs(4545));
    outputs(5978) <= layer4_outputs(1994);
    outputs(5979) <= layer4_outputs(694);
    outputs(5980) <= not(layer4_outputs(3596));
    outputs(5981) <= layer4_outputs(7460);
    outputs(5982) <= (layer4_outputs(809)) xor (layer4_outputs(1523));
    outputs(5983) <= (layer4_outputs(4812)) and (layer4_outputs(7339));
    outputs(5984) <= layer4_outputs(7187);
    outputs(5985) <= layer4_outputs(5137);
    outputs(5986) <= not(layer4_outputs(5898));
    outputs(5987) <= layer4_outputs(3963);
    outputs(5988) <= not(layer4_outputs(934));
    outputs(5989) <= (layer4_outputs(6982)) and not (layer4_outputs(531));
    outputs(5990) <= layer4_outputs(7569);
    outputs(5991) <= layer4_outputs(401);
    outputs(5992) <= not(layer4_outputs(4881));
    outputs(5993) <= layer4_outputs(4953);
    outputs(5994) <= not(layer4_outputs(4395));
    outputs(5995) <= (layer4_outputs(3495)) and not (layer4_outputs(2981));
    outputs(5996) <= not(layer4_outputs(4588));
    outputs(5997) <= not(layer4_outputs(2532));
    outputs(5998) <= not(layer4_outputs(4665));
    outputs(5999) <= layer4_outputs(7388);
    outputs(6000) <= not(layer4_outputs(780)) or (layer4_outputs(2907));
    outputs(6001) <= not((layer4_outputs(5077)) xor (layer4_outputs(7229)));
    outputs(6002) <= layer4_outputs(2248);
    outputs(6003) <= layer4_outputs(7523);
    outputs(6004) <= layer4_outputs(6548);
    outputs(6005) <= layer4_outputs(5089);
    outputs(6006) <= layer4_outputs(5327);
    outputs(6007) <= not(layer4_outputs(92));
    outputs(6008) <= not(layer4_outputs(2996));
    outputs(6009) <= not(layer4_outputs(1010));
    outputs(6010) <= not((layer4_outputs(5849)) xor (layer4_outputs(4061)));
    outputs(6011) <= layer4_outputs(1089);
    outputs(6012) <= not(layer4_outputs(804));
    outputs(6013) <= (layer4_outputs(1885)) and not (layer4_outputs(4876));
    outputs(6014) <= layer4_outputs(418);
    outputs(6015) <= (layer4_outputs(625)) and (layer4_outputs(1544));
    outputs(6016) <= layer4_outputs(3366);
    outputs(6017) <= not(layer4_outputs(3098)) or (layer4_outputs(5692));
    outputs(6018) <= not(layer4_outputs(5150));
    outputs(6019) <= not(layer4_outputs(2209));
    outputs(6020) <= layer4_outputs(285);
    outputs(6021) <= layer4_outputs(5483);
    outputs(6022) <= layer4_outputs(2744);
    outputs(6023) <= layer4_outputs(4025);
    outputs(6024) <= layer4_outputs(2344);
    outputs(6025) <= not(layer4_outputs(5161)) or (layer4_outputs(6367));
    outputs(6026) <= layer4_outputs(1065);
    outputs(6027) <= layer4_outputs(5440);
    outputs(6028) <= layer4_outputs(1812);
    outputs(6029) <= not((layer4_outputs(1573)) xor (layer4_outputs(1837)));
    outputs(6030) <= not(layer4_outputs(5721));
    outputs(6031) <= (layer4_outputs(7063)) xor (layer4_outputs(7391));
    outputs(6032) <= layer4_outputs(1838);
    outputs(6033) <= not(layer4_outputs(4441)) or (layer4_outputs(6138));
    outputs(6034) <= layer4_outputs(3028);
    outputs(6035) <= not(layer4_outputs(5672));
    outputs(6036) <= layer4_outputs(548);
    outputs(6037) <= (layer4_outputs(5267)) and not (layer4_outputs(6362));
    outputs(6038) <= not(layer4_outputs(4071));
    outputs(6039) <= (layer4_outputs(4676)) and (layer4_outputs(6204));
    outputs(6040) <= layer4_outputs(1346);
    outputs(6041) <= not(layer4_outputs(1177));
    outputs(6042) <= layer4_outputs(1308);
    outputs(6043) <= layer4_outputs(5087);
    outputs(6044) <= not(layer4_outputs(1226));
    outputs(6045) <= layer4_outputs(2484);
    outputs(6046) <= not((layer4_outputs(2885)) and (layer4_outputs(2779)));
    outputs(6047) <= (layer4_outputs(5046)) and not (layer4_outputs(5878));
    outputs(6048) <= not(layer4_outputs(3664));
    outputs(6049) <= not((layer4_outputs(450)) xor (layer4_outputs(1712)));
    outputs(6050) <= layer4_outputs(5469);
    outputs(6051) <= not(layer4_outputs(6532));
    outputs(6052) <= (layer4_outputs(1851)) xor (layer4_outputs(4464));
    outputs(6053) <= (layer4_outputs(1417)) and not (layer4_outputs(7123));
    outputs(6054) <= layer4_outputs(2852);
    outputs(6055) <= (layer4_outputs(5091)) or (layer4_outputs(7175));
    outputs(6056) <= not(layer4_outputs(6063));
    outputs(6057) <= layer4_outputs(1127);
    outputs(6058) <= not(layer4_outputs(799));
    outputs(6059) <= not((layer4_outputs(781)) xor (layer4_outputs(6614)));
    outputs(6060) <= not((layer4_outputs(2915)) xor (layer4_outputs(5509)));
    outputs(6061) <= layer4_outputs(3206);
    outputs(6062) <= layer4_outputs(64);
    outputs(6063) <= layer4_outputs(5131);
    outputs(6064) <= layer4_outputs(5309);
    outputs(6065) <= not(layer4_outputs(2708));
    outputs(6066) <= layer4_outputs(6021);
    outputs(6067) <= (layer4_outputs(4667)) and not (layer4_outputs(2949));
    outputs(6068) <= layer4_outputs(7608);
    outputs(6069) <= layer4_outputs(6467);
    outputs(6070) <= not(layer4_outputs(6336));
    outputs(6071) <= not((layer4_outputs(837)) xor (layer4_outputs(7636)));
    outputs(6072) <= layer4_outputs(4307);
    outputs(6073) <= not((layer4_outputs(1276)) xor (layer4_outputs(1788)));
    outputs(6074) <= (layer4_outputs(5235)) xor (layer4_outputs(501));
    outputs(6075) <= (layer4_outputs(2529)) and (layer4_outputs(2612));
    outputs(6076) <= layer4_outputs(151);
    outputs(6077) <= (layer4_outputs(458)) and (layer4_outputs(7483));
    outputs(6078) <= not(layer4_outputs(107)) or (layer4_outputs(3914));
    outputs(6079) <= layer4_outputs(5755);
    outputs(6080) <= not(layer4_outputs(4642));
    outputs(6081) <= not(layer4_outputs(2060));
    outputs(6082) <= not(layer4_outputs(4482));
    outputs(6083) <= not(layer4_outputs(3193));
    outputs(6084) <= not(layer4_outputs(7154));
    outputs(6085) <= layer4_outputs(6505);
    outputs(6086) <= not((layer4_outputs(2583)) or (layer4_outputs(4006)));
    outputs(6087) <= (layer4_outputs(6929)) and (layer4_outputs(3741));
    outputs(6088) <= layer4_outputs(6447);
    outputs(6089) <= (layer4_outputs(743)) and (layer4_outputs(4248));
    outputs(6090) <= not((layer4_outputs(4764)) or (layer4_outputs(4807)));
    outputs(6091) <= (layer4_outputs(4052)) and not (layer4_outputs(4768));
    outputs(6092) <= not(layer4_outputs(497));
    outputs(6093) <= not(layer4_outputs(3744));
    outputs(6094) <= (layer4_outputs(518)) or (layer4_outputs(5063));
    outputs(6095) <= layer4_outputs(665);
    outputs(6096) <= (layer4_outputs(1661)) and (layer4_outputs(6507));
    outputs(6097) <= layer4_outputs(4400);
    outputs(6098) <= layer4_outputs(3483);
    outputs(6099) <= layer4_outputs(6660);
    outputs(6100) <= layer4_outputs(5137);
    outputs(6101) <= layer4_outputs(81);
    outputs(6102) <= not(layer4_outputs(3837));
    outputs(6103) <= layer4_outputs(4340);
    outputs(6104) <= (layer4_outputs(1175)) xor (layer4_outputs(5502));
    outputs(6105) <= layer4_outputs(4913);
    outputs(6106) <= layer4_outputs(5954);
    outputs(6107) <= layer4_outputs(3347);
    outputs(6108) <= not(layer4_outputs(863));
    outputs(6109) <= not((layer4_outputs(6216)) and (layer4_outputs(2064)));
    outputs(6110) <= not((layer4_outputs(2504)) or (layer4_outputs(7211)));
    outputs(6111) <= not(layer4_outputs(6623));
    outputs(6112) <= layer4_outputs(5368);
    outputs(6113) <= not(layer4_outputs(365));
    outputs(6114) <= not((layer4_outputs(7270)) xor (layer4_outputs(6530)));
    outputs(6115) <= not(layer4_outputs(4));
    outputs(6116) <= not(layer4_outputs(5401));
    outputs(6117) <= layer4_outputs(2449);
    outputs(6118) <= layer4_outputs(1385);
    outputs(6119) <= not((layer4_outputs(7483)) xor (layer4_outputs(7418)));
    outputs(6120) <= not(layer4_outputs(857));
    outputs(6121) <= not((layer4_outputs(842)) xor (layer4_outputs(851)));
    outputs(6122) <= not(layer4_outputs(5620));
    outputs(6123) <= not(layer4_outputs(4515));
    outputs(6124) <= layer4_outputs(4488);
    outputs(6125) <= not(layer4_outputs(4120));
    outputs(6126) <= not(layer4_outputs(4046)) or (layer4_outputs(2792));
    outputs(6127) <= layer4_outputs(7345);
    outputs(6128) <= layer4_outputs(2487);
    outputs(6129) <= not((layer4_outputs(5405)) or (layer4_outputs(2194)));
    outputs(6130) <= (layer4_outputs(3605)) and (layer4_outputs(1643));
    outputs(6131) <= not(layer4_outputs(6902));
    outputs(6132) <= not(layer4_outputs(6715));
    outputs(6133) <= layer4_outputs(159);
    outputs(6134) <= (layer4_outputs(5335)) xor (layer4_outputs(3956));
    outputs(6135) <= layer4_outputs(856);
    outputs(6136) <= layer4_outputs(5981);
    outputs(6137) <= not((layer4_outputs(3523)) xor (layer4_outputs(1222)));
    outputs(6138) <= layer4_outputs(3606);
    outputs(6139) <= (layer4_outputs(6824)) and (layer4_outputs(7543));
    outputs(6140) <= (layer4_outputs(1642)) xor (layer4_outputs(4415));
    outputs(6141) <= layer4_outputs(3080);
    outputs(6142) <= layer4_outputs(6898);
    outputs(6143) <= layer4_outputs(4623);
    outputs(6144) <= (layer4_outputs(5826)) and not (layer4_outputs(7436));
    outputs(6145) <= not((layer4_outputs(1987)) and (layer4_outputs(7230)));
    outputs(6146) <= layer4_outputs(5325);
    outputs(6147) <= (layer4_outputs(2145)) xor (layer4_outputs(617));
    outputs(6148) <= layer4_outputs(4012);
    outputs(6149) <= layer4_outputs(3240);
    outputs(6150) <= not(layer4_outputs(862));
    outputs(6151) <= (layer4_outputs(2794)) and (layer4_outputs(7142));
    outputs(6152) <= layer4_outputs(3527);
    outputs(6153) <= layer4_outputs(7396);
    outputs(6154) <= not(layer4_outputs(1314));
    outputs(6155) <= not(layer4_outputs(1066));
    outputs(6156) <= (layer4_outputs(7414)) xor (layer4_outputs(5324));
    outputs(6157) <= (layer4_outputs(2496)) and not (layer4_outputs(3317));
    outputs(6158) <= layer4_outputs(20);
    outputs(6159) <= layer4_outputs(6222);
    outputs(6160) <= (layer4_outputs(2045)) xor (layer4_outputs(6830));
    outputs(6161) <= (layer4_outputs(2307)) xor (layer4_outputs(47));
    outputs(6162) <= not((layer4_outputs(6731)) xor (layer4_outputs(2267)));
    outputs(6163) <= layer4_outputs(5178);
    outputs(6164) <= not(layer4_outputs(3829));
    outputs(6165) <= layer4_outputs(4941);
    outputs(6166) <= layer4_outputs(7389);
    outputs(6167) <= not(layer4_outputs(979));
    outputs(6168) <= layer4_outputs(880);
    outputs(6169) <= not(layer4_outputs(3667)) or (layer4_outputs(6586));
    outputs(6170) <= not((layer4_outputs(6706)) xor (layer4_outputs(4996)));
    outputs(6171) <= layer4_outputs(1137);
    outputs(6172) <= (layer4_outputs(2360)) xor (layer4_outputs(5910));
    outputs(6173) <= layer4_outputs(1791);
    outputs(6174) <= not(layer4_outputs(603));
    outputs(6175) <= not((layer4_outputs(1959)) xor (layer4_outputs(4667)));
    outputs(6176) <= not(layer4_outputs(4061));
    outputs(6177) <= layer4_outputs(3289);
    outputs(6178) <= not(layer4_outputs(3790));
    outputs(6179) <= (layer4_outputs(1001)) xor (layer4_outputs(3663));
    outputs(6180) <= not((layer4_outputs(1925)) xor (layer4_outputs(2252)));
    outputs(6181) <= (layer4_outputs(1635)) and (layer4_outputs(2357));
    outputs(6182) <= not(layer4_outputs(727));
    outputs(6183) <= not(layer4_outputs(6822));
    outputs(6184) <= layer4_outputs(5239);
    outputs(6185) <= not(layer4_outputs(7160));
    outputs(6186) <= not(layer4_outputs(4814));
    outputs(6187) <= not(layer4_outputs(7350)) or (layer4_outputs(2725));
    outputs(6188) <= not((layer4_outputs(5543)) xor (layer4_outputs(3315)));
    outputs(6189) <= (layer4_outputs(6338)) and (layer4_outputs(2661));
    outputs(6190) <= layer4_outputs(7380);
    outputs(6191) <= (layer4_outputs(6511)) xor (layer4_outputs(3005));
    outputs(6192) <= (layer4_outputs(4302)) xor (layer4_outputs(6779));
    outputs(6193) <= not(layer4_outputs(5094)) or (layer4_outputs(5027));
    outputs(6194) <= (layer4_outputs(3525)) and not (layer4_outputs(4848));
    outputs(6195) <= layer4_outputs(4542);
    outputs(6196) <= (layer4_outputs(4142)) xor (layer4_outputs(6571));
    outputs(6197) <= not(layer4_outputs(2056));
    outputs(6198) <= (layer4_outputs(5906)) and not (layer4_outputs(4680));
    outputs(6199) <= not((layer4_outputs(4715)) or (layer4_outputs(3286)));
    outputs(6200) <= (layer4_outputs(3263)) or (layer4_outputs(5668));
    outputs(6201) <= layer4_outputs(6255);
    outputs(6202) <= not(layer4_outputs(26));
    outputs(6203) <= not(layer4_outputs(4305)) or (layer4_outputs(3548));
    outputs(6204) <= (layer4_outputs(3880)) or (layer4_outputs(585));
    outputs(6205) <= (layer4_outputs(1202)) xor (layer4_outputs(6200));
    outputs(6206) <= layer4_outputs(4954);
    outputs(6207) <= not((layer4_outputs(4925)) and (layer4_outputs(1640)));
    outputs(6208) <= not((layer4_outputs(909)) or (layer4_outputs(4740)));
    outputs(6209) <= (layer4_outputs(3955)) xor (layer4_outputs(4717));
    outputs(6210) <= layer4_outputs(7563);
    outputs(6211) <= (layer4_outputs(2937)) and (layer4_outputs(2089));
    outputs(6212) <= not(layer4_outputs(2590));
    outputs(6213) <= not(layer4_outputs(3434));
    outputs(6214) <= not((layer4_outputs(7410)) xor (layer4_outputs(1556)));
    outputs(6215) <= not((layer4_outputs(631)) or (layer4_outputs(5379)));
    outputs(6216) <= (layer4_outputs(567)) or (layer4_outputs(7215));
    outputs(6217) <= not((layer4_outputs(3602)) xor (layer4_outputs(3432)));
    outputs(6218) <= (layer4_outputs(7354)) and (layer4_outputs(5222));
    outputs(6219) <= layer4_outputs(2330);
    outputs(6220) <= not((layer4_outputs(4675)) or (layer4_outputs(4365)));
    outputs(6221) <= not((layer4_outputs(5782)) or (layer4_outputs(2494)));
    outputs(6222) <= layer4_outputs(6351);
    outputs(6223) <= not(layer4_outputs(4581));
    outputs(6224) <= not((layer4_outputs(3731)) and (layer4_outputs(904)));
    outputs(6225) <= layer4_outputs(7007);
    outputs(6226) <= (layer4_outputs(5041)) xor (layer4_outputs(1237));
    outputs(6227) <= layer4_outputs(1837);
    outputs(6228) <= (layer4_outputs(6110)) xor (layer4_outputs(6333));
    outputs(6229) <= layer4_outputs(508);
    outputs(6230) <= not((layer4_outputs(4995)) xor (layer4_outputs(3740)));
    outputs(6231) <= layer4_outputs(4189);
    outputs(6232) <= layer4_outputs(2085);
    outputs(6233) <= not(layer4_outputs(6392));
    outputs(6234) <= layer4_outputs(4969);
    outputs(6235) <= not(layer4_outputs(3942));
    outputs(6236) <= layer4_outputs(1814);
    outputs(6237) <= not(layer4_outputs(2988));
    outputs(6238) <= layer4_outputs(1627);
    outputs(6239) <= layer4_outputs(2829);
    outputs(6240) <= not(layer4_outputs(3427)) or (layer4_outputs(1559));
    outputs(6241) <= layer4_outputs(5566);
    outputs(6242) <= not((layer4_outputs(4039)) xor (layer4_outputs(1785)));
    outputs(6243) <= (layer4_outputs(6532)) and not (layer4_outputs(2590));
    outputs(6244) <= (layer4_outputs(6538)) xor (layer4_outputs(2001));
    outputs(6245) <= not((layer4_outputs(1015)) xor (layer4_outputs(669)));
    outputs(6246) <= (layer4_outputs(1722)) and (layer4_outputs(810));
    outputs(6247) <= (layer4_outputs(4352)) and (layer4_outputs(5597));
    outputs(6248) <= layer4_outputs(1927);
    outputs(6249) <= (layer4_outputs(6010)) and not (layer4_outputs(2259));
    outputs(6250) <= not((layer4_outputs(6774)) or (layer4_outputs(4328)));
    outputs(6251) <= not((layer4_outputs(3166)) xor (layer4_outputs(2275)));
    outputs(6252) <= not(layer4_outputs(4299));
    outputs(6253) <= (layer4_outputs(1292)) and (layer4_outputs(3152));
    outputs(6254) <= layer4_outputs(3162);
    outputs(6255) <= not(layer4_outputs(1973));
    outputs(6256) <= not((layer4_outputs(441)) xor (layer4_outputs(2031)));
    outputs(6257) <= not((layer4_outputs(555)) xor (layer4_outputs(5648)));
    outputs(6258) <= not((layer4_outputs(3889)) and (layer4_outputs(3167)));
    outputs(6259) <= not(layer4_outputs(2939));
    outputs(6260) <= (layer4_outputs(2383)) xor (layer4_outputs(3473));
    outputs(6261) <= (layer4_outputs(7577)) and not (layer4_outputs(7));
    outputs(6262) <= layer4_outputs(5093);
    outputs(6263) <= layer4_outputs(3582);
    outputs(6264) <= (layer4_outputs(442)) or (layer4_outputs(6252));
    outputs(6265) <= not(layer4_outputs(1511));
    outputs(6266) <= (layer4_outputs(8)) xor (layer4_outputs(4250));
    outputs(6267) <= (layer4_outputs(4085)) and not (layer4_outputs(6282));
    outputs(6268) <= not((layer4_outputs(2371)) or (layer4_outputs(4657)));
    outputs(6269) <= (layer4_outputs(6574)) xor (layer4_outputs(6445));
    outputs(6270) <= layer4_outputs(5240);
    outputs(6271) <= (layer4_outputs(783)) and not (layer4_outputs(1656));
    outputs(6272) <= layer4_outputs(1933);
    outputs(6273) <= layer4_outputs(1262);
    outputs(6274) <= (layer4_outputs(5277)) xor (layer4_outputs(6969));
    outputs(6275) <= not(layer4_outputs(4045));
    outputs(6276) <= not((layer4_outputs(5074)) xor (layer4_outputs(6203)));
    outputs(6277) <= not(layer4_outputs(2789));
    outputs(6278) <= not((layer4_outputs(6193)) xor (layer4_outputs(2814)));
    outputs(6279) <= (layer4_outputs(3628)) or (layer4_outputs(7255));
    outputs(6280) <= (layer4_outputs(6312)) or (layer4_outputs(5533));
    outputs(6281) <= (layer4_outputs(5008)) xor (layer4_outputs(3002));
    outputs(6282) <= layer4_outputs(4672);
    outputs(6283) <= layer4_outputs(6487);
    outputs(6284) <= (layer4_outputs(5200)) and not (layer4_outputs(5547));
    outputs(6285) <= (layer4_outputs(1811)) and (layer4_outputs(1194));
    outputs(6286) <= not((layer4_outputs(6372)) xor (layer4_outputs(7082)));
    outputs(6287) <= not(layer4_outputs(2249));
    outputs(6288) <= layer4_outputs(4524);
    outputs(6289) <= not(layer4_outputs(4652));
    outputs(6290) <= not(layer4_outputs(7048)) or (layer4_outputs(7300));
    outputs(6291) <= layer4_outputs(7532);
    outputs(6292) <= not(layer4_outputs(2648)) or (layer4_outputs(495));
    outputs(6293) <= (layer4_outputs(1948)) xor (layer4_outputs(1776));
    outputs(6294) <= not(layer4_outputs(511));
    outputs(6295) <= not((layer4_outputs(3047)) or (layer4_outputs(5538)));
    outputs(6296) <= not((layer4_outputs(4885)) or (layer4_outputs(5128)));
    outputs(6297) <= not(layer4_outputs(2770)) or (layer4_outputs(736));
    outputs(6298) <= not(layer4_outputs(5417));
    outputs(6299) <= layer4_outputs(6410);
    outputs(6300) <= layer4_outputs(3004);
    outputs(6301) <= not(layer4_outputs(5483));
    outputs(6302) <= (layer4_outputs(929)) and not (layer4_outputs(4733));
    outputs(6303) <= (layer4_outputs(4380)) and not (layer4_outputs(6295));
    outputs(6304) <= (layer4_outputs(5202)) xor (layer4_outputs(3770));
    outputs(6305) <= (layer4_outputs(7480)) or (layer4_outputs(5292));
    outputs(6306) <= layer4_outputs(2752);
    outputs(6307) <= layer4_outputs(3994);
    outputs(6308) <= not(layer4_outputs(2544));
    outputs(6309) <= not(layer4_outputs(4638));
    outputs(6310) <= not((layer4_outputs(3069)) xor (layer4_outputs(2866)));
    outputs(6311) <= not(layer4_outputs(2539)) or (layer4_outputs(3217));
    outputs(6312) <= not((layer4_outputs(1486)) xor (layer4_outputs(1663)));
    outputs(6313) <= not(layer4_outputs(1306)) or (layer4_outputs(6510));
    outputs(6314) <= not(layer4_outputs(930)) or (layer4_outputs(339));
    outputs(6315) <= layer4_outputs(2895);
    outputs(6316) <= (layer4_outputs(2585)) or (layer4_outputs(2437));
    outputs(6317) <= not(layer4_outputs(6792));
    outputs(6318) <= not(layer4_outputs(6070));
    outputs(6319) <= (layer4_outputs(1745)) and not (layer4_outputs(413));
    outputs(6320) <= not(layer4_outputs(6833));
    outputs(6321) <= (layer4_outputs(1727)) xor (layer4_outputs(7001));
    outputs(6322) <= (layer4_outputs(4754)) xor (layer4_outputs(3776));
    outputs(6323) <= not(layer4_outputs(5675));
    outputs(6324) <= not(layer4_outputs(5788));
    outputs(6325) <= not(layer4_outputs(4803));
    outputs(6326) <= not(layer4_outputs(2635));
    outputs(6327) <= (layer4_outputs(343)) xor (layer4_outputs(6475));
    outputs(6328) <= not(layer4_outputs(7652));
    outputs(6329) <= (layer4_outputs(4918)) xor (layer4_outputs(4175));
    outputs(6330) <= not(layer4_outputs(3348));
    outputs(6331) <= (layer4_outputs(3977)) xor (layer4_outputs(6612));
    outputs(6332) <= (layer4_outputs(4946)) and not (layer4_outputs(2200));
    outputs(6333) <= not(layer4_outputs(5180));
    outputs(6334) <= not(layer4_outputs(1289));
    outputs(6335) <= not((layer4_outputs(1700)) xor (layer4_outputs(7547)));
    outputs(6336) <= not((layer4_outputs(1323)) xor (layer4_outputs(649)));
    outputs(6337) <= layer4_outputs(746);
    outputs(6338) <= not(layer4_outputs(5408)) or (layer4_outputs(622));
    outputs(6339) <= layer4_outputs(2639);
    outputs(6340) <= not(layer4_outputs(4653));
    outputs(6341) <= layer4_outputs(901);
    outputs(6342) <= layer4_outputs(4294);
    outputs(6343) <= layer4_outputs(3983);
    outputs(6344) <= (layer4_outputs(7259)) xor (layer4_outputs(2418));
    outputs(6345) <= (layer4_outputs(1355)) and (layer4_outputs(705));
    outputs(6346) <= not(layer4_outputs(6900));
    outputs(6347) <= not(layer4_outputs(4701)) or (layer4_outputs(36));
    outputs(6348) <= layer4_outputs(5470);
    outputs(6349) <= not(layer4_outputs(1931)) or (layer4_outputs(5282));
    outputs(6350) <= not((layer4_outputs(5103)) xor (layer4_outputs(76)));
    outputs(6351) <= layer4_outputs(3788);
    outputs(6352) <= not((layer4_outputs(4123)) xor (layer4_outputs(6909)));
    outputs(6353) <= not((layer4_outputs(6953)) xor (layer4_outputs(141)));
    outputs(6354) <= (layer4_outputs(2630)) and (layer4_outputs(1083));
    outputs(6355) <= not(layer4_outputs(7587));
    outputs(6356) <= not(layer4_outputs(3517));
    outputs(6357) <= not(layer4_outputs(4074));
    outputs(6358) <= (layer4_outputs(997)) xor (layer4_outputs(2475));
    outputs(6359) <= not(layer4_outputs(4744));
    outputs(6360) <= not((layer4_outputs(6097)) xor (layer4_outputs(2433)));
    outputs(6361) <= layer4_outputs(4670);
    outputs(6362) <= not(layer4_outputs(6892));
    outputs(6363) <= layer4_outputs(263);
    outputs(6364) <= layer4_outputs(654);
    outputs(6365) <= layer4_outputs(4902);
    outputs(6366) <= layer4_outputs(6655);
    outputs(6367) <= (layer4_outputs(963)) xor (layer4_outputs(301));
    outputs(6368) <= not(layer4_outputs(1359)) or (layer4_outputs(6708));
    outputs(6369) <= not(layer4_outputs(5799));
    outputs(6370) <= not(layer4_outputs(3919));
    outputs(6371) <= not((layer4_outputs(4923)) xor (layer4_outputs(6328)));
    outputs(6372) <= not(layer4_outputs(3491));
    outputs(6373) <= not(layer4_outputs(2668));
    outputs(6374) <= (layer4_outputs(4663)) xor (layer4_outputs(3428));
    outputs(6375) <= not(layer4_outputs(571));
    outputs(6376) <= layer4_outputs(3943);
    outputs(6377) <= not(layer4_outputs(2202));
    outputs(6378) <= not(layer4_outputs(3422));
    outputs(6379) <= layer4_outputs(6889);
    outputs(6380) <= (layer4_outputs(5804)) or (layer4_outputs(5798));
    outputs(6381) <= (layer4_outputs(218)) and not (layer4_outputs(1199));
    outputs(6382) <= (layer4_outputs(4028)) xor (layer4_outputs(3476));
    outputs(6383) <= not((layer4_outputs(5328)) xor (layer4_outputs(5431)));
    outputs(6384) <= not((layer4_outputs(3259)) or (layer4_outputs(2732)));
    outputs(6385) <= not(layer4_outputs(2806));
    outputs(6386) <= layer4_outputs(7147);
    outputs(6387) <= layer4_outputs(6716);
    outputs(6388) <= layer4_outputs(4453);
    outputs(6389) <= layer4_outputs(5038);
    outputs(6390) <= (layer4_outputs(1675)) xor (layer4_outputs(5065));
    outputs(6391) <= (layer4_outputs(3484)) xor (layer4_outputs(6966));
    outputs(6392) <= layer4_outputs(6874);
    outputs(6393) <= layer4_outputs(3438);
    outputs(6394) <= not((layer4_outputs(2970)) and (layer4_outputs(4292)));
    outputs(6395) <= not((layer4_outputs(4020)) xor (layer4_outputs(16)));
    outputs(6396) <= not(layer4_outputs(2303));
    outputs(6397) <= layer4_outputs(5492);
    outputs(6398) <= not(layer4_outputs(7489));
    outputs(6399) <= not(layer4_outputs(6303)) or (layer4_outputs(7600));
    outputs(6400) <= layer4_outputs(6910);
    outputs(6401) <= layer4_outputs(3409);
    outputs(6402) <= layer4_outputs(7088);
    outputs(6403) <= (layer4_outputs(7273)) or (layer4_outputs(5425));
    outputs(6404) <= not((layer4_outputs(471)) xor (layer4_outputs(1639)));
    outputs(6405) <= not((layer4_outputs(2462)) xor (layer4_outputs(2169)));
    outputs(6406) <= layer4_outputs(3276);
    outputs(6407) <= layer4_outputs(7520);
    outputs(6408) <= not(layer4_outputs(6941));
    outputs(6409) <= not(layer4_outputs(2803));
    outputs(6410) <= not((layer4_outputs(2919)) and (layer4_outputs(5889)));
    outputs(6411) <= not((layer4_outputs(1501)) xor (layer4_outputs(5149)));
    outputs(6412) <= not((layer4_outputs(4413)) xor (layer4_outputs(2723)));
    outputs(6413) <= not(layer4_outputs(5466));
    outputs(6414) <= not(layer4_outputs(3425));
    outputs(6415) <= (layer4_outputs(709)) and (layer4_outputs(2341));
    outputs(6416) <= not((layer4_outputs(2395)) xor (layer4_outputs(3030)));
    outputs(6417) <= layer4_outputs(7579);
    outputs(6418) <= (layer4_outputs(2073)) xor (layer4_outputs(4677));
    outputs(6419) <= layer4_outputs(6233);
    outputs(6420) <= not(layer4_outputs(3256));
    outputs(6421) <= not(layer4_outputs(5190));
    outputs(6422) <= layer4_outputs(6041);
    outputs(6423) <= (layer4_outputs(5292)) and (layer4_outputs(1104));
    outputs(6424) <= (layer4_outputs(1316)) xor (layer4_outputs(2125));
    outputs(6425) <= not(layer4_outputs(7175));
    outputs(6426) <= (layer4_outputs(1288)) and (layer4_outputs(2020));
    outputs(6427) <= not(layer4_outputs(3849));
    outputs(6428) <= not(layer4_outputs(1451));
    outputs(6429) <= not(layer4_outputs(365));
    outputs(6430) <= not(layer4_outputs(3799)) or (layer4_outputs(4810));
    outputs(6431) <= (layer4_outputs(6631)) xor (layer4_outputs(4937));
    outputs(6432) <= layer4_outputs(949);
    outputs(6433) <= not(layer4_outputs(6383));
    outputs(6434) <= layer4_outputs(764);
    outputs(6435) <= (layer4_outputs(1384)) xor (layer4_outputs(6685));
    outputs(6436) <= (layer4_outputs(992)) xor (layer4_outputs(4711));
    outputs(6437) <= layer4_outputs(3722);
    outputs(6438) <= (layer4_outputs(6649)) and not (layer4_outputs(2080));
    outputs(6439) <= not(layer4_outputs(6774));
    outputs(6440) <= layer4_outputs(1995);
    outputs(6441) <= (layer4_outputs(989)) xor (layer4_outputs(6583));
    outputs(6442) <= not((layer4_outputs(4475)) xor (layer4_outputs(5881)));
    outputs(6443) <= layer4_outputs(901);
    outputs(6444) <= layer4_outputs(5368);
    outputs(6445) <= not(layer4_outputs(6244));
    outputs(6446) <= not(layer4_outputs(3969));
    outputs(6447) <= (layer4_outputs(599)) xor (layer4_outputs(3877));
    outputs(6448) <= not((layer4_outputs(2503)) xor (layer4_outputs(2986)));
    outputs(6449) <= not((layer4_outputs(5386)) xor (layer4_outputs(2315)));
    outputs(6450) <= not(layer4_outputs(1205)) or (layer4_outputs(699));
    outputs(6451) <= not((layer4_outputs(5926)) and (layer4_outputs(5691)));
    outputs(6452) <= (layer4_outputs(5278)) xor (layer4_outputs(4038));
    outputs(6453) <= (layer4_outputs(1335)) and not (layer4_outputs(3223));
    outputs(6454) <= layer4_outputs(1045);
    outputs(6455) <= layer4_outputs(7422);
    outputs(6456) <= not(layer4_outputs(6181));
    outputs(6457) <= not(layer4_outputs(1245));
    outputs(6458) <= (layer4_outputs(1958)) and not (layer4_outputs(4250));
    outputs(6459) <= not(layer4_outputs(3301));
    outputs(6460) <= (layer4_outputs(2004)) and not (layer4_outputs(3001));
    outputs(6461) <= not(layer4_outputs(1218));
    outputs(6462) <= not(layer4_outputs(1575));
    outputs(6463) <= layer4_outputs(4707);
    outputs(6464) <= layer4_outputs(6704);
    outputs(6465) <= not((layer4_outputs(2418)) xor (layer4_outputs(2765)));
    outputs(6466) <= layer4_outputs(3426);
    outputs(6467) <= layer4_outputs(5925);
    outputs(6468) <= not(layer4_outputs(554));
    outputs(6469) <= (layer4_outputs(3014)) xor (layer4_outputs(5980));
    outputs(6470) <= layer4_outputs(6272);
    outputs(6471) <= not((layer4_outputs(2139)) xor (layer4_outputs(4636)));
    outputs(6472) <= (layer4_outputs(27)) xor (layer4_outputs(2922));
    outputs(6473) <= layer4_outputs(2515);
    outputs(6474) <= not(layer4_outputs(2602));
    outputs(6475) <= (layer4_outputs(3449)) xor (layer4_outputs(6114));
    outputs(6476) <= not((layer4_outputs(6018)) xor (layer4_outputs(1115)));
    outputs(6477) <= not((layer4_outputs(7562)) xor (layer4_outputs(6784)));
    outputs(6478) <= (layer4_outputs(546)) xor (layer4_outputs(455));
    outputs(6479) <= layer4_outputs(7405);
    outputs(6480) <= layer4_outputs(520);
    outputs(6481) <= not((layer4_outputs(6658)) xor (layer4_outputs(2714)));
    outputs(6482) <= layer4_outputs(985);
    outputs(6483) <= layer4_outputs(2764);
    outputs(6484) <= layer4_outputs(4462);
    outputs(6485) <= (layer4_outputs(753)) and not (layer4_outputs(6939));
    outputs(6486) <= not(layer4_outputs(3419));
    outputs(6487) <= (layer4_outputs(2800)) xor (layer4_outputs(1369));
    outputs(6488) <= (layer4_outputs(2104)) and not (layer4_outputs(4241));
    outputs(6489) <= not(layer4_outputs(470));
    outputs(6490) <= layer4_outputs(4508);
    outputs(6491) <= not(layer4_outputs(4427));
    outputs(6492) <= layer4_outputs(4671);
    outputs(6493) <= not(layer4_outputs(1554));
    outputs(6494) <= (layer4_outputs(6402)) xor (layer4_outputs(313));
    outputs(6495) <= layer4_outputs(2521);
    outputs(6496) <= not(layer4_outputs(3603));
    outputs(6497) <= not(layer4_outputs(2926));
    outputs(6498) <= not(layer4_outputs(2673));
    outputs(6499) <= not((layer4_outputs(340)) xor (layer4_outputs(4821)));
    outputs(6500) <= not(layer4_outputs(7513));
    outputs(6501) <= layer4_outputs(6976);
    outputs(6502) <= layer4_outputs(709);
    outputs(6503) <= layer4_outputs(2151);
    outputs(6504) <= layer4_outputs(6642);
    outputs(6505) <= not(layer4_outputs(3849));
    outputs(6506) <= layer4_outputs(6866);
    outputs(6507) <= (layer4_outputs(825)) and not (layer4_outputs(490));
    outputs(6508) <= (layer4_outputs(7227)) xor (layer4_outputs(5130));
    outputs(6509) <= (layer4_outputs(7607)) and not (layer4_outputs(6660));
    outputs(6510) <= not(layer4_outputs(250));
    outputs(6511) <= not((layer4_outputs(539)) and (layer4_outputs(7054)));
    outputs(6512) <= layer4_outputs(5610);
    outputs(6513) <= not(layer4_outputs(1026));
    outputs(6514) <= not(layer4_outputs(5666));
    outputs(6515) <= layer4_outputs(7317);
    outputs(6516) <= not(layer4_outputs(234));
    outputs(6517) <= (layer4_outputs(1535)) xor (layer4_outputs(6514));
    outputs(6518) <= not(layer4_outputs(3342));
    outputs(6519) <= layer4_outputs(3217);
    outputs(6520) <= layer4_outputs(6920);
    outputs(6521) <= not(layer4_outputs(3826));
    outputs(6522) <= not(layer4_outputs(6927));
    outputs(6523) <= not(layer4_outputs(6366));
    outputs(6524) <= not((layer4_outputs(4310)) xor (layer4_outputs(5875)));
    outputs(6525) <= not((layer4_outputs(304)) or (layer4_outputs(577)));
    outputs(6526) <= (layer4_outputs(4988)) xor (layer4_outputs(786));
    outputs(6527) <= not(layer4_outputs(4180));
    outputs(6528) <= layer4_outputs(6294);
    outputs(6529) <= not((layer4_outputs(7194)) xor (layer4_outputs(2720)));
    outputs(6530) <= (layer4_outputs(1042)) and not (layer4_outputs(5625));
    outputs(6531) <= not((layer4_outputs(4017)) xor (layer4_outputs(4580)));
    outputs(6532) <= layer4_outputs(764);
    outputs(6533) <= layer4_outputs(1194);
    outputs(6534) <= (layer4_outputs(5949)) xor (layer4_outputs(794));
    outputs(6535) <= (layer4_outputs(1152)) or (layer4_outputs(5818));
    outputs(6536) <= layer4_outputs(4843);
    outputs(6537) <= (layer4_outputs(4684)) and (layer4_outputs(4461));
    outputs(6538) <= not(layer4_outputs(6661));
    outputs(6539) <= not(layer4_outputs(193));
    outputs(6540) <= (layer4_outputs(7325)) and (layer4_outputs(186));
    outputs(6541) <= not((layer4_outputs(7319)) xor (layer4_outputs(1266)));
    outputs(6542) <= layer4_outputs(3943);
    outputs(6543) <= (layer4_outputs(2285)) or (layer4_outputs(5838));
    outputs(6544) <= layer4_outputs(3379);
    outputs(6545) <= (layer4_outputs(2583)) and (layer4_outputs(5308));
    outputs(6546) <= not(layer4_outputs(3383));
    outputs(6547) <= layer4_outputs(7577);
    outputs(6548) <= not(layer4_outputs(5382));
    outputs(6549) <= not(layer4_outputs(7586));
    outputs(6550) <= layer4_outputs(206);
    outputs(6551) <= (layer4_outputs(2219)) xor (layer4_outputs(1002));
    outputs(6552) <= not(layer4_outputs(2592));
    outputs(6553) <= not(layer4_outputs(3541));
    outputs(6554) <= (layer4_outputs(6166)) xor (layer4_outputs(1422));
    outputs(6555) <= not(layer4_outputs(1337));
    outputs(6556) <= not((layer4_outputs(3572)) xor (layer4_outputs(4196)));
    outputs(6557) <= not((layer4_outputs(3342)) xor (layer4_outputs(7008)));
    outputs(6558) <= (layer4_outputs(6010)) and not (layer4_outputs(3105));
    outputs(6559) <= not(layer4_outputs(4188));
    outputs(6560) <= layer4_outputs(320);
    outputs(6561) <= layer4_outputs(7634);
    outputs(6562) <= layer4_outputs(4561);
    outputs(6563) <= (layer4_outputs(3329)) xor (layer4_outputs(3604));
    outputs(6564) <= layer4_outputs(1836);
    outputs(6565) <= (layer4_outputs(6564)) xor (layer4_outputs(582));
    outputs(6566) <= (layer4_outputs(5374)) xor (layer4_outputs(3793));
    outputs(6567) <= (layer4_outputs(2658)) and not (layer4_outputs(3511));
    outputs(6568) <= layer4_outputs(4169);
    outputs(6569) <= layer4_outputs(462);
    outputs(6570) <= layer4_outputs(1044);
    outputs(6571) <= (layer4_outputs(2342)) xor (layer4_outputs(3589));
    outputs(6572) <= not(layer4_outputs(2228));
    outputs(6573) <= not(layer4_outputs(1124));
    outputs(6574) <= not((layer4_outputs(3655)) xor (layer4_outputs(2283)));
    outputs(6575) <= not((layer4_outputs(6259)) xor (layer4_outputs(1153)));
    outputs(6576) <= not((layer4_outputs(5915)) xor (layer4_outputs(7236)));
    outputs(6577) <= not(layer4_outputs(5132));
    outputs(6578) <= not(layer4_outputs(2360)) or (layer4_outputs(4587));
    outputs(6579) <= (layer4_outputs(3326)) xor (layer4_outputs(5168));
    outputs(6580) <= (layer4_outputs(2181)) or (layer4_outputs(6612));
    outputs(6581) <= not(layer4_outputs(6392));
    outputs(6582) <= not((layer4_outputs(2673)) or (layer4_outputs(5780)));
    outputs(6583) <= not((layer4_outputs(4831)) xor (layer4_outputs(3729)));
    outputs(6584) <= (layer4_outputs(3436)) xor (layer4_outputs(5475));
    outputs(6585) <= layer4_outputs(719);
    outputs(6586) <= layer4_outputs(1092);
    outputs(6587) <= not(layer4_outputs(3190));
    outputs(6588) <= not(layer4_outputs(3337));
    outputs(6589) <= (layer4_outputs(1040)) xor (layer4_outputs(5866));
    outputs(6590) <= layer4_outputs(5247);
    outputs(6591) <= layer4_outputs(4761);
    outputs(6592) <= not(layer4_outputs(1755));
    outputs(6593) <= layer4_outputs(2779);
    outputs(6594) <= layer4_outputs(6222);
    outputs(6595) <= layer4_outputs(3893);
    outputs(6596) <= not(layer4_outputs(1895));
    outputs(6597) <= (layer4_outputs(6517)) xor (layer4_outputs(2286));
    outputs(6598) <= not(layer4_outputs(1771));
    outputs(6599) <= not(layer4_outputs(1039));
    outputs(6600) <= not(layer4_outputs(1212));
    outputs(6601) <= layer4_outputs(3244);
    outputs(6602) <= not((layer4_outputs(3259)) or (layer4_outputs(4548)));
    outputs(6603) <= not(layer4_outputs(3419));
    outputs(6604) <= not(layer4_outputs(1748));
    outputs(6605) <= layer4_outputs(5054);
    outputs(6606) <= not(layer4_outputs(3194));
    outputs(6607) <= not(layer4_outputs(3444));
    outputs(6608) <= (layer4_outputs(6552)) and not (layer4_outputs(5750));
    outputs(6609) <= (layer4_outputs(6671)) xor (layer4_outputs(5435));
    outputs(6610) <= (layer4_outputs(3351)) and not (layer4_outputs(5821));
    outputs(6611) <= layer4_outputs(7364);
    outputs(6612) <= not((layer4_outputs(7044)) xor (layer4_outputs(6899)));
    outputs(6613) <= (layer4_outputs(1582)) and (layer4_outputs(3009));
    outputs(6614) <= not(layer4_outputs(2646));
    outputs(6615) <= (layer4_outputs(3225)) xor (layer4_outputs(2631));
    outputs(6616) <= not(layer4_outputs(5972)) or (layer4_outputs(6424));
    outputs(6617) <= not(layer4_outputs(2278));
    outputs(6618) <= layer4_outputs(435);
    outputs(6619) <= not((layer4_outputs(3911)) xor (layer4_outputs(5512)));
    outputs(6620) <= layer4_outputs(5704);
    outputs(6621) <= layer4_outputs(6839);
    outputs(6622) <= layer4_outputs(3550);
    outputs(6623) <= not(layer4_outputs(2932)) or (layer4_outputs(2584));
    outputs(6624) <= layer4_outputs(3479);
    outputs(6625) <= not(layer4_outputs(671)) or (layer4_outputs(5681));
    outputs(6626) <= (layer4_outputs(4396)) xor (layer4_outputs(4122));
    outputs(6627) <= (layer4_outputs(6626)) and not (layer4_outputs(3700));
    outputs(6628) <= not((layer4_outputs(7502)) xor (layer4_outputs(3808)));
    outputs(6629) <= (layer4_outputs(2670)) and not (layer4_outputs(6467));
    outputs(6630) <= not((layer4_outputs(1264)) xor (layer4_outputs(3983)));
    outputs(6631) <= not(layer4_outputs(5466));
    outputs(6632) <= not((layer4_outputs(481)) xor (layer4_outputs(2767)));
    outputs(6633) <= not(layer4_outputs(6559));
    outputs(6634) <= (layer4_outputs(2084)) and not (layer4_outputs(2009));
    outputs(6635) <= layer4_outputs(2405);
    outputs(6636) <= layer4_outputs(4441);
    outputs(6637) <= not(layer4_outputs(862)) or (layer4_outputs(7612));
    outputs(6638) <= (layer4_outputs(5239)) and (layer4_outputs(3271));
    outputs(6639) <= (layer4_outputs(6301)) and not (layer4_outputs(432));
    outputs(6640) <= layer4_outputs(6147);
    outputs(6641) <= layer4_outputs(5474);
    outputs(6642) <= not(layer4_outputs(7261));
    outputs(6643) <= layer4_outputs(1870);
    outputs(6644) <= layer4_outputs(823);
    outputs(6645) <= not(layer4_outputs(5782));
    outputs(6646) <= not(layer4_outputs(6139));
    outputs(6647) <= not(layer4_outputs(5098));
    outputs(6648) <= layer4_outputs(4373);
    outputs(6649) <= not(layer4_outputs(1470)) or (layer4_outputs(939));
    outputs(6650) <= not((layer4_outputs(5611)) xor (layer4_outputs(131)));
    outputs(6651) <= not(layer4_outputs(7650));
    outputs(6652) <= not(layer4_outputs(3481));
    outputs(6653) <= layer4_outputs(1606);
    outputs(6654) <= (layer4_outputs(6775)) xor (layer4_outputs(873));
    outputs(6655) <= layer4_outputs(251);
    outputs(6656) <= layer4_outputs(2016);
    outputs(6657) <= not((layer4_outputs(4410)) or (layer4_outputs(80)));
    outputs(6658) <= layer4_outputs(3390);
    outputs(6659) <= not(layer4_outputs(7318));
    outputs(6660) <= layer4_outputs(3215);
    outputs(6661) <= not(layer4_outputs(3533));
    outputs(6662) <= not(layer4_outputs(1813));
    outputs(6663) <= not(layer4_outputs(4787));
    outputs(6664) <= layer4_outputs(4078);
    outputs(6665) <= layer4_outputs(4694);
    outputs(6666) <= not((layer4_outputs(5957)) and (layer4_outputs(2034)));
    outputs(6667) <= layer4_outputs(5120);
    outputs(6668) <= layer4_outputs(6851);
    outputs(6669) <= not(layer4_outputs(651));
    outputs(6670) <= layer4_outputs(1042);
    outputs(6671) <= (layer4_outputs(4062)) or (layer4_outputs(4934));
    outputs(6672) <= not(layer4_outputs(3826));
    outputs(6673) <= (layer4_outputs(5134)) and not (layer4_outputs(2069));
    outputs(6674) <= not(layer4_outputs(1520));
    outputs(6675) <= not(layer4_outputs(1143));
    outputs(6676) <= not((layer4_outputs(270)) xor (layer4_outputs(300)));
    outputs(6677) <= not(layer4_outputs(1307));
    outputs(6678) <= (layer4_outputs(2193)) xor (layer4_outputs(7633));
    outputs(6679) <= not(layer4_outputs(5773));
    outputs(6680) <= not(layer4_outputs(6017));
    outputs(6681) <= not((layer4_outputs(3475)) xor (layer4_outputs(4834)));
    outputs(6682) <= layer4_outputs(7243);
    outputs(6683) <= layer4_outputs(4169);
    outputs(6684) <= layer4_outputs(4218);
    outputs(6685) <= not(layer4_outputs(6857));
    outputs(6686) <= not((layer4_outputs(5442)) xor (layer4_outputs(318)));
    outputs(6687) <= (layer4_outputs(2370)) xor (layer4_outputs(537));
    outputs(6688) <= (layer4_outputs(7035)) or (layer4_outputs(4306));
    outputs(6689) <= not(layer4_outputs(1719));
    outputs(6690) <= (layer4_outputs(3294)) and (layer4_outputs(6962));
    outputs(6691) <= (layer4_outputs(3946)) xor (layer4_outputs(4652));
    outputs(6692) <= layer4_outputs(5833);
    outputs(6693) <= layer4_outputs(6079);
    outputs(6694) <= not(layer4_outputs(3688)) or (layer4_outputs(3616));
    outputs(6695) <= layer4_outputs(3215);
    outputs(6696) <= (layer4_outputs(5635)) and (layer4_outputs(667));
    outputs(6697) <= not((layer4_outputs(2184)) xor (layer4_outputs(6202)));
    outputs(6698) <= not((layer4_outputs(7633)) xor (layer4_outputs(7256)));
    outputs(6699) <= not(layer4_outputs(3465));
    outputs(6700) <= not((layer4_outputs(2848)) xor (layer4_outputs(4003)));
    outputs(6701) <= (layer4_outputs(1550)) and (layer4_outputs(2428));
    outputs(6702) <= layer4_outputs(1876);
    outputs(6703) <= not((layer4_outputs(6245)) xor (layer4_outputs(2893)));
    outputs(6704) <= not((layer4_outputs(5228)) xor (layer4_outputs(982)));
    outputs(6705) <= (layer4_outputs(4330)) xor (layer4_outputs(7532));
    outputs(6706) <= not((layer4_outputs(5761)) xor (layer4_outputs(2888)));
    outputs(6707) <= (layer4_outputs(5274)) and (layer4_outputs(6310));
    outputs(6708) <= (layer4_outputs(7003)) and not (layer4_outputs(2044));
    outputs(6709) <= not(layer4_outputs(4688)) or (layer4_outputs(3875));
    outputs(6710) <= not((layer4_outputs(7284)) xor (layer4_outputs(780)));
    outputs(6711) <= (layer4_outputs(5770)) or (layer4_outputs(4864));
    outputs(6712) <= layer4_outputs(1832);
    outputs(6713) <= (layer4_outputs(6438)) or (layer4_outputs(3238));
    outputs(6714) <= not(layer4_outputs(7658)) or (layer4_outputs(7263));
    outputs(6715) <= (layer4_outputs(1802)) xor (layer4_outputs(2570));
    outputs(6716) <= not(layer4_outputs(2582));
    outputs(6717) <= not(layer4_outputs(663));
    outputs(6718) <= not(layer4_outputs(7258));
    outputs(6719) <= (layer4_outputs(6471)) and not (layer4_outputs(794));
    outputs(6720) <= not(layer4_outputs(4098));
    outputs(6721) <= not(layer4_outputs(470));
    outputs(6722) <= not(layer4_outputs(974));
    outputs(6723) <= not(layer4_outputs(3590)) or (layer4_outputs(4679));
    outputs(6724) <= not(layer4_outputs(2454)) or (layer4_outputs(4706));
    outputs(6725) <= (layer4_outputs(2701)) xor (layer4_outputs(3839));
    outputs(6726) <= layer4_outputs(666);
    outputs(6727) <= not((layer4_outputs(5046)) and (layer4_outputs(447)));
    outputs(6728) <= not(layer4_outputs(149));
    outputs(6729) <= not((layer4_outputs(2085)) xor (layer4_outputs(7635)));
    outputs(6730) <= layer4_outputs(7493);
    outputs(6731) <= not(layer4_outputs(4362));
    outputs(6732) <= (layer4_outputs(701)) and not (layer4_outputs(2493));
    outputs(6733) <= layer4_outputs(1169);
    outputs(6734) <= not(layer4_outputs(5272));
    outputs(6735) <= layer4_outputs(5287);
    outputs(6736) <= (layer4_outputs(6347)) xor (layer4_outputs(6215));
    outputs(6737) <= layer4_outputs(1120);
    outputs(6738) <= not((layer4_outputs(4458)) xor (layer4_outputs(4839)));
    outputs(6739) <= not((layer4_outputs(2964)) xor (layer4_outputs(6047)));
    outputs(6740) <= not(layer4_outputs(2703));
    outputs(6741) <= (layer4_outputs(5714)) xor (layer4_outputs(3720));
    outputs(6742) <= not((layer4_outputs(3878)) or (layer4_outputs(3029)));
    outputs(6743) <= not((layer4_outputs(6062)) xor (layer4_outputs(6485)));
    outputs(6744) <= (layer4_outputs(1703)) and not (layer4_outputs(7434));
    outputs(6745) <= not(layer4_outputs(5758));
    outputs(6746) <= not(layer4_outputs(3821));
    outputs(6747) <= not(layer4_outputs(4848)) or (layer4_outputs(6938));
    outputs(6748) <= layer4_outputs(2802);
    outputs(6749) <= not(layer4_outputs(4784)) or (layer4_outputs(4402));
    outputs(6750) <= layer4_outputs(7439);
    outputs(6751) <= layer4_outputs(7265);
    outputs(6752) <= not(layer4_outputs(6448));
    outputs(6753) <= not(layer4_outputs(2065)) or (layer4_outputs(5752));
    outputs(6754) <= layer4_outputs(4690);
    outputs(6755) <= not((layer4_outputs(3651)) and (layer4_outputs(6425)));
    outputs(6756) <= layer4_outputs(7441);
    outputs(6757) <= (layer4_outputs(2135)) and not (layer4_outputs(3065));
    outputs(6758) <= not(layer4_outputs(4359));
    outputs(6759) <= (layer4_outputs(1731)) xor (layer4_outputs(3056));
    outputs(6760) <= (layer4_outputs(5023)) xor (layer4_outputs(2114));
    outputs(6761) <= not((layer4_outputs(5011)) xor (layer4_outputs(6262)));
    outputs(6762) <= not((layer4_outputs(4859)) or (layer4_outputs(4137)));
    outputs(6763) <= (layer4_outputs(273)) xor (layer4_outputs(2780));
    outputs(6764) <= (layer4_outputs(4661)) xor (layer4_outputs(5685));
    outputs(6765) <= layer4_outputs(1515);
    outputs(6766) <= (layer4_outputs(3744)) and not (layer4_outputs(2044));
    outputs(6767) <= not(layer4_outputs(6985));
    outputs(6768) <= (layer4_outputs(4159)) and not (layer4_outputs(3689));
    outputs(6769) <= not(layer4_outputs(1165));
    outputs(6770) <= (layer4_outputs(7292)) and not (layer4_outputs(2136));
    outputs(6771) <= (layer4_outputs(2628)) xor (layer4_outputs(3893));
    outputs(6772) <= layer4_outputs(5150);
    outputs(6773) <= layer4_outputs(3332);
    outputs(6774) <= not(layer4_outputs(6750)) or (layer4_outputs(2502));
    outputs(6775) <= (layer4_outputs(2478)) xor (layer4_outputs(6932));
    outputs(6776) <= not(layer4_outputs(4833));
    outputs(6777) <= layer4_outputs(5913);
    outputs(6778) <= not(layer4_outputs(3040)) or (layer4_outputs(6850));
    outputs(6779) <= layer4_outputs(3393);
    outputs(6780) <= not(layer4_outputs(124));
    outputs(6781) <= layer4_outputs(3361);
    outputs(6782) <= (layer4_outputs(1903)) or (layer4_outputs(2289));
    outputs(6783) <= layer4_outputs(1385);
    outputs(6784) <= not((layer4_outputs(6108)) xor (layer4_outputs(2695)));
    outputs(6785) <= layer4_outputs(6839);
    outputs(6786) <= (layer4_outputs(7537)) xor (layer4_outputs(3363));
    outputs(6787) <= (layer4_outputs(1681)) and not (layer4_outputs(6534));
    outputs(6788) <= not(layer4_outputs(6918));
    outputs(6789) <= not(layer4_outputs(4328));
    outputs(6790) <= not(layer4_outputs(5020));
    outputs(6791) <= not((layer4_outputs(5641)) and (layer4_outputs(198)));
    outputs(6792) <= not((layer4_outputs(2882)) xor (layer4_outputs(528)));
    outputs(6793) <= (layer4_outputs(3791)) xor (layer4_outputs(2907));
    outputs(6794) <= layer4_outputs(4);
    outputs(6795) <= not(layer4_outputs(2808)) or (layer4_outputs(5562));
    outputs(6796) <= not(layer4_outputs(6760));
    outputs(6797) <= not(layer4_outputs(7499)) or (layer4_outputs(6151));
    outputs(6798) <= not(layer4_outputs(2214));
    outputs(6799) <= layer4_outputs(985);
    outputs(6800) <= (layer4_outputs(4435)) and not (layer4_outputs(5576));
    outputs(6801) <= layer4_outputs(2401);
    outputs(6802) <= not(layer4_outputs(1523));
    outputs(6803) <= (layer4_outputs(3369)) xor (layer4_outputs(1943));
    outputs(6804) <= layer4_outputs(5310);
    outputs(6805) <= not((layer4_outputs(6472)) xor (layer4_outputs(5043)));
    outputs(6806) <= layer4_outputs(2578);
    outputs(6807) <= (layer4_outputs(7522)) xor (layer4_outputs(2733));
    outputs(6808) <= not(layer4_outputs(6119)) or (layer4_outputs(3182));
    outputs(6809) <= not(layer4_outputs(1379)) or (layer4_outputs(3830));
    outputs(6810) <= layer4_outputs(5847);
    outputs(6811) <= not(layer4_outputs(6864));
    outputs(6812) <= (layer4_outputs(6049)) xor (layer4_outputs(7530));
    outputs(6813) <= layer4_outputs(1284);
    outputs(6814) <= not(layer4_outputs(1013)) or (layer4_outputs(91));
    outputs(6815) <= not((layer4_outputs(2449)) xor (layer4_outputs(1562)));
    outputs(6816) <= not((layer4_outputs(6353)) xor (layer4_outputs(5193)));
    outputs(6817) <= (layer4_outputs(2514)) xor (layer4_outputs(921));
    outputs(6818) <= (layer4_outputs(3986)) and not (layer4_outputs(6838));
    outputs(6819) <= layer4_outputs(367);
    outputs(6820) <= layer4_outputs(1982);
    outputs(6821) <= not(layer4_outputs(3482));
    outputs(6822) <= layer4_outputs(7092);
    outputs(6823) <= layer4_outputs(4440);
    outputs(6824) <= not(layer4_outputs(7332));
    outputs(6825) <= layer4_outputs(4524);
    outputs(6826) <= (layer4_outputs(4572)) xor (layer4_outputs(779));
    outputs(6827) <= layer4_outputs(7379);
    outputs(6828) <= not(layer4_outputs(6163));
    outputs(6829) <= (layer4_outputs(990)) xor (layer4_outputs(1741));
    outputs(6830) <= layer4_outputs(3990);
    outputs(6831) <= layer4_outputs(494);
    outputs(6832) <= not((layer4_outputs(5943)) or (layer4_outputs(3404)));
    outputs(6833) <= not(layer4_outputs(2952));
    outputs(6834) <= not(layer4_outputs(1757));
    outputs(6835) <= (layer4_outputs(491)) and not (layer4_outputs(4860));
    outputs(6836) <= layer4_outputs(168);
    outputs(6837) <= (layer4_outputs(2992)) and not (layer4_outputs(3569));
    outputs(6838) <= not((layer4_outputs(3743)) or (layer4_outputs(6498)));
    outputs(6839) <= layer4_outputs(2595);
    outputs(6840) <= not((layer4_outputs(4418)) xor (layer4_outputs(5996)));
    outputs(6841) <= not(layer4_outputs(2621));
    outputs(6842) <= (layer4_outputs(2754)) xor (layer4_outputs(5153));
    outputs(6843) <= layer4_outputs(3921);
    outputs(6844) <= layer4_outputs(2350);
    outputs(6845) <= (layer4_outputs(6494)) xor (layer4_outputs(4875));
    outputs(6846) <= not(layer4_outputs(4152));
    outputs(6847) <= layer4_outputs(7357);
    outputs(6848) <= layer4_outputs(5920);
    outputs(6849) <= not((layer4_outputs(95)) xor (layer4_outputs(2867)));
    outputs(6850) <= not(layer4_outputs(6465));
    outputs(6851) <= not((layer4_outputs(2821)) and (layer4_outputs(505)));
    outputs(6852) <= (layer4_outputs(5709)) or (layer4_outputs(2605));
    outputs(6853) <= layer4_outputs(226);
    outputs(6854) <= layer4_outputs(4728);
    outputs(6855) <= (layer4_outputs(5351)) and not (layer4_outputs(1867));
    outputs(6856) <= not((layer4_outputs(3687)) and (layer4_outputs(2571)));
    outputs(6857) <= not(layer4_outputs(2586));
    outputs(6858) <= layer4_outputs(7346);
    outputs(6859) <= not((layer4_outputs(3503)) xor (layer4_outputs(4664)));
    outputs(6860) <= not((layer4_outputs(707)) xor (layer4_outputs(3260)));
    outputs(6861) <= not(layer4_outputs(4701));
    outputs(6862) <= (layer4_outputs(4200)) or (layer4_outputs(157));
    outputs(6863) <= not((layer4_outputs(3007)) xor (layer4_outputs(6374)));
    outputs(6864) <= layer4_outputs(7238);
    outputs(6865) <= (layer4_outputs(1084)) and not (layer4_outputs(2137));
    outputs(6866) <= (layer4_outputs(229)) and (layer4_outputs(7461));
    outputs(6867) <= (layer4_outputs(4026)) xor (layer4_outputs(6457));
    outputs(6868) <= not(layer4_outputs(6386));
    outputs(6869) <= not((layer4_outputs(1015)) or (layer4_outputs(4623)));
    outputs(6870) <= layer4_outputs(4456);
    outputs(6871) <= not((layer4_outputs(876)) xor (layer4_outputs(485)));
    outputs(6872) <= (layer4_outputs(5112)) xor (layer4_outputs(4523));
    outputs(6873) <= not((layer4_outputs(2192)) and (layer4_outputs(2287)));
    outputs(6874) <= layer4_outputs(3975);
    outputs(6875) <= layer4_outputs(4102);
    outputs(6876) <= layer4_outputs(6079);
    outputs(6877) <= not((layer4_outputs(7176)) or (layer4_outputs(5206)));
    outputs(6878) <= not(layer4_outputs(5974));
    outputs(6879) <= (layer4_outputs(1920)) xor (layer4_outputs(6953));
    outputs(6880) <= (layer4_outputs(2978)) and not (layer4_outputs(5256));
    outputs(6881) <= (layer4_outputs(1146)) and not (layer4_outputs(1691));
    outputs(6882) <= not((layer4_outputs(1868)) and (layer4_outputs(7021)));
    outputs(6883) <= (layer4_outputs(5636)) xor (layer4_outputs(3680));
    outputs(6884) <= not(layer4_outputs(2367));
    outputs(6885) <= layer4_outputs(5393);
    outputs(6886) <= not((layer4_outputs(427)) xor (layer4_outputs(5650)));
    outputs(6887) <= layer4_outputs(6649);
    outputs(6888) <= not(layer4_outputs(4149));
    outputs(6889) <= not(layer4_outputs(1963));
    outputs(6890) <= layer4_outputs(5325);
    outputs(6891) <= not(layer4_outputs(2034));
    outputs(6892) <= layer4_outputs(7013);
    outputs(6893) <= not((layer4_outputs(5500)) xor (layer4_outputs(35)));
    outputs(6894) <= (layer4_outputs(5380)) or (layer4_outputs(540));
    outputs(6895) <= not((layer4_outputs(4344)) xor (layer4_outputs(3675)));
    outputs(6896) <= not(layer4_outputs(5385));
    outputs(6897) <= (layer4_outputs(7474)) xor (layer4_outputs(2565));
    outputs(6898) <= layer4_outputs(7183);
    outputs(6899) <= not(layer4_outputs(222));
    outputs(6900) <= (layer4_outputs(935)) or (layer4_outputs(3453));
    outputs(6901) <= not(layer4_outputs(1298));
    outputs(6902) <= not(layer4_outputs(5576));
    outputs(6903) <= (layer4_outputs(3487)) and (layer4_outputs(3912));
    outputs(6904) <= not((layer4_outputs(5737)) and (layer4_outputs(1692)));
    outputs(6905) <= layer4_outputs(4529);
    outputs(6906) <= not(layer4_outputs(4268));
    outputs(6907) <= not(layer4_outputs(1099));
    outputs(6908) <= not(layer4_outputs(6288));
    outputs(6909) <= not((layer4_outputs(3694)) and (layer4_outputs(3047)));
    outputs(6910) <= not(layer4_outputs(4938));
    outputs(6911) <= layer4_outputs(6357);
    outputs(6912) <= not(layer4_outputs(611)) or (layer4_outputs(6123));
    outputs(6913) <= not(layer4_outputs(892));
    outputs(6914) <= not(layer4_outputs(3446));
    outputs(6915) <= layer4_outputs(5676);
    outputs(6916) <= layer4_outputs(1068);
    outputs(6917) <= (layer4_outputs(6560)) and not (layer4_outputs(4886));
    outputs(6918) <= layer4_outputs(4284);
    outputs(6919) <= not(layer4_outputs(1290));
    outputs(6920) <= not((layer4_outputs(3725)) xor (layer4_outputs(7231)));
    outputs(6921) <= (layer4_outputs(5560)) and (layer4_outputs(2282));
    outputs(6922) <= layer4_outputs(366);
    outputs(6923) <= not(layer4_outputs(7148));
    outputs(6924) <= (layer4_outputs(5162)) and not (layer4_outputs(1997));
    outputs(6925) <= (layer4_outputs(741)) and not (layer4_outputs(7356));
    outputs(6926) <= not(layer4_outputs(4776));
    outputs(6927) <= not((layer4_outputs(4544)) xor (layer4_outputs(7178)));
    outputs(6928) <= layer4_outputs(5526);
    outputs(6929) <= not(layer4_outputs(1428));
    outputs(6930) <= not(layer4_outputs(2425));
    outputs(6931) <= not((layer4_outputs(6340)) and (layer4_outputs(1282)));
    outputs(6932) <= not((layer4_outputs(1826)) and (layer4_outputs(7144)));
    outputs(6933) <= not(layer4_outputs(7310));
    outputs(6934) <= not(layer4_outputs(3639));
    outputs(6935) <= not((layer4_outputs(189)) or (layer4_outputs(5372)));
    outputs(6936) <= not(layer4_outputs(3248));
    outputs(6937) <= layer4_outputs(5443);
    outputs(6938) <= not(layer4_outputs(1314));
    outputs(6939) <= not(layer4_outputs(4377)) or (layer4_outputs(4758));
    outputs(6940) <= layer4_outputs(5801);
    outputs(6941) <= not(layer4_outputs(4746));
    outputs(6942) <= layer4_outputs(2995);
    outputs(6943) <= not(layer4_outputs(4502));
    outputs(6944) <= layer4_outputs(895);
    outputs(6945) <= not(layer4_outputs(3653));
    outputs(6946) <= not(layer4_outputs(2112));
    outputs(6947) <= not(layer4_outputs(2470));
    outputs(6948) <= not(layer4_outputs(4304));
    outputs(6949) <= layer4_outputs(2722);
    outputs(6950) <= (layer4_outputs(6315)) and (layer4_outputs(6821));
    outputs(6951) <= not((layer4_outputs(6321)) xor (layer4_outputs(569)));
    outputs(6952) <= (layer4_outputs(661)) xor (layer4_outputs(6780));
    outputs(6953) <= layer4_outputs(3686);
    outputs(6954) <= not((layer4_outputs(3820)) xor (layer4_outputs(3491)));
    outputs(6955) <= not(layer4_outputs(2643));
    outputs(6956) <= not(layer4_outputs(2630));
    outputs(6957) <= not(layer4_outputs(1421));
    outputs(6958) <= layer4_outputs(5810);
    outputs(6959) <= not(layer4_outputs(6979));
    outputs(6960) <= not((layer4_outputs(1227)) and (layer4_outputs(2562)));
    outputs(6961) <= (layer4_outputs(6035)) and (layer4_outputs(3704));
    outputs(6962) <= layer4_outputs(6443);
    outputs(6963) <= not((layer4_outputs(894)) or (layer4_outputs(223)));
    outputs(6964) <= not(layer4_outputs(6766));
    outputs(6965) <= layer4_outputs(5689);
    outputs(6966) <= (layer4_outputs(797)) and (layer4_outputs(6989));
    outputs(6967) <= not(layer4_outputs(2047));
    outputs(6968) <= not(layer4_outputs(4340));
    outputs(6969) <= not((layer4_outputs(4097)) xor (layer4_outputs(2541)));
    outputs(6970) <= (layer4_outputs(1208)) xor (layer4_outputs(1602));
    outputs(6971) <= not(layer4_outputs(4983));
    outputs(6972) <= layer4_outputs(6993);
    outputs(6973) <= not(layer4_outputs(6606));
    outputs(6974) <= layer4_outputs(5424);
    outputs(6975) <= (layer4_outputs(6726)) or (layer4_outputs(1147));
    outputs(6976) <= not(layer4_outputs(1513));
    outputs(6977) <= (layer4_outputs(5583)) and (layer4_outputs(6146));
    outputs(6978) <= not(layer4_outputs(3863));
    outputs(6979) <= not((layer4_outputs(7151)) xor (layer4_outputs(2593)));
    outputs(6980) <= not(layer4_outputs(1703));
    outputs(6981) <= not((layer4_outputs(2358)) or (layer4_outputs(1215)));
    outputs(6982) <= layer4_outputs(2441);
    outputs(6983) <= layer4_outputs(1098);
    outputs(6984) <= layer4_outputs(6936);
    outputs(6985) <= not(layer4_outputs(2074));
    outputs(6986) <= not(layer4_outputs(3851));
    outputs(6987) <= (layer4_outputs(5338)) xor (layer4_outputs(1887));
    outputs(6988) <= not(layer4_outputs(7527));
    outputs(6989) <= layer4_outputs(4164);
    outputs(6990) <= layer4_outputs(2353);
    outputs(6991) <= (layer4_outputs(1302)) xor (layer4_outputs(3401));
    outputs(6992) <= not(layer4_outputs(1781));
    outputs(6993) <= (layer4_outputs(661)) xor (layer4_outputs(4514));
    outputs(6994) <= layer4_outputs(7674);
    outputs(6995) <= not(layer4_outputs(4806));
    outputs(6996) <= not((layer4_outputs(2346)) xor (layer4_outputs(3764)));
    outputs(6997) <= not((layer4_outputs(946)) xor (layer4_outputs(1580)));
    outputs(6998) <= layer4_outputs(7260);
    outputs(6999) <= layer4_outputs(1687);
    outputs(7000) <= not((layer4_outputs(6106)) xor (layer4_outputs(4629)));
    outputs(7001) <= not(layer4_outputs(6901));
    outputs(7002) <= (layer4_outputs(174)) and (layer4_outputs(4692));
    outputs(7003) <= layer4_outputs(5346);
    outputs(7004) <= not(layer4_outputs(2142));
    outputs(7005) <= not(layer4_outputs(6364));
    outputs(7006) <= not(layer4_outputs(2002));
    outputs(7007) <= not(layer4_outputs(3064));
    outputs(7008) <= not(layer4_outputs(798));
    outputs(7009) <= not(layer4_outputs(6165));
    outputs(7010) <= not(layer4_outputs(3063));
    outputs(7011) <= not(layer4_outputs(2856));
    outputs(7012) <= not((layer4_outputs(93)) or (layer4_outputs(1906)));
    outputs(7013) <= layer4_outputs(7602);
    outputs(7014) <= layer4_outputs(4352);
    outputs(7015) <= (layer4_outputs(5893)) xor (layer4_outputs(295));
    outputs(7016) <= not(layer4_outputs(346));
    outputs(7017) <= layer4_outputs(197);
    outputs(7018) <= not(layer4_outputs(4942));
    outputs(7019) <= not(layer4_outputs(3119));
    outputs(7020) <= not((layer4_outputs(1334)) xor (layer4_outputs(7538)));
    outputs(7021) <= not(layer4_outputs(6694));
    outputs(7022) <= not((layer4_outputs(7377)) xor (layer4_outputs(645)));
    outputs(7023) <= not((layer4_outputs(4429)) xor (layer4_outputs(5233)));
    outputs(7024) <= layer4_outputs(416);
    outputs(7025) <= not(layer4_outputs(6955));
    outputs(7026) <= layer4_outputs(7280);
    outputs(7027) <= layer4_outputs(5611);
    outputs(7028) <= (layer4_outputs(6718)) and not (layer4_outputs(3352));
    outputs(7029) <= not(layer4_outputs(7486));
    outputs(7030) <= not((layer4_outputs(6551)) or (layer4_outputs(3842)));
    outputs(7031) <= layer4_outputs(2108);
    outputs(7032) <= (layer4_outputs(2229)) and (layer4_outputs(4425));
    outputs(7033) <= (layer4_outputs(3623)) and not (layer4_outputs(45));
    outputs(7034) <= layer4_outputs(6424);
    outputs(7035) <= not(layer4_outputs(3458));
    outputs(7036) <= layer4_outputs(4926);
    outputs(7037) <= layer4_outputs(4376);
    outputs(7038) <= layer4_outputs(6540);
    outputs(7039) <= not((layer4_outputs(6150)) and (layer4_outputs(3)));
    outputs(7040) <= (layer4_outputs(6360)) and (layer4_outputs(587));
    outputs(7041) <= layer4_outputs(3278);
    outputs(7042) <= not(layer4_outputs(1300));
    outputs(7043) <= (layer4_outputs(1298)) and not (layer4_outputs(5203));
    outputs(7044) <= (layer4_outputs(5397)) and not (layer4_outputs(1867));
    outputs(7045) <= not(layer4_outputs(7626));
    outputs(7046) <= not((layer4_outputs(313)) xor (layer4_outputs(4394)));
    outputs(7047) <= not((layer4_outputs(5204)) xor (layer4_outputs(3354)));
    outputs(7048) <= not(layer4_outputs(7037));
    outputs(7049) <= layer4_outputs(5322);
    outputs(7050) <= layer4_outputs(6707);
    outputs(7051) <= layer4_outputs(3834);
    outputs(7052) <= (layer4_outputs(4844)) and not (layer4_outputs(2408));
    outputs(7053) <= not(layer4_outputs(6166)) or (layer4_outputs(472));
    outputs(7054) <= not((layer4_outputs(2406)) or (layer4_outputs(7204)));
    outputs(7055) <= layer4_outputs(5563);
    outputs(7056) <= layer4_outputs(3819);
    outputs(7057) <= not((layer4_outputs(161)) or (layer4_outputs(2924)));
    outputs(7058) <= not(layer4_outputs(5180));
    outputs(7059) <= not(layer4_outputs(7372));
    outputs(7060) <= not((layer4_outputs(1516)) xor (layer4_outputs(6284)));
    outputs(7061) <= (layer4_outputs(7599)) and not (layer4_outputs(3020));
    outputs(7062) <= not((layer4_outputs(1713)) xor (layer4_outputs(7615)));
    outputs(7063) <= layer4_outputs(36);
    outputs(7064) <= not((layer4_outputs(5282)) xor (layer4_outputs(3857)));
    outputs(7065) <= not(layer4_outputs(5519));
    outputs(7066) <= not((layer4_outputs(4119)) xor (layer4_outputs(170)));
    outputs(7067) <= layer4_outputs(4321);
    outputs(7068) <= (layer4_outputs(6804)) xor (layer4_outputs(3288));
    outputs(7069) <= not(layer4_outputs(1631));
    outputs(7070) <= layer4_outputs(5490);
    outputs(7071) <= (layer4_outputs(7226)) xor (layer4_outputs(3265));
    outputs(7072) <= (layer4_outputs(7117)) and not (layer4_outputs(513));
    outputs(7073) <= layer4_outputs(4766);
    outputs(7074) <= layer4_outputs(5261);
    outputs(7075) <= layer4_outputs(5831);
    outputs(7076) <= not((layer4_outputs(4555)) xor (layer4_outputs(4392)));
    outputs(7077) <= layer4_outputs(2390);
    outputs(7078) <= layer4_outputs(6792);
    outputs(7079) <= not(layer4_outputs(590));
    outputs(7080) <= not(layer4_outputs(5813));
    outputs(7081) <= layer4_outputs(4861);
    outputs(7082) <= layer4_outputs(3609);
    outputs(7083) <= not((layer4_outputs(5612)) xor (layer4_outputs(5649)));
    outputs(7084) <= layer4_outputs(2456);
    outputs(7085) <= (layer4_outputs(2802)) and (layer4_outputs(436));
    outputs(7086) <= not((layer4_outputs(5229)) xor (layer4_outputs(163)));
    outputs(7087) <= not((layer4_outputs(750)) xor (layer4_outputs(4345)));
    outputs(7088) <= layer4_outputs(4924);
    outputs(7089) <= not(layer4_outputs(1877)) or (layer4_outputs(2832));
    outputs(7090) <= layer4_outputs(3417);
    outputs(7091) <= (layer4_outputs(3644)) or (layer4_outputs(4912));
    outputs(7092) <= (layer4_outputs(5315)) and (layer4_outputs(5184));
    outputs(7093) <= not(layer4_outputs(3625));
    outputs(7094) <= (layer4_outputs(6863)) xor (layer4_outputs(4580));
    outputs(7095) <= not((layer4_outputs(5953)) xor (layer4_outputs(2781)));
    outputs(7096) <= not((layer4_outputs(521)) and (layer4_outputs(6038)));
    outputs(7097) <= not((layer4_outputs(1597)) xor (layer4_outputs(3360)));
    outputs(7098) <= layer4_outputs(417);
    outputs(7099) <= (layer4_outputs(4941)) xor (layer4_outputs(1940));
    outputs(7100) <= not((layer4_outputs(4445)) xor (layer4_outputs(344)));
    outputs(7101) <= (layer4_outputs(7353)) and not (layer4_outputs(4657));
    outputs(7102) <= not((layer4_outputs(2068)) xor (layer4_outputs(1705)));
    outputs(7103) <= not((layer4_outputs(56)) and (layer4_outputs(5912)));
    outputs(7104) <= (layer4_outputs(6807)) xor (layer4_outputs(1668));
    outputs(7105) <= not(layer4_outputs(6772));
    outputs(7106) <= (layer4_outputs(6575)) or (layer4_outputs(5428));
    outputs(7107) <= not((layer4_outputs(6243)) xor (layer4_outputs(3675)));
    outputs(7108) <= layer4_outputs(4321);
    outputs(7109) <= not(layer4_outputs(3045));
    outputs(7110) <= (layer4_outputs(7446)) xor (layer4_outputs(2029));
    outputs(7111) <= layer4_outputs(1064);
    outputs(7112) <= layer4_outputs(356);
    outputs(7113) <= layer4_outputs(3226);
    outputs(7114) <= not(layer4_outputs(6954));
    outputs(7115) <= layer4_outputs(3492);
    outputs(7116) <= (layer4_outputs(6244)) and not (layer4_outputs(5293));
    outputs(7117) <= layer4_outputs(1996);
    outputs(7118) <= not(layer4_outputs(4450));
    outputs(7119) <= not((layer4_outputs(3113)) and (layer4_outputs(2631)));
    outputs(7120) <= layer4_outputs(5399);
    outputs(7121) <= layer4_outputs(5497);
    outputs(7122) <= (layer4_outputs(4259)) xor (layer4_outputs(87));
    outputs(7123) <= layer4_outputs(2832);
    outputs(7124) <= not((layer4_outputs(257)) and (layer4_outputs(5369)));
    outputs(7125) <= (layer4_outputs(6303)) xor (layer4_outputs(2572));
    outputs(7126) <= (layer4_outputs(1503)) and not (layer4_outputs(2313));
    outputs(7127) <= layer4_outputs(7504);
    outputs(7128) <= not(layer4_outputs(2091));
    outputs(7129) <= not(layer4_outputs(916));
    outputs(7130) <= (layer4_outputs(2793)) or (layer4_outputs(6652));
    outputs(7131) <= not((layer4_outputs(3676)) or (layer4_outputs(3420)));
    outputs(7132) <= not((layer4_outputs(3552)) xor (layer4_outputs(384)));
    outputs(7133) <= not(layer4_outputs(7573));
    outputs(7134) <= (layer4_outputs(5739)) or (layer4_outputs(3518));
    outputs(7135) <= not((layer4_outputs(6869)) or (layer4_outputs(832)));
    outputs(7136) <= not(layer4_outputs(6077)) or (layer4_outputs(3318));
    outputs(7137) <= layer4_outputs(5459);
    outputs(7138) <= layer4_outputs(5295);
    outputs(7139) <= not(layer4_outputs(7296));
    outputs(7140) <= (layer4_outputs(6359)) and (layer4_outputs(7198));
    outputs(7141) <= not(layer4_outputs(5531));
    outputs(7142) <= (layer4_outputs(3344)) and (layer4_outputs(4760));
    outputs(7143) <= (layer4_outputs(4583)) and (layer4_outputs(3524));
    outputs(7144) <= (layer4_outputs(719)) xor (layer4_outputs(79));
    outputs(7145) <= not(layer4_outputs(6473));
    outputs(7146) <= not(layer4_outputs(7390));
    outputs(7147) <= not(layer4_outputs(3624)) or (layer4_outputs(1673));
    outputs(7148) <= (layer4_outputs(5070)) xor (layer4_outputs(761));
    outputs(7149) <= layer4_outputs(5541);
    outputs(7150) <= not(layer4_outputs(3262));
    outputs(7151) <= (layer4_outputs(5528)) and (layer4_outputs(1940));
    outputs(7152) <= (layer4_outputs(1114)) and not (layer4_outputs(1516));
    outputs(7153) <= layer4_outputs(7205);
    outputs(7154) <= not(layer4_outputs(1512));
    outputs(7155) <= layer4_outputs(3620);
    outputs(7156) <= (layer4_outputs(4141)) and (layer4_outputs(4607));
    outputs(7157) <= not(layer4_outputs(1735));
    outputs(7158) <= not(layer4_outputs(6783));
    outputs(7159) <= not(layer4_outputs(586));
    outputs(7160) <= not((layer4_outputs(2190)) xor (layer4_outputs(5403)));
    outputs(7161) <= layer4_outputs(2884);
    outputs(7162) <= layer4_outputs(2393);
    outputs(7163) <= not((layer4_outputs(6025)) xor (layer4_outputs(7522)));
    outputs(7164) <= (layer4_outputs(6919)) xor (layer4_outputs(3405));
    outputs(7165) <= layer4_outputs(5145);
    outputs(7166) <= not((layer4_outputs(5938)) or (layer4_outputs(7119)));
    outputs(7167) <= not((layer4_outputs(7401)) xor (layer4_outputs(1423)));
    outputs(7168) <= not((layer4_outputs(5204)) or (layer4_outputs(4192)));
    outputs(7169) <= not(layer4_outputs(5037));
    outputs(7170) <= layer4_outputs(4267);
    outputs(7171) <= layer4_outputs(5524);
    outputs(7172) <= not(layer4_outputs(3451));
    outputs(7173) <= not((layer4_outputs(1604)) and (layer4_outputs(2945)));
    outputs(7174) <= (layer4_outputs(5807)) xor (layer4_outputs(7541));
    outputs(7175) <= not((layer4_outputs(1215)) xor (layer4_outputs(5680)));
    outputs(7176) <= not(layer4_outputs(2199));
    outputs(7177) <= layer4_outputs(2477);
    outputs(7178) <= not(layer4_outputs(3927)) or (layer4_outputs(4793));
    outputs(7179) <= not(layer4_outputs(6778));
    outputs(7180) <= layer4_outputs(7205);
    outputs(7181) <= layer4_outputs(5246);
    outputs(7182) <= (layer4_outputs(5299)) xor (layer4_outputs(5335));
    outputs(7183) <= not(layer4_outputs(6771));
    outputs(7184) <= (layer4_outputs(7600)) and not (layer4_outputs(6974));
    outputs(7185) <= not(layer4_outputs(2126));
    outputs(7186) <= not(layer4_outputs(6637));
    outputs(7187) <= not(layer4_outputs(7381));
    outputs(7188) <= layer4_outputs(1856);
    outputs(7189) <= not(layer4_outputs(5601));
    outputs(7190) <= layer4_outputs(6875);
    outputs(7191) <= (layer4_outputs(7465)) and (layer4_outputs(7029));
    outputs(7192) <= (layer4_outputs(7609)) and (layer4_outputs(2602));
    outputs(7193) <= (layer4_outputs(3021)) and not (layer4_outputs(4332));
    outputs(7194) <= not(layer4_outputs(6905));
    outputs(7195) <= not(layer4_outputs(6286));
    outputs(7196) <= not(layer4_outputs(2712));
    outputs(7197) <= not(layer4_outputs(6051));
    outputs(7198) <= not((layer4_outputs(6271)) or (layer4_outputs(6687)));
    outputs(7199) <= (layer4_outputs(5066)) xor (layer4_outputs(486));
    outputs(7200) <= layer4_outputs(4375);
    outputs(7201) <= not((layer4_outputs(4368)) or (layer4_outputs(5349)));
    outputs(7202) <= layer4_outputs(2374);
    outputs(7203) <= not((layer4_outputs(1917)) xor (layer4_outputs(6056)));
    outputs(7204) <= (layer4_outputs(395)) xor (layer4_outputs(1474));
    outputs(7205) <= not(layer4_outputs(532));
    outputs(7206) <= (layer4_outputs(2918)) and not (layer4_outputs(3356));
    outputs(7207) <= layer4_outputs(5852);
    outputs(7208) <= not((layer4_outputs(625)) xor (layer4_outputs(7015)));
    outputs(7209) <= layer4_outputs(1186);
    outputs(7210) <= layer4_outputs(653);
    outputs(7211) <= not(layer4_outputs(596));
    outputs(7212) <= (layer4_outputs(2971)) and not (layer4_outputs(5151));
    outputs(7213) <= not((layer4_outputs(1519)) xor (layer4_outputs(4751)));
    outputs(7214) <= (layer4_outputs(1046)) or (layer4_outputs(3956));
    outputs(7215) <= (layer4_outputs(4316)) and not (layer4_outputs(3672));
    outputs(7216) <= not((layer4_outputs(472)) xor (layer4_outputs(5715)));
    outputs(7217) <= not(layer4_outputs(7216)) or (layer4_outputs(6683));
    outputs(7218) <= not(layer4_outputs(1800)) or (layer4_outputs(1079));
    outputs(7219) <= (layer4_outputs(7003)) and (layer4_outputs(1030));
    outputs(7220) <= layer4_outputs(1966);
    outputs(7221) <= layer4_outputs(7077);
    outputs(7222) <= layer4_outputs(5968);
    outputs(7223) <= not(layer4_outputs(3392));
    outputs(7224) <= not((layer4_outputs(7264)) xor (layer4_outputs(7529)));
    outputs(7225) <= (layer4_outputs(598)) xor (layer4_outputs(3085));
    outputs(7226) <= not((layer4_outputs(4411)) and (layer4_outputs(4109)));
    outputs(7227) <= not(layer4_outputs(4717));
    outputs(7228) <= (layer4_outputs(6387)) and not (layer4_outputs(897));
    outputs(7229) <= not(layer4_outputs(5703));
    outputs(7230) <= layer4_outputs(426);
    outputs(7231) <= layer4_outputs(1534);
    outputs(7232) <= not(layer4_outputs(5260));
    outputs(7233) <= (layer4_outputs(6558)) xor (layer4_outputs(5937));
    outputs(7234) <= not(layer4_outputs(5473)) or (layer4_outputs(6969));
    outputs(7235) <= not(layer4_outputs(4869)) or (layer4_outputs(3397));
    outputs(7236) <= layer4_outputs(6061);
    outputs(7237) <= not(layer4_outputs(176));
    outputs(7238) <= not(layer4_outputs(321));
    outputs(7239) <= not((layer4_outputs(4314)) xor (layer4_outputs(90)));
    outputs(7240) <= not((layer4_outputs(5730)) xor (layer4_outputs(2023)));
    outputs(7241) <= (layer4_outputs(544)) xor (layer4_outputs(245));
    outputs(7242) <= not((layer4_outputs(4475)) xor (layer4_outputs(3590)));
    outputs(7243) <= layer4_outputs(6576);
    outputs(7244) <= (layer4_outputs(4239)) and not (layer4_outputs(7622));
    outputs(7245) <= layer4_outputs(5927);
    outputs(7246) <= not(layer4_outputs(2303));
    outputs(7247) <= layer4_outputs(3436);
    outputs(7248) <= not(layer4_outputs(4136));
    outputs(7249) <= layer4_outputs(2540);
    outputs(7250) <= layer4_outputs(706);
    outputs(7251) <= layer4_outputs(4274);
    outputs(7252) <= layer4_outputs(6115);
    outputs(7253) <= (layer4_outputs(4649)) xor (layer4_outputs(6207));
    outputs(7254) <= layer4_outputs(1605);
    outputs(7255) <= not((layer4_outputs(723)) xor (layer4_outputs(6240)));
    outputs(7256) <= (layer4_outputs(3560)) xor (layer4_outputs(3430));
    outputs(7257) <= (layer4_outputs(5742)) and (layer4_outputs(1164));
    outputs(7258) <= layer4_outputs(2246);
    outputs(7259) <= (layer4_outputs(5503)) and not (layer4_outputs(6072));
    outputs(7260) <= layer4_outputs(4095);
    outputs(7261) <= layer4_outputs(3224);
    outputs(7262) <= not(layer4_outputs(4852));
    outputs(7263) <= (layer4_outputs(3885)) and (layer4_outputs(2518));
    outputs(7264) <= layer4_outputs(4016);
    outputs(7265) <= not(layer4_outputs(5990));
    outputs(7266) <= not(layer4_outputs(4994));
    outputs(7267) <= not(layer4_outputs(4292));
    outputs(7268) <= layer4_outputs(4659);
    outputs(7269) <= (layer4_outputs(624)) or (layer4_outputs(6557));
    outputs(7270) <= not(layer4_outputs(2604));
    outputs(7271) <= not((layer4_outputs(7479)) xor (layer4_outputs(3545)));
    outputs(7272) <= layer4_outputs(3277);
    outputs(7273) <= layer4_outputs(3013);
    outputs(7274) <= (layer4_outputs(6727)) and not (layer4_outputs(4349));
    outputs(7275) <= layer4_outputs(4084);
    outputs(7276) <= layer4_outputs(975);
    outputs(7277) <= (layer4_outputs(4105)) xor (layer4_outputs(3746));
    outputs(7278) <= layer4_outputs(6058);
    outputs(7279) <= (layer4_outputs(919)) xor (layer4_outputs(7252));
    outputs(7280) <= layer4_outputs(1756);
    outputs(7281) <= (layer4_outputs(1994)) and not (layer4_outputs(5722));
    outputs(7282) <= (layer4_outputs(6938)) or (layer4_outputs(5746));
    outputs(7283) <= (layer4_outputs(1274)) or (layer4_outputs(7129));
    outputs(7284) <= not(layer4_outputs(471));
    outputs(7285) <= (layer4_outputs(2423)) and not (layer4_outputs(3004));
    outputs(7286) <= not(layer4_outputs(1775));
    outputs(7287) <= layer4_outputs(7138);
    outputs(7288) <= layer4_outputs(2780);
    outputs(7289) <= layer4_outputs(1505);
    outputs(7290) <= not((layer4_outputs(1122)) or (layer4_outputs(3827)));
    outputs(7291) <= not(layer4_outputs(5716));
    outputs(7292) <= not((layer4_outputs(7118)) or (layer4_outputs(1886)));
    outputs(7293) <= layer4_outputs(2982);
    outputs(7294) <= not(layer4_outputs(4118));
    outputs(7295) <= not(layer4_outputs(4354));
    outputs(7296) <= layer4_outputs(116);
    outputs(7297) <= not(layer4_outputs(5837));
    outputs(7298) <= layer4_outputs(2306);
    outputs(7299) <= (layer4_outputs(5334)) xor (layer4_outputs(3049));
    outputs(7300) <= (layer4_outputs(3525)) or (layer4_outputs(2902));
    outputs(7301) <= (layer4_outputs(236)) xor (layer4_outputs(5770));
    outputs(7302) <= not((layer4_outputs(3798)) or (layer4_outputs(1390)));
    outputs(7303) <= not(layer4_outputs(550));
    outputs(7304) <= layer4_outputs(104);
    outputs(7305) <= (layer4_outputs(4635)) and not (layer4_outputs(5400));
    outputs(7306) <= (layer4_outputs(6999)) xor (layer4_outputs(6270));
    outputs(7307) <= not(layer4_outputs(7232));
    outputs(7308) <= not(layer4_outputs(902));
    outputs(7309) <= not((layer4_outputs(3216)) xor (layer4_outputs(6292)));
    outputs(7310) <= layer4_outputs(5717);
    outputs(7311) <= not(layer4_outputs(6259));
    outputs(7312) <= not((layer4_outputs(7180)) xor (layer4_outputs(5481)));
    outputs(7313) <= (layer4_outputs(6082)) and not (layer4_outputs(1866));
    outputs(7314) <= (layer4_outputs(4046)) xor (layer4_outputs(1571));
    outputs(7315) <= (layer4_outputs(5506)) xor (layer4_outputs(1414));
    outputs(7316) <= (layer4_outputs(3780)) and (layer4_outputs(6047));
    outputs(7317) <= (layer4_outputs(1875)) and (layer4_outputs(6561));
    outputs(7318) <= layer4_outputs(6936);
    outputs(7319) <= not((layer4_outputs(6836)) xor (layer4_outputs(3736)));
    outputs(7320) <= not(layer4_outputs(4682));
    outputs(7321) <= not((layer4_outputs(1436)) or (layer4_outputs(1471)));
    outputs(7322) <= (layer4_outputs(6187)) and not (layer4_outputs(5217));
    outputs(7323) <= (layer4_outputs(6734)) xor (layer4_outputs(6377));
    outputs(7324) <= layer4_outputs(7068);
    outputs(7325) <= not((layer4_outputs(2718)) xor (layer4_outputs(5572)));
    outputs(7326) <= not(layer4_outputs(3010));
    outputs(7327) <= layer4_outputs(6585);
    outputs(7328) <= (layer4_outputs(4592)) and not (layer4_outputs(7160));
    outputs(7329) <= not((layer4_outputs(1955)) and (layer4_outputs(296)));
    outputs(7330) <= not(layer4_outputs(1538));
    outputs(7331) <= (layer4_outputs(3287)) and not (layer4_outputs(5191));
    outputs(7332) <= (layer4_outputs(1141)) and not (layer4_outputs(406));
    outputs(7333) <= layer4_outputs(5297);
    outputs(7334) <= layer4_outputs(4879);
    outputs(7335) <= not(layer4_outputs(5656));
    outputs(7336) <= (layer4_outputs(1917)) xor (layer4_outputs(1708));
    outputs(7337) <= (layer4_outputs(1043)) and not (layer4_outputs(1248));
    outputs(7338) <= (layer4_outputs(5904)) xor (layer4_outputs(249));
    outputs(7339) <= not((layer4_outputs(2916)) and (layer4_outputs(1528)));
    outputs(7340) <= layer4_outputs(4779);
    outputs(7341) <= not((layer4_outputs(5816)) xor (layer4_outputs(1444)));
    outputs(7342) <= not(layer4_outputs(6067)) or (layer4_outputs(1683));
    outputs(7343) <= layer4_outputs(2374);
    outputs(7344) <= not(layer4_outputs(6385));
    outputs(7345) <= layer4_outputs(942);
    outputs(7346) <= not(layer4_outputs(2496)) or (layer4_outputs(6654));
    outputs(7347) <= not((layer4_outputs(5747)) xor (layer4_outputs(2339)));
    outputs(7348) <= (layer4_outputs(5388)) xor (layer4_outputs(1581));
    outputs(7349) <= layer4_outputs(6720);
    outputs(7350) <= not(layer4_outputs(2244)) or (layer4_outputs(5746));
    outputs(7351) <= not(layer4_outputs(3555));
    outputs(7352) <= not(layer4_outputs(7206));
    outputs(7353) <= layer4_outputs(283);
    outputs(7354) <= not(layer4_outputs(4724));
    outputs(7355) <= layer4_outputs(649);
    outputs(7356) <= layer4_outputs(5645);
    outputs(7357) <= not((layer4_outputs(564)) or (layer4_outputs(1199)));
    outputs(7358) <= layer4_outputs(3594);
    outputs(7359) <= not(layer4_outputs(731));
    outputs(7360) <= (layer4_outputs(2354)) xor (layer4_outputs(1036));
    outputs(7361) <= layer4_outputs(144);
    outputs(7362) <= not(layer4_outputs(3143));
    outputs(7363) <= layer4_outputs(7478);
    outputs(7364) <= not(layer4_outputs(5462));
    outputs(7365) <= (layer4_outputs(572)) xor (layer4_outputs(4407));
    outputs(7366) <= not((layer4_outputs(760)) xor (layer4_outputs(6944)));
    outputs(7367) <= (layer4_outputs(374)) xor (layer4_outputs(3250));
    outputs(7368) <= layer4_outputs(7429);
    outputs(7369) <= (layer4_outputs(4005)) and (layer4_outputs(1647));
    outputs(7370) <= (layer4_outputs(4743)) and (layer4_outputs(1200));
    outputs(7371) <= (layer4_outputs(3000)) xor (layer4_outputs(6949));
    outputs(7372) <= not((layer4_outputs(6001)) xor (layer4_outputs(1593)));
    outputs(7373) <= not((layer4_outputs(769)) or (layer4_outputs(4379)));
    outputs(7374) <= (layer4_outputs(1819)) xor (layer4_outputs(4592));
    outputs(7375) <= layer4_outputs(6477);
    outputs(7376) <= not(layer4_outputs(4221));
    outputs(7377) <= (layer4_outputs(46)) xor (layer4_outputs(7471));
    outputs(7378) <= (layer4_outputs(961)) and not (layer4_outputs(6484));
    outputs(7379) <= not(layer4_outputs(6246));
    outputs(7380) <= not(layer4_outputs(5267));
    outputs(7381) <= layer4_outputs(7604);
    outputs(7382) <= not(layer4_outputs(4064));
    outputs(7383) <= layer4_outputs(5211);
    outputs(7384) <= (layer4_outputs(5344)) and (layer4_outputs(5052));
    outputs(7385) <= not(layer4_outputs(6036));
    outputs(7386) <= (layer4_outputs(1058)) and (layer4_outputs(253));
    outputs(7387) <= not(layer4_outputs(5918));
    outputs(7388) <= not((layer4_outputs(2739)) or (layer4_outputs(4469)));
    outputs(7389) <= layer4_outputs(2505);
    outputs(7390) <= not(layer4_outputs(2009));
    outputs(7391) <= not((layer4_outputs(3561)) or (layer4_outputs(1290)));
    outputs(7392) <= layer4_outputs(5160);
    outputs(7393) <= not(layer4_outputs(6724));
    outputs(7394) <= not(layer4_outputs(7373));
    outputs(7395) <= (layer4_outputs(3084)) and not (layer4_outputs(3661));
    outputs(7396) <= layer4_outputs(1272);
    outputs(7397) <= (layer4_outputs(6120)) and (layer4_outputs(549));
    outputs(7398) <= not(layer4_outputs(5789));
    outputs(7399) <= layer4_outputs(3330);
    outputs(7400) <= not(layer4_outputs(2773));
    outputs(7401) <= (layer4_outputs(3866)) xor (layer4_outputs(5595));
    outputs(7402) <= layer4_outputs(3605);
    outputs(7403) <= not((layer4_outputs(2987)) and (layer4_outputs(932)));
    outputs(7404) <= (layer4_outputs(4334)) and not (layer4_outputs(5349));
    outputs(7405) <= not((layer4_outputs(5196)) and (layer4_outputs(7390)));
    outputs(7406) <= not(layer4_outputs(1810));
    outputs(7407) <= layer4_outputs(694);
    outputs(7408) <= layer4_outputs(1514);
    outputs(7409) <= not(layer4_outputs(4627));
    outputs(7410) <= layer4_outputs(3613);
    outputs(7411) <= (layer4_outputs(282)) and (layer4_outputs(3250));
    outputs(7412) <= not(layer4_outputs(1135));
    outputs(7413) <= not(layer4_outputs(3670));
    outputs(7414) <= not(layer4_outputs(835));
    outputs(7415) <= not(layer4_outputs(778)) or (layer4_outputs(4268));
    outputs(7416) <= layer4_outputs(7580);
    outputs(7417) <= not(layer4_outputs(7022));
    outputs(7418) <= layer4_outputs(5937);
    outputs(7419) <= (layer4_outputs(4595)) xor (layer4_outputs(7005));
    outputs(7420) <= (layer4_outputs(813)) xor (layer4_outputs(7406));
    outputs(7421) <= not((layer4_outputs(7507)) xor (layer4_outputs(3892)));
    outputs(7422) <= not(layer4_outputs(3710));
    outputs(7423) <= layer4_outputs(125);
    outputs(7424) <= not(layer4_outputs(897));
    outputs(7425) <= (layer4_outputs(1548)) and (layer4_outputs(5859));
    outputs(7426) <= layer4_outputs(5566);
    outputs(7427) <= layer4_outputs(208);
    outputs(7428) <= not((layer4_outputs(4858)) xor (layer4_outputs(5963)));
    outputs(7429) <= layer4_outputs(7549);
    outputs(7430) <= layer4_outputs(4695);
    outputs(7431) <= layer4_outputs(1139);
    outputs(7432) <= not(layer4_outputs(281));
    outputs(7433) <= not(layer4_outputs(4227));
    outputs(7434) <= layer4_outputs(7138);
    outputs(7435) <= not((layer4_outputs(4438)) xor (layer4_outputs(1641)));
    outputs(7436) <= layer4_outputs(1145);
    outputs(7437) <= layer4_outputs(989);
    outputs(7438) <= (layer4_outputs(1064)) and (layer4_outputs(3984));
    outputs(7439) <= layer4_outputs(3490);
    outputs(7440) <= not(layer4_outputs(2695)) or (layer4_outputs(3846));
    outputs(7441) <= layer4_outputs(6173);
    outputs(7442) <= (layer4_outputs(1287)) xor (layer4_outputs(5883));
    outputs(7443) <= layer4_outputs(774);
    outputs(7444) <= not(layer4_outputs(412));
    outputs(7445) <= (layer4_outputs(6580)) xor (layer4_outputs(6986));
    outputs(7446) <= layer4_outputs(1003);
    outputs(7447) <= not(layer4_outputs(5682));
    outputs(7448) <= (layer4_outputs(4594)) and not (layer4_outputs(5687));
    outputs(7449) <= not(layer4_outputs(5042));
    outputs(7450) <= (layer4_outputs(728)) xor (layer4_outputs(7605));
    outputs(7451) <= not(layer4_outputs(4985));
    outputs(7452) <= layer4_outputs(1350);
    outputs(7453) <= not((layer4_outputs(5389)) xor (layer4_outputs(4389)));
    outputs(7454) <= (layer4_outputs(5650)) and not (layer4_outputs(7084));
    outputs(7455) <= (layer4_outputs(2197)) xor (layer4_outputs(6090));
    outputs(7456) <= not(layer4_outputs(1763));
    outputs(7457) <= (layer4_outputs(2608)) xor (layer4_outputs(17));
    outputs(7458) <= not((layer4_outputs(279)) xor (layer4_outputs(7076)));
    outputs(7459) <= (layer4_outputs(315)) xor (layer4_outputs(3349));
    outputs(7460) <= not((layer4_outputs(6833)) or (layer4_outputs(7344)));
    outputs(7461) <= layer4_outputs(90);
    outputs(7462) <= layer4_outputs(2189);
    outputs(7463) <= (layer4_outputs(42)) xor (layer4_outputs(935));
    outputs(7464) <= layer4_outputs(2505);
    outputs(7465) <= layer4_outputs(3447);
    outputs(7466) <= not(layer4_outputs(4272));
    outputs(7467) <= (layer4_outputs(3523)) xor (layer4_outputs(3536));
    outputs(7468) <= (layer4_outputs(981)) xor (layer4_outputs(4150));
    outputs(7469) <= not(layer4_outputs(2710)) or (layer4_outputs(38));
    outputs(7470) <= layer4_outputs(1988);
    outputs(7471) <= not((layer4_outputs(1280)) xor (layer4_outputs(3087)));
    outputs(7472) <= not(layer4_outputs(7344));
    outputs(7473) <= not(layer4_outputs(1728));
    outputs(7474) <= not(layer4_outputs(802));
    outputs(7475) <= not(layer4_outputs(5072));
    outputs(7476) <= (layer4_outputs(7383)) and (layer4_outputs(62));
    outputs(7477) <= layer4_outputs(4490);
    outputs(7478) <= not(layer4_outputs(6238));
    outputs(7479) <= not(layer4_outputs(3272));
    outputs(7480) <= layer4_outputs(7098);
    outputs(7481) <= not(layer4_outputs(6840)) or (layer4_outputs(3929));
    outputs(7482) <= layer4_outputs(768);
    outputs(7483) <= not(layer4_outputs(2497));
    outputs(7484) <= layer4_outputs(1475);
    outputs(7485) <= layer4_outputs(2849);
    outputs(7486) <= (layer4_outputs(3621)) or (layer4_outputs(7578));
    outputs(7487) <= (layer4_outputs(2790)) and (layer4_outputs(5307));
    outputs(7488) <= not(layer4_outputs(3821));
    outputs(7489) <= layer4_outputs(6135);
    outputs(7490) <= layer4_outputs(1254);
    outputs(7491) <= not(layer4_outputs(7315));
    outputs(7492) <= layer4_outputs(6830);
    outputs(7493) <= (layer4_outputs(75)) xor (layer4_outputs(1816));
    outputs(7494) <= not(layer4_outputs(5614));
    outputs(7495) <= not(layer4_outputs(523));
    outputs(7496) <= (layer4_outputs(1426)) or (layer4_outputs(1736));
    outputs(7497) <= (layer4_outputs(187)) or (layer4_outputs(5846));
    outputs(7498) <= not(layer4_outputs(7181));
    outputs(7499) <= (layer4_outputs(7599)) and not (layer4_outputs(921));
    outputs(7500) <= (layer4_outputs(4011)) and not (layer4_outputs(5740));
    outputs(7501) <= not((layer4_outputs(5883)) xor (layer4_outputs(4615)));
    outputs(7502) <= not(layer4_outputs(6235));
    outputs(7503) <= (layer4_outputs(716)) and not (layer4_outputs(2438));
    outputs(7504) <= layer4_outputs(2596);
    outputs(7505) <= layer4_outputs(5627);
    outputs(7506) <= (layer4_outputs(584)) and (layer4_outputs(5887));
    outputs(7507) <= (layer4_outputs(1934)) and not (layer4_outputs(2685));
    outputs(7508) <= (layer4_outputs(924)) xor (layer4_outputs(4506));
    outputs(7509) <= layer4_outputs(4454);
    outputs(7510) <= layer4_outputs(2138);
    outputs(7511) <= not(layer4_outputs(2574));
    outputs(7512) <= not((layer4_outputs(1329)) or (layer4_outputs(6206)));
    outputs(7513) <= not(layer4_outputs(6409));
    outputs(7514) <= (layer4_outputs(179)) and not (layer4_outputs(5862));
    outputs(7515) <= (layer4_outputs(4650)) xor (layer4_outputs(3085));
    outputs(7516) <= not((layer4_outputs(4327)) or (layer4_outputs(2065)));
    outputs(7517) <= not(layer4_outputs(6847));
    outputs(7518) <= layer4_outputs(284);
    outputs(7519) <= (layer4_outputs(2304)) and not (layer4_outputs(5572));
    outputs(7520) <= layer4_outputs(2510);
    outputs(7521) <= not((layer4_outputs(6579)) xor (layer4_outputs(6743)));
    outputs(7522) <= layer4_outputs(7147);
    outputs(7523) <= not((layer4_outputs(3598)) xor (layer4_outputs(2899)));
    outputs(7524) <= not(layer4_outputs(7329)) or (layer4_outputs(4076));
    outputs(7525) <= layer4_outputs(6670);
    outputs(7526) <= not(layer4_outputs(6369));
    outputs(7527) <= layer4_outputs(967);
    outputs(7528) <= not(layer4_outputs(1839));
    outputs(7529) <= layer4_outputs(2099);
    outputs(7530) <= not(layer4_outputs(7606));
    outputs(7531) <= layer4_outputs(7229);
    outputs(7532) <= not(layer4_outputs(1735));
    outputs(7533) <= layer4_outputs(585);
    outputs(7534) <= layer4_outputs(6711);
    outputs(7535) <= layer4_outputs(3998);
    outputs(7536) <= not(layer4_outputs(3070));
    outputs(7537) <= not(layer4_outputs(2987));
    outputs(7538) <= not((layer4_outputs(1566)) or (layer4_outputs(5118)));
    outputs(7539) <= (layer4_outputs(1450)) and (layer4_outputs(561));
    outputs(7540) <= layer4_outputs(4329);
    outputs(7541) <= layer4_outputs(13);
    outputs(7542) <= not(layer4_outputs(1440));
    outputs(7543) <= layer4_outputs(6456);
    outputs(7544) <= not((layer4_outputs(4500)) or (layer4_outputs(7323)));
    outputs(7545) <= layer4_outputs(6629);
    outputs(7546) <= not(layer4_outputs(7646)) or (layer4_outputs(3273));
    outputs(7547) <= not(layer4_outputs(664));
    outputs(7548) <= (layer4_outputs(7610)) or (layer4_outputs(1711));
    outputs(7549) <= not((layer4_outputs(3021)) xor (layer4_outputs(4628)));
    outputs(7550) <= layer4_outputs(7374);
    outputs(7551) <= not(layer4_outputs(4791));
    outputs(7552) <= layer4_outputs(7239);
    outputs(7553) <= not(layer4_outputs(3114));
    outputs(7554) <= not(layer4_outputs(6384));
    outputs(7555) <= (layer4_outputs(2735)) and (layer4_outputs(1221));
    outputs(7556) <= not(layer4_outputs(2031));
    outputs(7557) <= (layer4_outputs(393)) xor (layer4_outputs(5976));
    outputs(7558) <= layer4_outputs(1317);
    outputs(7559) <= layer4_outputs(3059);
    outputs(7560) <= layer4_outputs(2401);
    outputs(7561) <= not((layer4_outputs(5506)) or (layer4_outputs(3552)));
    outputs(7562) <= not(layer4_outputs(829));
    outputs(7563) <= not(layer4_outputs(3938));
    outputs(7564) <= layer4_outputs(3962);
    outputs(7565) <= not(layer4_outputs(805));
    outputs(7566) <= layer4_outputs(2467);
    outputs(7567) <= (layer4_outputs(7013)) and not (layer4_outputs(4907));
    outputs(7568) <= not(layer4_outputs(5856));
    outputs(7569) <= not((layer4_outputs(2167)) xor (layer4_outputs(3486)));
    outputs(7570) <= not((layer4_outputs(5835)) or (layer4_outputs(7459)));
    outputs(7571) <= layer4_outputs(5015);
    outputs(7572) <= layer4_outputs(4603);
    outputs(7573) <= layer4_outputs(6341);
    outputs(7574) <= layer4_outputs(4282);
    outputs(7575) <= not(layer4_outputs(6086));
    outputs(7576) <= (layer4_outputs(3558)) or (layer4_outputs(5406));
    outputs(7577) <= layer4_outputs(6975);
    outputs(7578) <= not(layer4_outputs(2430));
    outputs(7579) <= layer4_outputs(7168);
    outputs(7580) <= not((layer4_outputs(6504)) xor (layer4_outputs(6581)));
    outputs(7581) <= not((layer4_outputs(7136)) xor (layer4_outputs(5817)));
    outputs(7582) <= not(layer4_outputs(6069));
    outputs(7583) <= not(layer4_outputs(2495));
    outputs(7584) <= layer4_outputs(4965);
    outputs(7585) <= layer4_outputs(1192);
    outputs(7586) <= layer4_outputs(4936);
    outputs(7587) <= not(layer4_outputs(315));
    outputs(7588) <= not(layer4_outputs(7165));
    outputs(7589) <= layer4_outputs(3796);
    outputs(7590) <= not((layer4_outputs(5514)) or (layer4_outputs(2975)));
    outputs(7591) <= not(layer4_outputs(4655));
    outputs(7592) <= not(layer4_outputs(4631));
    outputs(7593) <= layer4_outputs(2941);
    outputs(7594) <= not(layer4_outputs(4377));
    outputs(7595) <= layer4_outputs(5526);
    outputs(7596) <= not((layer4_outputs(6342)) xor (layer4_outputs(7401)));
    outputs(7597) <= (layer4_outputs(4033)) and not (layer4_outputs(5873));
    outputs(7598) <= (layer4_outputs(4376)) and not (layer4_outputs(1447));
    outputs(7599) <= layer4_outputs(5445);
    outputs(7600) <= not((layer4_outputs(5088)) xor (layer4_outputs(1096)));
    outputs(7601) <= not(layer4_outputs(742));
    outputs(7602) <= not(layer4_outputs(2452));
    outputs(7603) <= not(layer4_outputs(7281));
    outputs(7604) <= not(layer4_outputs(4057));
    outputs(7605) <= not(layer4_outputs(3178)) or (layer4_outputs(1180));
    outputs(7606) <= (layer4_outputs(5989)) xor (layer4_outputs(2005));
    outputs(7607) <= layer4_outputs(3751);
    outputs(7608) <= not(layer4_outputs(1285));
    outputs(7609) <= not((layer4_outputs(5997)) or (layer4_outputs(1246)));
    outputs(7610) <= not(layer4_outputs(2685));
    outputs(7611) <= not(layer4_outputs(5766));
    outputs(7612) <= not((layer4_outputs(510)) or (layer4_outputs(4851)));
    outputs(7613) <= (layer4_outputs(4116)) and (layer4_outputs(3053));
    outputs(7614) <= not(layer4_outputs(3292));
    outputs(7615) <= layer4_outputs(5116);
    outputs(7616) <= not(layer4_outputs(3100)) or (layer4_outputs(1989));
    outputs(7617) <= (layer4_outputs(2899)) or (layer4_outputs(1743));
    outputs(7618) <= (layer4_outputs(1089)) xor (layer4_outputs(800));
    outputs(7619) <= not(layer4_outputs(5201));
    outputs(7620) <= not(layer4_outputs(896));
    outputs(7621) <= layer4_outputs(3148);
    outputs(7622) <= not(layer4_outputs(7022));
    outputs(7623) <= not(layer4_outputs(2839));
    outputs(7624) <= not(layer4_outputs(2234)) or (layer4_outputs(5637));
    outputs(7625) <= not(layer4_outputs(7586));
    outputs(7626) <= not(layer4_outputs(5260));
    outputs(7627) <= not(layer4_outputs(4688));
    outputs(7628) <= not((layer4_outputs(5867)) or (layer4_outputs(71)));
    outputs(7629) <= layer4_outputs(3717);
    outputs(7630) <= (layer4_outputs(5420)) and (layer4_outputs(4887));
    outputs(7631) <= not((layer4_outputs(5825)) and (layer4_outputs(3108)));
    outputs(7632) <= not(layer4_outputs(7427));
    outputs(7633) <= (layer4_outputs(2369)) xor (layer4_outputs(1689));
    outputs(7634) <= (layer4_outputs(5651)) and (layer4_outputs(5774));
    outputs(7635) <= not((layer4_outputs(4680)) xor (layer4_outputs(3766)));
    outputs(7636) <= not((layer4_outputs(1679)) and (layer4_outputs(98)));
    outputs(7637) <= (layer4_outputs(4830)) and (layer4_outputs(2450));
    outputs(7638) <= not((layer4_outputs(6158)) xor (layer4_outputs(4031)));
    outputs(7639) <= not((layer4_outputs(5606)) xor (layer4_outputs(1086)));
    outputs(7640) <= not(layer4_outputs(4752));
    outputs(7641) <= not(layer4_outputs(4422));
    outputs(7642) <= not(layer4_outputs(6250));
    outputs(7643) <= (layer4_outputs(1782)) xor (layer4_outputs(4330));
    outputs(7644) <= not(layer4_outputs(5682));
    outputs(7645) <= not(layer4_outputs(6297));
    outputs(7646) <= not((layer4_outputs(6667)) xor (layer4_outputs(4828)));
    outputs(7647) <= not(layer4_outputs(3357));
    outputs(7648) <= not((layer4_outputs(950)) xor (layer4_outputs(3717)));
    outputs(7649) <= (layer4_outputs(4289)) xor (layer4_outputs(3518));
    outputs(7650) <= layer4_outputs(2699);
    outputs(7651) <= not(layer4_outputs(4422));
    outputs(7652) <= not(layer4_outputs(1217));
    outputs(7653) <= (layer4_outputs(7043)) xor (layer4_outputs(4389));
    outputs(7654) <= not(layer4_outputs(2962));
    outputs(7655) <= not(layer4_outputs(2934));
    outputs(7656) <= not(layer4_outputs(348));
    outputs(7657) <= not(layer4_outputs(595)) or (layer4_outputs(1432));
    outputs(7658) <= layer4_outputs(1740);
    outputs(7659) <= layer4_outputs(2677);
    outputs(7660) <= not(layer4_outputs(2735)) or (layer4_outputs(6068));
    outputs(7661) <= not(layer4_outputs(69));
    outputs(7662) <= not(layer4_outputs(244));
    outputs(7663) <= layer4_outputs(160);
    outputs(7664) <= layer4_outputs(4311);
    outputs(7665) <= layer4_outputs(4565);
    outputs(7666) <= layer4_outputs(4234);
    outputs(7667) <= (layer4_outputs(2575)) xor (layer4_outputs(941));
    outputs(7668) <= layer4_outputs(7546);
    outputs(7669) <= layer4_outputs(2095);
    outputs(7670) <= layer4_outputs(1029);
    outputs(7671) <= not(layer4_outputs(5251));
    outputs(7672) <= (layer4_outputs(1716)) and not (layer4_outputs(6399));
    outputs(7673) <= layer4_outputs(6429);
    outputs(7674) <= layer4_outputs(6798);
    outputs(7675) <= (layer4_outputs(2620)) and not (layer4_outputs(1409));
    outputs(7676) <= not((layer4_outputs(3817)) xor (layer4_outputs(3576)));
    outputs(7677) <= layer4_outputs(7656);
    outputs(7678) <= (layer4_outputs(4748)) xor (layer4_outputs(4615));
    outputs(7679) <= not((layer4_outputs(6751)) xor (layer4_outputs(6349)));

end Behavioral;
