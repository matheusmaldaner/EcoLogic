library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(2559 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(2559 downto 0);
    signal layer1_outputs : std_logic_vector(2559 downto 0);
    signal layer2_outputs : std_logic_vector(2559 downto 0);
    signal layer3_outputs : std_logic_vector(2559 downto 0);
    signal layer4_outputs : std_logic_vector(2559 downto 0);
    signal layer5_outputs : std_logic_vector(2559 downto 0);
    signal layer6_outputs : std_logic_vector(2559 downto 0);

begin

    layer0_outputs(0) <= not(inputs(166)) or (inputs(45));
    layer0_outputs(1) <= '0';
    layer0_outputs(2) <= not(inputs(226));
    layer0_outputs(3) <= not(inputs(152));
    layer0_outputs(4) <= '0';
    layer0_outputs(5) <= not(inputs(87)) or (inputs(164));
    layer0_outputs(6) <= '0';
    layer0_outputs(7) <= not((inputs(34)) or (inputs(26)));
    layer0_outputs(8) <= not(inputs(250));
    layer0_outputs(9) <= inputs(2);
    layer0_outputs(10) <= not((inputs(81)) and (inputs(252)));
    layer0_outputs(11) <= '0';
    layer0_outputs(12) <= not(inputs(92)) or (inputs(142));
    layer0_outputs(13) <= not(inputs(18));
    layer0_outputs(14) <= inputs(104);
    layer0_outputs(15) <= not((inputs(56)) or (inputs(215)));
    layer0_outputs(16) <= not(inputs(114));
    layer0_outputs(17) <= inputs(82);
    layer0_outputs(18) <= (inputs(122)) and not (inputs(186));
    layer0_outputs(19) <= not(inputs(150)) or (inputs(26));
    layer0_outputs(20) <= not((inputs(188)) or (inputs(144)));
    layer0_outputs(21) <= '0';
    layer0_outputs(22) <= not((inputs(207)) and (inputs(65)));
    layer0_outputs(23) <= not(inputs(189));
    layer0_outputs(24) <= (inputs(251)) or (inputs(89));
    layer0_outputs(25) <= '0';
    layer0_outputs(26) <= (inputs(235)) xor (inputs(220));
    layer0_outputs(27) <= '0';
    layer0_outputs(28) <= inputs(75);
    layer0_outputs(29) <= inputs(161);
    layer0_outputs(30) <= (inputs(69)) or (inputs(22));
    layer0_outputs(31) <= not((inputs(224)) xor (inputs(76)));
    layer0_outputs(32) <= '1';
    layer0_outputs(33) <= inputs(148);
    layer0_outputs(34) <= inputs(74);
    layer0_outputs(35) <= not(inputs(171));
    layer0_outputs(36) <= '0';
    layer0_outputs(37) <= (inputs(100)) and (inputs(224));
    layer0_outputs(38) <= not((inputs(171)) or (inputs(101)));
    layer0_outputs(39) <= not((inputs(128)) or (inputs(248)));
    layer0_outputs(40) <= '0';
    layer0_outputs(41) <= (inputs(192)) and not (inputs(13));
    layer0_outputs(42) <= (inputs(91)) or (inputs(50));
    layer0_outputs(43) <= inputs(197);
    layer0_outputs(44) <= (inputs(9)) and not (inputs(27));
    layer0_outputs(45) <= not(inputs(71));
    layer0_outputs(46) <= inputs(189);
    layer0_outputs(47) <= not(inputs(220));
    layer0_outputs(48) <= inputs(189);
    layer0_outputs(49) <= inputs(151);
    layer0_outputs(50) <= '1';
    layer0_outputs(51) <= not((inputs(49)) and (inputs(153)));
    layer0_outputs(52) <= inputs(144);
    layer0_outputs(53) <= inputs(241);
    layer0_outputs(54) <= not(inputs(135));
    layer0_outputs(55) <= (inputs(156)) and not (inputs(196));
    layer0_outputs(56) <= not(inputs(99));
    layer0_outputs(57) <= not(inputs(161));
    layer0_outputs(58) <= not((inputs(0)) or (inputs(56)));
    layer0_outputs(59) <= not(inputs(4)) or (inputs(249));
    layer0_outputs(60) <= inputs(175);
    layer0_outputs(61) <= '1';
    layer0_outputs(62) <= '1';
    layer0_outputs(63) <= not(inputs(136));
    layer0_outputs(64) <= not((inputs(89)) and (inputs(22)));
    layer0_outputs(65) <= (inputs(196)) or (inputs(113));
    layer0_outputs(66) <= not((inputs(25)) or (inputs(94)));
    layer0_outputs(67) <= inputs(5);
    layer0_outputs(68) <= not((inputs(218)) or (inputs(190)));
    layer0_outputs(69) <= not(inputs(138)) or (inputs(150));
    layer0_outputs(70) <= (inputs(186)) and (inputs(250));
    layer0_outputs(71) <= not(inputs(6)) or (inputs(77));
    layer0_outputs(72) <= (inputs(189)) or (inputs(108));
    layer0_outputs(73) <= (inputs(4)) or (inputs(190));
    layer0_outputs(74) <= not((inputs(5)) and (inputs(26)));
    layer0_outputs(75) <= not(inputs(252)) or (inputs(11));
    layer0_outputs(76) <= not(inputs(235));
    layer0_outputs(77) <= inputs(46);
    layer0_outputs(78) <= inputs(34);
    layer0_outputs(79) <= (inputs(121)) and not (inputs(90));
    layer0_outputs(80) <= '0';
    layer0_outputs(81) <= (inputs(178)) or (inputs(50));
    layer0_outputs(82) <= not(inputs(107));
    layer0_outputs(83) <= inputs(26);
    layer0_outputs(84) <= '0';
    layer0_outputs(85) <= '0';
    layer0_outputs(86) <= not((inputs(12)) xor (inputs(6)));
    layer0_outputs(87) <= not(inputs(12));
    layer0_outputs(88) <= not(inputs(146));
    layer0_outputs(89) <= '0';
    layer0_outputs(90) <= inputs(44);
    layer0_outputs(91) <= not(inputs(84));
    layer0_outputs(92) <= '1';
    layer0_outputs(93) <= '1';
    layer0_outputs(94) <= not((inputs(220)) and (inputs(139)));
    layer0_outputs(95) <= inputs(230);
    layer0_outputs(96) <= not(inputs(197)) or (inputs(12));
    layer0_outputs(97) <= (inputs(117)) and not (inputs(13));
    layer0_outputs(98) <= not((inputs(169)) or (inputs(54)));
    layer0_outputs(99) <= not(inputs(134)) or (inputs(17));
    layer0_outputs(100) <= not((inputs(2)) or (inputs(187)));
    layer0_outputs(101) <= '1';
    layer0_outputs(102) <= '1';
    layer0_outputs(103) <= inputs(230);
    layer0_outputs(104) <= '1';
    layer0_outputs(105) <= inputs(85);
    layer0_outputs(106) <= not(inputs(102)) or (inputs(154));
    layer0_outputs(107) <= inputs(68);
    layer0_outputs(108) <= (inputs(198)) or (inputs(214));
    layer0_outputs(109) <= not(inputs(210));
    layer0_outputs(110) <= not((inputs(246)) or (inputs(100)));
    layer0_outputs(111) <= not(inputs(165));
    layer0_outputs(112) <= '0';
    layer0_outputs(113) <= not(inputs(82)) or (inputs(36));
    layer0_outputs(114) <= (inputs(252)) or (inputs(238));
    layer0_outputs(115) <= not(inputs(246));
    layer0_outputs(116) <= (inputs(174)) and not (inputs(70));
    layer0_outputs(117) <= (inputs(82)) or (inputs(238));
    layer0_outputs(118) <= not((inputs(90)) or (inputs(166)));
    layer0_outputs(119) <= inputs(143);
    layer0_outputs(120) <= '1';
    layer0_outputs(121) <= '1';
    layer0_outputs(122) <= (inputs(224)) or (inputs(246));
    layer0_outputs(123) <= (inputs(156)) or (inputs(10));
    layer0_outputs(124) <= not((inputs(126)) or (inputs(248)));
    layer0_outputs(125) <= inputs(174);
    layer0_outputs(126) <= not(inputs(91));
    layer0_outputs(127) <= not(inputs(145)) or (inputs(195));
    layer0_outputs(128) <= not(inputs(39));
    layer0_outputs(129) <= not(inputs(119)) or (inputs(107));
    layer0_outputs(130) <= (inputs(41)) and (inputs(125));
    layer0_outputs(131) <= inputs(100);
    layer0_outputs(132) <= '0';
    layer0_outputs(133) <= '0';
    layer0_outputs(134) <= (inputs(101)) and not (inputs(121));
    layer0_outputs(135) <= inputs(230);
    layer0_outputs(136) <= (inputs(102)) and (inputs(85));
    layer0_outputs(137) <= '1';
    layer0_outputs(138) <= (inputs(41)) or (inputs(5));
    layer0_outputs(139) <= inputs(93);
    layer0_outputs(140) <= inputs(14);
    layer0_outputs(141) <= (inputs(223)) xor (inputs(193));
    layer0_outputs(142) <= not((inputs(120)) xor (inputs(167)));
    layer0_outputs(143) <= (inputs(227)) and not (inputs(253));
    layer0_outputs(144) <= not(inputs(27)) or (inputs(152));
    layer0_outputs(145) <= (inputs(93)) and not (inputs(36));
    layer0_outputs(146) <= (inputs(198)) or (inputs(129));
    layer0_outputs(147) <= '0';
    layer0_outputs(148) <= '1';
    layer0_outputs(149) <= not((inputs(23)) and (inputs(10)));
    layer0_outputs(150) <= not((inputs(7)) and (inputs(118)));
    layer0_outputs(151) <= not(inputs(31));
    layer0_outputs(152) <= '0';
    layer0_outputs(153) <= (inputs(64)) and not (inputs(157));
    layer0_outputs(154) <= not((inputs(209)) or (inputs(2)));
    layer0_outputs(155) <= '0';
    layer0_outputs(156) <= not((inputs(28)) or (inputs(125)));
    layer0_outputs(157) <= (inputs(186)) or (inputs(77));
    layer0_outputs(158) <= (inputs(160)) or (inputs(129));
    layer0_outputs(159) <= '1';
    layer0_outputs(160) <= (inputs(75)) and not (inputs(224));
    layer0_outputs(161) <= not((inputs(42)) or (inputs(50)));
    layer0_outputs(162) <= inputs(19);
    layer0_outputs(163) <= inputs(116);
    layer0_outputs(164) <= (inputs(135)) and not (inputs(244));
    layer0_outputs(165) <= not((inputs(207)) or (inputs(241)));
    layer0_outputs(166) <= (inputs(0)) or (inputs(58));
    layer0_outputs(167) <= inputs(21);
    layer0_outputs(168) <= (inputs(111)) and (inputs(9));
    layer0_outputs(169) <= not(inputs(22));
    layer0_outputs(170) <= (inputs(188)) and not (inputs(48));
    layer0_outputs(171) <= inputs(41);
    layer0_outputs(172) <= not(inputs(231));
    layer0_outputs(173) <= (inputs(143)) and not (inputs(93));
    layer0_outputs(174) <= not(inputs(38));
    layer0_outputs(175) <= (inputs(88)) and (inputs(131));
    layer0_outputs(176) <= (inputs(28)) and (inputs(22));
    layer0_outputs(177) <= '1';
    layer0_outputs(178) <= (inputs(94)) or (inputs(108));
    layer0_outputs(179) <= not((inputs(93)) and (inputs(129)));
    layer0_outputs(180) <= '1';
    layer0_outputs(181) <= '0';
    layer0_outputs(182) <= not(inputs(92)) or (inputs(189));
    layer0_outputs(183) <= not(inputs(203));
    layer0_outputs(184) <= inputs(157);
    layer0_outputs(185) <= inputs(163);
    layer0_outputs(186) <= inputs(141);
    layer0_outputs(187) <= '0';
    layer0_outputs(188) <= '0';
    layer0_outputs(189) <= not((inputs(227)) or (inputs(37)));
    layer0_outputs(190) <= not(inputs(208)) or (inputs(66));
    layer0_outputs(191) <= not((inputs(76)) and (inputs(241)));
    layer0_outputs(192) <= not(inputs(101));
    layer0_outputs(193) <= not(inputs(4)) or (inputs(217));
    layer0_outputs(194) <= not((inputs(192)) or (inputs(33)));
    layer0_outputs(195) <= not(inputs(61));
    layer0_outputs(196) <= inputs(129);
    layer0_outputs(197) <= not(inputs(161));
    layer0_outputs(198) <= inputs(121);
    layer0_outputs(199) <= inputs(46);
    layer0_outputs(200) <= (inputs(123)) and not (inputs(41));
    layer0_outputs(201) <= not(inputs(29)) or (inputs(178));
    layer0_outputs(202) <= not(inputs(158));
    layer0_outputs(203) <= (inputs(7)) and (inputs(16));
    layer0_outputs(204) <= not(inputs(162));
    layer0_outputs(205) <= '0';
    layer0_outputs(206) <= inputs(226);
    layer0_outputs(207) <= not(inputs(234));
    layer0_outputs(208) <= not(inputs(26)) or (inputs(26));
    layer0_outputs(209) <= inputs(102);
    layer0_outputs(210) <= inputs(189);
    layer0_outputs(211) <= (inputs(71)) or (inputs(245));
    layer0_outputs(212) <= not((inputs(76)) or (inputs(165)));
    layer0_outputs(213) <= not((inputs(81)) and (inputs(228)));
    layer0_outputs(214) <= inputs(239);
    layer0_outputs(215) <= '0';
    layer0_outputs(216) <= not(inputs(255));
    layer0_outputs(217) <= inputs(229);
    layer0_outputs(218) <= '1';
    layer0_outputs(219) <= '1';
    layer0_outputs(220) <= not(inputs(23));
    layer0_outputs(221) <= (inputs(21)) and not (inputs(64));
    layer0_outputs(222) <= '1';
    layer0_outputs(223) <= inputs(191);
    layer0_outputs(224) <= (inputs(61)) and not (inputs(71));
    layer0_outputs(225) <= not(inputs(37)) or (inputs(0));
    layer0_outputs(226) <= '0';
    layer0_outputs(227) <= '0';
    layer0_outputs(228) <= not((inputs(74)) and (inputs(174)));
    layer0_outputs(229) <= not((inputs(70)) and (inputs(90)));
    layer0_outputs(230) <= not((inputs(166)) and (inputs(74)));
    layer0_outputs(231) <= '1';
    layer0_outputs(232) <= inputs(109);
    layer0_outputs(233) <= '0';
    layer0_outputs(234) <= (inputs(8)) or (inputs(94));
    layer0_outputs(235) <= '0';
    layer0_outputs(236) <= '1';
    layer0_outputs(237) <= (inputs(204)) and not (inputs(109));
    layer0_outputs(238) <= not(inputs(184));
    layer0_outputs(239) <= not(inputs(229));
    layer0_outputs(240) <= not(inputs(40)) or (inputs(221));
    layer0_outputs(241) <= not(inputs(76));
    layer0_outputs(242) <= inputs(90);
    layer0_outputs(243) <= inputs(247);
    layer0_outputs(244) <= not(inputs(96));
    layer0_outputs(245) <= not((inputs(107)) or (inputs(252)));
    layer0_outputs(246) <= not(inputs(180));
    layer0_outputs(247) <= (inputs(28)) or (inputs(52));
    layer0_outputs(248) <= not(inputs(231));
    layer0_outputs(249) <= '1';
    layer0_outputs(250) <= not((inputs(219)) and (inputs(145)));
    layer0_outputs(251) <= not(inputs(150));
    layer0_outputs(252) <= (inputs(250)) and not (inputs(149));
    layer0_outputs(253) <= inputs(25);
    layer0_outputs(254) <= not(inputs(158));
    layer0_outputs(255) <= inputs(175);
    layer0_outputs(256) <= '0';
    layer0_outputs(257) <= inputs(18);
    layer0_outputs(258) <= '1';
    layer0_outputs(259) <= not(inputs(219));
    layer0_outputs(260) <= not((inputs(16)) and (inputs(63)));
    layer0_outputs(261) <= inputs(122);
    layer0_outputs(262) <= (inputs(8)) xor (inputs(34));
    layer0_outputs(263) <= not((inputs(242)) and (inputs(143)));
    layer0_outputs(264) <= '0';
    layer0_outputs(265) <= not(inputs(229));
    layer0_outputs(266) <= not((inputs(202)) and (inputs(208)));
    layer0_outputs(267) <= '1';
    layer0_outputs(268) <= not(inputs(98));
    layer0_outputs(269) <= (inputs(17)) or (inputs(243));
    layer0_outputs(270) <= not(inputs(189));
    layer0_outputs(271) <= not(inputs(82));
    layer0_outputs(272) <= (inputs(212)) or (inputs(190));
    layer0_outputs(273) <= (inputs(140)) xor (inputs(26));
    layer0_outputs(274) <= inputs(106);
    layer0_outputs(275) <= not(inputs(15));
    layer0_outputs(276) <= not(inputs(255));
    layer0_outputs(277) <= inputs(134);
    layer0_outputs(278) <= not(inputs(164)) or (inputs(116));
    layer0_outputs(279) <= not(inputs(84));
    layer0_outputs(280) <= not(inputs(0)) or (inputs(17));
    layer0_outputs(281) <= not(inputs(206)) or (inputs(71));
    layer0_outputs(282) <= '0';
    layer0_outputs(283) <= inputs(9);
    layer0_outputs(284) <= not((inputs(133)) or (inputs(219)));
    layer0_outputs(285) <= not(inputs(146));
    layer0_outputs(286) <= (inputs(99)) xor (inputs(117));
    layer0_outputs(287) <= inputs(9);
    layer0_outputs(288) <= inputs(24);
    layer0_outputs(289) <= inputs(173);
    layer0_outputs(290) <= (inputs(134)) and (inputs(121));
    layer0_outputs(291) <= not(inputs(157));
    layer0_outputs(292) <= inputs(142);
    layer0_outputs(293) <= inputs(162);
    layer0_outputs(294) <= '0';
    layer0_outputs(295) <= '0';
    layer0_outputs(296) <= inputs(180);
    layer0_outputs(297) <= not((inputs(225)) and (inputs(166)));
    layer0_outputs(298) <= '1';
    layer0_outputs(299) <= not((inputs(226)) or (inputs(178)));
    layer0_outputs(300) <= inputs(208);
    layer0_outputs(301) <= inputs(92);
    layer0_outputs(302) <= not((inputs(250)) and (inputs(153)));
    layer0_outputs(303) <= (inputs(146)) and not (inputs(225));
    layer0_outputs(304) <= (inputs(61)) and not (inputs(240));
    layer0_outputs(305) <= inputs(196);
    layer0_outputs(306) <= not(inputs(168));
    layer0_outputs(307) <= not(inputs(110));
    layer0_outputs(308) <= not(inputs(188));
    layer0_outputs(309) <= not(inputs(144));
    layer0_outputs(310) <= inputs(163);
    layer0_outputs(311) <= (inputs(226)) and (inputs(115));
    layer0_outputs(312) <= (inputs(166)) and (inputs(17));
    layer0_outputs(313) <= not((inputs(51)) or (inputs(67)));
    layer0_outputs(314) <= not((inputs(104)) and (inputs(9)));
    layer0_outputs(315) <= not(inputs(129));
    layer0_outputs(316) <= not(inputs(71));
    layer0_outputs(317) <= not(inputs(48));
    layer0_outputs(318) <= not((inputs(155)) or (inputs(179)));
    layer0_outputs(319) <= not((inputs(110)) or (inputs(124)));
    layer0_outputs(320) <= '0';
    layer0_outputs(321) <= '1';
    layer0_outputs(322) <= inputs(113);
    layer0_outputs(323) <= inputs(65);
    layer0_outputs(324) <= (inputs(144)) or (inputs(245));
    layer0_outputs(325) <= not(inputs(42)) or (inputs(156));
    layer0_outputs(326) <= inputs(227);
    layer0_outputs(327) <= (inputs(181)) or (inputs(198));
    layer0_outputs(328) <= not(inputs(250)) or (inputs(17));
    layer0_outputs(329) <= inputs(176);
    layer0_outputs(330) <= not(inputs(162)) or (inputs(16));
    layer0_outputs(331) <= not(inputs(106));
    layer0_outputs(332) <= not(inputs(208)) or (inputs(233));
    layer0_outputs(333) <= '0';
    layer0_outputs(334) <= not(inputs(71)) or (inputs(203));
    layer0_outputs(335) <= (inputs(209)) or (inputs(235));
    layer0_outputs(336) <= inputs(106);
    layer0_outputs(337) <= not(inputs(238));
    layer0_outputs(338) <= inputs(70);
    layer0_outputs(339) <= not((inputs(40)) and (inputs(91)));
    layer0_outputs(340) <= (inputs(163)) and not (inputs(151));
    layer0_outputs(341) <= inputs(237);
    layer0_outputs(342) <= '1';
    layer0_outputs(343) <= '1';
    layer0_outputs(344) <= inputs(146);
    layer0_outputs(345) <= '1';
    layer0_outputs(346) <= (inputs(141)) and not (inputs(239));
    layer0_outputs(347) <= '1';
    layer0_outputs(348) <= not((inputs(136)) and (inputs(221)));
    layer0_outputs(349) <= inputs(50);
    layer0_outputs(350) <= (inputs(241)) and (inputs(160));
    layer0_outputs(351) <= not((inputs(84)) and (inputs(90)));
    layer0_outputs(352) <= inputs(26);
    layer0_outputs(353) <= inputs(77);
    layer0_outputs(354) <= inputs(109);
    layer0_outputs(355) <= '0';
    layer0_outputs(356) <= (inputs(232)) or (inputs(211));
    layer0_outputs(357) <= '0';
    layer0_outputs(358) <= not(inputs(92));
    layer0_outputs(359) <= '0';
    layer0_outputs(360) <= '1';
    layer0_outputs(361) <= '0';
    layer0_outputs(362) <= not(inputs(65));
    layer0_outputs(363) <= not(inputs(67)) or (inputs(33));
    layer0_outputs(364) <= not((inputs(84)) or (inputs(122)));
    layer0_outputs(365) <= (inputs(201)) and not (inputs(119));
    layer0_outputs(366) <= not((inputs(195)) or (inputs(165)));
    layer0_outputs(367) <= not(inputs(126)) or (inputs(3));
    layer0_outputs(368) <= '1';
    layer0_outputs(369) <= '0';
    layer0_outputs(370) <= inputs(147);
    layer0_outputs(371) <= '0';
    layer0_outputs(372) <= '0';
    layer0_outputs(373) <= not(inputs(15));
    layer0_outputs(374) <= inputs(154);
    layer0_outputs(375) <= (inputs(78)) or (inputs(141));
    layer0_outputs(376) <= not((inputs(227)) or (inputs(91)));
    layer0_outputs(377) <= inputs(158);
    layer0_outputs(378) <= not(inputs(77));
    layer0_outputs(379) <= (inputs(187)) and not (inputs(124));
    layer0_outputs(380) <= not(inputs(90));
    layer0_outputs(381) <= (inputs(146)) and not (inputs(80));
    layer0_outputs(382) <= not(inputs(159));
    layer0_outputs(383) <= '1';
    layer0_outputs(384) <= (inputs(136)) and not (inputs(98));
    layer0_outputs(385) <= inputs(38);
    layer0_outputs(386) <= '1';
    layer0_outputs(387) <= '0';
    layer0_outputs(388) <= not(inputs(167));
    layer0_outputs(389) <= not(inputs(1));
    layer0_outputs(390) <= '1';
    layer0_outputs(391) <= (inputs(148)) xor (inputs(103));
    layer0_outputs(392) <= inputs(102);
    layer0_outputs(393) <= inputs(133);
    layer0_outputs(394) <= not((inputs(12)) or (inputs(183)));
    layer0_outputs(395) <= not(inputs(12));
    layer0_outputs(396) <= not((inputs(118)) or (inputs(248)));
    layer0_outputs(397) <= inputs(248);
    layer0_outputs(398) <= '0';
    layer0_outputs(399) <= inputs(58);
    layer0_outputs(400) <= not(inputs(33)) or (inputs(93));
    layer0_outputs(401) <= not(inputs(165));
    layer0_outputs(402) <= (inputs(29)) or (inputs(239));
    layer0_outputs(403) <= '0';
    layer0_outputs(404) <= not(inputs(1)) or (inputs(104));
    layer0_outputs(405) <= inputs(209);
    layer0_outputs(406) <= '1';
    layer0_outputs(407) <= (inputs(127)) and (inputs(79));
    layer0_outputs(408) <= not(inputs(210)) or (inputs(120));
    layer0_outputs(409) <= not(inputs(132)) or (inputs(79));
    layer0_outputs(410) <= (inputs(4)) and not (inputs(82));
    layer0_outputs(411) <= inputs(143);
    layer0_outputs(412) <= (inputs(227)) or (inputs(212));
    layer0_outputs(413) <= inputs(213);
    layer0_outputs(414) <= not(inputs(109));
    layer0_outputs(415) <= not(inputs(40)) or (inputs(240));
    layer0_outputs(416) <= (inputs(141)) and not (inputs(253));
    layer0_outputs(417) <= inputs(245);
    layer0_outputs(418) <= '0';
    layer0_outputs(419) <= not(inputs(22));
    layer0_outputs(420) <= not(inputs(151)) or (inputs(17));
    layer0_outputs(421) <= '1';
    layer0_outputs(422) <= not((inputs(225)) xor (inputs(204)));
    layer0_outputs(423) <= inputs(108);
    layer0_outputs(424) <= inputs(3);
    layer0_outputs(425) <= '1';
    layer0_outputs(426) <= not(inputs(175));
    layer0_outputs(427) <= not(inputs(6)) or (inputs(33));
    layer0_outputs(428) <= not(inputs(125));
    layer0_outputs(429) <= '1';
    layer0_outputs(430) <= inputs(190);
    layer0_outputs(431) <= not((inputs(212)) or (inputs(174)));
    layer0_outputs(432) <= '1';
    layer0_outputs(433) <= '0';
    layer0_outputs(434) <= inputs(210);
    layer0_outputs(435) <= '1';
    layer0_outputs(436) <= (inputs(48)) and not (inputs(40));
    layer0_outputs(437) <= inputs(56);
    layer0_outputs(438) <= (inputs(140)) and (inputs(212));
    layer0_outputs(439) <= (inputs(75)) xor (inputs(253));
    layer0_outputs(440) <= (inputs(174)) and not (inputs(28));
    layer0_outputs(441) <= not(inputs(133));
    layer0_outputs(442) <= '1';
    layer0_outputs(443) <= not(inputs(165));
    layer0_outputs(444) <= not(inputs(184)) or (inputs(61));
    layer0_outputs(445) <= not((inputs(147)) or (inputs(203)));
    layer0_outputs(446) <= not(inputs(18));
    layer0_outputs(447) <= '0';
    layer0_outputs(448) <= not((inputs(191)) or (inputs(240)));
    layer0_outputs(449) <= inputs(67);
    layer0_outputs(450) <= (inputs(105)) or (inputs(135));
    layer0_outputs(451) <= inputs(136);
    layer0_outputs(452) <= (inputs(123)) or (inputs(172));
    layer0_outputs(453) <= (inputs(125)) and (inputs(114));
    layer0_outputs(454) <= '1';
    layer0_outputs(455) <= not(inputs(112));
    layer0_outputs(456) <= not(inputs(145));
    layer0_outputs(457) <= not(inputs(75));
    layer0_outputs(458) <= '1';
    layer0_outputs(459) <= inputs(117);
    layer0_outputs(460) <= inputs(182);
    layer0_outputs(461) <= not((inputs(168)) and (inputs(206)));
    layer0_outputs(462) <= not(inputs(25));
    layer0_outputs(463) <= inputs(107);
    layer0_outputs(464) <= not(inputs(218)) or (inputs(239));
    layer0_outputs(465) <= '1';
    layer0_outputs(466) <= not(inputs(16));
    layer0_outputs(467) <= not((inputs(27)) or (inputs(101)));
    layer0_outputs(468) <= (inputs(96)) and not (inputs(145));
    layer0_outputs(469) <= not(inputs(83));
    layer0_outputs(470) <= (inputs(82)) and (inputs(141));
    layer0_outputs(471) <= (inputs(7)) and (inputs(102));
    layer0_outputs(472) <= not((inputs(46)) and (inputs(94)));
    layer0_outputs(473) <= '1';
    layer0_outputs(474) <= not(inputs(155)) or (inputs(228));
    layer0_outputs(475) <= inputs(234);
    layer0_outputs(476) <= inputs(114);
    layer0_outputs(477) <= inputs(244);
    layer0_outputs(478) <= not((inputs(172)) xor (inputs(118)));
    layer0_outputs(479) <= not(inputs(61)) or (inputs(190));
    layer0_outputs(480) <= (inputs(190)) and not (inputs(249));
    layer0_outputs(481) <= not(inputs(225)) or (inputs(164));
    layer0_outputs(482) <= (inputs(12)) and not (inputs(236));
    layer0_outputs(483) <= not(inputs(107));
    layer0_outputs(484) <= (inputs(31)) xor (inputs(56));
    layer0_outputs(485) <= '1';
    layer0_outputs(486) <= (inputs(65)) xor (inputs(182));
    layer0_outputs(487) <= (inputs(149)) and not (inputs(32));
    layer0_outputs(488) <= not(inputs(174)) or (inputs(12));
    layer0_outputs(489) <= '0';
    layer0_outputs(490) <= not((inputs(62)) xor (inputs(124)));
    layer0_outputs(491) <= inputs(238);
    layer0_outputs(492) <= not(inputs(102)) or (inputs(17));
    layer0_outputs(493) <= inputs(19);
    layer0_outputs(494) <= '1';
    layer0_outputs(495) <= not(inputs(0));
    layer0_outputs(496) <= inputs(25);
    layer0_outputs(497) <= (inputs(149)) or (inputs(201));
    layer0_outputs(498) <= not((inputs(97)) or (inputs(63)));
    layer0_outputs(499) <= inputs(230);
    layer0_outputs(500) <= inputs(104);
    layer0_outputs(501) <= inputs(14);
    layer0_outputs(502) <= '1';
    layer0_outputs(503) <= '1';
    layer0_outputs(504) <= not(inputs(179)) or (inputs(74));
    layer0_outputs(505) <= not(inputs(25));
    layer0_outputs(506) <= not(inputs(110)) or (inputs(209));
    layer0_outputs(507) <= (inputs(116)) or (inputs(160));
    layer0_outputs(508) <= not((inputs(50)) and (inputs(97)));
    layer0_outputs(509) <= not(inputs(60));
    layer0_outputs(510) <= '0';
    layer0_outputs(511) <= '1';
    layer0_outputs(512) <= not(inputs(234));
    layer0_outputs(513) <= not(inputs(142));
    layer0_outputs(514) <= (inputs(64)) and (inputs(217));
    layer0_outputs(515) <= (inputs(120)) and not (inputs(181));
    layer0_outputs(516) <= '1';
    layer0_outputs(517) <= inputs(96);
    layer0_outputs(518) <= not(inputs(213)) or (inputs(30));
    layer0_outputs(519) <= not(inputs(25));
    layer0_outputs(520) <= not(inputs(232)) or (inputs(68));
    layer0_outputs(521) <= not(inputs(185)) or (inputs(47));
    layer0_outputs(522) <= (inputs(20)) and not (inputs(188));
    layer0_outputs(523) <= '0';
    layer0_outputs(524) <= (inputs(163)) and not (inputs(223));
    layer0_outputs(525) <= not(inputs(119)) or (inputs(154));
    layer0_outputs(526) <= not(inputs(68));
    layer0_outputs(527) <= not(inputs(194));
    layer0_outputs(528) <= not(inputs(22));
    layer0_outputs(529) <= not((inputs(218)) and (inputs(55)));
    layer0_outputs(530) <= inputs(102);
    layer0_outputs(531) <= inputs(206);
    layer0_outputs(532) <= not(inputs(72));
    layer0_outputs(533) <= (inputs(36)) and not (inputs(131));
    layer0_outputs(534) <= (inputs(180)) and (inputs(199));
    layer0_outputs(535) <= inputs(11);
    layer0_outputs(536) <= not(inputs(233));
    layer0_outputs(537) <= (inputs(2)) or (inputs(219));
    layer0_outputs(538) <= inputs(173);
    layer0_outputs(539) <= not(inputs(178));
    layer0_outputs(540) <= inputs(215);
    layer0_outputs(541) <= (inputs(39)) and not (inputs(57));
    layer0_outputs(542) <= not(inputs(59)) or (inputs(63));
    layer0_outputs(543) <= '0';
    layer0_outputs(544) <= (inputs(2)) and not (inputs(233));
    layer0_outputs(545) <= '1';
    layer0_outputs(546) <= not(inputs(60)) or (inputs(222));
    layer0_outputs(547) <= not(inputs(194)) or (inputs(167));
    layer0_outputs(548) <= (inputs(232)) and (inputs(219));
    layer0_outputs(549) <= not(inputs(25));
    layer0_outputs(550) <= inputs(247);
    layer0_outputs(551) <= (inputs(4)) and (inputs(39));
    layer0_outputs(552) <= (inputs(75)) and not (inputs(70));
    layer0_outputs(553) <= '1';
    layer0_outputs(554) <= not(inputs(40));
    layer0_outputs(555) <= '1';
    layer0_outputs(556) <= '0';
    layer0_outputs(557) <= not((inputs(66)) xor (inputs(240)));
    layer0_outputs(558) <= (inputs(114)) xor (inputs(79));
    layer0_outputs(559) <= not(inputs(179));
    layer0_outputs(560) <= inputs(165);
    layer0_outputs(561) <= (inputs(169)) or (inputs(216));
    layer0_outputs(562) <= not((inputs(197)) or (inputs(48)));
    layer0_outputs(563) <= not((inputs(230)) or (inputs(65)));
    layer0_outputs(564) <= '1';
    layer0_outputs(565) <= '0';
    layer0_outputs(566) <= (inputs(166)) and not (inputs(132));
    layer0_outputs(567) <= inputs(57);
    layer0_outputs(568) <= not(inputs(128));
    layer0_outputs(569) <= '0';
    layer0_outputs(570) <= '0';
    layer0_outputs(571) <= '1';
    layer0_outputs(572) <= not(inputs(123));
    layer0_outputs(573) <= '1';
    layer0_outputs(574) <= not(inputs(193)) or (inputs(144));
    layer0_outputs(575) <= (inputs(114)) and not (inputs(160));
    layer0_outputs(576) <= inputs(125);
    layer0_outputs(577) <= not(inputs(253));
    layer0_outputs(578) <= inputs(94);
    layer0_outputs(579) <= not((inputs(252)) or (inputs(166)));
    layer0_outputs(580) <= inputs(23);
    layer0_outputs(581) <= '0';
    layer0_outputs(582) <= (inputs(160)) and not (inputs(15));
    layer0_outputs(583) <= inputs(181);
    layer0_outputs(584) <= '0';
    layer0_outputs(585) <= (inputs(22)) or (inputs(138));
    layer0_outputs(586) <= not((inputs(10)) or (inputs(24)));
    layer0_outputs(587) <= not((inputs(151)) and (inputs(102)));
    layer0_outputs(588) <= '1';
    layer0_outputs(589) <= not(inputs(185)) or (inputs(88));
    layer0_outputs(590) <= '1';
    layer0_outputs(591) <= '1';
    layer0_outputs(592) <= (inputs(53)) or (inputs(152));
    layer0_outputs(593) <= (inputs(104)) and not (inputs(251));
    layer0_outputs(594) <= inputs(193);
    layer0_outputs(595) <= not((inputs(239)) or (inputs(96)));
    layer0_outputs(596) <= '0';
    layer0_outputs(597) <= '1';
    layer0_outputs(598) <= not(inputs(131));
    layer0_outputs(599) <= inputs(47);
    layer0_outputs(600) <= not(inputs(153));
    layer0_outputs(601) <= (inputs(8)) or (inputs(10));
    layer0_outputs(602) <= inputs(135);
    layer0_outputs(603) <= (inputs(66)) and not (inputs(191));
    layer0_outputs(604) <= not((inputs(227)) or (inputs(179)));
    layer0_outputs(605) <= '0';
    layer0_outputs(606) <= '0';
    layer0_outputs(607) <= '0';
    layer0_outputs(608) <= not(inputs(113));
    layer0_outputs(609) <= '1';
    layer0_outputs(610) <= (inputs(116)) and (inputs(70));
    layer0_outputs(611) <= (inputs(113)) and (inputs(75));
    layer0_outputs(612) <= (inputs(180)) and not (inputs(97));
    layer0_outputs(613) <= (inputs(190)) and not (inputs(244));
    layer0_outputs(614) <= not((inputs(35)) or (inputs(135)));
    layer0_outputs(615) <= not(inputs(99));
    layer0_outputs(616) <= '1';
    layer0_outputs(617) <= '0';
    layer0_outputs(618) <= inputs(67);
    layer0_outputs(619) <= inputs(69);
    layer0_outputs(620) <= not(inputs(148)) or (inputs(2));
    layer0_outputs(621) <= (inputs(225)) xor (inputs(81));
    layer0_outputs(622) <= not((inputs(90)) xor (inputs(89)));
    layer0_outputs(623) <= (inputs(248)) xor (inputs(239));
    layer0_outputs(624) <= '1';
    layer0_outputs(625) <= '0';
    layer0_outputs(626) <= not(inputs(83));
    layer0_outputs(627) <= '0';
    layer0_outputs(628) <= not(inputs(104));
    layer0_outputs(629) <= '1';
    layer0_outputs(630) <= (inputs(218)) and (inputs(117));
    layer0_outputs(631) <= (inputs(46)) or (inputs(123));
    layer0_outputs(632) <= not(inputs(92));
    layer0_outputs(633) <= '1';
    layer0_outputs(634) <= '0';
    layer0_outputs(635) <= (inputs(16)) and (inputs(88));
    layer0_outputs(636) <= not(inputs(156));
    layer0_outputs(637) <= '1';
    layer0_outputs(638) <= '0';
    layer0_outputs(639) <= '0';
    layer0_outputs(640) <= '0';
    layer0_outputs(641) <= '0';
    layer0_outputs(642) <= not(inputs(193));
    layer0_outputs(643) <= not(inputs(67));
    layer0_outputs(644) <= not(inputs(178));
    layer0_outputs(645) <= inputs(130);
    layer0_outputs(646) <= not(inputs(44));
    layer0_outputs(647) <= inputs(231);
    layer0_outputs(648) <= '0';
    layer0_outputs(649) <= inputs(87);
    layer0_outputs(650) <= (inputs(221)) or (inputs(252));
    layer0_outputs(651) <= (inputs(63)) or (inputs(222));
    layer0_outputs(652) <= (inputs(142)) and not (inputs(190));
    layer0_outputs(653) <= '1';
    layer0_outputs(654) <= (inputs(164)) and not (inputs(9));
    layer0_outputs(655) <= not(inputs(21));
    layer0_outputs(656) <= not(inputs(150));
    layer0_outputs(657) <= inputs(254);
    layer0_outputs(658) <= (inputs(243)) or (inputs(126));
    layer0_outputs(659) <= not((inputs(97)) or (inputs(155)));
    layer0_outputs(660) <= (inputs(221)) or (inputs(177));
    layer0_outputs(661) <= not(inputs(226)) or (inputs(75));
    layer0_outputs(662) <= not(inputs(132));
    layer0_outputs(663) <= '0';
    layer0_outputs(664) <= '0';
    layer0_outputs(665) <= '0';
    layer0_outputs(666) <= inputs(18);
    layer0_outputs(667) <= (inputs(88)) and not (inputs(175));
    layer0_outputs(668) <= not(inputs(57));
    layer0_outputs(669) <= (inputs(125)) and not (inputs(1));
    layer0_outputs(670) <= '0';
    layer0_outputs(671) <= not(inputs(207));
    layer0_outputs(672) <= inputs(78);
    layer0_outputs(673) <= (inputs(178)) or (inputs(82));
    layer0_outputs(674) <= (inputs(127)) or (inputs(159));
    layer0_outputs(675) <= not((inputs(221)) and (inputs(224)));
    layer0_outputs(676) <= inputs(106);
    layer0_outputs(677) <= inputs(229);
    layer0_outputs(678) <= (inputs(152)) and not (inputs(64));
    layer0_outputs(679) <= (inputs(246)) and not (inputs(81));
    layer0_outputs(680) <= (inputs(96)) and not (inputs(80));
    layer0_outputs(681) <= (inputs(216)) and not (inputs(101));
    layer0_outputs(682) <= not(inputs(145));
    layer0_outputs(683) <= inputs(82);
    layer0_outputs(684) <= inputs(160);
    layer0_outputs(685) <= (inputs(88)) and (inputs(81));
    layer0_outputs(686) <= not((inputs(110)) or (inputs(206)));
    layer0_outputs(687) <= not(inputs(237));
    layer0_outputs(688) <= '0';
    layer0_outputs(689) <= not(inputs(231));
    layer0_outputs(690) <= not(inputs(62)) or (inputs(11));
    layer0_outputs(691) <= (inputs(192)) or (inputs(161));
    layer0_outputs(692) <= '0';
    layer0_outputs(693) <= not(inputs(58)) or (inputs(161));
    layer0_outputs(694) <= not((inputs(53)) xor (inputs(94)));
    layer0_outputs(695) <= '0';
    layer0_outputs(696) <= not((inputs(60)) or (inputs(37)));
    layer0_outputs(697) <= '0';
    layer0_outputs(698) <= '0';
    layer0_outputs(699) <= inputs(237);
    layer0_outputs(700) <= not(inputs(164)) or (inputs(201));
    layer0_outputs(701) <= not((inputs(237)) or (inputs(122)));
    layer0_outputs(702) <= not(inputs(231)) or (inputs(229));
    layer0_outputs(703) <= '0';
    layer0_outputs(704) <= '1';
    layer0_outputs(705) <= (inputs(51)) or (inputs(100));
    layer0_outputs(706) <= not(inputs(44));
    layer0_outputs(707) <= inputs(24);
    layer0_outputs(708) <= '0';
    layer0_outputs(709) <= inputs(37);
    layer0_outputs(710) <= not((inputs(162)) xor (inputs(177)));
    layer0_outputs(711) <= not(inputs(1)) or (inputs(59));
    layer0_outputs(712) <= '1';
    layer0_outputs(713) <= not(inputs(150));
    layer0_outputs(714) <= '1';
    layer0_outputs(715) <= (inputs(218)) and not (inputs(134));
    layer0_outputs(716) <= '1';
    layer0_outputs(717) <= (inputs(181)) and not (inputs(47));
    layer0_outputs(718) <= not((inputs(114)) or (inputs(69)));
    layer0_outputs(719) <= '1';
    layer0_outputs(720) <= not((inputs(223)) or (inputs(51)));
    layer0_outputs(721) <= '1';
    layer0_outputs(722) <= not((inputs(243)) or (inputs(198)));
    layer0_outputs(723) <= (inputs(71)) or (inputs(217));
    layer0_outputs(724) <= '1';
    layer0_outputs(725) <= not(inputs(207));
    layer0_outputs(726) <= (inputs(242)) or (inputs(197));
    layer0_outputs(727) <= (inputs(53)) and (inputs(26));
    layer0_outputs(728) <= not((inputs(83)) or (inputs(37)));
    layer0_outputs(729) <= not((inputs(186)) and (inputs(173)));
    layer0_outputs(730) <= '1';
    layer0_outputs(731) <= not(inputs(160));
    layer0_outputs(732) <= (inputs(42)) or (inputs(95));
    layer0_outputs(733) <= inputs(184);
    layer0_outputs(734) <= not(inputs(35));
    layer0_outputs(735) <= not(inputs(79)) or (inputs(110));
    layer0_outputs(736) <= not(inputs(252));
    layer0_outputs(737) <= (inputs(155)) and not (inputs(240));
    layer0_outputs(738) <= (inputs(109)) or (inputs(203));
    layer0_outputs(739) <= (inputs(48)) or (inputs(151));
    layer0_outputs(740) <= (inputs(232)) and not (inputs(117));
    layer0_outputs(741) <= not(inputs(76));
    layer0_outputs(742) <= (inputs(4)) and not (inputs(81));
    layer0_outputs(743) <= not(inputs(162));
    layer0_outputs(744) <= not(inputs(18));
    layer0_outputs(745) <= not(inputs(211));
    layer0_outputs(746) <= not(inputs(126));
    layer0_outputs(747) <= not((inputs(183)) or (inputs(89)));
    layer0_outputs(748) <= not((inputs(113)) and (inputs(43)));
    layer0_outputs(749) <= not(inputs(244)) or (inputs(235));
    layer0_outputs(750) <= inputs(209);
    layer0_outputs(751) <= inputs(177);
    layer0_outputs(752) <= '1';
    layer0_outputs(753) <= (inputs(184)) or (inputs(229));
    layer0_outputs(754) <= '0';
    layer0_outputs(755) <= inputs(178);
    layer0_outputs(756) <= not((inputs(253)) and (inputs(108)));
    layer0_outputs(757) <= not((inputs(64)) and (inputs(26)));
    layer0_outputs(758) <= inputs(246);
    layer0_outputs(759) <= not(inputs(25)) or (inputs(54));
    layer0_outputs(760) <= not(inputs(105)) or (inputs(146));
    layer0_outputs(761) <= inputs(115);
    layer0_outputs(762) <= not((inputs(172)) or (inputs(107)));
    layer0_outputs(763) <= not(inputs(116)) or (inputs(56));
    layer0_outputs(764) <= (inputs(30)) or (inputs(160));
    layer0_outputs(765) <= '1';
    layer0_outputs(766) <= not(inputs(122));
    layer0_outputs(767) <= (inputs(130)) or (inputs(205));
    layer0_outputs(768) <= (inputs(227)) xor (inputs(215));
    layer0_outputs(769) <= inputs(180);
    layer0_outputs(770) <= '0';
    layer0_outputs(771) <= '0';
    layer0_outputs(772) <= '0';
    layer0_outputs(773) <= (inputs(93)) or (inputs(159));
    layer0_outputs(774) <= not(inputs(124));
    layer0_outputs(775) <= not(inputs(165));
    layer0_outputs(776) <= inputs(171);
    layer0_outputs(777) <= not(inputs(198)) or (inputs(144));
    layer0_outputs(778) <= not(inputs(157)) or (inputs(149));
    layer0_outputs(779) <= '0';
    layer0_outputs(780) <= not((inputs(118)) and (inputs(111)));
    layer0_outputs(781) <= '1';
    layer0_outputs(782) <= not(inputs(232));
    layer0_outputs(783) <= not((inputs(79)) or (inputs(212)));
    layer0_outputs(784) <= (inputs(0)) and (inputs(68));
    layer0_outputs(785) <= not((inputs(110)) and (inputs(73)));
    layer0_outputs(786) <= (inputs(231)) and (inputs(133));
    layer0_outputs(787) <= '0';
    layer0_outputs(788) <= inputs(31);
    layer0_outputs(789) <= not(inputs(187));
    layer0_outputs(790) <= '1';
    layer0_outputs(791) <= not(inputs(212)) or (inputs(44));
    layer0_outputs(792) <= (inputs(160)) or (inputs(147));
    layer0_outputs(793) <= (inputs(48)) or (inputs(170));
    layer0_outputs(794) <= not(inputs(207)) or (inputs(158));
    layer0_outputs(795) <= not(inputs(198)) or (inputs(146));
    layer0_outputs(796) <= not(inputs(233));
    layer0_outputs(797) <= '0';
    layer0_outputs(798) <= not((inputs(226)) and (inputs(214)));
    layer0_outputs(799) <= not(inputs(255));
    layer0_outputs(800) <= not(inputs(165));
    layer0_outputs(801) <= '1';
    layer0_outputs(802) <= not(inputs(96)) or (inputs(61));
    layer0_outputs(803) <= inputs(152);
    layer0_outputs(804) <= not(inputs(164));
    layer0_outputs(805) <= not(inputs(214)) or (inputs(98));
    layer0_outputs(806) <= '0';
    layer0_outputs(807) <= (inputs(232)) and not (inputs(242));
    layer0_outputs(808) <= (inputs(116)) or (inputs(76));
    layer0_outputs(809) <= (inputs(147)) or (inputs(180));
    layer0_outputs(810) <= '0';
    layer0_outputs(811) <= (inputs(55)) or (inputs(26));
    layer0_outputs(812) <= (inputs(69)) and not (inputs(167));
    layer0_outputs(813) <= '0';
    layer0_outputs(814) <= '0';
    layer0_outputs(815) <= (inputs(188)) and (inputs(120));
    layer0_outputs(816) <= not(inputs(194));
    layer0_outputs(817) <= inputs(140);
    layer0_outputs(818) <= inputs(102);
    layer0_outputs(819) <= inputs(56);
    layer0_outputs(820) <= inputs(243);
    layer0_outputs(821) <= '1';
    layer0_outputs(822) <= not(inputs(148)) or (inputs(42));
    layer0_outputs(823) <= not(inputs(231));
    layer0_outputs(824) <= not(inputs(126));
    layer0_outputs(825) <= '1';
    layer0_outputs(826) <= (inputs(34)) or (inputs(179));
    layer0_outputs(827) <= '0';
    layer0_outputs(828) <= not(inputs(133)) or (inputs(75));
    layer0_outputs(829) <= '0';
    layer0_outputs(830) <= not((inputs(250)) and (inputs(200)));
    layer0_outputs(831) <= not(inputs(27)) or (inputs(112));
    layer0_outputs(832) <= (inputs(73)) or (inputs(93));
    layer0_outputs(833) <= not((inputs(194)) and (inputs(128)));
    layer0_outputs(834) <= (inputs(169)) and not (inputs(66));
    layer0_outputs(835) <= inputs(43);
    layer0_outputs(836) <= not((inputs(238)) or (inputs(64)));
    layer0_outputs(837) <= (inputs(142)) and not (inputs(210));
    layer0_outputs(838) <= (inputs(103)) or (inputs(72));
    layer0_outputs(839) <= inputs(240);
    layer0_outputs(840) <= (inputs(101)) or (inputs(8));
    layer0_outputs(841) <= not(inputs(54)) or (inputs(189));
    layer0_outputs(842) <= not(inputs(252)) or (inputs(171));
    layer0_outputs(843) <= not(inputs(14)) or (inputs(40));
    layer0_outputs(844) <= (inputs(186)) and (inputs(232));
    layer0_outputs(845) <= not((inputs(193)) or (inputs(82)));
    layer0_outputs(846) <= '0';
    layer0_outputs(847) <= (inputs(83)) or (inputs(199));
    layer0_outputs(848) <= not(inputs(74));
    layer0_outputs(849) <= not(inputs(177));
    layer0_outputs(850) <= inputs(80);
    layer0_outputs(851) <= (inputs(209)) or (inputs(159));
    layer0_outputs(852) <= '0';
    layer0_outputs(853) <= not(inputs(76));
    layer0_outputs(854) <= not(inputs(103));
    layer0_outputs(855) <= (inputs(120)) and not (inputs(142));
    layer0_outputs(856) <= (inputs(109)) or (inputs(149));
    layer0_outputs(857) <= (inputs(156)) and not (inputs(29));
    layer0_outputs(858) <= '0';
    layer0_outputs(859) <= (inputs(231)) and not (inputs(105));
    layer0_outputs(860) <= '0';
    layer0_outputs(861) <= (inputs(163)) or (inputs(64));
    layer0_outputs(862) <= '1';
    layer0_outputs(863) <= inputs(138);
    layer0_outputs(864) <= '0';
    layer0_outputs(865) <= inputs(248);
    layer0_outputs(866) <= inputs(207);
    layer0_outputs(867) <= (inputs(68)) or (inputs(69));
    layer0_outputs(868) <= not((inputs(50)) or (inputs(240)));
    layer0_outputs(869) <= '0';
    layer0_outputs(870) <= not((inputs(143)) and (inputs(80)));
    layer0_outputs(871) <= '1';
    layer0_outputs(872) <= (inputs(32)) or (inputs(7));
    layer0_outputs(873) <= '0';
    layer0_outputs(874) <= not((inputs(163)) or (inputs(11)));
    layer0_outputs(875) <= not((inputs(23)) or (inputs(32)));
    layer0_outputs(876) <= '1';
    layer0_outputs(877) <= (inputs(158)) and not (inputs(238));
    layer0_outputs(878) <= not((inputs(45)) and (inputs(215)));
    layer0_outputs(879) <= not(inputs(142));
    layer0_outputs(880) <= '0';
    layer0_outputs(881) <= not(inputs(193)) or (inputs(31));
    layer0_outputs(882) <= not(inputs(98));
    layer0_outputs(883) <= '1';
    layer0_outputs(884) <= inputs(115);
    layer0_outputs(885) <= not(inputs(210));
    layer0_outputs(886) <= '1';
    layer0_outputs(887) <= '1';
    layer0_outputs(888) <= not((inputs(19)) or (inputs(134)));
    layer0_outputs(889) <= '0';
    layer0_outputs(890) <= not(inputs(49)) or (inputs(212));
    layer0_outputs(891) <= inputs(125);
    layer0_outputs(892) <= not(inputs(35));
    layer0_outputs(893) <= (inputs(193)) or (inputs(249));
    layer0_outputs(894) <= '0';
    layer0_outputs(895) <= (inputs(236)) and not (inputs(197));
    layer0_outputs(896) <= '0';
    layer0_outputs(897) <= '1';
    layer0_outputs(898) <= '1';
    layer0_outputs(899) <= not(inputs(23));
    layer0_outputs(900) <= not(inputs(59));
    layer0_outputs(901) <= '1';
    layer0_outputs(902) <= inputs(113);
    layer0_outputs(903) <= inputs(236);
    layer0_outputs(904) <= not(inputs(97));
    layer0_outputs(905) <= '0';
    layer0_outputs(906) <= '1';
    layer0_outputs(907) <= not((inputs(149)) xor (inputs(177)));
    layer0_outputs(908) <= (inputs(108)) and not (inputs(116));
    layer0_outputs(909) <= (inputs(250)) and (inputs(253));
    layer0_outputs(910) <= (inputs(199)) and not (inputs(43));
    layer0_outputs(911) <= '1';
    layer0_outputs(912) <= not(inputs(227));
    layer0_outputs(913) <= not(inputs(13)) or (inputs(168));
    layer0_outputs(914) <= (inputs(45)) or (inputs(6));
    layer0_outputs(915) <= not((inputs(132)) or (inputs(1)));
    layer0_outputs(916) <= not(inputs(108)) or (inputs(36));
    layer0_outputs(917) <= '0';
    layer0_outputs(918) <= (inputs(12)) and (inputs(222));
    layer0_outputs(919) <= '0';
    layer0_outputs(920) <= inputs(86);
    layer0_outputs(921) <= not((inputs(182)) or (inputs(148)));
    layer0_outputs(922) <= not(inputs(120));
    layer0_outputs(923) <= not(inputs(160)) or (inputs(253));
    layer0_outputs(924) <= not((inputs(191)) or (inputs(200)));
    layer0_outputs(925) <= '0';
    layer0_outputs(926) <= (inputs(141)) and not (inputs(154));
    layer0_outputs(927) <= (inputs(14)) and not (inputs(89));
    layer0_outputs(928) <= '1';
    layer0_outputs(929) <= not(inputs(98)) or (inputs(158));
    layer0_outputs(930) <= not(inputs(199)) or (inputs(225));
    layer0_outputs(931) <= '0';
    layer0_outputs(932) <= (inputs(31)) or (inputs(242));
    layer0_outputs(933) <= not(inputs(105));
    layer0_outputs(934) <= (inputs(41)) and (inputs(206));
    layer0_outputs(935) <= '1';
    layer0_outputs(936) <= (inputs(8)) and not (inputs(162));
    layer0_outputs(937) <= (inputs(213)) and not (inputs(45));
    layer0_outputs(938) <= not(inputs(237));
    layer0_outputs(939) <= not(inputs(104));
    layer0_outputs(940) <= not(inputs(58)) or (inputs(86));
    layer0_outputs(941) <= inputs(32);
    layer0_outputs(942) <= '0';
    layer0_outputs(943) <= (inputs(201)) or (inputs(188));
    layer0_outputs(944) <= inputs(192);
    layer0_outputs(945) <= not((inputs(78)) or (inputs(26)));
    layer0_outputs(946) <= not((inputs(37)) and (inputs(24)));
    layer0_outputs(947) <= inputs(149);
    layer0_outputs(948) <= (inputs(196)) and not (inputs(102));
    layer0_outputs(949) <= '0';
    layer0_outputs(950) <= (inputs(59)) or (inputs(74));
    layer0_outputs(951) <= inputs(53);
    layer0_outputs(952) <= '0';
    layer0_outputs(953) <= (inputs(192)) or (inputs(99));
    layer0_outputs(954) <= inputs(212);
    layer0_outputs(955) <= '0';
    layer0_outputs(956) <= not(inputs(22));
    layer0_outputs(957) <= inputs(25);
    layer0_outputs(958) <= (inputs(65)) and (inputs(89));
    layer0_outputs(959) <= (inputs(156)) or (inputs(77));
    layer0_outputs(960) <= (inputs(160)) or (inputs(115));
    layer0_outputs(961) <= (inputs(214)) or (inputs(24));
    layer0_outputs(962) <= '1';
    layer0_outputs(963) <= (inputs(102)) and not (inputs(191));
    layer0_outputs(964) <= not(inputs(105));
    layer0_outputs(965) <= not((inputs(214)) and (inputs(40)));
    layer0_outputs(966) <= not(inputs(33)) or (inputs(95));
    layer0_outputs(967) <= (inputs(169)) and not (inputs(5));
    layer0_outputs(968) <= '0';
    layer0_outputs(969) <= '0';
    layer0_outputs(970) <= not(inputs(117));
    layer0_outputs(971) <= not(inputs(192));
    layer0_outputs(972) <= inputs(21);
    layer0_outputs(973) <= (inputs(247)) or (inputs(241));
    layer0_outputs(974) <= '0';
    layer0_outputs(975) <= '0';
    layer0_outputs(976) <= inputs(17);
    layer0_outputs(977) <= not((inputs(29)) xor (inputs(54)));
    layer0_outputs(978) <= inputs(99);
    layer0_outputs(979) <= not((inputs(66)) or (inputs(101)));
    layer0_outputs(980) <= inputs(162);
    layer0_outputs(981) <= (inputs(249)) and not (inputs(70));
    layer0_outputs(982) <= not(inputs(52)) or (inputs(234));
    layer0_outputs(983) <= not(inputs(155));
    layer0_outputs(984) <= (inputs(220)) and not (inputs(31));
    layer0_outputs(985) <= not((inputs(36)) xor (inputs(2)));
    layer0_outputs(986) <= not((inputs(138)) and (inputs(16)));
    layer0_outputs(987) <= (inputs(2)) or (inputs(197));
    layer0_outputs(988) <= not(inputs(135));
    layer0_outputs(989) <= (inputs(53)) or (inputs(52));
    layer0_outputs(990) <= not(inputs(76)) or (inputs(47));
    layer0_outputs(991) <= (inputs(159)) xor (inputs(148));
    layer0_outputs(992) <= inputs(56);
    layer0_outputs(993) <= '0';
    layer0_outputs(994) <= not(inputs(10));
    layer0_outputs(995) <= inputs(223);
    layer0_outputs(996) <= '1';
    layer0_outputs(997) <= (inputs(109)) and (inputs(229));
    layer0_outputs(998) <= '0';
    layer0_outputs(999) <= not((inputs(30)) or (inputs(46)));
    layer0_outputs(1000) <= not(inputs(112));
    layer0_outputs(1001) <= (inputs(200)) xor (inputs(248));
    layer0_outputs(1002) <= not(inputs(225));
    layer0_outputs(1003) <= not(inputs(122)) or (inputs(238));
    layer0_outputs(1004) <= inputs(132);
    layer0_outputs(1005) <= '0';
    layer0_outputs(1006) <= '1';
    layer0_outputs(1007) <= inputs(14);
    layer0_outputs(1008) <= (inputs(213)) and (inputs(246));
    layer0_outputs(1009) <= '0';
    layer0_outputs(1010) <= '0';
    layer0_outputs(1011) <= '0';
    layer0_outputs(1012) <= '1';
    layer0_outputs(1013) <= not(inputs(144));
    layer0_outputs(1014) <= inputs(209);
    layer0_outputs(1015) <= '0';
    layer0_outputs(1016) <= not((inputs(42)) or (inputs(59)));
    layer0_outputs(1017) <= not((inputs(148)) or (inputs(6)));
    layer0_outputs(1018) <= not((inputs(200)) and (inputs(174)));
    layer0_outputs(1019) <= not(inputs(28)) or (inputs(163));
    layer0_outputs(1020) <= (inputs(88)) and not (inputs(50));
    layer0_outputs(1021) <= inputs(240);
    layer0_outputs(1022) <= not(inputs(104));
    layer0_outputs(1023) <= (inputs(179)) or (inputs(180));
    layer0_outputs(1024) <= not(inputs(168));
    layer0_outputs(1025) <= '1';
    layer0_outputs(1026) <= inputs(145);
    layer0_outputs(1027) <= (inputs(100)) and not (inputs(17));
    layer0_outputs(1028) <= inputs(183);
    layer0_outputs(1029) <= '0';
    layer0_outputs(1030) <= inputs(195);
    layer0_outputs(1031) <= (inputs(73)) xor (inputs(238));
    layer0_outputs(1032) <= not((inputs(18)) or (inputs(90)));
    layer0_outputs(1033) <= '0';
    layer0_outputs(1034) <= '0';
    layer0_outputs(1035) <= not(inputs(209));
    layer0_outputs(1036) <= inputs(91);
    layer0_outputs(1037) <= not(inputs(107)) or (inputs(193));
    layer0_outputs(1038) <= (inputs(161)) xor (inputs(69));
    layer0_outputs(1039) <= not(inputs(70));
    layer0_outputs(1040) <= inputs(216);
    layer0_outputs(1041) <= inputs(167);
    layer0_outputs(1042) <= not(inputs(132));
    layer0_outputs(1043) <= (inputs(67)) and not (inputs(202));
    layer0_outputs(1044) <= not((inputs(111)) or (inputs(168)));
    layer0_outputs(1045) <= '1';
    layer0_outputs(1046) <= '0';
    layer0_outputs(1047) <= not(inputs(127));
    layer0_outputs(1048) <= inputs(149);
    layer0_outputs(1049) <= inputs(52);
    layer0_outputs(1050) <= not(inputs(111));
    layer0_outputs(1051) <= (inputs(220)) and not (inputs(107));
    layer0_outputs(1052) <= not(inputs(195)) or (inputs(12));
    layer0_outputs(1053) <= inputs(80);
    layer0_outputs(1054) <= not(inputs(232));
    layer0_outputs(1055) <= not(inputs(131)) or (inputs(3));
    layer0_outputs(1056) <= (inputs(10)) and (inputs(15));
    layer0_outputs(1057) <= (inputs(4)) and not (inputs(102));
    layer0_outputs(1058) <= inputs(178);
    layer0_outputs(1059) <= inputs(87);
    layer0_outputs(1060) <= '1';
    layer0_outputs(1061) <= (inputs(252)) or (inputs(89));
    layer0_outputs(1062) <= (inputs(239)) and not (inputs(208));
    layer0_outputs(1063) <= not(inputs(112));
    layer0_outputs(1064) <= inputs(116);
    layer0_outputs(1065) <= inputs(35);
    layer0_outputs(1066) <= not((inputs(52)) and (inputs(53)));
    layer0_outputs(1067) <= (inputs(217)) or (inputs(175));
    layer0_outputs(1068) <= not(inputs(230)) or (inputs(53));
    layer0_outputs(1069) <= '1';
    layer0_outputs(1070) <= inputs(38);
    layer0_outputs(1071) <= not(inputs(165)) or (inputs(241));
    layer0_outputs(1072) <= (inputs(254)) and not (inputs(35));
    layer0_outputs(1073) <= '1';
    layer0_outputs(1074) <= not((inputs(245)) or (inputs(214)));
    layer0_outputs(1075) <= (inputs(63)) and not (inputs(174));
    layer0_outputs(1076) <= inputs(126);
    layer0_outputs(1077) <= not((inputs(78)) or (inputs(4)));
    layer0_outputs(1078) <= inputs(237);
    layer0_outputs(1079) <= inputs(2);
    layer0_outputs(1080) <= inputs(111);
    layer0_outputs(1081) <= inputs(131);
    layer0_outputs(1082) <= '0';
    layer0_outputs(1083) <= not((inputs(119)) or (inputs(103)));
    layer0_outputs(1084) <= not(inputs(248)) or (inputs(83));
    layer0_outputs(1085) <= not((inputs(144)) or (inputs(162)));
    layer0_outputs(1086) <= not((inputs(9)) or (inputs(156)));
    layer0_outputs(1087) <= not(inputs(136)) or (inputs(178));
    layer0_outputs(1088) <= inputs(151);
    layer0_outputs(1089) <= '0';
    layer0_outputs(1090) <= not((inputs(142)) or (inputs(173)));
    layer0_outputs(1091) <= '0';
    layer0_outputs(1092) <= not(inputs(24)) or (inputs(13));
    layer0_outputs(1093) <= '0';
    layer0_outputs(1094) <= not((inputs(141)) and (inputs(11)));
    layer0_outputs(1095) <= not(inputs(63)) or (inputs(23));
    layer0_outputs(1096) <= not(inputs(131));
    layer0_outputs(1097) <= inputs(218);
    layer0_outputs(1098) <= inputs(234);
    layer0_outputs(1099) <= (inputs(8)) and not (inputs(201));
    layer0_outputs(1100) <= not(inputs(195));
    layer0_outputs(1101) <= not(inputs(134));
    layer0_outputs(1102) <= inputs(111);
    layer0_outputs(1103) <= not((inputs(202)) and (inputs(160)));
    layer0_outputs(1104) <= (inputs(52)) or (inputs(117));
    layer0_outputs(1105) <= (inputs(150)) and not (inputs(173));
    layer0_outputs(1106) <= not(inputs(167));
    layer0_outputs(1107) <= not(inputs(202));
    layer0_outputs(1108) <= '0';
    layer0_outputs(1109) <= not(inputs(170));
    layer0_outputs(1110) <= not(inputs(62));
    layer0_outputs(1111) <= '0';
    layer0_outputs(1112) <= (inputs(254)) xor (inputs(127));
    layer0_outputs(1113) <= '0';
    layer0_outputs(1114) <= not(inputs(76)) or (inputs(129));
    layer0_outputs(1115) <= not(inputs(144));
    layer0_outputs(1116) <= not(inputs(95));
    layer0_outputs(1117) <= inputs(194);
    layer0_outputs(1118) <= not(inputs(242)) or (inputs(113));
    layer0_outputs(1119) <= '0';
    layer0_outputs(1120) <= not(inputs(108));
    layer0_outputs(1121) <= (inputs(99)) or (inputs(55));
    layer0_outputs(1122) <= inputs(9);
    layer0_outputs(1123) <= '1';
    layer0_outputs(1124) <= '1';
    layer0_outputs(1125) <= '0';
    layer0_outputs(1126) <= '0';
    layer0_outputs(1127) <= '1';
    layer0_outputs(1128) <= not(inputs(106)) or (inputs(112));
    layer0_outputs(1129) <= not(inputs(26)) or (inputs(150));
    layer0_outputs(1130) <= inputs(150);
    layer0_outputs(1131) <= inputs(196);
    layer0_outputs(1132) <= not(inputs(64)) or (inputs(37));
    layer0_outputs(1133) <= inputs(34);
    layer0_outputs(1134) <= not(inputs(62));
    layer0_outputs(1135) <= not(inputs(45));
    layer0_outputs(1136) <= (inputs(108)) and (inputs(70));
    layer0_outputs(1137) <= not(inputs(154));
    layer0_outputs(1138) <= not(inputs(56)) or (inputs(217));
    layer0_outputs(1139) <= not(inputs(56));
    layer0_outputs(1140) <= '0';
    layer0_outputs(1141) <= (inputs(161)) and not (inputs(29));
    layer0_outputs(1142) <= not((inputs(212)) and (inputs(21)));
    layer0_outputs(1143) <= (inputs(89)) or (inputs(113));
    layer0_outputs(1144) <= not(inputs(194));
    layer0_outputs(1145) <= not(inputs(148));
    layer0_outputs(1146) <= not(inputs(88));
    layer0_outputs(1147) <= not((inputs(106)) or (inputs(107)));
    layer0_outputs(1148) <= '0';
    layer0_outputs(1149) <= not((inputs(182)) or (inputs(185)));
    layer0_outputs(1150) <= (inputs(146)) and not (inputs(255));
    layer0_outputs(1151) <= not((inputs(27)) and (inputs(40)));
    layer0_outputs(1152) <= inputs(151);
    layer0_outputs(1153) <= not(inputs(216)) or (inputs(152));
    layer0_outputs(1154) <= not(inputs(184));
    layer0_outputs(1155) <= '0';
    layer0_outputs(1156) <= not(inputs(255));
    layer0_outputs(1157) <= not((inputs(202)) or (inputs(174)));
    layer0_outputs(1158) <= not(inputs(112));
    layer0_outputs(1159) <= '0';
    layer0_outputs(1160) <= not(inputs(104));
    layer0_outputs(1161) <= not(inputs(245));
    layer0_outputs(1162) <= (inputs(137)) or (inputs(47));
    layer0_outputs(1163) <= not((inputs(203)) xor (inputs(94)));
    layer0_outputs(1164) <= '0';
    layer0_outputs(1165) <= not(inputs(133)) or (inputs(9));
    layer0_outputs(1166) <= '0';
    layer0_outputs(1167) <= inputs(221);
    layer0_outputs(1168) <= not(inputs(105));
    layer0_outputs(1169) <= (inputs(0)) and not (inputs(128));
    layer0_outputs(1170) <= not(inputs(242));
    layer0_outputs(1171) <= inputs(255);
    layer0_outputs(1172) <= (inputs(125)) or (inputs(165));
    layer0_outputs(1173) <= (inputs(185)) and (inputs(144));
    layer0_outputs(1174) <= not((inputs(105)) or (inputs(44)));
    layer0_outputs(1175) <= (inputs(150)) and not (inputs(54));
    layer0_outputs(1176) <= not(inputs(121)) or (inputs(33));
    layer0_outputs(1177) <= not(inputs(143));
    layer0_outputs(1178) <= inputs(255);
    layer0_outputs(1179) <= not((inputs(61)) and (inputs(74)));
    layer0_outputs(1180) <= '0';
    layer0_outputs(1181) <= (inputs(235)) and not (inputs(118));
    layer0_outputs(1182) <= not(inputs(182));
    layer0_outputs(1183) <= (inputs(78)) and (inputs(10));
    layer0_outputs(1184) <= not((inputs(234)) and (inputs(133)));
    layer0_outputs(1185) <= inputs(230);
    layer0_outputs(1186) <= (inputs(115)) and not (inputs(41));
    layer0_outputs(1187) <= not((inputs(159)) and (inputs(199)));
    layer0_outputs(1188) <= not(inputs(202));
    layer0_outputs(1189) <= not(inputs(130));
    layer0_outputs(1190) <= inputs(233);
    layer0_outputs(1191) <= (inputs(37)) and not (inputs(221));
    layer0_outputs(1192) <= not(inputs(146));
    layer0_outputs(1193) <= inputs(222);
    layer0_outputs(1194) <= inputs(179);
    layer0_outputs(1195) <= not(inputs(76));
    layer0_outputs(1196) <= '0';
    layer0_outputs(1197) <= inputs(171);
    layer0_outputs(1198) <= (inputs(115)) and not (inputs(235));
    layer0_outputs(1199) <= '1';
    layer0_outputs(1200) <= not((inputs(189)) xor (inputs(145)));
    layer0_outputs(1201) <= (inputs(12)) and (inputs(106));
    layer0_outputs(1202) <= '0';
    layer0_outputs(1203) <= not(inputs(211));
    layer0_outputs(1204) <= '0';
    layer0_outputs(1205) <= not((inputs(217)) or (inputs(2)));
    layer0_outputs(1206) <= (inputs(210)) and not (inputs(56));
    layer0_outputs(1207) <= not((inputs(209)) and (inputs(156)));
    layer0_outputs(1208) <= not((inputs(55)) and (inputs(123)));
    layer0_outputs(1209) <= not(inputs(206)) or (inputs(24));
    layer0_outputs(1210) <= inputs(30);
    layer0_outputs(1211) <= not(inputs(6));
    layer0_outputs(1212) <= '1';
    layer0_outputs(1213) <= '0';
    layer0_outputs(1214) <= (inputs(145)) or (inputs(86));
    layer0_outputs(1215) <= not((inputs(171)) xor (inputs(92)));
    layer0_outputs(1216) <= '0';
    layer0_outputs(1217) <= '0';
    layer0_outputs(1218) <= not(inputs(128)) or (inputs(7));
    layer0_outputs(1219) <= inputs(85);
    layer0_outputs(1220) <= not((inputs(129)) and (inputs(129)));
    layer0_outputs(1221) <= not(inputs(9));
    layer0_outputs(1222) <= not(inputs(198));
    layer0_outputs(1223) <= inputs(22);
    layer0_outputs(1224) <= (inputs(200)) and (inputs(5));
    layer0_outputs(1225) <= inputs(1);
    layer0_outputs(1226) <= not(inputs(67));
    layer0_outputs(1227) <= inputs(55);
    layer0_outputs(1228) <= '0';
    layer0_outputs(1229) <= (inputs(200)) and not (inputs(244));
    layer0_outputs(1230) <= (inputs(121)) and not (inputs(200));
    layer0_outputs(1231) <= not(inputs(103));
    layer0_outputs(1232) <= not((inputs(131)) or (inputs(211)));
    layer0_outputs(1233) <= '1';
    layer0_outputs(1234) <= not(inputs(118)) or (inputs(234));
    layer0_outputs(1235) <= (inputs(169)) and not (inputs(61));
    layer0_outputs(1236) <= (inputs(183)) and not (inputs(96));
    layer0_outputs(1237) <= inputs(155);
    layer0_outputs(1238) <= (inputs(41)) or (inputs(34));
    layer0_outputs(1239) <= not(inputs(207));
    layer0_outputs(1240) <= (inputs(139)) and (inputs(228));
    layer0_outputs(1241) <= inputs(71);
    layer0_outputs(1242) <= not((inputs(150)) or (inputs(151)));
    layer0_outputs(1243) <= (inputs(135)) and not (inputs(0));
    layer0_outputs(1244) <= not(inputs(100));
    layer0_outputs(1245) <= '1';
    layer0_outputs(1246) <= not(inputs(17));
    layer0_outputs(1247) <= not(inputs(183));
    layer0_outputs(1248) <= (inputs(199)) or (inputs(95));
    layer0_outputs(1249) <= '0';
    layer0_outputs(1250) <= '0';
    layer0_outputs(1251) <= (inputs(178)) and not (inputs(229));
    layer0_outputs(1252) <= '0';
    layer0_outputs(1253) <= not(inputs(237));
    layer0_outputs(1254) <= '1';
    layer0_outputs(1255) <= not((inputs(47)) or (inputs(219)));
    layer0_outputs(1256) <= not(inputs(14)) or (inputs(226));
    layer0_outputs(1257) <= (inputs(19)) and not (inputs(146));
    layer0_outputs(1258) <= not(inputs(238));
    layer0_outputs(1259) <= not(inputs(33));
    layer0_outputs(1260) <= '0';
    layer0_outputs(1261) <= not(inputs(46)) or (inputs(175));
    layer0_outputs(1262) <= not(inputs(210)) or (inputs(237));
    layer0_outputs(1263) <= (inputs(59)) or (inputs(91));
    layer0_outputs(1264) <= not(inputs(12)) or (inputs(194));
    layer0_outputs(1265) <= not(inputs(189)) or (inputs(217));
    layer0_outputs(1266) <= not((inputs(66)) xor (inputs(69)));
    layer0_outputs(1267) <= not(inputs(195));
    layer0_outputs(1268) <= not((inputs(134)) and (inputs(147)));
    layer0_outputs(1269) <= (inputs(48)) and not (inputs(170));
    layer0_outputs(1270) <= '0';
    layer0_outputs(1271) <= (inputs(220)) or (inputs(236));
    layer0_outputs(1272) <= not(inputs(101)) or (inputs(17));
    layer0_outputs(1273) <= (inputs(158)) or (inputs(21));
    layer0_outputs(1274) <= not(inputs(167));
    layer0_outputs(1275) <= (inputs(210)) and (inputs(89));
    layer0_outputs(1276) <= (inputs(162)) or (inputs(175));
    layer0_outputs(1277) <= not(inputs(182));
    layer0_outputs(1278) <= '0';
    layer0_outputs(1279) <= not(inputs(228));
    layer0_outputs(1280) <= inputs(181);
    layer0_outputs(1281) <= not(inputs(131));
    layer0_outputs(1282) <= not(inputs(43));
    layer0_outputs(1283) <= (inputs(152)) and not (inputs(65));
    layer0_outputs(1284) <= not(inputs(63)) or (inputs(95));
    layer0_outputs(1285) <= not(inputs(185));
    layer0_outputs(1286) <= not(inputs(25)) or (inputs(98));
    layer0_outputs(1287) <= not(inputs(38));
    layer0_outputs(1288) <= '1';
    layer0_outputs(1289) <= '1';
    layer0_outputs(1290) <= (inputs(70)) and not (inputs(19));
    layer0_outputs(1291) <= inputs(127);
    layer0_outputs(1292) <= '0';
    layer0_outputs(1293) <= (inputs(200)) xor (inputs(39));
    layer0_outputs(1294) <= not(inputs(110));
    layer0_outputs(1295) <= '0';
    layer0_outputs(1296) <= '1';
    layer0_outputs(1297) <= not((inputs(19)) or (inputs(52)));
    layer0_outputs(1298) <= not(inputs(7));
    layer0_outputs(1299) <= '1';
    layer0_outputs(1300) <= inputs(126);
    layer0_outputs(1301) <= not((inputs(241)) and (inputs(185)));
    layer0_outputs(1302) <= not(inputs(70));
    layer0_outputs(1303) <= inputs(44);
    layer0_outputs(1304) <= not((inputs(49)) xor (inputs(78)));
    layer0_outputs(1305) <= inputs(103);
    layer0_outputs(1306) <= '0';
    layer0_outputs(1307) <= inputs(21);
    layer0_outputs(1308) <= '0';
    layer0_outputs(1309) <= '1';
    layer0_outputs(1310) <= (inputs(123)) and (inputs(185));
    layer0_outputs(1311) <= not(inputs(135));
    layer0_outputs(1312) <= not(inputs(175));
    layer0_outputs(1313) <= '0';
    layer0_outputs(1314) <= inputs(251);
    layer0_outputs(1315) <= '1';
    layer0_outputs(1316) <= inputs(115);
    layer0_outputs(1317) <= not((inputs(131)) and (inputs(239)));
    layer0_outputs(1318) <= (inputs(28)) xor (inputs(145));
    layer0_outputs(1319) <= inputs(165);
    layer0_outputs(1320) <= (inputs(174)) and (inputs(54));
    layer0_outputs(1321) <= not((inputs(238)) or (inputs(224)));
    layer0_outputs(1322) <= inputs(169);
    layer0_outputs(1323) <= '1';
    layer0_outputs(1324) <= not(inputs(154)) or (inputs(107));
    layer0_outputs(1325) <= (inputs(28)) and (inputs(182));
    layer0_outputs(1326) <= not((inputs(246)) or (inputs(132)));
    layer0_outputs(1327) <= not(inputs(223)) or (inputs(52));
    layer0_outputs(1328) <= not(inputs(40));
    layer0_outputs(1329) <= not(inputs(122));
    layer0_outputs(1330) <= not((inputs(83)) xor (inputs(219)));
    layer0_outputs(1331) <= inputs(134);
    layer0_outputs(1332) <= (inputs(117)) and not (inputs(231));
    layer0_outputs(1333) <= inputs(91);
    layer0_outputs(1334) <= (inputs(119)) or (inputs(146));
    layer0_outputs(1335) <= not((inputs(153)) and (inputs(226)));
    layer0_outputs(1336) <= not((inputs(15)) or (inputs(130)));
    layer0_outputs(1337) <= not(inputs(121));
    layer0_outputs(1338) <= '1';
    layer0_outputs(1339) <= (inputs(223)) and (inputs(220));
    layer0_outputs(1340) <= '0';
    layer0_outputs(1341) <= (inputs(117)) and not (inputs(92));
    layer0_outputs(1342) <= not(inputs(224)) or (inputs(46));
    layer0_outputs(1343) <= (inputs(171)) and not (inputs(92));
    layer0_outputs(1344) <= '1';
    layer0_outputs(1345) <= not((inputs(73)) xor (inputs(254)));
    layer0_outputs(1346) <= '1';
    layer0_outputs(1347) <= (inputs(139)) and (inputs(57));
    layer0_outputs(1348) <= (inputs(92)) and (inputs(84));
    layer0_outputs(1349) <= '1';
    layer0_outputs(1350) <= inputs(203);
    layer0_outputs(1351) <= '1';
    layer0_outputs(1352) <= '1';
    layer0_outputs(1353) <= '0';
    layer0_outputs(1354) <= not(inputs(203));
    layer0_outputs(1355) <= '1';
    layer0_outputs(1356) <= (inputs(179)) or (inputs(95));
    layer0_outputs(1357) <= not(inputs(102));
    layer0_outputs(1358) <= (inputs(69)) and not (inputs(237));
    layer0_outputs(1359) <= not(inputs(210)) or (inputs(249));
    layer0_outputs(1360) <= not((inputs(241)) and (inputs(45)));
    layer0_outputs(1361) <= (inputs(111)) and not (inputs(121));
    layer0_outputs(1362) <= '1';
    layer0_outputs(1363) <= not((inputs(138)) or (inputs(4)));
    layer0_outputs(1364) <= inputs(21);
    layer0_outputs(1365) <= not(inputs(108));
    layer0_outputs(1366) <= (inputs(141)) or (inputs(145));
    layer0_outputs(1367) <= not(inputs(155)) or (inputs(8));
    layer0_outputs(1368) <= (inputs(129)) xor (inputs(23));
    layer0_outputs(1369) <= inputs(151);
    layer0_outputs(1370) <= '1';
    layer0_outputs(1371) <= not(inputs(86));
    layer0_outputs(1372) <= '0';
    layer0_outputs(1373) <= not(inputs(252));
    layer0_outputs(1374) <= (inputs(67)) and (inputs(186));
    layer0_outputs(1375) <= not((inputs(110)) and (inputs(235)));
    layer0_outputs(1376) <= inputs(181);
    layer0_outputs(1377) <= not(inputs(141)) or (inputs(80));
    layer0_outputs(1378) <= inputs(216);
    layer0_outputs(1379) <= not(inputs(254)) or (inputs(6));
    layer0_outputs(1380) <= inputs(43);
    layer0_outputs(1381) <= inputs(105);
    layer0_outputs(1382) <= '0';
    layer0_outputs(1383) <= '1';
    layer0_outputs(1384) <= not(inputs(211)) or (inputs(103));
    layer0_outputs(1385) <= '0';
    layer0_outputs(1386) <= (inputs(39)) or (inputs(127));
    layer0_outputs(1387) <= inputs(77);
    layer0_outputs(1388) <= (inputs(159)) and not (inputs(81));
    layer0_outputs(1389) <= inputs(153);
    layer0_outputs(1390) <= inputs(127);
    layer0_outputs(1391) <= not(inputs(231));
    layer0_outputs(1392) <= (inputs(194)) or (inputs(66));
    layer0_outputs(1393) <= (inputs(56)) and (inputs(70));
    layer0_outputs(1394) <= inputs(41);
    layer0_outputs(1395) <= inputs(176);
    layer0_outputs(1396) <= '0';
    layer0_outputs(1397) <= not(inputs(9));
    layer0_outputs(1398) <= not(inputs(210));
    layer0_outputs(1399) <= not(inputs(65));
    layer0_outputs(1400) <= (inputs(39)) and (inputs(170));
    layer0_outputs(1401) <= '1';
    layer0_outputs(1402) <= not(inputs(21));
    layer0_outputs(1403) <= '0';
    layer0_outputs(1404) <= not(inputs(219)) or (inputs(63));
    layer0_outputs(1405) <= (inputs(30)) or (inputs(60));
    layer0_outputs(1406) <= not((inputs(175)) and (inputs(196)));
    layer0_outputs(1407) <= inputs(182);
    layer0_outputs(1408) <= (inputs(148)) or (inputs(117));
    layer0_outputs(1409) <= not((inputs(31)) or (inputs(168)));
    layer0_outputs(1410) <= inputs(254);
    layer0_outputs(1411) <= '1';
    layer0_outputs(1412) <= not(inputs(111));
    layer0_outputs(1413) <= not(inputs(33));
    layer0_outputs(1414) <= inputs(114);
    layer0_outputs(1415) <= inputs(17);
    layer0_outputs(1416) <= not((inputs(6)) or (inputs(75)));
    layer0_outputs(1417) <= '1';
    layer0_outputs(1418) <= '0';
    layer0_outputs(1419) <= inputs(140);
    layer0_outputs(1420) <= not((inputs(83)) and (inputs(241)));
    layer0_outputs(1421) <= '1';
    layer0_outputs(1422) <= '1';
    layer0_outputs(1423) <= not(inputs(192)) or (inputs(156));
    layer0_outputs(1424) <= (inputs(244)) and (inputs(36));
    layer0_outputs(1425) <= not(inputs(94));
    layer0_outputs(1426) <= not(inputs(95)) or (inputs(164));
    layer0_outputs(1427) <= inputs(33);
    layer0_outputs(1428) <= not(inputs(211));
    layer0_outputs(1429) <= (inputs(244)) and not (inputs(137));
    layer0_outputs(1430) <= '1';
    layer0_outputs(1431) <= not(inputs(105));
    layer0_outputs(1432) <= not(inputs(210)) or (inputs(157));
    layer0_outputs(1433) <= not(inputs(196));
    layer0_outputs(1434) <= '1';
    layer0_outputs(1435) <= (inputs(159)) and not (inputs(95));
    layer0_outputs(1436) <= inputs(148);
    layer0_outputs(1437) <= '1';
    layer0_outputs(1438) <= inputs(193);
    layer0_outputs(1439) <= not((inputs(202)) and (inputs(165)));
    layer0_outputs(1440) <= not(inputs(126));
    layer0_outputs(1441) <= '0';
    layer0_outputs(1442) <= (inputs(49)) and (inputs(188));
    layer0_outputs(1443) <= inputs(82);
    layer0_outputs(1444) <= (inputs(251)) and not (inputs(121));
    layer0_outputs(1445) <= (inputs(201)) and (inputs(236));
    layer0_outputs(1446) <= inputs(194);
    layer0_outputs(1447) <= not(inputs(148));
    layer0_outputs(1448) <= not(inputs(71)) or (inputs(0));
    layer0_outputs(1449) <= (inputs(46)) or (inputs(48));
    layer0_outputs(1450) <= (inputs(251)) xor (inputs(53));
    layer0_outputs(1451) <= '0';
    layer0_outputs(1452) <= inputs(121);
    layer0_outputs(1453) <= not(inputs(165));
    layer0_outputs(1454) <= (inputs(85)) and not (inputs(67));
    layer0_outputs(1455) <= not(inputs(238));
    layer0_outputs(1456) <= '0';
    layer0_outputs(1457) <= inputs(24);
    layer0_outputs(1458) <= not(inputs(133)) or (inputs(8));
    layer0_outputs(1459) <= not(inputs(76)) or (inputs(207));
    layer0_outputs(1460) <= not(inputs(160));
    layer0_outputs(1461) <= (inputs(237)) and not (inputs(51));
    layer0_outputs(1462) <= '0';
    layer0_outputs(1463) <= not(inputs(128));
    layer0_outputs(1464) <= (inputs(57)) or (inputs(115));
    layer0_outputs(1465) <= (inputs(83)) xor (inputs(113));
    layer0_outputs(1466) <= '1';
    layer0_outputs(1467) <= not(inputs(247));
    layer0_outputs(1468) <= (inputs(248)) or (inputs(158));
    layer0_outputs(1469) <= inputs(207);
    layer0_outputs(1470) <= '1';
    layer0_outputs(1471) <= not(inputs(161)) or (inputs(183));
    layer0_outputs(1472) <= inputs(120);
    layer0_outputs(1473) <= (inputs(65)) or (inputs(158));
    layer0_outputs(1474) <= (inputs(102)) and not (inputs(156));
    layer0_outputs(1475) <= inputs(208);
    layer0_outputs(1476) <= (inputs(99)) or (inputs(154));
    layer0_outputs(1477) <= not((inputs(220)) and (inputs(173)));
    layer0_outputs(1478) <= (inputs(202)) and (inputs(118));
    layer0_outputs(1479) <= inputs(14);
    layer0_outputs(1480) <= not((inputs(18)) or (inputs(120)));
    layer0_outputs(1481) <= inputs(110);
    layer0_outputs(1482) <= '0';
    layer0_outputs(1483) <= (inputs(244)) and (inputs(200));
    layer0_outputs(1484) <= not((inputs(205)) or (inputs(223)));
    layer0_outputs(1485) <= (inputs(44)) or (inputs(58));
    layer0_outputs(1486) <= inputs(99);
    layer0_outputs(1487) <= not((inputs(28)) or (inputs(34)));
    layer0_outputs(1488) <= not((inputs(71)) or (inputs(20)));
    layer0_outputs(1489) <= not(inputs(217)) or (inputs(233));
    layer0_outputs(1490) <= '0';
    layer0_outputs(1491) <= '0';
    layer0_outputs(1492) <= not(inputs(107));
    layer0_outputs(1493) <= not(inputs(201)) or (inputs(59));
    layer0_outputs(1494) <= inputs(199);
    layer0_outputs(1495) <= '0';
    layer0_outputs(1496) <= '0';
    layer0_outputs(1497) <= '1';
    layer0_outputs(1498) <= '0';
    layer0_outputs(1499) <= not(inputs(50));
    layer0_outputs(1500) <= not(inputs(231)) or (inputs(5));
    layer0_outputs(1501) <= not((inputs(155)) and (inputs(82)));
    layer0_outputs(1502) <= '0';
    layer0_outputs(1503) <= not(inputs(225));
    layer0_outputs(1504) <= (inputs(5)) or (inputs(109));
    layer0_outputs(1505) <= not(inputs(198));
    layer0_outputs(1506) <= not((inputs(110)) or (inputs(172)));
    layer0_outputs(1507) <= inputs(170);
    layer0_outputs(1508) <= '0';
    layer0_outputs(1509) <= inputs(119);
    layer0_outputs(1510) <= '0';
    layer0_outputs(1511) <= (inputs(38)) and not (inputs(88));
    layer0_outputs(1512) <= inputs(45);
    layer0_outputs(1513) <= '0';
    layer0_outputs(1514) <= not((inputs(210)) or (inputs(41)));
    layer0_outputs(1515) <= (inputs(89)) or (inputs(59));
    layer0_outputs(1516) <= not(inputs(136));
    layer0_outputs(1517) <= inputs(79);
    layer0_outputs(1518) <= not(inputs(12));
    layer0_outputs(1519) <= not(inputs(130));
    layer0_outputs(1520) <= not((inputs(89)) or (inputs(8)));
    layer0_outputs(1521) <= (inputs(26)) and (inputs(22));
    layer0_outputs(1522) <= inputs(85);
    layer0_outputs(1523) <= (inputs(108)) and not (inputs(4));
    layer0_outputs(1524) <= '1';
    layer0_outputs(1525) <= (inputs(219)) or (inputs(35));
    layer0_outputs(1526) <= not(inputs(76));
    layer0_outputs(1527) <= (inputs(23)) and not (inputs(199));
    layer0_outputs(1528) <= not(inputs(48));
    layer0_outputs(1529) <= inputs(163);
    layer0_outputs(1530) <= not((inputs(138)) or (inputs(20)));
    layer0_outputs(1531) <= not(inputs(4));
    layer0_outputs(1532) <= not(inputs(25)) or (inputs(219));
    layer0_outputs(1533) <= (inputs(171)) and not (inputs(111));
    layer0_outputs(1534) <= not(inputs(217)) or (inputs(158));
    layer0_outputs(1535) <= not(inputs(18));
    layer0_outputs(1536) <= (inputs(168)) and (inputs(111));
    layer0_outputs(1537) <= not(inputs(36)) or (inputs(14));
    layer0_outputs(1538) <= not((inputs(198)) or (inputs(183)));
    layer0_outputs(1539) <= not((inputs(79)) or (inputs(92)));
    layer0_outputs(1540) <= (inputs(85)) and not (inputs(78));
    layer0_outputs(1541) <= not(inputs(23));
    layer0_outputs(1542) <= not(inputs(85));
    layer0_outputs(1543) <= inputs(82);
    layer0_outputs(1544) <= inputs(247);
    layer0_outputs(1545) <= not(inputs(181)) or (inputs(28));
    layer0_outputs(1546) <= not(inputs(226));
    layer0_outputs(1547) <= '0';
    layer0_outputs(1548) <= '1';
    layer0_outputs(1549) <= not((inputs(177)) or (inputs(41)));
    layer0_outputs(1550) <= not(inputs(147));
    layer0_outputs(1551) <= '1';
    layer0_outputs(1552) <= not(inputs(156)) or (inputs(85));
    layer0_outputs(1553) <= not((inputs(113)) and (inputs(79)));
    layer0_outputs(1554) <= (inputs(208)) or (inputs(173));
    layer0_outputs(1555) <= (inputs(169)) and (inputs(137));
    layer0_outputs(1556) <= not(inputs(193));
    layer0_outputs(1557) <= not(inputs(232)) or (inputs(184));
    layer0_outputs(1558) <= inputs(248);
    layer0_outputs(1559) <= '0';
    layer0_outputs(1560) <= not((inputs(218)) or (inputs(157)));
    layer0_outputs(1561) <= (inputs(31)) or (inputs(225));
    layer0_outputs(1562) <= '1';
    layer0_outputs(1563) <= not((inputs(125)) or (inputs(187)));
    layer0_outputs(1564) <= (inputs(197)) and not (inputs(109));
    layer0_outputs(1565) <= inputs(218);
    layer0_outputs(1566) <= not((inputs(208)) or (inputs(140)));
    layer0_outputs(1567) <= not(inputs(103)) or (inputs(16));
    layer0_outputs(1568) <= (inputs(162)) and not (inputs(171));
    layer0_outputs(1569) <= not(inputs(110));
    layer0_outputs(1570) <= not(inputs(172));
    layer0_outputs(1571) <= '0';
    layer0_outputs(1572) <= not(inputs(56));
    layer0_outputs(1573) <= not((inputs(253)) and (inputs(144)));
    layer0_outputs(1574) <= not((inputs(223)) and (inputs(224)));
    layer0_outputs(1575) <= not((inputs(128)) or (inputs(142)));
    layer0_outputs(1576) <= not((inputs(85)) or (inputs(212)));
    layer0_outputs(1577) <= not(inputs(47));
    layer0_outputs(1578) <= '0';
    layer0_outputs(1579) <= '1';
    layer0_outputs(1580) <= (inputs(67)) and not (inputs(218));
    layer0_outputs(1581) <= (inputs(27)) and not (inputs(216));
    layer0_outputs(1582) <= not(inputs(29)) or (inputs(142));
    layer0_outputs(1583) <= not(inputs(84));
    layer0_outputs(1584) <= not(inputs(99));
    layer0_outputs(1585) <= not(inputs(78));
    layer0_outputs(1586) <= (inputs(229)) and not (inputs(234));
    layer0_outputs(1587) <= (inputs(130)) or (inputs(188));
    layer0_outputs(1588) <= not(inputs(245)) or (inputs(41));
    layer0_outputs(1589) <= '0';
    layer0_outputs(1590) <= not(inputs(252)) or (inputs(1));
    layer0_outputs(1591) <= '1';
    layer0_outputs(1592) <= not((inputs(105)) or (inputs(32)));
    layer0_outputs(1593) <= not(inputs(130));
    layer0_outputs(1594) <= '0';
    layer0_outputs(1595) <= '0';
    layer0_outputs(1596) <= not((inputs(9)) or (inputs(22)));
    layer0_outputs(1597) <= not((inputs(161)) or (inputs(162)));
    layer0_outputs(1598) <= not((inputs(16)) xor (inputs(48)));
    layer0_outputs(1599) <= inputs(83);
    layer0_outputs(1600) <= not((inputs(191)) or (inputs(207)));
    layer0_outputs(1601) <= not(inputs(71)) or (inputs(142));
    layer0_outputs(1602) <= '1';
    layer0_outputs(1603) <= not(inputs(68)) or (inputs(50));
    layer0_outputs(1604) <= inputs(217);
    layer0_outputs(1605) <= (inputs(92)) or (inputs(171));
    layer0_outputs(1606) <= not(inputs(78)) or (inputs(230));
    layer0_outputs(1607) <= inputs(147);
    layer0_outputs(1608) <= (inputs(177)) or (inputs(226));
    layer0_outputs(1609) <= not((inputs(122)) or (inputs(179)));
    layer0_outputs(1610) <= inputs(62);
    layer0_outputs(1611) <= '0';
    layer0_outputs(1612) <= (inputs(112)) or (inputs(113));
    layer0_outputs(1613) <= '1';
    layer0_outputs(1614) <= '1';
    layer0_outputs(1615) <= (inputs(83)) and (inputs(134));
    layer0_outputs(1616) <= (inputs(226)) and (inputs(124));
    layer0_outputs(1617) <= inputs(36);
    layer0_outputs(1618) <= inputs(197);
    layer0_outputs(1619) <= inputs(25);
    layer0_outputs(1620) <= '0';
    layer0_outputs(1621) <= not((inputs(141)) or (inputs(200)));
    layer0_outputs(1622) <= not(inputs(216)) or (inputs(198));
    layer0_outputs(1623) <= '1';
    layer0_outputs(1624) <= not((inputs(155)) or (inputs(94)));
    layer0_outputs(1625) <= '1';
    layer0_outputs(1626) <= inputs(104);
    layer0_outputs(1627) <= not(inputs(179)) or (inputs(138));
    layer0_outputs(1628) <= (inputs(22)) and not (inputs(55));
    layer0_outputs(1629) <= not((inputs(220)) xor (inputs(140)));
    layer0_outputs(1630) <= (inputs(16)) or (inputs(154));
    layer0_outputs(1631) <= (inputs(130)) xor (inputs(246));
    layer0_outputs(1632) <= '1';
    layer0_outputs(1633) <= inputs(73);
    layer0_outputs(1634) <= (inputs(123)) and (inputs(102));
    layer0_outputs(1635) <= not(inputs(91));
    layer0_outputs(1636) <= '1';
    layer0_outputs(1637) <= not(inputs(49));
    layer0_outputs(1638) <= not((inputs(218)) or (inputs(52)));
    layer0_outputs(1639) <= not((inputs(97)) or (inputs(170)));
    layer0_outputs(1640) <= not(inputs(105)) or (inputs(112));
    layer0_outputs(1641) <= '0';
    layer0_outputs(1642) <= (inputs(29)) and not (inputs(118));
    layer0_outputs(1643) <= '0';
    layer0_outputs(1644) <= '1';
    layer0_outputs(1645) <= not(inputs(123));
    layer0_outputs(1646) <= not(inputs(230)) or (inputs(223));
    layer0_outputs(1647) <= (inputs(120)) and not (inputs(156));
    layer0_outputs(1648) <= (inputs(238)) or (inputs(203));
    layer0_outputs(1649) <= not(inputs(100));
    layer0_outputs(1650) <= (inputs(198)) and (inputs(220));
    layer0_outputs(1651) <= inputs(101);
    layer0_outputs(1652) <= not(inputs(121)) or (inputs(230));
    layer0_outputs(1653) <= not(inputs(221));
    layer0_outputs(1654) <= not(inputs(167));
    layer0_outputs(1655) <= inputs(60);
    layer0_outputs(1656) <= not(inputs(56));
    layer0_outputs(1657) <= inputs(215);
    layer0_outputs(1658) <= not((inputs(156)) or (inputs(127)));
    layer0_outputs(1659) <= inputs(172);
    layer0_outputs(1660) <= not(inputs(42)) or (inputs(178));
    layer0_outputs(1661) <= (inputs(170)) and (inputs(107));
    layer0_outputs(1662) <= inputs(167);
    layer0_outputs(1663) <= not(inputs(204));
    layer0_outputs(1664) <= '0';
    layer0_outputs(1665) <= not(inputs(88)) or (inputs(168));
    layer0_outputs(1666) <= inputs(194);
    layer0_outputs(1667) <= '1';
    layer0_outputs(1668) <= (inputs(193)) and not (inputs(238));
    layer0_outputs(1669) <= not(inputs(147));
    layer0_outputs(1670) <= (inputs(208)) or (inputs(232));
    layer0_outputs(1671) <= '1';
    layer0_outputs(1672) <= (inputs(156)) or (inputs(222));
    layer0_outputs(1673) <= '1';
    layer0_outputs(1674) <= not(inputs(176));
    layer0_outputs(1675) <= not((inputs(147)) or (inputs(113)));
    layer0_outputs(1676) <= not(inputs(65));
    layer0_outputs(1677) <= (inputs(93)) or (inputs(44));
    layer0_outputs(1678) <= not(inputs(222));
    layer0_outputs(1679) <= inputs(120);
    layer0_outputs(1680) <= (inputs(195)) and not (inputs(183));
    layer0_outputs(1681) <= not(inputs(165));
    layer0_outputs(1682) <= not(inputs(112));
    layer0_outputs(1683) <= inputs(230);
    layer0_outputs(1684) <= inputs(3);
    layer0_outputs(1685) <= inputs(196);
    layer0_outputs(1686) <= not(inputs(239)) or (inputs(189));
    layer0_outputs(1687) <= not((inputs(253)) or (inputs(23)));
    layer0_outputs(1688) <= (inputs(31)) or (inputs(22));
    layer0_outputs(1689) <= (inputs(142)) xor (inputs(191));
    layer0_outputs(1690) <= (inputs(249)) or (inputs(109));
    layer0_outputs(1691) <= inputs(110);
    layer0_outputs(1692) <= '1';
    layer0_outputs(1693) <= inputs(49);
    layer0_outputs(1694) <= (inputs(212)) or (inputs(206));
    layer0_outputs(1695) <= (inputs(190)) or (inputs(145));
    layer0_outputs(1696) <= not((inputs(9)) xor (inputs(222)));
    layer0_outputs(1697) <= '0';
    layer0_outputs(1698) <= '0';
    layer0_outputs(1699) <= (inputs(51)) or (inputs(205));
    layer0_outputs(1700) <= not((inputs(196)) or (inputs(169)));
    layer0_outputs(1701) <= '1';
    layer0_outputs(1702) <= inputs(150);
    layer0_outputs(1703) <= (inputs(180)) and (inputs(64));
    layer0_outputs(1704) <= inputs(224);
    layer0_outputs(1705) <= (inputs(186)) and (inputs(210));
    layer0_outputs(1706) <= not((inputs(48)) and (inputs(73)));
    layer0_outputs(1707) <= not(inputs(84));
    layer0_outputs(1708) <= inputs(34);
    layer0_outputs(1709) <= '0';
    layer0_outputs(1710) <= '1';
    layer0_outputs(1711) <= '1';
    layer0_outputs(1712) <= (inputs(133)) and (inputs(240));
    layer0_outputs(1713) <= not((inputs(32)) or (inputs(73)));
    layer0_outputs(1714) <= (inputs(61)) or (inputs(63));
    layer0_outputs(1715) <= not(inputs(247));
    layer0_outputs(1716) <= not(inputs(143));
    layer0_outputs(1717) <= (inputs(195)) and not (inputs(88));
    layer0_outputs(1718) <= not(inputs(181));
    layer0_outputs(1719) <= not((inputs(219)) or (inputs(203)));
    layer0_outputs(1720) <= (inputs(31)) and (inputs(142));
    layer0_outputs(1721) <= '0';
    layer0_outputs(1722) <= not(inputs(101)) or (inputs(19));
    layer0_outputs(1723) <= (inputs(66)) and not (inputs(90));
    layer0_outputs(1724) <= not((inputs(7)) and (inputs(225)));
    layer0_outputs(1725) <= not((inputs(129)) or (inputs(116)));
    layer0_outputs(1726) <= not(inputs(98));
    layer0_outputs(1727) <= not(inputs(228));
    layer0_outputs(1728) <= '1';
    layer0_outputs(1729) <= not(inputs(85)) or (inputs(193));
    layer0_outputs(1730) <= '0';
    layer0_outputs(1731) <= not((inputs(192)) xor (inputs(192)));
    layer0_outputs(1732) <= not(inputs(201));
    layer0_outputs(1733) <= not(inputs(164)) or (inputs(33));
    layer0_outputs(1734) <= inputs(106);
    layer0_outputs(1735) <= '0';
    layer0_outputs(1736) <= not(inputs(130)) or (inputs(252));
    layer0_outputs(1737) <= not(inputs(223)) or (inputs(243));
    layer0_outputs(1738) <= '0';
    layer0_outputs(1739) <= not(inputs(45));
    layer0_outputs(1740) <= inputs(242);
    layer0_outputs(1741) <= '0';
    layer0_outputs(1742) <= (inputs(27)) and (inputs(66));
    layer0_outputs(1743) <= (inputs(223)) and (inputs(51));
    layer0_outputs(1744) <= (inputs(255)) xor (inputs(64));
    layer0_outputs(1745) <= not(inputs(228));
    layer0_outputs(1746) <= (inputs(58)) and (inputs(245));
    layer0_outputs(1747) <= (inputs(68)) and not (inputs(114));
    layer0_outputs(1748) <= not(inputs(179));
    layer0_outputs(1749) <= not(inputs(146)) or (inputs(251));
    layer0_outputs(1750) <= '1';
    layer0_outputs(1751) <= inputs(73);
    layer0_outputs(1752) <= not((inputs(189)) xor (inputs(254)));
    layer0_outputs(1753) <= '1';
    layer0_outputs(1754) <= inputs(109);
    layer0_outputs(1755) <= (inputs(119)) xor (inputs(117));
    layer0_outputs(1756) <= inputs(114);
    layer0_outputs(1757) <= '0';
    layer0_outputs(1758) <= inputs(181);
    layer0_outputs(1759) <= inputs(137);
    layer0_outputs(1760) <= not(inputs(250)) or (inputs(239));
    layer0_outputs(1761) <= inputs(153);
    layer0_outputs(1762) <= not(inputs(205)) or (inputs(14));
    layer0_outputs(1763) <= not(inputs(170));
    layer0_outputs(1764) <= not(inputs(143));
    layer0_outputs(1765) <= not(inputs(130));
    layer0_outputs(1766) <= '1';
    layer0_outputs(1767) <= not((inputs(163)) or (inputs(142)));
    layer0_outputs(1768) <= not(inputs(54));
    layer0_outputs(1769) <= inputs(227);
    layer0_outputs(1770) <= inputs(98);
    layer0_outputs(1771) <= not(inputs(22));
    layer0_outputs(1772) <= inputs(81);
    layer0_outputs(1773) <= not((inputs(42)) or (inputs(254)));
    layer0_outputs(1774) <= (inputs(237)) and (inputs(215));
    layer0_outputs(1775) <= inputs(176);
    layer0_outputs(1776) <= not(inputs(174));
    layer0_outputs(1777) <= '0';
    layer0_outputs(1778) <= not(inputs(179)) or (inputs(59));
    layer0_outputs(1779) <= inputs(149);
    layer0_outputs(1780) <= (inputs(161)) or (inputs(179));
    layer0_outputs(1781) <= '0';
    layer0_outputs(1782) <= '0';
    layer0_outputs(1783) <= (inputs(16)) and (inputs(166));
    layer0_outputs(1784) <= inputs(223);
    layer0_outputs(1785) <= inputs(173);
    layer0_outputs(1786) <= not(inputs(92)) or (inputs(100));
    layer0_outputs(1787) <= not((inputs(212)) or (inputs(204)));
    layer0_outputs(1788) <= (inputs(135)) and not (inputs(221));
    layer0_outputs(1789) <= (inputs(117)) and not (inputs(0));
    layer0_outputs(1790) <= not((inputs(134)) or (inputs(20)));
    layer0_outputs(1791) <= not(inputs(195));
    layer0_outputs(1792) <= not(inputs(66)) or (inputs(183));
    layer0_outputs(1793) <= (inputs(147)) or (inputs(149));
    layer0_outputs(1794) <= (inputs(86)) xor (inputs(159));
    layer0_outputs(1795) <= '1';
    layer0_outputs(1796) <= not(inputs(131)) or (inputs(138));
    layer0_outputs(1797) <= inputs(137);
    layer0_outputs(1798) <= '0';
    layer0_outputs(1799) <= not((inputs(220)) and (inputs(16)));
    layer0_outputs(1800) <= not(inputs(150)) or (inputs(141));
    layer0_outputs(1801) <= '0';
    layer0_outputs(1802) <= '0';
    layer0_outputs(1803) <= (inputs(232)) and not (inputs(1));
    layer0_outputs(1804) <= (inputs(39)) and not (inputs(192));
    layer0_outputs(1805) <= (inputs(19)) and not (inputs(53));
    layer0_outputs(1806) <= not((inputs(146)) or (inputs(171)));
    layer0_outputs(1807) <= '1';
    layer0_outputs(1808) <= not((inputs(128)) or (inputs(143)));
    layer0_outputs(1809) <= not((inputs(141)) and (inputs(211)));
    layer0_outputs(1810) <= (inputs(158)) or (inputs(196));
    layer0_outputs(1811) <= (inputs(225)) and (inputs(140));
    layer0_outputs(1812) <= (inputs(178)) and not (inputs(93));
    layer0_outputs(1813) <= not(inputs(169)) or (inputs(41));
    layer0_outputs(1814) <= not((inputs(139)) and (inputs(170)));
    layer0_outputs(1815) <= not((inputs(118)) or (inputs(234)));
    layer0_outputs(1816) <= '0';
    layer0_outputs(1817) <= inputs(13);
    layer0_outputs(1818) <= inputs(191);
    layer0_outputs(1819) <= not(inputs(45));
    layer0_outputs(1820) <= inputs(222);
    layer0_outputs(1821) <= not(inputs(147));
    layer0_outputs(1822) <= '1';
    layer0_outputs(1823) <= (inputs(147)) and not (inputs(154));
    layer0_outputs(1824) <= '0';
    layer0_outputs(1825) <= not(inputs(151));
    layer0_outputs(1826) <= inputs(103);
    layer0_outputs(1827) <= not((inputs(159)) and (inputs(120)));
    layer0_outputs(1828) <= not(inputs(2));
    layer0_outputs(1829) <= not(inputs(0)) or (inputs(222));
    layer0_outputs(1830) <= not(inputs(84)) or (inputs(49));
    layer0_outputs(1831) <= inputs(109);
    layer0_outputs(1832) <= not(inputs(81));
    layer0_outputs(1833) <= not(inputs(183));
    layer0_outputs(1834) <= inputs(136);
    layer0_outputs(1835) <= not((inputs(162)) and (inputs(223)));
    layer0_outputs(1836) <= not(inputs(24)) or (inputs(102));
    layer0_outputs(1837) <= (inputs(176)) and not (inputs(173));
    layer0_outputs(1838) <= not(inputs(149));
    layer0_outputs(1839) <= inputs(146);
    layer0_outputs(1840) <= '0';
    layer0_outputs(1841) <= '1';
    layer0_outputs(1842) <= not(inputs(248)) or (inputs(2));
    layer0_outputs(1843) <= (inputs(165)) and (inputs(4));
    layer0_outputs(1844) <= '0';
    layer0_outputs(1845) <= not(inputs(176)) or (inputs(22));
    layer0_outputs(1846) <= inputs(163);
    layer0_outputs(1847) <= inputs(220);
    layer0_outputs(1848) <= (inputs(85)) and not (inputs(159));
    layer0_outputs(1849) <= '1';
    layer0_outputs(1850) <= '0';
    layer0_outputs(1851) <= not(inputs(105)) or (inputs(213));
    layer0_outputs(1852) <= (inputs(123)) and not (inputs(198));
    layer0_outputs(1853) <= not(inputs(189)) or (inputs(162));
    layer0_outputs(1854) <= not(inputs(119));
    layer0_outputs(1855) <= (inputs(60)) and not (inputs(15));
    layer0_outputs(1856) <= (inputs(116)) or (inputs(45));
    layer0_outputs(1857) <= (inputs(157)) and not (inputs(168));
    layer0_outputs(1858) <= '0';
    layer0_outputs(1859) <= '0';
    layer0_outputs(1860) <= not(inputs(90));
    layer0_outputs(1861) <= '1';
    layer0_outputs(1862) <= not(inputs(166));
    layer0_outputs(1863) <= '1';
    layer0_outputs(1864) <= (inputs(180)) and not (inputs(241));
    layer0_outputs(1865) <= not(inputs(92)) or (inputs(30));
    layer0_outputs(1866) <= not(inputs(79));
    layer0_outputs(1867) <= '1';
    layer0_outputs(1868) <= not((inputs(211)) or (inputs(225)));
    layer0_outputs(1869) <= inputs(121);
    layer0_outputs(1870) <= not(inputs(233));
    layer0_outputs(1871) <= not(inputs(56));
    layer0_outputs(1872) <= (inputs(148)) or (inputs(98));
    layer0_outputs(1873) <= '0';
    layer0_outputs(1874) <= inputs(3);
    layer0_outputs(1875) <= (inputs(62)) and not (inputs(109));
    layer0_outputs(1876) <= (inputs(87)) xor (inputs(57));
    layer0_outputs(1877) <= (inputs(86)) and not (inputs(253));
    layer0_outputs(1878) <= not((inputs(83)) or (inputs(112)));
    layer0_outputs(1879) <= (inputs(176)) or (inputs(64));
    layer0_outputs(1880) <= '1';
    layer0_outputs(1881) <= '0';
    layer0_outputs(1882) <= not(inputs(117));
    layer0_outputs(1883) <= (inputs(92)) and not (inputs(188));
    layer0_outputs(1884) <= '0';
    layer0_outputs(1885) <= (inputs(77)) and (inputs(49));
    layer0_outputs(1886) <= (inputs(22)) xor (inputs(158));
    layer0_outputs(1887) <= '0';
    layer0_outputs(1888) <= not((inputs(166)) or (inputs(152)));
    layer0_outputs(1889) <= (inputs(195)) xor (inputs(14));
    layer0_outputs(1890) <= not(inputs(0)) or (inputs(49));
    layer0_outputs(1891) <= inputs(145);
    layer0_outputs(1892) <= '1';
    layer0_outputs(1893) <= not((inputs(113)) or (inputs(68)));
    layer0_outputs(1894) <= not((inputs(182)) or (inputs(221)));
    layer0_outputs(1895) <= (inputs(120)) and not (inputs(36));
    layer0_outputs(1896) <= inputs(100);
    layer0_outputs(1897) <= '1';
    layer0_outputs(1898) <= inputs(232);
    layer0_outputs(1899) <= not(inputs(127)) or (inputs(168));
    layer0_outputs(1900) <= '0';
    layer0_outputs(1901) <= '1';
    layer0_outputs(1902) <= inputs(84);
    layer0_outputs(1903) <= inputs(243);
    layer0_outputs(1904) <= not(inputs(190)) or (inputs(19));
    layer0_outputs(1905) <= '1';
    layer0_outputs(1906) <= inputs(177);
    layer0_outputs(1907) <= '0';
    layer0_outputs(1908) <= not(inputs(60)) or (inputs(205));
    layer0_outputs(1909) <= inputs(105);
    layer0_outputs(1910) <= not(inputs(207));
    layer0_outputs(1911) <= '1';
    layer0_outputs(1912) <= not((inputs(52)) or (inputs(131)));
    layer0_outputs(1913) <= '1';
    layer0_outputs(1914) <= not(inputs(79));
    layer0_outputs(1915) <= (inputs(71)) or (inputs(163));
    layer0_outputs(1916) <= '1';
    layer0_outputs(1917) <= not(inputs(172));
    layer0_outputs(1918) <= (inputs(207)) and (inputs(152));
    layer0_outputs(1919) <= (inputs(191)) and not (inputs(245));
    layer0_outputs(1920) <= '1';
    layer0_outputs(1921) <= '0';
    layer0_outputs(1922) <= not((inputs(220)) or (inputs(137)));
    layer0_outputs(1923) <= (inputs(18)) and not (inputs(203));
    layer0_outputs(1924) <= '0';
    layer0_outputs(1925) <= not((inputs(117)) or (inputs(128)));
    layer0_outputs(1926) <= not(inputs(161));
    layer0_outputs(1927) <= '1';
    layer0_outputs(1928) <= inputs(110);
    layer0_outputs(1929) <= '0';
    layer0_outputs(1930) <= inputs(124);
    layer0_outputs(1931) <= (inputs(46)) and (inputs(191));
    layer0_outputs(1932) <= not((inputs(92)) or (inputs(78)));
    layer0_outputs(1933) <= (inputs(35)) and not (inputs(57));
    layer0_outputs(1934) <= '1';
    layer0_outputs(1935) <= not(inputs(148)) or (inputs(13));
    layer0_outputs(1936) <= not((inputs(68)) or (inputs(126)));
    layer0_outputs(1937) <= (inputs(24)) and (inputs(114));
    layer0_outputs(1938) <= (inputs(89)) and (inputs(27));
    layer0_outputs(1939) <= not((inputs(109)) or (inputs(140)));
    layer0_outputs(1940) <= '1';
    layer0_outputs(1941) <= (inputs(163)) and not (inputs(39));
    layer0_outputs(1942) <= not(inputs(233)) or (inputs(112));
    layer0_outputs(1943) <= not((inputs(238)) and (inputs(235)));
    layer0_outputs(1944) <= inputs(173);
    layer0_outputs(1945) <= '1';
    layer0_outputs(1946) <= '1';
    layer0_outputs(1947) <= '0';
    layer0_outputs(1948) <= not(inputs(116));
    layer0_outputs(1949) <= inputs(112);
    layer0_outputs(1950) <= not(inputs(61));
    layer0_outputs(1951) <= '0';
    layer0_outputs(1952) <= inputs(214);
    layer0_outputs(1953) <= '1';
    layer0_outputs(1954) <= '0';
    layer0_outputs(1955) <= (inputs(254)) or (inputs(122));
    layer0_outputs(1956) <= not(inputs(7)) or (inputs(29));
    layer0_outputs(1957) <= inputs(164);
    layer0_outputs(1958) <= not((inputs(191)) or (inputs(206)));
    layer0_outputs(1959) <= not((inputs(188)) or (inputs(183)));
    layer0_outputs(1960) <= inputs(247);
    layer0_outputs(1961) <= (inputs(84)) and not (inputs(177));
    layer0_outputs(1962) <= inputs(155);
    layer0_outputs(1963) <= '1';
    layer0_outputs(1964) <= '1';
    layer0_outputs(1965) <= not(inputs(72)) or (inputs(251));
    layer0_outputs(1966) <= inputs(100);
    layer0_outputs(1967) <= not(inputs(173));
    layer0_outputs(1968) <= not((inputs(87)) and (inputs(143)));
    layer0_outputs(1969) <= not((inputs(185)) or (inputs(174)));
    layer0_outputs(1970) <= not(inputs(8));
    layer0_outputs(1971) <= not(inputs(119));
    layer0_outputs(1972) <= inputs(250);
    layer0_outputs(1973) <= not(inputs(34)) or (inputs(252));
    layer0_outputs(1974) <= (inputs(61)) and (inputs(92));
    layer0_outputs(1975) <= (inputs(132)) or (inputs(69));
    layer0_outputs(1976) <= '0';
    layer0_outputs(1977) <= (inputs(48)) and not (inputs(197));
    layer0_outputs(1978) <= '0';
    layer0_outputs(1979) <= not((inputs(126)) or (inputs(196)));
    layer0_outputs(1980) <= '1';
    layer0_outputs(1981) <= (inputs(46)) or (inputs(211));
    layer0_outputs(1982) <= '1';
    layer0_outputs(1983) <= not(inputs(83));
    layer0_outputs(1984) <= '0';
    layer0_outputs(1985) <= (inputs(25)) or (inputs(17));
    layer0_outputs(1986) <= inputs(166);
    layer0_outputs(1987) <= (inputs(233)) and not (inputs(81));
    layer0_outputs(1988) <= inputs(84);
    layer0_outputs(1989) <= not(inputs(37)) or (inputs(139));
    layer0_outputs(1990) <= not((inputs(173)) or (inputs(94)));
    layer0_outputs(1991) <= (inputs(78)) and not (inputs(37));
    layer0_outputs(1992) <= not((inputs(176)) or (inputs(125)));
    layer0_outputs(1993) <= not((inputs(85)) and (inputs(55)));
    layer0_outputs(1994) <= '1';
    layer0_outputs(1995) <= not(inputs(94));
    layer0_outputs(1996) <= (inputs(51)) and (inputs(251));
    layer0_outputs(1997) <= not(inputs(99));
    layer0_outputs(1998) <= inputs(36);
    layer0_outputs(1999) <= not((inputs(1)) or (inputs(235)));
    layer0_outputs(2000) <= not(inputs(174));
    layer0_outputs(2001) <= not((inputs(16)) or (inputs(217)));
    layer0_outputs(2002) <= not((inputs(62)) and (inputs(80)));
    layer0_outputs(2003) <= (inputs(106)) and not (inputs(13));
    layer0_outputs(2004) <= (inputs(21)) or (inputs(18));
    layer0_outputs(2005) <= (inputs(49)) or (inputs(123));
    layer0_outputs(2006) <= not((inputs(245)) and (inputs(0)));
    layer0_outputs(2007) <= inputs(167);
    layer0_outputs(2008) <= inputs(207);
    layer0_outputs(2009) <= '1';
    layer0_outputs(2010) <= (inputs(157)) or (inputs(133));
    layer0_outputs(2011) <= '1';
    layer0_outputs(2012) <= '1';
    layer0_outputs(2013) <= inputs(93);
    layer0_outputs(2014) <= '0';
    layer0_outputs(2015) <= '0';
    layer0_outputs(2016) <= not((inputs(43)) and (inputs(56)));
    layer0_outputs(2017) <= not((inputs(207)) or (inputs(220)));
    layer0_outputs(2018) <= not((inputs(63)) and (inputs(111)));
    layer0_outputs(2019) <= not(inputs(194));
    layer0_outputs(2020) <= (inputs(87)) and not (inputs(149));
    layer0_outputs(2021) <= not(inputs(134));
    layer0_outputs(2022) <= not(inputs(216));
    layer0_outputs(2023) <= (inputs(236)) or (inputs(235));
    layer0_outputs(2024) <= not(inputs(163));
    layer0_outputs(2025) <= not(inputs(127)) or (inputs(169));
    layer0_outputs(2026) <= not(inputs(2));
    layer0_outputs(2027) <= not(inputs(235)) or (inputs(157));
    layer0_outputs(2028) <= '1';
    layer0_outputs(2029) <= not(inputs(160));
    layer0_outputs(2030) <= not(inputs(139)) or (inputs(23));
    layer0_outputs(2031) <= '0';
    layer0_outputs(2032) <= inputs(194);
    layer0_outputs(2033) <= '0';
    layer0_outputs(2034) <= inputs(143);
    layer0_outputs(2035) <= inputs(94);
    layer0_outputs(2036) <= not((inputs(169)) or (inputs(55)));
    layer0_outputs(2037) <= (inputs(193)) or (inputs(114));
    layer0_outputs(2038) <= '1';
    layer0_outputs(2039) <= '1';
    layer0_outputs(2040) <= not(inputs(10)) or (inputs(250));
    layer0_outputs(2041) <= inputs(224);
    layer0_outputs(2042) <= not((inputs(2)) or (inputs(90)));
    layer0_outputs(2043) <= not(inputs(177)) or (inputs(139));
    layer0_outputs(2044) <= not(inputs(159));
    layer0_outputs(2045) <= (inputs(18)) and not (inputs(126));
    layer0_outputs(2046) <= not(inputs(60)) or (inputs(49));
    layer0_outputs(2047) <= not((inputs(60)) and (inputs(126)));
    layer0_outputs(2048) <= not(inputs(32));
    layer0_outputs(2049) <= not((inputs(254)) and (inputs(213)));
    layer0_outputs(2050) <= (inputs(191)) and not (inputs(72));
    layer0_outputs(2051) <= inputs(69);
    layer0_outputs(2052) <= not(inputs(155));
    layer0_outputs(2053) <= '0';
    layer0_outputs(2054) <= not(inputs(14));
    layer0_outputs(2055) <= (inputs(132)) and not (inputs(237));
    layer0_outputs(2056) <= not((inputs(42)) or (inputs(206)));
    layer0_outputs(2057) <= not(inputs(66));
    layer0_outputs(2058) <= not(inputs(119));
    layer0_outputs(2059) <= '0';
    layer0_outputs(2060) <= (inputs(140)) and not (inputs(215));
    layer0_outputs(2061) <= '1';
    layer0_outputs(2062) <= not(inputs(1));
    layer0_outputs(2063) <= inputs(32);
    layer0_outputs(2064) <= not(inputs(177));
    layer0_outputs(2065) <= not(inputs(39)) or (inputs(173));
    layer0_outputs(2066) <= inputs(105);
    layer0_outputs(2067) <= (inputs(149)) or (inputs(81));
    layer0_outputs(2068) <= (inputs(177)) or (inputs(233));
    layer0_outputs(2069) <= not(inputs(100));
    layer0_outputs(2070) <= (inputs(167)) or (inputs(135));
    layer0_outputs(2071) <= inputs(164);
    layer0_outputs(2072) <= not(inputs(97)) or (inputs(186));
    layer0_outputs(2073) <= not(inputs(74)) or (inputs(244));
    layer0_outputs(2074) <= not(inputs(140)) or (inputs(87));
    layer0_outputs(2075) <= '1';
    layer0_outputs(2076) <= not(inputs(25));
    layer0_outputs(2077) <= not(inputs(43));
    layer0_outputs(2078) <= inputs(210);
    layer0_outputs(2079) <= (inputs(100)) and not (inputs(48));
    layer0_outputs(2080) <= '0';
    layer0_outputs(2081) <= not(inputs(181));
    layer0_outputs(2082) <= not(inputs(185));
    layer0_outputs(2083) <= not(inputs(219));
    layer0_outputs(2084) <= not((inputs(203)) and (inputs(183)));
    layer0_outputs(2085) <= not((inputs(96)) or (inputs(152)));
    layer0_outputs(2086) <= '1';
    layer0_outputs(2087) <= not(inputs(19));
    layer0_outputs(2088) <= not(inputs(228)) or (inputs(51));
    layer0_outputs(2089) <= '1';
    layer0_outputs(2090) <= '1';
    layer0_outputs(2091) <= inputs(116);
    layer0_outputs(2092) <= not(inputs(107)) or (inputs(194));
    layer0_outputs(2093) <= (inputs(76)) and not (inputs(194));
    layer0_outputs(2094) <= not((inputs(164)) and (inputs(242)));
    layer0_outputs(2095) <= (inputs(19)) and (inputs(242));
    layer0_outputs(2096) <= not(inputs(183)) or (inputs(30));
    layer0_outputs(2097) <= inputs(235);
    layer0_outputs(2098) <= (inputs(125)) or (inputs(129));
    layer0_outputs(2099) <= not(inputs(174));
    layer0_outputs(2100) <= '0';
    layer0_outputs(2101) <= not((inputs(253)) or (inputs(153)));
    layer0_outputs(2102) <= '1';
    layer0_outputs(2103) <= '0';
    layer0_outputs(2104) <= not((inputs(167)) or (inputs(147)));
    layer0_outputs(2105) <= inputs(167);
    layer0_outputs(2106) <= inputs(249);
    layer0_outputs(2107) <= (inputs(0)) xor (inputs(3));
    layer0_outputs(2108) <= (inputs(245)) or (inputs(17));
    layer0_outputs(2109) <= not(inputs(203)) or (inputs(153));
    layer0_outputs(2110) <= (inputs(202)) or (inputs(162));
    layer0_outputs(2111) <= not(inputs(86));
    layer0_outputs(2112) <= not(inputs(249)) or (inputs(184));
    layer0_outputs(2113) <= inputs(82);
    layer0_outputs(2114) <= '1';
    layer0_outputs(2115) <= not(inputs(103));
    layer0_outputs(2116) <= not(inputs(90));
    layer0_outputs(2117) <= (inputs(252)) and (inputs(15));
    layer0_outputs(2118) <= not((inputs(231)) or (inputs(144)));
    layer0_outputs(2119) <= not(inputs(47));
    layer0_outputs(2120) <= inputs(30);
    layer0_outputs(2121) <= '0';
    layer0_outputs(2122) <= '0';
    layer0_outputs(2123) <= not(inputs(99)) or (inputs(190));
    layer0_outputs(2124) <= not(inputs(233));
    layer0_outputs(2125) <= (inputs(65)) and not (inputs(225));
    layer0_outputs(2126) <= (inputs(15)) xor (inputs(178));
    layer0_outputs(2127) <= not((inputs(137)) or (inputs(5)));
    layer0_outputs(2128) <= '0';
    layer0_outputs(2129) <= '0';
    layer0_outputs(2130) <= inputs(211);
    layer0_outputs(2131) <= not((inputs(120)) or (inputs(17)));
    layer0_outputs(2132) <= inputs(177);
    layer0_outputs(2133) <= not(inputs(161)) or (inputs(158));
    layer0_outputs(2134) <= '1';
    layer0_outputs(2135) <= (inputs(184)) and not (inputs(255));
    layer0_outputs(2136) <= not(inputs(3));
    layer0_outputs(2137) <= '0';
    layer0_outputs(2138) <= inputs(100);
    layer0_outputs(2139) <= '0';
    layer0_outputs(2140) <= (inputs(221)) or (inputs(164));
    layer0_outputs(2141) <= not(inputs(7));
    layer0_outputs(2142) <= (inputs(205)) and not (inputs(23));
    layer0_outputs(2143) <= '1';
    layer0_outputs(2144) <= (inputs(181)) and not (inputs(79));
    layer0_outputs(2145) <= '0';
    layer0_outputs(2146) <= not(inputs(138));
    layer0_outputs(2147) <= inputs(210);
    layer0_outputs(2148) <= (inputs(120)) or (inputs(247));
    layer0_outputs(2149) <= inputs(151);
    layer0_outputs(2150) <= inputs(127);
    layer0_outputs(2151) <= not((inputs(160)) xor (inputs(131)));
    layer0_outputs(2152) <= not(inputs(87));
    layer0_outputs(2153) <= (inputs(145)) or (inputs(190));
    layer0_outputs(2154) <= not(inputs(205)) or (inputs(110));
    layer0_outputs(2155) <= '1';
    layer0_outputs(2156) <= (inputs(213)) and not (inputs(11));
    layer0_outputs(2157) <= '1';
    layer0_outputs(2158) <= '0';
    layer0_outputs(2159) <= '0';
    layer0_outputs(2160) <= inputs(67);
    layer0_outputs(2161) <= not(inputs(151)) or (inputs(67));
    layer0_outputs(2162) <= inputs(35);
    layer0_outputs(2163) <= inputs(72);
    layer0_outputs(2164) <= '0';
    layer0_outputs(2165) <= (inputs(127)) xor (inputs(130));
    layer0_outputs(2166) <= not((inputs(172)) or (inputs(1)));
    layer0_outputs(2167) <= (inputs(122)) xor (inputs(81));
    layer0_outputs(2168) <= not(inputs(152)) or (inputs(28));
    layer0_outputs(2169) <= not(inputs(196)) or (inputs(111));
    layer0_outputs(2170) <= not(inputs(114)) or (inputs(5));
    layer0_outputs(2171) <= '1';
    layer0_outputs(2172) <= not((inputs(53)) and (inputs(106)));
    layer0_outputs(2173) <= '0';
    layer0_outputs(2174) <= (inputs(61)) or (inputs(163));
    layer0_outputs(2175) <= (inputs(206)) or (inputs(167));
    layer0_outputs(2176) <= not(inputs(183));
    layer0_outputs(2177) <= (inputs(137)) and not (inputs(143));
    layer0_outputs(2178) <= not((inputs(202)) and (inputs(29)));
    layer0_outputs(2179) <= not(inputs(169));
    layer0_outputs(2180) <= not((inputs(237)) or (inputs(17)));
    layer0_outputs(2181) <= not((inputs(35)) or (inputs(3)));
    layer0_outputs(2182) <= inputs(230);
    layer0_outputs(2183) <= not(inputs(103));
    layer0_outputs(2184) <= '1';
    layer0_outputs(2185) <= inputs(161);
    layer0_outputs(2186) <= (inputs(164)) or (inputs(113));
    layer0_outputs(2187) <= (inputs(3)) or (inputs(109));
    layer0_outputs(2188) <= not(inputs(135));
    layer0_outputs(2189) <= not(inputs(9));
    layer0_outputs(2190) <= inputs(68);
    layer0_outputs(2191) <= inputs(67);
    layer0_outputs(2192) <= not(inputs(79)) or (inputs(242));
    layer0_outputs(2193) <= not(inputs(1));
    layer0_outputs(2194) <= '0';
    layer0_outputs(2195) <= (inputs(145)) and not (inputs(137));
    layer0_outputs(2196) <= '1';
    layer0_outputs(2197) <= not(inputs(118));
    layer0_outputs(2198) <= (inputs(159)) and not (inputs(249));
    layer0_outputs(2199) <= (inputs(48)) and not (inputs(108));
    layer0_outputs(2200) <= (inputs(113)) or (inputs(139));
    layer0_outputs(2201) <= '0';
    layer0_outputs(2202) <= not(inputs(67));
    layer0_outputs(2203) <= not(inputs(7)) or (inputs(87));
    layer0_outputs(2204) <= inputs(236);
    layer0_outputs(2205) <= (inputs(239)) xor (inputs(175));
    layer0_outputs(2206) <= (inputs(244)) or (inputs(53));
    layer0_outputs(2207) <= not(inputs(75));
    layer0_outputs(2208) <= '1';
    layer0_outputs(2209) <= inputs(132);
    layer0_outputs(2210) <= (inputs(221)) and not (inputs(153));
    layer0_outputs(2211) <= inputs(166);
    layer0_outputs(2212) <= not(inputs(10)) or (inputs(209));
    layer0_outputs(2213) <= '1';
    layer0_outputs(2214) <= '1';
    layer0_outputs(2215) <= not(inputs(11)) or (inputs(95));
    layer0_outputs(2216) <= (inputs(145)) and (inputs(211));
    layer0_outputs(2217) <= (inputs(119)) xor (inputs(151));
    layer0_outputs(2218) <= (inputs(83)) and not (inputs(186));
    layer0_outputs(2219) <= not(inputs(127)) or (inputs(1));
    layer0_outputs(2220) <= '0';
    layer0_outputs(2221) <= not(inputs(247)) or (inputs(164));
    layer0_outputs(2222) <= not(inputs(33));
    layer0_outputs(2223) <= inputs(132);
    layer0_outputs(2224) <= not((inputs(202)) or (inputs(205)));
    layer0_outputs(2225) <= inputs(26);
    layer0_outputs(2226) <= (inputs(107)) and not (inputs(153));
    layer0_outputs(2227) <= (inputs(24)) or (inputs(47));
    layer0_outputs(2228) <= not(inputs(112));
    layer0_outputs(2229) <= inputs(138);
    layer0_outputs(2230) <= '1';
    layer0_outputs(2231) <= not((inputs(39)) and (inputs(45)));
    layer0_outputs(2232) <= (inputs(143)) or (inputs(94));
    layer0_outputs(2233) <= not(inputs(137));
    layer0_outputs(2234) <= not((inputs(129)) or (inputs(36)));
    layer0_outputs(2235) <= not(inputs(98));
    layer0_outputs(2236) <= inputs(157);
    layer0_outputs(2237) <= not((inputs(130)) and (inputs(77)));
    layer0_outputs(2238) <= not(inputs(84));
    layer0_outputs(2239) <= (inputs(228)) and not (inputs(182));
    layer0_outputs(2240) <= (inputs(127)) and not (inputs(220));
    layer0_outputs(2241) <= inputs(251);
    layer0_outputs(2242) <= '1';
    layer0_outputs(2243) <= (inputs(115)) or (inputs(117));
    layer0_outputs(2244) <= (inputs(103)) or (inputs(206));
    layer0_outputs(2245) <= not(inputs(86)) or (inputs(80));
    layer0_outputs(2246) <= not((inputs(96)) or (inputs(204)));
    layer0_outputs(2247) <= not(inputs(175));
    layer0_outputs(2248) <= (inputs(222)) xor (inputs(192));
    layer0_outputs(2249) <= '0';
    layer0_outputs(2250) <= '0';
    layer0_outputs(2251) <= not(inputs(255));
    layer0_outputs(2252) <= not(inputs(106)) or (inputs(75));
    layer0_outputs(2253) <= (inputs(150)) or (inputs(75));
    layer0_outputs(2254) <= not((inputs(1)) and (inputs(86)));
    layer0_outputs(2255) <= (inputs(39)) and not (inputs(183));
    layer0_outputs(2256) <= (inputs(186)) or (inputs(90));
    layer0_outputs(2257) <= not(inputs(154));
    layer0_outputs(2258) <= '1';
    layer0_outputs(2259) <= (inputs(30)) and (inputs(188));
    layer0_outputs(2260) <= inputs(70);
    layer0_outputs(2261) <= '0';
    layer0_outputs(2262) <= '0';
    layer0_outputs(2263) <= (inputs(82)) or (inputs(131));
    layer0_outputs(2264) <= (inputs(97)) and not (inputs(119));
    layer0_outputs(2265) <= '1';
    layer0_outputs(2266) <= (inputs(37)) or (inputs(171));
    layer0_outputs(2267) <= '0';
    layer0_outputs(2268) <= not(inputs(75));
    layer0_outputs(2269) <= (inputs(188)) xor (inputs(253));
    layer0_outputs(2270) <= not(inputs(192)) or (inputs(251));
    layer0_outputs(2271) <= (inputs(227)) and not (inputs(144));
    layer0_outputs(2272) <= '1';
    layer0_outputs(2273) <= '1';
    layer0_outputs(2274) <= not(inputs(91)) or (inputs(29));
    layer0_outputs(2275) <= '0';
    layer0_outputs(2276) <= (inputs(200)) and (inputs(115));
    layer0_outputs(2277) <= (inputs(15)) xor (inputs(79));
    layer0_outputs(2278) <= (inputs(89)) or (inputs(27));
    layer0_outputs(2279) <= (inputs(247)) or (inputs(72));
    layer0_outputs(2280) <= not((inputs(2)) or (inputs(224)));
    layer0_outputs(2281) <= (inputs(115)) and not (inputs(254));
    layer0_outputs(2282) <= '1';
    layer0_outputs(2283) <= not(inputs(109));
    layer0_outputs(2284) <= '1';
    layer0_outputs(2285) <= (inputs(50)) and not (inputs(138));
    layer0_outputs(2286) <= (inputs(170)) or (inputs(253));
    layer0_outputs(2287) <= (inputs(76)) and (inputs(55));
    layer0_outputs(2288) <= (inputs(156)) or (inputs(158));
    layer0_outputs(2289) <= not((inputs(220)) and (inputs(70)));
    layer0_outputs(2290) <= '0';
    layer0_outputs(2291) <= '1';
    layer0_outputs(2292) <= not(inputs(242)) or (inputs(57));
    layer0_outputs(2293) <= not((inputs(193)) xor (inputs(83)));
    layer0_outputs(2294) <= (inputs(31)) and not (inputs(229));
    layer0_outputs(2295) <= not(inputs(123));
    layer0_outputs(2296) <= '0';
    layer0_outputs(2297) <= not((inputs(245)) or (inputs(213)));
    layer0_outputs(2298) <= (inputs(119)) and not (inputs(63));
    layer0_outputs(2299) <= (inputs(205)) and (inputs(203));
    layer0_outputs(2300) <= not(inputs(217)) or (inputs(64));
    layer0_outputs(2301) <= not(inputs(249));
    layer0_outputs(2302) <= not((inputs(152)) or (inputs(151)));
    layer0_outputs(2303) <= not(inputs(192));
    layer0_outputs(2304) <= not((inputs(49)) xor (inputs(45)));
    layer0_outputs(2305) <= not(inputs(154));
    layer0_outputs(2306) <= not((inputs(12)) and (inputs(175)));
    layer0_outputs(2307) <= not(inputs(106)) or (inputs(216));
    layer0_outputs(2308) <= not(inputs(227));
    layer0_outputs(2309) <= '0';
    layer0_outputs(2310) <= not(inputs(6));
    layer0_outputs(2311) <= '0';
    layer0_outputs(2312) <= not((inputs(211)) or (inputs(200)));
    layer0_outputs(2313) <= not(inputs(47));
    layer0_outputs(2314) <= (inputs(104)) and not (inputs(139));
    layer0_outputs(2315) <= inputs(151);
    layer0_outputs(2316) <= (inputs(209)) and (inputs(219));
    layer0_outputs(2317) <= '1';
    layer0_outputs(2318) <= (inputs(248)) or (inputs(229));
    layer0_outputs(2319) <= inputs(23);
    layer0_outputs(2320) <= not(inputs(197));
    layer0_outputs(2321) <= '0';
    layer0_outputs(2322) <= '0';
    layer0_outputs(2323) <= not((inputs(198)) and (inputs(246)));
    layer0_outputs(2324) <= inputs(240);
    layer0_outputs(2325) <= '0';
    layer0_outputs(2326) <= (inputs(72)) and not (inputs(28));
    layer0_outputs(2327) <= '0';
    layer0_outputs(2328) <= (inputs(231)) or (inputs(213));
    layer0_outputs(2329) <= not(inputs(23));
    layer0_outputs(2330) <= not(inputs(3)) or (inputs(120));
    layer0_outputs(2331) <= not(inputs(14));
    layer0_outputs(2332) <= inputs(228);
    layer0_outputs(2333) <= not(inputs(59)) or (inputs(205));
    layer0_outputs(2334) <= not((inputs(120)) and (inputs(101)));
    layer0_outputs(2335) <= (inputs(32)) and (inputs(133));
    layer0_outputs(2336) <= '0';
    layer0_outputs(2337) <= (inputs(147)) or (inputs(88));
    layer0_outputs(2338) <= not(inputs(28));
    layer0_outputs(2339) <= not((inputs(57)) and (inputs(96)));
    layer0_outputs(2340) <= (inputs(100)) and (inputs(106));
    layer0_outputs(2341) <= inputs(91);
    layer0_outputs(2342) <= inputs(129);
    layer0_outputs(2343) <= '0';
    layer0_outputs(2344) <= '1';
    layer0_outputs(2345) <= '0';
    layer0_outputs(2346) <= not((inputs(204)) and (inputs(136)));
    layer0_outputs(2347) <= not(inputs(86));
    layer0_outputs(2348) <= '1';
    layer0_outputs(2349) <= (inputs(117)) or (inputs(66));
    layer0_outputs(2350) <= not(inputs(254)) or (inputs(203));
    layer0_outputs(2351) <= not((inputs(88)) or (inputs(85)));
    layer0_outputs(2352) <= not((inputs(176)) or (inputs(80)));
    layer0_outputs(2353) <= inputs(56);
    layer0_outputs(2354) <= not(inputs(195)) or (inputs(45));
    layer0_outputs(2355) <= '0';
    layer0_outputs(2356) <= (inputs(147)) and not (inputs(49));
    layer0_outputs(2357) <= '1';
    layer0_outputs(2358) <= not(inputs(255)) or (inputs(140));
    layer0_outputs(2359) <= (inputs(38)) or (inputs(178));
    layer0_outputs(2360) <= inputs(23);
    layer0_outputs(2361) <= (inputs(240)) and (inputs(103));
    layer0_outputs(2362) <= not((inputs(53)) or (inputs(98)));
    layer0_outputs(2363) <= not(inputs(209));
    layer0_outputs(2364) <= '0';
    layer0_outputs(2365) <= not(inputs(136)) or (inputs(163));
    layer0_outputs(2366) <= not(inputs(211)) or (inputs(61));
    layer0_outputs(2367) <= not(inputs(221));
    layer0_outputs(2368) <= inputs(246);
    layer0_outputs(2369) <= '0';
    layer0_outputs(2370) <= inputs(144);
    layer0_outputs(2371) <= '1';
    layer0_outputs(2372) <= inputs(222);
    layer0_outputs(2373) <= not(inputs(119)) or (inputs(49));
    layer0_outputs(2374) <= (inputs(71)) or (inputs(164));
    layer0_outputs(2375) <= not((inputs(223)) xor (inputs(190)));
    layer0_outputs(2376) <= not(inputs(106));
    layer0_outputs(2377) <= (inputs(133)) or (inputs(174));
    layer0_outputs(2378) <= '0';
    layer0_outputs(2379) <= not((inputs(31)) and (inputs(20)));
    layer0_outputs(2380) <= '0';
    layer0_outputs(2381) <= (inputs(211)) and not (inputs(195));
    layer0_outputs(2382) <= not(inputs(193)) or (inputs(160));
    layer0_outputs(2383) <= not(inputs(190));
    layer0_outputs(2384) <= inputs(204);
    layer0_outputs(2385) <= inputs(209);
    layer0_outputs(2386) <= (inputs(172)) and (inputs(247));
    layer0_outputs(2387) <= (inputs(7)) or (inputs(188));
    layer0_outputs(2388) <= inputs(0);
    layer0_outputs(2389) <= not(inputs(126));
    layer0_outputs(2390) <= not(inputs(145));
    layer0_outputs(2391) <= '1';
    layer0_outputs(2392) <= (inputs(85)) or (inputs(145));
    layer0_outputs(2393) <= not(inputs(204)) or (inputs(64));
    layer0_outputs(2394) <= '0';
    layer0_outputs(2395) <= '1';
    layer0_outputs(2396) <= not(inputs(177));
    layer0_outputs(2397) <= '1';
    layer0_outputs(2398) <= '0';
    layer0_outputs(2399) <= (inputs(123)) and not (inputs(245));
    layer0_outputs(2400) <= inputs(21);
    layer0_outputs(2401) <= not(inputs(192)) or (inputs(153));
    layer0_outputs(2402) <= (inputs(43)) and not (inputs(25));
    layer0_outputs(2403) <= (inputs(192)) and (inputs(1));
    layer0_outputs(2404) <= (inputs(216)) and (inputs(251));
    layer0_outputs(2405) <= (inputs(180)) and (inputs(93));
    layer0_outputs(2406) <= '0';
    layer0_outputs(2407) <= '1';
    layer0_outputs(2408) <= '1';
    layer0_outputs(2409) <= not(inputs(218)) or (inputs(169));
    layer0_outputs(2410) <= inputs(18);
    layer0_outputs(2411) <= not(inputs(228));
    layer0_outputs(2412) <= not((inputs(91)) or (inputs(239)));
    layer0_outputs(2413) <= not(inputs(77)) or (inputs(66));
    layer0_outputs(2414) <= inputs(232);
    layer0_outputs(2415) <= not((inputs(35)) or (inputs(51)));
    layer0_outputs(2416) <= not(inputs(154));
    layer0_outputs(2417) <= '1';
    layer0_outputs(2418) <= inputs(18);
    layer0_outputs(2419) <= inputs(25);
    layer0_outputs(2420) <= (inputs(99)) or (inputs(129));
    layer0_outputs(2421) <= not((inputs(108)) and (inputs(124)));
    layer0_outputs(2422) <= (inputs(51)) and not (inputs(116));
    layer0_outputs(2423) <= not(inputs(199));
    layer0_outputs(2424) <= '0';
    layer0_outputs(2425) <= '1';
    layer0_outputs(2426) <= '1';
    layer0_outputs(2427) <= inputs(192);
    layer0_outputs(2428) <= not(inputs(110));
    layer0_outputs(2429) <= not(inputs(129)) or (inputs(49));
    layer0_outputs(2430) <= not((inputs(249)) or (inputs(194)));
    layer0_outputs(2431) <= not(inputs(153)) or (inputs(12));
    layer0_outputs(2432) <= not((inputs(81)) or (inputs(108)));
    layer0_outputs(2433) <= '1';
    layer0_outputs(2434) <= inputs(207);
    layer0_outputs(2435) <= inputs(234);
    layer0_outputs(2436) <= not(inputs(78));
    layer0_outputs(2437) <= '0';
    layer0_outputs(2438) <= not((inputs(53)) or (inputs(64)));
    layer0_outputs(2439) <= not((inputs(73)) and (inputs(21)));
    layer0_outputs(2440) <= (inputs(219)) xor (inputs(208));
    layer0_outputs(2441) <= '0';
    layer0_outputs(2442) <= (inputs(219)) and (inputs(31));
    layer0_outputs(2443) <= '0';
    layer0_outputs(2444) <= not((inputs(86)) and (inputs(19)));
    layer0_outputs(2445) <= not(inputs(231));
    layer0_outputs(2446) <= '1';
    layer0_outputs(2447) <= (inputs(166)) and (inputs(109));
    layer0_outputs(2448) <= not((inputs(179)) or (inputs(239)));
    layer0_outputs(2449) <= (inputs(208)) and not (inputs(172));
    layer0_outputs(2450) <= (inputs(72)) or (inputs(232));
    layer0_outputs(2451) <= not(inputs(130));
    layer0_outputs(2452) <= (inputs(220)) or (inputs(187));
    layer0_outputs(2453) <= (inputs(127)) and not (inputs(251));
    layer0_outputs(2454) <= '0';
    layer0_outputs(2455) <= (inputs(16)) and (inputs(94));
    layer0_outputs(2456) <= not(inputs(51));
    layer0_outputs(2457) <= '1';
    layer0_outputs(2458) <= not(inputs(228));
    layer0_outputs(2459) <= inputs(14);
    layer0_outputs(2460) <= not((inputs(44)) or (inputs(154)));
    layer0_outputs(2461) <= inputs(121);
    layer0_outputs(2462) <= not(inputs(134));
    layer0_outputs(2463) <= '0';
    layer0_outputs(2464) <= not(inputs(124));
    layer0_outputs(2465) <= (inputs(67)) or (inputs(83));
    layer0_outputs(2466) <= inputs(39);
    layer0_outputs(2467) <= not(inputs(71));
    layer0_outputs(2468) <= (inputs(18)) or (inputs(5));
    layer0_outputs(2469) <= (inputs(162)) and not (inputs(95));
    layer0_outputs(2470) <= inputs(180);
    layer0_outputs(2471) <= (inputs(21)) xor (inputs(101));
    layer0_outputs(2472) <= inputs(35);
    layer0_outputs(2473) <= '1';
    layer0_outputs(2474) <= not(inputs(149)) or (inputs(136));
    layer0_outputs(2475) <= (inputs(195)) or (inputs(11));
    layer0_outputs(2476) <= not(inputs(6));
    layer0_outputs(2477) <= not(inputs(0));
    layer0_outputs(2478) <= '1';
    layer0_outputs(2479) <= not(inputs(20)) or (inputs(146));
    layer0_outputs(2480) <= (inputs(227)) and not (inputs(216));
    layer0_outputs(2481) <= not(inputs(188));
    layer0_outputs(2482) <= not(inputs(186));
    layer0_outputs(2483) <= inputs(106);
    layer0_outputs(2484) <= (inputs(107)) and (inputs(117));
    layer0_outputs(2485) <= not(inputs(61));
    layer0_outputs(2486) <= (inputs(254)) or (inputs(239));
    layer0_outputs(2487) <= not(inputs(79));
    layer0_outputs(2488) <= (inputs(163)) and not (inputs(3));
    layer0_outputs(2489) <= not(inputs(114));
    layer0_outputs(2490) <= not(inputs(41));
    layer0_outputs(2491) <= (inputs(144)) or (inputs(206));
    layer0_outputs(2492) <= (inputs(231)) and (inputs(109));
    layer0_outputs(2493) <= (inputs(241)) and not (inputs(33));
    layer0_outputs(2494) <= '1';
    layer0_outputs(2495) <= (inputs(178)) and not (inputs(15));
    layer0_outputs(2496) <= '1';
    layer0_outputs(2497) <= inputs(121);
    layer0_outputs(2498) <= '0';
    layer0_outputs(2499) <= not(inputs(168)) or (inputs(42));
    layer0_outputs(2500) <= inputs(195);
    layer0_outputs(2501) <= inputs(203);
    layer0_outputs(2502) <= (inputs(73)) and (inputs(173));
    layer0_outputs(2503) <= (inputs(179)) and not (inputs(223));
    layer0_outputs(2504) <= (inputs(139)) and (inputs(153));
    layer0_outputs(2505) <= not((inputs(234)) and (inputs(221)));
    layer0_outputs(2506) <= '1';
    layer0_outputs(2507) <= '1';
    layer0_outputs(2508) <= '1';
    layer0_outputs(2509) <= not(inputs(104));
    layer0_outputs(2510) <= (inputs(29)) and not (inputs(236));
    layer0_outputs(2511) <= (inputs(95)) and (inputs(35));
    layer0_outputs(2512) <= not(inputs(179));
    layer0_outputs(2513) <= not(inputs(204));
    layer0_outputs(2514) <= (inputs(85)) or (inputs(111));
    layer0_outputs(2515) <= inputs(72);
    layer0_outputs(2516) <= (inputs(232)) or (inputs(68));
    layer0_outputs(2517) <= '0';
    layer0_outputs(2518) <= not(inputs(21));
    layer0_outputs(2519) <= not(inputs(110));
    layer0_outputs(2520) <= inputs(227);
    layer0_outputs(2521) <= not((inputs(118)) and (inputs(32)));
    layer0_outputs(2522) <= not((inputs(231)) and (inputs(122)));
    layer0_outputs(2523) <= '0';
    layer0_outputs(2524) <= '0';
    layer0_outputs(2525) <= not((inputs(241)) and (inputs(253)));
    layer0_outputs(2526) <= (inputs(118)) and not (inputs(5));
    layer0_outputs(2527) <= not(inputs(15)) or (inputs(249));
    layer0_outputs(2528) <= not(inputs(75));
    layer0_outputs(2529) <= not((inputs(145)) or (inputs(130)));
    layer0_outputs(2530) <= not(inputs(4));
    layer0_outputs(2531) <= inputs(240);
    layer0_outputs(2532) <= '1';
    layer0_outputs(2533) <= (inputs(226)) and not (inputs(149));
    layer0_outputs(2534) <= '0';
    layer0_outputs(2535) <= (inputs(122)) or (inputs(168));
    layer0_outputs(2536) <= '1';
    layer0_outputs(2537) <= not(inputs(150)) or (inputs(228));
    layer0_outputs(2538) <= not(inputs(11)) or (inputs(24));
    layer0_outputs(2539) <= inputs(190);
    layer0_outputs(2540) <= (inputs(169)) or (inputs(102));
    layer0_outputs(2541) <= inputs(105);
    layer0_outputs(2542) <= inputs(152);
    layer0_outputs(2543) <= '1';
    layer0_outputs(2544) <= not(inputs(98));
    layer0_outputs(2545) <= '1';
    layer0_outputs(2546) <= (inputs(8)) or (inputs(77));
    layer0_outputs(2547) <= '1';
    layer0_outputs(2548) <= not(inputs(230)) or (inputs(167));
    layer0_outputs(2549) <= '1';
    layer0_outputs(2550) <= not(inputs(10)) or (inputs(226));
    layer0_outputs(2551) <= not((inputs(136)) and (inputs(27)));
    layer0_outputs(2552) <= not((inputs(115)) or (inputs(95)));
    layer0_outputs(2553) <= (inputs(114)) or (inputs(169));
    layer0_outputs(2554) <= inputs(196);
    layer0_outputs(2555) <= not(inputs(86)) or (inputs(187));
    layer0_outputs(2556) <= (inputs(152)) or (inputs(241));
    layer0_outputs(2557) <= not(inputs(137));
    layer0_outputs(2558) <= not((inputs(245)) or (inputs(104)));
    layer0_outputs(2559) <= not(inputs(162));
    layer1_outputs(0) <= '1';
    layer1_outputs(1) <= layer0_outputs(618);
    layer1_outputs(2) <= layer0_outputs(676);
    layer1_outputs(3) <= '1';
    layer1_outputs(4) <= not(layer0_outputs(444));
    layer1_outputs(5) <= (layer0_outputs(1763)) and (layer0_outputs(1052));
    layer1_outputs(6) <= '0';
    layer1_outputs(7) <= (layer0_outputs(1227)) and (layer0_outputs(257));
    layer1_outputs(8) <= not(layer0_outputs(1184));
    layer1_outputs(9) <= (layer0_outputs(1687)) and (layer0_outputs(1546));
    layer1_outputs(10) <= not((layer0_outputs(741)) or (layer0_outputs(2359)));
    layer1_outputs(11) <= '0';
    layer1_outputs(12) <= (layer0_outputs(140)) and (layer0_outputs(545));
    layer1_outputs(13) <= layer0_outputs(2231);
    layer1_outputs(14) <= not(layer0_outputs(107));
    layer1_outputs(15) <= (layer0_outputs(2339)) or (layer0_outputs(2408));
    layer1_outputs(16) <= layer0_outputs(1219);
    layer1_outputs(17) <= layer0_outputs(56);
    layer1_outputs(18) <= (layer0_outputs(1778)) and not (layer0_outputs(116));
    layer1_outputs(19) <= '1';
    layer1_outputs(20) <= layer0_outputs(1598);
    layer1_outputs(21) <= (layer0_outputs(2194)) and not (layer0_outputs(1827));
    layer1_outputs(22) <= '1';
    layer1_outputs(23) <= not(layer0_outputs(1367)) or (layer0_outputs(170));
    layer1_outputs(24) <= layer0_outputs(1557);
    layer1_outputs(25) <= not(layer0_outputs(1474));
    layer1_outputs(26) <= not(layer0_outputs(2263));
    layer1_outputs(27) <= not(layer0_outputs(1900)) or (layer0_outputs(2512));
    layer1_outputs(28) <= (layer0_outputs(1396)) and not (layer0_outputs(2213));
    layer1_outputs(29) <= layer0_outputs(419);
    layer1_outputs(30) <= '0';
    layer1_outputs(31) <= (layer0_outputs(415)) or (layer0_outputs(1066));
    layer1_outputs(32) <= layer0_outputs(1521);
    layer1_outputs(33) <= not((layer0_outputs(1475)) or (layer0_outputs(2373)));
    layer1_outputs(34) <= (layer0_outputs(1366)) or (layer0_outputs(583));
    layer1_outputs(35) <= '0';
    layer1_outputs(36) <= layer0_outputs(2154);
    layer1_outputs(37) <= '1';
    layer1_outputs(38) <= '0';
    layer1_outputs(39) <= (layer0_outputs(2168)) and not (layer0_outputs(505));
    layer1_outputs(40) <= '1';
    layer1_outputs(41) <= (layer0_outputs(1282)) and (layer0_outputs(746));
    layer1_outputs(42) <= '1';
    layer1_outputs(43) <= not((layer0_outputs(527)) or (layer0_outputs(2482)));
    layer1_outputs(44) <= '1';
    layer1_outputs(45) <= (layer0_outputs(2204)) and not (layer0_outputs(1661));
    layer1_outputs(46) <= '0';
    layer1_outputs(47) <= not(layer0_outputs(326));
    layer1_outputs(48) <= not(layer0_outputs(1198));
    layer1_outputs(49) <= not((layer0_outputs(134)) or (layer0_outputs(1067)));
    layer1_outputs(50) <= '1';
    layer1_outputs(51) <= (layer0_outputs(1162)) and (layer0_outputs(1966));
    layer1_outputs(52) <= '1';
    layer1_outputs(53) <= '0';
    layer1_outputs(54) <= '1';
    layer1_outputs(55) <= (layer0_outputs(2333)) and not (layer0_outputs(1283));
    layer1_outputs(56) <= layer0_outputs(77);
    layer1_outputs(57) <= not((layer0_outputs(2497)) or (layer0_outputs(1834)));
    layer1_outputs(58) <= (layer0_outputs(1238)) or (layer0_outputs(1637));
    layer1_outputs(59) <= not((layer0_outputs(2232)) or (layer0_outputs(438)));
    layer1_outputs(60) <= not((layer0_outputs(1121)) xor (layer0_outputs(557)));
    layer1_outputs(61) <= not(layer0_outputs(902));
    layer1_outputs(62) <= (layer0_outputs(13)) and not (layer0_outputs(1866));
    layer1_outputs(63) <= layer0_outputs(2108);
    layer1_outputs(64) <= '0';
    layer1_outputs(65) <= not(layer0_outputs(805)) or (layer0_outputs(524));
    layer1_outputs(66) <= (layer0_outputs(743)) or (layer0_outputs(1214));
    layer1_outputs(67) <= layer0_outputs(1736);
    layer1_outputs(68) <= (layer0_outputs(23)) and (layer0_outputs(1776));
    layer1_outputs(69) <= not(layer0_outputs(875)) or (layer0_outputs(1361));
    layer1_outputs(70) <= not(layer0_outputs(807));
    layer1_outputs(71) <= not((layer0_outputs(1925)) and (layer0_outputs(16)));
    layer1_outputs(72) <= not((layer0_outputs(2295)) and (layer0_outputs(1172)));
    layer1_outputs(73) <= not(layer0_outputs(1160));
    layer1_outputs(74) <= '1';
    layer1_outputs(75) <= not((layer0_outputs(1509)) and (layer0_outputs(2029)));
    layer1_outputs(76) <= layer0_outputs(1722);
    layer1_outputs(77) <= not(layer0_outputs(1432));
    layer1_outputs(78) <= not(layer0_outputs(788));
    layer1_outputs(79) <= '0';
    layer1_outputs(80) <= not((layer0_outputs(699)) or (layer0_outputs(673)));
    layer1_outputs(81) <= not(layer0_outputs(1824)) or (layer0_outputs(1582));
    layer1_outputs(82) <= layer0_outputs(1688);
    layer1_outputs(83) <= (layer0_outputs(1060)) and not (layer0_outputs(2162));
    layer1_outputs(84) <= '0';
    layer1_outputs(85) <= (layer0_outputs(1188)) and not (layer0_outputs(793));
    layer1_outputs(86) <= '0';
    layer1_outputs(87) <= not(layer0_outputs(2322)) or (layer0_outputs(1684));
    layer1_outputs(88) <= not(layer0_outputs(2162)) or (layer0_outputs(1635));
    layer1_outputs(89) <= (layer0_outputs(1005)) and (layer0_outputs(846));
    layer1_outputs(90) <= layer0_outputs(1281);
    layer1_outputs(91) <= (layer0_outputs(2067)) and not (layer0_outputs(1270));
    layer1_outputs(92) <= '1';
    layer1_outputs(93) <= not(layer0_outputs(1482)) or (layer0_outputs(752));
    layer1_outputs(94) <= not(layer0_outputs(1531));
    layer1_outputs(95) <= not(layer0_outputs(1572));
    layer1_outputs(96) <= '1';
    layer1_outputs(97) <= '1';
    layer1_outputs(98) <= (layer0_outputs(2423)) and not (layer0_outputs(43));
    layer1_outputs(99) <= (layer0_outputs(677)) and not (layer0_outputs(1759));
    layer1_outputs(100) <= '1';
    layer1_outputs(101) <= layer0_outputs(417);
    layer1_outputs(102) <= '0';
    layer1_outputs(103) <= (layer0_outputs(1013)) and (layer0_outputs(644));
    layer1_outputs(104) <= not(layer0_outputs(1300));
    layer1_outputs(105) <= not(layer0_outputs(932));
    layer1_outputs(106) <= layer0_outputs(1354);
    layer1_outputs(107) <= (layer0_outputs(2392)) and not (layer0_outputs(888));
    layer1_outputs(108) <= '0';
    layer1_outputs(109) <= not(layer0_outputs(927)) or (layer0_outputs(1337));
    layer1_outputs(110) <= '0';
    layer1_outputs(111) <= not(layer0_outputs(1647)) or (layer0_outputs(984));
    layer1_outputs(112) <= layer0_outputs(1481);
    layer1_outputs(113) <= layer0_outputs(1910);
    layer1_outputs(114) <= (layer0_outputs(1568)) and not (layer0_outputs(1185));
    layer1_outputs(115) <= (layer0_outputs(904)) or (layer0_outputs(1029));
    layer1_outputs(116) <= '1';
    layer1_outputs(117) <= '1';
    layer1_outputs(118) <= not(layer0_outputs(1522));
    layer1_outputs(119) <= layer0_outputs(2418);
    layer1_outputs(120) <= not(layer0_outputs(241));
    layer1_outputs(121) <= not((layer0_outputs(1684)) or (layer0_outputs(1987)));
    layer1_outputs(122) <= not(layer0_outputs(2323));
    layer1_outputs(123) <= layer0_outputs(517);
    layer1_outputs(124) <= not((layer0_outputs(2541)) or (layer0_outputs(469)));
    layer1_outputs(125) <= not((layer0_outputs(2109)) or (layer0_outputs(1124)));
    layer1_outputs(126) <= not(layer0_outputs(304));
    layer1_outputs(127) <= (layer0_outputs(2218)) and not (layer0_outputs(1925));
    layer1_outputs(128) <= (layer0_outputs(168)) and (layer0_outputs(2398));
    layer1_outputs(129) <= not(layer0_outputs(1117));
    layer1_outputs(130) <= not((layer0_outputs(28)) and (layer0_outputs(530)));
    layer1_outputs(131) <= layer0_outputs(70);
    layer1_outputs(132) <= not(layer0_outputs(2455)) or (layer0_outputs(1858));
    layer1_outputs(133) <= not(layer0_outputs(315)) or (layer0_outputs(1637));
    layer1_outputs(134) <= layer0_outputs(2319);
    layer1_outputs(135) <= not(layer0_outputs(207)) or (layer0_outputs(851));
    layer1_outputs(136) <= '1';
    layer1_outputs(137) <= not((layer0_outputs(225)) and (layer0_outputs(1364)));
    layer1_outputs(138) <= (layer0_outputs(833)) and not (layer0_outputs(2503));
    layer1_outputs(139) <= layer0_outputs(1564);
    layer1_outputs(140) <= not(layer0_outputs(1119)) or (layer0_outputs(1011));
    layer1_outputs(141) <= not(layer0_outputs(866)) or (layer0_outputs(711));
    layer1_outputs(142) <= not(layer0_outputs(274));
    layer1_outputs(143) <= '1';
    layer1_outputs(144) <= '0';
    layer1_outputs(145) <= '0';
    layer1_outputs(146) <= (layer0_outputs(2169)) and not (layer0_outputs(2299));
    layer1_outputs(147) <= not(layer0_outputs(436)) or (layer0_outputs(1302));
    layer1_outputs(148) <= not(layer0_outputs(563));
    layer1_outputs(149) <= not(layer0_outputs(613));
    layer1_outputs(150) <= (layer0_outputs(1693)) or (layer0_outputs(1783));
    layer1_outputs(151) <= not(layer0_outputs(204));
    layer1_outputs(152) <= '0';
    layer1_outputs(153) <= (layer0_outputs(689)) and not (layer0_outputs(743));
    layer1_outputs(154) <= '1';
    layer1_outputs(155) <= not((layer0_outputs(1180)) and (layer0_outputs(631)));
    layer1_outputs(156) <= not((layer0_outputs(1913)) xor (layer0_outputs(137)));
    layer1_outputs(157) <= layer0_outputs(1027);
    layer1_outputs(158) <= not((layer0_outputs(621)) or (layer0_outputs(930)));
    layer1_outputs(159) <= layer0_outputs(598);
    layer1_outputs(160) <= not(layer0_outputs(855)) or (layer0_outputs(2167));
    layer1_outputs(161) <= '1';
    layer1_outputs(162) <= (layer0_outputs(1359)) and (layer0_outputs(1043));
    layer1_outputs(163) <= not(layer0_outputs(445));
    layer1_outputs(164) <= not(layer0_outputs(117));
    layer1_outputs(165) <= '1';
    layer1_outputs(166) <= not((layer0_outputs(1626)) and (layer0_outputs(2243)));
    layer1_outputs(167) <= not((layer0_outputs(2378)) and (layer0_outputs(175)));
    layer1_outputs(168) <= '1';
    layer1_outputs(169) <= (layer0_outputs(2367)) and not (layer0_outputs(948));
    layer1_outputs(170) <= layer0_outputs(1488);
    layer1_outputs(171) <= '0';
    layer1_outputs(172) <= not(layer0_outputs(213));
    layer1_outputs(173) <= (layer0_outputs(1596)) and not (layer0_outputs(1562));
    layer1_outputs(174) <= (layer0_outputs(251)) and not (layer0_outputs(751));
    layer1_outputs(175) <= layer0_outputs(561);
    layer1_outputs(176) <= not(layer0_outputs(1284)) or (layer0_outputs(584));
    layer1_outputs(177) <= not(layer0_outputs(276));
    layer1_outputs(178) <= not(layer0_outputs(1310)) or (layer0_outputs(266));
    layer1_outputs(179) <= (layer0_outputs(1764)) and not (layer0_outputs(2210));
    layer1_outputs(180) <= (layer0_outputs(2231)) and not (layer0_outputs(2359));
    layer1_outputs(181) <= '1';
    layer1_outputs(182) <= not(layer0_outputs(1472));
    layer1_outputs(183) <= '1';
    layer1_outputs(184) <= (layer0_outputs(1423)) and not (layer0_outputs(1049));
    layer1_outputs(185) <= not(layer0_outputs(249)) or (layer0_outputs(1784));
    layer1_outputs(186) <= not(layer0_outputs(2233));
    layer1_outputs(187) <= not((layer0_outputs(1408)) or (layer0_outputs(1371)));
    layer1_outputs(188) <= (layer0_outputs(1660)) and not (layer0_outputs(1767));
    layer1_outputs(189) <= '1';
    layer1_outputs(190) <= layer0_outputs(885);
    layer1_outputs(191) <= not((layer0_outputs(495)) or (layer0_outputs(2133)));
    layer1_outputs(192) <= layer0_outputs(1843);
    layer1_outputs(193) <= not(layer0_outputs(238));
    layer1_outputs(194) <= (layer0_outputs(678)) and not (layer0_outputs(1075));
    layer1_outputs(195) <= not(layer0_outputs(1691));
    layer1_outputs(196) <= (layer0_outputs(674)) and (layer0_outputs(1617));
    layer1_outputs(197) <= (layer0_outputs(1985)) and not (layer0_outputs(943));
    layer1_outputs(198) <= (layer0_outputs(1663)) and (layer0_outputs(1530));
    layer1_outputs(199) <= not(layer0_outputs(1024));
    layer1_outputs(200) <= layer0_outputs(2138);
    layer1_outputs(201) <= (layer0_outputs(607)) or (layer0_outputs(288));
    layer1_outputs(202) <= not(layer0_outputs(1476));
    layer1_outputs(203) <= not((layer0_outputs(1501)) or (layer0_outputs(94)));
    layer1_outputs(204) <= (layer0_outputs(970)) xor (layer0_outputs(221));
    layer1_outputs(205) <= (layer0_outputs(903)) or (layer0_outputs(1474));
    layer1_outputs(206) <= layer0_outputs(548);
    layer1_outputs(207) <= (layer0_outputs(727)) or (layer0_outputs(39));
    layer1_outputs(208) <= layer0_outputs(2295);
    layer1_outputs(209) <= layer0_outputs(144);
    layer1_outputs(210) <= not(layer0_outputs(1611)) or (layer0_outputs(1797));
    layer1_outputs(211) <= not(layer0_outputs(1415)) or (layer0_outputs(2217));
    layer1_outputs(212) <= (layer0_outputs(2481)) and not (layer0_outputs(2388));
    layer1_outputs(213) <= (layer0_outputs(1251)) or (layer0_outputs(504));
    layer1_outputs(214) <= (layer0_outputs(1518)) and not (layer0_outputs(1733));
    layer1_outputs(215) <= not((layer0_outputs(138)) and (layer0_outputs(2000)));
    layer1_outputs(216) <= '0';
    layer1_outputs(217) <= layer0_outputs(92);
    layer1_outputs(218) <= not(layer0_outputs(1235));
    layer1_outputs(219) <= not(layer0_outputs(227)) or (layer0_outputs(500));
    layer1_outputs(220) <= '1';
    layer1_outputs(221) <= not(layer0_outputs(1239)) or (layer0_outputs(760));
    layer1_outputs(222) <= (layer0_outputs(1786)) and (layer0_outputs(1932));
    layer1_outputs(223) <= '0';
    layer1_outputs(224) <= '0';
    layer1_outputs(225) <= (layer0_outputs(744)) and not (layer0_outputs(1447));
    layer1_outputs(226) <= '0';
    layer1_outputs(227) <= (layer0_outputs(117)) or (layer0_outputs(72));
    layer1_outputs(228) <= not((layer0_outputs(811)) or (layer0_outputs(2088)));
    layer1_outputs(229) <= not(layer0_outputs(2063)) or (layer0_outputs(1224));
    layer1_outputs(230) <= '0';
    layer1_outputs(231) <= '0';
    layer1_outputs(232) <= (layer0_outputs(2317)) or (layer0_outputs(2252));
    layer1_outputs(233) <= not((layer0_outputs(525)) or (layer0_outputs(1507)));
    layer1_outputs(234) <= not(layer0_outputs(2375));
    layer1_outputs(235) <= not((layer0_outputs(864)) and (layer0_outputs(11)));
    layer1_outputs(236) <= (layer0_outputs(1518)) or (layer0_outputs(699));
    layer1_outputs(237) <= not(layer0_outputs(544)) or (layer0_outputs(292));
    layer1_outputs(238) <= layer0_outputs(619);
    layer1_outputs(239) <= (layer0_outputs(1565)) and not (layer0_outputs(1085));
    layer1_outputs(240) <= not(layer0_outputs(349));
    layer1_outputs(241) <= '1';
    layer1_outputs(242) <= not(layer0_outputs(1243));
    layer1_outputs(243) <= (layer0_outputs(1178)) and not (layer0_outputs(2441));
    layer1_outputs(244) <= not((layer0_outputs(876)) or (layer0_outputs(2258)));
    layer1_outputs(245) <= layer0_outputs(1172);
    layer1_outputs(246) <= not((layer0_outputs(498)) xor (layer0_outputs(1958)));
    layer1_outputs(247) <= not(layer0_outputs(251));
    layer1_outputs(248) <= (layer0_outputs(1424)) and not (layer0_outputs(1063));
    layer1_outputs(249) <= (layer0_outputs(753)) or (layer0_outputs(2002));
    layer1_outputs(250) <= '0';
    layer1_outputs(251) <= '0';
    layer1_outputs(252) <= '1';
    layer1_outputs(253) <= not(layer0_outputs(2172)) or (layer0_outputs(569));
    layer1_outputs(254) <= not(layer0_outputs(327));
    layer1_outputs(255) <= '0';
    layer1_outputs(256) <= not((layer0_outputs(1301)) and (layer0_outputs(399)));
    layer1_outputs(257) <= layer0_outputs(239);
    layer1_outputs(258) <= '0';
    layer1_outputs(259) <= (layer0_outputs(1422)) or (layer0_outputs(458));
    layer1_outputs(260) <= layer0_outputs(1651);
    layer1_outputs(261) <= (layer0_outputs(1386)) and not (layer0_outputs(1728));
    layer1_outputs(262) <= not(layer0_outputs(2039)) or (layer0_outputs(836));
    layer1_outputs(263) <= (layer0_outputs(1071)) and not (layer0_outputs(1487));
    layer1_outputs(264) <= (layer0_outputs(753)) and not (layer0_outputs(912));
    layer1_outputs(265) <= '0';
    layer1_outputs(266) <= not(layer0_outputs(240));
    layer1_outputs(267) <= layer0_outputs(2267);
    layer1_outputs(268) <= layer0_outputs(272);
    layer1_outputs(269) <= '0';
    layer1_outputs(270) <= layer0_outputs(990);
    layer1_outputs(271) <= (layer0_outputs(1966)) or (layer0_outputs(2223));
    layer1_outputs(272) <= layer0_outputs(2320);
    layer1_outputs(273) <= layer0_outputs(1597);
    layer1_outputs(274) <= not(layer0_outputs(962)) or (layer0_outputs(2166));
    layer1_outputs(275) <= not((layer0_outputs(1247)) or (layer0_outputs(2030)));
    layer1_outputs(276) <= not(layer0_outputs(124));
    layer1_outputs(277) <= '0';
    layer1_outputs(278) <= layer0_outputs(1147);
    layer1_outputs(279) <= '0';
    layer1_outputs(280) <= layer0_outputs(1895);
    layer1_outputs(281) <= layer0_outputs(2254);
    layer1_outputs(282) <= not(layer0_outputs(2384));
    layer1_outputs(283) <= (layer0_outputs(2302)) and not (layer0_outputs(1463));
    layer1_outputs(284) <= '0';
    layer1_outputs(285) <= not(layer0_outputs(1381)) or (layer0_outputs(1832));
    layer1_outputs(286) <= layer0_outputs(179);
    layer1_outputs(287) <= not(layer0_outputs(375)) or (layer0_outputs(49));
    layer1_outputs(288) <= not((layer0_outputs(2387)) and (layer0_outputs(1149)));
    layer1_outputs(289) <= '1';
    layer1_outputs(290) <= not((layer0_outputs(1911)) and (layer0_outputs(230)));
    layer1_outputs(291) <= layer0_outputs(2032);
    layer1_outputs(292) <= not(layer0_outputs(1624)) or (layer0_outputs(360));
    layer1_outputs(293) <= not(layer0_outputs(199));
    layer1_outputs(294) <= not(layer0_outputs(536));
    layer1_outputs(295) <= not((layer0_outputs(28)) xor (layer0_outputs(2477)));
    layer1_outputs(296) <= not((layer0_outputs(56)) or (layer0_outputs(2094)));
    layer1_outputs(297) <= (layer0_outputs(2188)) and not (layer0_outputs(2284));
    layer1_outputs(298) <= layer0_outputs(1195);
    layer1_outputs(299) <= layer0_outputs(244);
    layer1_outputs(300) <= (layer0_outputs(1169)) and (layer0_outputs(2443));
    layer1_outputs(301) <= layer0_outputs(1820);
    layer1_outputs(302) <= '1';
    layer1_outputs(303) <= '0';
    layer1_outputs(304) <= not(layer0_outputs(718));
    layer1_outputs(305) <= '0';
    layer1_outputs(306) <= not(layer0_outputs(1745)) or (layer0_outputs(66));
    layer1_outputs(307) <= not(layer0_outputs(1755));
    layer1_outputs(308) <= not((layer0_outputs(1185)) or (layer0_outputs(2463)));
    layer1_outputs(309) <= layer0_outputs(339);
    layer1_outputs(310) <= not(layer0_outputs(13));
    layer1_outputs(311) <= '1';
    layer1_outputs(312) <= not(layer0_outputs(1439));
    layer1_outputs(313) <= (layer0_outputs(2555)) and not (layer0_outputs(216));
    layer1_outputs(314) <= layer0_outputs(1062);
    layer1_outputs(315) <= not((layer0_outputs(1342)) or (layer0_outputs(488)));
    layer1_outputs(316) <= (layer0_outputs(882)) or (layer0_outputs(2551));
    layer1_outputs(317) <= layer0_outputs(184);
    layer1_outputs(318) <= not((layer0_outputs(1449)) or (layer0_outputs(1153)));
    layer1_outputs(319) <= not(layer0_outputs(2248)) or (layer0_outputs(671));
    layer1_outputs(320) <= '0';
    layer1_outputs(321) <= '1';
    layer1_outputs(322) <= layer0_outputs(2286);
    layer1_outputs(323) <= not(layer0_outputs(2024)) or (layer0_outputs(794));
    layer1_outputs(324) <= layer0_outputs(2130);
    layer1_outputs(325) <= not(layer0_outputs(1773));
    layer1_outputs(326) <= not(layer0_outputs(1404));
    layer1_outputs(327) <= layer0_outputs(1345);
    layer1_outputs(328) <= (layer0_outputs(657)) and not (layer0_outputs(731));
    layer1_outputs(329) <= not(layer0_outputs(708));
    layer1_outputs(330) <= '1';
    layer1_outputs(331) <= not((layer0_outputs(1886)) or (layer0_outputs(2226)));
    layer1_outputs(332) <= not(layer0_outputs(1760)) or (layer0_outputs(2530));
    layer1_outputs(333) <= layer0_outputs(999);
    layer1_outputs(334) <= (layer0_outputs(1974)) and not (layer0_outputs(1149));
    layer1_outputs(335) <= not(layer0_outputs(1311));
    layer1_outputs(336) <= not(layer0_outputs(1024)) or (layer0_outputs(1877));
    layer1_outputs(337) <= '1';
    layer1_outputs(338) <= not(layer0_outputs(435)) or (layer0_outputs(654));
    layer1_outputs(339) <= not((layer0_outputs(2372)) or (layer0_outputs(1751)));
    layer1_outputs(340) <= (layer0_outputs(2529)) and not (layer0_outputs(558));
    layer1_outputs(341) <= not(layer0_outputs(2243));
    layer1_outputs(342) <= '0';
    layer1_outputs(343) <= (layer0_outputs(1967)) and not (layer0_outputs(1395));
    layer1_outputs(344) <= layer0_outputs(286);
    layer1_outputs(345) <= '0';
    layer1_outputs(346) <= layer0_outputs(1629);
    layer1_outputs(347) <= not(layer0_outputs(2301));
    layer1_outputs(348) <= '0';
    layer1_outputs(349) <= (layer0_outputs(920)) xor (layer0_outputs(152));
    layer1_outputs(350) <= layer0_outputs(1028);
    layer1_outputs(351) <= not((layer0_outputs(2490)) and (layer0_outputs(2376)));
    layer1_outputs(352) <= not(layer0_outputs(2046));
    layer1_outputs(353) <= not((layer0_outputs(284)) or (layer0_outputs(2117)));
    layer1_outputs(354) <= not(layer0_outputs(709));
    layer1_outputs(355) <= not((layer0_outputs(1685)) or (layer0_outputs(2550)));
    layer1_outputs(356) <= layer0_outputs(140);
    layer1_outputs(357) <= not(layer0_outputs(10)) or (layer0_outputs(153));
    layer1_outputs(358) <= not((layer0_outputs(219)) xor (layer0_outputs(1116)));
    layer1_outputs(359) <= (layer0_outputs(2160)) and not (layer0_outputs(538));
    layer1_outputs(360) <= (layer0_outputs(817)) xor (layer0_outputs(577));
    layer1_outputs(361) <= not(layer0_outputs(664)) or (layer0_outputs(201));
    layer1_outputs(362) <= layer0_outputs(450);
    layer1_outputs(363) <= not((layer0_outputs(106)) and (layer0_outputs(1854)));
    layer1_outputs(364) <= (layer0_outputs(1000)) and not (layer0_outputs(217));
    layer1_outputs(365) <= '0';
    layer1_outputs(366) <= not(layer0_outputs(2381)) or (layer0_outputs(1313));
    layer1_outputs(367) <= not(layer0_outputs(1480)) or (layer0_outputs(1257));
    layer1_outputs(368) <= '0';
    layer1_outputs(369) <= '0';
    layer1_outputs(370) <= layer0_outputs(1304);
    layer1_outputs(371) <= (layer0_outputs(923)) or (layer0_outputs(1208));
    layer1_outputs(372) <= not(layer0_outputs(1100)) or (layer0_outputs(792));
    layer1_outputs(373) <= '1';
    layer1_outputs(374) <= not((layer0_outputs(1030)) or (layer0_outputs(53)));
    layer1_outputs(375) <= not(layer0_outputs(868));
    layer1_outputs(376) <= '0';
    layer1_outputs(377) <= layer0_outputs(1369);
    layer1_outputs(378) <= layer0_outputs(1585);
    layer1_outputs(379) <= layer0_outputs(796);
    layer1_outputs(380) <= (layer0_outputs(30)) or (layer0_outputs(580));
    layer1_outputs(381) <= layer0_outputs(2510);
    layer1_outputs(382) <= layer0_outputs(690);
    layer1_outputs(383) <= '0';
    layer1_outputs(384) <= not(layer0_outputs(350)) or (layer0_outputs(1835));
    layer1_outputs(385) <= '1';
    layer1_outputs(386) <= not(layer0_outputs(269));
    layer1_outputs(387) <= not(layer0_outputs(229)) or (layer0_outputs(2399));
    layer1_outputs(388) <= '1';
    layer1_outputs(389) <= not(layer0_outputs(2414));
    layer1_outputs(390) <= '1';
    layer1_outputs(391) <= layer0_outputs(1790);
    layer1_outputs(392) <= '0';
    layer1_outputs(393) <= not(layer0_outputs(2037)) or (layer0_outputs(2456));
    layer1_outputs(394) <= not(layer0_outputs(2116));
    layer1_outputs(395) <= (layer0_outputs(2010)) and not (layer0_outputs(1014));
    layer1_outputs(396) <= not((layer0_outputs(642)) and (layer0_outputs(2083)));
    layer1_outputs(397) <= not(layer0_outputs(1333));
    layer1_outputs(398) <= not(layer0_outputs(1090));
    layer1_outputs(399) <= not(layer0_outputs(667));
    layer1_outputs(400) <= not((layer0_outputs(465)) or (layer0_outputs(694)));
    layer1_outputs(401) <= not((layer0_outputs(1431)) and (layer0_outputs(1810)));
    layer1_outputs(402) <= not((layer0_outputs(1867)) or (layer0_outputs(2245)));
    layer1_outputs(403) <= not(layer0_outputs(1443));
    layer1_outputs(404) <= '0';
    layer1_outputs(405) <= (layer0_outputs(2220)) and not (layer0_outputs(306));
    layer1_outputs(406) <= (layer0_outputs(2487)) and not (layer0_outputs(1577));
    layer1_outputs(407) <= not(layer0_outputs(1010)) or (layer0_outputs(1585));
    layer1_outputs(408) <= not((layer0_outputs(1406)) or (layer0_outputs(1456)));
    layer1_outputs(409) <= layer0_outputs(645);
    layer1_outputs(410) <= layer0_outputs(2440);
    layer1_outputs(411) <= (layer0_outputs(2097)) and not (layer0_outputs(1471));
    layer1_outputs(412) <= '0';
    layer1_outputs(413) <= (layer0_outputs(2219)) and not (layer0_outputs(870));
    layer1_outputs(414) <= layer0_outputs(611);
    layer1_outputs(415) <= '1';
    layer1_outputs(416) <= not((layer0_outputs(2127)) or (layer0_outputs(630)));
    layer1_outputs(417) <= not((layer0_outputs(860)) and (layer0_outputs(1418)));
    layer1_outputs(418) <= not(layer0_outputs(1131));
    layer1_outputs(419) <= '0';
    layer1_outputs(420) <= layer0_outputs(1076);
    layer1_outputs(421) <= '1';
    layer1_outputs(422) <= not((layer0_outputs(867)) and (layer0_outputs(2026)));
    layer1_outputs(423) <= layer0_outputs(816);
    layer1_outputs(424) <= not((layer0_outputs(245)) and (layer0_outputs(723)));
    layer1_outputs(425) <= (layer0_outputs(1228)) and not (layer0_outputs(2317));
    layer1_outputs(426) <= (layer0_outputs(2090)) xor (layer0_outputs(586));
    layer1_outputs(427) <= not(layer0_outputs(438));
    layer1_outputs(428) <= not(layer0_outputs(1870));
    layer1_outputs(429) <= not((layer0_outputs(2486)) or (layer0_outputs(2190)));
    layer1_outputs(430) <= not(layer0_outputs(1365));
    layer1_outputs(431) <= '1';
    layer1_outputs(432) <= '0';
    layer1_outputs(433) <= not(layer0_outputs(1539));
    layer1_outputs(434) <= not(layer0_outputs(782));
    layer1_outputs(435) <= '1';
    layer1_outputs(436) <= not((layer0_outputs(2415)) and (layer0_outputs(1170)));
    layer1_outputs(437) <= not((layer0_outputs(1740)) or (layer0_outputs(354)));
    layer1_outputs(438) <= '0';
    layer1_outputs(439) <= '1';
    layer1_outputs(440) <= layer0_outputs(1452);
    layer1_outputs(441) <= not(layer0_outputs(481)) or (layer0_outputs(1528));
    layer1_outputs(442) <= not(layer0_outputs(1956));
    layer1_outputs(443) <= (layer0_outputs(184)) or (layer0_outputs(1542));
    layer1_outputs(444) <= not(layer0_outputs(1516)) or (layer0_outputs(1805));
    layer1_outputs(445) <= not(layer0_outputs(1904));
    layer1_outputs(446) <= not(layer0_outputs(1653));
    layer1_outputs(447) <= not((layer0_outputs(136)) or (layer0_outputs(220)));
    layer1_outputs(448) <= (layer0_outputs(62)) xor (layer0_outputs(176));
    layer1_outputs(449) <= not((layer0_outputs(1048)) or (layer0_outputs(1171)));
    layer1_outputs(450) <= not((layer0_outputs(951)) and (layer0_outputs(1686)));
    layer1_outputs(451) <= (layer0_outputs(718)) and (layer0_outputs(1287));
    layer1_outputs(452) <= not(layer0_outputs(317)) or (layer0_outputs(1152));
    layer1_outputs(453) <= not(layer0_outputs(504));
    layer1_outputs(454) <= not(layer0_outputs(1002)) or (layer0_outputs(1517));
    layer1_outputs(455) <= not(layer0_outputs(534));
    layer1_outputs(456) <= (layer0_outputs(1086)) and not (layer0_outputs(52));
    layer1_outputs(457) <= layer0_outputs(212);
    layer1_outputs(458) <= (layer0_outputs(1316)) and (layer0_outputs(725));
    layer1_outputs(459) <= not(layer0_outputs(1420)) or (layer0_outputs(536));
    layer1_outputs(460) <= not(layer0_outputs(2434));
    layer1_outputs(461) <= '1';
    layer1_outputs(462) <= layer0_outputs(599);
    layer1_outputs(463) <= (layer0_outputs(994)) or (layer0_outputs(424));
    layer1_outputs(464) <= '0';
    layer1_outputs(465) <= layer0_outputs(2410);
    layer1_outputs(466) <= (layer0_outputs(2478)) and not (layer0_outputs(1110));
    layer1_outputs(467) <= (layer0_outputs(621)) and not (layer0_outputs(126));
    layer1_outputs(468) <= not(layer0_outputs(1299));
    layer1_outputs(469) <= layer0_outputs(856);
    layer1_outputs(470) <= '0';
    layer1_outputs(471) <= not(layer0_outputs(2117)) or (layer0_outputs(2508));
    layer1_outputs(472) <= not(layer0_outputs(2381));
    layer1_outputs(473) <= not(layer0_outputs(1903)) or (layer0_outputs(409));
    layer1_outputs(474) <= not((layer0_outputs(834)) or (layer0_outputs(381)));
    layer1_outputs(475) <= '0';
    layer1_outputs(476) <= (layer0_outputs(1074)) and (layer0_outputs(1111));
    layer1_outputs(477) <= layer0_outputs(2419);
    layer1_outputs(478) <= not(layer0_outputs(1839));
    layer1_outputs(479) <= layer0_outputs(1210);
    layer1_outputs(480) <= not(layer0_outputs(73));
    layer1_outputs(481) <= layer0_outputs(2084);
    layer1_outputs(482) <= not(layer0_outputs(1886));
    layer1_outputs(483) <= layer0_outputs(854);
    layer1_outputs(484) <= (layer0_outputs(1673)) and (layer0_outputs(1695));
    layer1_outputs(485) <= layer0_outputs(2489);
    layer1_outputs(486) <= not((layer0_outputs(520)) and (layer0_outputs(1164)));
    layer1_outputs(487) <= (layer0_outputs(374)) or (layer0_outputs(2491));
    layer1_outputs(488) <= (layer0_outputs(70)) and not (layer0_outputs(494));
    layer1_outputs(489) <= (layer0_outputs(921)) and not (layer0_outputs(1756));
    layer1_outputs(490) <= not((layer0_outputs(123)) or (layer0_outputs(2388)));
    layer1_outputs(491) <= (layer0_outputs(1811)) or (layer0_outputs(1618));
    layer1_outputs(492) <= not(layer0_outputs(672));
    layer1_outputs(493) <= (layer0_outputs(130)) and not (layer0_outputs(1927));
    layer1_outputs(494) <= (layer0_outputs(1425)) or (layer0_outputs(506));
    layer1_outputs(495) <= not(layer0_outputs(1828));
    layer1_outputs(496) <= (layer0_outputs(2079)) and (layer0_outputs(2477));
    layer1_outputs(497) <= (layer0_outputs(2001)) and (layer0_outputs(1868));
    layer1_outputs(498) <= not((layer0_outputs(874)) and (layer0_outputs(617)));
    layer1_outputs(499) <= (layer0_outputs(1789)) or (layer0_outputs(1543));
    layer1_outputs(500) <= layer0_outputs(1515);
    layer1_outputs(501) <= (layer0_outputs(1129)) and not (layer0_outputs(1593));
    layer1_outputs(502) <= (layer0_outputs(1255)) and not (layer0_outputs(1998));
    layer1_outputs(503) <= not(layer0_outputs(1517)) or (layer0_outputs(2499));
    layer1_outputs(504) <= '1';
    layer1_outputs(505) <= (layer0_outputs(879)) or (layer0_outputs(304));
    layer1_outputs(506) <= (layer0_outputs(1231)) and not (layer0_outputs(2148));
    layer1_outputs(507) <= '0';
    layer1_outputs(508) <= not(layer0_outputs(560));
    layer1_outputs(509) <= '0';
    layer1_outputs(510) <= '1';
    layer1_outputs(511) <= not((layer0_outputs(707)) or (layer0_outputs(1222)));
    layer1_outputs(512) <= not((layer0_outputs(1917)) or (layer0_outputs(662)));
    layer1_outputs(513) <= layer0_outputs(848);
    layer1_outputs(514) <= not((layer0_outputs(2448)) or (layer0_outputs(1817)));
    layer1_outputs(515) <= '1';
    layer1_outputs(516) <= (layer0_outputs(716)) or (layer0_outputs(1514));
    layer1_outputs(517) <= (layer0_outputs(839)) and (layer0_outputs(490));
    layer1_outputs(518) <= not((layer0_outputs(954)) and (layer0_outputs(2112)));
    layer1_outputs(519) <= not(layer0_outputs(950)) or (layer0_outputs(746));
    layer1_outputs(520) <= layer0_outputs(859);
    layer1_outputs(521) <= not(layer0_outputs(645)) or (layer0_outputs(2483));
    layer1_outputs(522) <= '0';
    layer1_outputs(523) <= not(layer0_outputs(1026));
    layer1_outputs(524) <= (layer0_outputs(1079)) and not (layer0_outputs(773));
    layer1_outputs(525) <= layer0_outputs(1141);
    layer1_outputs(526) <= not(layer0_outputs(1971));
    layer1_outputs(527) <= layer0_outputs(1621);
    layer1_outputs(528) <= '0';
    layer1_outputs(529) <= '0';
    layer1_outputs(530) <= not(layer0_outputs(1370));
    layer1_outputs(531) <= layer0_outputs(1889);
    layer1_outputs(532) <= '0';
    layer1_outputs(533) <= not(layer0_outputs(1896));
    layer1_outputs(534) <= layer0_outputs(2552);
    layer1_outputs(535) <= '0';
    layer1_outputs(536) <= not(layer0_outputs(1078)) or (layer0_outputs(578));
    layer1_outputs(537) <= '0';
    layer1_outputs(538) <= (layer0_outputs(1144)) and (layer0_outputs(1298));
    layer1_outputs(539) <= '1';
    layer1_outputs(540) <= not((layer0_outputs(1489)) or (layer0_outputs(404)));
    layer1_outputs(541) <= (layer0_outputs(1299)) or (layer0_outputs(1421));
    layer1_outputs(542) <= '0';
    layer1_outputs(543) <= not(layer0_outputs(1631));
    layer1_outputs(544) <= not(layer0_outputs(566));
    layer1_outputs(545) <= '0';
    layer1_outputs(546) <= not(layer0_outputs(1940)) or (layer0_outputs(87));
    layer1_outputs(547) <= '0';
    layer1_outputs(548) <= layer0_outputs(604);
    layer1_outputs(549) <= (layer0_outputs(2332)) or (layer0_outputs(909));
    layer1_outputs(550) <= not(layer0_outputs(1607));
    layer1_outputs(551) <= (layer0_outputs(1544)) or (layer0_outputs(2227));
    layer1_outputs(552) <= layer0_outputs(1864);
    layer1_outputs(553) <= not(layer0_outputs(970));
    layer1_outputs(554) <= not(layer0_outputs(586)) or (layer0_outputs(1053));
    layer1_outputs(555) <= (layer0_outputs(599)) or (layer0_outputs(1163));
    layer1_outputs(556) <= not((layer0_outputs(2312)) and (layer0_outputs(1175)));
    layer1_outputs(557) <= '1';
    layer1_outputs(558) <= (layer0_outputs(2131)) and not (layer0_outputs(90));
    layer1_outputs(559) <= not((layer0_outputs(1862)) or (layer0_outputs(1743)));
    layer1_outputs(560) <= (layer0_outputs(837)) and (layer0_outputs(787));
    layer1_outputs(561) <= layer0_outputs(844);
    layer1_outputs(562) <= not(layer0_outputs(713));
    layer1_outputs(563) <= not((layer0_outputs(1852)) or (layer0_outputs(18)));
    layer1_outputs(564) <= layer0_outputs(895);
    layer1_outputs(565) <= layer0_outputs(722);
    layer1_outputs(566) <= not(layer0_outputs(1789));
    layer1_outputs(567) <= (layer0_outputs(2182)) and not (layer0_outputs(372));
    layer1_outputs(568) <= (layer0_outputs(1325)) and not (layer0_outputs(1389));
    layer1_outputs(569) <= not(layer0_outputs(2095));
    layer1_outputs(570) <= not(layer0_outputs(2180)) or (layer0_outputs(1899));
    layer1_outputs(571) <= (layer0_outputs(2009)) or (layer0_outputs(1934));
    layer1_outputs(572) <= not(layer0_outputs(511)) or (layer0_outputs(432));
    layer1_outputs(573) <= layer0_outputs(2070);
    layer1_outputs(574) <= (layer0_outputs(2060)) and (layer0_outputs(1008));
    layer1_outputs(575) <= not((layer0_outputs(2442)) and (layer0_outputs(1308)));
    layer1_outputs(576) <= '1';
    layer1_outputs(577) <= not(layer0_outputs(1514));
    layer1_outputs(578) <= not(layer0_outputs(388));
    layer1_outputs(579) <= (layer0_outputs(157)) and not (layer0_outputs(2047));
    layer1_outputs(580) <= not(layer0_outputs(2136));
    layer1_outputs(581) <= '1';
    layer1_outputs(582) <= '1';
    layer1_outputs(583) <= '0';
    layer1_outputs(584) <= not(layer0_outputs(738)) or (layer0_outputs(2229));
    layer1_outputs(585) <= '0';
    layer1_outputs(586) <= (layer0_outputs(1179)) and (layer0_outputs(726));
    layer1_outputs(587) <= layer0_outputs(2392);
    layer1_outputs(588) <= layer0_outputs(2224);
    layer1_outputs(589) <= not((layer0_outputs(508)) and (layer0_outputs(1642)));
    layer1_outputs(590) <= '0';
    layer1_outputs(591) <= layer0_outputs(1054);
    layer1_outputs(592) <= layer0_outputs(680);
    layer1_outputs(593) <= not(layer0_outputs(186));
    layer1_outputs(594) <= not((layer0_outputs(1742)) and (layer0_outputs(2488)));
    layer1_outputs(595) <= (layer0_outputs(2431)) and (layer0_outputs(1552));
    layer1_outputs(596) <= layer0_outputs(1051);
    layer1_outputs(597) <= '0';
    layer1_outputs(598) <= (layer0_outputs(1781)) and not (layer0_outputs(728));
    layer1_outputs(599) <= not((layer0_outputs(1402)) and (layer0_outputs(2313)));
    layer1_outputs(600) <= not(layer0_outputs(2124)) or (layer0_outputs(789));
    layer1_outputs(601) <= layer0_outputs(381);
    layer1_outputs(602) <= layer0_outputs(1458);
    layer1_outputs(603) <= '1';
    layer1_outputs(604) <= (layer0_outputs(728)) and not (layer0_outputs(1831));
    layer1_outputs(605) <= '0';
    layer1_outputs(606) <= not(layer0_outputs(47));
    layer1_outputs(607) <= '1';
    layer1_outputs(608) <= not(layer0_outputs(311)) or (layer0_outputs(2212));
    layer1_outputs(609) <= not((layer0_outputs(1403)) and (layer0_outputs(2250)));
    layer1_outputs(610) <= (layer0_outputs(559)) or (layer0_outputs(1560));
    layer1_outputs(611) <= (layer0_outputs(1566)) and not (layer0_outputs(826));
    layer1_outputs(612) <= layer0_outputs(1278);
    layer1_outputs(613) <= '0';
    layer1_outputs(614) <= '1';
    layer1_outputs(615) <= (layer0_outputs(1392)) or (layer0_outputs(1561));
    layer1_outputs(616) <= not(layer0_outputs(696));
    layer1_outputs(617) <= not((layer0_outputs(1503)) or (layer0_outputs(982)));
    layer1_outputs(618) <= not((layer0_outputs(1587)) or (layer0_outputs(2501)));
    layer1_outputs(619) <= '1';
    layer1_outputs(620) <= not(layer0_outputs(440));
    layer1_outputs(621) <= not(layer0_outputs(75));
    layer1_outputs(622) <= '1';
    layer1_outputs(623) <= not(layer0_outputs(190)) or (layer0_outputs(2384));
    layer1_outputs(624) <= (layer0_outputs(185)) or (layer0_outputs(977));
    layer1_outputs(625) <= not(layer0_outputs(1719)) or (layer0_outputs(210));
    layer1_outputs(626) <= not((layer0_outputs(2394)) and (layer0_outputs(433)));
    layer1_outputs(627) <= not((layer0_outputs(1259)) and (layer0_outputs(1186)));
    layer1_outputs(628) <= (layer0_outputs(1428)) and not (layer0_outputs(2170));
    layer1_outputs(629) <= not(layer0_outputs(1468));
    layer1_outputs(630) <= (layer0_outputs(1608)) or (layer0_outputs(2040));
    layer1_outputs(631) <= not(layer0_outputs(2185));
    layer1_outputs(632) <= '0';
    layer1_outputs(633) <= (layer0_outputs(507)) and not (layer0_outputs(1909));
    layer1_outputs(634) <= '0';
    layer1_outputs(635) <= layer0_outputs(890);
    layer1_outputs(636) <= '1';
    layer1_outputs(637) <= not(layer0_outputs(1435));
    layer1_outputs(638) <= (layer0_outputs(1706)) and not (layer0_outputs(1050));
    layer1_outputs(639) <= not(layer0_outputs(160));
    layer1_outputs(640) <= not((layer0_outputs(894)) and (layer0_outputs(1225)));
    layer1_outputs(641) <= not(layer0_outputs(978));
    layer1_outputs(642) <= not((layer0_outputs(1205)) and (layer0_outputs(71)));
    layer1_outputs(643) <= layer0_outputs(1583);
    layer1_outputs(644) <= layer0_outputs(956);
    layer1_outputs(645) <= layer0_outputs(2439);
    layer1_outputs(646) <= not(layer0_outputs(1856)) or (layer0_outputs(1248));
    layer1_outputs(647) <= '1';
    layer1_outputs(648) <= '1';
    layer1_outputs(649) <= not((layer0_outputs(2301)) and (layer0_outputs(1177)));
    layer1_outputs(650) <= (layer0_outputs(2290)) and (layer0_outputs(112));
    layer1_outputs(651) <= not((layer0_outputs(340)) or (layer0_outputs(411)));
    layer1_outputs(652) <= not(layer0_outputs(824));
    layer1_outputs(653) <= not(layer0_outputs(2147));
    layer1_outputs(654) <= '0';
    layer1_outputs(655) <= not(layer0_outputs(1654));
    layer1_outputs(656) <= not(layer0_outputs(1413));
    layer1_outputs(657) <= not(layer0_outputs(1241)) or (layer0_outputs(668));
    layer1_outputs(658) <= not(layer0_outputs(1387));
    layer1_outputs(659) <= (layer0_outputs(2389)) and (layer0_outputs(1001));
    layer1_outputs(660) <= (layer0_outputs(1576)) and (layer0_outputs(631));
    layer1_outputs(661) <= '0';
    layer1_outputs(662) <= layer0_outputs(2257);
    layer1_outputs(663) <= (layer0_outputs(1879)) and (layer0_outputs(1615));
    layer1_outputs(664) <= '1';
    layer1_outputs(665) <= not(layer0_outputs(1263));
    layer1_outputs(666) <= layer0_outputs(86);
    layer1_outputs(667) <= not(layer0_outputs(220));
    layer1_outputs(668) <= (layer0_outputs(1887)) and (layer0_outputs(2305));
    layer1_outputs(669) <= not(layer0_outputs(2497)) or (layer0_outputs(1443));
    layer1_outputs(670) <= not((layer0_outputs(2187)) or (layer0_outputs(1605)));
    layer1_outputs(671) <= not(layer0_outputs(1433)) or (layer0_outputs(1240));
    layer1_outputs(672) <= '0';
    layer1_outputs(673) <= '1';
    layer1_outputs(674) <= not((layer0_outputs(1295)) and (layer0_outputs(2150)));
    layer1_outputs(675) <= '0';
    layer1_outputs(676) <= '0';
    layer1_outputs(677) <= not(layer0_outputs(1211));
    layer1_outputs(678) <= not(layer0_outputs(228));
    layer1_outputs(679) <= not((layer0_outputs(1399)) and (layer0_outputs(748)));
    layer1_outputs(680) <= not((layer0_outputs(1451)) and (layer0_outputs(760)));
    layer1_outputs(681) <= not((layer0_outputs(1788)) and (layer0_outputs(729)));
    layer1_outputs(682) <= '1';
    layer1_outputs(683) <= not(layer0_outputs(609));
    layer1_outputs(684) <= layer0_outputs(1952);
    layer1_outputs(685) <= not((layer0_outputs(444)) and (layer0_outputs(814)));
    layer1_outputs(686) <= (layer0_outputs(1019)) and (layer0_outputs(2313));
    layer1_outputs(687) <= '0';
    layer1_outputs(688) <= (layer0_outputs(1271)) and not (layer0_outputs(897));
    layer1_outputs(689) <= layer0_outputs(1830);
    layer1_outputs(690) <= (layer0_outputs(1720)) and not (layer0_outputs(710));
    layer1_outputs(691) <= not(layer0_outputs(106)) or (layer0_outputs(879));
    layer1_outputs(692) <= '1';
    layer1_outputs(693) <= '1';
    layer1_outputs(694) <= layer0_outputs(1276);
    layer1_outputs(695) <= not((layer0_outputs(1878)) and (layer0_outputs(820)));
    layer1_outputs(696) <= '1';
    layer1_outputs(697) <= (layer0_outputs(332)) and not (layer0_outputs(2447));
    layer1_outputs(698) <= not((layer0_outputs(530)) or (layer0_outputs(2437)));
    layer1_outputs(699) <= not(layer0_outputs(1885)) or (layer0_outputs(2075));
    layer1_outputs(700) <= (layer0_outputs(235)) or (layer0_outputs(2170));
    layer1_outputs(701) <= not(layer0_outputs(2556));
    layer1_outputs(702) <= '1';
    layer1_outputs(703) <= (layer0_outputs(1110)) and (layer0_outputs(801));
    layer1_outputs(704) <= not(layer0_outputs(2376));
    layer1_outputs(705) <= (layer0_outputs(495)) and (layer0_outputs(1265));
    layer1_outputs(706) <= not((layer0_outputs(2307)) or (layer0_outputs(1350)));
    layer1_outputs(707) <= not((layer0_outputs(1534)) or (layer0_outputs(805)));
    layer1_outputs(708) <= not(layer0_outputs(2085)) or (layer0_outputs(2289));
    layer1_outputs(709) <= '0';
    layer1_outputs(710) <= '1';
    layer1_outputs(711) <= (layer0_outputs(947)) or (layer0_outputs(1022));
    layer1_outputs(712) <= (layer0_outputs(1306)) and (layer0_outputs(948));
    layer1_outputs(713) <= not(layer0_outputs(47)) or (layer0_outputs(2004));
    layer1_outputs(714) <= not(layer0_outputs(2152)) or (layer0_outputs(240));
    layer1_outputs(715) <= '1';
    layer1_outputs(716) <= not(layer0_outputs(154)) or (layer0_outputs(2040));
    layer1_outputs(717) <= (layer0_outputs(376)) or (layer0_outputs(2397));
    layer1_outputs(718) <= not(layer0_outputs(2360));
    layer1_outputs(719) <= not(layer0_outputs(243));
    layer1_outputs(720) <= layer0_outputs(303);
    layer1_outputs(721) <= '1';
    layer1_outputs(722) <= layer0_outputs(2520);
    layer1_outputs(723) <= layer0_outputs(1771);
    layer1_outputs(724) <= (layer0_outputs(963)) and not (layer0_outputs(1264));
    layer1_outputs(725) <= not((layer0_outputs(1266)) and (layer0_outputs(626)));
    layer1_outputs(726) <= not(layer0_outputs(509));
    layer1_outputs(727) <= (layer0_outputs(1866)) and not (layer0_outputs(301));
    layer1_outputs(728) <= '0';
    layer1_outputs(729) <= layer0_outputs(1527);
    layer1_outputs(730) <= (layer0_outputs(784)) and (layer0_outputs(967));
    layer1_outputs(731) <= not((layer0_outputs(2142)) and (layer0_outputs(2120)));
    layer1_outputs(732) <= (layer0_outputs(2402)) and not (layer0_outputs(1490));
    layer1_outputs(733) <= not(layer0_outputs(1143)) or (layer0_outputs(548));
    layer1_outputs(734) <= (layer0_outputs(2406)) and not (layer0_outputs(831));
    layer1_outputs(735) <= not(layer0_outputs(677));
    layer1_outputs(736) <= not(layer0_outputs(1202)) or (layer0_outputs(2486));
    layer1_outputs(737) <= '0';
    layer1_outputs(738) <= not(layer0_outputs(1896)) or (layer0_outputs(1434));
    layer1_outputs(739) <= layer0_outputs(338);
    layer1_outputs(740) <= not(layer0_outputs(452)) or (layer0_outputs(2371));
    layer1_outputs(741) <= '1';
    layer1_outputs(742) <= layer0_outputs(91);
    layer1_outputs(743) <= layer0_outputs(1788);
    layer1_outputs(744) <= (layer0_outputs(2016)) and not (layer0_outputs(1691));
    layer1_outputs(745) <= (layer0_outputs(2044)) and not (layer0_outputs(2322));
    layer1_outputs(746) <= not((layer0_outputs(2399)) and (layer0_outputs(2262)));
    layer1_outputs(747) <= not((layer0_outputs(1357)) and (layer0_outputs(2197)));
    layer1_outputs(748) <= not(layer0_outputs(1061));
    layer1_outputs(749) <= layer0_outputs(1096);
    layer1_outputs(750) <= '1';
    layer1_outputs(751) <= not(layer0_outputs(463));
    layer1_outputs(752) <= '0';
    layer1_outputs(753) <= not(layer0_outputs(143)) or (layer0_outputs(2160));
    layer1_outputs(754) <= not(layer0_outputs(196)) or (layer0_outputs(2008));
    layer1_outputs(755) <= not(layer0_outputs(2186));
    layer1_outputs(756) <= '1';
    layer1_outputs(757) <= (layer0_outputs(116)) or (layer0_outputs(2058));
    layer1_outputs(758) <= not(layer0_outputs(2140)) or (layer0_outputs(1366));
    layer1_outputs(759) <= (layer0_outputs(171)) or (layer0_outputs(212));
    layer1_outputs(760) <= (layer0_outputs(757)) or (layer0_outputs(502));
    layer1_outputs(761) <= (layer0_outputs(388)) or (layer0_outputs(1991));
    layer1_outputs(762) <= (layer0_outputs(512)) and (layer0_outputs(2209));
    layer1_outputs(763) <= (layer0_outputs(647)) or (layer0_outputs(1109));
    layer1_outputs(764) <= (layer0_outputs(2470)) and not (layer0_outputs(121));
    layer1_outputs(765) <= not((layer0_outputs(2063)) and (layer0_outputs(2279)));
    layer1_outputs(766) <= '0';
    layer1_outputs(767) <= layer0_outputs(2111);
    layer1_outputs(768) <= not(layer0_outputs(229)) or (layer0_outputs(1095));
    layer1_outputs(769) <= not(layer0_outputs(835));
    layer1_outputs(770) <= (layer0_outputs(2202)) and not (layer0_outputs(2316));
    layer1_outputs(771) <= (layer0_outputs(2315)) and not (layer0_outputs(336));
    layer1_outputs(772) <= not(layer0_outputs(1083)) or (layer0_outputs(2109));
    layer1_outputs(773) <= not(layer0_outputs(1769));
    layer1_outputs(774) <= not(layer0_outputs(277));
    layer1_outputs(775) <= not((layer0_outputs(441)) and (layer0_outputs(590)));
    layer1_outputs(776) <= layer0_outputs(1658);
    layer1_outputs(777) <= (layer0_outputs(2086)) and not (layer0_outputs(2223));
    layer1_outputs(778) <= not(layer0_outputs(1830)) or (layer0_outputs(691));
    layer1_outputs(779) <= not(layer0_outputs(476));
    layer1_outputs(780) <= (layer0_outputs(2409)) or (layer0_outputs(2330));
    layer1_outputs(781) <= not(layer0_outputs(151)) or (layer0_outputs(2377));
    layer1_outputs(782) <= (layer0_outputs(1140)) and (layer0_outputs(355));
    layer1_outputs(783) <= not(layer0_outputs(1032)) or (layer0_outputs(336));
    layer1_outputs(784) <= (layer0_outputs(1292)) and (layer0_outputs(685));
    layer1_outputs(785) <= not(layer0_outputs(1745)) or (layer0_outputs(2195));
    layer1_outputs(786) <= layer0_outputs(1567);
    layer1_outputs(787) <= (layer0_outputs(1341)) and not (layer0_outputs(1390));
    layer1_outputs(788) <= not(layer0_outputs(2279)) or (layer0_outputs(832));
    layer1_outputs(789) <= '0';
    layer1_outputs(790) <= '0';
    layer1_outputs(791) <= not(layer0_outputs(1220));
    layer1_outputs(792) <= not((layer0_outputs(1357)) or (layer0_outputs(2427)));
    layer1_outputs(793) <= not((layer0_outputs(1088)) or (layer0_outputs(1703)));
    layer1_outputs(794) <= layer0_outputs(1818);
    layer1_outputs(795) <= '1';
    layer1_outputs(796) <= layer0_outputs(776);
    layer1_outputs(797) <= '0';
    layer1_outputs(798) <= '1';
    layer1_outputs(799) <= layer0_outputs(2004);
    layer1_outputs(800) <= not(layer0_outputs(1591));
    layer1_outputs(801) <= '1';
    layer1_outputs(802) <= (layer0_outputs(2091)) xor (layer0_outputs(585));
    layer1_outputs(803) <= '1';
    layer1_outputs(804) <= not(layer0_outputs(1990));
    layer1_outputs(805) <= not(layer0_outputs(1534)) or (layer0_outputs(474));
    layer1_outputs(806) <= '0';
    layer1_outputs(807) <= '1';
    layer1_outputs(808) <= layer0_outputs(1670);
    layer1_outputs(809) <= not((layer0_outputs(2050)) xor (layer0_outputs(547)));
    layer1_outputs(810) <= '0';
    layer1_outputs(811) <= (layer0_outputs(969)) and not (layer0_outputs(1765));
    layer1_outputs(812) <= '0';
    layer1_outputs(813) <= not((layer0_outputs(1080)) and (layer0_outputs(1253)));
    layer1_outputs(814) <= '1';
    layer1_outputs(815) <= layer0_outputs(1683);
    layer1_outputs(816) <= (layer0_outputs(2299)) and not (layer0_outputs(508));
    layer1_outputs(817) <= (layer0_outputs(2374)) or (layer0_outputs(2078));
    layer1_outputs(818) <= '1';
    layer1_outputs(819) <= (layer0_outputs(2247)) and not (layer0_outputs(767));
    layer1_outputs(820) <= not(layer0_outputs(0));
    layer1_outputs(821) <= layer0_outputs(1567);
    layer1_outputs(822) <= not(layer0_outputs(44)) or (layer0_outputs(755));
    layer1_outputs(823) <= '0';
    layer1_outputs(824) <= not((layer0_outputs(26)) or (layer0_outputs(198)));
    layer1_outputs(825) <= '1';
    layer1_outputs(826) <= layer0_outputs(953);
    layer1_outputs(827) <= not(layer0_outputs(987));
    layer1_outputs(828) <= (layer0_outputs(574)) or (layer0_outputs(2434));
    layer1_outputs(829) <= layer0_outputs(804);
    layer1_outputs(830) <= (layer0_outputs(582)) and not (layer0_outputs(1679));
    layer1_outputs(831) <= not((layer0_outputs(1154)) or (layer0_outputs(589)));
    layer1_outputs(832) <= layer0_outputs(132);
    layer1_outputs(833) <= '0';
    layer1_outputs(834) <= not(layer0_outputs(916)) or (layer0_outputs(1182));
    layer1_outputs(835) <= layer0_outputs(554);
    layer1_outputs(836) <= not((layer0_outputs(96)) or (layer0_outputs(1373)));
    layer1_outputs(837) <= not((layer0_outputs(2356)) or (layer0_outputs(1494)));
    layer1_outputs(838) <= layer0_outputs(144);
    layer1_outputs(839) <= not(layer0_outputs(2235));
    layer1_outputs(840) <= not(layer0_outputs(1888));
    layer1_outputs(841) <= layer0_outputs(2516);
    layer1_outputs(842) <= not(layer0_outputs(228)) or (layer0_outputs(1104));
    layer1_outputs(843) <= '1';
    layer1_outputs(844) <= layer0_outputs(2280);
    layer1_outputs(845) <= not((layer0_outputs(8)) or (layer0_outputs(1538)));
    layer1_outputs(846) <= layer0_outputs(1256);
    layer1_outputs(847) <= (layer0_outputs(740)) and not (layer0_outputs(2416));
    layer1_outputs(848) <= (layer0_outputs(674)) or (layer0_outputs(1857));
    layer1_outputs(849) <= not(layer0_outputs(1394));
    layer1_outputs(850) <= (layer0_outputs(885)) xor (layer0_outputs(1671));
    layer1_outputs(851) <= (layer0_outputs(312)) and not (layer0_outputs(790));
    layer1_outputs(852) <= not(layer0_outputs(1467)) or (layer0_outputs(29));
    layer1_outputs(853) <= layer0_outputs(682);
    layer1_outputs(854) <= not((layer0_outputs(2546)) and (layer0_outputs(1122)));
    layer1_outputs(855) <= not(layer0_outputs(700));
    layer1_outputs(856) <= (layer0_outputs(1758)) and (layer0_outputs(2185));
    layer1_outputs(857) <= not(layer0_outputs(293));
    layer1_outputs(858) <= '0';
    layer1_outputs(859) <= layer0_outputs(1707);
    layer1_outputs(860) <= layer0_outputs(366);
    layer1_outputs(861) <= (layer0_outputs(1556)) and not (layer0_outputs(1106));
    layer1_outputs(862) <= '1';
    layer1_outputs(863) <= '1';
    layer1_outputs(864) <= not(layer0_outputs(2483)) or (layer0_outputs(25));
    layer1_outputs(865) <= '1';
    layer1_outputs(866) <= '1';
    layer1_outputs(867) <= not(layer0_outputs(1282)) or (layer0_outputs(166));
    layer1_outputs(868) <= (layer0_outputs(487)) or (layer0_outputs(1267));
    layer1_outputs(869) <= not((layer0_outputs(1242)) or (layer0_outputs(357)));
    layer1_outputs(870) <= not(layer0_outputs(253));
    layer1_outputs(871) <= not((layer0_outputs(2361)) xor (layer0_outputs(2341)));
    layer1_outputs(872) <= '1';
    layer1_outputs(873) <= (layer0_outputs(483)) and (layer0_outputs(2498));
    layer1_outputs(874) <= (layer0_outputs(413)) and (layer0_outputs(1326));
    layer1_outputs(875) <= '0';
    layer1_outputs(876) <= (layer0_outputs(1429)) and not (layer0_outputs(1074));
    layer1_outputs(877) <= not((layer0_outputs(698)) or (layer0_outputs(2270)));
    layer1_outputs(878) <= (layer0_outputs(910)) and not (layer0_outputs(2459));
    layer1_outputs(879) <= not(layer0_outputs(443)) or (layer0_outputs(1415));
    layer1_outputs(880) <= not(layer0_outputs(1547)) or (layer0_outputs(545));
    layer1_outputs(881) <= (layer0_outputs(610)) or (layer0_outputs(938));
    layer1_outputs(882) <= not(layer0_outputs(828));
    layer1_outputs(883) <= not((layer0_outputs(1875)) or (layer0_outputs(67)));
    layer1_outputs(884) <= '1';
    layer1_outputs(885) <= not(layer0_outputs(992));
    layer1_outputs(886) <= layer0_outputs(131);
    layer1_outputs(887) <= '0';
    layer1_outputs(888) <= '0';
    layer1_outputs(889) <= layer0_outputs(1344);
    layer1_outputs(890) <= '0';
    layer1_outputs(891) <= '1';
    layer1_outputs(892) <= not(layer0_outputs(2469));
    layer1_outputs(893) <= (layer0_outputs(1893)) xor (layer0_outputs(1556));
    layer1_outputs(894) <= not(layer0_outputs(831));
    layer1_outputs(895) <= not((layer0_outputs(419)) and (layer0_outputs(385)));
    layer1_outputs(896) <= '1';
    layer1_outputs(897) <= layer0_outputs(1372);
    layer1_outputs(898) <= '0';
    layer1_outputs(899) <= not(layer0_outputs(769));
    layer1_outputs(900) <= not(layer0_outputs(1244)) or (layer0_outputs(2144));
    layer1_outputs(901) <= (layer0_outputs(364)) and not (layer0_outputs(420));
    layer1_outputs(902) <= (layer0_outputs(786)) or (layer0_outputs(857));
    layer1_outputs(903) <= not(layer0_outputs(1484)) or (layer0_outputs(1098));
    layer1_outputs(904) <= not(layer0_outputs(2238)) or (layer0_outputs(139));
    layer1_outputs(905) <= '1';
    layer1_outputs(906) <= not(layer0_outputs(1787)) or (layer0_outputs(225));
    layer1_outputs(907) <= '0';
    layer1_outputs(908) <= not(layer0_outputs(995));
    layer1_outputs(909) <= not((layer0_outputs(1669)) or (layer0_outputs(164)));
    layer1_outputs(910) <= not(layer0_outputs(1027));
    layer1_outputs(911) <= '0';
    layer1_outputs(912) <= (layer0_outputs(30)) and not (layer0_outputs(1986));
    layer1_outputs(913) <= layer0_outputs(237);
    layer1_outputs(914) <= layer0_outputs(1695);
    layer1_outputs(915) <= layer0_outputs(26);
    layer1_outputs(916) <= not((layer0_outputs(2282)) or (layer0_outputs(2421)));
    layer1_outputs(917) <= layer0_outputs(1722);
    layer1_outputs(918) <= '0';
    layer1_outputs(919) <= not(layer0_outputs(625)) or (layer0_outputs(1250));
    layer1_outputs(920) <= layer0_outputs(1373);
    layer1_outputs(921) <= '0';
    layer1_outputs(922) <= not((layer0_outputs(737)) and (layer0_outputs(745)));
    layer1_outputs(923) <= not(layer0_outputs(2454)) or (layer0_outputs(771));
    layer1_outputs(924) <= (layer0_outputs(1222)) and not (layer0_outputs(769));
    layer1_outputs(925) <= (layer0_outputs(243)) and (layer0_outputs(615));
    layer1_outputs(926) <= (layer0_outputs(664)) and (layer0_outputs(1508));
    layer1_outputs(927) <= layer0_outputs(1758);
    layer1_outputs(928) <= not(layer0_outputs(449));
    layer1_outputs(929) <= not(layer0_outputs(2027));
    layer1_outputs(930) <= (layer0_outputs(2247)) and (layer0_outputs(1737));
    layer1_outputs(931) <= layer0_outputs(1214);
    layer1_outputs(932) <= (layer0_outputs(692)) and not (layer0_outputs(2083));
    layer1_outputs(933) <= (layer0_outputs(1326)) and not (layer0_outputs(863));
    layer1_outputs(934) <= not(layer0_outputs(594));
    layer1_outputs(935) <= layer0_outputs(2324);
    layer1_outputs(936) <= not(layer0_outputs(982)) or (layer0_outputs(847));
    layer1_outputs(937) <= layer0_outputs(479);
    layer1_outputs(938) <= (layer0_outputs(1283)) and not (layer0_outputs(458));
    layer1_outputs(939) <= not((layer0_outputs(563)) and (layer0_outputs(1888)));
    layer1_outputs(940) <= not(layer0_outputs(1850));
    layer1_outputs(941) <= not((layer0_outputs(2285)) or (layer0_outputs(1061)));
    layer1_outputs(942) <= (layer0_outputs(1378)) or (layer0_outputs(679));
    layer1_outputs(943) <= not(layer0_outputs(245));
    layer1_outputs(944) <= '1';
    layer1_outputs(945) <= not(layer0_outputs(462));
    layer1_outputs(946) <= not(layer0_outputs(829));
    layer1_outputs(947) <= layer0_outputs(1744);
    layer1_outputs(948) <= not(layer0_outputs(308)) or (layer0_outputs(906));
    layer1_outputs(949) <= (layer0_outputs(1496)) and (layer0_outputs(1747));
    layer1_outputs(950) <= not((layer0_outputs(19)) or (layer0_outputs(300)));
    layer1_outputs(951) <= not((layer0_outputs(1019)) xor (layer0_outputs(908)));
    layer1_outputs(952) <= layer0_outputs(1495);
    layer1_outputs(953) <= not(layer0_outputs(1291));
    layer1_outputs(954) <= not((layer0_outputs(2515)) or (layer0_outputs(893)));
    layer1_outputs(955) <= (layer0_outputs(2464)) and not (layer0_outputs(2468));
    layer1_outputs(956) <= '0';
    layer1_outputs(957) <= layer0_outputs(2540);
    layer1_outputs(958) <= not(layer0_outputs(892));
    layer1_outputs(959) <= (layer0_outputs(723)) or (layer0_outputs(739));
    layer1_outputs(960) <= '0';
    layer1_outputs(961) <= not(layer0_outputs(2238));
    layer1_outputs(962) <= not(layer0_outputs(2326)) or (layer0_outputs(255));
    layer1_outputs(963) <= not((layer0_outputs(478)) or (layer0_outputs(540)));
    layer1_outputs(964) <= not(layer0_outputs(82));
    layer1_outputs(965) <= (layer0_outputs(1029)) or (layer0_outputs(1835));
    layer1_outputs(966) <= layer0_outputs(819);
    layer1_outputs(967) <= (layer0_outputs(1223)) and not (layer0_outputs(492));
    layer1_outputs(968) <= not((layer0_outputs(9)) and (layer0_outputs(372)));
    layer1_outputs(969) <= '0';
    layer1_outputs(970) <= '1';
    layer1_outputs(971) <= layer0_outputs(1037);
    layer1_outputs(972) <= (layer0_outputs(1301)) and (layer0_outputs(1418));
    layer1_outputs(973) <= '0';
    layer1_outputs(974) <= '0';
    layer1_outputs(975) <= not(layer0_outputs(2537));
    layer1_outputs(976) <= (layer0_outputs(550)) and not (layer0_outputs(2081));
    layer1_outputs(977) <= not(layer0_outputs(2424)) or (layer0_outputs(148));
    layer1_outputs(978) <= not((layer0_outputs(2191)) and (layer0_outputs(93)));
    layer1_outputs(979) <= not(layer0_outputs(1297)) or (layer0_outputs(2260));
    layer1_outputs(980) <= (layer0_outputs(2282)) or (layer0_outputs(1331));
    layer1_outputs(981) <= (layer0_outputs(2401)) and not (layer0_outputs(1098));
    layer1_outputs(982) <= '1';
    layer1_outputs(983) <= (layer0_outputs(554)) and not (layer0_outputs(1473));
    layer1_outputs(984) <= layer0_outputs(1868);
    layer1_outputs(985) <= not((layer0_outputs(1086)) and (layer0_outputs(439)));
    layer1_outputs(986) <= not((layer0_outputs(265)) or (layer0_outputs(1041)));
    layer1_outputs(987) <= not(layer0_outputs(968));
    layer1_outputs(988) <= not(layer0_outputs(1881)) or (layer0_outputs(2081));
    layer1_outputs(989) <= layer0_outputs(2304);
    layer1_outputs(990) <= (layer0_outputs(2298)) and (layer0_outputs(778));
    layer1_outputs(991) <= not((layer0_outputs(794)) or (layer0_outputs(609)));
    layer1_outputs(992) <= '1';
    layer1_outputs(993) <= (layer0_outputs(1994)) or (layer0_outputs(594));
    layer1_outputs(994) <= layer0_outputs(362);
    layer1_outputs(995) <= layer0_outputs(2548);
    layer1_outputs(996) <= '1';
    layer1_outputs(997) <= '0';
    layer1_outputs(998) <= not(layer0_outputs(1575));
    layer1_outputs(999) <= not(layer0_outputs(1662));
    layer1_outputs(1000) <= not(layer0_outputs(1762));
    layer1_outputs(1001) <= not(layer0_outputs(2352)) or (layer0_outputs(2163));
    layer1_outputs(1002) <= '0';
    layer1_outputs(1003) <= not(layer0_outputs(2325)) or (layer0_outputs(946));
    layer1_outputs(1004) <= (layer0_outputs(2098)) and not (layer0_outputs(1596));
    layer1_outputs(1005) <= (layer0_outputs(1549)) or (layer0_outputs(1986));
    layer1_outputs(1006) <= not((layer0_outputs(1101)) and (layer0_outputs(2135)));
    layer1_outputs(1007) <= (layer0_outputs(1979)) and not (layer0_outputs(302));
    layer1_outputs(1008) <= layer0_outputs(1305);
    layer1_outputs(1009) <= (layer0_outputs(2386)) and not (layer0_outputs(1050));
    layer1_outputs(1010) <= not((layer0_outputs(1168)) and (layer0_outputs(358)));
    layer1_outputs(1011) <= '0';
    layer1_outputs(1012) <= '0';
    layer1_outputs(1013) <= (layer0_outputs(1906)) and (layer0_outputs(977));
    layer1_outputs(1014) <= not((layer0_outputs(961)) or (layer0_outputs(59)));
    layer1_outputs(1015) <= not((layer0_outputs(276)) xor (layer0_outputs(1989)));
    layer1_outputs(1016) <= '0';
    layer1_outputs(1017) <= '0';
    layer1_outputs(1018) <= not(layer0_outputs(1192)) or (layer0_outputs(1319));
    layer1_outputs(1019) <= layer0_outputs(2148);
    layer1_outputs(1020) <= (layer0_outputs(1123)) or (layer0_outputs(2545));
    layer1_outputs(1021) <= layer0_outputs(914);
    layer1_outputs(1022) <= (layer0_outputs(120)) or (layer0_outputs(1532));
    layer1_outputs(1023) <= not(layer0_outputs(768)) or (layer0_outputs(1791));
    layer1_outputs(1024) <= not(layer0_outputs(1544)) or (layer0_outputs(214));
    layer1_outputs(1025) <= '1';
    layer1_outputs(1026) <= (layer0_outputs(1134)) xor (layer0_outputs(918));
    layer1_outputs(1027) <= layer0_outputs(598);
    layer1_outputs(1028) <= not(layer0_outputs(472)) or (layer0_outputs(2363));
    layer1_outputs(1029) <= not(layer0_outputs(1804));
    layer1_outputs(1030) <= (layer0_outputs(1743)) and not (layer0_outputs(1355));
    layer1_outputs(1031) <= not(layer0_outputs(54));
    layer1_outputs(1032) <= not(layer0_outputs(1383));
    layer1_outputs(1033) <= not((layer0_outputs(593)) or (layer0_outputs(1586)));
    layer1_outputs(1034) <= (layer0_outputs(762)) and not (layer0_outputs(2258));
    layer1_outputs(1035) <= (layer0_outputs(991)) or (layer0_outputs(1408));
    layer1_outputs(1036) <= (layer0_outputs(734)) and not (layer0_outputs(936));
    layer1_outputs(1037) <= (layer0_outputs(1891)) and not (layer0_outputs(2361));
    layer1_outputs(1038) <= not(layer0_outputs(2253));
    layer1_outputs(1039) <= not(layer0_outputs(736)) or (layer0_outputs(2023));
    layer1_outputs(1040) <= layer0_outputs(1981);
    layer1_outputs(1041) <= (layer0_outputs(185)) xor (layer0_outputs(1115));
    layer1_outputs(1042) <= not(layer0_outputs(1898));
    layer1_outputs(1043) <= layer0_outputs(223);
    layer1_outputs(1044) <= layer0_outputs(549);
    layer1_outputs(1045) <= (layer0_outputs(647)) and not (layer0_outputs(1410));
    layer1_outputs(1046) <= '1';
    layer1_outputs(1047) <= (layer0_outputs(2191)) and not (layer0_outputs(1073));
    layer1_outputs(1048) <= not(layer0_outputs(1320)) or (layer0_outputs(1843));
    layer1_outputs(1049) <= not((layer0_outputs(298)) or (layer0_outputs(2280)));
    layer1_outputs(1050) <= (layer0_outputs(76)) or (layer0_outputs(2144));
    layer1_outputs(1051) <= not((layer0_outputs(191)) or (layer0_outputs(1844)));
    layer1_outputs(1052) <= not(layer0_outputs(675));
    layer1_outputs(1053) <= (layer0_outputs(1957)) or (layer0_outputs(809));
    layer1_outputs(1054) <= '0';
    layer1_outputs(1055) <= layer0_outputs(823);
    layer1_outputs(1056) <= (layer0_outputs(384)) and not (layer0_outputs(1431));
    layer1_outputs(1057) <= layer0_outputs(1058);
    layer1_outputs(1058) <= not(layer0_outputs(1842)) or (layer0_outputs(1689));
    layer1_outputs(1059) <= (layer0_outputs(1537)) and (layer0_outputs(1117));
    layer1_outputs(1060) <= (layer0_outputs(1388)) or (layer0_outputs(796));
    layer1_outputs(1061) <= (layer0_outputs(2056)) and not (layer0_outputs(1137));
    layer1_outputs(1062) <= '0';
    layer1_outputs(1063) <= not(layer0_outputs(1442)) or (layer0_outputs(1234));
    layer1_outputs(1064) <= not(layer0_outputs(1616)) or (layer0_outputs(1423));
    layer1_outputs(1065) <= '1';
    layer1_outputs(1066) <= not(layer0_outputs(2054));
    layer1_outputs(1067) <= (layer0_outputs(46)) or (layer0_outputs(1312));
    layer1_outputs(1068) <= (layer0_outputs(2202)) and not (layer0_outputs(2015));
    layer1_outputs(1069) <= '1';
    layer1_outputs(1070) <= (layer0_outputs(1609)) and not (layer0_outputs(791));
    layer1_outputs(1071) <= (layer0_outputs(1002)) and (layer0_outputs(957));
    layer1_outputs(1072) <= '0';
    layer1_outputs(1073) <= not(layer0_outputs(2383)) or (layer0_outputs(37));
    layer1_outputs(1074) <= not((layer0_outputs(105)) or (layer0_outputs(2091)));
    layer1_outputs(1075) <= (layer0_outputs(2328)) and (layer0_outputs(538));
    layer1_outputs(1076) <= (layer0_outputs(2184)) or (layer0_outputs(1963));
    layer1_outputs(1077) <= '1';
    layer1_outputs(1078) <= (layer0_outputs(493)) and not (layer0_outputs(65));
    layer1_outputs(1079) <= '1';
    layer1_outputs(1080) <= (layer0_outputs(2432)) or (layer0_outputs(3));
    layer1_outputs(1081) <= layer0_outputs(878);
    layer1_outputs(1082) <= '0';
    layer1_outputs(1083) <= not((layer0_outputs(748)) and (layer0_outputs(1977)));
    layer1_outputs(1084) <= '0';
    layer1_outputs(1085) <= not(layer0_outputs(2182)) or (layer0_outputs(1858));
    layer1_outputs(1086) <= '1';
    layer1_outputs(1087) <= '0';
    layer1_outputs(1088) <= (layer0_outputs(1498)) and (layer0_outputs(2340));
    layer1_outputs(1089) <= layer0_outputs(1252);
    layer1_outputs(1090) <= '0';
    layer1_outputs(1091) <= (layer0_outputs(1795)) and not (layer0_outputs(2515));
    layer1_outputs(1092) <= (layer0_outputs(2533)) and (layer0_outputs(383));
    layer1_outputs(1093) <= '1';
    layer1_outputs(1094) <= not(layer0_outputs(777));
    layer1_outputs(1095) <= not(layer0_outputs(1340));
    layer1_outputs(1096) <= not(layer0_outputs(1906));
    layer1_outputs(1097) <= (layer0_outputs(1928)) or (layer0_outputs(2098));
    layer1_outputs(1098) <= (layer0_outputs(915)) and (layer0_outputs(1130));
    layer1_outputs(1099) <= (layer0_outputs(2456)) and not (layer0_outputs(914));
    layer1_outputs(1100) <= '1';
    layer1_outputs(1101) <= (layer0_outputs(2187)) and not (layer0_outputs(93));
    layer1_outputs(1102) <= '1';
    layer1_outputs(1103) <= (layer0_outputs(657)) and (layer0_outputs(1293));
    layer1_outputs(1104) <= not((layer0_outputs(1392)) or (layer0_outputs(394)));
    layer1_outputs(1105) <= '0';
    layer1_outputs(1106) <= not(layer0_outputs(628));
    layer1_outputs(1107) <= not((layer0_outputs(1630)) or (layer0_outputs(2052)));
    layer1_outputs(1108) <= not(layer0_outputs(1174)) or (layer0_outputs(487));
    layer1_outputs(1109) <= not((layer0_outputs(1486)) and (layer0_outputs(1479)));
    layer1_outputs(1110) <= not(layer0_outputs(2204)) or (layer0_outputs(348));
    layer1_outputs(1111) <= (layer0_outputs(2402)) or (layer0_outputs(713));
    layer1_outputs(1112) <= not(layer0_outputs(2127)) or (layer0_outputs(421));
    layer1_outputs(1113) <= (layer0_outputs(1241)) and not (layer0_outputs(1624));
    layer1_outputs(1114) <= layer0_outputs(100);
    layer1_outputs(1115) <= '1';
    layer1_outputs(1116) <= not(layer0_outputs(522)) or (layer0_outputs(237));
    layer1_outputs(1117) <= '0';
    layer1_outputs(1118) <= (layer0_outputs(2511)) and not (layer0_outputs(1471));
    layer1_outputs(1119) <= not(layer0_outputs(862));
    layer1_outputs(1120) <= '0';
    layer1_outputs(1121) <= not(layer0_outputs(459)) or (layer0_outputs(1020));
    layer1_outputs(1122) <= layer0_outputs(38);
    layer1_outputs(1123) <= (layer0_outputs(1970)) or (layer0_outputs(766));
    layer1_outputs(1124) <= not(layer0_outputs(470)) or (layer0_outputs(2379));
    layer1_outputs(1125) <= not(layer0_outputs(1948));
    layer1_outputs(1126) <= layer0_outputs(1878);
    layer1_outputs(1127) <= not(layer0_outputs(2390));
    layer1_outputs(1128) <= not((layer0_outputs(391)) and (layer0_outputs(1145)));
    layer1_outputs(1129) <= '0';
    layer1_outputs(1130) <= '0';
    layer1_outputs(1131) <= (layer0_outputs(675)) and (layer0_outputs(1763));
    layer1_outputs(1132) <= '0';
    layer1_outputs(1133) <= not(layer0_outputs(268)) or (layer0_outputs(2195));
    layer1_outputs(1134) <= not(layer0_outputs(412));
    layer1_outputs(1135) <= layer0_outputs(2225);
    layer1_outputs(1136) <= '1';
    layer1_outputs(1137) <= not((layer0_outputs(1391)) or (layer0_outputs(2013)));
    layer1_outputs(1138) <= not(layer0_outputs(758));
    layer1_outputs(1139) <= not(layer0_outputs(1820));
    layer1_outputs(1140) <= not(layer0_outputs(129));
    layer1_outputs(1141) <= not(layer0_outputs(1106));
    layer1_outputs(1142) <= not(layer0_outputs(1064));
    layer1_outputs(1143) <= not(layer0_outputs(2519)) or (layer0_outputs(1191));
    layer1_outputs(1144) <= (layer0_outputs(1091)) and not (layer0_outputs(704));
    layer1_outputs(1145) <= not((layer0_outputs(473)) or (layer0_outputs(1179)));
    layer1_outputs(1146) <= layer0_outputs(296);
    layer1_outputs(1147) <= layer0_outputs(1748);
    layer1_outputs(1148) <= '1';
    layer1_outputs(1149) <= not((layer0_outputs(1065)) and (layer0_outputs(610)));
    layer1_outputs(1150) <= '0';
    layer1_outputs(1151) <= not(layer0_outputs(1093)) or (layer0_outputs(392));
    layer1_outputs(1152) <= (layer0_outputs(2329)) and not (layer0_outputs(941));
    layer1_outputs(1153) <= layer0_outputs(2439);
    layer1_outputs(1154) <= not(layer0_outputs(1856)) or (layer0_outputs(877));
    layer1_outputs(1155) <= not(layer0_outputs(567)) or (layer0_outputs(2476));
    layer1_outputs(1156) <= not(layer0_outputs(1550));
    layer1_outputs(1157) <= not(layer0_outputs(2387));
    layer1_outputs(1158) <= not((layer0_outputs(1383)) and (layer0_outputs(158)));
    layer1_outputs(1159) <= '0';
    layer1_outputs(1160) <= not(layer0_outputs(670)) or (layer0_outputs(1362));
    layer1_outputs(1161) <= (layer0_outputs(1831)) and not (layer0_outputs(2481));
    layer1_outputs(1162) <= (layer0_outputs(262)) and not (layer0_outputs(2082));
    layer1_outputs(1163) <= (layer0_outputs(2445)) and not (layer0_outputs(1659));
    layer1_outputs(1164) <= not((layer0_outputs(2068)) xor (layer0_outputs(2021)));
    layer1_outputs(1165) <= '1';
    layer1_outputs(1166) <= layer0_outputs(2065);
    layer1_outputs(1167) <= not(layer0_outputs(2303));
    layer1_outputs(1168) <= not(layer0_outputs(1649)) or (layer0_outputs(2037));
    layer1_outputs(1169) <= not((layer0_outputs(1914)) and (layer0_outputs(2269)));
    layer1_outputs(1170) <= not((layer0_outputs(1793)) and (layer0_outputs(2221)));
    layer1_outputs(1171) <= (layer0_outputs(1806)) and not (layer0_outputs(1273));
    layer1_outputs(1172) <= (layer0_outputs(2338)) and not (layer0_outputs(1274));
    layer1_outputs(1173) <= not((layer0_outputs(848)) and (layer0_outputs(1261)));
    layer1_outputs(1174) <= '1';
    layer1_outputs(1175) <= not(layer0_outputs(1005)) or (layer0_outputs(2043));
    layer1_outputs(1176) <= not(layer0_outputs(1895));
    layer1_outputs(1177) <= not(layer0_outputs(2003));
    layer1_outputs(1178) <= not((layer0_outputs(1992)) or (layer0_outputs(342)));
    layer1_outputs(1179) <= (layer0_outputs(1259)) and not (layer0_outputs(99));
    layer1_outputs(1180) <= layer0_outputs(1865);
    layer1_outputs(1181) <= not(layer0_outputs(2283)) or (layer0_outputs(2553));
    layer1_outputs(1182) <= layer0_outputs(288);
    layer1_outputs(1183) <= not((layer0_outputs(636)) and (layer0_outputs(437)));
    layer1_outputs(1184) <= (layer0_outputs(1794)) and not (layer0_outputs(2479));
    layer1_outputs(1185) <= not(layer0_outputs(1979)) or (layer0_outputs(652));
    layer1_outputs(1186) <= (layer0_outputs(2255)) and (layer0_outputs(1082));
    layer1_outputs(1187) <= not(layer0_outputs(803)) or (layer0_outputs(686));
    layer1_outputs(1188) <= '1';
    layer1_outputs(1189) <= not(layer0_outputs(1680));
    layer1_outputs(1190) <= layer0_outputs(950);
    layer1_outputs(1191) <= layer0_outputs(2302);
    layer1_outputs(1192) <= not(layer0_outputs(1767));
    layer1_outputs(1193) <= not(layer0_outputs(1943)) or (layer0_outputs(1327));
    layer1_outputs(1194) <= not(layer0_outputs(533));
    layer1_outputs(1195) <= not((layer0_outputs(1330)) and (layer0_outputs(1324)));
    layer1_outputs(1196) <= '0';
    layer1_outputs(1197) <= not(layer0_outputs(81));
    layer1_outputs(1198) <= (layer0_outputs(2285)) and (layer0_outputs(501));
    layer1_outputs(1199) <= '1';
    layer1_outputs(1200) <= not(layer0_outputs(833));
    layer1_outputs(1201) <= (layer0_outputs(1694)) and not (layer0_outputs(2503));
    layer1_outputs(1202) <= (layer0_outputs(937)) and (layer0_outputs(519));
    layer1_outputs(1203) <= layer0_outputs(1099);
    layer1_outputs(1204) <= not((layer0_outputs(2029)) and (layer0_outputs(1047)));
    layer1_outputs(1205) <= not(layer0_outputs(1837));
    layer1_outputs(1206) <= not((layer0_outputs(1126)) and (layer0_outputs(1057)));
    layer1_outputs(1207) <= not(layer0_outputs(673));
    layer1_outputs(1208) <= not(layer0_outputs(2429)) or (layer0_outputs(1376));
    layer1_outputs(1209) <= layer0_outputs(194);
    layer1_outputs(1210) <= not(layer0_outputs(2539));
    layer1_outputs(1211) <= (layer0_outputs(1225)) and not (layer0_outputs(1907));
    layer1_outputs(1212) <= (layer0_outputs(2241)) and not (layer0_outputs(2525));
    layer1_outputs(1213) <= '1';
    layer1_outputs(1214) <= layer0_outputs(956);
    layer1_outputs(1215) <= '0';
    layer1_outputs(1216) <= not(layer0_outputs(95));
    layer1_outputs(1217) <= (layer0_outputs(905)) or (layer0_outputs(923));
    layer1_outputs(1218) <= (layer0_outputs(1947)) and not (layer0_outputs(661));
    layer1_outputs(1219) <= '0';
    layer1_outputs(1220) <= '0';
    layer1_outputs(1221) <= layer0_outputs(1746);
    layer1_outputs(1222) <= '1';
    layer1_outputs(1223) <= not(layer0_outputs(1030));
    layer1_outputs(1224) <= (layer0_outputs(2442)) and (layer0_outputs(2275));
    layer1_outputs(1225) <= not(layer0_outputs(1038));
    layer1_outputs(1226) <= not(layer0_outputs(341)) or (layer0_outputs(1512));
    layer1_outputs(1227) <= not(layer0_outputs(2041));
    layer1_outputs(1228) <= '0';
    layer1_outputs(1229) <= not(layer0_outputs(2278));
    layer1_outputs(1230) <= '1';
    layer1_outputs(1231) <= (layer0_outputs(501)) and (layer0_outputs(1612));
    layer1_outputs(1232) <= not(layer0_outputs(1277));
    layer1_outputs(1233) <= not((layer0_outputs(213)) or (layer0_outputs(2527)));
    layer1_outputs(1234) <= '1';
    layer1_outputs(1235) <= not(layer0_outputs(1949));
    layer1_outputs(1236) <= '0';
    layer1_outputs(1237) <= not(layer0_outputs(595));
    layer1_outputs(1238) <= '1';
    layer1_outputs(1239) <= (layer0_outputs(1039)) and not (layer0_outputs(2465));
    layer1_outputs(1240) <= '1';
    layer1_outputs(1241) <= not(layer0_outputs(1139)) or (layer0_outputs(2151));
    layer1_outputs(1242) <= (layer0_outputs(2532)) xor (layer0_outputs(968));
    layer1_outputs(1243) <= not(layer0_outputs(1965));
    layer1_outputs(1244) <= '1';
    layer1_outputs(1245) <= '0';
    layer1_outputs(1246) <= not((layer0_outputs(1457)) or (layer0_outputs(850)));
    layer1_outputs(1247) <= (layer0_outputs(1458)) and not (layer0_outputs(2342));
    layer1_outputs(1248) <= not((layer0_outputs(1511)) or (layer0_outputs(899)));
    layer1_outputs(1249) <= '1';
    layer1_outputs(1250) <= not((layer0_outputs(1065)) or (layer0_outputs(2161)));
    layer1_outputs(1251) <= (layer0_outputs(1335)) and not (layer0_outputs(150));
    layer1_outputs(1252) <= (layer0_outputs(1087)) and not (layer0_outputs(1509));
    layer1_outputs(1253) <= '1';
    layer1_outputs(1254) <= (layer0_outputs(1647)) and (layer0_outputs(2218));
    layer1_outputs(1255) <= '1';
    layer1_outputs(1256) <= '1';
    layer1_outputs(1257) <= not(layer0_outputs(1974));
    layer1_outputs(1258) <= (layer0_outputs(768)) and (layer0_outputs(133));
    layer1_outputs(1259) <= not(layer0_outputs(448)) or (layer0_outputs(623));
    layer1_outputs(1260) <= '1';
    layer1_outputs(1261) <= layer0_outputs(1051);
    layer1_outputs(1262) <= not(layer0_outputs(1151)) or (layer0_outputs(1852));
    layer1_outputs(1263) <= layer0_outputs(2356);
    layer1_outputs(1264) <= not(layer0_outputs(978)) or (layer0_outputs(807));
    layer1_outputs(1265) <= (layer0_outputs(1145)) and not (layer0_outputs(1750));
    layer1_outputs(1266) <= not((layer0_outputs(2444)) or (layer0_outputs(907)));
    layer1_outputs(1267) <= not(layer0_outputs(1102));
    layer1_outputs(1268) <= '0';
    layer1_outputs(1269) <= (layer0_outputs(1678)) and not (layer0_outputs(1023));
    layer1_outputs(1270) <= layer0_outputs(901);
    layer1_outputs(1271) <= not(layer0_outputs(58));
    layer1_outputs(1272) <= not(layer0_outputs(1452)) or (layer0_outputs(957));
    layer1_outputs(1273) <= layer0_outputs(917);
    layer1_outputs(1274) <= layer0_outputs(207);
    layer1_outputs(1275) <= '0';
    layer1_outputs(1276) <= not((layer0_outputs(250)) and (layer0_outputs(2347)));
    layer1_outputs(1277) <= (layer0_outputs(1781)) and not (layer0_outputs(2047));
    layer1_outputs(1278) <= layer0_outputs(449);
    layer1_outputs(1279) <= not(layer0_outputs(1674)) or (layer0_outputs(1666));
    layer1_outputs(1280) <= not((layer0_outputs(1035)) and (layer0_outputs(1883)));
    layer1_outputs(1281) <= layer0_outputs(2283);
    layer1_outputs(1282) <= not((layer0_outputs(2417)) or (layer0_outputs(1208)));
    layer1_outputs(1283) <= not((layer0_outputs(1469)) xor (layer0_outputs(2200)));
    layer1_outputs(1284) <= '0';
    layer1_outputs(1285) <= '0';
    layer1_outputs(1286) <= '0';
    layer1_outputs(1287) <= not(layer0_outputs(1527));
    layer1_outputs(1288) <= layer0_outputs(1948);
    layer1_outputs(1289) <= not(layer0_outputs(2092));
    layer1_outputs(1290) <= not(layer0_outputs(496)) or (layer0_outputs(1604));
    layer1_outputs(1291) <= '1';
    layer1_outputs(1292) <= (layer0_outputs(1717)) and not (layer0_outputs(1580));
    layer1_outputs(1293) <= not(layer0_outputs(1407));
    layer1_outputs(1294) <= not(layer0_outputs(1879)) or (layer0_outputs(2024));
    layer1_outputs(1295) <= '1';
    layer1_outputs(1296) <= layer0_outputs(1558);
    layer1_outputs(1297) <= layer0_outputs(2003);
    layer1_outputs(1298) <= not(layer0_outputs(1654));
    layer1_outputs(1299) <= (layer0_outputs(2292)) and not (layer0_outputs(701));
    layer1_outputs(1300) <= '1';
    layer1_outputs(1301) <= layer0_outputs(431);
    layer1_outputs(1302) <= not(layer0_outputs(192)) or (layer0_outputs(719));
    layer1_outputs(1303) <= '1';
    layer1_outputs(1304) <= layer0_outputs(1386);
    layer1_outputs(1305) <= not(layer0_outputs(764));
    layer1_outputs(1306) <= (layer0_outputs(573)) or (layer0_outputs(2549));
    layer1_outputs(1307) <= '1';
    layer1_outputs(1308) <= (layer0_outputs(892)) and not (layer0_outputs(1133));
    layer1_outputs(1309) <= layer0_outputs(36);
    layer1_outputs(1310) <= (layer0_outputs(1432)) and not (layer0_outputs(620));
    layer1_outputs(1311) <= layer0_outputs(158);
    layer1_outputs(1312) <= (layer0_outputs(1759)) and not (layer0_outputs(2256));
    layer1_outputs(1313) <= layer0_outputs(72);
    layer1_outputs(1314) <= not(layer0_outputs(2538)) or (layer0_outputs(216));
    layer1_outputs(1315) <= not(layer0_outputs(620));
    layer1_outputs(1316) <= not((layer0_outputs(125)) or (layer0_outputs(1607)));
    layer1_outputs(1317) <= layer0_outputs(2362);
    layer1_outputs(1318) <= '0';
    layer1_outputs(1319) <= '0';
    layer1_outputs(1320) <= (layer0_outputs(1436)) and not (layer0_outputs(1056));
    layer1_outputs(1321) <= (layer0_outputs(305)) and not (layer0_outputs(835));
    layer1_outputs(1322) <= (layer0_outputs(648)) and not (layer0_outputs(1528));
    layer1_outputs(1323) <= '0';
    layer1_outputs(1324) <= (layer0_outputs(1802)) and (layer0_outputs(1295));
    layer1_outputs(1325) <= (layer0_outputs(19)) and (layer0_outputs(2351));
    layer1_outputs(1326) <= '0';
    layer1_outputs(1327) <= (layer0_outputs(961)) and (layer0_outputs(995));
    layer1_outputs(1328) <= not(layer0_outputs(146));
    layer1_outputs(1329) <= not(layer0_outputs(2134)) or (layer0_outputs(291));
    layer1_outputs(1330) <= '1';
    layer1_outputs(1331) <= (layer0_outputs(590)) and not (layer0_outputs(217));
    layer1_outputs(1332) <= not(layer0_outputs(142));
    layer1_outputs(1333) <= (layer0_outputs(1235)) or (layer0_outputs(1929));
    layer1_outputs(1334) <= (layer0_outputs(1405)) and (layer0_outputs(756));
    layer1_outputs(1335) <= not((layer0_outputs(1626)) or (layer0_outputs(2430)));
    layer1_outputs(1336) <= layer0_outputs(1939);
    layer1_outputs(1337) <= (layer0_outputs(1146)) and not (layer0_outputs(58));
    layer1_outputs(1338) <= not(layer0_outputs(960));
    layer1_outputs(1339) <= not(layer0_outputs(702));
    layer1_outputs(1340) <= not(layer0_outputs(1266));
    layer1_outputs(1341) <= not(layer0_outputs(1787));
    layer1_outputs(1342) <= (layer0_outputs(503)) or (layer0_outputs(2425));
    layer1_outputs(1343) <= (layer0_outputs(1089)) and (layer0_outputs(2441));
    layer1_outputs(1344) <= not((layer0_outputs(2095)) and (layer0_outputs(635)));
    layer1_outputs(1345) <= (layer0_outputs(2346)) and not (layer0_outputs(467));
    layer1_outputs(1346) <= not(layer0_outputs(1715));
    layer1_outputs(1347) <= layer0_outputs(2422);
    layer1_outputs(1348) <= '0';
    layer1_outputs(1349) <= '1';
    layer1_outputs(1350) <= not(layer0_outputs(1503)) or (layer0_outputs(88));
    layer1_outputs(1351) <= layer0_outputs(1220);
    layer1_outputs(1352) <= (layer0_outputs(580)) and not (layer0_outputs(1239));
    layer1_outputs(1353) <= not((layer0_outputs(925)) and (layer0_outputs(361)));
    layer1_outputs(1354) <= layer0_outputs(1018);
    layer1_outputs(1355) <= '0';
    layer1_outputs(1356) <= (layer0_outputs(570)) and not (layer0_outputs(368));
    layer1_outputs(1357) <= '0';
    layer1_outputs(1358) <= '1';
    layer1_outputs(1359) <= not(layer0_outputs(2395)) or (layer0_outputs(150));
    layer1_outputs(1360) <= not(layer0_outputs(1876)) or (layer0_outputs(734));
    layer1_outputs(1361) <= '1';
    layer1_outputs(1362) <= layer0_outputs(1634);
    layer1_outputs(1363) <= layer0_outputs(162);
    layer1_outputs(1364) <= '0';
    layer1_outputs(1365) <= layer0_outputs(1774);
    layer1_outputs(1366) <= not(layer0_outputs(518));
    layer1_outputs(1367) <= not(layer0_outputs(109));
    layer1_outputs(1368) <= not((layer0_outputs(2071)) and (layer0_outputs(2446)));
    layer1_outputs(1369) <= (layer0_outputs(46)) and not (layer0_outputs(2082));
    layer1_outputs(1370) <= not(layer0_outputs(1754));
    layer1_outputs(1371) <= not(layer0_outputs(2318));
    layer1_outputs(1372) <= not((layer0_outputs(426)) xor (layer0_outputs(1112)));
    layer1_outputs(1373) <= (layer0_outputs(900)) and (layer0_outputs(883));
    layer1_outputs(1374) <= not(layer0_outputs(2072)) or (layer0_outputs(1975));
    layer1_outputs(1375) <= '1';
    layer1_outputs(1376) <= not(layer0_outputs(1601)) or (layer0_outputs(568));
    layer1_outputs(1377) <= (layer0_outputs(652)) and not (layer0_outputs(873));
    layer1_outputs(1378) <= not(layer0_outputs(1855));
    layer1_outputs(1379) <= (layer0_outputs(2545)) or (layer0_outputs(1937));
    layer1_outputs(1380) <= (layer0_outputs(1076)) or (layer0_outputs(1021));
    layer1_outputs(1381) <= layer0_outputs(1294);
    layer1_outputs(1382) <= not((layer0_outputs(2176)) or (layer0_outputs(2084)));
    layer1_outputs(1383) <= not(layer0_outputs(556));
    layer1_outputs(1384) <= not((layer0_outputs(1954)) or (layer0_outputs(2360)));
    layer1_outputs(1385) <= not(layer0_outputs(2484)) or (layer0_outputs(2533));
    layer1_outputs(1386) <= not((layer0_outputs(662)) or (layer0_outputs(1701)));
    layer1_outputs(1387) <= not(layer0_outputs(130));
    layer1_outputs(1388) <= (layer0_outputs(448)) and not (layer0_outputs(2554));
    layer1_outputs(1389) <= not(layer0_outputs(55));
    layer1_outputs(1390) <= (layer0_outputs(2499)) and not (layer0_outputs(2007));
    layer1_outputs(1391) <= '0';
    layer1_outputs(1392) <= not((layer0_outputs(467)) and (layer0_outputs(1570)));
    layer1_outputs(1393) <= not(layer0_outputs(1775)) or (layer0_outputs(1445));
    layer1_outputs(1394) <= '0';
    layer1_outputs(1395) <= not(layer0_outputs(1316));
    layer1_outputs(1396) <= not((layer0_outputs(20)) or (layer0_outputs(1136)));
    layer1_outputs(1397) <= '0';
    layer1_outputs(1398) <= (layer0_outputs(2404)) and (layer0_outputs(2557));
    layer1_outputs(1399) <= layer0_outputs(2339);
    layer1_outputs(1400) <= (layer0_outputs(1887)) and not (layer0_outputs(263));
    layer1_outputs(1401) <= not(layer0_outputs(1915));
    layer1_outputs(1402) <= not((layer0_outputs(18)) xor (layer0_outputs(2341)));
    layer1_outputs(1403) <= not(layer0_outputs(397)) or (layer0_outputs(447));
    layer1_outputs(1404) <= not(layer0_outputs(21)) or (layer0_outputs(514));
    layer1_outputs(1405) <= layer0_outputs(110);
    layer1_outputs(1406) <= not(layer0_outputs(38));
    layer1_outputs(1407) <= '0';
    layer1_outputs(1408) <= not((layer0_outputs(201)) xor (layer0_outputs(248)));
    layer1_outputs(1409) <= (layer0_outputs(493)) and not (layer0_outputs(190));
    layer1_outputs(1410) <= not((layer0_outputs(2332)) or (layer0_outputs(822)));
    layer1_outputs(1411) <= layer0_outputs(34);
    layer1_outputs(1412) <= (layer0_outputs(142)) and (layer0_outputs(1690));
    layer1_outputs(1413) <= (layer0_outputs(986)) or (layer0_outputs(1457));
    layer1_outputs(1414) <= (layer0_outputs(2296)) and not (layer0_outputs(588));
    layer1_outputs(1415) <= not(layer0_outputs(1640));
    layer1_outputs(1416) <= not(layer0_outputs(632)) or (layer0_outputs(1481));
    layer1_outputs(1417) <= layer0_outputs(1039);
    layer1_outputs(1418) <= layer0_outputs(2133);
    layer1_outputs(1419) <= not((layer0_outputs(1193)) or (layer0_outputs(2260)));
    layer1_outputs(1420) <= '1';
    layer1_outputs(1421) <= '0';
    layer1_outputs(1422) <= '1';
    layer1_outputs(1423) <= not((layer0_outputs(2300)) and (layer0_outputs(1552)));
    layer1_outputs(1424) <= '1';
    layer1_outputs(1425) <= not((layer0_outputs(407)) and (layer0_outputs(1723)));
    layer1_outputs(1426) <= '1';
    layer1_outputs(1427) <= not(layer0_outputs(2154));
    layer1_outputs(1428) <= not(layer0_outputs(1640));
    layer1_outputs(1429) <= not(layer0_outputs(2)) or (layer0_outputs(1190));
    layer1_outputs(1430) <= '0';
    layer1_outputs(1431) <= not(layer0_outputs(395));
    layer1_outputs(1432) <= not(layer0_outputs(878)) or (layer0_outputs(1739));
    layer1_outputs(1433) <= not(layer0_outputs(416));
    layer1_outputs(1434) <= layer0_outputs(66);
    layer1_outputs(1435) <= (layer0_outputs(2126)) or (layer0_outputs(1402));
    layer1_outputs(1436) <= (layer0_outputs(2179)) and not (layer0_outputs(1280));
    layer1_outputs(1437) <= (layer0_outputs(2216)) and not (layer0_outputs(2001));
    layer1_outputs(1438) <= not(layer0_outputs(2201)) or (layer0_outputs(74));
    layer1_outputs(1439) <= not(layer0_outputs(1449)) or (layer0_outputs(1702));
    layer1_outputs(1440) <= not(layer0_outputs(1155)) or (layer0_outputs(1988));
    layer1_outputs(1441) <= not(layer0_outputs(31));
    layer1_outputs(1442) <= (layer0_outputs(2066)) and not (layer0_outputs(478));
    layer1_outputs(1443) <= not(layer0_outputs(2248));
    layer1_outputs(1444) <= layer0_outputs(774);
    layer1_outputs(1445) <= not(layer0_outputs(993));
    layer1_outputs(1446) <= '1';
    layer1_outputs(1447) <= not((layer0_outputs(1977)) or (layer0_outputs(989)));
    layer1_outputs(1448) <= layer0_outputs(316);
    layer1_outputs(1449) <= '1';
    layer1_outputs(1450) <= not(layer0_outputs(308)) or (layer0_outputs(684));
    layer1_outputs(1451) <= '1';
    layer1_outputs(1452) <= not(layer0_outputs(1044)) or (layer0_outputs(1244));
    layer1_outputs(1453) <= not(layer0_outputs(1123)) or (layer0_outputs(1485));
    layer1_outputs(1454) <= (layer0_outputs(247)) or (layer0_outputs(486));
    layer1_outputs(1455) <= (layer0_outputs(1389)) and not (layer0_outputs(1321));
    layer1_outputs(1456) <= (layer0_outputs(2273)) or (layer0_outputs(825));
    layer1_outputs(1457) <= not((layer0_outputs(527)) or (layer0_outputs(870)));
    layer1_outputs(1458) <= '1';
    layer1_outputs(1459) <= not(layer0_outputs(1459));
    layer1_outputs(1460) <= '1';
    layer1_outputs(1461) <= not(layer0_outputs(1803));
    layer1_outputs(1462) <= not((layer0_outputs(290)) and (layer0_outputs(765)));
    layer1_outputs(1463) <= '0';
    layer1_outputs(1464) <= '0';
    layer1_outputs(1465) <= '1';
    layer1_outputs(1466) <= layer0_outputs(2349);
    layer1_outputs(1467) <= '1';
    layer1_outputs(1468) <= layer0_outputs(81);
    layer1_outputs(1469) <= '1';
    layer1_outputs(1470) <= layer0_outputs(2175);
    layer1_outputs(1471) <= not((layer0_outputs(568)) and (layer0_outputs(1992)));
    layer1_outputs(1472) <= '1';
    layer1_outputs(1473) <= not(layer0_outputs(1633)) or (layer0_outputs(1779));
    layer1_outputs(1474) <= (layer0_outputs(1543)) and not (layer0_outputs(485));
    layer1_outputs(1475) <= layer0_outputs(1397);
    layer1_outputs(1476) <= not(layer0_outputs(2019)) or (layer0_outputs(973));
    layer1_outputs(1477) <= not((layer0_outputs(1935)) and (layer0_outputs(171)));
    layer1_outputs(1478) <= not(layer0_outputs(1754));
    layer1_outputs(1479) <= '0';
    layer1_outputs(1480) <= not((layer0_outputs(2147)) or (layer0_outputs(1606)));
    layer1_outputs(1481) <= not((layer0_outputs(808)) or (layer0_outputs(176)));
    layer1_outputs(1482) <= not((layer0_outputs(1217)) and (layer0_outputs(1180)));
    layer1_outputs(1483) <= not(layer0_outputs(1285));
    layer1_outputs(1484) <= layer0_outputs(402);
    layer1_outputs(1485) <= (layer0_outputs(958)) and not (layer0_outputs(2534));
    layer1_outputs(1486) <= not((layer0_outputs(1017)) and (layer0_outputs(313)));
    layer1_outputs(1487) <= (layer0_outputs(577)) and (layer0_outputs(331));
    layer1_outputs(1488) <= (layer0_outputs(1705)) and (layer0_outputs(2129));
    layer1_outputs(1489) <= not((layer0_outputs(2076)) and (layer0_outputs(1819)));
    layer1_outputs(1490) <= (layer0_outputs(802)) or (layer0_outputs(101));
    layer1_outputs(1491) <= layer0_outputs(1154);
    layer1_outputs(1492) <= not(layer0_outputs(2400)) or (layer0_outputs(335));
    layer1_outputs(1493) <= not(layer0_outputs(1584));
    layer1_outputs(1494) <= (layer0_outputs(2331)) or (layer0_outputs(1105));
    layer1_outputs(1495) <= not((layer0_outputs(2206)) or (layer0_outputs(75)));
    layer1_outputs(1496) <= not(layer0_outputs(2288));
    layer1_outputs(1497) <= not(layer0_outputs(161));
    layer1_outputs(1498) <= not(layer0_outputs(549)) or (layer0_outputs(2371));
    layer1_outputs(1499) <= (layer0_outputs(1339)) and not (layer0_outputs(187));
    layer1_outputs(1500) <= layer0_outputs(575);
    layer1_outputs(1501) <= (layer0_outputs(335)) and (layer0_outputs(2199));
    layer1_outputs(1502) <= (layer0_outputs(2451)) and (layer0_outputs(1823));
    layer1_outputs(1503) <= '1';
    layer1_outputs(1504) <= not((layer0_outputs(322)) and (layer0_outputs(931)));
    layer1_outputs(1505) <= not(layer0_outputs(1232)) or (layer0_outputs(367));
    layer1_outputs(1506) <= (layer0_outputs(1104)) and not (layer0_outputs(1972));
    layer1_outputs(1507) <= not((layer0_outputs(284)) and (layer0_outputs(183)));
    layer1_outputs(1508) <= (layer0_outputs(816)) and (layer0_outputs(248));
    layer1_outputs(1509) <= not(layer0_outputs(2366));
    layer1_outputs(1510) <= not(layer0_outputs(1710)) or (layer0_outputs(2329));
    layer1_outputs(1511) <= (layer0_outputs(399)) or (layer0_outputs(1953));
    layer1_outputs(1512) <= layer0_outputs(867);
    layer1_outputs(1513) <= not(layer0_outputs(1277)) or (layer0_outputs(293));
    layer1_outputs(1514) <= (layer0_outputs(1575)) and not (layer0_outputs(118));
    layer1_outputs(1515) <= (layer0_outputs(2368)) or (layer0_outputs(337));
    layer1_outputs(1516) <= (layer0_outputs(1260)) and not (layer0_outputs(1911));
    layer1_outputs(1517) <= '1';
    layer1_outputs(1518) <= '0';
    layer1_outputs(1519) <= layer0_outputs(2382);
    layer1_outputs(1520) <= layer0_outputs(477);
    layer1_outputs(1521) <= '1';
    layer1_outputs(1522) <= not((layer0_outputs(122)) and (layer0_outputs(224)));
    layer1_outputs(1523) <= not(layer0_outputs(2062)) or (layer0_outputs(2542));
    layer1_outputs(1524) <= '1';
    layer1_outputs(1525) <= '0';
    layer1_outputs(1526) <= (layer0_outputs(329)) and not (layer0_outputs(767));
    layer1_outputs(1527) <= '0';
    layer1_outputs(1528) <= not((layer0_outputs(1704)) and (layer0_outputs(2240)));
    layer1_outputs(1529) <= layer0_outputs(178);
    layer1_outputs(1530) <= layer0_outputs(818);
    layer1_outputs(1531) <= (layer0_outputs(2036)) and not (layer0_outputs(1151));
    layer1_outputs(1532) <= layer0_outputs(824);
    layer1_outputs(1533) <= (layer0_outputs(856)) or (layer0_outputs(1007));
    layer1_outputs(1534) <= not(layer0_outputs(1375)) or (layer0_outputs(1480));
    layer1_outputs(1535) <= not(layer0_outputs(1242));
    layer1_outputs(1536) <= layer0_outputs(865);
    layer1_outputs(1537) <= (layer0_outputs(1798)) and not (layer0_outputs(1669));
    layer1_outputs(1538) <= (layer0_outputs(1662)) and (layer0_outputs(720));
    layer1_outputs(1539) <= (layer0_outputs(603)) or (layer0_outputs(1894));
    layer1_outputs(1540) <= (layer0_outputs(107)) or (layer0_outputs(553));
    layer1_outputs(1541) <= layer0_outputs(904);
    layer1_outputs(1542) <= not(layer0_outputs(297)) or (layer0_outputs(651));
    layer1_outputs(1543) <= not(layer0_outputs(2233));
    layer1_outputs(1544) <= layer0_outputs(1526);
    layer1_outputs(1545) <= (layer0_outputs(1671)) and (layer0_outputs(1689));
    layer1_outputs(1546) <= (layer0_outputs(812)) or (layer0_outputs(97));
    layer1_outputs(1547) <= not(layer0_outputs(1358));
    layer1_outputs(1548) <= not((layer0_outputs(611)) and (layer0_outputs(2362)));
    layer1_outputs(1549) <= (layer0_outputs(2353)) and (layer0_outputs(1437));
    layer1_outputs(1550) <= not(layer0_outputs(84)) or (layer0_outputs(421));
    layer1_outputs(1551) <= layer0_outputs(370);
    layer1_outputs(1552) <= '1';
    layer1_outputs(1553) <= '1';
    layer1_outputs(1554) <= (layer0_outputs(1909)) and (layer0_outputs(729));
    layer1_outputs(1555) <= layer0_outputs(37);
    layer1_outputs(1556) <= not(layer0_outputs(2268));
    layer1_outputs(1557) <= not((layer0_outputs(175)) or (layer0_outputs(2467)));
    layer1_outputs(1558) <= layer0_outputs(1237);
    layer1_outputs(1559) <= layer0_outputs(683);
    layer1_outputs(1560) <= not(layer0_outputs(1793));
    layer1_outputs(1561) <= not(layer0_outputs(2239));
    layer1_outputs(1562) <= '1';
    layer1_outputs(1563) <= '0';
    layer1_outputs(1564) <= '1';
    layer1_outputs(1565) <= (layer0_outputs(2327)) and (layer0_outputs(1322));
    layer1_outputs(1566) <= (layer0_outputs(1161)) and not (layer0_outputs(1094));
    layer1_outputs(1567) <= '1';
    layer1_outputs(1568) <= (layer0_outputs(846)) and (layer0_outputs(740));
    layer1_outputs(1569) <= layer0_outputs(45);
    layer1_outputs(1570) <= '0';
    layer1_outputs(1571) <= layer0_outputs(7);
    layer1_outputs(1572) <= '0';
    layer1_outputs(1573) <= (layer0_outputs(1045)) or (layer0_outputs(2348));
    layer1_outputs(1574) <= not((layer0_outputs(1446)) or (layer0_outputs(2156)));
    layer1_outputs(1575) <= (layer0_outputs(971)) and not (layer0_outputs(1194));
    layer1_outputs(1576) <= not(layer0_outputs(320)) or (layer0_outputs(1365));
    layer1_outputs(1577) <= '1';
    layer1_outputs(1578) <= '0';
    layer1_outputs(1579) <= layer0_outputs(534);
    layer1_outputs(1580) <= not(layer0_outputs(849));
    layer1_outputs(1581) <= '1';
    layer1_outputs(1582) <= not(layer0_outputs(1682)) or (layer0_outputs(2093));
    layer1_outputs(1583) <= (layer0_outputs(1476)) or (layer0_outputs(1833));
    layer1_outputs(1584) <= not((layer0_outputs(955)) or (layer0_outputs(1713)));
    layer1_outputs(1585) <= (layer0_outputs(181)) and not (layer0_outputs(2288));
    layer1_outputs(1586) <= not((layer0_outputs(2403)) xor (layer0_outputs(2416)));
    layer1_outputs(1587) <= '1';
    layer1_outputs(1588) <= '1';
    layer1_outputs(1589) <= layer0_outputs(933);
    layer1_outputs(1590) <= not(layer0_outputs(1980));
    layer1_outputs(1591) <= layer0_outputs(1167);
    layer1_outputs(1592) <= (layer0_outputs(1529)) and (layer0_outputs(1126));
    layer1_outputs(1593) <= not((layer0_outputs(299)) or (layer0_outputs(792)));
    layer1_outputs(1594) <= not(layer0_outputs(1092));
    layer1_outputs(1595) <= layer0_outputs(1686);
    layer1_outputs(1596) <= '0';
    layer1_outputs(1597) <= layer0_outputs(1869);
    layer1_outputs(1598) <= layer0_outputs(115);
    layer1_outputs(1599) <= not(layer0_outputs(2292));
    layer1_outputs(1600) <= '1';
    layer1_outputs(1601) <= layer0_outputs(2263);
    layer1_outputs(1602) <= (layer0_outputs(1387)) and not (layer0_outputs(2222));
    layer1_outputs(1603) <= (layer0_outputs(14)) or (layer0_outputs(1677));
    layer1_outputs(1604) <= '0';
    layer1_outputs(1605) <= '0';
    layer1_outputs(1606) <= not(layer0_outputs(1714));
    layer1_outputs(1607) <= not(layer0_outputs(319));
    layer1_outputs(1608) <= not(layer0_outputs(1137));
    layer1_outputs(1609) <= (layer0_outputs(126)) and not (layer0_outputs(576));
    layer1_outputs(1610) <= layer0_outputs(2076);
    layer1_outputs(1611) <= not(layer0_outputs(945));
    layer1_outputs(1612) <= not(layer0_outputs(172));
    layer1_outputs(1613) <= (layer0_outputs(2550)) and not (layer0_outputs(2217));
    layer1_outputs(1614) <= layer0_outputs(2163);
    layer1_outputs(1615) <= not((layer0_outputs(2425)) and (layer0_outputs(1175)));
    layer1_outputs(1616) <= not(layer0_outputs(1571)) or (layer0_outputs(2265));
    layer1_outputs(1617) <= (layer0_outputs(246)) and not (layer0_outputs(411));
    layer1_outputs(1618) <= not(layer0_outputs(113)) or (layer0_outputs(1285));
    layer1_outputs(1619) <= not(layer0_outputs(742));
    layer1_outputs(1620) <= layer0_outputs(2189);
    layer1_outputs(1621) <= not((layer0_outputs(2203)) or (layer0_outputs(1576)));
    layer1_outputs(1622) <= (layer0_outputs(1245)) and (layer0_outputs(2427));
    layer1_outputs(1623) <= (layer0_outputs(991)) and not (layer0_outputs(1784));
    layer1_outputs(1624) <= layer0_outputs(539);
    layer1_outputs(1625) <= not(layer0_outputs(2323));
    layer1_outputs(1626) <= '0';
    layer1_outputs(1627) <= (layer0_outputs(408)) and not (layer0_outputs(2244));
    layer1_outputs(1628) <= (layer0_outputs(1328)) and not (layer0_outputs(283));
    layer1_outputs(1629) <= layer0_outputs(475);
    layer1_outputs(1630) <= not(layer0_outputs(2511));
    layer1_outputs(1631) <= '1';
    layer1_outputs(1632) <= '1';
    layer1_outputs(1633) <= '1';
    layer1_outputs(1634) <= '0';
    layer1_outputs(1635) <= (layer0_outputs(1709)) and (layer0_outputs(312));
    layer1_outputs(1636) <= (layer0_outputs(1281)) and (layer0_outputs(481));
    layer1_outputs(1637) <= (layer0_outputs(287)) and not (layer0_outputs(976));
    layer1_outputs(1638) <= not(layer0_outputs(33));
    layer1_outputs(1639) <= not(layer0_outputs(1752)) or (layer0_outputs(365));
    layer1_outputs(1640) <= (layer0_outputs(1904)) or (layer0_outputs(1332));
    layer1_outputs(1641) <= not(layer0_outputs(95)) or (layer0_outputs(1348));
    layer1_outputs(1642) <= (layer0_outputs(497)) and not (layer0_outputs(1215));
    layer1_outputs(1643) <= not((layer0_outputs(868)) or (layer0_outputs(700)));
    layer1_outputs(1644) <= (layer0_outputs(2386)) or (layer0_outputs(351));
    layer1_outputs(1645) <= not(layer0_outputs(12));
    layer1_outputs(1646) <= (layer0_outputs(535)) and not (layer0_outputs(571));
    layer1_outputs(1647) <= '0';
    layer1_outputs(1648) <= not((layer0_outputs(1088)) or (layer0_outputs(2436)));
    layer1_outputs(1649) <= not(layer0_outputs(1542));
    layer1_outputs(1650) <= layer0_outputs(921);
    layer1_outputs(1651) <= '0';
    layer1_outputs(1652) <= not((layer0_outputs(1304)) and (layer0_outputs(965)));
    layer1_outputs(1653) <= not((layer0_outputs(560)) or (layer0_outputs(882)));
    layer1_outputs(1654) <= (layer0_outputs(210)) and not (layer0_outputs(464));
    layer1_outputs(1655) <= not(layer0_outputs(689)) or (layer0_outputs(2242));
    layer1_outputs(1656) <= (layer0_outputs(2331)) and not (layer0_outputs(1902));
    layer1_outputs(1657) <= (layer0_outputs(1063)) and (layer0_outputs(1519));
    layer1_outputs(1658) <= not(layer0_outputs(1785));
    layer1_outputs(1659) <= '0';
    layer1_outputs(1660) <= (layer0_outputs(2198)) and not (layer0_outputs(842));
    layer1_outputs(1661) <= layer0_outputs(1207);
    layer1_outputs(1662) <= not(layer0_outputs(866)) or (layer0_outputs(2319));
    layer1_outputs(1663) <= not(layer0_outputs(1725)) or (layer0_outputs(423));
    layer1_outputs(1664) <= (layer0_outputs(1569)) and not (layer0_outputs(1273));
    layer1_outputs(1665) <= not(layer0_outputs(331)) or (layer0_outputs(1044));
    layer1_outputs(1666) <= layer0_outputs(2123);
    layer1_outputs(1667) <= not((layer0_outputs(1875)) and (layer0_outputs(34)));
    layer1_outputs(1668) <= '1';
    layer1_outputs(1669) <= not((layer0_outputs(1558)) and (layer0_outputs(942)));
    layer1_outputs(1670) <= not((layer0_outputs(119)) or (layer0_outputs(2470)));
    layer1_outputs(1671) <= '1';
    layer1_outputs(1672) <= layer0_outputs(257);
    layer1_outputs(1673) <= not((layer0_outputs(267)) or (layer0_outputs(315)));
    layer1_outputs(1674) <= (layer0_outputs(1286)) and not (layer0_outputs(1826));
    layer1_outputs(1675) <= not(layer0_outputs(1157)) or (layer0_outputs(1450));
    layer1_outputs(1676) <= (layer0_outputs(1267)) and not (layer0_outputs(1525));
    layer1_outputs(1677) <= (layer0_outputs(929)) and (layer0_outputs(1081));
    layer1_outputs(1678) <= (layer0_outputs(306)) and not (layer0_outputs(1177));
    layer1_outputs(1679) <= not(layer0_outputs(178));
    layer1_outputs(1680) <= '1';
    layer1_outputs(1681) <= not(layer0_outputs(197));
    layer1_outputs(1682) <= not(layer0_outputs(528));
    layer1_outputs(1683) <= (layer0_outputs(1058)) and not (layer0_outputs(1829));
    layer1_outputs(1684) <= (layer0_outputs(2505)) xor (layer0_outputs(1791));
    layer1_outputs(1685) <= '0';
    layer1_outputs(1686) <= (layer0_outputs(1539)) or (layer0_outputs(2069));
    layer1_outputs(1687) <= '0';
    layer1_outputs(1688) <= (layer0_outputs(2334)) xor (layer0_outputs(1536));
    layer1_outputs(1689) <= not((layer0_outputs(273)) and (layer0_outputs(87)));
    layer1_outputs(1690) <= '1';
    layer1_outputs(1691) <= '1';
    layer1_outputs(1692) <= not((layer0_outputs(2336)) xor (layer0_outputs(845)));
    layer1_outputs(1693) <= not(layer0_outputs(668)) or (layer0_outputs(1619));
    layer1_outputs(1694) <= layer0_outputs(259);
    layer1_outputs(1695) <= layer0_outputs(450);
    layer1_outputs(1696) <= layer0_outputs(1808);
    layer1_outputs(1697) <= '0';
    layer1_outputs(1698) <= '1';
    layer1_outputs(1699) <= '0';
    layer1_outputs(1700) <= '1';
    layer1_outputs(1701) <= not(layer0_outputs(1716)) or (layer0_outputs(1975));
    layer1_outputs(1702) <= (layer0_outputs(1535)) xor (layer0_outputs(114));
    layer1_outputs(1703) <= layer0_outputs(1247);
    layer1_outputs(1704) <= (layer0_outputs(1132)) and not (layer0_outputs(492));
    layer1_outputs(1705) <= '0';
    layer1_outputs(1706) <= not(layer0_outputs(466)) or (layer0_outputs(1380));
    layer1_outputs(1707) <= not(layer0_outputs(1541));
    layer1_outputs(1708) <= not((layer0_outputs(1451)) and (layer0_outputs(1319)));
    layer1_outputs(1709) <= '0';
    layer1_outputs(1710) <= not(layer0_outputs(756));
    layer1_outputs(1711) <= not((layer0_outputs(595)) or (layer0_outputs(2139)));
    layer1_outputs(1712) <= (layer0_outputs(2310)) and (layer0_outputs(400));
    layer1_outputs(1713) <= not(layer0_outputs(324));
    layer1_outputs(1714) <= layer0_outputs(1221);
    layer1_outputs(1715) <= not((layer0_outputs(2157)) and (layer0_outputs(605)));
    layer1_outputs(1716) <= not(layer0_outputs(161)) or (layer0_outputs(1416));
    layer1_outputs(1717) <= layer0_outputs(726);
    layer1_outputs(1718) <= (layer0_outputs(1269)) and not (layer0_outputs(2174));
    layer1_outputs(1719) <= '1';
    layer1_outputs(1720) <= not(layer0_outputs(60));
    layer1_outputs(1721) <= layer0_outputs(138);
    layer1_outputs(1722) <= not(layer0_outputs(600));
    layer1_outputs(1723) <= (layer0_outputs(300)) and (layer0_outputs(1434));
    layer1_outputs(1724) <= (layer0_outputs(1199)) or (layer0_outputs(1118));
    layer1_outputs(1725) <= not(layer0_outputs(1628));
    layer1_outputs(1726) <= (layer0_outputs(270)) and (layer0_outputs(1696));
    layer1_outputs(1727) <= layer0_outputs(1837);
    layer1_outputs(1728) <= not(layer0_outputs(847)) or (layer0_outputs(188));
    layer1_outputs(1729) <= not(layer0_outputs(551)) or (layer0_outputs(2016));
    layer1_outputs(1730) <= '1';
    layer1_outputs(1731) <= (layer0_outputs(2264)) and not (layer0_outputs(1506));
    layer1_outputs(1732) <= (layer0_outputs(918)) and (layer0_outputs(837));
    layer1_outputs(1733) <= layer0_outputs(972);
    layer1_outputs(1734) <= layer0_outputs(1231);
    layer1_outputs(1735) <= '0';
    layer1_outputs(1736) <= (layer0_outputs(1930)) and not (layer0_outputs(2125));
    layer1_outputs(1737) <= not(layer0_outputs(2005)) or (layer0_outputs(523));
    layer1_outputs(1738) <= layer0_outputs(42);
    layer1_outputs(1739) <= not(layer0_outputs(226)) or (layer0_outputs(1405));
    layer1_outputs(1740) <= (layer0_outputs(1195)) and not (layer0_outputs(971));
    layer1_outputs(1741) <= not(layer0_outputs(278));
    layer1_outputs(1742) <= not(layer0_outputs(1675));
    layer1_outputs(1743) <= (layer0_outputs(418)) and (layer0_outputs(1489));
    layer1_outputs(1744) <= not(layer0_outputs(2252));
    layer1_outputs(1745) <= layer0_outputs(1652);
    layer1_outputs(1746) <= layer0_outputs(1142);
    layer1_outputs(1747) <= not(layer0_outputs(1015)) or (layer0_outputs(1437));
    layer1_outputs(1748) <= layer0_outputs(1700);
    layer1_outputs(1749) <= layer0_outputs(111);
    layer1_outputs(1750) <= not(layer0_outputs(1656));
    layer1_outputs(1751) <= layer0_outputs(707);
    layer1_outputs(1752) <= not((layer0_outputs(2034)) or (layer0_outputs(656)));
    layer1_outputs(1753) <= '0';
    layer1_outputs(1754) <= not(layer0_outputs(920));
    layer1_outputs(1755) <= layer0_outputs(1361);
    layer1_outputs(1756) <= not((layer0_outputs(1338)) and (layer0_outputs(1224)));
    layer1_outputs(1757) <= layer0_outputs(2017);
    layer1_outputs(1758) <= not(layer0_outputs(389)) or (layer0_outputs(480));
    layer1_outputs(1759) <= not(layer0_outputs(1533)) or (layer0_outputs(78));
    layer1_outputs(1760) <= layer0_outputs(2559);
    layer1_outputs(1761) <= '1';
    layer1_outputs(1762) <= layer0_outputs(1942);
    layer1_outputs(1763) <= not(layer0_outputs(57)) or (layer0_outputs(2400));
    layer1_outputs(1764) <= '0';
    layer1_outputs(1765) <= (layer0_outputs(966)) and not (layer0_outputs(992));
    layer1_outputs(1766) <= not(layer0_outputs(2527)) or (layer0_outputs(67));
    layer1_outputs(1767) <= '1';
    layer1_outputs(1768) <= '0';
    layer1_outputs(1769) <= not(layer0_outputs(1226)) or (layer0_outputs(1150));
    layer1_outputs(1770) <= not(layer0_outputs(1785));
    layer1_outputs(1771) <= '1';
    layer1_outputs(1772) <= (layer0_outputs(124)) and (layer0_outputs(264));
    layer1_outputs(1773) <= layer0_outputs(206);
    layer1_outputs(1774) <= '0';
    layer1_outputs(1775) <= not((layer0_outputs(1941)) and (layer0_outputs(604)));
    layer1_outputs(1776) <= '1';
    layer1_outputs(1777) <= '1';
    layer1_outputs(1778) <= '1';
    layer1_outputs(1779) <= '1';
    layer1_outputs(1780) <= layer0_outputs(858);
    layer1_outputs(1781) <= not(layer0_outputs(1012)) or (layer0_outputs(1211));
    layer1_outputs(1782) <= '1';
    layer1_outputs(1783) <= not(layer0_outputs(351));
    layer1_outputs(1784) <= (layer0_outputs(2270)) or (layer0_outputs(1799));
    layer1_outputs(1785) <= (layer0_outputs(643)) or (layer0_outputs(430));
    layer1_outputs(1786) <= '0';
    layer1_outputs(1787) <= not((layer0_outputs(1502)) and (layer0_outputs(1871)));
    layer1_outputs(1788) <= layer0_outputs(118);
    layer1_outputs(1789) <= not((layer0_outputs(68)) or (layer0_outputs(424)));
    layer1_outputs(1790) <= (layer0_outputs(2385)) or (layer0_outputs(51));
    layer1_outputs(1791) <= not(layer0_outputs(471));
    layer1_outputs(1792) <= '1';
    layer1_outputs(1793) <= not((layer0_outputs(1144)) or (layer0_outputs(1230)));
    layer1_outputs(1794) <= layer0_outputs(2239);
    layer1_outputs(1795) <= not(layer0_outputs(1125)) or (layer0_outputs(1644));
    layer1_outputs(1796) <= not(layer0_outputs(958)) or (layer0_outputs(1072));
    layer1_outputs(1797) <= '1';
    layer1_outputs(1798) <= layer0_outputs(2055);
    layer1_outputs(1799) <= not((layer0_outputs(2106)) and (layer0_outputs(299)));
    layer1_outputs(1800) <= layer0_outputs(1223);
    layer1_outputs(1801) <= (layer0_outputs(260)) xor (layer0_outputs(562));
    layer1_outputs(1802) <= layer0_outputs(1592);
    layer1_outputs(1803) <= (layer0_outputs(1071)) and not (layer0_outputs(1957));
    layer1_outputs(1804) <= (layer0_outputs(2449)) and not (layer0_outputs(324));
    layer1_outputs(1805) <= not((layer0_outputs(1990)) or (layer0_outputs(401)));
    layer1_outputs(1806) <= not(layer0_outputs(1612));
    layer1_outputs(1807) <= '0';
    layer1_outputs(1808) <= (layer0_outputs(2397)) and not (layer0_outputs(114));
    layer1_outputs(1809) <= layer0_outputs(1294);
    layer1_outputs(1810) <= not((layer0_outputs(2205)) or (layer0_outputs(246)));
    layer1_outputs(1811) <= (layer0_outputs(702)) and not (layer0_outputs(35));
    layer1_outputs(1812) <= not(layer0_outputs(1936)) or (layer0_outputs(1293));
    layer1_outputs(1813) <= layer0_outputs(1778);
    layer1_outputs(1814) <= not(layer0_outputs(1815));
    layer1_outputs(1815) <= '1';
    layer1_outputs(1816) <= not(layer0_outputs(1429));
    layer1_outputs(1817) <= '0';
    layer1_outputs(1818) <= layer0_outputs(2277);
    layer1_outputs(1819) <= not((layer0_outputs(759)) or (layer0_outputs(646)));
    layer1_outputs(1820) <= not((layer0_outputs(940)) and (layer0_outputs(1739)));
    layer1_outputs(1821) <= (layer0_outputs(344)) and (layer0_outputs(842));
    layer1_outputs(1822) <= '0';
    layer1_outputs(1823) <= (layer0_outputs(2057)) and not (layer0_outputs(132));
    layer1_outputs(1824) <= '1';
    layer1_outputs(1825) <= layer0_outputs(2370);
    layer1_outputs(1826) <= not((layer0_outputs(2228)) or (layer0_outputs(2390)));
    layer1_outputs(1827) <= not((layer0_outputs(1923)) or (layer0_outputs(901)));
    layer1_outputs(1828) <= layer0_outputs(2281);
    layer1_outputs(1829) <= layer0_outputs(984);
    layer1_outputs(1830) <= (layer0_outputs(1809)) and (layer0_outputs(1336));
    layer1_outputs(1831) <= not((layer0_outputs(2428)) xor (layer0_outputs(917)));
    layer1_outputs(1832) <= not((layer0_outputs(1861)) or (layer0_outputs(1046)));
    layer1_outputs(1833) <= layer0_outputs(143);
    layer1_outputs(1834) <= not(layer0_outputs(1846));
    layer1_outputs(1835) <= not((layer0_outputs(1553)) or (layer0_outputs(1477)));
    layer1_outputs(1836) <= '1';
    layer1_outputs(1837) <= layer0_outputs(2105);
    layer1_outputs(1838) <= not(layer0_outputs(2093)) or (layer0_outputs(849));
    layer1_outputs(1839) <= not(layer0_outputs(572)) or (layer0_outputs(1504));
    layer1_outputs(1840) <= (layer0_outputs(314)) and (layer0_outputs(1031));
    layer1_outputs(1841) <= not(layer0_outputs(526));
    layer1_outputs(1842) <= not(layer0_outputs(483));
    layer1_outputs(1843) <= (layer0_outputs(2467)) or (layer0_outputs(2535));
    layer1_outputs(1844) <= (layer0_outputs(1206)) and (layer0_outputs(541));
    layer1_outputs(1845) <= not(layer0_outputs(2466));
    layer1_outputs(1846) <= not(layer0_outputs(546));
    layer1_outputs(1847) <= (layer0_outputs(2192)) and (layer0_outputs(60));
    layer1_outputs(1848) <= (layer0_outputs(2305)) and not (layer0_outputs(1738));
    layer1_outputs(1849) <= '1';
    layer1_outputs(1850) <= not(layer0_outputs(135));
    layer1_outputs(1851) <= not((layer0_outputs(730)) and (layer0_outputs(908)));
    layer1_outputs(1852) <= not(layer0_outputs(1347));
    layer1_outputs(1853) <= not(layer0_outputs(2326));
    layer1_outputs(1854) <= layer0_outputs(384);
    layer1_outputs(1855) <= not(layer0_outputs(2559));
    layer1_outputs(1856) <= '1';
    layer1_outputs(1857) <= '0';
    layer1_outputs(1858) <= not(layer0_outputs(2145)) or (layer0_outputs(1317));
    layer1_outputs(1859) <= '0';
    layer1_outputs(1860) <= not((layer0_outputs(2168)) and (layer0_outputs(119)));
    layer1_outputs(1861) <= layer0_outputs(1937);
    layer1_outputs(1862) <= not((layer0_outputs(79)) and (layer0_outputs(2491)));
    layer1_outputs(1863) <= (layer0_outputs(417)) or (layer0_outputs(751));
    layer1_outputs(1864) <= (layer0_outputs(2088)) and not (layer0_outputs(1891));
    layer1_outputs(1865) <= not((layer0_outputs(980)) or (layer0_outputs(5)));
    layer1_outputs(1866) <= not(layer0_outputs(720));
    layer1_outputs(1867) <= '0';
    layer1_outputs(1868) <= layer0_outputs(2542);
    layer1_outputs(1869) <= (layer0_outputs(1753)) and not (layer0_outputs(933));
    layer1_outputs(1870) <= layer0_outputs(151);
    layer1_outputs(1871) <= '1';
    layer1_outputs(1872) <= not((layer0_outputs(953)) or (layer0_outputs(200)));
    layer1_outputs(1873) <= '1';
    layer1_outputs(1874) <= (layer0_outputs(1822)) or (layer0_outputs(254));
    layer1_outputs(1875) <= not((layer0_outputs(1515)) and (layer0_outputs(2115)));
    layer1_outputs(1876) <= layer0_outputs(1229);
    layer1_outputs(1877) <= not(layer0_outputs(1668));
    layer1_outputs(1878) <= layer0_outputs(197);
    layer1_outputs(1879) <= not(layer0_outputs(317)) or (layer0_outputs(619));
    layer1_outputs(1880) <= layer0_outputs(323);
    layer1_outputs(1881) <= (layer0_outputs(69)) and not (layer0_outputs(1037));
    layer1_outputs(1882) <= (layer0_outputs(572)) and not (layer0_outputs(2097));
    layer1_outputs(1883) <= not((layer0_outputs(323)) and (layer0_outputs(327)));
    layer1_outputs(1884) <= (layer0_outputs(1638)) and not (layer0_outputs(1322));
    layer1_outputs(1885) <= not(layer0_outputs(1332));
    layer1_outputs(1886) <= layer0_outputs(2357);
    layer1_outputs(1887) <= (layer0_outputs(2125)) and not (layer0_outputs(1025));
    layer1_outputs(1888) <= not((layer0_outputs(1940)) or (layer0_outputs(2054)));
    layer1_outputs(1889) <= '0';
    layer1_outputs(1890) <= not((layer0_outputs(1197)) or (layer0_outputs(1659)));
    layer1_outputs(1891) <= (layer0_outputs(2465)) or (layer0_outputs(1464));
    layer1_outputs(1892) <= layer0_outputs(1433);
    layer1_outputs(1893) <= layer0_outputs(261);
    layer1_outputs(1894) <= '0';
    layer1_outputs(1895) <= '1';
    layer1_outputs(1896) <= not(layer0_outputs(2558)) or (layer0_outputs(1435));
    layer1_outputs(1897) <= not(layer0_outputs(2246)) or (layer0_outputs(2492));
    layer1_outputs(1898) <= (layer0_outputs(2219)) and not (layer0_outputs(1727));
    layer1_outputs(1899) <= (layer0_outputs(685)) xor (layer0_outputs(2463));
    layer1_outputs(1900) <= '1';
    layer1_outputs(1901) <= (layer0_outputs(693)) or (layer0_outputs(1170));
    layer1_outputs(1902) <= '1';
    layer1_outputs(1903) <= (layer0_outputs(1794)) xor (layer0_outputs(169));
    layer1_outputs(1904) <= '1';
    layer1_outputs(1905) <= not((layer0_outputs(2432)) or (layer0_outputs(1279)));
    layer1_outputs(1906) <= '1';
    layer1_outputs(1907) <= not((layer0_outputs(1999)) or (layer0_outputs(1436)));
    layer1_outputs(1908) <= not(layer0_outputs(687));
    layer1_outputs(1909) <= layer0_outputs(1971);
    layer1_outputs(1910) <= not(layer0_outputs(791)) or (layer0_outputs(1812));
    layer1_outputs(1911) <= layer0_outputs(836);
    layer1_outputs(1912) <= not((layer0_outputs(439)) or (layer0_outputs(1646)));
    layer1_outputs(1913) <= (layer0_outputs(353)) and not (layer0_outputs(2368));
    layer1_outputs(1914) <= not(layer0_outputs(2181));
    layer1_outputs(1915) <= (layer0_outputs(2225)) and (layer0_outputs(1590));
    layer1_outputs(1916) <= '1';
    layer1_outputs(1917) <= (layer0_outputs(1860)) xor (layer0_outputs(193));
    layer1_outputs(1918) <= '1';
    layer1_outputs(1919) <= '0';
    layer1_outputs(1920) <= layer0_outputs(1708);
    layer1_outputs(1921) <= layer0_outputs(2297);
    layer1_outputs(1922) <= '1';
    layer1_outputs(1923) <= '1';
    layer1_outputs(1924) <= not((layer0_outputs(1734)) or (layer0_outputs(2120)));
    layer1_outputs(1925) <= (layer0_outputs(428)) and not (layer0_outputs(1335));
    layer1_outputs(1926) <= (layer0_outputs(585)) and not (layer0_outputs(1280));
    layer1_outputs(1927) <= (layer0_outputs(517)) and not (layer0_outputs(1682));
    layer1_outputs(1928) <= not((layer0_outputs(1694)) or (layer0_outputs(997)));
    layer1_outputs(1929) <= (layer0_outputs(2290)) and not (layer0_outputs(886));
    layer1_outputs(1930) <= '1';
    layer1_outputs(1931) <= '0';
    layer1_outputs(1932) <= (layer0_outputs(457)) and not (layer0_outputs(2188));
    layer1_outputs(1933) <= '0';
    layer1_outputs(1934) <= not(layer0_outputs(380)) or (layer0_outputs(944));
    layer1_outputs(1935) <= not((layer0_outputs(349)) or (layer0_outputs(149)));
    layer1_outputs(1936) <= not(layer0_outputs(41)) or (layer0_outputs(601));
    layer1_outputs(1937) <= layer0_outputs(1440);
    layer1_outputs(1938) <= not(layer0_outputs(853));
    layer1_outputs(1939) <= not(layer0_outputs(884)) or (layer0_outputs(2101));
    layer1_outputs(1940) <= (layer0_outputs(2176)) and not (layer0_outputs(1681));
    layer1_outputs(1941) <= '1';
    layer1_outputs(1942) <= '0';
    layer1_outputs(1943) <= not((layer0_outputs(1455)) and (layer0_outputs(828)));
    layer1_outputs(1944) <= not(layer0_outputs(1219));
    layer1_outputs(1945) <= (layer0_outputs(1796)) and not (layer0_outputs(287));
    layer1_outputs(1946) <= layer0_outputs(741);
    layer1_outputs(1947) <= (layer0_outputs(32)) and (layer0_outputs(141));
    layer1_outputs(1948) <= (layer0_outputs(1419)) or (layer0_outputs(1237));
    layer1_outputs(1949) <= not((layer0_outputs(520)) or (layer0_outputs(795)));
    layer1_outputs(1950) <= '0';
    layer1_outputs(1951) <= '0';
    layer1_outputs(1952) <= layer0_outputs(1657);
    layer1_outputs(1953) <= layer0_outputs(63);
    layer1_outputs(1954) <= not(layer0_outputs(1052));
    layer1_outputs(1955) <= not(layer0_outputs(2208)) or (layer0_outputs(1158));
    layer1_outputs(1956) <= not(layer0_outputs(1638));
    layer1_outputs(1957) <= layer0_outputs(2151);
    layer1_outputs(1958) <= not((layer0_outputs(318)) and (layer0_outputs(1107)));
    layer1_outputs(1959) <= '1';
    layer1_outputs(1960) <= layer0_outputs(2056);
    layer1_outputs(1961) <= (layer0_outputs(1323)) and not (layer0_outputs(244));
    layer1_outputs(1962) <= not(layer0_outputs(2337)) or (layer0_outputs(1246));
    layer1_outputs(1963) <= '0';
    layer1_outputs(1964) <= not(layer0_outputs(163)) or (layer0_outputs(691));
    layer1_outputs(1965) <= not(layer0_outputs(891)) or (layer0_outputs(1699));
    layer1_outputs(1966) <= layer0_outputs(16);
    layer1_outputs(1967) <= '1';
    layer1_outputs(1968) <= not(layer0_outputs(1860));
    layer1_outputs(1969) <= '0';
    layer1_outputs(1970) <= not(layer0_outputs(2141));
    layer1_outputs(1971) <= layer0_outputs(329);
    layer1_outputs(1972) <= (layer0_outputs(1325)) and (layer0_outputs(1719));
    layer1_outputs(1973) <= not(layer0_outputs(1554));
    layer1_outputs(1974) <= not((layer0_outputs(660)) or (layer0_outputs(1413)));
    layer1_outputs(1975) <= (layer0_outputs(1216)) and not (layer0_outputs(587));
    layer1_outputs(1976) <= '0';
    layer1_outputs(1977) <= not((layer0_outputs(1)) and (layer0_outputs(333)));
    layer1_outputs(1978) <= not(layer0_outputs(2045)) or (layer0_outputs(2022));
    layer1_outputs(1979) <= '0';
    layer1_outputs(1980) <= (layer0_outputs(1334)) and not (layer0_outputs(823));
    layer1_outputs(1981) <= '1';
    layer1_outputs(1982) <= '0';
    layer1_outputs(1983) <= '0';
    layer1_outputs(1984) <= not(layer0_outputs(1124)) or (layer0_outputs(2245));
    layer1_outputs(1985) <= (layer0_outputs(2536)) and not (layer0_outputs(2551));
    layer1_outputs(1986) <= (layer0_outputs(874)) and not (layer0_outputs(1100));
    layer1_outputs(1987) <= '1';
    layer1_outputs(1988) <= not((layer0_outputs(71)) or (layer0_outputs(946)));
    layer1_outputs(1989) <= (layer0_outputs(131)) and not (layer0_outputs(491));
    layer1_outputs(1990) <= not((layer0_outputs(639)) or (layer0_outputs(1440)));
    layer1_outputs(1991) <= not(layer0_outputs(2406)) or (layer0_outputs(2183));
    layer1_outputs(1992) <= layer0_outputs(370);
    layer1_outputs(1993) <= (layer0_outputs(1414)) or (layer0_outputs(1622));
    layer1_outputs(1994) <= not(layer0_outputs(2514)) or (layer0_outputs(420));
    layer1_outputs(1995) <= not(layer0_outputs(2060)) or (layer0_outputs(1676));
    layer1_outputs(1996) <= '1';
    layer1_outputs(1997) <= not((layer0_outputs(650)) or (layer0_outputs(498)));
    layer1_outputs(1998) <= not(layer0_outputs(1102)) or (layer0_outputs(164));
    layer1_outputs(1999) <= '1';
    layer1_outputs(2000) <= '1';
    layer1_outputs(2001) <= not(layer0_outputs(1468));
    layer1_outputs(2002) <= not(layer0_outputs(2150)) or (layer0_outputs(309));
    layer1_outputs(2003) <= layer0_outputs(2124);
    layer1_outputs(2004) <= not(layer0_outputs(1655));
    layer1_outputs(2005) <= not(layer0_outputs(1636));
    layer1_outputs(2006) <= not(layer0_outputs(1761));
    layer1_outputs(2007) <= '1';
    layer1_outputs(2008) <= not(layer0_outputs(1959)) or (layer0_outputs(54));
    layer1_outputs(2009) <= layer0_outputs(428);
    layer1_outputs(2010) <= (layer0_outputs(597)) or (layer0_outputs(1711));
    layer1_outputs(2011) <= not(layer0_outputs(1120));
    layer1_outputs(2012) <= not((layer0_outputs(250)) and (layer0_outputs(451)));
    layer1_outputs(2013) <= not(layer0_outputs(665)) or (layer0_outputs(1470));
    layer1_outputs(2014) <= not((layer0_outputs(1563)) or (layer0_outputs(1581)));
    layer1_outputs(2015) <= (layer0_outputs(1679)) and not (layer0_outputs(983));
    layer1_outputs(2016) <= '0';
    layer1_outputs(2017) <= not((layer0_outputs(195)) and (layer0_outputs(1028)));
    layer1_outputs(2018) <= (layer0_outputs(1944)) and not (layer0_outputs(265));
    layer1_outputs(2019) <= not(layer0_outputs(544)) or (layer0_outputs(145));
    layer1_outputs(2020) <= (layer0_outputs(2071)) and not (layer0_outputs(1961));
    layer1_outputs(2021) <= not(layer0_outputs(1693));
    layer1_outputs(2022) <= not((layer0_outputs(1307)) xor (layer0_outputs(683)));
    layer1_outputs(2023) <= '0';
    layer1_outputs(2024) <= (layer0_outputs(1189)) and (layer0_outputs(1561));
    layer1_outputs(2025) <= layer0_outputs(1448);
    layer1_outputs(2026) <= '0';
    layer1_outputs(2027) <= '1';
    layer1_outputs(2028) <= not(layer0_outputs(1206)) or (layer0_outputs(275));
    layer1_outputs(2029) <= not(layer0_outputs(65));
    layer1_outputs(2030) <= not((layer0_outputs(1333)) or (layer0_outputs(90)));
    layer1_outputs(2031) <= (layer0_outputs(1577)) and not (layer0_outputs(1096));
    layer1_outputs(2032) <= layer0_outputs(2051);
    layer1_outputs(2033) <= not(layer0_outputs(929)) or (layer0_outputs(1114));
    layer1_outputs(2034) <= not((layer0_outputs(706)) and (layer0_outputs(1819)));
    layer1_outputs(2035) <= layer0_outputs(2110);
    layer1_outputs(2036) <= not(layer0_outputs(515)) or (layer0_outputs(2107));
    layer1_outputs(2037) <= '0';
    layer1_outputs(2038) <= not(layer0_outputs(1118)) or (layer0_outputs(2520));
    layer1_outputs(2039) <= not(layer0_outputs(68));
    layer1_outputs(2040) <= (layer0_outputs(387)) and not (layer0_outputs(2457));
    layer1_outputs(2041) <= not(layer0_outputs(2113)) or (layer0_outputs(1931));
    layer1_outputs(2042) <= (layer0_outputs(661)) and (layer0_outputs(402));
    layer1_outputs(2043) <= layer0_outputs(43);
    layer1_outputs(2044) <= not(layer0_outputs(939)) or (layer0_outputs(234));
    layer1_outputs(2045) <= '0';
    layer1_outputs(2046) <= not(layer0_outputs(1173)) or (layer0_outputs(2017));
    layer1_outputs(2047) <= not(layer0_outputs(1664)) or (layer0_outputs(380));
    layer1_outputs(2048) <= (layer0_outputs(1839)) and not (layer0_outputs(2464));
    layer1_outputs(2049) <= not(layer0_outputs(1923));
    layer1_outputs(2050) <= '1';
    layer1_outputs(2051) <= (layer0_outputs(1272)) and not (layer0_outputs(818));
    layer1_outputs(2052) <= not((layer0_outputs(949)) and (layer0_outputs(593)));
    layer1_outputs(2053) <= (layer0_outputs(980)) or (layer0_outputs(2240));
    layer1_outputs(2054) <= (layer0_outputs(2025)) or (layer0_outputs(754));
    layer1_outputs(2055) <= '1';
    layer1_outputs(2056) <= layer0_outputs(1633);
    layer1_outputs(2057) <= (layer0_outputs(775)) or (layer0_outputs(165));
    layer1_outputs(2058) <= (layer0_outputs(2226)) or (layer0_outputs(2023));
    layer1_outputs(2059) <= '0';
    layer1_outputs(2060) <= not((layer0_outputs(2111)) or (layer0_outputs(1042)));
    layer1_outputs(2061) <= not(layer0_outputs(1595)) or (layer0_outputs(2012));
    layer1_outputs(2062) <= (layer0_outputs(1810)) and not (layer0_outputs(2484));
    layer1_outputs(2063) <= not(layer0_outputs(680)) or (layer0_outputs(2193));
    layer1_outputs(2064) <= '0';
    layer1_outputs(2065) <= not((layer0_outputs(1505)) or (layer0_outputs(2472)));
    layer1_outputs(2066) <= layer0_outputs(253);
    layer1_outputs(2067) <= not((layer0_outputs(167)) and (layer0_outputs(209)));
    layer1_outputs(2068) <= layer0_outputs(108);
    layer1_outputs(2069) <= layer0_outputs(1667);
    layer1_outputs(2070) <= not((layer0_outputs(83)) or (layer0_outputs(732)));
    layer1_outputs(2071) <= '0';
    layer1_outputs(2072) <= not((layer0_outputs(2026)) and (layer0_outputs(459)));
    layer1_outputs(2073) <= not(layer0_outputs(401));
    layer1_outputs(2074) <= (layer0_outputs(2146)) or (layer0_outputs(1501));
    layer1_outputs(2075) <= layer0_outputs(529);
    layer1_outputs(2076) <= '0';
    layer1_outputs(2077) <= (layer0_outputs(1678)) and (layer0_outputs(400));
    layer1_outputs(2078) <= '0';
    layer1_outputs(2079) <= '0';
    layer1_outputs(2080) <= '1';
    layer1_outputs(2081) <= (layer0_outputs(1562)) and (layer0_outputs(1680));
    layer1_outputs(2082) <= layer0_outputs(154);
    layer1_outputs(2083) <= layer0_outputs(125);
    layer1_outputs(2084) <= '1';
    layer1_outputs(2085) <= not(layer0_outputs(1707));
    layer1_outputs(2086) <= (layer0_outputs(2118)) and not (layer0_outputs(2153));
    layer1_outputs(2087) <= not(layer0_outputs(347));
    layer1_outputs(2088) <= layer0_outputs(172);
    layer1_outputs(2089) <= not((layer0_outputs(208)) or (layer0_outputs(600)));
    layer1_outputs(2090) <= '0';
    layer1_outputs(2091) <= not(layer0_outputs(301));
    layer1_outputs(2092) <= (layer0_outputs(1412)) and not (layer0_outputs(988));
    layer1_outputs(2093) <= (layer0_outputs(2221)) and (layer0_outputs(1122));
    layer1_outputs(2094) <= '1';
    layer1_outputs(2095) <= not(layer0_outputs(1882));
    layer1_outputs(2096) <= layer0_outputs(408);
    layer1_outputs(2097) <= (layer0_outputs(2370)) and not (layer0_outputs(1832));
    layer1_outputs(2098) <= (layer0_outputs(1427)) and (layer0_outputs(1708));
    layer1_outputs(2099) <= not(layer0_outputs(1049));
    layer1_outputs(2100) <= not((layer0_outputs(1968)) or (layer0_outputs(1090)));
    layer1_outputs(2101) <= (layer0_outputs(1905)) or (layer0_outputs(2284));
    layer1_outputs(2102) <= '0';
    layer1_outputs(2103) <= (layer0_outputs(1815)) and not (layer0_outputs(1097));
    layer1_outputs(2104) <= (layer0_outputs(922)) and (layer0_outputs(2509));
    layer1_outputs(2105) <= '1';
    layer1_outputs(2106) <= (layer0_outputs(202)) and (layer0_outputs(694));
    layer1_outputs(2107) <= (layer0_outputs(2053)) xor (layer0_outputs(1674));
    layer1_outputs(2108) <= not(layer0_outputs(1036));
    layer1_outputs(2109) <= '1';
    layer1_outputs(2110) <= not(layer0_outputs(1765)) or (layer0_outputs(2458));
    layer1_outputs(2111) <= not(layer0_outputs(1652));
    layer1_outputs(2112) <= layer0_outputs(434);
    layer1_outputs(2113) <= not(layer0_outputs(1771)) or (layer0_outputs(198));
    layer1_outputs(2114) <= (layer0_outputs(592)) and not (layer0_outputs(669));
    layer1_outputs(2115) <= not(layer0_outputs(2235));
    layer1_outputs(2116) <= (layer0_outputs(1870)) and not (layer0_outputs(1419));
    layer1_outputs(2117) <= not(layer0_outputs(222));
    layer1_outputs(2118) <= not(layer0_outputs(393));
    layer1_outputs(2119) <= layer0_outputs(1271);
    layer1_outputs(2120) <= not(layer0_outputs(1493)) or (layer0_outputs(964));
    layer1_outputs(2121) <= not(layer0_outputs(1672));
    layer1_outputs(2122) <= '0';
    layer1_outputs(2123) <= not(layer0_outputs(763)) or (layer0_outputs(33));
    layer1_outputs(2124) <= not(layer0_outputs(1203));
    layer1_outputs(2125) <= not(layer0_outputs(2487));
    layer1_outputs(2126) <= '0';
    layer1_outputs(2127) <= layer0_outputs(1448);
    layer1_outputs(2128) <= not(layer0_outputs(650));
    layer1_outputs(2129) <= (layer0_outputs(759)) and not (layer0_outputs(352));
    layer1_outputs(2130) <= layer0_outputs(1569);
    layer1_outputs(2131) <= '0';
    layer1_outputs(2132) <= not(layer0_outputs(1466)) or (layer0_outputs(2196));
    layer1_outputs(2133) <= not(layer0_outputs(2141)) or (layer0_outputs(1248));
    layer1_outputs(2134) <= layer0_outputs(2335);
    layer1_outputs(2135) <= not(layer0_outputs(784));
    layer1_outputs(2136) <= '0';
    layer1_outputs(2137) <= layer0_outputs(537);
    layer1_outputs(2138) <= not(layer0_outputs(613)) or (layer0_outputs(367));
    layer1_outputs(2139) <= '0';
    layer1_outputs(2140) <= layer0_outputs(1955);
    layer1_outputs(2141) <= layer0_outputs(346);
    layer1_outputs(2142) <= '0';
    layer1_outputs(2143) <= (layer0_outputs(2100)) and not (layer0_outputs(2116));
    layer1_outputs(2144) <= not(layer0_outputs(2447)) or (layer0_outputs(2155));
    layer1_outputs(2145) <= layer0_outputs(2268);
    layer1_outputs(2146) <= (layer0_outputs(512)) and not (layer0_outputs(1256));
    layer1_outputs(2147) <= (layer0_outputs(1323)) or (layer0_outputs(128));
    layer1_outputs(2148) <= '1';
    layer1_outputs(2149) <= not(layer0_outputs(1070)) or (layer0_outputs(343));
    layer1_outputs(2150) <= '0';
    layer1_outputs(2151) <= not((layer0_outputs(271)) or (layer0_outputs(2393)));
    layer1_outputs(2152) <= (layer0_outputs(1107)) and not (layer0_outputs(705));
    layer1_outputs(2153) <= not(layer0_outputs(2000)) or (layer0_outputs(211));
    layer1_outputs(2154) <= not(layer0_outputs(2366)) or (layer0_outputs(1064));
    layer1_outputs(2155) <= not(layer0_outputs(1291)) or (layer0_outputs(423));
    layer1_outputs(2156) <= layer0_outputs(452);
    layer1_outputs(2157) <= not((layer0_outputs(924)) and (layer0_outputs(2038)));
    layer1_outputs(2158) <= '1';
    layer1_outputs(2159) <= (layer0_outputs(543)) and (layer0_outputs(2378));
    layer1_outputs(2160) <= layer0_outputs(2405);
    layer1_outputs(2161) <= not((layer0_outputs(1890)) and (layer0_outputs(1526)));
    layer1_outputs(2162) <= layer0_outputs(960);
    layer1_outputs(2163) <= (layer0_outputs(456)) or (layer0_outputs(1460));
    layer1_outputs(2164) <= layer0_outputs(24);
    layer1_outputs(2165) <= not(layer0_outputs(1747));
    layer1_outputs(2166) <= not(layer0_outputs(2500));
    layer1_outputs(2167) <= '1';
    layer1_outputs(2168) <= not(layer0_outputs(443));
    layer1_outputs(2169) <= '0';
    layer1_outputs(2170) <= not((layer0_outputs(1343)) and (layer0_outputs(1187)));
    layer1_outputs(2171) <= layer0_outputs(1003);
    layer1_outputs(2172) <= '0';
    layer1_outputs(2173) <= not(layer0_outputs(513)) or (layer0_outputs(2266));
    layer1_outputs(2174) <= not(layer0_outputs(2493));
    layer1_outputs(2175) <= not((layer0_outputs(2224)) or (layer0_outputs(1731)));
    layer1_outputs(2176) <= (layer0_outputs(887)) and (layer0_outputs(2446));
    layer1_outputs(2177) <= '0';
    layer1_outputs(2178) <= not(layer0_outputs(2544));
    layer1_outputs(2179) <= layer0_outputs(2132);
    layer1_outputs(2180) <= layer0_outputs(281);
    layer1_outputs(2181) <= not(layer0_outputs(307));
    layer1_outputs(2182) <= not((layer0_outputs(497)) or (layer0_outputs(460)));
    layer1_outputs(2183) <= not((layer0_outputs(382)) or (layer0_outputs(1836)));
    layer1_outputs(2184) <= (layer0_outputs(2495)) or (layer0_outputs(761));
    layer1_outputs(2185) <= not((layer0_outputs(981)) or (layer0_outputs(430)));
    layer1_outputs(2186) <= (layer0_outputs(1178)) and not (layer0_outputs(92));
    layer1_outputs(2187) <= not((layer0_outputs(1116)) and (layer0_outputs(2528)));
    layer1_outputs(2188) <= layer0_outputs(167);
    layer1_outputs(2189) <= '0';
    layer1_outputs(2190) <= '0';
    layer1_outputs(2191) <= not(layer0_outputs(1391));
    layer1_outputs(2192) <= layer0_outputs(1439);
    layer1_outputs(2193) <= (layer0_outputs(41)) and not (layer0_outputs(2010));
    layer1_outputs(2194) <= not((layer0_outputs(1749)) and (layer0_outputs(2293)));
    layer1_outputs(2195) <= layer0_outputs(1816);
    layer1_outputs(2196) <= not((layer0_outputs(602)) and (layer0_outputs(1814)));
    layer1_outputs(2197) <= layer0_outputs(1792);
    layer1_outputs(2198) <= (layer0_outputs(1303)) and not (layer0_outputs(451));
    layer1_outputs(2199) <= '1';
    layer1_outputs(2200) <= (layer0_outputs(1982)) or (layer0_outputs(1710));
    layer1_outputs(2201) <= not(layer0_outputs(2453)) or (layer0_outputs(646));
    layer1_outputs(2202) <= (layer0_outputs(2177)) and (layer0_outputs(482));
    layer1_outputs(2203) <= not(layer0_outputs(1618));
    layer1_outputs(2204) <= (layer0_outputs(482)) or (layer0_outputs(798));
    layer1_outputs(2205) <= not(layer0_outputs(1582));
    layer1_outputs(2206) <= '1';
    layer1_outputs(2207) <= layer0_outputs(1492);
    layer1_outputs(2208) <= layer0_outputs(821);
    layer1_outputs(2209) <= not((layer0_outputs(1072)) or (layer0_outputs(1675)));
    layer1_outputs(2210) <= '1';
    layer1_outputs(2211) <= not(layer0_outputs(555)) or (layer0_outputs(830));
    layer1_outputs(2212) <= not(layer0_outputs(719));
    layer1_outputs(2213) <= not((layer0_outputs(2379)) or (layer0_outputs(2318)));
    layer1_outputs(2214) <= not(layer0_outputs(1068)) or (layer0_outputs(671));
    layer1_outputs(2215) <= not(layer0_outputs(1580));
    layer1_outputs(2216) <= '1';
    layer1_outputs(2217) <= not((layer0_outputs(1599)) and (layer0_outputs(241)));
    layer1_outputs(2218) <= '0';
    layer1_outputs(2219) <= not((layer0_outputs(2014)) and (layer0_outputs(475)));
    layer1_outputs(2220) <= '1';
    layer1_outputs(2221) <= not((layer0_outputs(1486)) and (layer0_outputs(226)));
    layer1_outputs(2222) <= not((layer0_outputs(2156)) and (layer0_outputs(1176)));
    layer1_outputs(2223) <= (layer0_outputs(122)) and not (layer0_outputs(705));
    layer1_outputs(2224) <= (layer0_outputs(1377)) xor (layer0_outputs(1663));
    layer1_outputs(2225) <= (layer0_outputs(861)) or (layer0_outputs(872));
    layer1_outputs(2226) <= '0';
    layer1_outputs(2227) <= not(layer0_outputs(2422));
    layer1_outputs(2228) <= not((layer0_outputs(1205)) or (layer0_outputs(2411)));
    layer1_outputs(2229) <= (layer0_outputs(2466)) or (layer0_outputs(1374));
    layer1_outputs(2230) <= (layer0_outputs(1972)) or (layer0_outputs(1989));
    layer1_outputs(2231) <= not(layer0_outputs(1627));
    layer1_outputs(2232) <= (layer0_outputs(1384)) and not (layer0_outputs(1666));
    layer1_outputs(2233) <= not((layer0_outputs(332)) and (layer0_outputs(881)));
    layer1_outputs(2234) <= layer0_outputs(1685);
    layer1_outputs(2235) <= not((layer0_outputs(1960)) or (layer0_outputs(1825)));
    layer1_outputs(2236) <= (layer0_outputs(529)) and not (layer0_outputs(1847));
    layer1_outputs(2237) <= '0';
    layer1_outputs(2238) <= layer0_outputs(103);
    layer1_outputs(2239) <= not(layer0_outputs(1934));
    layer1_outputs(2240) <= not(layer0_outputs(629));
    layer1_outputs(2241) <= '1';
    layer1_outputs(2242) <= (layer0_outputs(2184)) or (layer0_outputs(1603));
    layer1_outputs(2243) <= layer0_outputs(1619);
    layer1_outputs(2244) <= '0';
    layer1_outputs(2245) <= not((layer0_outputs(869)) and (layer0_outputs(2013)));
    layer1_outputs(2246) <= layer0_outputs(209);
    layer1_outputs(2247) <= layer0_outputs(1007);
    layer1_outputs(2248) <= not(layer0_outputs(1272));
    layer1_outputs(2249) <= (layer0_outputs(1056)) and (layer0_outputs(1578));
    layer1_outputs(2250) <= not((layer0_outputs(721)) or (layer0_outputs(1653)));
    layer1_outputs(2251) <= '0';
    layer1_outputs(2252) <= not((layer0_outputs(1625)) or (layer0_outputs(2485)));
    layer1_outputs(2253) <= layer0_outputs(1770);
    layer1_outputs(2254) <= not(layer0_outputs(800));
    layer1_outputs(2255) <= (layer0_outputs(749)) or (layer0_outputs(1138));
    layer1_outputs(2256) <= '1';
    layer1_outputs(2257) <= '0';
    layer1_outputs(2258) <= not((layer0_outputs(1532)) and (layer0_outputs(1378)));
    layer1_outputs(2259) <= (layer0_outputs(2181)) xor (layer0_outputs(465));
    layer1_outputs(2260) <= (layer0_outputs(1444)) or (layer0_outputs(86));
    layer1_outputs(2261) <= (layer0_outputs(516)) or (layer0_outputs(2039));
    layer1_outputs(2262) <= '1';
    layer1_outputs(2263) <= (layer0_outputs(499)) and not (layer0_outputs(2411));
    layer1_outputs(2264) <= '1';
    layer1_outputs(2265) <= not((layer0_outputs(531)) or (layer0_outputs(457)));
    layer1_outputs(2266) <= not((layer0_outputs(1665)) or (layer0_outputs(812)));
    layer1_outputs(2267) <= '1';
    layer1_outputs(2268) <= layer0_outputs(434);
    layer1_outputs(2269) <= layer0_outputs(979);
    layer1_outputs(2270) <= layer0_outputs(289);
    layer1_outputs(2271) <= not(layer0_outputs(1553));
    layer1_outputs(2272) <= layer0_outputs(2211);
    layer1_outputs(2273) <= not(layer0_outputs(2490));
    layer1_outputs(2274) <= not((layer0_outputs(477)) and (layer0_outputs(25)));
    layer1_outputs(2275) <= '1';
    layer1_outputs(2276) <= not(layer0_outputs(221)) or (layer0_outputs(2206));
    layer1_outputs(2277) <= (layer0_outputs(1922)) and (layer0_outputs(1645));
    layer1_outputs(2278) <= '1';
    layer1_outputs(2279) <= not(layer0_outputs(2251));
    layer1_outputs(2280) <= (layer0_outputs(2412)) and not (layer0_outputs(789));
    layer1_outputs(2281) <= layer0_outputs(1200);
    layer1_outputs(2282) <= '0';
    layer1_outputs(2283) <= (layer0_outputs(1115)) and (layer0_outputs(615));
    layer1_outputs(2284) <= not((layer0_outputs(2255)) or (layer0_outputs(105)));
    layer1_outputs(2285) <= (layer0_outputs(285)) and not (layer0_outputs(1864));
    layer1_outputs(2286) <= (layer0_outputs(855)) and not (layer0_outputs(1181));
    layer1_outputs(2287) <= '1';
    layer1_outputs(2288) <= not(layer0_outputs(783));
    layer1_outputs(2289) <= not(layer0_outputs(1359));
    layer1_outputs(2290) <= '0';
    layer1_outputs(2291) <= not((layer0_outputs(2119)) and (layer0_outputs(1446)));
    layer1_outputs(2292) <= '0';
    layer1_outputs(2293) <= not((layer0_outputs(1821)) and (layer0_outputs(1042)));
    layer1_outputs(2294) <= '1';
    layer1_outputs(2295) <= not((layer0_outputs(1059)) or (layer0_outputs(715)));
    layer1_outputs(2296) <= (layer0_outputs(2383)) and (layer0_outputs(1112));
    layer1_outputs(2297) <= not((layer0_outputs(247)) and (layer0_outputs(2512)));
    layer1_outputs(2298) <= '1';
    layer1_outputs(2299) <= not((layer0_outputs(944)) or (layer0_outputs(1523)));
    layer1_outputs(2300) <= (layer0_outputs(1529)) and (layer0_outputs(1920));
    layer1_outputs(2301) <= '1';
    layer1_outputs(2302) <= layer0_outputs(608);
    layer1_outputs(2303) <= (layer0_outputs(1243)) or (layer0_outputs(1000));
    layer1_outputs(2304) <= not(layer0_outputs(395));
    layer1_outputs(2305) <= (layer0_outputs(1872)) or (layer0_outputs(1912));
    layer1_outputs(2306) <= '1';
    layer1_outputs(2307) <= '0';
    layer1_outputs(2308) <= not(layer0_outputs(328)) or (layer0_outputs(2435));
    layer1_outputs(2309) <= (layer0_outputs(330)) or (layer0_outputs(484));
    layer1_outputs(2310) <= not(layer0_outputs(2451)) or (layer0_outputs(1964));
    layer1_outputs(2311) <= (layer0_outputs(311)) xor (layer0_outputs(1318));
    layer1_outputs(2312) <= not(layer0_outputs(1356));
    layer1_outputs(2313) <= '1';
    layer1_outputs(2314) <= (layer0_outputs(659)) and not (layer0_outputs(1507));
    layer1_outputs(2315) <= not(layer0_outputs(398)) or (layer0_outputs(801));
    layer1_outputs(2316) <= layer0_outputs(414);
    layer1_outputs(2317) <= '1';
    layer1_outputs(2318) <= layer0_outputs(1414);
    layer1_outputs(2319) <= '1';
    layer1_outputs(2320) <= (layer0_outputs(2092)) and (layer0_outputs(1932));
    layer1_outputs(2321) <= (layer0_outputs(1915)) and (layer0_outputs(1938));
    layer1_outputs(2322) <= '1';
    layer1_outputs(2323) <= not((layer0_outputs(1358)) and (layer0_outputs(1183)));
    layer1_outputs(2324) <= not(layer0_outputs(1942)) or (layer0_outputs(2074));
    layer1_outputs(2325) <= (layer0_outputs(1727)) and not (layer0_outputs(266));
    layer1_outputs(2326) <= layer0_outputs(139);
    layer1_outputs(2327) <= not(layer0_outputs(2115)) or (layer0_outputs(252));
    layer1_outputs(2328) <= not(layer0_outputs(1004)) or (layer0_outputs(1331));
    layer1_outputs(2329) <= not(layer0_outputs(2138));
    layer1_outputs(2330) <= not(layer0_outputs(840)) or (layer0_outputs(979));
    layer1_outputs(2331) <= layer0_outputs(103);
    layer1_outputs(2332) <= '1';
    layer1_outputs(2333) <= '0';
    layer1_outputs(2334) <= not((layer0_outputs(200)) and (layer0_outputs(1698)));
    layer1_outputs(2335) <= (layer0_outputs(1848)) or (layer0_outputs(303));
    layer1_outputs(2336) <= (layer0_outputs(1460)) and (layer0_outputs(2118));
    layer1_outputs(2337) <= not(layer0_outputs(2227));
    layer1_outputs(2338) <= (layer0_outputs(455)) and (layer0_outputs(954));
    layer1_outputs(2339) <= (layer0_outputs(2049)) and (layer0_outputs(989));
    layer1_outputs(2340) <= (layer0_outputs(396)) and not (layer0_outputs(196));
    layer1_outputs(2341) <= '1';
    layer1_outputs(2342) <= not(layer0_outputs(310));
    layer1_outputs(2343) <= not((layer0_outputs(589)) or (layer0_outputs(2458)));
    layer1_outputs(2344) <= '1';
    layer1_outputs(2345) <= '1';
    layer1_outputs(2346) <= not((layer0_outputs(1523)) or (layer0_outputs(1573)));
    layer1_outputs(2347) <= not(layer0_outputs(48));
    layer1_outputs(2348) <= (layer0_outputs(537)) or (layer0_outputs(2452));
    layer1_outputs(2349) <= '0';
    layer1_outputs(2350) <= (layer0_outputs(1454)) and (layer0_outputs(410));
    layer1_outputs(2351) <= not(layer0_outputs(2035));
    layer1_outputs(2352) <= layer0_outputs(1453);
    layer1_outputs(2353) <= not(layer0_outputs(1152));
    layer1_outputs(2354) <= not((layer0_outputs(2032)) or (layer0_outputs(1790)));
    layer1_outputs(2355) <= not(layer0_outputs(2393)) or (layer0_outputs(356));
    layer1_outputs(2356) <= layer0_outputs(1648);
    layer1_outputs(2357) <= not((layer0_outputs(2513)) and (layer0_outputs(636)));
    layer1_outputs(2358) <= layer0_outputs(340);
    layer1_outputs(2359) <= (layer0_outputs(2166)) and not (layer0_outputs(1512));
    layer1_outputs(2360) <= not(layer0_outputs(1757)) or (layer0_outputs(2408));
    layer1_outputs(2361) <= layer0_outputs(1885);
    layer1_outputs(2362) <= not(layer0_outputs(612)) or (layer0_outputs(2209));
    layer1_outputs(2363) <= '1';
    layer1_outputs(2364) <= (layer0_outputs(2079)) and not (layer0_outputs(1910));
    layer1_outputs(2365) <= not(layer0_outputs(1600)) or (layer0_outputs(926));
    layer1_outputs(2366) <= '1';
    layer1_outputs(2367) <= layer0_outputs(1997);
    layer1_outputs(2368) <= '1';
    layer1_outputs(2369) <= (layer0_outputs(4)) and not (layer0_outputs(941));
    layer1_outputs(2370) <= (layer0_outputs(1442)) and (layer0_outputs(214));
    layer1_outputs(2371) <= not((layer0_outputs(542)) and (layer0_outputs(2420)));
    layer1_outputs(2372) <= not(layer0_outputs(490)) or (layer0_outputs(532));
    layer1_outputs(2373) <= '1';
    layer1_outputs(2374) <= '1';
    layer1_outputs(2375) <= layer0_outputs(1627);
    layer1_outputs(2376) <= (layer0_outputs(1738)) and (layer0_outputs(233));
    layer1_outputs(2377) <= not(layer0_outputs(1516));
    layer1_outputs(2378) <= layer0_outputs(2189);
    layer1_outputs(2379) <= layer0_outputs(2438);
    layer1_outputs(2380) <= not((layer0_outputs(632)) and (layer0_outputs(1714)));
    layer1_outputs(2381) <= '0';
    layer1_outputs(2382) <= not(layer0_outputs(781));
    layer1_outputs(2383) <= (layer0_outputs(1884)) and not (layer0_outputs(1376));
    layer1_outputs(2384) <= not((layer0_outputs(2480)) or (layer0_outputs(2002)));
    layer1_outputs(2385) <= '0';
    layer1_outputs(2386) <= (layer0_outputs(1723)) and not (layer0_outputs(1573));
    layer1_outputs(2387) <= not(layer0_outputs(2273));
    layer1_outputs(2388) <= '0';
    layer1_outputs(2389) <= not(layer0_outputs(533));
    layer1_outputs(2390) <= '0';
    layer1_outputs(2391) <= (layer0_outputs(2374)) and not (layer0_outputs(2472));
    layer1_outputs(2392) <= not(layer0_outputs(2485)) or (layer0_outputs(2308));
    layer1_outputs(2393) <= '1';
    layer1_outputs(2394) <= (layer0_outputs(1236)) or (layer0_outputs(1926));
    layer1_outputs(2395) <= (layer0_outputs(1404)) or (layer0_outputs(1462));
    layer1_outputs(2396) <= '1';
    layer1_outputs(2397) <= not(layer0_outputs(539));
    layer1_outputs(2398) <= (layer0_outputs(177)) and not (layer0_outputs(302));
    layer1_outputs(2399) <= (layer0_outputs(1500)) and (layer0_outputs(1588));
    layer1_outputs(2400) <= '1';
    layer1_outputs(2401) <= not(layer0_outputs(809));
    layer1_outputs(2402) <= not((layer0_outputs(1993)) and (layer0_outputs(778)));
    layer1_outputs(2403) <= not(layer0_outputs(1704)) or (layer0_outputs(1559));
    layer1_outputs(2404) <= not(layer0_outputs(1829));
    layer1_outputs(2405) <= not(layer0_outputs(770)) or (layer0_outputs(321));
    layer1_outputs(2406) <= not(layer0_outputs(2462));
    layer1_outputs(2407) <= not(layer0_outputs(14));
    layer1_outputs(2408) <= (layer0_outputs(2271)) or (layer0_outputs(1312));
    layer1_outputs(2409) <= '0';
    layer1_outputs(2410) <= not(layer0_outputs(838)) or (layer0_outputs(2526));
    layer1_outputs(2411) <= layer0_outputs(518);
    layer1_outputs(2412) <= not((layer0_outputs(1958)) and (layer0_outputs(1375)));
    layer1_outputs(2413) <= '0';
    layer1_outputs(2414) <= not(layer0_outputs(1545)) or (layer0_outputs(128));
    layer1_outputs(2415) <= '1';
    layer1_outputs(2416) <= '1';
    layer1_outputs(2417) <= not(layer0_outputs(1416));
    layer1_outputs(2418) <= '0';
    layer1_outputs(2419) <= not((layer0_outputs(1813)) and (layer0_outputs(413)));
    layer1_outputs(2420) <= layer0_outputs(2104);
    layer1_outputs(2421) <= (layer0_outputs(274)) or (layer0_outputs(907));
    layer1_outputs(2422) <= (layer0_outputs(194)) and not (layer0_outputs(583));
    layer1_outputs(2423) <= '0';
    layer1_outputs(2424) <= (layer0_outputs(1428)) and (layer0_outputs(2005));
    layer1_outputs(2425) <= not((layer0_outputs(2128)) and (layer0_outputs(1313)));
    layer1_outputs(2426) <= '1';
    layer1_outputs(2427) <= '1';
    layer1_outputs(2428) <= not((layer0_outputs(1838)) and (layer0_outputs(1718)));
    layer1_outputs(2429) <= layer0_outputs(49);
    layer1_outputs(2430) <= not((layer0_outputs(279)) or (layer0_outputs(666)));
    layer1_outputs(2431) <= not(layer0_outputs(353)) or (layer0_outputs(1645));
    layer1_outputs(2432) <= not((layer0_outputs(273)) or (layer0_outputs(2509)));
    layer1_outputs(2433) <= not((layer0_outputs(180)) or (layer0_outputs(1851)));
    layer1_outputs(2434) <= '0';
    layer1_outputs(2435) <= not((layer0_outputs(1268)) and (layer0_outputs(2236)));
    layer1_outputs(2436) <= '1';
    layer1_outputs(2437) <= (layer0_outputs(403)) and not (layer0_outputs(1288));
    layer1_outputs(2438) <= layer0_outputs(2354);
    layer1_outputs(2439) <= not((layer0_outputs(551)) and (layer0_outputs(2183)));
    layer1_outputs(2440) <= not(layer0_outputs(2159)) or (layer0_outputs(730));
    layer1_outputs(2441) <= not((layer0_outputs(1729)) and (layer0_outputs(469)));
    layer1_outputs(2442) <= not((layer0_outputs(24)) and (layer0_outputs(1751)));
    layer1_outputs(2443) <= '1';
    layer1_outputs(2444) <= (layer0_outputs(2020)) and (layer0_outputs(2048));
    layer1_outputs(2445) <= '0';
    layer1_outputs(2446) <= (layer0_outputs(1818)) and not (layer0_outputs(2546));
    layer1_outputs(2447) <= '1';
    layer1_outputs(2448) <= (layer0_outputs(2207)) and not (layer0_outputs(1610));
    layer1_outputs(2449) <= not((layer0_outputs(1417)) or (layer0_outputs(360)));
    layer1_outputs(2450) <= '1';
    layer1_outputs(2451) <= not(layer0_outputs(1401)) or (layer0_outputs(561));
    layer1_outputs(2452) <= '0';
    layer1_outputs(2453) <= '0';
    layer1_outputs(2454) <= '1';
    layer1_outputs(2455) <= not(layer0_outputs(2314));
    layer1_outputs(2456) <= (layer0_outputs(2340)) or (layer0_outputs(191));
    layer1_outputs(2457) <= '0';
    layer1_outputs(2458) <= (layer0_outputs(1780)) or (layer0_outputs(391));
    layer1_outputs(2459) <= not((layer0_outputs(2471)) and (layer0_outputs(2099)));
    layer1_outputs(2460) <= not(layer0_outputs(280));
    layer1_outputs(2461) <= layer0_outputs(1055);
    layer1_outputs(2462) <= layer0_outputs(2522);
    layer1_outputs(2463) <= layer0_outputs(939);
    layer1_outputs(2464) <= (layer0_outputs(1399)) and not (layer0_outputs(725));
    layer1_outputs(2465) <= not((layer0_outputs(275)) or (layer0_outputs(48)));
    layer1_outputs(2466) <= '0';
    layer1_outputs(2467) <= not(layer0_outputs(2155)) or (layer0_outputs(485));
    layer1_outputs(2468) <= (layer0_outputs(2244)) and not (layer0_outputs(1139));
    layer1_outputs(2469) <= not(layer0_outputs(852)) or (layer0_outputs(2090));
    layer1_outputs(2470) <= '0';
    layer1_outputs(2471) <= not((layer0_outputs(815)) and (layer0_outputs(2149)));
    layer1_outputs(2472) <= layer0_outputs(541);
    layer1_outputs(2473) <= not(layer0_outputs(1409));
    layer1_outputs(2474) <= not(layer0_outputs(242));
    layer1_outputs(2475) <= (layer0_outputs(532)) and not (layer0_outputs(2213));
    layer1_outputs(2476) <= not(layer0_outputs(1917)) or (layer0_outputs(1279));
    layer1_outputs(2477) <= not((layer0_outputs(1135)) and (layer0_outputs(378)));
    layer1_outputs(2478) <= not(layer0_outputs(1091)) or (layer0_outputs(127));
    layer1_outputs(2479) <= (layer0_outputs(2455)) and not (layer0_outputs(2207));
    layer1_outputs(2480) <= (layer0_outputs(1379)) and (layer0_outputs(472));
    layer1_outputs(2481) <= '0';
    layer1_outputs(2482) <= not(layer0_outputs(1681));
    layer1_outputs(2483) <= not(layer0_outputs(1114)) or (layer0_outputs(2241));
    layer1_outputs(2484) <= layer0_outputs(893);
    layer1_outputs(2485) <= '1';
    layer1_outputs(2486) <= '0';
    layer1_outputs(2487) <= (layer0_outputs(294)) and not (layer0_outputs(1905));
    layer1_outputs(2488) <= (layer0_outputs(1016)) or (layer0_outputs(2042));
    layer1_outputs(2489) <= not(layer0_outputs(468));
    layer1_outputs(2490) <= '0';
    layer1_outputs(2491) <= '1';
    layer1_outputs(2492) <= not(layer0_outputs(1744)) or (layer0_outputs(1157));
    layer1_outputs(2493) <= '0';
    layer1_outputs(2494) <= not(layer0_outputs(1201)) or (layer0_outputs(1863));
    layer1_outputs(2495) <= layer0_outputs(1218);
    layer1_outputs(2496) <= '1';
    layer1_outputs(2497) <= (layer0_outputs(1329)) and not (layer0_outputs(717));
    layer1_outputs(2498) <= '0';
    layer1_outputs(2499) <= not((layer0_outputs(2234)) and (layer0_outputs(1726)));
    layer1_outputs(2500) <= layer0_outputs(799);
    layer1_outputs(2501) <= '1';
    layer1_outputs(2502) <= not(layer0_outputs(89)) or (layer0_outputs(1113));
    layer1_outputs(2503) <= '0';
    layer1_outputs(2504) <= not((layer0_outputs(347)) xor (layer0_outputs(109)));
    layer1_outputs(2505) <= (layer0_outputs(607)) and (layer0_outputs(1946));
    layer1_outputs(2506) <= not(layer0_outputs(1263)) or (layer0_outputs(1461));
    layer1_outputs(2507) <= '1';
    layer1_outputs(2508) <= layer0_outputs(1381);
    layer1_outputs(2509) <= layer0_outputs(1609);
    layer1_outputs(2510) <= layer0_outputs(2186);
    layer1_outputs(2511) <= not(layer0_outputs(1606)) or (layer0_outputs(2373));
    layer1_outputs(2512) <= not((layer0_outputs(1634)) or (layer0_outputs(2096)));
    layer1_outputs(2513) <= not(layer0_outputs(2064));
    layer1_outputs(2514) <= '1';
    layer1_outputs(2515) <= not((layer0_outputs(2312)) and (layer0_outputs(891)));
    layer1_outputs(2516) <= not((layer0_outputs(1274)) xor (layer0_outputs(455)));
    layer1_outputs(2517) <= not(layer0_outputs(1382)) or (layer0_outputs(358));
    layer1_outputs(2518) <= '1';
    layer1_outputs(2519) <= layer0_outputs(42);
    layer1_outputs(2520) <= not((layer0_outputs(153)) or (layer0_outputs(2385)));
    layer1_outputs(2521) <= layer0_outputs(1390);
    layer1_outputs(2522) <= layer0_outputs(1649);
    layer1_outputs(2523) <= not((layer0_outputs(1683)) or (layer0_outputs(256)));
    layer1_outputs(2524) <= layer0_outputs(488);
    layer1_outputs(2525) <= (layer0_outputs(374)) and (layer0_outputs(134));
    layer1_outputs(2526) <= not(layer0_outputs(1128));
    layer1_outputs(2527) <= (layer0_outputs(2543)) or (layer0_outputs(2507));
    layer1_outputs(2528) <= not(layer0_outputs(1651)) or (layer0_outputs(441));
    layer1_outputs(2529) <= '0';
    layer1_outputs(2530) <= '1';
    layer1_outputs(2531) <= not(layer0_outputs(268)) or (layer0_outputs(521));
    layer1_outputs(2532) <= (layer0_outputs(1203)) and not (layer0_outputs(2132));
    layer1_outputs(2533) <= not(layer0_outputs(2405));
    layer1_outputs(2534) <= layer0_outputs(1635);
    layer1_outputs(2535) <= (layer0_outputs(362)) and not (layer0_outputs(446));
    layer1_outputs(2536) <= not((layer0_outputs(461)) or (layer0_outputs(2396)));
    layer1_outputs(2537) <= layer0_outputs(2461);
    layer1_outputs(2538) <= (layer0_outputs(1097)) or (layer0_outputs(1846));
    layer1_outputs(2539) <= (layer0_outputs(854)) and (layer0_outputs(1026));
    layer1_outputs(2540) <= (layer0_outputs(1639)) and (layer0_outputs(2552));
    layer1_outputs(2541) <= '1';
    layer1_outputs(2542) <= not(layer0_outputs(802)) or (layer0_outputs(412));
    layer1_outputs(2543) <= (layer0_outputs(414)) and (layer0_outputs(202));
    layer1_outputs(2544) <= '1';
    layer1_outputs(2545) <= not((layer0_outputs(2087)) xor (layer0_outputs(2043)));
    layer1_outputs(2546) <= not((layer0_outputs(2267)) xor (layer0_outputs(780)));
    layer1_outputs(2547) <= layer0_outputs(1725);
    layer1_outputs(2548) <= (layer0_outputs(1368)) or (layer0_outputs(821));
    layer1_outputs(2549) <= not((layer0_outputs(2286)) or (layer0_outputs(1160)));
    layer1_outputs(2550) <= not(layer0_outputs(902));
    layer1_outputs(2551) <= (layer0_outputs(658)) and not (layer0_outputs(509));
    layer1_outputs(2552) <= (layer0_outputs(2008)) and (layer0_outputs(2025));
    layer1_outputs(2553) <= not(layer0_outputs(1525));
    layer1_outputs(2554) <= layer0_outputs(39);
    layer1_outputs(2555) <= '0';
    layer1_outputs(2556) <= (layer0_outputs(1276)) or (layer0_outputs(174));
    layer1_outputs(2557) <= (layer0_outputs(736)) and not (layer0_outputs(1484));
    layer1_outputs(2558) <= layer0_outputs(909);
    layer1_outputs(2559) <= (layer0_outputs(1540)) or (layer0_outputs(2358));
    layer2_outputs(0) <= layer1_outputs(1645);
    layer2_outputs(1) <= not(layer1_outputs(1811));
    layer2_outputs(2) <= not((layer1_outputs(920)) or (layer1_outputs(7)));
    layer2_outputs(3) <= not(layer1_outputs(199));
    layer2_outputs(4) <= not((layer1_outputs(4)) and (layer1_outputs(1071)));
    layer2_outputs(5) <= layer1_outputs(1247);
    layer2_outputs(6) <= not(layer1_outputs(6));
    layer2_outputs(7) <= layer1_outputs(893);
    layer2_outputs(8) <= '1';
    layer2_outputs(9) <= '0';
    layer2_outputs(10) <= not((layer1_outputs(1452)) and (layer1_outputs(503)));
    layer2_outputs(11) <= layer1_outputs(580);
    layer2_outputs(12) <= not(layer1_outputs(1378));
    layer2_outputs(13) <= not((layer1_outputs(830)) or (layer1_outputs(245)));
    layer2_outputs(14) <= layer1_outputs(1825);
    layer2_outputs(15) <= not((layer1_outputs(2067)) xor (layer1_outputs(1995)));
    layer2_outputs(16) <= layer1_outputs(1652);
    layer2_outputs(17) <= not(layer1_outputs(273));
    layer2_outputs(18) <= (layer1_outputs(1419)) or (layer1_outputs(775));
    layer2_outputs(19) <= layer1_outputs(1401);
    layer2_outputs(20) <= '0';
    layer2_outputs(21) <= '0';
    layer2_outputs(22) <= layer1_outputs(1372);
    layer2_outputs(23) <= not((layer1_outputs(1984)) and (layer1_outputs(1142)));
    layer2_outputs(24) <= (layer1_outputs(917)) and not (layer1_outputs(692));
    layer2_outputs(25) <= (layer1_outputs(1812)) and not (layer1_outputs(174));
    layer2_outputs(26) <= not(layer1_outputs(1950)) or (layer1_outputs(1739));
    layer2_outputs(27) <= layer1_outputs(118);
    layer2_outputs(28) <= layer1_outputs(499);
    layer2_outputs(29) <= not(layer1_outputs(740));
    layer2_outputs(30) <= (layer1_outputs(75)) and (layer1_outputs(1027));
    layer2_outputs(31) <= '1';
    layer2_outputs(32) <= layer1_outputs(374);
    layer2_outputs(33) <= (layer1_outputs(1028)) and not (layer1_outputs(817));
    layer2_outputs(34) <= '0';
    layer2_outputs(35) <= (layer1_outputs(1478)) and not (layer1_outputs(1453));
    layer2_outputs(36) <= layer1_outputs(1060);
    layer2_outputs(37) <= '0';
    layer2_outputs(38) <= (layer1_outputs(988)) or (layer1_outputs(1762));
    layer2_outputs(39) <= '0';
    layer2_outputs(40) <= not((layer1_outputs(602)) or (layer1_outputs(1009)));
    layer2_outputs(41) <= (layer1_outputs(2232)) and not (layer1_outputs(947));
    layer2_outputs(42) <= (layer1_outputs(2223)) and not (layer1_outputs(849));
    layer2_outputs(43) <= not(layer1_outputs(2546)) or (layer1_outputs(2311));
    layer2_outputs(44) <= not((layer1_outputs(730)) or (layer1_outputs(1250)));
    layer2_outputs(45) <= not(layer1_outputs(2423)) or (layer1_outputs(651));
    layer2_outputs(46) <= (layer1_outputs(545)) and (layer1_outputs(1774));
    layer2_outputs(47) <= (layer1_outputs(1285)) and (layer1_outputs(1599));
    layer2_outputs(48) <= '0';
    layer2_outputs(49) <= (layer1_outputs(1099)) and not (layer1_outputs(50));
    layer2_outputs(50) <= layer1_outputs(822);
    layer2_outputs(51) <= not(layer1_outputs(1056));
    layer2_outputs(52) <= not((layer1_outputs(1371)) or (layer1_outputs(660)));
    layer2_outputs(53) <= (layer1_outputs(936)) xor (layer1_outputs(2065));
    layer2_outputs(54) <= not((layer1_outputs(421)) or (layer1_outputs(2294)));
    layer2_outputs(55) <= layer1_outputs(1035);
    layer2_outputs(56) <= (layer1_outputs(1443)) or (layer1_outputs(581));
    layer2_outputs(57) <= layer1_outputs(498);
    layer2_outputs(58) <= (layer1_outputs(657)) and not (layer1_outputs(1150));
    layer2_outputs(59) <= not((layer1_outputs(2158)) and (layer1_outputs(2027)));
    layer2_outputs(60) <= (layer1_outputs(2414)) and not (layer1_outputs(2284));
    layer2_outputs(61) <= (layer1_outputs(1807)) and (layer1_outputs(1673));
    layer2_outputs(62) <= not(layer1_outputs(1795));
    layer2_outputs(63) <= (layer1_outputs(1627)) or (layer1_outputs(2318));
    layer2_outputs(64) <= not(layer1_outputs(982)) or (layer1_outputs(143));
    layer2_outputs(65) <= not(layer1_outputs(2201));
    layer2_outputs(66) <= (layer1_outputs(2412)) xor (layer1_outputs(2525));
    layer2_outputs(67) <= not(layer1_outputs(259));
    layer2_outputs(68) <= (layer1_outputs(2540)) and not (layer1_outputs(2058));
    layer2_outputs(69) <= not(layer1_outputs(810)) or (layer1_outputs(473));
    layer2_outputs(70) <= (layer1_outputs(1928)) and (layer1_outputs(2481));
    layer2_outputs(71) <= not(layer1_outputs(1046)) or (layer1_outputs(2178));
    layer2_outputs(72) <= (layer1_outputs(1569)) and (layer1_outputs(1331));
    layer2_outputs(73) <= not(layer1_outputs(699));
    layer2_outputs(74) <= '1';
    layer2_outputs(75) <= (layer1_outputs(140)) or (layer1_outputs(183));
    layer2_outputs(76) <= not(layer1_outputs(2124));
    layer2_outputs(77) <= '1';
    layer2_outputs(78) <= not(layer1_outputs(826));
    layer2_outputs(79) <= (layer1_outputs(1298)) xor (layer1_outputs(1995));
    layer2_outputs(80) <= (layer1_outputs(1985)) and not (layer1_outputs(1193));
    layer2_outputs(81) <= '0';
    layer2_outputs(82) <= (layer1_outputs(541)) and (layer1_outputs(650));
    layer2_outputs(83) <= (layer1_outputs(486)) and (layer1_outputs(1731));
    layer2_outputs(84) <= not((layer1_outputs(169)) and (layer1_outputs(465)));
    layer2_outputs(85) <= (layer1_outputs(1864)) xor (layer1_outputs(244));
    layer2_outputs(86) <= (layer1_outputs(483)) and not (layer1_outputs(2537));
    layer2_outputs(87) <= not((layer1_outputs(2503)) and (layer1_outputs(634)));
    layer2_outputs(88) <= (layer1_outputs(2349)) and not (layer1_outputs(385));
    layer2_outputs(89) <= not(layer1_outputs(341));
    layer2_outputs(90) <= not((layer1_outputs(390)) or (layer1_outputs(2372)));
    layer2_outputs(91) <= layer1_outputs(2327);
    layer2_outputs(92) <= not(layer1_outputs(151)) or (layer1_outputs(1525));
    layer2_outputs(93) <= not(layer1_outputs(2266));
    layer2_outputs(94) <= (layer1_outputs(486)) or (layer1_outputs(377));
    layer2_outputs(95) <= not((layer1_outputs(2188)) or (layer1_outputs(2098)));
    layer2_outputs(96) <= layer1_outputs(2060);
    layer2_outputs(97) <= '0';
    layer2_outputs(98) <= layer1_outputs(1862);
    layer2_outputs(99) <= layer1_outputs(2146);
    layer2_outputs(100) <= (layer1_outputs(854)) and not (layer1_outputs(2307));
    layer2_outputs(101) <= not(layer1_outputs(719)) or (layer1_outputs(1471));
    layer2_outputs(102) <= (layer1_outputs(1946)) and (layer1_outputs(237));
    layer2_outputs(103) <= layer1_outputs(703);
    layer2_outputs(104) <= '0';
    layer2_outputs(105) <= not(layer1_outputs(1477));
    layer2_outputs(106) <= not(layer1_outputs(1943));
    layer2_outputs(107) <= not(layer1_outputs(108)) or (layer1_outputs(827));
    layer2_outputs(108) <= not(layer1_outputs(131));
    layer2_outputs(109) <= not((layer1_outputs(249)) and (layer1_outputs(1591)));
    layer2_outputs(110) <= not(layer1_outputs(1290));
    layer2_outputs(111) <= '1';
    layer2_outputs(112) <= (layer1_outputs(1001)) and (layer1_outputs(490));
    layer2_outputs(113) <= not(layer1_outputs(1179));
    layer2_outputs(114) <= layer1_outputs(616);
    layer2_outputs(115) <= (layer1_outputs(2515)) or (layer1_outputs(147));
    layer2_outputs(116) <= layer1_outputs(418);
    layer2_outputs(117) <= not(layer1_outputs(20));
    layer2_outputs(118) <= not(layer1_outputs(1835)) or (layer1_outputs(285));
    layer2_outputs(119) <= not(layer1_outputs(1855));
    layer2_outputs(120) <= (layer1_outputs(1555)) or (layer1_outputs(1390));
    layer2_outputs(121) <= layer1_outputs(733);
    layer2_outputs(122) <= not(layer1_outputs(721)) or (layer1_outputs(1424));
    layer2_outputs(123) <= not((layer1_outputs(673)) and (layer1_outputs(1820)));
    layer2_outputs(124) <= '0';
    layer2_outputs(125) <= not(layer1_outputs(1481)) or (layer1_outputs(1557));
    layer2_outputs(126) <= not((layer1_outputs(811)) xor (layer1_outputs(1029)));
    layer2_outputs(127) <= not(layer1_outputs(1555)) or (layer1_outputs(2095));
    layer2_outputs(128) <= not(layer1_outputs(2145)) or (layer1_outputs(2245));
    layer2_outputs(129) <= layer1_outputs(710);
    layer2_outputs(130) <= layer1_outputs(2356);
    layer2_outputs(131) <= not(layer1_outputs(232));
    layer2_outputs(132) <= layer1_outputs(1679);
    layer2_outputs(133) <= not(layer1_outputs(2325)) or (layer1_outputs(25));
    layer2_outputs(134) <= '0';
    layer2_outputs(135) <= not(layer1_outputs(1758)) or (layer1_outputs(813));
    layer2_outputs(136) <= (layer1_outputs(621)) and not (layer1_outputs(2372));
    layer2_outputs(137) <= not(layer1_outputs(538));
    layer2_outputs(138) <= layer1_outputs(961);
    layer2_outputs(139) <= not(layer1_outputs(2191));
    layer2_outputs(140) <= not(layer1_outputs(710)) or (layer1_outputs(1481));
    layer2_outputs(141) <= '1';
    layer2_outputs(142) <= not(layer1_outputs(859)) or (layer1_outputs(1171));
    layer2_outputs(143) <= (layer1_outputs(2001)) or (layer1_outputs(2473));
    layer2_outputs(144) <= (layer1_outputs(1472)) or (layer1_outputs(981));
    layer2_outputs(145) <= not((layer1_outputs(541)) and (layer1_outputs(2459)));
    layer2_outputs(146) <= not(layer1_outputs(663)) or (layer1_outputs(1000));
    layer2_outputs(147) <= (layer1_outputs(2388)) and (layer1_outputs(1563));
    layer2_outputs(148) <= layer1_outputs(2082);
    layer2_outputs(149) <= (layer1_outputs(1821)) and not (layer1_outputs(1830));
    layer2_outputs(150) <= (layer1_outputs(534)) and (layer1_outputs(175));
    layer2_outputs(151) <= not(layer1_outputs(1035));
    layer2_outputs(152) <= layer1_outputs(653);
    layer2_outputs(153) <= (layer1_outputs(789)) and not (layer1_outputs(1503));
    layer2_outputs(154) <= not(layer1_outputs(1284)) or (layer1_outputs(170));
    layer2_outputs(155) <= not(layer1_outputs(2519));
    layer2_outputs(156) <= layer1_outputs(861);
    layer2_outputs(157) <= layer1_outputs(2041);
    layer2_outputs(158) <= not(layer1_outputs(1171));
    layer2_outputs(159) <= (layer1_outputs(315)) and (layer1_outputs(974));
    layer2_outputs(160) <= '0';
    layer2_outputs(161) <= (layer1_outputs(364)) and not (layer1_outputs(601));
    layer2_outputs(162) <= not(layer1_outputs(1134));
    layer2_outputs(163) <= layer1_outputs(1856);
    layer2_outputs(164) <= '0';
    layer2_outputs(165) <= layer1_outputs(240);
    layer2_outputs(166) <= '0';
    layer2_outputs(167) <= (layer1_outputs(643)) and (layer1_outputs(942));
    layer2_outputs(168) <= not(layer1_outputs(1298));
    layer2_outputs(169) <= not(layer1_outputs(2547));
    layer2_outputs(170) <= (layer1_outputs(2488)) and not (layer1_outputs(1846));
    layer2_outputs(171) <= (layer1_outputs(1939)) and not (layer1_outputs(194));
    layer2_outputs(172) <= layer1_outputs(659);
    layer2_outputs(173) <= '1';
    layer2_outputs(174) <= layer1_outputs(2378);
    layer2_outputs(175) <= layer1_outputs(1738);
    layer2_outputs(176) <= not(layer1_outputs(1436));
    layer2_outputs(177) <= layer1_outputs(1959);
    layer2_outputs(178) <= layer1_outputs(1126);
    layer2_outputs(179) <= not(layer1_outputs(1552));
    layer2_outputs(180) <= layer1_outputs(2510);
    layer2_outputs(181) <= '1';
    layer2_outputs(182) <= layer1_outputs(1670);
    layer2_outputs(183) <= not(layer1_outputs(1638));
    layer2_outputs(184) <= '0';
    layer2_outputs(185) <= (layer1_outputs(2)) and not (layer1_outputs(1479));
    layer2_outputs(186) <= not(layer1_outputs(2282)) or (layer1_outputs(316));
    layer2_outputs(187) <= (layer1_outputs(2272)) or (layer1_outputs(2070));
    layer2_outputs(188) <= layer1_outputs(2550);
    layer2_outputs(189) <= not(layer1_outputs(2309)) or (layer1_outputs(1351));
    layer2_outputs(190) <= '1';
    layer2_outputs(191) <= (layer1_outputs(2224)) or (layer1_outputs(2123));
    layer2_outputs(192) <= not(layer1_outputs(1269)) or (layer1_outputs(1200));
    layer2_outputs(193) <= (layer1_outputs(391)) and (layer1_outputs(2290));
    layer2_outputs(194) <= not((layer1_outputs(1664)) and (layer1_outputs(1221)));
    layer2_outputs(195) <= layer1_outputs(743);
    layer2_outputs(196) <= layer1_outputs(264);
    layer2_outputs(197) <= not(layer1_outputs(2214)) or (layer1_outputs(2190));
    layer2_outputs(198) <= '1';
    layer2_outputs(199) <= not((layer1_outputs(1659)) or (layer1_outputs(1147)));
    layer2_outputs(200) <= layer1_outputs(1589);
    layer2_outputs(201) <= (layer1_outputs(258)) and (layer1_outputs(2040));
    layer2_outputs(202) <= not((layer1_outputs(2298)) or (layer1_outputs(571)));
    layer2_outputs(203) <= layer1_outputs(633);
    layer2_outputs(204) <= (layer1_outputs(1193)) or (layer1_outputs(2257));
    layer2_outputs(205) <= '1';
    layer2_outputs(206) <= (layer1_outputs(338)) and not (layer1_outputs(367));
    layer2_outputs(207) <= (layer1_outputs(294)) and not (layer1_outputs(1246));
    layer2_outputs(208) <= '1';
    layer2_outputs(209) <= (layer1_outputs(871)) and (layer1_outputs(1323));
    layer2_outputs(210) <= (layer1_outputs(1751)) and not (layer1_outputs(1017));
    layer2_outputs(211) <= (layer1_outputs(1730)) or (layer1_outputs(1057));
    layer2_outputs(212) <= (layer1_outputs(546)) and not (layer1_outputs(1706));
    layer2_outputs(213) <= not(layer1_outputs(2053));
    layer2_outputs(214) <= not((layer1_outputs(1259)) and (layer1_outputs(396)));
    layer2_outputs(215) <= layer1_outputs(1865);
    layer2_outputs(216) <= '0';
    layer2_outputs(217) <= not((layer1_outputs(998)) or (layer1_outputs(244)));
    layer2_outputs(218) <= layer1_outputs(1160);
    layer2_outputs(219) <= '1';
    layer2_outputs(220) <= '1';
    layer2_outputs(221) <= not(layer1_outputs(1814));
    layer2_outputs(222) <= not(layer1_outputs(2149)) or (layer1_outputs(757));
    layer2_outputs(223) <= not((layer1_outputs(1111)) or (layer1_outputs(768)));
    layer2_outputs(224) <= not(layer1_outputs(701)) or (layer1_outputs(2179));
    layer2_outputs(225) <= layer1_outputs(1476);
    layer2_outputs(226) <= '1';
    layer2_outputs(227) <= not((layer1_outputs(2045)) and (layer1_outputs(1929)));
    layer2_outputs(228) <= layer1_outputs(1947);
    layer2_outputs(229) <= layer1_outputs(197);
    layer2_outputs(230) <= '0';
    layer2_outputs(231) <= '1';
    layer2_outputs(232) <= not(layer1_outputs(180)) or (layer1_outputs(918));
    layer2_outputs(233) <= (layer1_outputs(2115)) and not (layer1_outputs(1584));
    layer2_outputs(234) <= layer1_outputs(195);
    layer2_outputs(235) <= '1';
    layer2_outputs(236) <= not(layer1_outputs(2558));
    layer2_outputs(237) <= not(layer1_outputs(2020));
    layer2_outputs(238) <= (layer1_outputs(585)) and (layer1_outputs(1888));
    layer2_outputs(239) <= '0';
    layer2_outputs(240) <= not((layer1_outputs(1542)) or (layer1_outputs(120)));
    layer2_outputs(241) <= (layer1_outputs(1522)) xor (layer1_outputs(1482));
    layer2_outputs(242) <= layer1_outputs(2039);
    layer2_outputs(243) <= not(layer1_outputs(1898));
    layer2_outputs(244) <= '0';
    layer2_outputs(245) <= '1';
    layer2_outputs(246) <= '0';
    layer2_outputs(247) <= '1';
    layer2_outputs(248) <= layer1_outputs(966);
    layer2_outputs(249) <= not(layer1_outputs(1602)) or (layer1_outputs(1030));
    layer2_outputs(250) <= not(layer1_outputs(2326));
    layer2_outputs(251) <= layer1_outputs(2422);
    layer2_outputs(252) <= layer1_outputs(2483);
    layer2_outputs(253) <= not(layer1_outputs(1939)) or (layer1_outputs(1179));
    layer2_outputs(254) <= not(layer1_outputs(851));
    layer2_outputs(255) <= (layer1_outputs(157)) and (layer1_outputs(1710));
    layer2_outputs(256) <= layer1_outputs(1965);
    layer2_outputs(257) <= not(layer1_outputs(2555)) or (layer1_outputs(1759));
    layer2_outputs(258) <= layer1_outputs(1288);
    layer2_outputs(259) <= (layer1_outputs(611)) and (layer1_outputs(2314));
    layer2_outputs(260) <= not(layer1_outputs(2499));
    layer2_outputs(261) <= (layer1_outputs(1927)) and (layer1_outputs(1900));
    layer2_outputs(262) <= not((layer1_outputs(1938)) and (layer1_outputs(962)));
    layer2_outputs(263) <= '1';
    layer2_outputs(264) <= not((layer1_outputs(2067)) xor (layer1_outputs(1205)));
    layer2_outputs(265) <= not(layer1_outputs(2214)) or (layer1_outputs(1682));
    layer2_outputs(266) <= not(layer1_outputs(504)) or (layer1_outputs(2469));
    layer2_outputs(267) <= layer1_outputs(1988);
    layer2_outputs(268) <= layer1_outputs(2387);
    layer2_outputs(269) <= not(layer1_outputs(2181));
    layer2_outputs(270) <= not(layer1_outputs(430));
    layer2_outputs(271) <= (layer1_outputs(1972)) or (layer1_outputs(1921));
    layer2_outputs(272) <= not(layer1_outputs(391));
    layer2_outputs(273) <= not(layer1_outputs(1374));
    layer2_outputs(274) <= layer1_outputs(831);
    layer2_outputs(275) <= (layer1_outputs(450)) and not (layer1_outputs(1));
    layer2_outputs(276) <= layer1_outputs(2328);
    layer2_outputs(277) <= (layer1_outputs(166)) and not (layer1_outputs(2029));
    layer2_outputs(278) <= not((layer1_outputs(68)) or (layer1_outputs(1130)));
    layer2_outputs(279) <= not((layer1_outputs(1372)) or (layer1_outputs(1450)));
    layer2_outputs(280) <= not(layer1_outputs(2414));
    layer2_outputs(281) <= not(layer1_outputs(537)) or (layer1_outputs(1955));
    layer2_outputs(282) <= layer1_outputs(2354);
    layer2_outputs(283) <= (layer1_outputs(671)) and (layer1_outputs(1623));
    layer2_outputs(284) <= layer1_outputs(2012);
    layer2_outputs(285) <= (layer1_outputs(1767)) xor (layer1_outputs(1417));
    layer2_outputs(286) <= (layer1_outputs(9)) and (layer1_outputs(2481));
    layer2_outputs(287) <= (layer1_outputs(1740)) and not (layer1_outputs(179));
    layer2_outputs(288) <= not(layer1_outputs(1190)) or (layer1_outputs(646));
    layer2_outputs(289) <= '0';
    layer2_outputs(290) <= '0';
    layer2_outputs(291) <= not((layer1_outputs(1451)) or (layer1_outputs(1560)));
    layer2_outputs(292) <= not((layer1_outputs(2379)) and (layer1_outputs(978)));
    layer2_outputs(293) <= not(layer1_outputs(1759));
    layer2_outputs(294) <= not(layer1_outputs(586)) or (layer1_outputs(2386));
    layer2_outputs(295) <= layer1_outputs(2248);
    layer2_outputs(296) <= (layer1_outputs(706)) and not (layer1_outputs(2547));
    layer2_outputs(297) <= (layer1_outputs(1402)) or (layer1_outputs(58));
    layer2_outputs(298) <= layer1_outputs(555);
    layer2_outputs(299) <= not((layer1_outputs(1451)) and (layer1_outputs(2524)));
    layer2_outputs(300) <= (layer1_outputs(1761)) and (layer1_outputs(1531));
    layer2_outputs(301) <= not(layer1_outputs(1241)) or (layer1_outputs(839));
    layer2_outputs(302) <= '0';
    layer2_outputs(303) <= (layer1_outputs(1646)) xor (layer1_outputs(303));
    layer2_outputs(304) <= (layer1_outputs(1265)) and (layer1_outputs(1687));
    layer2_outputs(305) <= layer1_outputs(1797);
    layer2_outputs(306) <= not(layer1_outputs(639)) or (layer1_outputs(1545));
    layer2_outputs(307) <= '1';
    layer2_outputs(308) <= (layer1_outputs(246)) and not (layer1_outputs(912));
    layer2_outputs(309) <= not(layer1_outputs(975));
    layer2_outputs(310) <= not(layer1_outputs(125)) or (layer1_outputs(717));
    layer2_outputs(311) <= (layer1_outputs(2418)) and not (layer1_outputs(319));
    layer2_outputs(312) <= not(layer1_outputs(1870));
    layer2_outputs(313) <= layer1_outputs(1589);
    layer2_outputs(314) <= (layer1_outputs(1456)) and not (layer1_outputs(1944));
    layer2_outputs(315) <= not((layer1_outputs(1443)) and (layer1_outputs(1114)));
    layer2_outputs(316) <= (layer1_outputs(2261)) or (layer1_outputs(2176));
    layer2_outputs(317) <= (layer1_outputs(637)) and not (layer1_outputs(2419));
    layer2_outputs(318) <= '0';
    layer2_outputs(319) <= (layer1_outputs(759)) and not (layer1_outputs(773));
    layer2_outputs(320) <= (layer1_outputs(2458)) and not (layer1_outputs(340));
    layer2_outputs(321) <= layer1_outputs(1280);
    layer2_outputs(322) <= (layer1_outputs(1717)) and not (layer1_outputs(2403));
    layer2_outputs(323) <= layer1_outputs(1176);
    layer2_outputs(324) <= not(layer1_outputs(1765)) or (layer1_outputs(1135));
    layer2_outputs(325) <= not(layer1_outputs(617));
    layer2_outputs(326) <= (layer1_outputs(219)) and not (layer1_outputs(2255));
    layer2_outputs(327) <= (layer1_outputs(1311)) and not (layer1_outputs(19));
    layer2_outputs(328) <= not(layer1_outputs(1820));
    layer2_outputs(329) <= not(layer1_outputs(2389));
    layer2_outputs(330) <= not(layer1_outputs(2461)) or (layer1_outputs(2524));
    layer2_outputs(331) <= not(layer1_outputs(1202));
    layer2_outputs(332) <= (layer1_outputs(320)) and not (layer1_outputs(1079));
    layer2_outputs(333) <= '1';
    layer2_outputs(334) <= (layer1_outputs(2163)) and not (layer1_outputs(1053));
    layer2_outputs(335) <= (layer1_outputs(864)) xor (layer1_outputs(1370));
    layer2_outputs(336) <= not((layer1_outputs(1926)) and (layer1_outputs(595)));
    layer2_outputs(337) <= not(layer1_outputs(378)) or (layer1_outputs(1235));
    layer2_outputs(338) <= (layer1_outputs(902)) and not (layer1_outputs(2186));
    layer2_outputs(339) <= (layer1_outputs(28)) xor (layer1_outputs(2022));
    layer2_outputs(340) <= not(layer1_outputs(526)) or (layer1_outputs(1340));
    layer2_outputs(341) <= not(layer1_outputs(2229));
    layer2_outputs(342) <= not(layer1_outputs(6));
    layer2_outputs(343) <= not(layer1_outputs(655));
    layer2_outputs(344) <= not(layer1_outputs(796)) or (layer1_outputs(2492));
    layer2_outputs(345) <= (layer1_outputs(2365)) and (layer1_outputs(393));
    layer2_outputs(346) <= not(layer1_outputs(1208));
    layer2_outputs(347) <= not(layer1_outputs(442));
    layer2_outputs(348) <= not(layer1_outputs(1050));
    layer2_outputs(349) <= layer1_outputs(2102);
    layer2_outputs(350) <= not((layer1_outputs(1464)) and (layer1_outputs(1894)));
    layer2_outputs(351) <= not(layer1_outputs(2187));
    layer2_outputs(352) <= layer1_outputs(701);
    layer2_outputs(353) <= not(layer1_outputs(46));
    layer2_outputs(354) <= not((layer1_outputs(303)) and (layer1_outputs(737)));
    layer2_outputs(355) <= (layer1_outputs(1385)) or (layer1_outputs(1106));
    layer2_outputs(356) <= not(layer1_outputs(2097)) or (layer1_outputs(1306));
    layer2_outputs(357) <= not(layer1_outputs(2279));
    layer2_outputs(358) <= (layer1_outputs(1335)) and not (layer1_outputs(2197));
    layer2_outputs(359) <= (layer1_outputs(981)) and not (layer1_outputs(2542));
    layer2_outputs(360) <= not((layer1_outputs(612)) and (layer1_outputs(1570)));
    layer2_outputs(361) <= '1';
    layer2_outputs(362) <= (layer1_outputs(328)) or (layer1_outputs(17));
    layer2_outputs(363) <= not(layer1_outputs(2003));
    layer2_outputs(364) <= not(layer1_outputs(1755)) or (layer1_outputs(2527));
    layer2_outputs(365) <= not(layer1_outputs(2351));
    layer2_outputs(366) <= not(layer1_outputs(1069)) or (layer1_outputs(606));
    layer2_outputs(367) <= layer1_outputs(1833);
    layer2_outputs(368) <= not(layer1_outputs(1806));
    layer2_outputs(369) <= not(layer1_outputs(2344)) or (layer1_outputs(113));
    layer2_outputs(370) <= '0';
    layer2_outputs(371) <= not(layer1_outputs(2409)) or (layer1_outputs(1981));
    layer2_outputs(372) <= not(layer1_outputs(715)) or (layer1_outputs(40));
    layer2_outputs(373) <= not(layer1_outputs(479)) or (layer1_outputs(275));
    layer2_outputs(374) <= not(layer1_outputs(641)) or (layer1_outputs(271));
    layer2_outputs(375) <= '1';
    layer2_outputs(376) <= (layer1_outputs(911)) and not (layer1_outputs(1260));
    layer2_outputs(377) <= (layer1_outputs(1996)) and not (layer1_outputs(1399));
    layer2_outputs(378) <= layer1_outputs(1259);
    layer2_outputs(379) <= not(layer1_outputs(2127));
    layer2_outputs(380) <= layer1_outputs(424);
    layer2_outputs(381) <= not(layer1_outputs(862)) or (layer1_outputs(1955));
    layer2_outputs(382) <= layer1_outputs(1484);
    layer2_outputs(383) <= (layer1_outputs(1685)) and not (layer1_outputs(1188));
    layer2_outputs(384) <= not(layer1_outputs(2383)) or (layer1_outputs(1244));
    layer2_outputs(385) <= (layer1_outputs(1688)) and not (layer1_outputs(286));
    layer2_outputs(386) <= '0';
    layer2_outputs(387) <= layer1_outputs(779);
    layer2_outputs(388) <= not(layer1_outputs(917));
    layer2_outputs(389) <= layer1_outputs(2556);
    layer2_outputs(390) <= layer1_outputs(433);
    layer2_outputs(391) <= '1';
    layer2_outputs(392) <= not((layer1_outputs(2353)) and (layer1_outputs(1911)));
    layer2_outputs(393) <= not(layer1_outputs(2463));
    layer2_outputs(394) <= (layer1_outputs(203)) or (layer1_outputs(1637));
    layer2_outputs(395) <= not(layer1_outputs(1043)) or (layer1_outputs(836));
    layer2_outputs(396) <= not((layer1_outputs(614)) or (layer1_outputs(1826)));
    layer2_outputs(397) <= not(layer1_outputs(1111));
    layer2_outputs(398) <= '1';
    layer2_outputs(399) <= (layer1_outputs(647)) and not (layer1_outputs(2428));
    layer2_outputs(400) <= not((layer1_outputs(1701)) or (layer1_outputs(830)));
    layer2_outputs(401) <= not(layer1_outputs(1907));
    layer2_outputs(402) <= not((layer1_outputs(2430)) and (layer1_outputs(424)));
    layer2_outputs(403) <= (layer1_outputs(21)) and not (layer1_outputs(1756));
    layer2_outputs(404) <= not(layer1_outputs(1778)) or (layer1_outputs(1644));
    layer2_outputs(405) <= (layer1_outputs(1848)) or (layer1_outputs(63));
    layer2_outputs(406) <= (layer1_outputs(367)) and not (layer1_outputs(269));
    layer2_outputs(407) <= not(layer1_outputs(1698)) or (layer1_outputs(0));
    layer2_outputs(408) <= (layer1_outputs(178)) or (layer1_outputs(173));
    layer2_outputs(409) <= not((layer1_outputs(969)) and (layer1_outputs(2057)));
    layer2_outputs(410) <= (layer1_outputs(1815)) and not (layer1_outputs(2384));
    layer2_outputs(411) <= layer1_outputs(599);
    layer2_outputs(412) <= '1';
    layer2_outputs(413) <= not((layer1_outputs(819)) or (layer1_outputs(2293)));
    layer2_outputs(414) <= not((layer1_outputs(716)) or (layer1_outputs(780)));
    layer2_outputs(415) <= not(layer1_outputs(2231)) or (layer1_outputs(1469));
    layer2_outputs(416) <= not((layer1_outputs(967)) or (layer1_outputs(2464)));
    layer2_outputs(417) <= layer1_outputs(2209);
    layer2_outputs(418) <= '0';
    layer2_outputs(419) <= not(layer1_outputs(75));
    layer2_outputs(420) <= not(layer1_outputs(913));
    layer2_outputs(421) <= not((layer1_outputs(1528)) or (layer1_outputs(686)));
    layer2_outputs(422) <= (layer1_outputs(1859)) and (layer1_outputs(819));
    layer2_outputs(423) <= '0';
    layer2_outputs(424) <= not(layer1_outputs(800));
    layer2_outputs(425) <= '0';
    layer2_outputs(426) <= not(layer1_outputs(871));
    layer2_outputs(427) <= (layer1_outputs(2032)) or (layer1_outputs(356));
    layer2_outputs(428) <= (layer1_outputs(398)) and (layer1_outputs(213));
    layer2_outputs(429) <= '1';
    layer2_outputs(430) <= (layer1_outputs(2131)) and not (layer1_outputs(2363));
    layer2_outputs(431) <= not((layer1_outputs(1130)) and (layer1_outputs(968)));
    layer2_outputs(432) <= not((layer1_outputs(1142)) or (layer1_outputs(2521)));
    layer2_outputs(433) <= (layer1_outputs(725)) and not (layer1_outputs(2398));
    layer2_outputs(434) <= (layer1_outputs(1234)) or (layer1_outputs(637));
    layer2_outputs(435) <= not(layer1_outputs(1617)) or (layer1_outputs(1872));
    layer2_outputs(436) <= not((layer1_outputs(997)) and (layer1_outputs(1665)));
    layer2_outputs(437) <= (layer1_outputs(2486)) and not (layer1_outputs(154));
    layer2_outputs(438) <= (layer1_outputs(35)) and not (layer1_outputs(1238));
    layer2_outputs(439) <= not(layer1_outputs(499));
    layer2_outputs(440) <= '0';
    layer2_outputs(441) <= not((layer1_outputs(1644)) or (layer1_outputs(1727)));
    layer2_outputs(442) <= (layer1_outputs(150)) and not (layer1_outputs(1072));
    layer2_outputs(443) <= not(layer1_outputs(2228));
    layer2_outputs(444) <= '0';
    layer2_outputs(445) <= (layer1_outputs(1898)) or (layer1_outputs(2112));
    layer2_outputs(446) <= '0';
    layer2_outputs(447) <= (layer1_outputs(1667)) and not (layer1_outputs(1341));
    layer2_outputs(448) <= (layer1_outputs(1640)) or (layer1_outputs(840));
    layer2_outputs(449) <= '0';
    layer2_outputs(450) <= (layer1_outputs(849)) and (layer1_outputs(2163));
    layer2_outputs(451) <= (layer1_outputs(1091)) and not (layer1_outputs(1498));
    layer2_outputs(452) <= '1';
    layer2_outputs(453) <= '0';
    layer2_outputs(454) <= (layer1_outputs(705)) or (layer1_outputs(624));
    layer2_outputs(455) <= layer1_outputs(638);
    layer2_outputs(456) <= (layer1_outputs(825)) and not (layer1_outputs(138));
    layer2_outputs(457) <= (layer1_outputs(2331)) and (layer1_outputs(1045));
    layer2_outputs(458) <= '1';
    layer2_outputs(459) <= (layer1_outputs(1368)) and (layer1_outputs(2217));
    layer2_outputs(460) <= (layer1_outputs(2558)) and not (layer1_outputs(898));
    layer2_outputs(461) <= (layer1_outputs(2124)) or (layer1_outputs(1340));
    layer2_outputs(462) <= not(layer1_outputs(924)) or (layer1_outputs(820));
    layer2_outputs(463) <= not(layer1_outputs(2142)) or (layer1_outputs(794));
    layer2_outputs(464) <= not((layer1_outputs(1267)) and (layer1_outputs(2420)));
    layer2_outputs(465) <= not(layer1_outputs(1137));
    layer2_outputs(466) <= (layer1_outputs(476)) and not (layer1_outputs(1962));
    layer2_outputs(467) <= layer1_outputs(2264);
    layer2_outputs(468) <= not((layer1_outputs(2474)) or (layer1_outputs(2097)));
    layer2_outputs(469) <= (layer1_outputs(816)) and not (layer1_outputs(361));
    layer2_outputs(470) <= not((layer1_outputs(877)) and (layer1_outputs(732)));
    layer2_outputs(471) <= not(layer1_outputs(2068)) or (layer1_outputs(1092));
    layer2_outputs(472) <= (layer1_outputs(2209)) and (layer1_outputs(1415));
    layer2_outputs(473) <= '0';
    layer2_outputs(474) <= (layer1_outputs(71)) and not (layer1_outputs(2271));
    layer2_outputs(475) <= not((layer1_outputs(1839)) or (layer1_outputs(487)));
    layer2_outputs(476) <= (layer1_outputs(403)) and not (layer1_outputs(1989));
    layer2_outputs(477) <= (layer1_outputs(2461)) and not (layer1_outputs(1628));
    layer2_outputs(478) <= '1';
    layer2_outputs(479) <= '1';
    layer2_outputs(480) <= '0';
    layer2_outputs(481) <= layer1_outputs(1883);
    layer2_outputs(482) <= (layer1_outputs(1544)) and not (layer1_outputs(2194));
    layer2_outputs(483) <= not(layer1_outputs(63)) or (layer1_outputs(1525));
    layer2_outputs(484) <= not(layer1_outputs(860)) or (layer1_outputs(1763));
    layer2_outputs(485) <= '1';
    layer2_outputs(486) <= (layer1_outputs(645)) and not (layer1_outputs(1412));
    layer2_outputs(487) <= not((layer1_outputs(1380)) or (layer1_outputs(2034)));
    layer2_outputs(488) <= not(layer1_outputs(2385)) or (layer1_outputs(1553));
    layer2_outputs(489) <= (layer1_outputs(748)) or (layer1_outputs(847));
    layer2_outputs(490) <= layer1_outputs(1489);
    layer2_outputs(491) <= (layer1_outputs(1087)) and not (layer1_outputs(1606));
    layer2_outputs(492) <= not(layer1_outputs(1063));
    layer2_outputs(493) <= not(layer1_outputs(287));
    layer2_outputs(494) <= not((layer1_outputs(1992)) and (layer1_outputs(1155)));
    layer2_outputs(495) <= not(layer1_outputs(1953)) or (layer1_outputs(455));
    layer2_outputs(496) <= not(layer1_outputs(1997));
    layer2_outputs(497) <= (layer1_outputs(1597)) and not (layer1_outputs(644));
    layer2_outputs(498) <= layer1_outputs(714);
    layer2_outputs(499) <= not(layer1_outputs(446)) or (layer1_outputs(1520));
    layer2_outputs(500) <= '1';
    layer2_outputs(501) <= layer1_outputs(539);
    layer2_outputs(502) <= not(layer1_outputs(396)) or (layer1_outputs(1607));
    layer2_outputs(503) <= not(layer1_outputs(2009));
    layer2_outputs(504) <= layer1_outputs(1648);
    layer2_outputs(505) <= not(layer1_outputs(938));
    layer2_outputs(506) <= layer1_outputs(257);
    layer2_outputs(507) <= '1';
    layer2_outputs(508) <= not(layer1_outputs(2261));
    layer2_outputs(509) <= layer1_outputs(1005);
    layer2_outputs(510) <= (layer1_outputs(2443)) xor (layer1_outputs(48));
    layer2_outputs(511) <= layer1_outputs(2402);
    layer2_outputs(512) <= (layer1_outputs(1407)) and not (layer1_outputs(2344));
    layer2_outputs(513) <= not(layer1_outputs(1508));
    layer2_outputs(514) <= (layer1_outputs(409)) and not (layer1_outputs(1868));
    layer2_outputs(515) <= not((layer1_outputs(1145)) and (layer1_outputs(916)));
    layer2_outputs(516) <= layer1_outputs(2535);
    layer2_outputs(517) <= layer1_outputs(2477);
    layer2_outputs(518) <= layer1_outputs(1450);
    layer2_outputs(519) <= layer1_outputs(751);
    layer2_outputs(520) <= not(layer1_outputs(1760)) or (layer1_outputs(1339));
    layer2_outputs(521) <= layer1_outputs(2086);
    layer2_outputs(522) <= layer1_outputs(2202);
    layer2_outputs(523) <= (layer1_outputs(1582)) or (layer1_outputs(1869));
    layer2_outputs(524) <= (layer1_outputs(1015)) and (layer1_outputs(414));
    layer2_outputs(525) <= layer1_outputs(941);
    layer2_outputs(526) <= layer1_outputs(1966);
    layer2_outputs(527) <= not(layer1_outputs(1194)) or (layer1_outputs(1143));
    layer2_outputs(528) <= '1';
    layer2_outputs(529) <= '1';
    layer2_outputs(530) <= not(layer1_outputs(1366));
    layer2_outputs(531) <= (layer1_outputs(471)) or (layer1_outputs(2077));
    layer2_outputs(532) <= not(layer1_outputs(1395)) or (layer1_outputs(381));
    layer2_outputs(533) <= not((layer1_outputs(815)) and (layer1_outputs(985)));
    layer2_outputs(534) <= (layer1_outputs(786)) and not (layer1_outputs(1847));
    layer2_outputs(535) <= '0';
    layer2_outputs(536) <= not((layer1_outputs(1935)) or (layer1_outputs(1594)));
    layer2_outputs(537) <= not(layer1_outputs(731));
    layer2_outputs(538) <= layer1_outputs(1313);
    layer2_outputs(539) <= '1';
    layer2_outputs(540) <= layer1_outputs(2153);
    layer2_outputs(541) <= not((layer1_outputs(1131)) and (layer1_outputs(2420)));
    layer2_outputs(542) <= layer1_outputs(1287);
    layer2_outputs(543) <= not((layer1_outputs(1168)) or (layer1_outputs(904)));
    layer2_outputs(544) <= (layer1_outputs(196)) or (layer1_outputs(2194));
    layer2_outputs(545) <= '1';
    layer2_outputs(546) <= (layer1_outputs(1376)) and not (layer1_outputs(999));
    layer2_outputs(547) <= (layer1_outputs(1354)) xor (layer1_outputs(829));
    layer2_outputs(548) <= not((layer1_outputs(1978)) or (layer1_outputs(2283)));
    layer2_outputs(549) <= (layer1_outputs(1970)) and not (layer1_outputs(1932));
    layer2_outputs(550) <= not(layer1_outputs(1823));
    layer2_outputs(551) <= not(layer1_outputs(2429)) or (layer1_outputs(1997));
    layer2_outputs(552) <= '1';
    layer2_outputs(553) <= '1';
    layer2_outputs(554) <= (layer1_outputs(2405)) and not (layer1_outputs(2542));
    layer2_outputs(555) <= not(layer1_outputs(1650)) or (layer1_outputs(1741));
    layer2_outputs(556) <= not(layer1_outputs(1603)) or (layer1_outputs(2082));
    layer2_outputs(557) <= not((layer1_outputs(176)) or (layer1_outputs(1041)));
    layer2_outputs(558) <= (layer1_outputs(1919)) and not (layer1_outputs(2094));
    layer2_outputs(559) <= (layer1_outputs(1311)) and not (layer1_outputs(1621));
    layer2_outputs(560) <= '1';
    layer2_outputs(561) <= (layer1_outputs(76)) and not (layer1_outputs(1154));
    layer2_outputs(562) <= not((layer1_outputs(757)) and (layer1_outputs(1128)));
    layer2_outputs(563) <= (layer1_outputs(1984)) and not (layer1_outputs(1649));
    layer2_outputs(564) <= layer1_outputs(1126);
    layer2_outputs(565) <= not(layer1_outputs(283));
    layer2_outputs(566) <= not((layer1_outputs(1788)) or (layer1_outputs(1070)));
    layer2_outputs(567) <= (layer1_outputs(1138)) and not (layer1_outputs(1912));
    layer2_outputs(568) <= (layer1_outputs(1271)) and not (layer1_outputs(1314));
    layer2_outputs(569) <= not((layer1_outputs(700)) and (layer1_outputs(506)));
    layer2_outputs(570) <= layer1_outputs(1475);
    layer2_outputs(571) <= (layer1_outputs(2316)) and not (layer1_outputs(2168));
    layer2_outputs(572) <= not(layer1_outputs(1497));
    layer2_outputs(573) <= '1';
    layer2_outputs(574) <= not((layer1_outputs(190)) and (layer1_outputs(1539)));
    layer2_outputs(575) <= '0';
    layer2_outputs(576) <= not((layer1_outputs(2329)) and (layer1_outputs(347)));
    layer2_outputs(577) <= not(layer1_outputs(363));
    layer2_outputs(578) <= '0';
    layer2_outputs(579) <= '0';
    layer2_outputs(580) <= (layer1_outputs(2548)) or (layer1_outputs(1567));
    layer2_outputs(581) <= not(layer1_outputs(2444));
    layer2_outputs(582) <= not(layer1_outputs(1541)) or (layer1_outputs(2005));
    layer2_outputs(583) <= (layer1_outputs(2421)) or (layer1_outputs(1593));
    layer2_outputs(584) <= '0';
    layer2_outputs(585) <= not((layer1_outputs(543)) or (layer1_outputs(684)));
    layer2_outputs(586) <= not(layer1_outputs(508));
    layer2_outputs(587) <= '0';
    layer2_outputs(588) <= not(layer1_outputs(89));
    layer2_outputs(589) <= not((layer1_outputs(1218)) and (layer1_outputs(11)));
    layer2_outputs(590) <= layer1_outputs(254);
    layer2_outputs(591) <= not(layer1_outputs(520)) or (layer1_outputs(1297));
    layer2_outputs(592) <= layer1_outputs(1928);
    layer2_outputs(593) <= not(layer1_outputs(129)) or (layer1_outputs(1121));
    layer2_outputs(594) <= (layer1_outputs(611)) or (layer1_outputs(2112));
    layer2_outputs(595) <= not((layer1_outputs(2504)) and (layer1_outputs(579)));
    layer2_outputs(596) <= not((layer1_outputs(1365)) and (layer1_outputs(1025)));
    layer2_outputs(597) <= layer1_outputs(2348);
    layer2_outputs(598) <= not((layer1_outputs(1613)) and (layer1_outputs(2284)));
    layer2_outputs(599) <= (layer1_outputs(1109)) and not (layer1_outputs(1946));
    layer2_outputs(600) <= not(layer1_outputs(2377));
    layer2_outputs(601) <= (layer1_outputs(16)) or (layer1_outputs(936));
    layer2_outputs(602) <= layer1_outputs(2119);
    layer2_outputs(603) <= not(layer1_outputs(1047)) or (layer1_outputs(148));
    layer2_outputs(604) <= '1';
    layer2_outputs(605) <= layer1_outputs(1760);
    layer2_outputs(606) <= '0';
    layer2_outputs(607) <= layer1_outputs(1620);
    layer2_outputs(608) <= '1';
    layer2_outputs(609) <= not(layer1_outputs(2051));
    layer2_outputs(610) <= not(layer1_outputs(2440)) or (layer1_outputs(440));
    layer2_outputs(611) <= not(layer1_outputs(2312));
    layer2_outputs(612) <= not(layer1_outputs(1147)) or (layer1_outputs(215));
    layer2_outputs(613) <= (layer1_outputs(1528)) and (layer1_outputs(153));
    layer2_outputs(614) <= (layer1_outputs(378)) and not (layer1_outputs(1416));
    layer2_outputs(615) <= (layer1_outputs(1828)) xor (layer1_outputs(2015));
    layer2_outputs(616) <= not(layer1_outputs(482)) or (layer1_outputs(1637));
    layer2_outputs(617) <= '1';
    layer2_outputs(618) <= not(layer1_outputs(2108));
    layer2_outputs(619) <= not(layer1_outputs(2459));
    layer2_outputs(620) <= not(layer1_outputs(2185)) or (layer1_outputs(1529));
    layer2_outputs(621) <= not(layer1_outputs(2292));
    layer2_outputs(622) <= not(layer1_outputs(2520)) or (layer1_outputs(2098));
    layer2_outputs(623) <= '0';
    layer2_outputs(624) <= (layer1_outputs(984)) and not (layer1_outputs(2234));
    layer2_outputs(625) <= not(layer1_outputs(2114));
    layer2_outputs(626) <= (layer1_outputs(496)) xor (layer1_outputs(1551));
    layer2_outputs(627) <= not(layer1_outputs(103));
    layer2_outputs(628) <= '1';
    layer2_outputs(629) <= layer1_outputs(1231);
    layer2_outputs(630) <= not(layer1_outputs(1913)) or (layer1_outputs(1904));
    layer2_outputs(631) <= layer1_outputs(2316);
    layer2_outputs(632) <= layer1_outputs(2454);
    layer2_outputs(633) <= '1';
    layer2_outputs(634) <= not(layer1_outputs(2281)) or (layer1_outputs(1332));
    layer2_outputs(635) <= (layer1_outputs(405)) and not (layer1_outputs(2435));
    layer2_outputs(636) <= not((layer1_outputs(1180)) and (layer1_outputs(1944)));
    layer2_outputs(637) <= layer1_outputs(1207);
    layer2_outputs(638) <= (layer1_outputs(1793)) and not (layer1_outputs(77));
    layer2_outputs(639) <= not(layer1_outputs(356));
    layer2_outputs(640) <= '0';
    layer2_outputs(641) <= '1';
    layer2_outputs(642) <= '1';
    layer2_outputs(643) <= layer1_outputs(827);
    layer2_outputs(644) <= '1';
    layer2_outputs(645) <= not((layer1_outputs(28)) and (layer1_outputs(510)));
    layer2_outputs(646) <= (layer1_outputs(1974)) or (layer1_outputs(2198));
    layer2_outputs(647) <= not((layer1_outputs(2397)) and (layer1_outputs(2109)));
    layer2_outputs(648) <= not(layer1_outputs(879));
    layer2_outputs(649) <= layer1_outputs(1276);
    layer2_outputs(650) <= not((layer1_outputs(880)) and (layer1_outputs(468)));
    layer2_outputs(651) <= layer1_outputs(2359);
    layer2_outputs(652) <= not(layer1_outputs(111));
    layer2_outputs(653) <= not(layer1_outputs(1971));
    layer2_outputs(654) <= (layer1_outputs(2497)) and not (layer1_outputs(1010));
    layer2_outputs(655) <= (layer1_outputs(2277)) and (layer1_outputs(184));
    layer2_outputs(656) <= (layer1_outputs(1978)) and not (layer1_outputs(1094));
    layer2_outputs(657) <= not(layer1_outputs(177)) or (layer1_outputs(2265));
    layer2_outputs(658) <= layer1_outputs(2141);
    layer2_outputs(659) <= layer1_outputs(198);
    layer2_outputs(660) <= not((layer1_outputs(937)) and (layer1_outputs(1492)));
    layer2_outputs(661) <= not(layer1_outputs(217)) or (layer1_outputs(2366));
    layer2_outputs(662) <= not(layer1_outputs(544)) or (layer1_outputs(1317));
    layer2_outputs(663) <= not(layer1_outputs(558)) or (layer1_outputs(1520));
    layer2_outputs(664) <= '0';
    layer2_outputs(665) <= layer1_outputs(236);
    layer2_outputs(666) <= (layer1_outputs(2221)) and not (layer1_outputs(1878));
    layer2_outputs(667) <= layer1_outputs(1255);
    layer2_outputs(668) <= not((layer1_outputs(784)) and (layer1_outputs(1990)));
    layer2_outputs(669) <= not(layer1_outputs(1614));
    layer2_outputs(670) <= not(layer1_outputs(1656));
    layer2_outputs(671) <= (layer1_outputs(816)) and (layer1_outputs(734));
    layer2_outputs(672) <= not((layer1_outputs(185)) or (layer1_outputs(330)));
    layer2_outputs(673) <= not(layer1_outputs(1615));
    layer2_outputs(674) <= not((layer1_outputs(256)) and (layer1_outputs(1642)));
    layer2_outputs(675) <= not((layer1_outputs(2012)) or (layer1_outputs(1156)));
    layer2_outputs(676) <= (layer1_outputs(1770)) and not (layer1_outputs(1028));
    layer2_outputs(677) <= '0';
    layer2_outputs(678) <= '1';
    layer2_outputs(679) <= layer1_outputs(2077);
    layer2_outputs(680) <= not((layer1_outputs(1923)) or (layer1_outputs(2355)));
    layer2_outputs(681) <= layer1_outputs(931);
    layer2_outputs(682) <= (layer1_outputs(1301)) and not (layer1_outputs(2513));
    layer2_outputs(683) <= layer1_outputs(1794);
    layer2_outputs(684) <= '0';
    layer2_outputs(685) <= not((layer1_outputs(507)) and (layer1_outputs(806)));
    layer2_outputs(686) <= not(layer1_outputs(456));
    layer2_outputs(687) <= (layer1_outputs(1630)) or (layer1_outputs(1266));
    layer2_outputs(688) <= layer1_outputs(1877);
    layer2_outputs(689) <= layer1_outputs(1376);
    layer2_outputs(690) <= '0';
    layer2_outputs(691) <= (layer1_outputs(1605)) and not (layer1_outputs(90));
    layer2_outputs(692) <= (layer1_outputs(1428)) and (layer1_outputs(1832));
    layer2_outputs(693) <= not(layer1_outputs(2053));
    layer2_outputs(694) <= (layer1_outputs(255)) and (layer1_outputs(135));
    layer2_outputs(695) <= layer1_outputs(1494);
    layer2_outputs(696) <= not(layer1_outputs(2054));
    layer2_outputs(697) <= (layer1_outputs(1720)) and not (layer1_outputs(2288));
    layer2_outputs(698) <= not(layer1_outputs(1434));
    layer2_outputs(699) <= '0';
    layer2_outputs(700) <= not(layer1_outputs(563));
    layer2_outputs(701) <= not((layer1_outputs(542)) and (layer1_outputs(762)));
    layer2_outputs(702) <= '1';
    layer2_outputs(703) <= '1';
    layer2_outputs(704) <= not((layer1_outputs(892)) and (layer1_outputs(584)));
    layer2_outputs(705) <= layer1_outputs(1532);
    layer2_outputs(706) <= not(layer1_outputs(20));
    layer2_outputs(707) <= not(layer1_outputs(1905));
    layer2_outputs(708) <= not((layer1_outputs(1052)) or (layer1_outputs(2050)));
    layer2_outputs(709) <= layer1_outputs(2448);
    layer2_outputs(710) <= (layer1_outputs(1290)) and (layer1_outputs(464));
    layer2_outputs(711) <= not((layer1_outputs(695)) and (layer1_outputs(2203)));
    layer2_outputs(712) <= not(layer1_outputs(1163));
    layer2_outputs(713) <= '1';
    layer2_outputs(714) <= '0';
    layer2_outputs(715) <= not(layer1_outputs(1945));
    layer2_outputs(716) <= not(layer1_outputs(635)) or (layer1_outputs(1536));
    layer2_outputs(717) <= (layer1_outputs(1042)) or (layer1_outputs(1410));
    layer2_outputs(718) <= (layer1_outputs(501)) or (layer1_outputs(2406));
    layer2_outputs(719) <= (layer1_outputs(1987)) or (layer1_outputs(2530));
    layer2_outputs(720) <= not(layer1_outputs(1862));
    layer2_outputs(721) <= not((layer1_outputs(2132)) or (layer1_outputs(2178)));
    layer2_outputs(722) <= (layer1_outputs(1003)) and (layer1_outputs(1067));
    layer2_outputs(723) <= not(layer1_outputs(1541)) or (layer1_outputs(2553));
    layer2_outputs(724) <= (layer1_outputs(416)) and (layer1_outputs(2215));
    layer2_outputs(725) <= not(layer1_outputs(2509));
    layer2_outputs(726) <= not((layer1_outputs(2270)) and (layer1_outputs(1118)));
    layer2_outputs(727) <= (layer1_outputs(713)) and not (layer1_outputs(542));
    layer2_outputs(728) <= not((layer1_outputs(1629)) or (layer1_outputs(910)));
    layer2_outputs(729) <= not((layer1_outputs(2217)) or (layer1_outputs(1169)));
    layer2_outputs(730) <= (layer1_outputs(665)) and not (layer1_outputs(1172));
    layer2_outputs(731) <= (layer1_outputs(692)) and not (layer1_outputs(262));
    layer2_outputs(732) <= not(layer1_outputs(1514));
    layer2_outputs(733) <= not(layer1_outputs(788)) or (layer1_outputs(1429));
    layer2_outputs(734) <= (layer1_outputs(400)) and not (layer1_outputs(1580));
    layer2_outputs(735) <= '1';
    layer2_outputs(736) <= (layer1_outputs(2434)) or (layer1_outputs(2118));
    layer2_outputs(737) <= (layer1_outputs(1593)) and not (layer1_outputs(181));
    layer2_outputs(738) <= layer1_outputs(267);
    layer2_outputs(739) <= (layer1_outputs(1272)) or (layer1_outputs(772));
    layer2_outputs(740) <= not(layer1_outputs(2032));
    layer2_outputs(741) <= (layer1_outputs(928)) and (layer1_outputs(2091));
    layer2_outputs(742) <= not(layer1_outputs(45));
    layer2_outputs(743) <= layer1_outputs(1461);
    layer2_outputs(744) <= (layer1_outputs(1409)) and not (layer1_outputs(1215));
    layer2_outputs(745) <= '0';
    layer2_outputs(746) <= not(layer1_outputs(525));
    layer2_outputs(747) <= '0';
    layer2_outputs(748) <= not(layer1_outputs(2110));
    layer2_outputs(749) <= '0';
    layer2_outputs(750) <= '0';
    layer2_outputs(751) <= layer1_outputs(566);
    layer2_outputs(752) <= '1';
    layer2_outputs(753) <= not(layer1_outputs(1457)) or (layer1_outputs(2135));
    layer2_outputs(754) <= '0';
    layer2_outputs(755) <= (layer1_outputs(1071)) and not (layer1_outputs(576));
    layer2_outputs(756) <= not(layer1_outputs(829));
    layer2_outputs(757) <= layer1_outputs(1973);
    layer2_outputs(758) <= (layer1_outputs(1369)) and not (layer1_outputs(27));
    layer2_outputs(759) <= not((layer1_outputs(312)) or (layer1_outputs(1252)));
    layer2_outputs(760) <= (layer1_outputs(376)) and (layer1_outputs(152));
    layer2_outputs(761) <= (layer1_outputs(2464)) and not (layer1_outputs(1256));
    layer2_outputs(762) <= '0';
    layer2_outputs(763) <= (layer1_outputs(747)) and not (layer1_outputs(1625));
    layer2_outputs(764) <= layer1_outputs(958);
    layer2_outputs(765) <= '0';
    layer2_outputs(766) <= not(layer1_outputs(1609)) or (layer1_outputs(2155));
    layer2_outputs(767) <= '0';
    layer2_outputs(768) <= (layer1_outputs(2016)) and not (layer1_outputs(1029));
    layer2_outputs(769) <= (layer1_outputs(314)) xor (layer1_outputs(553));
    layer2_outputs(770) <= '1';
    layer2_outputs(771) <= not(layer1_outputs(755));
    layer2_outputs(772) <= layer1_outputs(834);
    layer2_outputs(773) <= layer1_outputs(77);
    layer2_outputs(774) <= not(layer1_outputs(3)) or (layer1_outputs(2500));
    layer2_outputs(775) <= (layer1_outputs(2182)) and not (layer1_outputs(2008));
    layer2_outputs(776) <= (layer1_outputs(845)) and not (layer1_outputs(61));
    layer2_outputs(777) <= (layer1_outputs(2392)) and not (layer1_outputs(1636));
    layer2_outputs(778) <= not((layer1_outputs(1387)) and (layer1_outputs(225)));
    layer2_outputs(779) <= layer1_outputs(1073);
    layer2_outputs(780) <= (layer1_outputs(2528)) and not (layer1_outputs(147));
    layer2_outputs(781) <= not(layer1_outputs(491)) or (layer1_outputs(2235));
    layer2_outputs(782) <= not(layer1_outputs(1058));
    layer2_outputs(783) <= not(layer1_outputs(1227)) or (layer1_outputs(727));
    layer2_outputs(784) <= not(layer1_outputs(2358));
    layer2_outputs(785) <= layer1_outputs(2341);
    layer2_outputs(786) <= '0';
    layer2_outputs(787) <= not(layer1_outputs(1353));
    layer2_outputs(788) <= layer1_outputs(549);
    layer2_outputs(789) <= (layer1_outputs(4)) and not (layer1_outputs(2489));
    layer2_outputs(790) <= not(layer1_outputs(58));
    layer2_outputs(791) <= (layer1_outputs(494)) and (layer1_outputs(317));
    layer2_outputs(792) <= not(layer1_outputs(26)) or (layer1_outputs(1888));
    layer2_outputs(793) <= layer1_outputs(1366);
    layer2_outputs(794) <= (layer1_outputs(789)) and (layer1_outputs(972));
    layer2_outputs(795) <= not(layer1_outputs(345)) or (layer1_outputs(1086));
    layer2_outputs(796) <= not(layer1_outputs(105));
    layer2_outputs(797) <= (layer1_outputs(19)) or (layer1_outputs(1791));
    layer2_outputs(798) <= '1';
    layer2_outputs(799) <= (layer1_outputs(1188)) or (layer1_outputs(1020));
    layer2_outputs(800) <= (layer1_outputs(1711)) and not (layer1_outputs(2362));
    layer2_outputs(801) <= (layer1_outputs(53)) or (layer1_outputs(1581));
    layer2_outputs(802) <= layer1_outputs(25);
    layer2_outputs(803) <= (layer1_outputs(1436)) and not (layer1_outputs(2395));
    layer2_outputs(804) <= not((layer1_outputs(892)) and (layer1_outputs(1388)));
    layer2_outputs(805) <= (layer1_outputs(672)) or (layer1_outputs(648));
    layer2_outputs(806) <= (layer1_outputs(2201)) and not (layer1_outputs(2246));
    layer2_outputs(807) <= layer1_outputs(2075);
    layer2_outputs(808) <= (layer1_outputs(922)) or (layer1_outputs(2168));
    layer2_outputs(809) <= not(layer1_outputs(824)) or (layer1_outputs(703));
    layer2_outputs(810) <= not((layer1_outputs(1018)) or (layer1_outputs(2050)));
    layer2_outputs(811) <= '1';
    layer2_outputs(812) <= (layer1_outputs(624)) and not (layer1_outputs(1583));
    layer2_outputs(813) <= not((layer1_outputs(1800)) and (layer1_outputs(473)));
    layer2_outputs(814) <= (layer1_outputs(2522)) or (layer1_outputs(1642));
    layer2_outputs(815) <= (layer1_outputs(1895)) or (layer1_outputs(1757));
    layer2_outputs(816) <= not(layer1_outputs(59)) or (layer1_outputs(1769));
    layer2_outputs(817) <= '0';
    layer2_outputs(818) <= layer1_outputs(65);
    layer2_outputs(819) <= not((layer1_outputs(1532)) xor (layer1_outputs(1930)));
    layer2_outputs(820) <= '1';
    layer2_outputs(821) <= (layer1_outputs(1178)) or (layer1_outputs(799));
    layer2_outputs(822) <= not(layer1_outputs(1167));
    layer2_outputs(823) <= '1';
    layer2_outputs(824) <= not((layer1_outputs(1375)) or (layer1_outputs(1690)));
    layer2_outputs(825) <= not(layer1_outputs(2551));
    layer2_outputs(826) <= '0';
    layer2_outputs(827) <= (layer1_outputs(432)) and (layer1_outputs(2023));
    layer2_outputs(828) <= (layer1_outputs(261)) and not (layer1_outputs(292));
    layer2_outputs(829) <= (layer1_outputs(1196)) and not (layer1_outputs(1350));
    layer2_outputs(830) <= layer1_outputs(1316);
    layer2_outputs(831) <= layer1_outputs(1042);
    layer2_outputs(832) <= layer1_outputs(808);
    layer2_outputs(833) <= (layer1_outputs(2054)) and not (layer1_outputs(1566));
    layer2_outputs(834) <= layer1_outputs(1283);
    layer2_outputs(835) <= (layer1_outputs(219)) or (layer1_outputs(404));
    layer2_outputs(836) <= '1';
    layer2_outputs(837) <= not((layer1_outputs(180)) and (layer1_outputs(47)));
    layer2_outputs(838) <= not(layer1_outputs(2497));
    layer2_outputs(839) <= '1';
    layer2_outputs(840) <= (layer1_outputs(2057)) and not (layer1_outputs(1336));
    layer2_outputs(841) <= layer1_outputs(764);
    layer2_outputs(842) <= not(layer1_outputs(112));
    layer2_outputs(843) <= '0';
    layer2_outputs(844) <= '1';
    layer2_outputs(845) <= (layer1_outputs(1279)) or (layer1_outputs(733));
    layer2_outputs(846) <= not(layer1_outputs(2074));
    layer2_outputs(847) <= layer1_outputs(1386);
    layer2_outputs(848) <= layer1_outputs(333);
    layer2_outputs(849) <= (layer1_outputs(966)) and not (layer1_outputs(1007));
    layer2_outputs(850) <= not((layer1_outputs(835)) or (layer1_outputs(2048)));
    layer2_outputs(851) <= not(layer1_outputs(2177)) or (layer1_outputs(1175));
    layer2_outputs(852) <= (layer1_outputs(617)) and (layer1_outputs(583));
    layer2_outputs(853) <= not(layer1_outputs(934)) or (layer1_outputs(2228));
    layer2_outputs(854) <= (layer1_outputs(1638)) and (layer1_outputs(76));
    layer2_outputs(855) <= not(layer1_outputs(1195)) or (layer1_outputs(780));
    layer2_outputs(856) <= not(layer1_outputs(1654));
    layer2_outputs(857) <= '0';
    layer2_outputs(858) <= layer1_outputs(266);
    layer2_outputs(859) <= '1';
    layer2_outputs(860) <= (layer1_outputs(1448)) xor (layer1_outputs(2330));
    layer2_outputs(861) <= '0';
    layer2_outputs(862) <= layer1_outputs(784);
    layer2_outputs(863) <= not(layer1_outputs(1966));
    layer2_outputs(864) <= (layer1_outputs(1501)) and (layer1_outputs(1516));
    layer2_outputs(865) <= not(layer1_outputs(1069)) or (layer1_outputs(18));
    layer2_outputs(866) <= (layer1_outputs(2034)) or (layer1_outputs(2187));
    layer2_outputs(867) <= '0';
    layer2_outputs(868) <= not((layer1_outputs(54)) or (layer1_outputs(1093)));
    layer2_outputs(869) <= '0';
    layer2_outputs(870) <= '1';
    layer2_outputs(871) <= not(layer1_outputs(431)) or (layer1_outputs(1746));
    layer2_outputs(872) <= not(layer1_outputs(29));
    layer2_outputs(873) <= not((layer1_outputs(2185)) and (layer1_outputs(30)));
    layer2_outputs(874) <= '0';
    layer2_outputs(875) <= layer1_outputs(1031);
    layer2_outputs(876) <= '0';
    layer2_outputs(877) <= not(layer1_outputs(1037));
    layer2_outputs(878) <= '0';
    layer2_outputs(879) <= (layer1_outputs(1475)) xor (layer1_outputs(1105));
    layer2_outputs(880) <= not(layer1_outputs(1187));
    layer2_outputs(881) <= (layer1_outputs(2063)) or (layer1_outputs(2138));
    layer2_outputs(882) <= not(layer1_outputs(521));
    layer2_outputs(883) <= layer1_outputs(2038);
    layer2_outputs(884) <= (layer1_outputs(1088)) and not (layer1_outputs(2356));
    layer2_outputs(885) <= not(layer1_outputs(355));
    layer2_outputs(886) <= '1';
    layer2_outputs(887) <= not((layer1_outputs(227)) or (layer1_outputs(1956)));
    layer2_outputs(888) <= not(layer1_outputs(2388)) or (layer1_outputs(1404));
    layer2_outputs(889) <= not(layer1_outputs(1500));
    layer2_outputs(890) <= (layer1_outputs(2143)) and not (layer1_outputs(1067));
    layer2_outputs(891) <= layer1_outputs(1672);
    layer2_outputs(892) <= not((layer1_outputs(1044)) or (layer1_outputs(1841)));
    layer2_outputs(893) <= '0';
    layer2_outputs(894) <= not((layer1_outputs(915)) or (layer1_outputs(1994)));
    layer2_outputs(895) <= (layer1_outputs(2444)) and (layer1_outputs(2492));
    layer2_outputs(896) <= not(layer1_outputs(928));
    layer2_outputs(897) <= not((layer1_outputs(799)) and (layer1_outputs(2460)));
    layer2_outputs(898) <= layer1_outputs(2511);
    layer2_outputs(899) <= layer1_outputs(2096);
    layer2_outputs(900) <= layer1_outputs(1175);
    layer2_outputs(901) <= not(layer1_outputs(1658)) or (layer1_outputs(1551));
    layer2_outputs(902) <= not(layer1_outputs(960));
    layer2_outputs(903) <= not(layer1_outputs(188));
    layer2_outputs(904) <= layer1_outputs(656);
    layer2_outputs(905) <= (layer1_outputs(1792)) and (layer1_outputs(1486));
    layer2_outputs(906) <= not((layer1_outputs(1097)) or (layer1_outputs(1508)));
    layer2_outputs(907) <= not((layer1_outputs(1214)) and (layer1_outputs(139)));
    layer2_outputs(908) <= not(layer1_outputs(1504)) or (layer1_outputs(536));
    layer2_outputs(909) <= (layer1_outputs(233)) or (layer1_outputs(1695));
    layer2_outputs(910) <= not(layer1_outputs(359));
    layer2_outputs(911) <= layer1_outputs(625);
    layer2_outputs(912) <= '0';
    layer2_outputs(913) <= layer1_outputs(212);
    layer2_outputs(914) <= '0';
    layer2_outputs(915) <= '0';
    layer2_outputs(916) <= (layer1_outputs(584)) and (layer1_outputs(363));
    layer2_outputs(917) <= not((layer1_outputs(255)) and (layer1_outputs(1950)));
    layer2_outputs(918) <= not((layer1_outputs(2089)) and (layer1_outputs(1010)));
    layer2_outputs(919) <= layer1_outputs(1354);
    layer2_outputs(920) <= not(layer1_outputs(808));
    layer2_outputs(921) <= layer1_outputs(2431);
    layer2_outputs(922) <= (layer1_outputs(460)) and not (layer1_outputs(1217));
    layer2_outputs(923) <= not(layer1_outputs(1362));
    layer2_outputs(924) <= (layer1_outputs(557)) and not (layer1_outputs(1306));
    layer2_outputs(925) <= not((layer1_outputs(366)) or (layer1_outputs(1452)));
    layer2_outputs(926) <= layer1_outputs(1665);
    layer2_outputs(927) <= (layer1_outputs(374)) or (layer1_outputs(1317));
    layer2_outputs(928) <= '1';
    layer2_outputs(929) <= (layer1_outputs(119)) or (layer1_outputs(2367));
    layer2_outputs(930) <= (layer1_outputs(2051)) and not (layer1_outputs(200));
    layer2_outputs(931) <= (layer1_outputs(2260)) and not (layer1_outputs(1697));
    layer2_outputs(932) <= (layer1_outputs(1237)) or (layer1_outputs(708));
    layer2_outputs(933) <= (layer1_outputs(2103)) and not (layer1_outputs(1507));
    layer2_outputs(934) <= not(layer1_outputs(804));
    layer2_outputs(935) <= (layer1_outputs(530)) and not (layer1_outputs(1619));
    layer2_outputs(936) <= not(layer1_outputs(1833)) or (layer1_outputs(527));
    layer2_outputs(937) <= not((layer1_outputs(53)) and (layer1_outputs(209)));
    layer2_outputs(938) <= not(layer1_outputs(387));
    layer2_outputs(939) <= (layer1_outputs(2381)) and (layer1_outputs(517));
    layer2_outputs(940) <= '0';
    layer2_outputs(941) <= (layer1_outputs(1602)) and not (layer1_outputs(1702));
    layer2_outputs(942) <= not((layer1_outputs(2328)) and (layer1_outputs(485)));
    layer2_outputs(943) <= not((layer1_outputs(2358)) and (layer1_outputs(555)));
    layer2_outputs(944) <= '0';
    layer2_outputs(945) <= layer1_outputs(1371);
    layer2_outputs(946) <= not((layer1_outputs(550)) or (layer1_outputs(2533)));
    layer2_outputs(947) <= (layer1_outputs(383)) and not (layer1_outputs(1349));
    layer2_outputs(948) <= '1';
    layer2_outputs(949) <= (layer1_outputs(711)) and not (layer1_outputs(2411));
    layer2_outputs(950) <= not(layer1_outputs(422));
    layer2_outputs(951) <= not(layer1_outputs(2154));
    layer2_outputs(952) <= (layer1_outputs(583)) and not (layer1_outputs(946));
    layer2_outputs(953) <= not(layer1_outputs(1489)) or (layer1_outputs(1682));
    layer2_outputs(954) <= not((layer1_outputs(501)) or (layer1_outputs(2306)));
    layer2_outputs(955) <= not(layer1_outputs(608));
    layer2_outputs(956) <= (layer1_outputs(753)) and not (layer1_outputs(309));
    layer2_outputs(957) <= layer1_outputs(287);
    layer2_outputs(958) <= not(layer1_outputs(794)) or (layer1_outputs(1233));
    layer2_outputs(959) <= not(layer1_outputs(1053)) or (layer1_outputs(2100));
    layer2_outputs(960) <= '0';
    layer2_outputs(961) <= '0';
    layer2_outputs(962) <= not(layer1_outputs(261));
    layer2_outputs(963) <= layer1_outputs(2320);
    layer2_outputs(964) <= (layer1_outputs(1349)) or (layer1_outputs(2415));
    layer2_outputs(965) <= (layer1_outputs(2)) or (layer1_outputs(1893));
    layer2_outputs(966) <= layer1_outputs(859);
    layer2_outputs(967) <= layer1_outputs(386);
    layer2_outputs(968) <= layer1_outputs(1574);
    layer2_outputs(969) <= '0';
    layer2_outputs(970) <= not(layer1_outputs(2285));
    layer2_outputs(971) <= (layer1_outputs(2495)) or (layer1_outputs(672));
    layer2_outputs(972) <= (layer1_outputs(2465)) and not (layer1_outputs(1470));
    layer2_outputs(973) <= not(layer1_outputs(122));
    layer2_outputs(974) <= (layer1_outputs(1135)) and not (layer1_outputs(354));
    layer2_outputs(975) <= layer1_outputs(1771);
    layer2_outputs(976) <= layer1_outputs(268);
    layer2_outputs(977) <= not(layer1_outputs(2299));
    layer2_outputs(978) <= not(layer1_outputs(1094)) or (layer1_outputs(1447));
    layer2_outputs(979) <= (layer1_outputs(2274)) and (layer1_outputs(627));
    layer2_outputs(980) <= layer1_outputs(2482);
    layer2_outputs(981) <= not(layer1_outputs(2044));
    layer2_outputs(982) <= (layer1_outputs(412)) and not (layer1_outputs(1123));
    layer2_outputs(983) <= (layer1_outputs(1299)) and not (layer1_outputs(919));
    layer2_outputs(984) <= not((layer1_outputs(1120)) and (layer1_outputs(226)));
    layer2_outputs(985) <= not((layer1_outputs(1894)) or (layer1_outputs(1892)));
    layer2_outputs(986) <= layer1_outputs(455);
    layer2_outputs(987) <= '1';
    layer2_outputs(988) <= (layer1_outputs(1373)) and not (layer1_outputs(1853));
    layer2_outputs(989) <= layer1_outputs(1118);
    layer2_outputs(990) <= '0';
    layer2_outputs(991) <= layer1_outputs(1630);
    layer2_outputs(992) <= (layer1_outputs(662)) or (layer1_outputs(986));
    layer2_outputs(993) <= not(layer1_outputs(590)) or (layer1_outputs(2393));
    layer2_outputs(994) <= not(layer1_outputs(1558)) or (layer1_outputs(1079));
    layer2_outputs(995) <= (layer1_outputs(133)) or (layer1_outputs(1799));
    layer2_outputs(996) <= layer1_outputs(1355);
    layer2_outputs(997) <= '1';
    layer2_outputs(998) <= (layer1_outputs(2277)) and not (layer1_outputs(13));
    layer2_outputs(999) <= (layer1_outputs(1850)) or (layer1_outputs(193));
    layer2_outputs(1000) <= (layer1_outputs(1226)) and (layer1_outputs(1960));
    layer2_outputs(1001) <= (layer1_outputs(812)) and (layer1_outputs(680));
    layer2_outputs(1002) <= not((layer1_outputs(955)) and (layer1_outputs(354)));
    layer2_outputs(1003) <= (layer1_outputs(1783)) and not (layer1_outputs(1291));
    layer2_outputs(1004) <= '1';
    layer2_outputs(1005) <= not(layer1_outputs(2326));
    layer2_outputs(1006) <= (layer1_outputs(438)) and (layer1_outputs(535));
    layer2_outputs(1007) <= '0';
    layer2_outputs(1008) <= (layer1_outputs(995)) and not (layer1_outputs(267));
    layer2_outputs(1009) <= '0';
    layer2_outputs(1010) <= not(layer1_outputs(2253)) or (layer1_outputs(1140));
    layer2_outputs(1011) <= layer1_outputs(2002);
    layer2_outputs(1012) <= (layer1_outputs(2068)) or (layer1_outputs(428));
    layer2_outputs(1013) <= not(layer1_outputs(2184));
    layer2_outputs(1014) <= layer1_outputs(1304);
    layer2_outputs(1015) <= not(layer1_outputs(942));
    layer2_outputs(1016) <= (layer1_outputs(101)) or (layer1_outputs(909));
    layer2_outputs(1017) <= not(layer1_outputs(472)) or (layer1_outputs(1432));
    layer2_outputs(1018) <= layer1_outputs(1643);
    layer2_outputs(1019) <= (layer1_outputs(8)) xor (layer1_outputs(15));
    layer2_outputs(1020) <= layer1_outputs(395);
    layer2_outputs(1021) <= layer1_outputs(1930);
    layer2_outputs(1022) <= (layer1_outputs(1006)) and not (layer1_outputs(734));
    layer2_outputs(1023) <= '1';
    layer2_outputs(1024) <= not((layer1_outputs(94)) xor (layer1_outputs(776)));
    layer2_outputs(1025) <= not(layer1_outputs(2474));
    layer2_outputs(1026) <= not(layer1_outputs(2025)) or (layer1_outputs(2085));
    layer2_outputs(1027) <= not(layer1_outputs(689)) or (layer1_outputs(1622));
    layer2_outputs(1028) <= layer1_outputs(242);
    layer2_outputs(1029) <= (layer1_outputs(1568)) or (layer1_outputs(815));
    layer2_outputs(1030) <= '0';
    layer2_outputs(1031) <= not((layer1_outputs(1096)) and (layer1_outputs(964)));
    layer2_outputs(1032) <= (layer1_outputs(1217)) and (layer1_outputs(502));
    layer2_outputs(1033) <= not(layer1_outputs(598)) or (layer1_outputs(1498));
    layer2_outputs(1034) <= layer1_outputs(1624);
    layer2_outputs(1035) <= '0';
    layer2_outputs(1036) <= '0';
    layer2_outputs(1037) <= '0';
    layer2_outputs(1038) <= '1';
    layer2_outputs(1039) <= not(layer1_outputs(2042)) or (layer1_outputs(1434));
    layer2_outputs(1040) <= not(layer1_outputs(633));
    layer2_outputs(1041) <= not((layer1_outputs(1917)) or (layer1_outputs(1539)));
    layer2_outputs(1042) <= (layer1_outputs(1707)) xor (layer1_outputs(868));
    layer2_outputs(1043) <= not((layer1_outputs(1904)) or (layer1_outputs(996)));
    layer2_outputs(1044) <= not((layer1_outputs(1948)) xor (layer1_outputs(1851)));
    layer2_outputs(1045) <= not(layer1_outputs(128)) or (layer1_outputs(1101));
    layer2_outputs(1046) <= (layer1_outputs(1994)) and (layer1_outputs(1823));
    layer2_outputs(1047) <= (layer1_outputs(1225)) and (layer1_outputs(1251));
    layer2_outputs(1048) <= not(layer1_outputs(2104)) or (layer1_outputs(2117));
    layer2_outputs(1049) <= '1';
    layer2_outputs(1050) <= not(layer1_outputs(2429));
    layer2_outputs(1051) <= (layer1_outputs(556)) and not (layer1_outputs(778));
    layer2_outputs(1052) <= (layer1_outputs(258)) and not (layer1_outputs(351));
    layer2_outputs(1053) <= '1';
    layer2_outputs(1054) <= layer1_outputs(1403);
    layer2_outputs(1055) <= not(layer1_outputs(1034)) or (layer1_outputs(2055));
    layer2_outputs(1056) <= not((layer1_outputs(938)) and (layer1_outputs(1951)));
    layer2_outputs(1057) <= not(layer1_outputs(1913)) or (layer1_outputs(1781));
    layer2_outputs(1058) <= layer1_outputs(914);
    layer2_outputs(1059) <= (layer1_outputs(2025)) or (layer1_outputs(1734));
    layer2_outputs(1060) <= '0';
    layer2_outputs(1061) <= (layer1_outputs(426)) and not (layer1_outputs(723));
    layer2_outputs(1062) <= (layer1_outputs(1499)) or (layer1_outputs(1594));
    layer2_outputs(1063) <= not(layer1_outputs(783)) or (layer1_outputs(2539));
    layer2_outputs(1064) <= not(layer1_outputs(578)) or (layer1_outputs(600));
    layer2_outputs(1065) <= not(layer1_outputs(1499)) or (layer1_outputs(5));
    layer2_outputs(1066) <= layer1_outputs(1742);
    layer2_outputs(1067) <= (layer1_outputs(607)) and (layer1_outputs(2247));
    layer2_outputs(1068) <= not(layer1_outputs(2323));
    layer2_outputs(1069) <= not(layer1_outputs(1048)) or (layer1_outputs(508));
    layer2_outputs(1070) <= not(layer1_outputs(1818));
    layer2_outputs(1071) <= not(layer1_outputs(229));
    layer2_outputs(1072) <= layer1_outputs(1315);
    layer2_outputs(1073) <= (layer1_outputs(1582)) and not (layer1_outputs(2443));
    layer2_outputs(1074) <= '1';
    layer2_outputs(1075) <= (layer1_outputs(2478)) or (layer1_outputs(795));
    layer2_outputs(1076) <= not(layer1_outputs(1704));
    layer2_outputs(1077) <= not((layer1_outputs(1907)) or (layer1_outputs(2085)));
    layer2_outputs(1078) <= (layer1_outputs(781)) or (layer1_outputs(2270));
    layer2_outputs(1079) <= not((layer1_outputs(980)) or (layer1_outputs(2224)));
    layer2_outputs(1080) <= (layer1_outputs(447)) and not (layer1_outputs(720));
    layer2_outputs(1081) <= '1';
    layer2_outputs(1082) <= '0';
    layer2_outputs(1083) <= (layer1_outputs(112)) and not (layer1_outputs(1523));
    layer2_outputs(1084) <= (layer1_outputs(115)) and (layer1_outputs(187));
    layer2_outputs(1085) <= (layer1_outputs(1569)) or (layer1_outputs(1189));
    layer2_outputs(1086) <= (layer1_outputs(895)) and not (layer1_outputs(1408));
    layer2_outputs(1087) <= (layer1_outputs(1810)) and not (layer1_outputs(1813));
    layer2_outputs(1088) <= not(layer1_outputs(599));
    layer2_outputs(1089) <= '0';
    layer2_outputs(1090) <= '0';
    layer2_outputs(1091) <= '0';
    layer2_outputs(1092) <= layer1_outputs(748);
    layer2_outputs(1093) <= not(layer1_outputs(1580));
    layer2_outputs(1094) <= not(layer1_outputs(458));
    layer2_outputs(1095) <= not((layer1_outputs(1893)) and (layer1_outputs(1277)));
    layer2_outputs(1096) <= (layer1_outputs(1181)) or (layer1_outputs(793));
    layer2_outputs(1097) <= not(layer1_outputs(151));
    layer2_outputs(1098) <= not((layer1_outputs(1189)) or (layer1_outputs(2106)));
    layer2_outputs(1099) <= layer1_outputs(2510);
    layer2_outputs(1100) <= (layer1_outputs(585)) and (layer1_outputs(11));
    layer2_outputs(1101) <= '1';
    layer2_outputs(1102) <= (layer1_outputs(1543)) or (layer1_outputs(2501));
    layer2_outputs(1103) <= (layer1_outputs(44)) and (layer1_outputs(769));
    layer2_outputs(1104) <= layer1_outputs(2491);
    layer2_outputs(1105) <= not(layer1_outputs(704));
    layer2_outputs(1106) <= not(layer1_outputs(2130)) or (layer1_outputs(1441));
    layer2_outputs(1107) <= layer1_outputs(353);
    layer2_outputs(1108) <= (layer1_outputs(2100)) and (layer1_outputs(1931));
    layer2_outputs(1109) <= layer1_outputs(1559);
    layer2_outputs(1110) <= (layer1_outputs(2180)) and not (layer1_outputs(2280));
    layer2_outputs(1111) <= not(layer1_outputs(802));
    layer2_outputs(1112) <= not(layer1_outputs(516));
    layer2_outputs(1113) <= (layer1_outputs(73)) or (layer1_outputs(280));
    layer2_outputs(1114) <= '0';
    layer2_outputs(1115) <= (layer1_outputs(1357)) and not (layer1_outputs(117));
    layer2_outputs(1116) <= not(layer1_outputs(2390)) or (layer1_outputs(1661));
    layer2_outputs(1117) <= '0';
    layer2_outputs(1118) <= not(layer1_outputs(1198)) or (layer1_outputs(408));
    layer2_outputs(1119) <= '0';
    layer2_outputs(1120) <= '1';
    layer2_outputs(1121) <= not((layer1_outputs(698)) and (layer1_outputs(1288)));
    layer2_outputs(1122) <= not((layer1_outputs(2029)) and (layer1_outputs(1197)));
    layer2_outputs(1123) <= (layer1_outputs(1002)) and (layer1_outputs(305));
    layer2_outputs(1124) <= not(layer1_outputs(222));
    layer2_outputs(1125) <= layer1_outputs(658);
    layer2_outputs(1126) <= '1';
    layer2_outputs(1127) <= layer1_outputs(943);
    layer2_outputs(1128) <= not((layer1_outputs(98)) or (layer1_outputs(49)));
    layer2_outputs(1129) <= (layer1_outputs(1699)) and not (layer1_outputs(1108));
    layer2_outputs(1130) <= '0';
    layer2_outputs(1131) <= not(layer1_outputs(565));
    layer2_outputs(1132) <= not(layer1_outputs(2327)) or (layer1_outputs(663));
    layer2_outputs(1133) <= not((layer1_outputs(554)) and (layer1_outputs(380)));
    layer2_outputs(1134) <= layer1_outputs(205);
    layer2_outputs(1135) <= (layer1_outputs(935)) and (layer1_outputs(64));
    layer2_outputs(1136) <= not(layer1_outputs(1204));
    layer2_outputs(1137) <= layer1_outputs(134);
    layer2_outputs(1138) <= '1';
    layer2_outputs(1139) <= not(layer1_outputs(2231));
    layer2_outputs(1140) <= (layer1_outputs(177)) or (layer1_outputs(1758));
    layer2_outputs(1141) <= not(layer1_outputs(121));
    layer2_outputs(1142) <= not(layer1_outputs(1422));
    layer2_outputs(1143) <= not(layer1_outputs(522)) or (layer1_outputs(189));
    layer2_outputs(1144) <= not(layer1_outputs(689));
    layer2_outputs(1145) <= (layer1_outputs(1473)) and (layer1_outputs(445));
    layer2_outputs(1146) <= '1';
    layer2_outputs(1147) <= (layer1_outputs(370)) and (layer1_outputs(631));
    layer2_outputs(1148) <= (layer1_outputs(2470)) and not (layer1_outputs(1989));
    layer2_outputs(1149) <= (layer1_outputs(2437)) and not (layer1_outputs(2348));
    layer2_outputs(1150) <= '0';
    layer2_outputs(1151) <= '1';
    layer2_outputs(1152) <= (layer1_outputs(352)) and not (layer1_outputs(1716));
    layer2_outputs(1153) <= not((layer1_outputs(2049)) and (layer1_outputs(1628)));
    layer2_outputs(1154) <= layer1_outputs(2362);
    layer2_outputs(1155) <= not(layer1_outputs(190)) or (layer1_outputs(1110));
    layer2_outputs(1156) <= layer1_outputs(2049);
    layer2_outputs(1157) <= (layer1_outputs(2445)) and not (layer1_outputs(1799));
    layer2_outputs(1158) <= not((layer1_outputs(1599)) or (layer1_outputs(331)));
    layer2_outputs(1159) <= '1';
    layer2_outputs(1160) <= (layer1_outputs(205)) and not (layer1_outputs(1328));
    layer2_outputs(1161) <= layer1_outputs(1009);
    layer2_outputs(1162) <= not(layer1_outputs(2204));
    layer2_outputs(1163) <= not(layer1_outputs(1752));
    layer2_outputs(1164) <= layer1_outputs(927);
    layer2_outputs(1165) <= (layer1_outputs(2069)) and not (layer1_outputs(1808));
    layer2_outputs(1166) <= not(layer1_outputs(344));
    layer2_outputs(1167) <= not((layer1_outputs(31)) and (layer1_outputs(840)));
    layer2_outputs(1168) <= (layer1_outputs(1753)) and not (layer1_outputs(40));
    layer2_outputs(1169) <= (layer1_outputs(1382)) and not (layer1_outputs(1993));
    layer2_outputs(1170) <= not(layer1_outputs(573));
    layer2_outputs(1171) <= (layer1_outputs(2010)) and (layer1_outputs(1037));
    layer2_outputs(1172) <= not(layer1_outputs(276));
    layer2_outputs(1173) <= not(layer1_outputs(1073)) or (layer1_outputs(1517));
    layer2_outputs(1174) <= not(layer1_outputs(2468)) or (layer1_outputs(740));
    layer2_outputs(1175) <= layer1_outputs(1415);
    layer2_outputs(1176) <= (layer1_outputs(1459)) or (layer1_outputs(379));
    layer2_outputs(1177) <= layer1_outputs(2333);
    layer2_outputs(1178) <= layer1_outputs(1912);
    layer2_outputs(1179) <= '1';
    layer2_outputs(1180) <= not(layer1_outputs(284));
    layer2_outputs(1181) <= not(layer1_outputs(1954)) or (layer1_outputs(107));
    layer2_outputs(1182) <= not((layer1_outputs(276)) and (layer1_outputs(994)));
    layer2_outputs(1183) <= layer1_outputs(466);
    layer2_outputs(1184) <= layer1_outputs(779);
    layer2_outputs(1185) <= '1';
    layer2_outputs(1186) <= (layer1_outputs(32)) and not (layer1_outputs(2028));
    layer2_outputs(1187) <= (layer1_outputs(1385)) and not (layer1_outputs(1040));
    layer2_outputs(1188) <= layer1_outputs(667);
    layer2_outputs(1189) <= (layer1_outputs(1892)) or (layer1_outputs(1330));
    layer2_outputs(1190) <= layer1_outputs(1652);
    layer2_outputs(1191) <= layer1_outputs(1096);
    layer2_outputs(1192) <= not((layer1_outputs(1004)) or (layer1_outputs(1243)));
    layer2_outputs(1193) <= '1';
    layer2_outputs(1194) <= '0';
    layer2_outputs(1195) <= (layer1_outputs(12)) or (layer1_outputs(456));
    layer2_outputs(1196) <= layer1_outputs(1977);
    layer2_outputs(1197) <= '1';
    layer2_outputs(1198) <= not(layer1_outputs(2324)) or (layer1_outputs(1312));
    layer2_outputs(1199) <= layer1_outputs(1134);
    layer2_outputs(1200) <= not((layer1_outputs(155)) or (layer1_outputs(1490)));
    layer2_outputs(1201) <= '1';
    layer2_outputs(1202) <= not((layer1_outputs(379)) and (layer1_outputs(59)));
    layer2_outputs(1203) <= not(layer1_outputs(178)) or (layer1_outputs(2134));
    layer2_outputs(1204) <= (layer1_outputs(1377)) and not (layer1_outputs(46));
    layer2_outputs(1205) <= not(layer1_outputs(630)) or (layer1_outputs(1607));
    layer2_outputs(1206) <= '0';
    layer2_outputs(1207) <= '1';
    layer2_outputs(1208) <= '0';
    layer2_outputs(1209) <= not((layer1_outputs(1666)) and (layer1_outputs(2230)));
    layer2_outputs(1210) <= (layer1_outputs(598)) or (layer1_outputs(1424));
    layer2_outputs(1211) <= (layer1_outputs(2150)) and not (layer1_outputs(896));
    layer2_outputs(1212) <= (layer1_outputs(410)) and not (layer1_outputs(1767));
    layer2_outputs(1213) <= '1';
    layer2_outputs(1214) <= '0';
    layer2_outputs(1215) <= (layer1_outputs(1827)) and (layer1_outputs(2183));
    layer2_outputs(1216) <= layer1_outputs(1542);
    layer2_outputs(1217) <= '1';
    layer2_outputs(1218) <= '0';
    layer2_outputs(1219) <= not(layer1_outputs(1546));
    layer2_outputs(1220) <= not(layer1_outputs(1325));
    layer2_outputs(1221) <= (layer1_outputs(2283)) and not (layer1_outputs(792));
    layer2_outputs(1222) <= (layer1_outputs(1897)) and not (layer1_outputs(853));
    layer2_outputs(1223) <= '0';
    layer2_outputs(1224) <= (layer1_outputs(956)) and not (layer1_outputs(23));
    layer2_outputs(1225) <= '1';
    layer2_outputs(1226) <= not((layer1_outputs(785)) or (layer1_outputs(2551)));
    layer2_outputs(1227) <= '1';
    layer2_outputs(1228) <= (layer1_outputs(1559)) xor (layer1_outputs(2527));
    layer2_outputs(1229) <= layer1_outputs(2534);
    layer2_outputs(1230) <= not(layer1_outputs(1506));
    layer2_outputs(1231) <= '0';
    layer2_outputs(1232) <= '1';
    layer2_outputs(1233) <= (layer1_outputs(1855)) and (layer1_outputs(635));
    layer2_outputs(1234) <= '1';
    layer2_outputs(1235) <= not((layer1_outputs(1847)) and (layer1_outputs(412)));
    layer2_outputs(1236) <= not(layer1_outputs(2342)) or (layer1_outputs(514));
    layer2_outputs(1237) <= '1';
    layer2_outputs(1238) <= layer1_outputs(1305);
    layer2_outputs(1239) <= (layer1_outputs(653)) and not (layer1_outputs(1337));
    layer2_outputs(1240) <= layer1_outputs(192);
    layer2_outputs(1241) <= '0';
    layer2_outputs(1242) <= '1';
    layer2_outputs(1243) <= not((layer1_outputs(739)) or (layer1_outputs(1692)));
    layer2_outputs(1244) <= (layer1_outputs(2545)) and not (layer1_outputs(768));
    layer2_outputs(1245) <= (layer1_outputs(2415)) and not (layer1_outputs(1157));
    layer2_outputs(1246) <= '1';
    layer2_outputs(1247) <= (layer1_outputs(1050)) and (layer1_outputs(301));
    layer2_outputs(1248) <= '1';
    layer2_outputs(1249) <= not(layer1_outputs(729)) or (layer1_outputs(629));
    layer2_outputs(1250) <= layer1_outputs(864);
    layer2_outputs(1251) <= not(layer1_outputs(1619));
    layer2_outputs(1252) <= layer1_outputs(142);
    layer2_outputs(1253) <= not((layer1_outputs(1952)) or (layer1_outputs(410)));
    layer2_outputs(1254) <= not(layer1_outputs(897)) or (layer1_outputs(1257));
    layer2_outputs(1255) <= (layer1_outputs(2044)) and not (layer1_outputs(1211));
    layer2_outputs(1256) <= '0';
    layer2_outputs(1257) <= not(layer1_outputs(1246));
    layer2_outputs(1258) <= layer1_outputs(1885);
    layer2_outputs(1259) <= '1';
    layer2_outputs(1260) <= not(layer1_outputs(2236)) or (layer1_outputs(1341));
    layer2_outputs(1261) <= not(layer1_outputs(2017)) or (layer1_outputs(2073));
    layer2_outputs(1262) <= not((layer1_outputs(1730)) or (layer1_outputs(1124)));
    layer2_outputs(1263) <= '0';
    layer2_outputs(1264) <= (layer1_outputs(300)) and (layer1_outputs(1286));
    layer2_outputs(1265) <= '1';
    layer2_outputs(1266) <= layer1_outputs(1293);
    layer2_outputs(1267) <= not(layer1_outputs(2449)) or (layer1_outputs(137));
    layer2_outputs(1268) <= not(layer1_outputs(2030));
    layer2_outputs(1269) <= not(layer1_outputs(448)) or (layer1_outputs(2208));
    layer2_outputs(1270) <= not((layer1_outputs(2373)) and (layer1_outputs(1639)));
    layer2_outputs(1271) <= not(layer1_outputs(844)) or (layer1_outputs(114));
    layer2_outputs(1272) <= (layer1_outputs(2491)) xor (layer1_outputs(2552));
    layer2_outputs(1273) <= not((layer1_outputs(1729)) or (layer1_outputs(1573)));
    layer2_outputs(1274) <= layer1_outputs(749);
    layer2_outputs(1275) <= (layer1_outputs(1496)) and not (layer1_outputs(796));
    layer2_outputs(1276) <= (layer1_outputs(93)) or (layer1_outputs(220));
    layer2_outputs(1277) <= not(layer1_outputs(2553));
    layer2_outputs(1278) <= not(layer1_outputs(91)) or (layer1_outputs(1173));
    layer2_outputs(1279) <= '1';
    layer2_outputs(1280) <= layer1_outputs(1737);
    layer2_outputs(1281) <= not((layer1_outputs(315)) and (layer1_outputs(762)));
    layer2_outputs(1282) <= not(layer1_outputs(2376)) or (layer1_outputs(1465));
    layer2_outputs(1283) <= '1';
    layer2_outputs(1284) <= (layer1_outputs(1170)) and not (layer1_outputs(2435));
    layer2_outputs(1285) <= not((layer1_outputs(464)) and (layer1_outputs(1284)));
    layer2_outputs(1286) <= not(layer1_outputs(1645)) or (layer1_outputs(1721));
    layer2_outputs(1287) <= layer1_outputs(1312);
    layer2_outputs(1288) <= (layer1_outputs(182)) and not (layer1_outputs(335));
    layer2_outputs(1289) <= (layer1_outputs(574)) and not (layer1_outputs(746));
    layer2_outputs(1290) <= not(layer1_outputs(1330)) or (layer1_outputs(1393));
    layer2_outputs(1291) <= not(layer1_outputs(929));
    layer2_outputs(1292) <= not(layer1_outputs(123)) or (layer1_outputs(1356));
    layer2_outputs(1293) <= (layer1_outputs(965)) or (layer1_outputs(459));
    layer2_outputs(1294) <= not(layer1_outputs(282));
    layer2_outputs(1295) <= (layer1_outputs(1521)) and not (layer1_outputs(109));
    layer2_outputs(1296) <= (layer1_outputs(2451)) or (layer1_outputs(55));
    layer2_outputs(1297) <= not(layer1_outputs(2192));
    layer2_outputs(1298) <= '1';
    layer2_outputs(1299) <= (layer1_outputs(2246)) or (layer1_outputs(826));
    layer2_outputs(1300) <= not(layer1_outputs(2018)) or (layer1_outputs(1139));
    layer2_outputs(1301) <= not(layer1_outputs(1323));
    layer2_outputs(1302) <= (layer1_outputs(754)) and not (layer1_outputs(1045));
    layer2_outputs(1303) <= not((layer1_outputs(1177)) or (layer1_outputs(1780)));
    layer2_outputs(1304) <= (layer1_outputs(901)) or (layer1_outputs(1145));
    layer2_outputs(1305) <= '1';
    layer2_outputs(1306) <= '1';
    layer2_outputs(1307) <= not(layer1_outputs(604)) or (layer1_outputs(2125));
    layer2_outputs(1308) <= (layer1_outputs(2239)) and not (layer1_outputs(1426));
    layer2_outputs(1309) <= '1';
    layer2_outputs(1310) <= (layer1_outputs(260)) and (layer1_outputs(2339));
    layer2_outputs(1311) <= '0';
    layer2_outputs(1312) <= not(layer1_outputs(336)) or (layer1_outputs(1725));
    layer2_outputs(1313) <= layer1_outputs(2129);
    layer2_outputs(1314) <= '1';
    layer2_outputs(1315) <= (layer1_outputs(1764)) and (layer1_outputs(1161));
    layer2_outputs(1316) <= not(layer1_outputs(1137));
    layer2_outputs(1317) <= not(layer1_outputs(1300)) or (layer1_outputs(2278));
    layer2_outputs(1318) <= layer1_outputs(1678);
    layer2_outputs(1319) <= '1';
    layer2_outputs(1320) <= layer1_outputs(304);
    layer2_outputs(1321) <= (layer1_outputs(1867)) and (layer1_outputs(926));
    layer2_outputs(1322) <= (layer1_outputs(673)) or (layer1_outputs(738));
    layer2_outputs(1323) <= '0';
    layer2_outputs(1324) <= (layer1_outputs(1755)) or (layer1_outputs(423));
    layer2_outputs(1325) <= not((layer1_outputs(1632)) or (layer1_outputs(1576)));
    layer2_outputs(1326) <= (layer1_outputs(2205)) or (layer1_outputs(1526));
    layer2_outputs(1327) <= (layer1_outputs(2431)) and (layer1_outputs(137));
    layer2_outputs(1328) <= not(layer1_outputs(246));
    layer2_outputs(1329) <= (layer1_outputs(452)) and (layer1_outputs(1123));
    layer2_outputs(1330) <= '0';
    layer2_outputs(1331) <= not((layer1_outputs(241)) or (layer1_outputs(130)));
    layer2_outputs(1332) <= (layer1_outputs(1055)) and not (layer1_outputs(1346));
    layer2_outputs(1333) <= layer1_outputs(2119);
    layer2_outputs(1334) <= not(layer1_outputs(394));
    layer2_outputs(1335) <= '1';
    layer2_outputs(1336) <= (layer1_outputs(338)) and not (layer1_outputs(2533));
    layer2_outputs(1337) <= '0';
    layer2_outputs(1338) <= not(layer1_outputs(2535));
    layer2_outputs(1339) <= layer1_outputs(106);
    layer2_outputs(1340) <= (layer1_outputs(2387)) and (layer1_outputs(1897));
    layer2_outputs(1341) <= not((layer1_outputs(690)) or (layer1_outputs(2038)));
    layer2_outputs(1342) <= (layer1_outputs(2543)) or (layer1_outputs(2549));
    layer2_outputs(1343) <= layer1_outputs(642);
    layer2_outputs(1344) <= not((layer1_outputs(1348)) and (layer1_outputs(1474)));
    layer2_outputs(1345) <= not((layer1_outputs(2105)) xor (layer1_outputs(858)));
    layer2_outputs(1346) <= (layer1_outputs(404)) and not (layer1_outputs(1342));
    layer2_outputs(1347) <= not(layer1_outputs(1737)) or (layer1_outputs(211));
    layer2_outputs(1348) <= not(layer1_outputs(979));
    layer2_outputs(1349) <= (layer1_outputs(2337)) and (layer1_outputs(1634));
    layer2_outputs(1350) <= '1';
    layer2_outputs(1351) <= (layer1_outputs(2099)) and not (layer1_outputs(2086));
    layer2_outputs(1352) <= '0';
    layer2_outputs(1353) <= (layer1_outputs(360)) and not (layer1_outputs(1136));
    layer2_outputs(1354) <= not(layer1_outputs(2222)) or (layer1_outputs(580));
    layer2_outputs(1355) <= not(layer1_outputs(1008));
    layer2_outputs(1356) <= not(layer1_outputs(560));
    layer2_outputs(1357) <= (layer1_outputs(884)) or (layer1_outputs(2148));
    layer2_outputs(1358) <= layer1_outputs(1774);
    layer2_outputs(1359) <= not(layer1_outputs(275)) or (layer1_outputs(1795));
    layer2_outputs(1360) <= not(layer1_outputs(322));
    layer2_outputs(1361) <= (layer1_outputs(754)) or (layer1_outputs(679));
    layer2_outputs(1362) <= '0';
    layer2_outputs(1363) <= not(layer1_outputs(1681)) or (layer1_outputs(1212));
    layer2_outputs(1364) <= (layer1_outputs(2131)) and (layer1_outputs(752));
    layer2_outputs(1365) <= '0';
    layer2_outputs(1366) <= '1';
    layer2_outputs(1367) <= not(layer1_outputs(1477));
    layer2_outputs(1368) <= '1';
    layer2_outputs(1369) <= layer1_outputs(1127);
    layer2_outputs(1370) <= not((layer1_outputs(2343)) and (layer1_outputs(600)));
    layer2_outputs(1371) <= layer1_outputs(2145);
    layer2_outputs(1372) <= not((layer1_outputs(1878)) or (layer1_outputs(400)));
    layer2_outputs(1373) <= '1';
    layer2_outputs(1374) <= layer1_outputs(1745);
    layer2_outputs(1375) <= not((layer1_outputs(1421)) or (layer1_outputs(850)));
    layer2_outputs(1376) <= not((layer1_outputs(1485)) and (layer1_outputs(873)));
    layer2_outputs(1377) <= '0';
    layer2_outputs(1378) <= layer1_outputs(184);
    layer2_outputs(1379) <= layer1_outputs(1321);
    layer2_outputs(1380) <= (layer1_outputs(1860)) and (layer1_outputs(1816));
    layer2_outputs(1381) <= layer1_outputs(1263);
    layer2_outputs(1382) <= not(layer1_outputs(2382)) or (layer1_outputs(66));
    layer2_outputs(1383) <= not(layer1_outputs(533));
    layer2_outputs(1384) <= (layer1_outputs(1316)) xor (layer1_outputs(1771));
    layer2_outputs(1385) <= (layer1_outputs(401)) and not (layer1_outputs(886));
    layer2_outputs(1386) <= '0';
    layer2_outputs(1387) <= not(layer1_outputs(399));
    layer2_outputs(1388) <= '0';
    layer2_outputs(1389) <= not((layer1_outputs(783)) or (layer1_outputs(1416)));
    layer2_outputs(1390) <= layer1_outputs(1078);
    layer2_outputs(1391) <= '0';
    layer2_outputs(1392) <= '1';
    layer2_outputs(1393) <= '0';
    layer2_outputs(1394) <= not(layer1_outputs(1953)) or (layer1_outputs(370));
    layer2_outputs(1395) <= '1';
    layer2_outputs(1396) <= not((layer1_outputs(1264)) and (layer1_outputs(2340)));
    layer2_outputs(1397) <= not((layer1_outputs(2536)) and (layer1_outputs(1303)));
    layer2_outputs(1398) <= not(layer1_outputs(32));
    layer2_outputs(1399) <= (layer1_outputs(1733)) and (layer1_outputs(1158));
    layer2_outputs(1400) <= layer1_outputs(1233);
    layer2_outputs(1401) <= layer1_outputs(2361);
    layer2_outputs(1402) <= (layer1_outputs(838)) or (layer1_outputs(2072));
    layer2_outputs(1403) <= (layer1_outputs(1226)) or (layer1_outputs(952));
    layer2_outputs(1404) <= not(layer1_outputs(1184)) or (layer1_outputs(2165));
    layer2_outputs(1405) <= '1';
    layer2_outputs(1406) <= layer1_outputs(2121);
    layer2_outputs(1407) <= (layer1_outputs(1925)) and (layer1_outputs(2532));
    layer2_outputs(1408) <= layer1_outputs(1604);
    layer2_outputs(1409) <= '1';
    layer2_outputs(1410) <= '1';
    layer2_outputs(1411) <= (layer1_outputs(675)) or (layer1_outputs(2006));
    layer2_outputs(1412) <= (layer1_outputs(2404)) or (layer1_outputs(481));
    layer2_outputs(1413) <= not((layer1_outputs(1163)) and (layer1_outputs(114)));
    layer2_outputs(1414) <= '1';
    layer2_outputs(1415) <= (layer1_outputs(191)) and not (layer1_outputs(1716));
    layer2_outputs(1416) <= not(layer1_outputs(1529));
    layer2_outputs(1417) <= (layer1_outputs(1549)) and not (layer1_outputs(1289));
    layer2_outputs(1418) <= (layer1_outputs(2093)) and not (layer1_outputs(1718));
    layer2_outputs(1419) <= '1';
    layer2_outputs(1420) <= (layer1_outputs(1148)) and (layer1_outputs(1917));
    layer2_outputs(1421) <= layer1_outputs(1493);
    layer2_outputs(1422) <= '1';
    layer2_outputs(1423) <= not(layer1_outputs(149)) or (layer1_outputs(2015));
    layer2_outputs(1424) <= not(layer1_outputs(1691)) or (layer1_outputs(414));
    layer2_outputs(1425) <= not(layer1_outputs(1830));
    layer2_outputs(1426) <= not(layer1_outputs(1153)) or (layer1_outputs(2088));
    layer2_outputs(1427) <= '1';
    layer2_outputs(1428) <= layer1_outputs(169);
    layer2_outputs(1429) <= (layer1_outputs(1641)) and not (layer1_outputs(802));
    layer2_outputs(1430) <= not((layer1_outputs(431)) and (layer1_outputs(2253)));
    layer2_outputs(1431) <= (layer1_outputs(373)) and (layer1_outputs(1586));
    layer2_outputs(1432) <= (layer1_outputs(903)) and not (layer1_outputs(1663));
    layer2_outputs(1433) <= (layer1_outputs(1229)) or (layer1_outputs(1987));
    layer2_outputs(1434) <= not(layer1_outputs(723));
    layer2_outputs(1435) <= not(layer1_outputs(1214));
    layer2_outputs(1436) <= not(layer1_outputs(770));
    layer2_outputs(1437) <= layer1_outputs(61);
    layer2_outputs(1438) <= layer1_outputs(2160);
    layer2_outputs(1439) <= layer1_outputs(1516);
    layer2_outputs(1440) <= (layer1_outputs(2479)) and (layer1_outputs(1831));
    layer2_outputs(1441) <= (layer1_outputs(1840)) xor (layer1_outputs(296));
    layer2_outputs(1442) <= (layer1_outputs(1957)) and (layer1_outputs(1864));
    layer2_outputs(1443) <= not((layer1_outputs(2312)) xor (layer1_outputs(2013)));
    layer2_outputs(1444) <= '0';
    layer2_outputs(1445) <= '1';
    layer2_outputs(1446) <= layer1_outputs(2500);
    layer2_outputs(1447) <= layer1_outputs(202);
    layer2_outputs(1448) <= (layer1_outputs(256)) and not (layer1_outputs(2432));
    layer2_outputs(1449) <= (layer1_outputs(1110)) or (layer1_outputs(81));
    layer2_outputs(1450) <= (layer1_outputs(1790)) and (layer1_outputs(791));
    layer2_outputs(1451) <= '0';
    layer2_outputs(1452) <= '0';
    layer2_outputs(1453) <= not((layer1_outputs(2234)) or (layer1_outputs(1509)));
    layer2_outputs(1454) <= (layer1_outputs(476)) and (layer1_outputs(446));
    layer2_outputs(1455) <= not(layer1_outputs(1636));
    layer2_outputs(1456) <= not(layer1_outputs(41));
    layer2_outputs(1457) <= layer1_outputs(848);
    layer2_outputs(1458) <= '1';
    layer2_outputs(1459) <= not((layer1_outputs(263)) xor (layer1_outputs(737)));
    layer2_outputs(1460) <= not(layer1_outputs(85));
    layer2_outputs(1461) <= not((layer1_outputs(2069)) and (layer1_outputs(1007)));
    layer2_outputs(1462) <= not((layer1_outputs(206)) or (layer1_outputs(985)));
    layer2_outputs(1463) <= not(layer1_outputs(833)) or (layer1_outputs(1911));
    layer2_outputs(1464) <= '1';
    layer2_outputs(1465) <= not(layer1_outputs(2113));
    layer2_outputs(1466) <= (layer1_outputs(2472)) or (layer1_outputs(5));
    layer2_outputs(1467) <= (layer1_outputs(1444)) and (layer1_outputs(222));
    layer2_outputs(1468) <= not(layer1_outputs(283)) or (layer1_outputs(1510));
    layer2_outputs(1469) <= not((layer1_outputs(1798)) and (layer1_outputs(965)));
    layer2_outputs(1470) <= (layer1_outputs(47)) and not (layer1_outputs(99));
    layer2_outputs(1471) <= (layer1_outputs(321)) or (layer1_outputs(2287));
    layer2_outputs(1472) <= '0';
    layer2_outputs(1473) <= (layer1_outputs(2384)) and not (layer1_outputs(2132));
    layer2_outputs(1474) <= not(layer1_outputs(1413)) or (layer1_outputs(36));
    layer2_outputs(1475) <= (layer1_outputs(2296)) or (layer1_outputs(1952));
    layer2_outputs(1476) <= not(layer1_outputs(1182));
    layer2_outputs(1477) <= not((layer1_outputs(790)) and (layer1_outputs(2531)));
    layer2_outputs(1478) <= '1';
    layer2_outputs(1479) <= layer1_outputs(1232);
    layer2_outputs(1480) <= '1';
    layer2_outputs(1481) <= not((layer1_outputs(310)) and (layer1_outputs(1584)));
    layer2_outputs(1482) <= '0';
    layer2_outputs(1483) <= (layer1_outputs(1754)) and not (layer1_outputs(2501));
    layer2_outputs(1484) <= not((layer1_outputs(2239)) and (layer1_outputs(1578)));
    layer2_outputs(1485) <= not((layer1_outputs(878)) and (layer1_outputs(78)));
    layer2_outputs(1486) <= layer1_outputs(1396);
    layer2_outputs(1487) <= layer1_outputs(1751);
    layer2_outputs(1488) <= layer1_outputs(135);
    layer2_outputs(1489) <= not(layer1_outputs(1051));
    layer2_outputs(1490) <= '0';
    layer2_outputs(1491) <= (layer1_outputs(385)) and not (layer1_outputs(1017));
    layer2_outputs(1492) <= '0';
    layer2_outputs(1493) <= layer1_outputs(2007);
    layer2_outputs(1494) <= not((layer1_outputs(1474)) and (layer1_outputs(328)));
    layer2_outputs(1495) <= (layer1_outputs(1109)) and not (layer1_outputs(1903));
    layer2_outputs(1496) <= '0';
    layer2_outputs(1497) <= not((layer1_outputs(1240)) or (layer1_outputs(905)));
    layer2_outputs(1498) <= (layer1_outputs(1914)) and (layer1_outputs(398));
    layer2_outputs(1499) <= (layer1_outputs(2251)) or (layer1_outputs(1120));
    layer2_outputs(1500) <= not(layer1_outputs(1176));
    layer2_outputs(1501) <= not((layer1_outputs(290)) or (layer1_outputs(207)));
    layer2_outputs(1502) <= (layer1_outputs(1229)) and (layer1_outputs(24));
    layer2_outputs(1503) <= (layer1_outputs(2507)) or (layer1_outputs(1918));
    layer2_outputs(1504) <= not(layer1_outputs(1689));
    layer2_outputs(1505) <= (layer1_outputs(118)) and (layer1_outputs(350));
    layer2_outputs(1506) <= (layer1_outputs(1291)) xor (layer1_outputs(626));
    layer2_outputs(1507) <= '0';
    layer2_outputs(1508) <= not(layer1_outputs(867));
    layer2_outputs(1509) <= not(layer1_outputs(2465)) or (layer1_outputs(469));
    layer2_outputs(1510) <= not(layer1_outputs(2152)) or (layer1_outputs(713));
    layer2_outputs(1511) <= not(layer1_outputs(1343));
    layer2_outputs(1512) <= layer1_outputs(1896);
    layer2_outputs(1513) <= layer1_outputs(142);
    layer2_outputs(1514) <= (layer1_outputs(2207)) and (layer1_outputs(2171));
    layer2_outputs(1515) <= not(layer1_outputs(1657));
    layer2_outputs(1516) <= layer1_outputs(1125);
    layer2_outputs(1517) <= (layer1_outputs(720)) and not (layer1_outputs(549));
    layer2_outputs(1518) <= '1';
    layer2_outputs(1519) <= not(layer1_outputs(1065)) or (layer1_outputs(523));
    layer2_outputs(1520) <= '1';
    layer2_outputs(1521) <= (layer1_outputs(2526)) and not (layer1_outputs(1608));
    layer2_outputs(1522) <= layer1_outputs(1674);
    layer2_outputs(1523) <= not(layer1_outputs(1387));
    layer2_outputs(1524) <= '0';
    layer2_outputs(1525) <= not(layer1_outputs(1724));
    layer2_outputs(1526) <= '0';
    layer2_outputs(1527) <= (layer1_outputs(1282)) and not (layer1_outputs(2528));
    layer2_outputs(1528) <= not(layer1_outputs(13)) or (layer1_outputs(1195));
    layer2_outputs(1529) <= not((layer1_outputs(1733)) and (layer1_outputs(2076)));
    layer2_outputs(1530) <= layer1_outputs(271);
    layer2_outputs(1531) <= not((layer1_outputs(2060)) or (layer1_outputs(361)));
    layer2_outputs(1532) <= (layer1_outputs(133)) and not (layer1_outputs(2221));
    layer2_outputs(1533) <= (layer1_outputs(660)) and not (layer1_outputs(2509));
    layer2_outputs(1534) <= (layer1_outputs(2033)) xor (layer1_outputs(259));
    layer2_outputs(1535) <= not(layer1_outputs(1368));
    layer2_outputs(1536) <= '0';
    layer2_outputs(1537) <= (layer1_outputs(1871)) or (layer1_outputs(515));
    layer2_outputs(1538) <= layer1_outputs(1156);
    layer2_outputs(1539) <= layer1_outputs(1367);
    layer2_outputs(1540) <= layer1_outputs(1243);
    layer2_outputs(1541) <= (layer1_outputs(878)) xor (layer1_outputs(788));
    layer2_outputs(1542) <= not((layer1_outputs(934)) and (layer1_outputs(146)));
    layer2_outputs(1543) <= '1';
    layer2_outputs(1544) <= not(layer1_outputs(2254));
    layer2_outputs(1545) <= not(layer1_outputs(1431)) or (layer1_outputs(277));
    layer2_outputs(1546) <= '0';
    layer2_outputs(1547) <= '1';
    layer2_outputs(1548) <= '0';
    layer2_outputs(1549) <= not(layer1_outputs(2263));
    layer2_outputs(1550) <= (layer1_outputs(1209)) and (layer1_outputs(627));
    layer2_outputs(1551) <= layer1_outputs(2129);
    layer2_outputs(1552) <= (layer1_outputs(182)) or (layer1_outputs(1346));
    layer2_outputs(1553) <= not(layer1_outputs(767)) or (layer1_outputs(228));
    layer2_outputs(1554) <= (layer1_outputs(2190)) or (layer1_outputs(159));
    layer2_outputs(1555) <= '0';
    layer2_outputs(1556) <= (layer1_outputs(1332)) and (layer1_outputs(1843));
    layer2_outputs(1557) <= not(layer1_outputs(350)) or (layer1_outputs(2289));
    layer2_outputs(1558) <= '0';
    layer2_outputs(1559) <= '0';
    layer2_outputs(1560) <= '1';
    layer2_outputs(1561) <= '1';
    layer2_outputs(1562) <= not((layer1_outputs(552)) and (layer1_outputs(569)));
    layer2_outputs(1563) <= layer1_outputs(1024);
    layer2_outputs(1564) <= not(layer1_outputs(274));
    layer2_outputs(1565) <= '0';
    layer2_outputs(1566) <= not((layer1_outputs(1549)) or (layer1_outputs(1461)));
    layer2_outputs(1567) <= not(layer1_outputs(2394));
    layer2_outputs(1568) <= not(layer1_outputs(588)) or (layer1_outputs(623));
    layer2_outputs(1569) <= (layer1_outputs(570)) and not (layer1_outputs(224));
    layer2_outputs(1570) <= layer1_outputs(1185);
    layer2_outputs(1571) <= '0';
    layer2_outputs(1572) <= layer1_outputs(429);
    layer2_outputs(1573) <= not(layer1_outputs(357)) or (layer1_outputs(1324));
    layer2_outputs(1574) <= (layer1_outputs(2035)) and (layer1_outputs(425));
    layer2_outputs(1575) <= not((layer1_outputs(1442)) and (layer1_outputs(33)));
    layer2_outputs(1576) <= not(layer1_outputs(1726));
    layer2_outputs(1577) <= not((layer1_outputs(1038)) or (layer1_outputs(228)));
    layer2_outputs(1578) <= not((layer1_outputs(564)) and (layer1_outputs(1784)));
    layer2_outputs(1579) <= not(layer1_outputs(1159)) or (layer1_outputs(696));
    layer2_outputs(1580) <= layer1_outputs(2136);
    layer2_outputs(1581) <= not((layer1_outputs(775)) and (layer1_outputs(497)));
    layer2_outputs(1582) <= (layer1_outputs(313)) and (layer1_outputs(1040));
    layer2_outputs(1583) <= '1';
    layer2_outputs(1584) <= (layer1_outputs(2079)) or (layer1_outputs(1782));
    layer2_outputs(1585) <= '1';
    layer2_outputs(1586) <= not(layer1_outputs(1326)) or (layer1_outputs(2061));
    layer2_outputs(1587) <= layer1_outputs(505);
    layer2_outputs(1588) <= (layer1_outputs(463)) xor (layer1_outputs(1327));
    layer2_outputs(1589) <= not((layer1_outputs(922)) and (layer1_outputs(1248)));
    layer2_outputs(1590) <= not(layer1_outputs(1617));
    layer2_outputs(1591) <= not((layer1_outputs(479)) xor (layer1_outputs(2333)));
    layer2_outputs(1592) <= '0';
    layer2_outputs(1593) <= not(layer1_outputs(610));
    layer2_outputs(1594) <= (layer1_outputs(2182)) and (layer1_outputs(1653));
    layer2_outputs(1595) <= '0';
    layer2_outputs(1596) <= layer1_outputs(1113);
    layer2_outputs(1597) <= not(layer1_outputs(912));
    layer2_outputs(1598) <= not(layer1_outputs(613)) or (layer1_outputs(571));
    layer2_outputs(1599) <= layer1_outputs(90);
    layer2_outputs(1600) <= not(layer1_outputs(1044)) or (layer1_outputs(95));
    layer2_outputs(1601) <= layer1_outputs(348);
    layer2_outputs(1602) <= layer1_outputs(2346);
    layer2_outputs(1603) <= layer1_outputs(850);
    layer2_outputs(1604) <= not(layer1_outputs(968)) or (layer1_outputs(1274));
    layer2_outputs(1605) <= (layer1_outputs(1985)) and (layer1_outputs(2297));
    layer2_outputs(1606) <= (layer1_outputs(2237)) and not (layer1_outputs(1598));
    layer2_outputs(1607) <= not(layer1_outputs(2336));
    layer2_outputs(1608) <= not(layer1_outputs(346));
    layer2_outputs(1609) <= '0';
    layer2_outputs(1610) <= '1';
    layer2_outputs(1611) <= layer1_outputs(449);
    layer2_outputs(1612) <= not(layer1_outputs(2211));
    layer2_outputs(1613) <= not(layer1_outputs(2462)) or (layer1_outputs(484));
    layer2_outputs(1614) <= layer1_outputs(1742);
    layer2_outputs(1615) <= '1';
    layer2_outputs(1616) <= not((layer1_outputs(957)) and (layer1_outputs(885)));
    layer2_outputs(1617) <= not(layer1_outputs(202));
    layer2_outputs(1618) <= (layer1_outputs(889)) or (layer1_outputs(1024));
    layer2_outputs(1619) <= not(layer1_outputs(1083));
    layer2_outputs(1620) <= not(layer1_outputs(1641)) or (layer1_outputs(1971));
    layer2_outputs(1621) <= not(layer1_outputs(861));
    layer2_outputs(1622) <= (layer1_outputs(1785)) and (layer1_outputs(559));
    layer2_outputs(1623) <= (layer1_outputs(156)) or (layer1_outputs(2495));
    layer2_outputs(1624) <= not((layer1_outputs(907)) or (layer1_outputs(27)));
    layer2_outputs(1625) <= not(layer1_outputs(1908));
    layer2_outputs(1626) <= (layer1_outputs(1409)) and not (layer1_outputs(1844));
    layer2_outputs(1627) <= '1';
    layer2_outputs(1628) <= (layer1_outputs(2499)) and (layer1_outputs(876));
    layer2_outputs(1629) <= not(layer1_outputs(2075));
    layer2_outputs(1630) <= not(layer1_outputs(2442));
    layer2_outputs(1631) <= not(layer1_outputs(1881)) or (layer1_outputs(2393));
    layer2_outputs(1632) <= not((layer1_outputs(2161)) or (layer1_outputs(1263)));
    layer2_outputs(1633) <= not((layer1_outputs(1585)) or (layer1_outputs(375)));
    layer2_outputs(1634) <= not((layer1_outputs(1194)) or (layer1_outputs(2438)));
    layer2_outputs(1635) <= not((layer1_outputs(1245)) and (layer1_outputs(2376)));
    layer2_outputs(1636) <= (layer1_outputs(1102)) or (layer1_outputs(2144));
    layer2_outputs(1637) <= not(layer1_outputs(2172));
    layer2_outputs(1638) <= not((layer1_outputs(630)) or (layer1_outputs(1662)));
    layer2_outputs(1639) <= (layer1_outputs(2128)) and not (layer1_outputs(1639));
    layer2_outputs(1640) <= '0';
    layer2_outputs(1641) <= (layer1_outputs(1397)) and (layer1_outputs(2433));
    layer2_outputs(1642) <= '1';
    layer2_outputs(1643) <= '0';
    layer2_outputs(1644) <= not(layer1_outputs(1901)) or (layer1_outputs(639));
    layer2_outputs(1645) <= (layer1_outputs(215)) and not (layer1_outputs(697));
    layer2_outputs(1646) <= (layer1_outputs(1133)) or (layer1_outputs(1435));
    layer2_outputs(1647) <= not(layer1_outputs(1261));
    layer2_outputs(1648) <= layer1_outputs(1406);
    layer2_outputs(1649) <= layer1_outputs(1331);
    layer2_outputs(1650) <= not(layer1_outputs(377));
    layer2_outputs(1651) <= (layer1_outputs(1575)) and not (layer1_outputs(2030));
    layer2_outputs(1652) <= not(layer1_outputs(1218)) or (layer1_outputs(434));
    layer2_outputs(1653) <= '1';
    layer2_outputs(1654) <= not(layer1_outputs(444));
    layer2_outputs(1655) <= '1';
    layer2_outputs(1656) <= (layer1_outputs(1186)) and (layer1_outputs(1457));
    layer2_outputs(1657) <= not((layer1_outputs(1223)) xor (layer1_outputs(1777)));
    layer2_outputs(1658) <= not(layer1_outputs(2518));
    layer2_outputs(1659) <= layer1_outputs(841);
    layer2_outputs(1660) <= '1';
    layer2_outputs(1661) <= layer1_outputs(1241);
    layer2_outputs(1662) <= layer1_outputs(577);
    layer2_outputs(1663) <= not(layer1_outputs(1162)) or (layer1_outputs(626));
    layer2_outputs(1664) <= not((layer1_outputs(1992)) xor (layer1_outputs(1015)));
    layer2_outputs(1665) <= (layer1_outputs(647)) xor (layer1_outputs(2516));
    layer2_outputs(1666) <= layer1_outputs(428);
    layer2_outputs(1667) <= not((layer1_outputs(1547)) or (layer1_outputs(1089)));
    layer2_outputs(1668) <= '0';
    layer2_outputs(1669) <= '1';
    layer2_outputs(1670) <= (layer1_outputs(1206)) or (layer1_outputs(1873));
    layer2_outputs(1671) <= (layer1_outputs(1891)) and not (layer1_outputs(1544));
    layer2_outputs(1672) <= not(layer1_outputs(1670)) or (layer1_outputs(519));
    layer2_outputs(1673) <= not((layer1_outputs(1122)) or (layer1_outputs(638)));
    layer2_outputs(1674) <= not((layer1_outputs(1514)) or (layer1_outputs(964)));
    layer2_outputs(1675) <= layer1_outputs(12);
    layer2_outputs(1676) <= not(layer1_outputs(2286));
    layer2_outputs(1677) <= (layer1_outputs(2480)) and not (layer1_outputs(141));
    layer2_outputs(1678) <= not(layer1_outputs(1252));
    layer2_outputs(1679) <= not(layer1_outputs(242)) or (layer1_outputs(1741));
    layer2_outputs(1680) <= not((layer1_outputs(1327)) and (layer1_outputs(2076)));
    layer2_outputs(1681) <= (layer1_outputs(607)) and not (layer1_outputs(254));
    layer2_outputs(1682) <= not(layer1_outputs(243));
    layer2_outputs(1683) <= '0';
    layer2_outputs(1684) <= (layer1_outputs(1031)) or (layer1_outputs(2540));
    layer2_outputs(1685) <= '1';
    layer2_outputs(1686) <= (layer1_outputs(2252)) and not (layer1_outputs(2369));
    layer2_outputs(1687) <= not((layer1_outputs(1806)) or (layer1_outputs(2374)));
    layer2_outputs(1688) <= '0';
    layer2_outputs(1689) <= not(layer1_outputs(1915));
    layer2_outputs(1690) <= '1';
    layer2_outputs(1691) <= (layer1_outputs(1524)) and not (layer1_outputs(1177));
    layer2_outputs(1692) <= not(layer1_outputs(1834)) or (layer1_outputs(1961));
    layer2_outputs(1693) <= (layer1_outputs(1706)) and (layer1_outputs(758));
    layer2_outputs(1694) <= (layer1_outputs(591)) and not (layer1_outputs(1942));
    layer2_outputs(1695) <= not((layer1_outputs(1473)) or (layer1_outputs(1059)));
    layer2_outputs(1696) <= not(layer1_outputs(1863));
    layer2_outputs(1697) <= layer1_outputs(39);
    layer2_outputs(1698) <= layer1_outputs(2043);
    layer2_outputs(1699) <= (layer1_outputs(1352)) and not (layer1_outputs(919));
    layer2_outputs(1700) <= '0';
    layer2_outputs(1701) <= layer1_outputs(257);
    layer2_outputs(1702) <= layer1_outputs(238);
    layer2_outputs(1703) <= not(layer1_outputs(1501)) or (layer1_outputs(567));
    layer2_outputs(1704) <= not((layer1_outputs(1866)) or (layer1_outputs(615)));
    layer2_outputs(1705) <= not(layer1_outputs(1940));
    layer2_outputs(1706) <= layer1_outputs(1487);
    layer2_outputs(1707) <= (layer1_outputs(1115)) and (layer1_outputs(1471));
    layer2_outputs(1708) <= not(layer1_outputs(129));
    layer2_outputs(1709) <= (layer1_outputs(1280)) and (layer1_outputs(1679));
    layer2_outputs(1710) <= not(layer1_outputs(313));
    layer2_outputs(1711) <= not(layer1_outputs(667));
    layer2_outputs(1712) <= not(layer1_outputs(2031));
    layer2_outputs(1713) <= not((layer1_outputs(263)) or (layer1_outputs(2011)));
    layer2_outputs(1714) <= '1';
    layer2_outputs(1715) <= '0';
    layer2_outputs(1716) <= (layer1_outputs(726)) or (layer1_outputs(954));
    layer2_outputs(1717) <= not((layer1_outputs(1909)) or (layer1_outputs(43)));
    layer2_outputs(1718) <= not(layer1_outputs(1275)) or (layer1_outputs(492));
    layer2_outputs(1719) <= (layer1_outputs(1714)) and (layer1_outputs(753));
    layer2_outputs(1720) <= '1';
    layer2_outputs(1721) <= (layer1_outputs(1956)) and not (layer1_outputs(704));
    layer2_outputs(1722) <= '0';
    layer2_outputs(1723) <= not((layer1_outputs(305)) and (layer1_outputs(1647)));
    layer2_outputs(1724) <= (layer1_outputs(2513)) and (layer1_outputs(1814));
    layer2_outputs(1725) <= '1';
    layer2_outputs(1726) <= not(layer1_outputs(2271)) or (layer1_outputs(2480));
    layer2_outputs(1727) <= not((layer1_outputs(372)) or (layer1_outputs(1057)));
    layer2_outputs(1728) <= not(layer1_outputs(848)) or (layer1_outputs(854));
    layer2_outputs(1729) <= layer1_outputs(2330);
    layer2_outputs(1730) <= '0';
    layer2_outputs(1731) <= layer1_outputs(1595);
    layer2_outputs(1732) <= (layer1_outputs(1728)) and not (layer1_outputs(1389));
    layer2_outputs(1733) <= not(layer1_outputs(975)) or (layer1_outputs(842));
    layer2_outputs(1734) <= (layer1_outputs(2122)) and (layer1_outputs(1414));
    layer2_outputs(1735) <= layer1_outputs(1998);
    layer2_outputs(1736) <= not(layer1_outputs(480)) or (layer1_outputs(760));
    layer2_outputs(1737) <= not(layer1_outputs(602));
    layer2_outputs(1738) <= '1';
    layer2_outputs(1739) <= (layer1_outputs(1722)) and (layer1_outputs(1183));
    layer2_outputs(1740) <= '1';
    layer2_outputs(1741) <= not(layer1_outputs(1216)) or (layer1_outputs(1656));
    layer2_outputs(1742) <= (layer1_outputs(906)) and not (layer1_outputs(1964));
    layer2_outputs(1743) <= not((layer1_outputs(2003)) and (layer1_outputs(1363)));
    layer2_outputs(1744) <= layer1_outputs(1334);
    layer2_outputs(1745) <= (layer1_outputs(776)) and not (layer1_outputs(899));
    layer2_outputs(1746) <= (layer1_outputs(2380)) and not (layer1_outputs(1578));
    layer2_outputs(1747) <= not((layer1_outputs(52)) and (layer1_outputs(80)));
    layer2_outputs(1748) <= (layer1_outputs(1550)) and (layer1_outputs(1487));
    layer2_outputs(1749) <= not(layer1_outputs(2120));
    layer2_outputs(1750) <= '0';
    layer2_outputs(1751) <= layer1_outputs(2262);
    layer2_outputs(1752) <= (layer1_outputs(1386)) and not (layer1_outputs(1615));
    layer2_outputs(1753) <= layer1_outputs(2140);
    layer2_outputs(1754) <= not(layer1_outputs(107)) or (layer1_outputs(443));
    layer2_outputs(1755) <= not((layer1_outputs(2107)) or (layer1_outputs(2238)));
    layer2_outputs(1756) <= not((layer1_outputs(411)) and (layer1_outputs(2419)));
    layer2_outputs(1757) <= '1';
    layer2_outputs(1758) <= '0';
    layer2_outputs(1759) <= not(layer1_outputs(1215)) or (layer1_outputs(1247));
    layer2_outputs(1760) <= not(layer1_outputs(1714)) or (layer1_outputs(1693));
    layer2_outputs(1761) <= not(layer1_outputs(1099));
    layer2_outputs(1762) <= (layer1_outputs(1012)) and (layer1_outputs(191));
    layer2_outputs(1763) <= not((layer1_outputs(2244)) and (layer1_outputs(489)));
    layer2_outputs(1764) <= (layer1_outputs(1151)) and not (layer1_outputs(1121));
    layer2_outputs(1765) <= '1';
    layer2_outputs(1766) <= '0';
    layer2_outputs(1767) <= (layer1_outputs(1713)) and (layer1_outputs(351));
    layer2_outputs(1768) <= not(layer1_outputs(160));
    layer2_outputs(1769) <= not(layer1_outputs(1761));
    layer2_outputs(1770) <= not(layer1_outputs(1848)) or (layer1_outputs(1860));
    layer2_outputs(1771) <= not(layer1_outputs(832));
    layer2_outputs(1772) <= not(layer1_outputs(512));
    layer2_outputs(1773) <= not(layer1_outputs(1261)) or (layer1_outputs(1143));
    layer2_outputs(1774) <= '1';
    layer2_outputs(1775) <= layer1_outputs(1466);
    layer2_outputs(1776) <= '0';
    layer2_outputs(1777) <= (layer1_outputs(1658)) or (layer1_outputs(1805));
    layer2_outputs(1778) <= layer1_outputs(831);
    layer2_outputs(1779) <= layer1_outputs(1502);
    layer2_outputs(1780) <= (layer1_outputs(937)) or (layer1_outputs(2047));
    layer2_outputs(1781) <= (layer1_outputs(2374)) xor (layer1_outputs(1803));
    layer2_outputs(1782) <= not(layer1_outputs(457));
    layer2_outputs(1783) <= not((layer1_outputs(1530)) and (layer1_outputs(1899)));
    layer2_outputs(1784) <= '1';
    layer2_outputs(1785) <= layer1_outputs(1146);
    layer2_outputs(1786) <= not(layer1_outputs(2537));
    layer2_outputs(1787) <= layer1_outputs(491);
    layer2_outputs(1788) <= not(layer1_outputs(484)) or (layer1_outputs(1776));
    layer2_outputs(1789) <= layer1_outputs(2181);
    layer2_outputs(1790) <= not(layer1_outputs(998));
    layer2_outputs(1791) <= '1';
    layer2_outputs(1792) <= layer1_outputs(563);
    layer2_outputs(1793) <= (layer1_outputs(1842)) and (layer1_outputs(2302));
    layer2_outputs(1794) <= '1';
    layer2_outputs(1795) <= not((layer1_outputs(2157)) or (layer1_outputs(1809)));
    layer2_outputs(1796) <= '1';
    layer2_outputs(1797) <= not(layer1_outputs(900));
    layer2_outputs(1798) <= (layer1_outputs(1083)) or (layer1_outputs(962));
    layer2_outputs(1799) <= not((layer1_outputs(293)) xor (layer1_outputs(2546)));
    layer2_outputs(1800) <= (layer1_outputs(1344)) and not (layer1_outputs(1968));
    layer2_outputs(1801) <= layer1_outputs(587);
    layer2_outputs(1802) <= not(layer1_outputs(213));
    layer2_outputs(1803) <= '1';
    layer2_outputs(1804) <= (layer1_outputs(597)) and not (layer1_outputs(2485));
    layer2_outputs(1805) <= not((layer1_outputs(553)) and (layer1_outputs(2227)));
    layer2_outputs(1806) <= not(layer1_outputs(2196)) or (layer1_outputs(440));
    layer2_outputs(1807) <= not((layer1_outputs(881)) and (layer1_outputs(1210)));
    layer2_outputs(1808) <= (layer1_outputs(312)) and not (layer1_outputs(805));
    layer2_outputs(1809) <= not(layer1_outputs(1606));
    layer2_outputs(1810) <= not(layer1_outputs(1810)) or (layer1_outputs(221));
    layer2_outputs(1811) <= (layer1_outputs(2529)) and not (layer1_outputs(1902));
    layer2_outputs(1812) <= (layer1_outputs(384)) or (layer1_outputs(2544));
    layer2_outputs(1813) <= '0';
    layer2_outputs(1814) <= layer1_outputs(10);
    layer2_outputs(1815) <= not((layer1_outputs(643)) or (layer1_outputs(2056)));
    layer2_outputs(1816) <= not((layer1_outputs(1723)) or (layer1_outputs(1914)));
    layer2_outputs(1817) <= not(layer1_outputs(1350)) or (layer1_outputs(2118));
    layer2_outputs(1818) <= layer1_outputs(1200);
    layer2_outputs(1819) <= (layer1_outputs(1352)) and not (layer1_outputs(668));
    layer2_outputs(1820) <= layer1_outputs(1819);
    layer2_outputs(1821) <= (layer1_outputs(164)) and (layer1_outputs(2230));
    layer2_outputs(1822) <= (layer1_outputs(150)) and (layer1_outputs(1999));
    layer2_outputs(1823) <= not((layer1_outputs(1691)) or (layer1_outputs(2147)));
    layer2_outputs(1824) <= (layer1_outputs(605)) and not (layer1_outputs(2167));
    layer2_outputs(1825) <= layer1_outputs(1809);
    layer2_outputs(1826) <= not((layer1_outputs(1032)) and (layer1_outputs(2009)));
    layer2_outputs(1827) <= layer1_outputs(727);
    layer2_outputs(1828) <= not((layer1_outputs(989)) or (layer1_outputs(471)));
    layer2_outputs(1829) <= not(layer1_outputs(1949));
    layer2_outputs(1830) <= layer1_outputs(1935);
    layer2_outputs(1831) <= (layer1_outputs(2554)) or (layer1_outputs(1063));
    layer2_outputs(1832) <= '1';
    layer2_outputs(1833) <= layer1_outputs(2088);
    layer2_outputs(1834) <= (layer1_outputs(2438)) and (layer1_outputs(2146));
    layer2_outputs(1835) <= not(layer1_outputs(1626)) or (layer1_outputs(302));
    layer2_outputs(1836) <= (layer1_outputs(1512)) or (layer1_outputs(1660));
    layer2_outputs(1837) <= not((layer1_outputs(1794)) or (layer1_outputs(218)));
    layer2_outputs(1838) <= not(layer1_outputs(1943));
    layer2_outputs(1839) <= '1';
    layer2_outputs(1840) <= (layer1_outputs(1060)) and not (layer1_outputs(785));
    layer2_outputs(1841) <= layer1_outputs(1796);
    layer2_outputs(1842) <= not(layer1_outputs(295)) or (layer1_outputs(176));
    layer2_outputs(1843) <= layer1_outputs(71);
    layer2_outputs(1844) <= '0';
    layer2_outputs(1845) <= (layer1_outputs(1962)) or (layer1_outputs(1811));
    layer2_outputs(1846) <= not(layer1_outputs(409));
    layer2_outputs(1847) <= (layer1_outputs(1139)) and (layer1_outputs(718));
    layer2_outputs(1848) <= not(layer1_outputs(372));
    layer2_outputs(1849) <= layer1_outputs(699);
    layer2_outputs(1850) <= not((layer1_outputs(652)) xor (layer1_outputs(564)));
    layer2_outputs(1851) <= (layer1_outputs(236)) and (layer1_outputs(2476));
    layer2_outputs(1852) <= layer1_outputs(967);
    layer2_outputs(1853) <= layer1_outputs(1318);
    layer2_outputs(1854) <= not(layer1_outputs(1920)) or (layer1_outputs(485));
    layer2_outputs(1855) <= (layer1_outputs(2157)) and (layer1_outputs(286));
    layer2_outputs(1856) <= not(layer1_outputs(1623));
    layer2_outputs(1857) <= not((layer1_outputs(529)) and (layer1_outputs(2078)));
    layer2_outputs(1858) <= '1';
    layer2_outputs(1859) <= not((layer1_outputs(475)) and (layer1_outputs(1397)));
    layer2_outputs(1860) <= (layer1_outputs(870)) or (layer1_outputs(1951));
    layer2_outputs(1861) <= not(layer1_outputs(294));
    layer2_outputs(1862) <= (layer1_outputs(1278)) and not (layer1_outputs(1167));
    layer2_outputs(1863) <= layer1_outputs(1098);
    layer2_outputs(1864) <= not(layer1_outputs(2205)) or (layer1_outputs(950));
    layer2_outputs(1865) <= layer1_outputs(1075);
    layer2_outputs(1866) <= '1';
    layer2_outputs(1867) <= (layer1_outputs(302)) and (layer1_outputs(1601));
    layer2_outputs(1868) <= (layer1_outputs(1746)) and (layer1_outputs(1756));
    layer2_outputs(1869) <= not(layer1_outputs(2364)) or (layer1_outputs(18));
    layer2_outputs(1870) <= not((layer1_outputs(1744)) or (layer1_outputs(971)));
    layer2_outputs(1871) <= not(layer1_outputs(1209)) or (layer1_outputs(1732));
    layer2_outputs(1872) <= '1';
    layer2_outputs(1873) <= layer1_outputs(1853);
    layer2_outputs(1874) <= not(layer1_outputs(1683));
    layer2_outputs(1875) <= not(layer1_outputs(429)) or (layer1_outputs(893));
    layer2_outputs(1876) <= (layer1_outputs(1773)) and (layer1_outputs(953));
    layer2_outputs(1877) <= (layer1_outputs(2010)) and not (layer1_outputs(631));
    layer2_outputs(1878) <= not((layer1_outputs(2021)) or (layer1_outputs(2398)));
    layer2_outputs(1879) <= not(layer1_outputs(817));
    layer2_outputs(1880) <= not(layer1_outputs(852)) or (layer1_outputs(1223));
    layer2_outputs(1881) <= not((layer1_outputs(360)) and (layer1_outputs(67)));
    layer2_outputs(1882) <= not(layer1_outputs(2367));
    layer2_outputs(1883) <= '0';
    layer2_outputs(1884) <= not(layer1_outputs(1264));
    layer2_outputs(1885) <= not((layer1_outputs(524)) and (layer1_outputs(1260)));
    layer2_outputs(1886) <= not(layer1_outputs(1423));
    layer2_outputs(1887) <= (layer1_outputs(393)) or (layer1_outputs(2315));
    layer2_outputs(1888) <= (layer1_outputs(1975)) and (layer1_outputs(1337));
    layer2_outputs(1889) <= not((layer1_outputs(1924)) or (layer1_outputs(2048)));
    layer2_outputs(1890) <= not((layer1_outputs(559)) xor (layer1_outputs(1065)));
    layer2_outputs(1891) <= (layer1_outputs(641)) and (layer1_outputs(1834));
    layer2_outputs(1892) <= not((layer1_outputs(2308)) and (layer1_outputs(2410)));
    layer2_outputs(1893) <= '1';
    layer2_outputs(1894) <= '0';
    layer2_outputs(1895) <= not(layer1_outputs(1983)) or (layer1_outputs(1739));
    layer2_outputs(1896) <= '0';
    layer2_outputs(1897) <= not((layer1_outputs(2155)) or (layer1_outputs(1495)));
    layer2_outputs(1898) <= (layer1_outputs(1920)) and not (layer1_outputs(2206));
    layer2_outputs(1899) <= '0';
    layer2_outputs(1900) <= not(layer1_outputs(1250)) or (layer1_outputs(371));
    layer2_outputs(1901) <= layer1_outputs(1560);
    layer2_outputs(1902) <= (layer1_outputs(2033)) and not (layer1_outputs(976));
    layer2_outputs(1903) <= not(layer1_outputs(451)) or (layer1_outputs(2188));
    layer2_outputs(1904) <= (layer1_outputs(1103)) and not (layer1_outputs(700));
    layer2_outputs(1905) <= '1';
    layer2_outputs(1906) <= (layer1_outputs(1769)) and not (layer1_outputs(851));
    layer2_outputs(1907) <= not((layer1_outputs(251)) and (layer1_outputs(823)));
    layer2_outputs(1908) <= not(layer1_outputs(51)) or (layer1_outputs(1562));
    layer2_outputs(1909) <= not(layer1_outputs(1128));
    layer2_outputs(1910) <= not(layer1_outputs(791));
    layer2_outputs(1911) <= (layer1_outputs(326)) and not (layer1_outputs(1762));
    layer2_outputs(1912) <= not((layer1_outputs(1212)) and (layer1_outputs(1554)));
    layer2_outputs(1913) <= (layer1_outputs(2371)) and not (layer1_outputs(1986));
    layer2_outputs(1914) <= (layer1_outputs(1695)) and (layer1_outputs(2120));
    layer2_outputs(1915) <= '0';
    layer2_outputs(1916) <= not(layer1_outputs(56)) or (layer1_outputs(1692));
    layer2_outputs(1917) <= not(layer1_outputs(2446));
    layer2_outputs(1918) <= not((layer1_outputs(1768)) and (layer1_outputs(2385)));
    layer2_outputs(1919) <= layer1_outputs(1310);
    layer2_outputs(1920) <= '1';
    layer2_outputs(1921) <= not(layer1_outputs(1455));
    layer2_outputs(1922) <= '1';
    layer2_outputs(1923) <= not(layer1_outputs(2220));
    layer2_outputs(1924) <= (layer1_outputs(2000)) or (layer1_outputs(1272));
    layer2_outputs(1925) <= not(layer1_outputs(1557));
    layer2_outputs(1926) <= (layer1_outputs(945)) or (layer1_outputs(1750));
    layer2_outputs(1927) <= layer1_outputs(1168);
    layer2_outputs(1928) <= '1';
    layer2_outputs(1929) <= (layer1_outputs(1719)) and not (layer1_outputs(999));
    layer2_outputs(1930) <= not((layer1_outputs(1803)) and (layer1_outputs(2166)));
    layer2_outputs(1931) <= (layer1_outputs(2407)) or (layer1_outputs(2114));
    layer2_outputs(1932) <= not(layer1_outputs(2320));
    layer2_outputs(1933) <= not(layer1_outputs(2439)) or (layer1_outputs(1014));
    layer2_outputs(1934) <= not(layer1_outputs(2262));
    layer2_outputs(1935) <= '0';
    layer2_outputs(1936) <= not(layer1_outputs(857));
    layer2_outputs(1937) <= (layer1_outputs(1285)) and (layer1_outputs(1709));
    layer2_outputs(1938) <= '0';
    layer2_outputs(1939) <= not((layer1_outputs(2318)) or (layer1_outputs(344)));
    layer2_outputs(1940) <= layer1_outputs(1910);
    layer2_outputs(1941) <= (layer1_outputs(2392)) and not (layer1_outputs(623));
    layer2_outputs(1942) <= layer1_outputs(509);
    layer2_outputs(1943) <= '0';
    layer2_outputs(1944) <= '1';
    layer2_outputs(1945) <= (layer1_outputs(423)) xor (layer1_outputs(1460));
    layer2_outputs(1946) <= layer1_outputs(382);
    layer2_outputs(1947) <= not((layer1_outputs(1531)) and (layer1_outputs(2142)));
    layer2_outputs(1948) <= '0';
    layer2_outputs(1949) <= not((layer1_outputs(2006)) and (layer1_outputs(1854)));
    layer2_outputs(1950) <= layer1_outputs(566);
    layer2_outputs(1951) <= '0';
    layer2_outputs(1952) <= not(layer1_outputs(241));
    layer2_outputs(1953) <= (layer1_outputs(1173)) and not (layer1_outputs(23));
    layer2_outputs(1954) <= '0';
    layer2_outputs(1955) <= not(layer1_outputs(365));
    layer2_outputs(1956) <= (layer1_outputs(453)) and (layer1_outputs(1633));
    layer2_outputs(1957) <= '1';
    layer2_outputs(1958) <= not(layer1_outputs(1575));
    layer2_outputs(1959) <= not((layer1_outputs(1505)) or (layer1_outputs(272)));
    layer2_outputs(1960) <= not(layer1_outputs(904));
    layer2_outputs(1961) <= not((layer1_outputs(842)) and (layer1_outputs(2099)));
    layer2_outputs(1962) <= not((layer1_outputs(1152)) and (layer1_outputs(1388)));
    layer2_outputs(1963) <= (layer1_outputs(2276)) and not (layer1_outputs(1158));
    layer2_outputs(1964) <= layer1_outputs(127);
    layer2_outputs(1965) <= (layer1_outputs(1369)) and not (layer1_outputs(889));
    layer2_outputs(1966) <= (layer1_outputs(1703)) and not (layer1_outputs(1513));
    layer2_outputs(1967) <= not((layer1_outputs(1702)) or (layer1_outputs(336)));
    layer2_outputs(1968) <= not(layer1_outputs(561));
    layer2_outputs(1969) <= not(layer1_outputs(1491)) or (layer1_outputs(362));
    layer2_outputs(1970) <= '1';
    layer2_outputs(1971) <= not((layer1_outputs(403)) and (layer1_outputs(856)));
    layer2_outputs(1972) <= layer1_outputs(1329);
    layer2_outputs(1973) <= not(layer1_outputs(51)) or (layer1_outputs(1510));
    layer2_outputs(1974) <= not(layer1_outputs(1533));
    layer2_outputs(1975) <= layer1_outputs(1293);
    layer2_outputs(1976) <= (layer1_outputs(1203)) and not (layer1_outputs(1524));
    layer2_outputs(1977) <= layer1_outputs(1062);
    layer2_outputs(1978) <= not((layer1_outputs(1379)) or (layer1_outputs(1977)));
    layer2_outputs(1979) <= not(layer1_outputs(1748));
    layer2_outputs(1980) <= not(layer1_outputs(1268)) or (layer1_outputs(1432));
    layer2_outputs(1981) <= (layer1_outputs(2199)) or (layer1_outputs(1964));
    layer2_outputs(1982) <= (layer1_outputs(996)) and not (layer1_outputs(2166));
    layer2_outputs(1983) <= layer1_outputs(227);
    layer2_outputs(1984) <= (layer1_outputs(765)) and not (layer1_outputs(26));
    layer2_outputs(1985) <= layer1_outputs(681);
    layer2_outputs(1986) <= (layer1_outputs(2494)) and (layer1_outputs(722));
    layer2_outputs(1987) <= layer1_outputs(433);
    layer2_outputs(1988) <= not((layer1_outputs(422)) or (layer1_outputs(7)));
    layer2_outputs(1989) <= '0';
    layer2_outputs(1990) <= not(layer1_outputs(208));
    layer2_outputs(1991) <= '1';
    layer2_outputs(1992) <= layer1_outputs(2104);
    layer2_outputs(1993) <= not(layer1_outputs(2337));
    layer2_outputs(1994) <= (layer1_outputs(502)) and not (layer1_outputs(78));
    layer2_outputs(1995) <= layer1_outputs(1845);
    layer2_outputs(1996) <= '0';
    layer2_outputs(1997) <= not(layer1_outputs(511)) or (layer1_outputs(896));
    layer2_outputs(1998) <= not(layer1_outputs(2335)) or (layer1_outputs(891));
    layer2_outputs(1999) <= (layer1_outputs(56)) and (layer1_outputs(1880));
    layer2_outputs(2000) <= '1';
    layer2_outputs(2001) <= not((layer1_outputs(902)) and (layer1_outputs(941)));
    layer2_outputs(2002) <= '0';
    layer2_outputs(2003) <= '0';
    layer2_outputs(2004) <= '0';
    layer2_outputs(2005) <= not((layer1_outputs(828)) xor (layer1_outputs(459)));
    layer2_outputs(2006) <= not(layer1_outputs(2456));
    layer2_outputs(2007) <= (layer1_outputs(2406)) or (layer1_outputs(2123));
    layer2_outputs(2008) <= (layer1_outputs(1091)) and not (layer1_outputs(2151));
    layer2_outputs(2009) <= (layer1_outputs(2504)) and (layer1_outputs(610));
    layer2_outputs(2010) <= '0';
    layer2_outputs(2011) <= (layer1_outputs(2206)) and not (layer1_outputs(765));
    layer2_outputs(2012) <= layer1_outputs(2160);
    layer2_outputs(2013) <= not(layer1_outputs(2315));
    layer2_outputs(2014) <= not(layer1_outputs(477));
    layer2_outputs(2015) <= not(layer1_outputs(2539)) or (layer1_outputs(1011));
    layer2_outputs(2016) <= '1';
    layer2_outputs(2017) <= layer1_outputs(677);
    layer2_outputs(2018) <= not(layer1_outputs(1011)) or (layer1_outputs(2192));
    layer2_outputs(2019) <= '0';
    layer2_outputs(2020) <= '1';
    layer2_outputs(2021) <= '0';
    layer2_outputs(2022) <= (layer1_outputs(2019)) and not (layer1_outputs(2268));
    layer2_outputs(2023) <= not(layer1_outputs(2490)) or (layer1_outputs(1077));
    layer2_outputs(2024) <= not((layer1_outputs(1113)) or (layer1_outputs(200)));
    layer2_outputs(2025) <= '0';
    layer2_outputs(2026) <= not(layer1_outputs(450));
    layer2_outputs(2027) <= (layer1_outputs(656)) or (layer1_outputs(1292));
    layer2_outputs(2028) <= '1';
    layer2_outputs(2029) <= not(layer1_outputs(262));
    layer2_outputs(2030) <= '1';
    layer2_outputs(2031) <= layer1_outputs(925);
    layer2_outputs(2032) <= not((layer1_outputs(1085)) or (layer1_outputs(729)));
    layer2_outputs(2033) <= layer1_outputs(1981);
    layer2_outputs(2034) <= '1';
    layer2_outputs(2035) <= not((layer1_outputs(1591)) and (layer1_outputs(216)));
    layer2_outputs(2036) <= not(layer1_outputs(1289)) or (layer1_outputs(2028));
    layer2_outputs(2037) <= (layer1_outputs(397)) and (layer1_outputs(686));
    layer2_outputs(2038) <= '0';
    layer2_outputs(2039) <= not(layer1_outputs(1740)) or (layer1_outputs(1367));
    layer2_outputs(2040) <= not(layer1_outputs(223)) or (layer1_outputs(576));
    layer2_outputs(2041) <= not((layer1_outputs(2137)) or (layer1_outputs(2156)));
    layer2_outputs(2042) <= layer1_outputs(2407);
    layer2_outputs(2043) <= '1';
    layer2_outputs(2044) <= layer1_outputs(513);
    layer2_outputs(2045) <= not(layer1_outputs(170));
    layer2_outputs(2046) <= layer1_outputs(2269);
    layer2_outputs(2047) <= layer1_outputs(2014);
    layer2_outputs(2048) <= not(layer1_outputs(251)) or (layer1_outputs(2489));
    layer2_outputs(2049) <= '0';
    layer2_outputs(2050) <= (layer1_outputs(1887)) and not (layer1_outputs(805));
    layer2_outputs(2051) <= not(layer1_outputs(2422));
    layer2_outputs(2052) <= not(layer1_outputs(2001));
    layer2_outputs(2053) <= not(layer1_outputs(2476));
    layer2_outputs(2054) <= layer1_outputs(1325);
    layer2_outputs(2055) <= not((layer1_outputs(149)) and (layer1_outputs(1080)));
    layer2_outputs(2056) <= (layer1_outputs(2349)) and not (layer1_outputs(1886));
    layer2_outputs(2057) <= (layer1_outputs(427)) or (layer1_outputs(620));
    layer2_outputs(2058) <= not((layer1_outputs(88)) xor (layer1_outputs(1012)));
    layer2_outputs(2059) <= not(layer1_outputs(1611));
    layer2_outputs(2060) <= (layer1_outputs(644)) or (layer1_outputs(855));
    layer2_outputs(2061) <= '0';
    layer2_outputs(2062) <= (layer1_outputs(91)) and (layer1_outputs(1463));
    layer2_outputs(2063) <= layer1_outputs(474);
    layer2_outputs(2064) <= (layer1_outputs(1378)) or (layer1_outputs(158));
    layer2_outputs(2065) <= not(layer1_outputs(803)) or (layer1_outputs(760));
    layer2_outputs(2066) <= (layer1_outputs(1647)) and (layer1_outputs(445));
    layer2_outputs(2067) <= not(layer1_outputs(2108)) or (layer1_outputs(1225));
    layer2_outputs(2068) <= '1';
    layer2_outputs(2069) <= '0';
    layer2_outputs(2070) <= (layer1_outputs(2305)) and not (layer1_outputs(903));
    layer2_outputs(2071) <= not(layer1_outputs(513));
    layer2_outputs(2072) <= not(layer1_outputs(1435));
    layer2_outputs(2073) <= not((layer1_outputs(210)) or (layer1_outputs(1778)));
    layer2_outputs(2074) <= not(layer1_outputs(31)) or (layer1_outputs(474));
    layer2_outputs(2075) <= not(layer1_outputs(901)) or (layer1_outputs(531));
    layer2_outputs(2076) <= not(layer1_outputs(1554));
    layer2_outputs(2077) <= (layer1_outputs(1104)) and not (layer1_outputs(604));
    layer2_outputs(2078) <= '0';
    layer2_outputs(2079) <= not(layer1_outputs(1356)) or (layer1_outputs(1728));
    layer2_outputs(2080) <= not(layer1_outputs(2550));
    layer2_outputs(2081) <= layer1_outputs(2391);
    layer2_outputs(2082) <= '0';
    layer2_outputs(2083) <= layer1_outputs(2091);
    layer2_outputs(2084) <= not(layer1_outputs(1837));
    layer2_outputs(2085) <= not((layer1_outputs(642)) and (layer1_outputs(2479)));
    layer2_outputs(2086) <= (layer1_outputs(73)) and not (layer1_outputs(2345));
    layer2_outputs(2087) <= '1';
    layer2_outputs(2088) <= '0';
    layer2_outputs(2089) <= not(layer1_outputs(2036)) or (layer1_outputs(2441));
    layer2_outputs(2090) <= layer1_outputs(1162);
    layer2_outputs(2091) <= layer1_outputs(548);
    layer2_outputs(2092) <= '0';
    layer2_outputs(2093) <= not(layer1_outputs(1519)) or (layer1_outputs(742));
    layer2_outputs(2094) <= not((layer1_outputs(1224)) and (layer1_outputs(2212)));
    layer2_outputs(2095) <= (layer1_outputs(1129)) and not (layer1_outputs(2158));
    layer2_outputs(2096) <= not(layer1_outputs(525));
    layer2_outputs(2097) <= not((layer1_outputs(1333)) xor (layer1_outputs(2425)));
    layer2_outputs(2098) <= '1';
    layer2_outputs(2099) <= layer1_outputs(2265);
    layer2_outputs(2100) <= '0';
    layer2_outputs(2101) <= '1';
    layer2_outputs(2102) <= not((layer1_outputs(845)) or (layer1_outputs(1664)));
    layer2_outputs(2103) <= (layer1_outputs(916)) and not (layer1_outputs(2203));
    layer2_outputs(2104) <= layer1_outputs(772);
    layer2_outputs(2105) <= not(layer1_outputs(2004));
    layer2_outputs(2106) <= layer1_outputs(573);
    layer2_outputs(2107) <= (layer1_outputs(1460)) or (layer1_outputs(1784));
    layer2_outputs(2108) <= not((layer1_outputs(2508)) and (layer1_outputs(1170)));
    layer2_outputs(2109) <= (layer1_outputs(1026)) and (layer1_outputs(333));
    layer2_outputs(2110) <= not(layer1_outputs(735)) or (layer1_outputs(1610));
    layer2_outputs(2111) <= '1';
    layer2_outputs(2112) <= layer1_outputs(2448);
    layer2_outputs(2113) <= (layer1_outputs(593)) and not (layer1_outputs(9));
    layer2_outputs(2114) <= not((layer1_outputs(2000)) or (layer1_outputs(1517)));
    layer2_outputs(2115) <= not(layer1_outputs(592)) or (layer1_outputs(1766));
    layer2_outputs(2116) <= '1';
    layer2_outputs(2117) <= layer1_outputs(1347);
    layer2_outputs(2118) <= '1';
    layer2_outputs(2119) <= not((layer1_outputs(843)) or (layer1_outputs(1039)));
    layer2_outputs(2120) <= layer1_outputs(1239);
    layer2_outputs(2121) <= layer1_outputs(2243);
    layer2_outputs(2122) <= not(layer1_outputs(519));
    layer2_outputs(2123) <= not(layer1_outputs(1940));
    layer2_outputs(2124) <= layer1_outputs(1890);
    layer2_outputs(2125) <= '0';
    layer2_outputs(2126) <= (layer1_outputs(478)) and (layer1_outputs(621));
    layer2_outputs(2127) <= (layer1_outputs(1439)) and (layer1_outputs(1152));
    layer2_outputs(2128) <= not(layer1_outputs(1747)) or (layer1_outputs(2467));
    layer2_outputs(2129) <= (layer1_outputs(98)) or (layer1_outputs(2350));
    layer2_outputs(2130) <= (layer1_outputs(1519)) or (layer1_outputs(298));
    layer2_outputs(2131) <= (layer1_outputs(2070)) and not (layer1_outputs(1191));
    layer2_outputs(2132) <= not(layer1_outputs(670));
    layer2_outputs(2133) <= not((layer1_outputs(1616)) or (layer1_outputs(1797)));
    layer2_outputs(2134) <= not(layer1_outputs(2062));
    layer2_outputs(2135) <= not(layer1_outputs(1320));
    layer2_outputs(2136) <= not(layer1_outputs(813));
    layer2_outputs(2137) <= '0';
    layer2_outputs(2138) <= (layer1_outputs(1684)) or (layer1_outputs(1526));
    layer2_outputs(2139) <= not(layer1_outputs(2152)) or (layer1_outputs(323));
    layer2_outputs(2140) <= layer1_outputs(1958);
    layer2_outputs(2141) <= '1';
    layer2_outputs(2142) <= layer1_outputs(1535);
    layer2_outputs(2143) <= not(layer1_outputs(1696));
    layer2_outputs(2144) <= layer1_outputs(558);
    layer2_outputs(2145) <= '0';
    layer2_outputs(2146) <= '0';
    layer2_outputs(2147) <= layer1_outputs(2225);
    layer2_outputs(2148) <= not(layer1_outputs(62));
    layer2_outputs(2149) <= not((layer1_outputs(382)) or (layer1_outputs(465)));
    layer2_outputs(2150) <= '1';
    layer2_outputs(2151) <= not(layer1_outputs(1021));
    layer2_outputs(2152) <= layer1_outputs(735);
    layer2_outputs(2153) <= not(layer1_outputs(304));
    layer2_outputs(2154) <= layer1_outputs(1622);
    layer2_outputs(2155) <= not(layer1_outputs(577)) or (layer1_outputs(127));
    layer2_outputs(2156) <= (layer1_outputs(1336)) and not (layer1_outputs(1433));
    layer2_outputs(2157) <= not((layer1_outputs(1885)) or (layer1_outputs(318)));
    layer2_outputs(2158) <= not(layer1_outputs(1036)) or (layer1_outputs(2424));
    layer2_outputs(2159) <= not(layer1_outputs(57)) or (layer1_outputs(1732));
    layer2_outputs(2160) <= not(layer1_outputs(270));
    layer2_outputs(2161) <= not(layer1_outputs(2487)) or (layer1_outputs(288));
    layer2_outputs(2162) <= (layer1_outputs(195)) and not (layer1_outputs(1160));
    layer2_outputs(2163) <= layer1_outputs(749);
    layer2_outputs(2164) <= not(layer1_outputs(526));
    layer2_outputs(2165) <= not((layer1_outputs(337)) or (layer1_outputs(539)));
    layer2_outputs(2166) <= layer1_outputs(2043);
    layer2_outputs(2167) <= layer1_outputs(2018);
    layer2_outputs(2168) <= not(layer1_outputs(1383));
    layer2_outputs(2169) <= layer1_outputs(2210);
    layer2_outputs(2170) <= not((layer1_outputs(628)) and (layer1_outputs(1237)));
    layer2_outputs(2171) <= '0';
    layer2_outputs(2172) <= (layer1_outputs(1677)) or (layer1_outputs(1653));
    layer2_outputs(2173) <= layer1_outputs(380);
    layer2_outputs(2174) <= '1';
    layer2_outputs(2175) <= layer1_outputs(1598);
    layer2_outputs(2176) <= layer1_outputs(2297);
    layer2_outputs(2177) <= not(layer1_outputs(480));
    layer2_outputs(2178) <= (layer1_outputs(939)) and not (layer1_outputs(1556));
    layer2_outputs(2179) <= (layer1_outputs(695)) and not (layer1_outputs(1146));
    layer2_outputs(2180) <= (layer1_outputs(1902)) and (layer1_outputs(2375));
    layer2_outputs(2181) <= '0';
    layer2_outputs(2182) <= not(layer1_outputs(406)) or (layer1_outputs(1736));
    layer2_outputs(2183) <= '1';
    layer2_outputs(2184) <= not(layer1_outputs(1791));
    layer2_outputs(2185) <= '0';
    layer2_outputs(2186) <= layer1_outputs(69);
    layer2_outputs(2187) <= layer1_outputs(2090);
    layer2_outputs(2188) <= '1';
    layer2_outputs(2189) <= (layer1_outputs(1708)) or (layer1_outputs(1165));
    layer2_outputs(2190) <= not(layer1_outputs(1654)) or (layer1_outputs(970));
    layer2_outputs(2191) <= '0';
    layer2_outputs(2192) <= not(layer1_outputs(777)) or (layer1_outputs(1231));
    layer2_outputs(2193) <= '1';
    layer2_outputs(2194) <= layer1_outputs(1776);
    layer2_outputs(2195) <= '0';
    layer2_outputs(2196) <= '0';
    layer2_outputs(2197) <= layer1_outputs(1049);
    layer2_outputs(2198) <= '1';
    layer2_outputs(2199) <= '0';
    layer2_outputs(2200) <= layer1_outputs(1882);
    layer2_outputs(2201) <= layer1_outputs(2092);
    layer2_outputs(2202) <= not((layer1_outputs(2174)) xor (layer1_outputs(1308)));
    layer2_outputs(2203) <= not((layer1_outputs(1497)) and (layer1_outputs(2291)));
    layer2_outputs(2204) <= not((layer1_outputs(2211)) and (layer1_outputs(2066)));
    layer2_outputs(2205) <= layer1_outputs(101);
    layer2_outputs(2206) <= layer1_outputs(1785);
    layer2_outputs(2207) <= '1';
    layer2_outputs(2208) <= not(layer1_outputs(2484));
    layer2_outputs(2209) <= (layer1_outputs(69)) and not (layer1_outputs(16));
    layer2_outputs(2210) <= (layer1_outputs(188)) and (layer1_outputs(1802));
    layer2_outputs(2211) <= layer1_outputs(1816);
    layer2_outputs(2212) <= (layer1_outputs(2353)) and not (layer1_outputs(1511));
    layer2_outputs(2213) <= not(layer1_outputs(2218)) or (layer1_outputs(1815));
    layer2_outputs(2214) <= '1';
    layer2_outputs(2215) <= (layer1_outputs(1228)) and not (layer1_outputs(1019));
    layer2_outputs(2216) <= not((layer1_outputs(1222)) or (layer1_outputs(1199)));
    layer2_outputs(2217) <= not(layer1_outputs(2377)) or (layer1_outputs(2267));
    layer2_outputs(2218) <= not(layer1_outputs(767)) or (layer1_outputs(741));
    layer2_outputs(2219) <= not(layer1_outputs(1039));
    layer2_outputs(2220) <= not(layer1_outputs(201));
    layer2_outputs(2221) <= '1';
    layer2_outputs(2222) <= (layer1_outputs(1908)) or (layer1_outputs(341));
    layer2_outputs(2223) <= not(layer1_outputs(389));
    layer2_outputs(2224) <= layer1_outputs(113);
    layer2_outputs(2225) <= not(layer1_outputs(2401));
    layer2_outputs(2226) <= (layer1_outputs(3)) or (layer1_outputs(1924));
    layer2_outputs(2227) <= '1';
    layer2_outputs(2228) <= not(layer1_outputs(1972)) or (layer1_outputs(1240));
    layer2_outputs(2229) <= (layer1_outputs(1480)) and (layer1_outputs(1804));
    layer2_outputs(2230) <= not(layer1_outputs(1495)) or (layer1_outputs(1923));
    layer2_outputs(2231) <= layer1_outputs(1161);
    layer2_outputs(2232) <= not(layer1_outputs(57));
    layer2_outputs(2233) <= '0';
    layer2_outputs(2234) <= not((layer1_outputs(324)) or (layer1_outputs(1694)));
    layer2_outputs(2235) <= layer1_outputs(1798);
    layer2_outputs(2236) <= '0';
    layer2_outputs(2237) <= layer1_outputs(2335);
    layer2_outputs(2238) <= not(layer1_outputs(1919)) or (layer1_outputs(994));
    layer2_outputs(2239) <= '0';
    layer2_outputs(2240) <= '0';
    layer2_outputs(2241) <= layer1_outputs(899);
    layer2_outputs(2242) <= (layer1_outputs(1116)) and not (layer1_outputs(882));
    layer2_outputs(2243) <= (layer1_outputs(2408)) or (layer1_outputs(774));
    layer2_outputs(2244) <= not((layer1_outputs(1257)) or (layer1_outputs(517)));
    layer2_outputs(2245) <= not(layer1_outputs(2295));
    layer2_outputs(2246) <= (layer1_outputs(2113)) and (layer1_outputs(427));
    layer2_outputs(2247) <= '1';
    layer2_outputs(2248) <= '0';
    layer2_outputs(2249) <= layer1_outputs(2279);
    layer2_outputs(2250) <= '1';
    layer2_outputs(2251) <= (layer1_outputs(2199)) or (layer1_outputs(612));
    layer2_outputs(2252) <= (layer1_outputs(732)) and not (layer1_outputs(253));
    layer2_outputs(2253) <= (layer1_outputs(2147)) or (layer1_outputs(608));
    layer2_outputs(2254) <= (layer1_outputs(1596)) and not (layer1_outputs(1404));
    layer2_outputs(2255) <= not(layer1_outputs(1211));
    layer2_outputs(2256) <= (layer1_outputs(595)) and (layer1_outputs(707));
    layer2_outputs(2257) <= not((layer1_outputs(1006)) and (layer1_outputs(761)));
    layer2_outputs(2258) <= '0';
    layer2_outputs(2259) <= not((layer1_outputs(1870)) or (layer1_outputs(277)));
    layer2_outputs(2260) <= not((layer1_outputs(1766)) and (layer1_outputs(1358)));
    layer2_outputs(2261) <= layer1_outputs(2196);
    layer2_outputs(2262) <= not((layer1_outputs(2411)) or (layer1_outputs(747)));
    layer2_outputs(2263) <= (layer1_outputs(1056)) and (layer1_outputs(1933));
    layer2_outputs(2264) <= not(layer1_outputs(666));
    layer2_outputs(2265) <= not(layer1_outputs(2115)) or (layer1_outputs(1066));
    layer2_outputs(2266) <= (layer1_outputs(1571)) and not (layer1_outputs(2273));
    layer2_outputs(2267) <= not(layer1_outputs(273));
    layer2_outputs(2268) <= '0';
    layer2_outputs(2269) <= not(layer1_outputs(70));
    layer2_outputs(2270) <= layer1_outputs(521);
    layer2_outputs(2271) <= not(layer1_outputs(2394));
    layer2_outputs(2272) <= not(layer1_outputs(495)) or (layer1_outputs(1687));
    layer2_outputs(2273) <= (layer1_outputs(2409)) and (layer1_outputs(279));
    layer2_outputs(2274) <= (layer1_outputs(873)) and not (layer1_outputs(371));
    layer2_outputs(2275) <= layer1_outputs(34);
    layer2_outputs(2276) <= not(layer1_outputs(669));
    layer2_outputs(2277) <= '0';
    layer2_outputs(2278) <= layer1_outputs(1561);
    layer2_outputs(2279) <= not((layer1_outputs(1292)) or (layer1_outputs(1192)));
    layer2_outputs(2280) <= not(layer1_outputs(2408));
    layer2_outputs(2281) <= (layer1_outputs(1320)) or (layer1_outputs(1112));
    layer2_outputs(2282) <= (layer1_outputs(2045)) and (layer1_outputs(1572));
    layer2_outputs(2283) <= '1';
    layer2_outputs(2284) <= layer1_outputs(886);
    layer2_outputs(2285) <= (layer1_outputs(570)) and not (layer1_outputs(824));
    layer2_outputs(2286) <= (layer1_outputs(1796)) and not (layer1_outputs(1561));
    layer2_outputs(2287) <= '0';
    layer2_outputs(2288) <= '1';
    layer2_outputs(2289) <= layer1_outputs(120);
    layer2_outputs(2290) <= not(layer1_outputs(951)) or (layer1_outputs(1757));
    layer2_outputs(2291) <= not(layer1_outputs(961));
    layer2_outputs(2292) <= '1';
    layer2_outputs(2293) <= (layer1_outputs(1478)) or (layer1_outputs(48));
    layer2_outputs(2294) <= not(layer1_outputs(1398)) or (layer1_outputs(619));
    layer2_outputs(2295) <= (layer1_outputs(616)) and not (layer1_outputs(2453));
    layer2_outputs(2296) <= (layer1_outputs(1876)) and not (layer1_outputs(1133));
    layer2_outputs(2297) <= not(layer1_outputs(1074));
    layer2_outputs(2298) <= layer1_outputs(1958);
    layer2_outputs(2299) <= not(layer1_outputs(1390));
    layer2_outputs(2300) <= '1';
    layer2_outputs(2301) <= layer1_outputs(1157);
    layer2_outputs(2302) <= not((layer1_outputs(72)) and (layer1_outputs(2531)));
    layer2_outputs(2303) <= not(layer1_outputs(172)) or (layer1_outputs(1515));
    layer2_outputs(2304) <= (layer1_outputs(1916)) and not (layer1_outputs(726));
    layer2_outputs(2305) <= layer1_outputs(496);
    layer2_outputs(2306) <= '1';
    layer2_outputs(2307) <= layer1_outputs(301);
    layer2_outputs(2308) <= (layer1_outputs(869)) and not (layer1_outputs(307));
    layer2_outputs(2309) <= '0';
    layer2_outputs(2310) <= (layer1_outputs(2161)) and not (layer1_outputs(1398));
    layer2_outputs(2311) <= layer1_outputs(1381);
    layer2_outputs(2312) <= '1';
    layer2_outputs(2313) <= (layer1_outputs(1033)) and not (layer1_outputs(2485));
    layer2_outputs(2314) <= not(layer1_outputs(1852));
    layer2_outputs(2315) <= not(layer1_outputs(103)) or (layer1_outputs(2022));
    layer2_outputs(2316) <= (layer1_outputs(685)) and (layer1_outputs(2432));
    layer2_outputs(2317) <= (layer1_outputs(2363)) and (layer1_outputs(2466));
    layer2_outputs(2318) <= not(layer1_outputs(2447));
    layer2_outputs(2319) <= '0';
    layer2_outputs(2320) <= not(layer1_outputs(291));
    layer2_outputs(2321) <= '1';
    layer2_outputs(2322) <= '1';
    layer2_outputs(2323) <= '0';
    layer2_outputs(2324) <= '0';
    layer2_outputs(2325) <= not(layer1_outputs(327));
    layer2_outputs(2326) <= (layer1_outputs(139)) and not (layer1_outputs(500));
    layer2_outputs(2327) <= (layer1_outputs(1140)) and not (layer1_outputs(2084));
    layer2_outputs(2328) <= not(layer1_outputs(1456)) or (layer1_outputs(104));
    layer2_outputs(2329) <= not(layer1_outputs(1164));
    layer2_outputs(2330) <= (layer1_outputs(1055)) and (layer1_outputs(2475));
    layer2_outputs(2331) <= not((layer1_outputs(281)) or (layer1_outputs(1846)));
    layer2_outputs(2332) <= (layer1_outputs(1829)) and (layer1_outputs(652));
    layer2_outputs(2333) <= not(layer1_outputs(89)) or (layer1_outputs(2306));
    layer2_outputs(2334) <= (layer1_outputs(2052)) or (layer1_outputs(992));
    layer2_outputs(2335) <= layer1_outputs(326);
    layer2_outputs(2336) <= (layer1_outputs(1127)) and (layer1_outputs(2418));
    layer2_outputs(2337) <= (layer1_outputs(1245)) and not (layer1_outputs(2467));
    layer2_outputs(2338) <= layer1_outputs(2556);
    layer2_outputs(2339) <= not(layer1_outputs(1586));
    layer2_outputs(2340) <= not(layer1_outputs(646));
    layer2_outputs(2341) <= layer1_outputs(2458);
    layer2_outputs(2342) <= (layer1_outputs(1023)) or (layer1_outputs(560));
    layer2_outputs(2343) <= (layer1_outputs(809)) or (layer1_outputs(877));
    layer2_outputs(2344) <= layer1_outputs(2522);
    layer2_outputs(2345) <= layer1_outputs(1828);
    layer2_outputs(2346) <= not((layer1_outputs(875)) and (layer1_outputs(1711)));
    layer2_outputs(2347) <= (layer1_outputs(2361)) and not (layer1_outputs(218));
    layer2_outputs(2348) <= layer1_outputs(711);
    layer2_outputs(2349) <= not((layer1_outputs(1116)) and (layer1_outputs(1054)));
    layer2_outputs(2350) <= '0';
    layer2_outputs(2351) <= (layer1_outputs(2323)) and (layer1_outputs(384));
    layer2_outputs(2352) <= (layer1_outputs(2471)) or (layer1_outputs(325));
    layer2_outputs(2353) <= not(layer1_outputs(2258));
    layer2_outputs(2354) <= not((layer1_outputs(2341)) xor (layer1_outputs(2538)));
    layer2_outputs(2355) <= not((layer1_outputs(99)) and (layer1_outputs(567)));
    layer2_outputs(2356) <= layer1_outputs(183);
    layer2_outputs(2357) <= (layer1_outputs(950)) and not (layer1_outputs(443));
    layer2_outputs(2358) <= layer1_outputs(1937);
    layer2_outputs(2359) <= '1';
    layer2_outputs(2360) <= not((layer1_outputs(88)) and (layer1_outputs(1601)));
    layer2_outputs(2361) <= not((layer1_outputs(1407)) or (layer1_outputs(2502)));
    layer2_outputs(2362) <= not(layer1_outputs(1934));
    layer2_outputs(2363) <= not(layer1_outputs(820));
    layer2_outputs(2364) <= not(layer1_outputs(2346));
    layer2_outputs(2365) <= not((layer1_outputs(931)) or (layer1_outputs(2083)));
    layer2_outputs(2366) <= not(layer1_outputs(618)) or (layer1_outputs(345));
    layer2_outputs(2367) <= '0';
    layer2_outputs(2368) <= (layer1_outputs(148)) and not (layer1_outputs(248));
    layer2_outputs(2369) <= layer1_outputs(562);
    layer2_outputs(2370) <= not(layer1_outputs(1507));
    layer2_outputs(2371) <= not((layer1_outputs(535)) or (layer1_outputs(126)));
    layer2_outputs(2372) <= '1';
    layer2_outputs(2373) <= not((layer1_outputs(927)) and (layer1_outputs(511)));
    layer2_outputs(2374) <= not((layer1_outputs(1230)) and (layer1_outputs(462)));
    layer2_outputs(2375) <= (layer1_outputs(2197)) or (layer1_outputs(2080));
    layer2_outputs(2376) <= '1';
    layer2_outputs(2377) <= not(layer1_outputs(330));
    layer2_outputs(2378) <= (layer1_outputs(2292)) and not (layer1_outputs(983));
    layer2_outputs(2379) <= (layer1_outputs(1817)) and not (layer1_outputs(572));
    layer2_outputs(2380) <= '0';
    layer2_outputs(2381) <= not(layer1_outputs(1106));
    layer2_outputs(2382) <= not(layer1_outputs(132)) or (layer1_outputs(654));
    layer2_outputs(2383) <= (layer1_outputs(1008)) or (layer1_outputs(138));
    layer2_outputs(2384) <= (layer1_outputs(2505)) and not (layer1_outputs(589));
    layer2_outputs(2385) <= not(layer1_outputs(751));
    layer2_outputs(2386) <= not((layer1_outputs(1197)) and (layer1_outputs(14)));
    layer2_outputs(2387) <= (layer1_outputs(1462)) and (layer1_outputs(1483));
    layer2_outputs(2388) <= not((layer1_outputs(1005)) xor (layer1_outputs(1671)));
    layer2_outputs(2389) <= not((layer1_outputs(434)) and (layer1_outputs(821)));
    layer2_outputs(2390) <= (layer1_outputs(1359)) and not (layer1_outputs(1748));
    layer2_outputs(2391) <= '0';
    layer2_outputs(2392) <= '0';
    layer2_outputs(2393) <= (layer1_outputs(2071)) and not (layer1_outputs(2468));
    layer2_outputs(2394) <= not(layer1_outputs(1648)) or (layer1_outputs(83));
    layer2_outputs(2395) <= not(layer1_outputs(1718)) or (layer1_outputs(746));
    layer2_outputs(2396) <= layer1_outputs(291);
    layer2_outputs(2397) <= (layer1_outputs(1384)) and not (layer1_outputs(1034));
    layer2_outputs(2398) <= not(layer1_outputs(2002)) or (layer1_outputs(201));
    layer2_outputs(2399) <= not((layer1_outputs(1141)) or (layer1_outputs(2300)));
    layer2_outputs(2400) <= not(layer1_outputs(1401));
    layer2_outputs(2401) <= '0';
    layer2_outputs(2402) <= (layer1_outputs(1749)) or (layer1_outputs(2126));
    layer2_outputs(2403) <= not((layer1_outputs(132)) and (layer1_outputs(1681)));
    layer2_outputs(2404) <= '0';
    layer2_outputs(2405) <= not((layer1_outputs(1896)) and (layer1_outputs(763)));
    layer2_outputs(2406) <= layer1_outputs(437);
    layer2_outputs(2407) <= layer1_outputs(1649);
    layer2_outputs(2408) <= layer1_outputs(995);
    layer2_outputs(2409) <= not((layer1_outputs(2063)) or (layer1_outputs(1521)));
    layer2_outputs(2410) <= layer1_outputs(2138);
    layer2_outputs(2411) <= not(layer1_outputs(2236)) or (layer1_outputs(1829));
    layer2_outputs(2412) <= not(layer1_outputs(786));
    layer2_outputs(2413) <= (layer1_outputs(2460)) and (layer1_outputs(1458));
    layer2_outputs(2414) <= layer1_outputs(651);
    layer2_outputs(2415) <= not(layer1_outputs(2232)) or (layer1_outputs(1547));
    layer2_outputs(2416) <= (layer1_outputs(1018)) and not (layer1_outputs(879));
    layer2_outputs(2417) <= (layer1_outputs(522)) and (layer1_outputs(186));
    layer2_outputs(2418) <= (layer1_outputs(2304)) and not (layer1_outputs(1027));
    layer2_outputs(2419) <= not((layer1_outputs(2256)) or (layer1_outputs(1782)));
    layer2_outputs(2420) <= (layer1_outputs(366)) or (layer1_outputs(1267));
    layer2_outputs(2421) <= (layer1_outputs(207)) and (layer1_outputs(2520));
    layer2_outputs(2422) <= not(layer1_outputs(693)) or (layer1_outputs(1838));
    layer2_outputs(2423) <= '0';
    layer2_outputs(2424) <= layer1_outputs(206);
    layer2_outputs(2425) <= not(layer1_outputs(2484));
    layer2_outputs(2426) <= (layer1_outputs(2257)) and (layer1_outputs(2304));
    layer2_outputs(2427) <= layer1_outputs(551);
    layer2_outputs(2428) <= not(layer1_outputs(1153));
    layer2_outputs(2429) <= (layer1_outputs(1344)) and not (layer1_outputs(1043));
    layer2_outputs(2430) <= not((layer1_outputs(531)) or (layer1_outputs(804)));
    layer2_outputs(2431) <= (layer1_outputs(245)) and not (layer1_outputs(1470));
    layer2_outputs(2432) <= '0';
    layer2_outputs(2433) <= not(layer1_outputs(2512));
    layer2_outputs(2434) <= not(layer1_outputs(1600)) or (layer1_outputs(2135));
    layer2_outputs(2435) <= '0';
    layer2_outputs(2436) <= (layer1_outputs(1592)) and (layer1_outputs(1805));
    layer2_outputs(2437) <= (layer1_outputs(2039)) and not (layer1_outputs(988));
    layer2_outputs(2438) <= not(layer1_outputs(2173));
    layer2_outputs(2439) <= not(layer1_outputs(2081)) or (layer1_outputs(821));
    layer2_outputs(2440) <= layer1_outputs(1418);
    layer2_outputs(2441) <= '1';
    layer2_outputs(2442) <= '0';
    layer2_outputs(2443) <= not((layer1_outputs(690)) and (layer1_outputs(856)));
    layer2_outputs(2444) <= not(layer1_outputs(2521));
    layer2_outputs(2445) <= not(layer1_outputs(2023)) or (layer1_outputs(1411));
    layer2_outputs(2446) <= not(layer1_outputs(2506));
    layer2_outputs(2447) <= (layer1_outputs(1430)) and not (layer1_outputs(2332));
    layer2_outputs(2448) <= '1';
    layer2_outputs(2449) <= '0';
    layer2_outputs(2450) <= layer1_outputs(1266);
    layer2_outputs(2451) <= not((layer1_outputs(2056)) or (layer1_outputs(835)));
    layer2_outputs(2452) <= layer1_outputs(1877);
    layer2_outputs(2453) <= '0';
    layer2_outputs(2454) <= not((layer1_outputs(963)) or (layer1_outputs(163)));
    layer2_outputs(2455) <= (layer1_outputs(332)) and not (layer1_outputs(2017));
    layer2_outputs(2456) <= '0';
    layer2_outputs(2457) <= (layer1_outputs(2310)) or (layer1_outputs(0));
    layer2_outputs(2458) <= not(layer1_outputs(454)) or (layer1_outputs(2175));
    layer2_outputs(2459) <= not(layer1_outputs(1535)) or (layer1_outputs(1033));
    layer2_outputs(2460) <= layer1_outputs(2282);
    layer2_outputs(2461) <= not(layer1_outputs(349)) or (layer1_outputs(231));
    layer2_outputs(2462) <= '0';
    layer2_outputs(2463) <= layer1_outputs(953);
    layer2_outputs(2464) <= (layer1_outputs(1169)) and not (layer1_outputs(1454));
    layer2_outputs(2465) <= not((layer1_outputs(1074)) or (layer1_outputs(697)));
    layer2_outputs(2466) <= '0';
    layer2_outputs(2467) <= not(layer1_outputs(296)) or (layer1_outputs(407));
    layer2_outputs(2468) <= '1';
    layer2_outputs(2469) <= '1';
    layer2_outputs(2470) <= (layer1_outputs(855)) and (layer1_outputs(1207));
    layer2_outputs(2471) <= (layer1_outputs(335)) and not (layer1_outputs(862));
    layer2_outputs(2472) <= '1';
    layer2_outputs(2473) <= not(layer1_outputs(130)) or (layer1_outputs(1884));
    layer2_outputs(2474) <= (layer1_outputs(1624)) and not (layer1_outputs(229));
    layer2_outputs(2475) <= (layer1_outputs(2193)) and (layer1_outputs(172));
    layer2_outputs(2476) <= not(layer1_outputs(1357)) or (layer1_outputs(2559));
    layer2_outputs(2477) <= (layer1_outputs(489)) and not (layer1_outputs(2370));
    layer2_outputs(2478) <= (layer1_outputs(468)) and not (layer1_outputs(136));
    layer2_outputs(2479) <= not(layer1_outputs(728)) or (layer1_outputs(1089));
    layer2_outputs(2480) <= not(layer1_outputs(1783));
    layer2_outputs(2481) <= (layer1_outputs(1345)) and (layer1_outputs(518));
    layer2_outputs(2482) <= (layer1_outputs(425)) and not (layer1_outputs(1668));
    layer2_outputs(2483) <= (layer1_outputs(1149)) and (layer1_outputs(2350));
    layer2_outputs(2484) <= not(layer1_outputs(947)) or (layer1_outputs(2046));
    layer2_outputs(2485) <= not((layer1_outputs(544)) and (layer1_outputs(221)));
    layer2_outputs(2486) <= not((layer1_outputs(1550)) or (layer1_outputs(1610)));
    layer2_outputs(2487) <= layer1_outputs(1254);
    layer2_outputs(2488) <= (layer1_outputs(1414)) and (layer1_outputs(495));
    layer2_outputs(2489) <= not((layer1_outputs(1954)) and (layer1_outputs(1970)));
    layer2_outputs(2490) <= '1';
    layer2_outputs(2491) <= (layer1_outputs(265)) xor (layer1_outputs(1779));
    layer2_outputs(2492) <= not((layer1_outputs(1190)) and (layer1_outputs(2035)));
    layer2_outputs(2493) <= '1';
    layer2_outputs(2494) <= '1';
    layer2_outputs(2495) <= not(layer1_outputs(930)) or (layer1_outputs(2357));
    layer2_outputs(2496) <= not((layer1_outputs(230)) and (layer1_outputs(2233)));
    layer2_outputs(2497) <= (layer1_outputs(782)) and not (layer1_outputs(1446));
    layer2_outputs(2498) <= '1';
    layer2_outputs(2499) <= not(layer1_outputs(2508));
    layer2_outputs(2500) <= (layer1_outputs(1268)) and not (layer1_outputs(2216));
    layer2_outputs(2501) <= not(layer1_outputs(1296));
    layer2_outputs(2502) <= not(layer1_outputs(394)) or (layer1_outputs(801));
    layer2_outputs(2503) <= not((layer1_outputs(375)) and (layer1_outputs(1827)));
    layer2_outputs(2504) <= not((layer1_outputs(339)) and (layer1_outputs(214)));
    layer2_outputs(2505) <= not(layer1_outputs(146));
    layer2_outputs(2506) <= '1';
    layer2_outputs(2507) <= '0';
    layer2_outputs(2508) <= layer1_outputs(2515);
    layer2_outputs(2509) <= (layer1_outputs(231)) and not (layer1_outputs(983));
    layer2_outputs(2510) <= not((layer1_outputs(278)) xor (layer1_outputs(1837)));
    layer2_outputs(2511) <= '0';
    layer2_outputs(2512) <= (layer1_outputs(987)) or (layer1_outputs(1476));
    layer2_outputs(2513) <= not(layer1_outputs(1712)) or (layer1_outputs(82));
    layer2_outputs(2514) <= not(layer1_outputs(2426));
    layer2_outputs(2515) <= (layer1_outputs(2042)) and (layer1_outputs(209));
    layer2_outputs(2516) <= layer1_outputs(2233);
    layer2_outputs(2517) <= not(layer1_outputs(2143)) or (layer1_outputs(232));
    layer2_outputs(2518) <= layer1_outputs(1455);
    layer2_outputs(2519) <= not(layer1_outputs(266)) or (layer1_outputs(2559));
    layer2_outputs(2520) <= (layer1_outputs(1515)) and not (layer1_outputs(1675));
    layer2_outputs(2521) <= not(layer1_outputs(2317));
    layer2_outputs(2522) <= not(layer1_outputs(492)) or (layer1_outputs(2417));
    layer2_outputs(2523) <= not(layer1_outputs(447)) or (layer1_outputs(705));
    layer2_outputs(2524) <= not((layer1_outputs(1248)) xor (layer1_outputs(1720)));
    layer2_outputs(2525) <= not((layer1_outputs(1663)) and (layer1_outputs(1889)));
    layer2_outputs(2526) <= not(layer1_outputs(1191));
    layer2_outputs(2527) <= not((layer1_outputs(685)) or (layer1_outputs(1370)));
    layer2_outputs(2528) <= (layer1_outputs(1192)) and (layer1_outputs(908));
    layer2_outputs(2529) <= not(layer1_outputs(1172));
    layer2_outputs(2530) <= '1';
    layer2_outputs(2531) <= '0';
    layer2_outputs(2532) <= (layer1_outputs(1315)) and (layer1_outputs(74));
    layer2_outputs(2533) <= (layer1_outputs(1533)) and (layer1_outputs(318));
    layer2_outputs(2534) <= (layer1_outputs(1563)) and not (layer1_outputs(1295));
    layer2_outputs(2535) <= not(layer1_outputs(834)) or (layer1_outputs(243));
    layer2_outputs(2536) <= not((layer1_outputs(308)) or (layer1_outputs(2347)));
    layer2_outputs(2537) <= (layer1_outputs(654)) and not (layer1_outputs(2021));
    layer2_outputs(2538) <= not(layer1_outputs(990)) or (layer1_outputs(483));
    layer2_outputs(2539) <= not((layer1_outputs(2321)) or (layer1_outputs(187)));
    layer2_outputs(2540) <= not((layer1_outputs(1075)) or (layer1_outputs(306)));
    layer2_outputs(2541) <= not(layer1_outputs(846));
    layer2_outputs(2542) <= (layer1_outputs(2072)) and not (layer1_outputs(1500));
    layer2_outputs(2543) <= layer1_outputs(1754);
    layer2_outputs(2544) <= not(layer1_outputs(2347));
    layer2_outputs(2545) <= layer1_outputs(1843);
    layer2_outputs(2546) <= (layer1_outputs(436)) and (layer1_outputs(841));
    layer2_outputs(2547) <= layer1_outputs(2007);
    layer2_outputs(2548) <= not(layer1_outputs(2360));
    layer2_outputs(2549) <= (layer1_outputs(2355)) and not (layer1_outputs(1262));
    layer2_outputs(2550) <= not(layer1_outputs(2494));
    layer2_outputs(2551) <= (layer1_outputs(1874)) and not (layer1_outputs(289));
    layer2_outputs(2552) <= not((layer1_outputs(2452)) and (layer1_outputs(212)));
    layer2_outputs(2553) <= '0';
    layer2_outputs(2554) <= layer1_outputs(1269);
    layer2_outputs(2555) <= layer1_outputs(24);
    layer2_outputs(2556) <= not(layer1_outputs(1534));
    layer2_outputs(2557) <= (layer1_outputs(2177)) and not (layer1_outputs(1402));
    layer2_outputs(2558) <= (layer1_outputs(655)) and not (layer1_outputs(29));
    layer2_outputs(2559) <= not(layer1_outputs(157));
    layer3_outputs(0) <= layer2_outputs(2257);
    layer3_outputs(1) <= not((layer2_outputs(1238)) or (layer2_outputs(1765)));
    layer3_outputs(2) <= not(layer2_outputs(1289)) or (layer2_outputs(412));
    layer3_outputs(3) <= '0';
    layer3_outputs(4) <= not(layer2_outputs(1452));
    layer3_outputs(5) <= (layer2_outputs(1621)) or (layer2_outputs(2307));
    layer3_outputs(6) <= not(layer2_outputs(2177));
    layer3_outputs(7) <= not(layer2_outputs(1448)) or (layer2_outputs(1253));
    layer3_outputs(8) <= not((layer2_outputs(2265)) and (layer2_outputs(329)));
    layer3_outputs(9) <= not((layer2_outputs(925)) and (layer2_outputs(970)));
    layer3_outputs(10) <= not(layer2_outputs(1247));
    layer3_outputs(11) <= not((layer2_outputs(861)) xor (layer2_outputs(844)));
    layer3_outputs(12) <= not(layer2_outputs(1636));
    layer3_outputs(13) <= (layer2_outputs(87)) or (layer2_outputs(789));
    layer3_outputs(14) <= layer2_outputs(2048);
    layer3_outputs(15) <= '0';
    layer3_outputs(16) <= '1';
    layer3_outputs(17) <= '0';
    layer3_outputs(18) <= (layer2_outputs(627)) and not (layer2_outputs(1614));
    layer3_outputs(19) <= not(layer2_outputs(2086)) or (layer2_outputs(243));
    layer3_outputs(20) <= layer2_outputs(1995);
    layer3_outputs(21) <= not((layer2_outputs(1754)) and (layer2_outputs(1985)));
    layer3_outputs(22) <= (layer2_outputs(1492)) and not (layer2_outputs(945));
    layer3_outputs(23) <= (layer2_outputs(859)) and not (layer2_outputs(63));
    layer3_outputs(24) <= '1';
    layer3_outputs(25) <= layer2_outputs(2495);
    layer3_outputs(26) <= layer2_outputs(930);
    layer3_outputs(27) <= not(layer2_outputs(2545)) or (layer2_outputs(788));
    layer3_outputs(28) <= not(layer2_outputs(2070));
    layer3_outputs(29) <= (layer2_outputs(2170)) xor (layer2_outputs(2008));
    layer3_outputs(30) <= not(layer2_outputs(697)) or (layer2_outputs(1865));
    layer3_outputs(31) <= not(layer2_outputs(2071)) or (layer2_outputs(1054));
    layer3_outputs(32) <= not((layer2_outputs(334)) and (layer2_outputs(1442)));
    layer3_outputs(33) <= layer2_outputs(1320);
    layer3_outputs(34) <= not((layer2_outputs(1956)) and (layer2_outputs(252)));
    layer3_outputs(35) <= layer2_outputs(1443);
    layer3_outputs(36) <= not((layer2_outputs(2546)) or (layer2_outputs(237)));
    layer3_outputs(37) <= (layer2_outputs(2084)) and not (layer2_outputs(238));
    layer3_outputs(38) <= '1';
    layer3_outputs(39) <= not(layer2_outputs(290)) or (layer2_outputs(1095));
    layer3_outputs(40) <= '1';
    layer3_outputs(41) <= not(layer2_outputs(1973)) or (layer2_outputs(256));
    layer3_outputs(42) <= not(layer2_outputs(2096));
    layer3_outputs(43) <= not(layer2_outputs(355)) or (layer2_outputs(1474));
    layer3_outputs(44) <= not(layer2_outputs(2072));
    layer3_outputs(45) <= not(layer2_outputs(2094));
    layer3_outputs(46) <= not((layer2_outputs(1662)) and (layer2_outputs(69)));
    layer3_outputs(47) <= layer2_outputs(1607);
    layer3_outputs(48) <= not(layer2_outputs(929));
    layer3_outputs(49) <= (layer2_outputs(1144)) and (layer2_outputs(2452));
    layer3_outputs(50) <= not(layer2_outputs(2139));
    layer3_outputs(51) <= (layer2_outputs(849)) or (layer2_outputs(807));
    layer3_outputs(52) <= layer2_outputs(514);
    layer3_outputs(53) <= not(layer2_outputs(557)) or (layer2_outputs(370));
    layer3_outputs(54) <= layer2_outputs(65);
    layer3_outputs(55) <= (layer2_outputs(1908)) and (layer2_outputs(1150));
    layer3_outputs(56) <= not(layer2_outputs(1272));
    layer3_outputs(57) <= (layer2_outputs(1693)) and not (layer2_outputs(2345));
    layer3_outputs(58) <= '1';
    layer3_outputs(59) <= not(layer2_outputs(1710)) or (layer2_outputs(1810));
    layer3_outputs(60) <= (layer2_outputs(791)) and (layer2_outputs(874));
    layer3_outputs(61) <= layer2_outputs(1457);
    layer3_outputs(62) <= (layer2_outputs(1733)) and (layer2_outputs(998));
    layer3_outputs(63) <= (layer2_outputs(1550)) and (layer2_outputs(1208));
    layer3_outputs(64) <= '0';
    layer3_outputs(65) <= '1';
    layer3_outputs(66) <= not(layer2_outputs(128)) or (layer2_outputs(870));
    layer3_outputs(67) <= layer2_outputs(2164);
    layer3_outputs(68) <= layer2_outputs(13);
    layer3_outputs(69) <= not((layer2_outputs(1203)) or (layer2_outputs(1097)));
    layer3_outputs(70) <= layer2_outputs(2358);
    layer3_outputs(71) <= '1';
    layer3_outputs(72) <= not(layer2_outputs(1625)) or (layer2_outputs(92));
    layer3_outputs(73) <= not(layer2_outputs(725)) or (layer2_outputs(510));
    layer3_outputs(74) <= not((layer2_outputs(1085)) or (layer2_outputs(2067)));
    layer3_outputs(75) <= not(layer2_outputs(1737)) or (layer2_outputs(2368));
    layer3_outputs(76) <= (layer2_outputs(2407)) and (layer2_outputs(2217));
    layer3_outputs(77) <= layer2_outputs(946);
    layer3_outputs(78) <= not((layer2_outputs(2165)) and (layer2_outputs(1393)));
    layer3_outputs(79) <= not(layer2_outputs(2181)) or (layer2_outputs(2119));
    layer3_outputs(80) <= (layer2_outputs(2375)) and not (layer2_outputs(676));
    layer3_outputs(81) <= layer2_outputs(1530);
    layer3_outputs(82) <= (layer2_outputs(1964)) and (layer2_outputs(1746));
    layer3_outputs(83) <= not((layer2_outputs(1576)) or (layer2_outputs(772)));
    layer3_outputs(84) <= '0';
    layer3_outputs(85) <= (layer2_outputs(1646)) and not (layer2_outputs(1822));
    layer3_outputs(86) <= '1';
    layer3_outputs(87) <= layer2_outputs(25);
    layer3_outputs(88) <= layer2_outputs(1447);
    layer3_outputs(89) <= not((layer2_outputs(273)) and (layer2_outputs(924)));
    layer3_outputs(90) <= not(layer2_outputs(260));
    layer3_outputs(91) <= layer2_outputs(1065);
    layer3_outputs(92) <= not(layer2_outputs(2167));
    layer3_outputs(93) <= (layer2_outputs(269)) and not (layer2_outputs(908));
    layer3_outputs(94) <= not((layer2_outputs(1221)) and (layer2_outputs(1894)));
    layer3_outputs(95) <= not(layer2_outputs(2141));
    layer3_outputs(96) <= (layer2_outputs(616)) and not (layer2_outputs(730));
    layer3_outputs(97) <= (layer2_outputs(944)) and not (layer2_outputs(1491));
    layer3_outputs(98) <= not(layer2_outputs(1689));
    layer3_outputs(99) <= not(layer2_outputs(2460)) or (layer2_outputs(1766));
    layer3_outputs(100) <= '1';
    layer3_outputs(101) <= not(layer2_outputs(2028)) or (layer2_outputs(2500));
    layer3_outputs(102) <= not(layer2_outputs(283));
    layer3_outputs(103) <= not(layer2_outputs(295)) or (layer2_outputs(2508));
    layer3_outputs(104) <= not(layer2_outputs(86));
    layer3_outputs(105) <= (layer2_outputs(234)) and not (layer2_outputs(1068));
    layer3_outputs(106) <= not(layer2_outputs(319)) or (layer2_outputs(880));
    layer3_outputs(107) <= '0';
    layer3_outputs(108) <= (layer2_outputs(2535)) and (layer2_outputs(2440));
    layer3_outputs(109) <= not(layer2_outputs(740)) or (layer2_outputs(1098));
    layer3_outputs(110) <= not((layer2_outputs(1111)) or (layer2_outputs(1319)));
    layer3_outputs(111) <= (layer2_outputs(1496)) and not (layer2_outputs(231));
    layer3_outputs(112) <= not(layer2_outputs(352));
    layer3_outputs(113) <= (layer2_outputs(281)) or (layer2_outputs(927));
    layer3_outputs(114) <= (layer2_outputs(423)) and (layer2_outputs(916));
    layer3_outputs(115) <= not((layer2_outputs(229)) or (layer2_outputs(2540)));
    layer3_outputs(116) <= layer2_outputs(880);
    layer3_outputs(117) <= (layer2_outputs(2126)) and not (layer2_outputs(2111));
    layer3_outputs(118) <= not((layer2_outputs(1331)) or (layer2_outputs(582)));
    layer3_outputs(119) <= (layer2_outputs(1044)) or (layer2_outputs(1990));
    layer3_outputs(120) <= not(layer2_outputs(671)) or (layer2_outputs(454));
    layer3_outputs(121) <= '0';
    layer3_outputs(122) <= layer2_outputs(2191);
    layer3_outputs(123) <= not(layer2_outputs(489));
    layer3_outputs(124) <= not(layer2_outputs(1018));
    layer3_outputs(125) <= not(layer2_outputs(189));
    layer3_outputs(126) <= not(layer2_outputs(2478));
    layer3_outputs(127) <= (layer2_outputs(724)) and not (layer2_outputs(1703));
    layer3_outputs(128) <= '1';
    layer3_outputs(129) <= not(layer2_outputs(578)) or (layer2_outputs(1155));
    layer3_outputs(130) <= '0';
    layer3_outputs(131) <= not(layer2_outputs(2356));
    layer3_outputs(132) <= (layer2_outputs(1493)) or (layer2_outputs(118));
    layer3_outputs(133) <= not((layer2_outputs(2411)) or (layer2_outputs(130)));
    layer3_outputs(134) <= (layer2_outputs(1418)) and not (layer2_outputs(267));
    layer3_outputs(135) <= layer2_outputs(253);
    layer3_outputs(136) <= '0';
    layer3_outputs(137) <= layer2_outputs(819);
    layer3_outputs(138) <= not((layer2_outputs(228)) and (layer2_outputs(113)));
    layer3_outputs(139) <= (layer2_outputs(1835)) and not (layer2_outputs(433));
    layer3_outputs(140) <= layer2_outputs(837);
    layer3_outputs(141) <= (layer2_outputs(775)) and (layer2_outputs(23));
    layer3_outputs(142) <= '1';
    layer3_outputs(143) <= (layer2_outputs(1274)) and not (layer2_outputs(1088));
    layer3_outputs(144) <= not(layer2_outputs(2163)) or (layer2_outputs(922));
    layer3_outputs(145) <= (layer2_outputs(2465)) or (layer2_outputs(663));
    layer3_outputs(146) <= layer2_outputs(1175);
    layer3_outputs(147) <= '0';
    layer3_outputs(148) <= (layer2_outputs(1327)) and not (layer2_outputs(2147));
    layer3_outputs(149) <= not(layer2_outputs(1038));
    layer3_outputs(150) <= layer2_outputs(1505);
    layer3_outputs(151) <= not(layer2_outputs(2353));
    layer3_outputs(152) <= not((layer2_outputs(2190)) or (layer2_outputs(588)));
    layer3_outputs(153) <= not((layer2_outputs(710)) or (layer2_outputs(2384)));
    layer3_outputs(154) <= layer2_outputs(1161);
    layer3_outputs(155) <= (layer2_outputs(828)) xor (layer2_outputs(2430));
    layer3_outputs(156) <= '1';
    layer3_outputs(157) <= (layer2_outputs(310)) and not (layer2_outputs(1966));
    layer3_outputs(158) <= (layer2_outputs(2062)) and (layer2_outputs(1371));
    layer3_outputs(159) <= not(layer2_outputs(2272));
    layer3_outputs(160) <= not(layer2_outputs(865));
    layer3_outputs(161) <= '0';
    layer3_outputs(162) <= (layer2_outputs(901)) and not (layer2_outputs(1521));
    layer3_outputs(163) <= not(layer2_outputs(2402)) or (layer2_outputs(149));
    layer3_outputs(164) <= not(layer2_outputs(481));
    layer3_outputs(165) <= (layer2_outputs(1942)) and (layer2_outputs(1602));
    layer3_outputs(166) <= not((layer2_outputs(1430)) or (layer2_outputs(995)));
    layer3_outputs(167) <= (layer2_outputs(2221)) or (layer2_outputs(1827));
    layer3_outputs(168) <= not((layer2_outputs(1563)) or (layer2_outputs(1749)));
    layer3_outputs(169) <= (layer2_outputs(2245)) and (layer2_outputs(808));
    layer3_outputs(170) <= layer2_outputs(1860);
    layer3_outputs(171) <= not((layer2_outputs(2251)) xor (layer2_outputs(1009)));
    layer3_outputs(172) <= not(layer2_outputs(2553)) or (layer2_outputs(1608));
    layer3_outputs(173) <= '0';
    layer3_outputs(174) <= not((layer2_outputs(837)) or (layer2_outputs(31)));
    layer3_outputs(175) <= not(layer2_outputs(2399)) or (layer2_outputs(1674));
    layer3_outputs(176) <= not(layer2_outputs(867)) or (layer2_outputs(815));
    layer3_outputs(177) <= (layer2_outputs(183)) or (layer2_outputs(464));
    layer3_outputs(178) <= '0';
    layer3_outputs(179) <= not(layer2_outputs(1214));
    layer3_outputs(180) <= not(layer2_outputs(1516));
    layer3_outputs(181) <= layer2_outputs(2121);
    layer3_outputs(182) <= not(layer2_outputs(1913)) or (layer2_outputs(2081));
    layer3_outputs(183) <= not(layer2_outputs(1667)) or (layer2_outputs(194));
    layer3_outputs(184) <= (layer2_outputs(2321)) and (layer2_outputs(872));
    layer3_outputs(185) <= (layer2_outputs(95)) and not (layer2_outputs(1712));
    layer3_outputs(186) <= (layer2_outputs(2459)) and not (layer2_outputs(1878));
    layer3_outputs(187) <= (layer2_outputs(667)) or (layer2_outputs(1997));
    layer3_outputs(188) <= not(layer2_outputs(158));
    layer3_outputs(189) <= (layer2_outputs(166)) and not (layer2_outputs(1023));
    layer3_outputs(190) <= '1';
    layer3_outputs(191) <= not(layer2_outputs(1221));
    layer3_outputs(192) <= not(layer2_outputs(731)) or (layer2_outputs(1410));
    layer3_outputs(193) <= (layer2_outputs(1941)) or (layer2_outputs(1318));
    layer3_outputs(194) <= layer2_outputs(582);
    layer3_outputs(195) <= not(layer2_outputs(1717));
    layer3_outputs(196) <= layer2_outputs(972);
    layer3_outputs(197) <= not(layer2_outputs(28)) or (layer2_outputs(1656));
    layer3_outputs(198) <= layer2_outputs(470);
    layer3_outputs(199) <= layer2_outputs(730);
    layer3_outputs(200) <= not(layer2_outputs(1943)) or (layer2_outputs(1598));
    layer3_outputs(201) <= (layer2_outputs(877)) and (layer2_outputs(1644));
    layer3_outputs(202) <= (layer2_outputs(404)) and not (layer2_outputs(891));
    layer3_outputs(203) <= not(layer2_outputs(1823));
    layer3_outputs(204) <= not(layer2_outputs(1520)) or (layer2_outputs(186));
    layer3_outputs(205) <= '0';
    layer3_outputs(206) <= (layer2_outputs(2469)) or (layer2_outputs(2387));
    layer3_outputs(207) <= (layer2_outputs(1804)) and (layer2_outputs(274));
    layer3_outputs(208) <= not(layer2_outputs(1763)) or (layer2_outputs(1338));
    layer3_outputs(209) <= not(layer2_outputs(2246)) or (layer2_outputs(1692));
    layer3_outputs(210) <= (layer2_outputs(607)) xor (layer2_outputs(1788));
    layer3_outputs(211) <= (layer2_outputs(1818)) and not (layer2_outputs(869));
    layer3_outputs(212) <= not(layer2_outputs(336)) or (layer2_outputs(1024));
    layer3_outputs(213) <= layer2_outputs(881);
    layer3_outputs(214) <= layer2_outputs(380);
    layer3_outputs(215) <= not(layer2_outputs(1424)) or (layer2_outputs(1091));
    layer3_outputs(216) <= layer2_outputs(273);
    layer3_outputs(217) <= (layer2_outputs(2343)) and (layer2_outputs(2406));
    layer3_outputs(218) <= not(layer2_outputs(938));
    layer3_outputs(219) <= layer2_outputs(1134);
    layer3_outputs(220) <= not(layer2_outputs(321));
    layer3_outputs(221) <= not(layer2_outputs(1530)) or (layer2_outputs(1779));
    layer3_outputs(222) <= not(layer2_outputs(148)) or (layer2_outputs(1905));
    layer3_outputs(223) <= (layer2_outputs(1469)) and (layer2_outputs(1176));
    layer3_outputs(224) <= not(layer2_outputs(1727));
    layer3_outputs(225) <= layer2_outputs(1370);
    layer3_outputs(226) <= '1';
    layer3_outputs(227) <= (layer2_outputs(1403)) or (layer2_outputs(2447));
    layer3_outputs(228) <= not((layer2_outputs(851)) or (layer2_outputs(1653)));
    layer3_outputs(229) <= (layer2_outputs(1316)) and not (layer2_outputs(1208));
    layer3_outputs(230) <= not(layer2_outputs(1145));
    layer3_outputs(231) <= '0';
    layer3_outputs(232) <= (layer2_outputs(2408)) and not (layer2_outputs(733));
    layer3_outputs(233) <= layer2_outputs(619);
    layer3_outputs(234) <= '0';
    layer3_outputs(235) <= not(layer2_outputs(1425));
    layer3_outputs(236) <= not(layer2_outputs(1946));
    layer3_outputs(237) <= (layer2_outputs(1954)) and not (layer2_outputs(227));
    layer3_outputs(238) <= layer2_outputs(125);
    layer3_outputs(239) <= not(layer2_outputs(1239));
    layer3_outputs(240) <= (layer2_outputs(1457)) and not (layer2_outputs(1537));
    layer3_outputs(241) <= layer2_outputs(2153);
    layer3_outputs(242) <= not((layer2_outputs(664)) or (layer2_outputs(432)));
    layer3_outputs(243) <= (layer2_outputs(1237)) or (layer2_outputs(2334));
    layer3_outputs(244) <= layer2_outputs(2258);
    layer3_outputs(245) <= (layer2_outputs(308)) and (layer2_outputs(652));
    layer3_outputs(246) <= not(layer2_outputs(1162));
    layer3_outputs(247) <= (layer2_outputs(2167)) or (layer2_outputs(625));
    layer3_outputs(248) <= not(layer2_outputs(24)) or (layer2_outputs(1187));
    layer3_outputs(249) <= (layer2_outputs(2483)) and not (layer2_outputs(2300));
    layer3_outputs(250) <= not(layer2_outputs(50)) or (layer2_outputs(794));
    layer3_outputs(251) <= not((layer2_outputs(522)) or (layer2_outputs(2246)));
    layer3_outputs(252) <= '1';
    layer3_outputs(253) <= not((layer2_outputs(1593)) or (layer2_outputs(1608)));
    layer3_outputs(254) <= '1';
    layer3_outputs(255) <= not(layer2_outputs(2404)) or (layer2_outputs(607));
    layer3_outputs(256) <= not(layer2_outputs(2466));
    layer3_outputs(257) <= not(layer2_outputs(285));
    layer3_outputs(258) <= layer2_outputs(1013);
    layer3_outputs(259) <= layer2_outputs(1025);
    layer3_outputs(260) <= '1';
    layer3_outputs(261) <= (layer2_outputs(555)) and not (layer2_outputs(1061));
    layer3_outputs(262) <= '1';
    layer3_outputs(263) <= (layer2_outputs(1643)) and not (layer2_outputs(1138));
    layer3_outputs(264) <= not(layer2_outputs(399));
    layer3_outputs(265) <= layer2_outputs(2556);
    layer3_outputs(266) <= not(layer2_outputs(1348));
    layer3_outputs(267) <= not(layer2_outputs(459));
    layer3_outputs(268) <= '0';
    layer3_outputs(269) <= (layer2_outputs(282)) and not (layer2_outputs(1497));
    layer3_outputs(270) <= (layer2_outputs(1663)) or (layer2_outputs(77));
    layer3_outputs(271) <= not(layer2_outputs(898));
    layer3_outputs(272) <= (layer2_outputs(1895)) or (layer2_outputs(1201));
    layer3_outputs(273) <= not(layer2_outputs(1083));
    layer3_outputs(274) <= layer2_outputs(323);
    layer3_outputs(275) <= (layer2_outputs(1)) and (layer2_outputs(464));
    layer3_outputs(276) <= not(layer2_outputs(2363));
    layer3_outputs(277) <= layer2_outputs(1024);
    layer3_outputs(278) <= '0';
    layer3_outputs(279) <= not(layer2_outputs(238)) or (layer2_outputs(1619));
    layer3_outputs(280) <= (layer2_outputs(1476)) and not (layer2_outputs(2026));
    layer3_outputs(281) <= not(layer2_outputs(589)) or (layer2_outputs(2176));
    layer3_outputs(282) <= (layer2_outputs(1798)) and (layer2_outputs(2014));
    layer3_outputs(283) <= (layer2_outputs(1524)) and not (layer2_outputs(1197));
    layer3_outputs(284) <= layer2_outputs(1468);
    layer3_outputs(285) <= not(layer2_outputs(508));
    layer3_outputs(286) <= (layer2_outputs(1890)) and (layer2_outputs(699));
    layer3_outputs(287) <= not((layer2_outputs(112)) or (layer2_outputs(137)));
    layer3_outputs(288) <= layer2_outputs(33);
    layer3_outputs(289) <= layer2_outputs(1255);
    layer3_outputs(290) <= not(layer2_outputs(448)) or (layer2_outputs(611));
    layer3_outputs(291) <= not(layer2_outputs(1385));
    layer3_outputs(292) <= not(layer2_outputs(1706));
    layer3_outputs(293) <= not(layer2_outputs(1605));
    layer3_outputs(294) <= '1';
    layer3_outputs(295) <= not(layer2_outputs(329)) or (layer2_outputs(820));
    layer3_outputs(296) <= not(layer2_outputs(1611)) or (layer2_outputs(53));
    layer3_outputs(297) <= '1';
    layer3_outputs(298) <= (layer2_outputs(1684)) or (layer2_outputs(2123));
    layer3_outputs(299) <= '0';
    layer3_outputs(300) <= (layer2_outputs(1129)) and not (layer2_outputs(719));
    layer3_outputs(301) <= '0';
    layer3_outputs(302) <= '0';
    layer3_outputs(303) <= layer2_outputs(1673);
    layer3_outputs(304) <= not((layer2_outputs(584)) and (layer2_outputs(954)));
    layer3_outputs(305) <= not((layer2_outputs(1755)) or (layer2_outputs(1512)));
    layer3_outputs(306) <= not(layer2_outputs(1402));
    layer3_outputs(307) <= layer2_outputs(1124);
    layer3_outputs(308) <= (layer2_outputs(1785)) and not (layer2_outputs(326));
    layer3_outputs(309) <= layer2_outputs(912);
    layer3_outputs(310) <= not(layer2_outputs(1059));
    layer3_outputs(311) <= layer2_outputs(551);
    layer3_outputs(312) <= (layer2_outputs(88)) and not (layer2_outputs(154));
    layer3_outputs(313) <= layer2_outputs(2476);
    layer3_outputs(314) <= (layer2_outputs(1312)) and not (layer2_outputs(377));
    layer3_outputs(315) <= (layer2_outputs(904)) and (layer2_outputs(1074));
    layer3_outputs(316) <= layer2_outputs(1973);
    layer3_outputs(317) <= (layer2_outputs(777)) and (layer2_outputs(871));
    layer3_outputs(318) <= not(layer2_outputs(1276));
    layer3_outputs(319) <= not(layer2_outputs(2269)) or (layer2_outputs(1083));
    layer3_outputs(320) <= not((layer2_outputs(1272)) or (layer2_outputs(1418)));
    layer3_outputs(321) <= not((layer2_outputs(1006)) and (layer2_outputs(2197)));
    layer3_outputs(322) <= layer2_outputs(2280);
    layer3_outputs(323) <= not(layer2_outputs(1876));
    layer3_outputs(324) <= not(layer2_outputs(1554));
    layer3_outputs(325) <= not(layer2_outputs(1969));
    layer3_outputs(326) <= not(layer2_outputs(695));
    layer3_outputs(327) <= layer2_outputs(2261);
    layer3_outputs(328) <= (layer2_outputs(67)) and not (layer2_outputs(962));
    layer3_outputs(329) <= not((layer2_outputs(2414)) or (layer2_outputs(271)));
    layer3_outputs(330) <= not((layer2_outputs(1797)) xor (layer2_outputs(2352)));
    layer3_outputs(331) <= (layer2_outputs(2536)) and not (layer2_outputs(125));
    layer3_outputs(332) <= not((layer2_outputs(324)) xor (layer2_outputs(1565)));
    layer3_outputs(333) <= not(layer2_outputs(1084)) or (layer2_outputs(809));
    layer3_outputs(334) <= not(layer2_outputs(1706));
    layer3_outputs(335) <= '0';
    layer3_outputs(336) <= layer2_outputs(1518);
    layer3_outputs(337) <= layer2_outputs(1621);
    layer3_outputs(338) <= (layer2_outputs(2148)) and not (layer2_outputs(435));
    layer3_outputs(339) <= (layer2_outputs(1895)) or (layer2_outputs(1916));
    layer3_outputs(340) <= layer2_outputs(446);
    layer3_outputs(341) <= not((layer2_outputs(2328)) or (layer2_outputs(1660)));
    layer3_outputs(342) <= not(layer2_outputs(974));
    layer3_outputs(343) <= not(layer2_outputs(2104));
    layer3_outputs(344) <= not((layer2_outputs(2039)) or (layer2_outputs(2517)));
    layer3_outputs(345) <= not((layer2_outputs(2021)) and (layer2_outputs(1149)));
    layer3_outputs(346) <= layer2_outputs(2225);
    layer3_outputs(347) <= layer2_outputs(2271);
    layer3_outputs(348) <= (layer2_outputs(327)) and not (layer2_outputs(1004));
    layer3_outputs(349) <= not((layer2_outputs(1487)) or (layer2_outputs(144)));
    layer3_outputs(350) <= (layer2_outputs(2155)) and not (layer2_outputs(350));
    layer3_outputs(351) <= (layer2_outputs(1008)) and not (layer2_outputs(1389));
    layer3_outputs(352) <= (layer2_outputs(895)) and (layer2_outputs(1902));
    layer3_outputs(353) <= layer2_outputs(1172);
    layer3_outputs(354) <= not((layer2_outputs(2534)) and (layer2_outputs(400)));
    layer3_outputs(355) <= not(layer2_outputs(2396));
    layer3_outputs(356) <= '0';
    layer3_outputs(357) <= not(layer2_outputs(769));
    layer3_outputs(358) <= (layer2_outputs(2126)) or (layer2_outputs(2501));
    layer3_outputs(359) <= layer2_outputs(2493);
    layer3_outputs(360) <= '1';
    layer3_outputs(361) <= (layer2_outputs(460)) and not (layer2_outputs(2005));
    layer3_outputs(362) <= '0';
    layer3_outputs(363) <= layer2_outputs(1266);
    layer3_outputs(364) <= not(layer2_outputs(1001)) or (layer2_outputs(1831));
    layer3_outputs(365) <= not((layer2_outputs(1409)) or (layer2_outputs(741)));
    layer3_outputs(366) <= not(layer2_outputs(419)) or (layer2_outputs(1379));
    layer3_outputs(367) <= layer2_outputs(901);
    layer3_outputs(368) <= not((layer2_outputs(2176)) and (layer2_outputs(2037)));
    layer3_outputs(369) <= not((layer2_outputs(1691)) and (layer2_outputs(1790)));
    layer3_outputs(370) <= '0';
    layer3_outputs(371) <= layer2_outputs(110);
    layer3_outputs(372) <= '0';
    layer3_outputs(373) <= layer2_outputs(1435);
    layer3_outputs(374) <= not((layer2_outputs(1564)) or (layer2_outputs(636)));
    layer3_outputs(375) <= layer2_outputs(1986);
    layer3_outputs(376) <= (layer2_outputs(368)) and not (layer2_outputs(244));
    layer3_outputs(377) <= (layer2_outputs(1293)) or (layer2_outputs(123));
    layer3_outputs(378) <= (layer2_outputs(2475)) or (layer2_outputs(2438));
    layer3_outputs(379) <= not(layer2_outputs(968));
    layer3_outputs(380) <= layer2_outputs(1787);
    layer3_outputs(381) <= not(layer2_outputs(1639));
    layer3_outputs(382) <= not((layer2_outputs(1238)) and (layer2_outputs(1505)));
    layer3_outputs(383) <= '0';
    layer3_outputs(384) <= (layer2_outputs(178)) and not (layer2_outputs(619));
    layer3_outputs(385) <= layer2_outputs(2235);
    layer3_outputs(386) <= layer2_outputs(1067);
    layer3_outputs(387) <= layer2_outputs(777);
    layer3_outputs(388) <= not(layer2_outputs(1233));
    layer3_outputs(389) <= (layer2_outputs(132)) and not (layer2_outputs(2474));
    layer3_outputs(390) <= (layer2_outputs(90)) and not (layer2_outputs(2137));
    layer3_outputs(391) <= not((layer2_outputs(1925)) and (layer2_outputs(883)));
    layer3_outputs(392) <= not((layer2_outputs(1724)) and (layer2_outputs(1598)));
    layer3_outputs(393) <= not(layer2_outputs(2158));
    layer3_outputs(394) <= (layer2_outputs(925)) and not (layer2_outputs(756));
    layer3_outputs(395) <= (layer2_outputs(249)) and not (layer2_outputs(970));
    layer3_outputs(396) <= not(layer2_outputs(1940));
    layer3_outputs(397) <= layer2_outputs(394);
    layer3_outputs(398) <= (layer2_outputs(2152)) or (layer2_outputs(1303));
    layer3_outputs(399) <= (layer2_outputs(1037)) xor (layer2_outputs(149));
    layer3_outputs(400) <= layer2_outputs(1692);
    layer3_outputs(401) <= '0';
    layer3_outputs(402) <= (layer2_outputs(1157)) and not (layer2_outputs(1347));
    layer3_outputs(403) <= not((layer2_outputs(1387)) or (layer2_outputs(1825)));
    layer3_outputs(404) <= not(layer2_outputs(2160)) or (layer2_outputs(2401));
    layer3_outputs(405) <= not(layer2_outputs(1187));
    layer3_outputs(406) <= not((layer2_outputs(215)) or (layer2_outputs(1632)));
    layer3_outputs(407) <= not(layer2_outputs(404));
    layer3_outputs(408) <= not((layer2_outputs(2420)) or (layer2_outputs(1918)));
    layer3_outputs(409) <= not(layer2_outputs(2043));
    layer3_outputs(410) <= (layer2_outputs(1881)) and (layer2_outputs(1740));
    layer3_outputs(411) <= (layer2_outputs(696)) and (layer2_outputs(1169));
    layer3_outputs(412) <= not((layer2_outputs(844)) or (layer2_outputs(2296)));
    layer3_outputs(413) <= not(layer2_outputs(2538)) or (layer2_outputs(583));
    layer3_outputs(414) <= layer2_outputs(591);
    layer3_outputs(415) <= not(layer2_outputs(426)) or (layer2_outputs(2146));
    layer3_outputs(416) <= not((layer2_outputs(2360)) or (layer2_outputs(2064)));
    layer3_outputs(417) <= (layer2_outputs(2047)) and (layer2_outputs(2166));
    layer3_outputs(418) <= (layer2_outputs(2059)) or (layer2_outputs(1837));
    layer3_outputs(419) <= (layer2_outputs(493)) and (layer2_outputs(266));
    layer3_outputs(420) <= not(layer2_outputs(1668)) or (layer2_outputs(1884));
    layer3_outputs(421) <= not(layer2_outputs(1310));
    layer3_outputs(422) <= (layer2_outputs(401)) and not (layer2_outputs(215));
    layer3_outputs(423) <= (layer2_outputs(1057)) and (layer2_outputs(2225));
    layer3_outputs(424) <= '0';
    layer3_outputs(425) <= not(layer2_outputs(1599));
    layer3_outputs(426) <= (layer2_outputs(692)) and not (layer2_outputs(36));
    layer3_outputs(427) <= layer2_outputs(444);
    layer3_outputs(428) <= not(layer2_outputs(677));
    layer3_outputs(429) <= '0';
    layer3_outputs(430) <= (layer2_outputs(1555)) and not (layer2_outputs(1900));
    layer3_outputs(431) <= (layer2_outputs(1181)) and not (layer2_outputs(838));
    layer3_outputs(432) <= layer2_outputs(465);
    layer3_outputs(433) <= '1';
    layer3_outputs(434) <= (layer2_outputs(1649)) and not (layer2_outputs(2280));
    layer3_outputs(435) <= not(layer2_outputs(119));
    layer3_outputs(436) <= not(layer2_outputs(259));
    layer3_outputs(437) <= not((layer2_outputs(799)) or (layer2_outputs(470)));
    layer3_outputs(438) <= (layer2_outputs(1)) and (layer2_outputs(259));
    layer3_outputs(439) <= (layer2_outputs(1743)) and not (layer2_outputs(2210));
    layer3_outputs(440) <= (layer2_outputs(601)) and not (layer2_outputs(1871));
    layer3_outputs(441) <= not(layer2_outputs(1539));
    layer3_outputs(442) <= not(layer2_outputs(825));
    layer3_outputs(443) <= '1';
    layer3_outputs(444) <= not(layer2_outputs(1901));
    layer3_outputs(445) <= (layer2_outputs(2014)) and not (layer2_outputs(715));
    layer3_outputs(446) <= (layer2_outputs(2189)) and (layer2_outputs(2546));
    layer3_outputs(447) <= not((layer2_outputs(2376)) xor (layer2_outputs(2123)));
    layer3_outputs(448) <= not(layer2_outputs(2143));
    layer3_outputs(449) <= '0';
    layer3_outputs(450) <= (layer2_outputs(1868)) and not (layer2_outputs(1390));
    layer3_outputs(451) <= not((layer2_outputs(1449)) or (layer2_outputs(1410)));
    layer3_outputs(452) <= not(layer2_outputs(6));
    layer3_outputs(453) <= layer2_outputs(694);
    layer3_outputs(454) <= (layer2_outputs(35)) or (layer2_outputs(1590));
    layer3_outputs(455) <= not(layer2_outputs(757)) or (layer2_outputs(599));
    layer3_outputs(456) <= not(layer2_outputs(168));
    layer3_outputs(457) <= not((layer2_outputs(375)) or (layer2_outputs(560)));
    layer3_outputs(458) <= layer2_outputs(2053);
    layer3_outputs(459) <= not(layer2_outputs(1206)) or (layer2_outputs(1196));
    layer3_outputs(460) <= layer2_outputs(1983);
    layer3_outputs(461) <= not((layer2_outputs(314)) xor (layer2_outputs(1298)));
    layer3_outputs(462) <= not(layer2_outputs(1219));
    layer3_outputs(463) <= layer2_outputs(278);
    layer3_outputs(464) <= not((layer2_outputs(1709)) and (layer2_outputs(2358)));
    layer3_outputs(465) <= '1';
    layer3_outputs(466) <= (layer2_outputs(232)) and not (layer2_outputs(65));
    layer3_outputs(467) <= layer2_outputs(2348);
    layer3_outputs(468) <= (layer2_outputs(1639)) and (layer2_outputs(1347));
    layer3_outputs(469) <= not((layer2_outputs(1651)) and (layer2_outputs(1954)));
    layer3_outputs(470) <= not(layer2_outputs(941));
    layer3_outputs(471) <= (layer2_outputs(575)) and (layer2_outputs(1264));
    layer3_outputs(472) <= (layer2_outputs(119)) and not (layer2_outputs(1864));
    layer3_outputs(473) <= not((layer2_outputs(254)) or (layer2_outputs(553)));
    layer3_outputs(474) <= not(layer2_outputs(2267)) or (layer2_outputs(967));
    layer3_outputs(475) <= not(layer2_outputs(691)) or (layer2_outputs(2218));
    layer3_outputs(476) <= not((layer2_outputs(2050)) and (layer2_outputs(786)));
    layer3_outputs(477) <= layer2_outputs(2543);
    layer3_outputs(478) <= not(layer2_outputs(760));
    layer3_outputs(479) <= layer2_outputs(1115);
    layer3_outputs(480) <= '1';
    layer3_outputs(481) <= not(layer2_outputs(466)) or (layer2_outputs(542));
    layer3_outputs(482) <= layer2_outputs(2299);
    layer3_outputs(483) <= not(layer2_outputs(920));
    layer3_outputs(484) <= not((layer2_outputs(1057)) and (layer2_outputs(1252)));
    layer3_outputs(485) <= layer2_outputs(1760);
    layer3_outputs(486) <= layer2_outputs(1078);
    layer3_outputs(487) <= layer2_outputs(1588);
    layer3_outputs(488) <= not(layer2_outputs(903));
    layer3_outputs(489) <= layer2_outputs(534);
    layer3_outputs(490) <= not(layer2_outputs(1767)) or (layer2_outputs(142));
    layer3_outputs(491) <= layer2_outputs(2089);
    layer3_outputs(492) <= not((layer2_outputs(1526)) and (layer2_outputs(1451)));
    layer3_outputs(493) <= layer2_outputs(2022);
    layer3_outputs(494) <= not(layer2_outputs(591));
    layer3_outputs(495) <= not(layer2_outputs(159)) or (layer2_outputs(2150));
    layer3_outputs(496) <= (layer2_outputs(2373)) and not (layer2_outputs(2211));
    layer3_outputs(497) <= layer2_outputs(664);
    layer3_outputs(498) <= '1';
    layer3_outputs(499) <= (layer2_outputs(2482)) and not (layer2_outputs(798));
    layer3_outputs(500) <= not((layer2_outputs(1760)) or (layer2_outputs(1059)));
    layer3_outputs(501) <= (layer2_outputs(396)) and not (layer2_outputs(2118));
    layer3_outputs(502) <= not(layer2_outputs(1232));
    layer3_outputs(503) <= layer2_outputs(2371);
    layer3_outputs(504) <= (layer2_outputs(1077)) and (layer2_outputs(260));
    layer3_outputs(505) <= not(layer2_outputs(1149)) or (layer2_outputs(1356));
    layer3_outputs(506) <= not((layer2_outputs(374)) or (layer2_outputs(188)));
    layer3_outputs(507) <= '0';
    layer3_outputs(508) <= layer2_outputs(1788);
    layer3_outputs(509) <= (layer2_outputs(1850)) or (layer2_outputs(1631));
    layer3_outputs(510) <= not((layer2_outputs(1148)) and (layer2_outputs(202)));
    layer3_outputs(511) <= layer2_outputs(447);
    layer3_outputs(512) <= (layer2_outputs(2254)) and (layer2_outputs(2078));
    layer3_outputs(513) <= (layer2_outputs(2352)) and not (layer2_outputs(614));
    layer3_outputs(514) <= '0';
    layer3_outputs(515) <= layer2_outputs(2519);
    layer3_outputs(516) <= layer2_outputs(433);
    layer3_outputs(517) <= layer2_outputs(624);
    layer3_outputs(518) <= '1';
    layer3_outputs(519) <= not(layer2_outputs(1792));
    layer3_outputs(520) <= (layer2_outputs(1486)) and not (layer2_outputs(2329));
    layer3_outputs(521) <= layer2_outputs(80);
    layer3_outputs(522) <= not((layer2_outputs(978)) and (layer2_outputs(1906)));
    layer3_outputs(523) <= not(layer2_outputs(1732)) or (layer2_outputs(367));
    layer3_outputs(524) <= (layer2_outputs(1127)) or (layer2_outputs(1158));
    layer3_outputs(525) <= layer2_outputs(1096);
    layer3_outputs(526) <= '0';
    layer3_outputs(527) <= not((layer2_outputs(1173)) or (layer2_outputs(2226)));
    layer3_outputs(528) <= (layer2_outputs(677)) and (layer2_outputs(765));
    layer3_outputs(529) <= (layer2_outputs(649)) xor (layer2_outputs(1741));
    layer3_outputs(530) <= not(layer2_outputs(136)) or (layer2_outputs(2023));
    layer3_outputs(531) <= layer2_outputs(806);
    layer3_outputs(532) <= '0';
    layer3_outputs(533) <= (layer2_outputs(1624)) and (layer2_outputs(1602));
    layer3_outputs(534) <= not(layer2_outputs(1802)) or (layer2_outputs(1440));
    layer3_outputs(535) <= (layer2_outputs(385)) and not (layer2_outputs(1380));
    layer3_outputs(536) <= layer2_outputs(520);
    layer3_outputs(537) <= '1';
    layer3_outputs(538) <= '0';
    layer3_outputs(539) <= (layer2_outputs(2194)) or (layer2_outputs(1714));
    layer3_outputs(540) <= (layer2_outputs(2439)) or (layer2_outputs(931));
    layer3_outputs(541) <= layer2_outputs(751);
    layer3_outputs(542) <= layer2_outputs(569);
    layer3_outputs(543) <= (layer2_outputs(1043)) and (layer2_outputs(1943));
    layer3_outputs(544) <= not(layer2_outputs(913)) or (layer2_outputs(597));
    layer3_outputs(545) <= (layer2_outputs(1855)) and not (layer2_outputs(346));
    layer3_outputs(546) <= '1';
    layer3_outputs(547) <= not((layer2_outputs(441)) or (layer2_outputs(1968)));
    layer3_outputs(548) <= layer2_outputs(364);
    layer3_outputs(549) <= '1';
    layer3_outputs(550) <= not(layer2_outputs(1659));
    layer3_outputs(551) <= not(layer2_outputs(1786));
    layer3_outputs(552) <= (layer2_outputs(1371)) and not (layer2_outputs(1630));
    layer3_outputs(553) <= not(layer2_outputs(1068)) or (layer2_outputs(2045));
    layer3_outputs(554) <= not(layer2_outputs(1387));
    layer3_outputs(555) <= layer2_outputs(2556);
    layer3_outputs(556) <= not(layer2_outputs(647));
    layer3_outputs(557) <= (layer2_outputs(949)) and not (layer2_outputs(1555));
    layer3_outputs(558) <= layer2_outputs(2446);
    layer3_outputs(559) <= '1';
    layer3_outputs(560) <= not(layer2_outputs(640));
    layer3_outputs(561) <= not((layer2_outputs(1318)) or (layer2_outputs(2203)));
    layer3_outputs(562) <= not(layer2_outputs(1118)) or (layer2_outputs(1256));
    layer3_outputs(563) <= '0';
    layer3_outputs(564) <= not(layer2_outputs(2308)) or (layer2_outputs(1046));
    layer3_outputs(565) <= (layer2_outputs(613)) xor (layer2_outputs(831));
    layer3_outputs(566) <= layer2_outputs(989);
    layer3_outputs(567) <= not(layer2_outputs(1026));
    layer3_outputs(568) <= not((layer2_outputs(1842)) or (layer2_outputs(1126)));
    layer3_outputs(569) <= '1';
    layer3_outputs(570) <= (layer2_outputs(1212)) and not (layer2_outputs(2457));
    layer3_outputs(571) <= (layer2_outputs(2330)) and not (layer2_outputs(1652));
    layer3_outputs(572) <= not((layer2_outputs(961)) and (layer2_outputs(2236)));
    layer3_outputs(573) <= (layer2_outputs(994)) and not (layer2_outputs(1355));
    layer3_outputs(574) <= layer2_outputs(637);
    layer3_outputs(575) <= (layer2_outputs(612)) and (layer2_outputs(369));
    layer3_outputs(576) <= not(layer2_outputs(858));
    layer3_outputs(577) <= not(layer2_outputs(986)) or (layer2_outputs(1301));
    layer3_outputs(578) <= (layer2_outputs(2179)) and not (layer2_outputs(519));
    layer3_outputs(579) <= layer2_outputs(1958);
    layer3_outputs(580) <= (layer2_outputs(1496)) and not (layer2_outputs(2147));
    layer3_outputs(581) <= (layer2_outputs(1506)) or (layer2_outputs(158));
    layer3_outputs(582) <= (layer2_outputs(54)) and not (layer2_outputs(429));
    layer3_outputs(583) <= not(layer2_outputs(27));
    layer3_outputs(584) <= not(layer2_outputs(152));
    layer3_outputs(585) <= not(layer2_outputs(1537));
    layer3_outputs(586) <= not(layer2_outputs(696));
    layer3_outputs(587) <= (layer2_outputs(1212)) and not (layer2_outputs(1155));
    layer3_outputs(588) <= (layer2_outputs(396)) and not (layer2_outputs(996));
    layer3_outputs(589) <= layer2_outputs(532);
    layer3_outputs(590) <= (layer2_outputs(1092)) or (layer2_outputs(813));
    layer3_outputs(591) <= (layer2_outputs(145)) and (layer2_outputs(821));
    layer3_outputs(592) <= not((layer2_outputs(1065)) and (layer2_outputs(1514)));
    layer3_outputs(593) <= '1';
    layer3_outputs(594) <= '1';
    layer3_outputs(595) <= (layer2_outputs(2484)) and not (layer2_outputs(1620));
    layer3_outputs(596) <= layer2_outputs(2136);
    layer3_outputs(597) <= (layer2_outputs(1742)) and (layer2_outputs(166));
    layer3_outputs(598) <= (layer2_outputs(2038)) and (layer2_outputs(2317));
    layer3_outputs(599) <= (layer2_outputs(246)) xor (layer2_outputs(398));
    layer3_outputs(600) <= not(layer2_outputs(299));
    layer3_outputs(601) <= (layer2_outputs(1789)) and (layer2_outputs(435));
    layer3_outputs(602) <= not(layer2_outputs(2048));
    layer3_outputs(603) <= not(layer2_outputs(2462));
    layer3_outputs(604) <= not(layer2_outputs(2439)) or (layer2_outputs(133));
    layer3_outputs(605) <= not(layer2_outputs(1852));
    layer3_outputs(606) <= not((layer2_outputs(2076)) xor (layer2_outputs(1053)));
    layer3_outputs(607) <= '1';
    layer3_outputs(608) <= layer2_outputs(1416);
    layer3_outputs(609) <= not(layer2_outputs(462)) or (layer2_outputs(296));
    layer3_outputs(610) <= (layer2_outputs(635)) and not (layer2_outputs(661));
    layer3_outputs(611) <= layer2_outputs(1847);
    layer3_outputs(612) <= not((layer2_outputs(2287)) and (layer2_outputs(2062)));
    layer3_outputs(613) <= not((layer2_outputs(2131)) and (layer2_outputs(2555)));
    layer3_outputs(614) <= '0';
    layer3_outputs(615) <= (layer2_outputs(556)) and not (layer2_outputs(675));
    layer3_outputs(616) <= not(layer2_outputs(1454)) or (layer2_outputs(1159));
    layer3_outputs(617) <= (layer2_outputs(2331)) or (layer2_outputs(494));
    layer3_outputs(618) <= not((layer2_outputs(546)) and (layer2_outputs(952)));
    layer3_outputs(619) <= (layer2_outputs(553)) or (layer2_outputs(838));
    layer3_outputs(620) <= (layer2_outputs(773)) and (layer2_outputs(1038));
    layer3_outputs(621) <= (layer2_outputs(617)) xor (layer2_outputs(1252));
    layer3_outputs(622) <= not(layer2_outputs(55)) or (layer2_outputs(1382));
    layer3_outputs(623) <= '1';
    layer3_outputs(624) <= (layer2_outputs(1663)) or (layer2_outputs(1758));
    layer3_outputs(625) <= (layer2_outputs(2481)) or (layer2_outputs(1412));
    layer3_outputs(626) <= '1';
    layer3_outputs(627) <= not((layer2_outputs(876)) or (layer2_outputs(811)));
    layer3_outputs(628) <= not((layer2_outputs(2428)) and (layer2_outputs(2078)));
    layer3_outputs(629) <= not((layer2_outputs(148)) and (layer2_outputs(347)));
    layer3_outputs(630) <= (layer2_outputs(1076)) or (layer2_outputs(1828));
    layer3_outputs(631) <= '1';
    layer3_outputs(632) <= layer2_outputs(1137);
    layer3_outputs(633) <= not(layer2_outputs(1747));
    layer3_outputs(634) <= (layer2_outputs(371)) and not (layer2_outputs(1573));
    layer3_outputs(635) <= (layer2_outputs(1551)) and not (layer2_outputs(153));
    layer3_outputs(636) <= not(layer2_outputs(1250)) or (layer2_outputs(1045));
    layer3_outputs(637) <= (layer2_outputs(359)) and not (layer2_outputs(1206));
    layer3_outputs(638) <= (layer2_outputs(2266)) and (layer2_outputs(1317));
    layer3_outputs(639) <= (layer2_outputs(1684)) and not (layer2_outputs(1066));
    layer3_outputs(640) <= (layer2_outputs(979)) and (layer2_outputs(1876));
    layer3_outputs(641) <= (layer2_outputs(2370)) and (layer2_outputs(1707));
    layer3_outputs(642) <= layer2_outputs(1342);
    layer3_outputs(643) <= not(layer2_outputs(495)) or (layer2_outputs(2341));
    layer3_outputs(644) <= not(layer2_outputs(1400)) or (layer2_outputs(1683));
    layer3_outputs(645) <= (layer2_outputs(2223)) and not (layer2_outputs(1462));
    layer3_outputs(646) <= '1';
    layer3_outputs(647) <= '0';
    layer3_outputs(648) <= not(layer2_outputs(469)) or (layer2_outputs(1314));
    layer3_outputs(649) <= not(layer2_outputs(1551)) or (layer2_outputs(891));
    layer3_outputs(650) <= (layer2_outputs(563)) and not (layer2_outputs(2080));
    layer3_outputs(651) <= not(layer2_outputs(978));
    layer3_outputs(652) <= not(layer2_outputs(2522));
    layer3_outputs(653) <= (layer2_outputs(2479)) or (layer2_outputs(2467));
    layer3_outputs(654) <= layer2_outputs(1234);
    layer3_outputs(655) <= (layer2_outputs(1091)) or (layer2_outputs(1029));
    layer3_outputs(656) <= (layer2_outputs(2204)) or (layer2_outputs(1023));
    layer3_outputs(657) <= (layer2_outputs(1744)) or (layer2_outputs(2331));
    layer3_outputs(658) <= not(layer2_outputs(751));
    layer3_outputs(659) <= (layer2_outputs(965)) and not (layer2_outputs(326));
    layer3_outputs(660) <= not(layer2_outputs(265)) or (layer2_outputs(1566));
    layer3_outputs(661) <= not(layer2_outputs(79));
    layer3_outputs(662) <= (layer2_outputs(2012)) or (layer2_outputs(420));
    layer3_outputs(663) <= (layer2_outputs(343)) and not (layer2_outputs(176));
    layer3_outputs(664) <= not(layer2_outputs(242));
    layer3_outputs(665) <= not(layer2_outputs(823)) or (layer2_outputs(705));
    layer3_outputs(666) <= (layer2_outputs(897)) or (layer2_outputs(1846));
    layer3_outputs(667) <= not((layer2_outputs(866)) and (layer2_outputs(1921)));
    layer3_outputs(668) <= (layer2_outputs(1236)) and (layer2_outputs(170));
    layer3_outputs(669) <= not((layer2_outputs(2530)) or (layer2_outputs(531)));
    layer3_outputs(670) <= not(layer2_outputs(836)) or (layer2_outputs(1435));
    layer3_outputs(671) <= not(layer2_outputs(1439)) or (layer2_outputs(190));
    layer3_outputs(672) <= layer2_outputs(154);
    layer3_outputs(673) <= (layer2_outputs(262)) and (layer2_outputs(2191));
    layer3_outputs(674) <= '0';
    layer3_outputs(675) <= '1';
    layer3_outputs(676) <= not(layer2_outputs(1362));
    layer3_outputs(677) <= not(layer2_outputs(2323)) or (layer2_outputs(1541));
    layer3_outputs(678) <= '0';
    layer3_outputs(679) <= '0';
    layer3_outputs(680) <= (layer2_outputs(2206)) and not (layer2_outputs(1422));
    layer3_outputs(681) <= (layer2_outputs(610)) and (layer2_outputs(2196));
    layer3_outputs(682) <= not(layer2_outputs(471)) or (layer2_outputs(888));
    layer3_outputs(683) <= (layer2_outputs(51)) or (layer2_outputs(2332));
    layer3_outputs(684) <= not(layer2_outputs(864));
    layer3_outputs(685) <= '0';
    layer3_outputs(686) <= not((layer2_outputs(1391)) and (layer2_outputs(1527)));
    layer3_outputs(687) <= (layer2_outputs(780)) xor (layer2_outputs(1342));
    layer3_outputs(688) <= not((layer2_outputs(538)) or (layer2_outputs(2303)));
    layer3_outputs(689) <= (layer2_outputs(755)) and not (layer2_outputs(2232));
    layer3_outputs(690) <= not(layer2_outputs(1619));
    layer3_outputs(691) <= (layer2_outputs(1372)) and not (layer2_outputs(2299));
    layer3_outputs(692) <= '1';
    layer3_outputs(693) <= not((layer2_outputs(1279)) xor (layer2_outputs(1440)));
    layer3_outputs(694) <= not((layer2_outputs(2412)) xor (layer2_outputs(83)));
    layer3_outputs(695) <= '1';
    layer3_outputs(696) <= layer2_outputs(332);
    layer3_outputs(697) <= (layer2_outputs(2162)) and not (layer2_outputs(189));
    layer3_outputs(698) <= not((layer2_outputs(2390)) or (layer2_outputs(1605)));
    layer3_outputs(699) <= '0';
    layer3_outputs(700) <= layer2_outputs(1697);
    layer3_outputs(701) <= not((layer2_outputs(325)) or (layer2_outputs(583)));
    layer3_outputs(702) <= '1';
    layer3_outputs(703) <= layer2_outputs(2477);
    layer3_outputs(704) <= (layer2_outputs(1328)) and not (layer2_outputs(122));
    layer3_outputs(705) <= not(layer2_outputs(1470));
    layer3_outputs(706) <= (layer2_outputs(1427)) or (layer2_outputs(993));
    layer3_outputs(707) <= layer2_outputs(1174);
    layer3_outputs(708) <= (layer2_outputs(2154)) and not (layer2_outputs(344));
    layer3_outputs(709) <= (layer2_outputs(2286)) and not (layer2_outputs(1164));
    layer3_outputs(710) <= not(layer2_outputs(1132));
    layer3_outputs(711) <= '1';
    layer3_outputs(712) <= (layer2_outputs(1712)) and not (layer2_outputs(482));
    layer3_outputs(713) <= layer2_outputs(1177);
    layer3_outputs(714) <= '1';
    layer3_outputs(715) <= not((layer2_outputs(2344)) and (layer2_outputs(1082)));
    layer3_outputs(716) <= layer2_outputs(392);
    layer3_outputs(717) <= not(layer2_outputs(1544));
    layer3_outputs(718) <= not(layer2_outputs(58));
    layer3_outputs(719) <= (layer2_outputs(322)) and not (layer2_outputs(2188));
    layer3_outputs(720) <= layer2_outputs(1646);
    layer3_outputs(721) <= not(layer2_outputs(2060)) or (layer2_outputs(36));
    layer3_outputs(722) <= '1';
    layer3_outputs(723) <= layer2_outputs(1533);
    layer3_outputs(724) <= (layer2_outputs(2281)) or (layer2_outputs(1569));
    layer3_outputs(725) <= not(layer2_outputs(1269)) or (layer2_outputs(505));
    layer3_outputs(726) <= (layer2_outputs(2114)) and (layer2_outputs(70));
    layer3_outputs(727) <= not(layer2_outputs(2457));
    layer3_outputs(728) <= '0';
    layer3_outputs(729) <= (layer2_outputs(446)) and (layer2_outputs(1483));
    layer3_outputs(730) <= (layer2_outputs(2337)) and (layer2_outputs(2274));
    layer3_outputs(731) <= '0';
    layer3_outputs(732) <= layer2_outputs(2477);
    layer3_outputs(733) <= not((layer2_outputs(545)) or (layer2_outputs(797)));
    layer3_outputs(734) <= not(layer2_outputs(153));
    layer3_outputs(735) <= (layer2_outputs(1708)) xor (layer2_outputs(1352));
    layer3_outputs(736) <= '1';
    layer3_outputs(737) <= layer2_outputs(1694);
    layer3_outputs(738) <= layer2_outputs(1332);
    layer3_outputs(739) <= (layer2_outputs(1814)) and not (layer2_outputs(801));
    layer3_outputs(740) <= not(layer2_outputs(1434)) or (layer2_outputs(320));
    layer3_outputs(741) <= (layer2_outputs(963)) and (layer2_outputs(1957));
    layer3_outputs(742) <= not(layer2_outputs(785));
    layer3_outputs(743) <= '0';
    layer3_outputs(744) <= layer2_outputs(2396);
    layer3_outputs(745) <= not(layer2_outputs(1169)) or (layer2_outputs(1603));
    layer3_outputs(746) <= layer2_outputs(2424);
    layer3_outputs(747) <= layer2_outputs(1802);
    layer3_outputs(748) <= not(layer2_outputs(298));
    layer3_outputs(749) <= layer2_outputs(1183);
    layer3_outputs(750) <= not((layer2_outputs(1993)) xor (layer2_outputs(746)));
    layer3_outputs(751) <= '1';
    layer3_outputs(752) <= (layer2_outputs(1365)) and not (layer2_outputs(2372));
    layer3_outputs(753) <= not(layer2_outputs(1275));
    layer3_outputs(754) <= not(layer2_outputs(934));
    layer3_outputs(755) <= layer2_outputs(596);
    layer3_outputs(756) <= not(layer2_outputs(983)) or (layer2_outputs(1058));
    layer3_outputs(757) <= (layer2_outputs(474)) xor (layer2_outputs(1791));
    layer3_outputs(758) <= (layer2_outputs(2264)) and not (layer2_outputs(1829));
    layer3_outputs(759) <= not(layer2_outputs(1231)) or (layer2_outputs(1193));
    layer3_outputs(760) <= not((layer2_outputs(1764)) and (layer2_outputs(117)));
    layer3_outputs(761) <= (layer2_outputs(543)) and not (layer2_outputs(368));
    layer3_outputs(762) <= '0';
    layer3_outputs(763) <= not(layer2_outputs(1487)) or (layer2_outputs(2454));
    layer3_outputs(764) <= '0';
    layer3_outputs(765) <= (layer2_outputs(1947)) and not (layer2_outputs(1141));
    layer3_outputs(766) <= layer2_outputs(2427);
    layer3_outputs(767) <= (layer2_outputs(436)) or (layer2_outputs(364));
    layer3_outputs(768) <= layer2_outputs(210);
    layer3_outputs(769) <= (layer2_outputs(529)) or (layer2_outputs(165));
    layer3_outputs(770) <= not(layer2_outputs(398));
    layer3_outputs(771) <= not(layer2_outputs(665));
    layer3_outputs(772) <= (layer2_outputs(73)) and not (layer2_outputs(2033));
    layer3_outputs(773) <= (layer2_outputs(896)) and not (layer2_outputs(1755));
    layer3_outputs(774) <= not((layer2_outputs(1587)) and (layer2_outputs(2311)));
    layer3_outputs(775) <= not(layer2_outputs(1394)) or (layer2_outputs(1926));
    layer3_outputs(776) <= (layer2_outputs(392)) and not (layer2_outputs(853));
    layer3_outputs(777) <= not(layer2_outputs(411)) or (layer2_outputs(380));
    layer3_outputs(778) <= (layer2_outputs(1129)) and (layer2_outputs(1592));
    layer3_outputs(779) <= not(layer2_outputs(626)) or (layer2_outputs(2156));
    layer3_outputs(780) <= not(layer2_outputs(2434)) or (layer2_outputs(648));
    layer3_outputs(781) <= not((layer2_outputs(14)) or (layer2_outputs(711)));
    layer3_outputs(782) <= (layer2_outputs(761)) and (layer2_outputs(2263));
    layer3_outputs(783) <= '0';
    layer3_outputs(784) <= layer2_outputs(2310);
    layer3_outputs(785) <= not((layer2_outputs(1999)) or (layer2_outputs(697)));
    layer3_outputs(786) <= not((layer2_outputs(19)) or (layer2_outputs(2539)));
    layer3_outputs(787) <= not(layer2_outputs(2033)) or (layer2_outputs(1482));
    layer3_outputs(788) <= not(layer2_outputs(1500)) or (layer2_outputs(1086));
    layer3_outputs(789) <= not(layer2_outputs(2456)) or (layer2_outputs(1726));
    layer3_outputs(790) <= layer2_outputs(345);
    layer3_outputs(791) <= '0';
    layer3_outputs(792) <= (layer2_outputs(2458)) and not (layer2_outputs(1697));
    layer3_outputs(793) <= not(layer2_outputs(810)) or (layer2_outputs(2247));
    layer3_outputs(794) <= not(layer2_outputs(2480));
    layer3_outputs(795) <= '0';
    layer3_outputs(796) <= '0';
    layer3_outputs(797) <= (layer2_outputs(1958)) or (layer2_outputs(2326));
    layer3_outputs(798) <= '0';
    layer3_outputs(799) <= not((layer2_outputs(2429)) and (layer2_outputs(1341)));
    layer3_outputs(800) <= not(layer2_outputs(954)) or (layer2_outputs(878));
    layer3_outputs(801) <= not(layer2_outputs(17)) or (layer2_outputs(1125));
    layer3_outputs(802) <= (layer2_outputs(914)) and not (layer2_outputs(736));
    layer3_outputs(803) <= not((layer2_outputs(758)) or (layer2_outputs(1936)));
    layer3_outputs(804) <= (layer2_outputs(324)) and (layer2_outputs(2513));
    layer3_outputs(805) <= (layer2_outputs(2520)) and not (layer2_outputs(2132));
    layer3_outputs(806) <= not(layer2_outputs(2153));
    layer3_outputs(807) <= (layer2_outputs(1404)) and (layer2_outputs(911));
    layer3_outputs(808) <= (layer2_outputs(1455)) and not (layer2_outputs(1872));
    layer3_outputs(809) <= '1';
    layer3_outputs(810) <= (layer2_outputs(107)) and not (layer2_outputs(505));
    layer3_outputs(811) <= not(layer2_outputs(1586));
    layer3_outputs(812) <= (layer2_outputs(2367)) and not (layer2_outputs(489));
    layer3_outputs(813) <= not((layer2_outputs(2492)) and (layer2_outputs(1139)));
    layer3_outputs(814) <= layer2_outputs(2338);
    layer3_outputs(815) <= not(layer2_outputs(71));
    layer3_outputs(816) <= not(layer2_outputs(2006));
    layer3_outputs(817) <= not(layer2_outputs(7));
    layer3_outputs(818) <= not(layer2_outputs(2390));
    layer3_outputs(819) <= '1';
    layer3_outputs(820) <= layer2_outputs(2391);
    layer3_outputs(821) <= (layer2_outputs(1471)) and not (layer2_outputs(1312));
    layer3_outputs(822) <= layer2_outputs(875);
    layer3_outputs(823) <= layer2_outputs(1359);
    layer3_outputs(824) <= '1';
    layer3_outputs(825) <= (layer2_outputs(2534)) and not (layer2_outputs(1478));
    layer3_outputs(826) <= '1';
    layer3_outputs(827) <= layer2_outputs(934);
    layer3_outputs(828) <= not(layer2_outputs(192)) or (layer2_outputs(1152));
    layer3_outputs(829) <= layer2_outputs(1527);
    layer3_outputs(830) <= not((layer2_outputs(1888)) and (layer2_outputs(224)));
    layer3_outputs(831) <= (layer2_outputs(1549)) and not (layer2_outputs(513));
    layer3_outputs(832) <= '0';
    layer3_outputs(833) <= '1';
    layer3_outputs(834) <= (layer2_outputs(958)) and not (layer2_outputs(683));
    layer3_outputs(835) <= (layer2_outputs(185)) and not (layer2_outputs(321));
    layer3_outputs(836) <= not(layer2_outputs(1792));
    layer3_outputs(837) <= (layer2_outputs(1606)) and not (layer2_outputs(135));
    layer3_outputs(838) <= '1';
    layer3_outputs(839) <= layer2_outputs(201);
    layer3_outputs(840) <= not(layer2_outputs(2214));
    layer3_outputs(841) <= (layer2_outputs(787)) xor (layer2_outputs(1903));
    layer3_outputs(842) <= '1';
    layer3_outputs(843) <= not(layer2_outputs(137)) or (layer2_outputs(91));
    layer3_outputs(844) <= (layer2_outputs(341)) and not (layer2_outputs(1886));
    layer3_outputs(845) <= layer2_outputs(1404);
    layer3_outputs(846) <= not((layer2_outputs(327)) xor (layer2_outputs(2523)));
    layer3_outputs(847) <= not((layer2_outputs(673)) and (layer2_outputs(1687)));
    layer3_outputs(848) <= not(layer2_outputs(2252)) or (layer2_outputs(871));
    layer3_outputs(849) <= '0';
    layer3_outputs(850) <= (layer2_outputs(2455)) and not (layer2_outputs(1423));
    layer3_outputs(851) <= layer2_outputs(179);
    layer3_outputs(852) <= not(layer2_outputs(1920)) or (layer2_outputs(155));
    layer3_outputs(853) <= not(layer2_outputs(810));
    layer3_outputs(854) <= not((layer2_outputs(1258)) or (layer2_outputs(2193)));
    layer3_outputs(855) <= not(layer2_outputs(1080));
    layer3_outputs(856) <= (layer2_outputs(1408)) and (layer2_outputs(1449));
    layer3_outputs(857) <= layer2_outputs(1514);
    layer3_outputs(858) <= not(layer2_outputs(61));
    layer3_outputs(859) <= not(layer2_outputs(1381));
    layer3_outputs(860) <= layer2_outputs(2051);
    layer3_outputs(861) <= (layer2_outputs(2392)) and (layer2_outputs(762));
    layer3_outputs(862) <= '0';
    layer3_outputs(863) <= not(layer2_outputs(69)) or (layer2_outputs(1331));
    layer3_outputs(864) <= '0';
    layer3_outputs(865) <= not((layer2_outputs(90)) and (layer2_outputs(287)));
    layer3_outputs(866) <= not(layer2_outputs(1113)) or (layer2_outputs(1441));
    layer3_outputs(867) <= '1';
    layer3_outputs(868) <= not(layer2_outputs(1009)) or (layer2_outputs(865));
    layer3_outputs(869) <= (layer2_outputs(1987)) or (layer2_outputs(199));
    layer3_outputs(870) <= layer2_outputs(169);
    layer3_outputs(871) <= '1';
    layer3_outputs(872) <= (layer2_outputs(1183)) and (layer2_outputs(2121));
    layer3_outputs(873) <= not(layer2_outputs(1882)) or (layer2_outputs(1846));
    layer3_outputs(874) <= not(layer2_outputs(2112));
    layer3_outputs(875) <= layer2_outputs(1284);
    layer3_outputs(876) <= (layer2_outputs(1911)) and (layer2_outputs(2019));
    layer3_outputs(877) <= (layer2_outputs(2290)) and not (layer2_outputs(1885));
    layer3_outputs(878) <= (layer2_outputs(1430)) and (layer2_outputs(1094));
    layer3_outputs(879) <= layer2_outputs(515);
    layer3_outputs(880) <= layer2_outputs(879);
    layer3_outputs(881) <= not(layer2_outputs(816)) or (layer2_outputs(753));
    layer3_outputs(882) <= not(layer2_outputs(1665));
    layer3_outputs(883) <= (layer2_outputs(1769)) and not (layer2_outputs(719));
    layer3_outputs(884) <= '1';
    layer3_outputs(885) <= not(layer2_outputs(1669)) or (layer2_outputs(705));
    layer3_outputs(886) <= layer2_outputs(638);
    layer3_outputs(887) <= not((layer2_outputs(16)) and (layer2_outputs(434)));
    layer3_outputs(888) <= not((layer2_outputs(574)) or (layer2_outputs(1930)));
    layer3_outputs(889) <= not(layer2_outputs(2203)) or (layer2_outputs(2035));
    layer3_outputs(890) <= layer2_outputs(965);
    layer3_outputs(891) <= not(layer2_outputs(2542));
    layer3_outputs(892) <= not(layer2_outputs(921)) or (layer2_outputs(771));
    layer3_outputs(893) <= (layer2_outputs(1306)) or (layer2_outputs(539));
    layer3_outputs(894) <= '0';
    layer3_outputs(895) <= (layer2_outputs(1218)) and not (layer2_outputs(1104));
    layer3_outputs(896) <= not(layer2_outputs(2032));
    layer3_outputs(897) <= (layer2_outputs(303)) and (layer2_outputs(935));
    layer3_outputs(898) <= not((layer2_outputs(12)) xor (layer2_outputs(2011)));
    layer3_outputs(899) <= not((layer2_outputs(1849)) or (layer2_outputs(902)));
    layer3_outputs(900) <= '1';
    layer3_outputs(901) <= not((layer2_outputs(776)) or (layer2_outputs(1840)));
    layer3_outputs(902) <= not(layer2_outputs(301));
    layer3_outputs(903) <= (layer2_outputs(1439)) and (layer2_outputs(491));
    layer3_outputs(904) <= '1';
    layer3_outputs(905) <= (layer2_outputs(1938)) and (layer2_outputs(2516));
    layer3_outputs(906) <= not((layer2_outputs(921)) and (layer2_outputs(1808)));
    layer3_outputs(907) <= (layer2_outputs(1284)) and (layer2_outputs(1071));
    layer3_outputs(908) <= (layer2_outputs(893)) and not (layer2_outputs(545));
    layer3_outputs(909) <= (layer2_outputs(1267)) and not (layer2_outputs(2362));
    layer3_outputs(910) <= not((layer2_outputs(1817)) or (layer2_outputs(1967)));
    layer3_outputs(911) <= (layer2_outputs(738)) and not (layer2_outputs(1494));
    layer3_outputs(912) <= layer2_outputs(571);
    layer3_outputs(913) <= layer2_outputs(2319);
    layer3_outputs(914) <= layer2_outputs(2532);
    layer3_outputs(915) <= not((layer2_outputs(1739)) or (layer2_outputs(1243)));
    layer3_outputs(916) <= (layer2_outputs(686)) and not (layer2_outputs(812));
    layer3_outputs(917) <= '1';
    layer3_outputs(918) <= not((layer2_outputs(742)) or (layer2_outputs(977)));
    layer3_outputs(919) <= not(layer2_outputs(214));
    layer3_outputs(920) <= (layer2_outputs(1140)) and not (layer2_outputs(20));
    layer3_outputs(921) <= '1';
    layer3_outputs(922) <= '0';
    layer3_outputs(923) <= (layer2_outputs(2216)) and not (layer2_outputs(1893));
    layer3_outputs(924) <= not(layer2_outputs(562)) or (layer2_outputs(1069));
    layer3_outputs(925) <= layer2_outputs(313);
    layer3_outputs(926) <= not((layer2_outputs(548)) and (layer2_outputs(1935)));
    layer3_outputs(927) <= not((layer2_outputs(1986)) and (layer2_outputs(1092)));
    layer3_outputs(928) <= not(layer2_outputs(1904)) or (layer2_outputs(608));
    layer3_outputs(929) <= not((layer2_outputs(568)) or (layer2_outputs(611)));
    layer3_outputs(930) <= not(layer2_outputs(1250));
    layer3_outputs(931) <= layer2_outputs(275);
    layer3_outputs(932) <= not(layer2_outputs(279));
    layer3_outputs(933) <= '0';
    layer3_outputs(934) <= (layer2_outputs(1090)) and (layer2_outputs(827));
    layer3_outputs(935) <= not((layer2_outputs(728)) or (layer2_outputs(1671)));
    layer3_outputs(936) <= not(layer2_outputs(570));
    layer3_outputs(937) <= not(layer2_outputs(1082)) or (layer2_outputs(416));
    layer3_outputs(938) <= (layer2_outputs(1518)) and (layer2_outputs(1897));
    layer3_outputs(939) <= (layer2_outputs(1313)) and not (layer2_outputs(248));
    layer3_outputs(940) <= '1';
    layer3_outputs(941) <= not(layer2_outputs(286)) or (layer2_outputs(620));
    layer3_outputs(942) <= (layer2_outputs(472)) and not (layer2_outputs(2100));
    layer3_outputs(943) <= not(layer2_outputs(2501));
    layer3_outputs(944) <= not(layer2_outputs(2276));
    layer3_outputs(945) <= (layer2_outputs(1267)) or (layer2_outputs(1566));
    layer3_outputs(946) <= not(layer2_outputs(271));
    layer3_outputs(947) <= not((layer2_outputs(61)) xor (layer2_outputs(1010)));
    layer3_outputs(948) <= layer2_outputs(1635);
    layer3_outputs(949) <= (layer2_outputs(718)) or (layer2_outputs(1352));
    layer3_outputs(950) <= (layer2_outputs(2143)) or (layer2_outputs(1421));
    layer3_outputs(951) <= (layer2_outputs(2344)) and not (layer2_outputs(233));
    layer3_outputs(952) <= not(layer2_outputs(1316));
    layer3_outputs(953) <= layer2_outputs(200);
    layer3_outputs(954) <= not(layer2_outputs(1165));
    layer3_outputs(955) <= not((layer2_outputs(300)) or (layer2_outputs(658)));
    layer3_outputs(956) <= not(layer2_outputs(243)) or (layer2_outputs(171));
    layer3_outputs(957) <= (layer2_outputs(1482)) and not (layer2_outputs(1227));
    layer3_outputs(958) <= (layer2_outputs(1947)) and (layer2_outputs(1261));
    layer3_outputs(959) <= not((layer2_outputs(1290)) and (layer2_outputs(2360)));
    layer3_outputs(960) <= not((layer2_outputs(845)) or (layer2_outputs(1724)));
    layer3_outputs(961) <= not(layer2_outputs(683));
    layer3_outputs(962) <= not(layer2_outputs(509)) or (layer2_outputs(1163));
    layer3_outputs(963) <= not(layer2_outputs(1013));
    layer3_outputs(964) <= (layer2_outputs(1582)) and not (layer2_outputs(1946));
    layer3_outputs(965) <= not((layer2_outputs(115)) xor (layer2_outputs(766)));
    layer3_outputs(966) <= not((layer2_outputs(2417)) and (layer2_outputs(1658)));
    layer3_outputs(967) <= layer2_outputs(675);
    layer3_outputs(968) <= not(layer2_outputs(2046));
    layer3_outputs(969) <= not(layer2_outputs(2044));
    layer3_outputs(970) <= (layer2_outputs(1718)) or (layer2_outputs(1116));
    layer3_outputs(971) <= '1';
    layer3_outputs(972) <= not(layer2_outputs(1897));
    layer3_outputs(973) <= not((layer2_outputs(1297)) or (layer2_outputs(620)));
    layer3_outputs(974) <= layer2_outputs(2497);
    layer3_outputs(975) <= layer2_outputs(1875);
    layer3_outputs(976) <= layer2_outputs(1927);
    layer3_outputs(977) <= (layer2_outputs(1277)) or (layer2_outputs(22));
    layer3_outputs(978) <= not(layer2_outputs(1948)) or (layer2_outputs(1333));
    layer3_outputs(979) <= layer2_outputs(354);
    layer3_outputs(980) <= not(layer2_outputs(1848));
    layer3_outputs(981) <= not(layer2_outputs(1060)) or (layer2_outputs(1726));
    layer3_outputs(982) <= layer2_outputs(55);
    layer3_outputs(983) <= '0';
    layer3_outputs(984) <= not(layer2_outputs(286)) or (layer2_outputs(129));
    layer3_outputs(985) <= '1';
    layer3_outputs(986) <= not(layer2_outputs(856));
    layer3_outputs(987) <= not(layer2_outputs(773)) or (layer2_outputs(1585));
    layer3_outputs(988) <= not(layer2_outputs(2107));
    layer3_outputs(989) <= not((layer2_outputs(2179)) and (layer2_outputs(116)));
    layer3_outputs(990) <= not(layer2_outputs(2216)) or (layer2_outputs(1291));
    layer3_outputs(991) <= '1';
    layer3_outputs(992) <= not(layer2_outputs(537)) or (layer2_outputs(608));
    layer3_outputs(993) <= '0';
    layer3_outputs(994) <= not(layer2_outputs(1517));
    layer3_outputs(995) <= not(layer2_outputs(72));
    layer3_outputs(996) <= not(layer2_outputs(1606)) or (layer2_outputs(993));
    layer3_outputs(997) <= layer2_outputs(457);
    layer3_outputs(998) <= not(layer2_outputs(556)) or (layer2_outputs(2113));
    layer3_outputs(999) <= not(layer2_outputs(662)) or (layer2_outputs(1383));
    layer3_outputs(1000) <= (layer2_outputs(108)) or (layer2_outputs(549));
    layer3_outputs(1001) <= not(layer2_outputs(2109));
    layer3_outputs(1002) <= not(layer2_outputs(2433)) or (layer2_outputs(138));
    layer3_outputs(1003) <= layer2_outputs(1288);
    layer3_outputs(1004) <= (layer2_outputs(1581)) or (layer2_outputs(2017));
    layer3_outputs(1005) <= '0';
    layer3_outputs(1006) <= (layer2_outputs(2548)) and (layer2_outputs(1722));
    layer3_outputs(1007) <= '0';
    layer3_outputs(1008) <= not(layer2_outputs(1075));
    layer3_outputs(1009) <= (layer2_outputs(634)) or (layer2_outputs(1975));
    layer3_outputs(1010) <= (layer2_outputs(358)) or (layer2_outputs(1654));
    layer3_outputs(1011) <= not(layer2_outputs(912));
    layer3_outputs(1012) <= not(layer2_outputs(399));
    layer3_outputs(1013) <= '1';
    layer3_outputs(1014) <= '1';
    layer3_outputs(1015) <= (layer2_outputs(1796)) or (layer2_outputs(948));
    layer3_outputs(1016) <= not(layer2_outputs(767)) or (layer2_outputs(1189));
    layer3_outputs(1017) <= (layer2_outputs(1354)) and not (layer2_outputs(272));
    layer3_outputs(1018) <= (layer2_outputs(783)) or (layer2_outputs(1610));
    layer3_outputs(1019) <= not((layer2_outputs(1475)) or (layer2_outputs(1314)));
    layer3_outputs(1020) <= (layer2_outputs(1816)) and (layer2_outputs(1821));
    layer3_outputs(1021) <= not(layer2_outputs(1562)) or (layer2_outputs(91));
    layer3_outputs(1022) <= not(layer2_outputs(1529));
    layer3_outputs(1023) <= layer2_outputs(280);
    layer3_outputs(1024) <= not((layer2_outputs(391)) or (layer2_outputs(1360)));
    layer3_outputs(1025) <= '0';
    layer3_outputs(1026) <= not(layer2_outputs(2083));
    layer3_outputs(1027) <= (layer2_outputs(747)) and not (layer2_outputs(270));
    layer3_outputs(1028) <= not((layer2_outputs(483)) xor (layer2_outputs(2487)));
    layer3_outputs(1029) <= layer2_outputs(1523);
    layer3_outputs(1030) <= (layer2_outputs(1851)) and not (layer2_outputs(1771));
    layer3_outputs(1031) <= (layer2_outputs(1711)) and (layer2_outputs(699));
    layer3_outputs(1032) <= not(layer2_outputs(1834)) or (layer2_outputs(1841));
    layer3_outputs(1033) <= not(layer2_outputs(1198)) or (layer2_outputs(850));
    layer3_outputs(1034) <= not(layer2_outputs(1778));
    layer3_outputs(1035) <= not(layer2_outputs(476));
    layer3_outputs(1036) <= not(layer2_outputs(679));
    layer3_outputs(1037) <= layer2_outputs(716);
    layer3_outputs(1038) <= not(layer2_outputs(196)) or (layer2_outputs(1201));
    layer3_outputs(1039) <= not(layer2_outputs(1545));
    layer3_outputs(1040) <= not(layer2_outputs(442)) or (layer2_outputs(1311));
    layer3_outputs(1041) <= layer2_outputs(550);
    layer3_outputs(1042) <= not((layer2_outputs(73)) and (layer2_outputs(852)));
    layer3_outputs(1043) <= not(layer2_outputs(1529)) or (layer2_outputs(1265));
    layer3_outputs(1044) <= (layer2_outputs(2201)) and not (layer2_outputs(2005));
    layer3_outputs(1045) <= not(layer2_outputs(2125)) or (layer2_outputs(734));
    layer3_outputs(1046) <= not(layer2_outputs(997));
    layer3_outputs(1047) <= not(layer2_outputs(957));
    layer3_outputs(1048) <= (layer2_outputs(187)) and not (layer2_outputs(1570));
    layer3_outputs(1049) <= not(layer2_outputs(1931)) or (layer2_outputs(43));
    layer3_outputs(1050) <= not((layer2_outputs(1538)) or (layer2_outputs(200)));
    layer3_outputs(1051) <= '0';
    layer3_outputs(1052) <= (layer2_outputs(1437)) and (layer2_outputs(2421));
    layer3_outputs(1053) <= (layer2_outputs(1866)) and not (layer2_outputs(2508));
    layer3_outputs(1054) <= layer2_outputs(2428);
    layer3_outputs(1055) <= (layer2_outputs(1327)) and not (layer2_outputs(704));
    layer3_outputs(1056) <= (layer2_outputs(1385)) and not (layer2_outputs(1553));
    layer3_outputs(1057) <= '1';
    layer3_outputs(1058) <= (layer2_outputs(1345)) and not (layer2_outputs(1945));
    layer3_outputs(1059) <= '1';
    layer3_outputs(1060) <= not(layer2_outputs(2413));
    layer3_outputs(1061) <= not(layer2_outputs(280));
    layer3_outputs(1062) <= not(layer2_outputs(1541)) or (layer2_outputs(2443));
    layer3_outputs(1063) <= layer2_outputs(1575);
    layer3_outputs(1064) <= not(layer2_outputs(2327));
    layer3_outputs(1065) <= not(layer2_outputs(1245));
    layer3_outputs(1066) <= not(layer2_outputs(655));
    layer3_outputs(1067) <= not(layer2_outputs(872));
    layer3_outputs(1068) <= not(layer2_outputs(1110));
    layer3_outputs(1069) <= (layer2_outputs(1722)) and not (layer2_outputs(181));
    layer3_outputs(1070) <= '1';
    layer3_outputs(1071) <= layer2_outputs(1753);
    layer3_outputs(1072) <= not((layer2_outputs(2184)) or (layer2_outputs(1097)));
    layer3_outputs(1073) <= '0';
    layer3_outputs(1074) <= layer2_outputs(1392);
    layer3_outputs(1075) <= layer2_outputs(195);
    layer3_outputs(1076) <= layer2_outputs(1041);
    layer3_outputs(1077) <= '1';
    layer3_outputs(1078) <= not((layer2_outputs(0)) or (layer2_outputs(892)));
    layer3_outputs(1079) <= '1';
    layer3_outputs(1080) <= '1';
    layer3_outputs(1081) <= not(layer2_outputs(2085));
    layer3_outputs(1082) <= not((layer2_outputs(2511)) and (layer2_outputs(2168)));
    layer3_outputs(1083) <= '0';
    layer3_outputs(1084) <= layer2_outputs(1069);
    layer3_outputs(1085) <= not(layer2_outputs(2419));
    layer3_outputs(1086) <= '0';
    layer3_outputs(1087) <= layer2_outputs(1657);
    layer3_outputs(1088) <= '0';
    layer3_outputs(1089) <= '0';
    layer3_outputs(1090) <= not((layer2_outputs(1493)) or (layer2_outputs(278)));
    layer3_outputs(1091) <= layer2_outputs(1085);
    layer3_outputs(1092) <= layer2_outputs(702);
    layer3_outputs(1093) <= not(layer2_outputs(1914)) or (layer2_outputs(2479));
    layer3_outputs(1094) <= not(layer2_outputs(15)) or (layer2_outputs(1955));
    layer3_outputs(1095) <= layer2_outputs(1940);
    layer3_outputs(1096) <= layer2_outputs(1775);
    layer3_outputs(1097) <= '1';
    layer3_outputs(1098) <= not(layer2_outputs(2480)) or (layer2_outputs(1890));
    layer3_outputs(1099) <= (layer2_outputs(2512)) xor (layer2_outputs(407));
    layer3_outputs(1100) <= (layer2_outputs(113)) or (layer2_outputs(698));
    layer3_outputs(1101) <= '1';
    layer3_outputs(1102) <= layer2_outputs(708);
    layer3_outputs(1103) <= not((layer2_outputs(1900)) or (layer2_outputs(394)));
    layer3_outputs(1104) <= not(layer2_outputs(609));
    layer3_outputs(1105) <= (layer2_outputs(1513)) xor (layer2_outputs(1655));
    layer3_outputs(1106) <= not(layer2_outputs(1061)) or (layer2_outputs(1815));
    layer3_outputs(1107) <= (layer2_outputs(2010)) and not (layer2_outputs(1281));
    layer3_outputs(1108) <= not((layer2_outputs(241)) and (layer2_outputs(1773)));
    layer3_outputs(1109) <= not(layer2_outputs(2392)) or (layer2_outputs(820));
    layer3_outputs(1110) <= not((layer2_outputs(676)) and (layer2_outputs(2040)));
    layer3_outputs(1111) <= not(layer2_outputs(700));
    layer3_outputs(1112) <= not(layer2_outputs(765)) or (layer2_outputs(458));
    layer3_outputs(1113) <= (layer2_outputs(408)) or (layer2_outputs(984));
    layer3_outputs(1114) <= (layer2_outputs(1950)) and (layer2_outputs(659));
    layer3_outputs(1115) <= not((layer2_outputs(657)) or (layer2_outputs(803)));
    layer3_outputs(1116) <= not(layer2_outputs(77)) or (layer2_outputs(682));
    layer3_outputs(1117) <= (layer2_outputs(414)) and (layer2_outputs(437));
    layer3_outputs(1118) <= layer2_outputs(171);
    layer3_outputs(1119) <= layer2_outputs(1094);
    layer3_outputs(1120) <= (layer2_outputs(1216)) xor (layer2_outputs(263));
    layer3_outputs(1121) <= not(layer2_outputs(101));
    layer3_outputs(1122) <= layer2_outputs(162);
    layer3_outputs(1123) <= '1';
    layer3_outputs(1124) <= (layer2_outputs(2157)) or (layer2_outputs(461));
    layer3_outputs(1125) <= layer2_outputs(988);
    layer3_outputs(1126) <= '0';
    layer3_outputs(1127) <= not(layer2_outputs(986));
    layer3_outputs(1128) <= not((layer2_outputs(2459)) or (layer2_outputs(284)));
    layer3_outputs(1129) <= '0';
    layer3_outputs(1130) <= (layer2_outputs(388)) and not (layer2_outputs(2187));
    layer3_outputs(1131) <= not(layer2_outputs(186));
    layer3_outputs(1132) <= not((layer2_outputs(1855)) or (layer2_outputs(150)));
    layer3_outputs(1133) <= (layer2_outputs(613)) or (layer2_outputs(731));
    layer3_outputs(1134) <= (layer2_outputs(2371)) and not (layer2_outputs(1055));
    layer3_outputs(1135) <= (layer2_outputs(1333)) and (layer2_outputs(193));
    layer3_outputs(1136) <= not(layer2_outputs(996));
    layer3_outputs(1137) <= layer2_outputs(2105);
    layer3_outputs(1138) <= '0';
    layer3_outputs(1139) <= (layer2_outputs(376)) and not (layer2_outputs(377));
    layer3_outputs(1140) <= not(layer2_outputs(540));
    layer3_outputs(1141) <= not(layer2_outputs(1618));
    layer3_outputs(1142) <= (layer2_outputs(602)) and (layer2_outputs(1535));
    layer3_outputs(1143) <= layer2_outputs(156);
    layer3_outputs(1144) <= layer2_outputs(1535);
    layer3_outputs(1145) <= layer2_outputs(2416);
    layer3_outputs(1146) <= '0';
    layer3_outputs(1147) <= '1';
    layer3_outputs(1148) <= not(layer2_outputs(990)) or (layer2_outputs(1623));
    layer3_outputs(1149) <= not(layer2_outputs(2467)) or (layer2_outputs(1774));
    layer3_outputs(1150) <= not(layer2_outputs(746));
    layer3_outputs(1151) <= not(layer2_outputs(779));
    layer3_outputs(1152) <= (layer2_outputs(204)) or (layer2_outputs(1224));
    layer3_outputs(1153) <= '1';
    layer3_outputs(1154) <= not((layer2_outputs(678)) or (layer2_outputs(1366)));
    layer3_outputs(1155) <= layer2_outputs(648);
    layer3_outputs(1156) <= not(layer2_outputs(885)) or (layer2_outputs(1835));
    layer3_outputs(1157) <= layer2_outputs(1100);
    layer3_outputs(1158) <= not((layer2_outputs(1949)) or (layer2_outputs(1441)));
    layer3_outputs(1159) <= not(layer2_outputs(1255));
    layer3_outputs(1160) <= not(layer2_outputs(233)) or (layer2_outputs(1796));
    layer3_outputs(1161) <= '0';
    layer3_outputs(1162) <= not(layer2_outputs(2368));
    layer3_outputs(1163) <= layer2_outputs(586);
    layer3_outputs(1164) <= '0';
    layer3_outputs(1165) <= layer2_outputs(2275);
    layer3_outputs(1166) <= not(layer2_outputs(1191));
    layer3_outputs(1167) <= layer2_outputs(654);
    layer3_outputs(1168) <= not((layer2_outputs(1012)) and (layer2_outputs(2031)));
    layer3_outputs(1169) <= not(layer2_outputs(1062));
    layer3_outputs(1170) <= not(layer2_outputs(1695));
    layer3_outputs(1171) <= layer2_outputs(1806);
    layer3_outputs(1172) <= not(layer2_outputs(629));
    layer3_outputs(1173) <= (layer2_outputs(857)) and not (layer2_outputs(685));
    layer3_outputs(1174) <= (layer2_outputs(71)) and not (layer2_outputs(1361));
    layer3_outputs(1175) <= not((layer2_outputs(45)) or (layer2_outputs(1690)));
    layer3_outputs(1176) <= '1';
    layer3_outputs(1177) <= not((layer2_outputs(1905)) and (layer2_outputs(89)));
    layer3_outputs(1178) <= '1';
    layer3_outputs(1179) <= not(layer2_outputs(1323));
    layer3_outputs(1180) <= not(layer2_outputs(1820)) or (layer2_outputs(649));
    layer3_outputs(1181) <= (layer2_outputs(701)) or (layer2_outputs(1386));
    layer3_outputs(1182) <= (layer2_outputs(1215)) or (layer2_outputs(75));
    layer3_outputs(1183) <= (layer2_outputs(214)) and (layer2_outputs(2041));
    layer3_outputs(1184) <= not(layer2_outputs(410)) or (layer2_outputs(1661));
    layer3_outputs(1185) <= (layer2_outputs(1962)) or (layer2_outputs(1019));
    layer3_outputs(1186) <= (layer2_outputs(2468)) and (layer2_outputs(261));
    layer3_outputs(1187) <= '0';
    layer3_outputs(1188) <= not((layer2_outputs(537)) or (layer2_outputs(2314)));
    layer3_outputs(1189) <= not(layer2_outputs(1205)) or (layer2_outputs(1071));
    layer3_outputs(1190) <= not(layer2_outputs(2291));
    layer3_outputs(1191) <= (layer2_outputs(2460)) and not (layer2_outputs(242));
    layer3_outputs(1192) <= not(layer2_outputs(884));
    layer3_outputs(1193) <= '1';
    layer3_outputs(1194) <= layer2_outputs(2522);
    layer3_outputs(1195) <= '1';
    layer3_outputs(1196) <= not(layer2_outputs(2511)) or (layer2_outputs(2547));
    layer3_outputs(1197) <= not(layer2_outputs(2110)) or (layer2_outputs(744));
    layer3_outputs(1198) <= (layer2_outputs(2536)) and not (layer2_outputs(103));
    layer3_outputs(1199) <= not(layer2_outputs(1732)) or (layer2_outputs(2357));
    layer3_outputs(1200) <= not(layer2_outputs(2057)) or (layer2_outputs(395));
    layer3_outputs(1201) <= not(layer2_outputs(41));
    layer3_outputs(1202) <= not(layer2_outputs(1363));
    layer3_outputs(1203) <= (layer2_outputs(2401)) and not (layer2_outputs(485));
    layer3_outputs(1204) <= not((layer2_outputs(361)) and (layer2_outputs(1595)));
    layer3_outputs(1205) <= '0';
    layer3_outputs(1206) <= layer2_outputs(1400);
    layer3_outputs(1207) <= not(layer2_outputs(458));
    layer3_outputs(1208) <= layer2_outputs(1467);
    layer3_outputs(1209) <= '1';
    layer3_outputs(1210) <= (layer2_outputs(2524)) and (layer2_outputs(1364));
    layer3_outputs(1211) <= layer2_outputs(1128);
    layer3_outputs(1212) <= '0';
    layer3_outputs(1213) <= '0';
    layer3_outputs(1214) <= (layer2_outputs(1970)) and not (layer2_outputs(338));
    layer3_outputs(1215) <= (layer2_outputs(2472)) and not (layer2_outputs(567));
    layer3_outputs(1216) <= (layer2_outputs(2263)) and not (layer2_outputs(2198));
    layer3_outputs(1217) <= not(layer2_outputs(2463));
    layer3_outputs(1218) <= layer2_outputs(1899);
    layer3_outputs(1219) <= not(layer2_outputs(1112)) or (layer2_outputs(1757));
    layer3_outputs(1220) <= not(layer2_outputs(2152));
    layer3_outputs(1221) <= layer2_outputs(1077);
    layer3_outputs(1222) <= not((layer2_outputs(1017)) or (layer2_outputs(1589)));
    layer3_outputs(1223) <= not(layer2_outputs(23));
    layer3_outputs(1224) <= (layer2_outputs(554)) or (layer2_outputs(2029));
    layer3_outputs(1225) <= (layer2_outputs(1757)) or (layer2_outputs(1350));
    layer3_outputs(1226) <= (layer2_outputs(2515)) or (layer2_outputs(13));
    layer3_outputs(1227) <= layer2_outputs(1628);
    layer3_outputs(1228) <= '0';
    layer3_outputs(1229) <= layer2_outputs(2172);
    layer3_outputs(1230) <= not(layer2_outputs(449)) or (layer2_outputs(632));
    layer3_outputs(1231) <= not(layer2_outputs(1334));
    layer3_outputs(1232) <= not((layer2_outputs(1133)) xor (layer2_outputs(1959)));
    layer3_outputs(1233) <= (layer2_outputs(604)) or (layer2_outputs(2503));
    layer3_outputs(1234) <= layer2_outputs(474);
    layer3_outputs(1235) <= not(layer2_outputs(2037));
    layer3_outputs(1236) <= not(layer2_outputs(1298));
    layer3_outputs(1237) <= (layer2_outputs(783)) and (layer2_outputs(1230));
    layer3_outputs(1238) <= (layer2_outputs(1461)) and not (layer2_outputs(670));
    layer3_outputs(1239) <= not((layer2_outputs(1465)) or (layer2_outputs(1522)));
    layer3_outputs(1240) <= not(layer2_outputs(385)) or (layer2_outputs(289));
    layer3_outputs(1241) <= '0';
    layer3_outputs(1242) <= (layer2_outputs(2129)) and not (layer2_outputs(1036));
    layer3_outputs(1243) <= layer2_outputs(780);
    layer3_outputs(1244) <= not(layer2_outputs(1064)) or (layer2_outputs(1239));
    layer3_outputs(1245) <= not(layer2_outputs(999)) or (layer2_outputs(504));
    layer3_outputs(1246) <= (layer2_outputs(781)) and (layer2_outputs(2554));
    layer3_outputs(1247) <= not((layer2_outputs(614)) or (layer2_outputs(450)));
    layer3_outputs(1248) <= layer2_outputs(691);
    layer3_outputs(1249) <= not(layer2_outputs(250)) or (layer2_outputs(1460));
    layer3_outputs(1250) <= layer2_outputs(76);
    layer3_outputs(1251) <= (layer2_outputs(2237)) and (layer2_outputs(547));
    layer3_outputs(1252) <= not(layer2_outputs(387));
    layer3_outputs(1253) <= not(layer2_outputs(2124));
    layer3_outputs(1254) <= layer2_outputs(1995);
    layer3_outputs(1255) <= (layer2_outputs(2446)) xor (layer2_outputs(1256));
    layer3_outputs(1256) <= (layer2_outputs(2328)) and not (layer2_outputs(2047));
    layer3_outputs(1257) <= (layer2_outputs(2311)) and (layer2_outputs(1005));
    layer3_outputs(1258) <= not(layer2_outputs(402));
    layer3_outputs(1259) <= not((layer2_outputs(588)) or (layer2_outputs(1543)));
    layer3_outputs(1260) <= '0';
    layer3_outputs(1261) <= '1';
    layer3_outputs(1262) <= layer2_outputs(2315);
    layer3_outputs(1263) <= not(layer2_outputs(1481)) or (layer2_outputs(225));
    layer3_outputs(1264) <= '1';
    layer3_outputs(1265) <= (layer2_outputs(240)) and (layer2_outputs(2455));
    layer3_outputs(1266) <= '0';
    layer3_outputs(1267) <= (layer2_outputs(1842)) and not (layer2_outputs(2310));
    layer3_outputs(1268) <= layer2_outputs(2438);
    layer3_outputs(1269) <= not(layer2_outputs(1735));
    layer3_outputs(1270) <= not(layer2_outputs(1375));
    layer3_outputs(1271) <= not((layer2_outputs(307)) or (layer2_outputs(1480)));
    layer3_outputs(1272) <= (layer2_outputs(2001)) and (layer2_outputs(331));
    layer3_outputs(1273) <= not((layer2_outputs(1679)) xor (layer2_outputs(568)));
    layer3_outputs(1274) <= '0';
    layer3_outputs(1275) <= layer2_outputs(1799);
    layer3_outputs(1276) <= not((layer2_outputs(32)) or (layer2_outputs(1963)));
    layer3_outputs(1277) <= not(layer2_outputs(849)) or (layer2_outputs(1270));
    layer3_outputs(1278) <= '1';
    layer3_outputs(1279) <= '0';
    layer3_outputs(1280) <= layer2_outputs(679);
    layer3_outputs(1281) <= (layer2_outputs(353)) or (layer2_outputs(2183));
    layer3_outputs(1282) <= (layer2_outputs(1332)) and not (layer2_outputs(1502));
    layer3_outputs(1283) <= layer2_outputs(1188);
    layer3_outputs(1284) <= not((layer2_outputs(212)) or (layer2_outputs(1512)));
    layer3_outputs(1285) <= '1';
    layer3_outputs(1286) <= not((layer2_outputs(2103)) and (layer2_outputs(30)));
    layer3_outputs(1287) <= not(layer2_outputs(1244)) or (layer2_outputs(1207));
    layer3_outputs(1288) <= not(layer2_outputs(506));
    layer3_outputs(1289) <= '1';
    layer3_outputs(1290) <= (layer2_outputs(2555)) and not (layer2_outputs(1016));
    layer3_outputs(1291) <= not(layer2_outputs(1513)) or (layer2_outputs(468));
    layer3_outputs(1292) <= (layer2_outputs(1446)) or (layer2_outputs(2421));
    layer3_outputs(1293) <= layer2_outputs(239);
    layer3_outputs(1294) <= '1';
    layer3_outputs(1295) <= not(layer2_outputs(2100)) or (layer2_outputs(1680));
    layer3_outputs(1296) <= layer2_outputs(236);
    layer3_outputs(1297) <= not(layer2_outputs(6));
    layer3_outputs(1298) <= (layer2_outputs(1234)) or (layer2_outputs(2042));
    layer3_outputs(1299) <= not(layer2_outputs(1051));
    layer3_outputs(1300) <= not((layer2_outputs(501)) and (layer2_outputs(1982)));
    layer3_outputs(1301) <= not((layer2_outputs(1994)) and (layer2_outputs(2095)));
    layer3_outputs(1302) <= '1';
    layer3_outputs(1303) <= not(layer2_outputs(2359)) or (layer2_outputs(742));
    layer3_outputs(1304) <= layer2_outputs(2444);
    layer3_outputs(1305) <= not(layer2_outputs(303)) or (layer2_outputs(2490));
    layer3_outputs(1306) <= not(layer2_outputs(2224));
    layer3_outputs(1307) <= not(layer2_outputs(2369)) or (layer2_outputs(1884));
    layer3_outputs(1308) <= (layer2_outputs(2173)) or (layer2_outputs(2214));
    layer3_outputs(1309) <= not(layer2_outputs(1614));
    layer3_outputs(1310) <= '0';
    layer3_outputs(1311) <= layer2_outputs(2408);
    layer3_outputs(1312) <= (layer2_outputs(2169)) or (layer2_outputs(226));
    layer3_outputs(1313) <= not(layer2_outputs(2541));
    layer3_outputs(1314) <= not(layer2_outputs(1908));
    layer3_outputs(1315) <= (layer2_outputs(276)) and not (layer2_outputs(956));
    layer3_outputs(1316) <= not(layer2_outputs(472));
    layer3_outputs(1317) <= layer2_outputs(139);
    layer3_outputs(1318) <= '0';
    layer3_outputs(1319) <= (layer2_outputs(1665)) xor (layer2_outputs(1160));
    layer3_outputs(1320) <= layer2_outputs(982);
    layer3_outputs(1321) <= not(layer2_outputs(2052)) or (layer2_outputs(666));
    layer3_outputs(1322) <= not((layer2_outputs(1306)) or (layer2_outputs(1910)));
    layer3_outputs(1323) <= not((layer2_outputs(1473)) and (layer2_outputs(1721)));
    layer3_outputs(1324) <= '0';
    layer3_outputs(1325) <= not((layer2_outputs(1075)) xor (layer2_outputs(2252)));
    layer3_outputs(1326) <= not(layer2_outputs(199));
    layer3_outputs(1327) <= not((layer2_outputs(2127)) or (layer2_outputs(2317)));
    layer3_outputs(1328) <= not((layer2_outputs(220)) or (layer2_outputs(1832)));
    layer3_outputs(1329) <= not(layer2_outputs(1299));
    layer3_outputs(1330) <= (layer2_outputs(76)) and not (layer2_outputs(779));
    layer3_outputs(1331) <= layer2_outputs(1847);
    layer3_outputs(1332) <= not(layer2_outputs(2374)) or (layer2_outputs(62));
    layer3_outputs(1333) <= (layer2_outputs(1431)) or (layer2_outputs(2532));
    layer3_outputs(1334) <= not(layer2_outputs(665));
    layer3_outputs(1335) <= (layer2_outputs(2427)) and not (layer2_outputs(1109));
    layer3_outputs(1336) <= (layer2_outputs(1099)) and not (layer2_outputs(105));
    layer3_outputs(1337) <= (layer2_outputs(452)) and (layer2_outputs(467));
    layer3_outputs(1338) <= not((layer2_outputs(1686)) and (layer2_outputs(998)));
    layer3_outputs(1339) <= not((layer2_outputs(809)) and (layer2_outputs(2068)));
    layer3_outputs(1340) <= layer2_outputs(1348);
    layer3_outputs(1341) <= not(layer2_outputs(2424));
    layer3_outputs(1342) <= (layer2_outputs(1110)) and not (layer2_outputs(791));
    layer3_outputs(1343) <= (layer2_outputs(1503)) or (layer2_outputs(1033));
    layer3_outputs(1344) <= layer2_outputs(1398);
    layer3_outputs(1345) <= not(layer2_outputs(899));
    layer3_outputs(1346) <= not(layer2_outputs(397)) or (layer2_outputs(2507));
    layer3_outputs(1347) <= not(layer2_outputs(2038)) or (layer2_outputs(1997));
    layer3_outputs(1348) <= not(layer2_outputs(1489));
    layer3_outputs(1349) <= not((layer2_outputs(1337)) and (layer2_outputs(1823)));
    layer3_outputs(1350) <= not(layer2_outputs(1378));
    layer3_outputs(1351) <= '0';
    layer3_outputs(1352) <= '0';
    layer3_outputs(1353) <= layer2_outputs(1308);
    layer3_outputs(1354) <= (layer2_outputs(1635)) xor (layer2_outputs(1330));
    layer3_outputs(1355) <= (layer2_outputs(2096)) and (layer2_outputs(605));
    layer3_outputs(1356) <= layer2_outputs(4);
    layer3_outputs(1357) <= not(layer2_outputs(847));
    layer3_outputs(1358) <= '0';
    layer3_outputs(1359) <= (layer2_outputs(98)) or (layer2_outputs(958));
    layer3_outputs(1360) <= '1';
    layer3_outputs(1361) <= not((layer2_outputs(1991)) or (layer2_outputs(177)));
    layer3_outputs(1362) <= not(layer2_outputs(2405));
    layer3_outputs(1363) <= not(layer2_outputs(2444));
    layer3_outputs(1364) <= layer2_outputs(1050);
    layer3_outputs(1365) <= not(layer2_outputs(923)) or (layer2_outputs(2277));
    layer3_outputs(1366) <= layer2_outputs(2221);
    layer3_outputs(1367) <= '0';
    layer3_outputs(1368) <= layer2_outputs(2478);
    layer3_outputs(1369) <= not(layer2_outputs(547)) or (layer2_outputs(1353));
    layer3_outputs(1370) <= (layer2_outputs(1822)) and (layer2_outputs(898));
    layer3_outputs(1371) <= '0';
    layer3_outputs(1372) <= (layer2_outputs(2407)) and not (layer2_outputs(1956));
    layer3_outputs(1373) <= not(layer2_outputs(1979));
    layer3_outputs(1374) <= (layer2_outputs(441)) xor (layer2_outputs(2210));
    layer3_outputs(1375) <= layer2_outputs(1158);
    layer3_outputs(1376) <= layer2_outputs(974);
    layer3_outputs(1377) <= '0';
    layer3_outputs(1378) <= not(layer2_outputs(2397)) or (layer2_outputs(593));
    layer3_outputs(1379) <= not(layer2_outputs(2136));
    layer3_outputs(1380) <= not(layer2_outputs(1678));
    layer3_outputs(1381) <= '0';
    layer3_outputs(1382) <= layer2_outputs(973);
    layer3_outputs(1383) <= layer2_outputs(1434);
    layer3_outputs(1384) <= not(layer2_outputs(362));
    layer3_outputs(1385) <= not(layer2_outputs(681));
    layer3_outputs(1386) <= (layer2_outputs(1979)) and (layer2_outputs(340));
    layer3_outputs(1387) <= (layer2_outputs(2375)) and (layer2_outputs(2487));
    layer3_outputs(1388) <= not(layer2_outputs(2142));
    layer3_outputs(1389) <= layer2_outputs(531);
    layer3_outputs(1390) <= not(layer2_outputs(2084)) or (layer2_outputs(2296));
    layer3_outputs(1391) <= not((layer2_outputs(1286)) and (layer2_outputs(169)));
    layer3_outputs(1392) <= '1';
    layer3_outputs(1393) <= layer2_outputs(2542);
    layer3_outputs(1394) <= not(layer2_outputs(2175));
    layer3_outputs(1395) <= not(layer2_outputs(2447));
    layer3_outputs(1396) <= '1';
    layer3_outputs(1397) <= not(layer2_outputs(1935));
    layer3_outputs(1398) <= not(layer2_outputs(530));
    layer3_outputs(1399) <= not(layer2_outputs(2400));
    layer3_outputs(1400) <= not((layer2_outputs(102)) and (layer2_outputs(1466)));
    layer3_outputs(1401) <= not((layer2_outputs(1114)) and (layer2_outputs(1989)));
    layer3_outputs(1402) <= not(layer2_outputs(1177));
    layer3_outputs(1403) <= layer2_outputs(585);
    layer3_outputs(1404) <= (layer2_outputs(1889)) and not (layer2_outputs(2507));
    layer3_outputs(1405) <= (layer2_outputs(141)) and not (layer2_outputs(1751));
    layer3_outputs(1406) <= (layer2_outputs(1399)) and not (layer2_outputs(2089));
    layer3_outputs(1407) <= not((layer2_outputs(973)) or (layer2_outputs(2423)));
    layer3_outputs(1408) <= not(layer2_outputs(1501));
    layer3_outputs(1409) <= (layer2_outputs(1988)) and not (layer2_outputs(444));
    layer3_outputs(1410) <= '1';
    layer3_outputs(1411) <= not(layer2_outputs(2544)) or (layer2_outputs(576));
    layer3_outputs(1412) <= (layer2_outputs(1699)) and (layer2_outputs(2492));
    layer3_outputs(1413) <= (layer2_outputs(564)) and not (layer2_outputs(1020));
    layer3_outputs(1414) <= not(layer2_outputs(2363)) or (layer2_outputs(2387));
    layer3_outputs(1415) <= not((layer2_outputs(2506)) and (layer2_outputs(2541)));
    layer3_outputs(1416) <= not(layer2_outputs(2345));
    layer3_outputs(1417) <= not((layer2_outputs(427)) or (layer2_outputs(180)));
    layer3_outputs(1418) <= not(layer2_outputs(629));
    layer3_outputs(1419) <= not(layer2_outputs(351)) or (layer2_outputs(1036));
    layer3_outputs(1420) <= layer2_outputs(1504);
    layer3_outputs(1421) <= (layer2_outputs(1135)) and not (layer2_outputs(1874));
    layer3_outputs(1422) <= layer2_outputs(1809);
    layer3_outputs(1423) <= layer2_outputs(251);
    layer3_outputs(1424) <= '0';
    layer3_outputs(1425) <= (layer2_outputs(207)) or (layer2_outputs(1004));
    layer3_outputs(1426) <= not((layer2_outputs(2102)) or (layer2_outputs(2117)));
    layer3_outputs(1427) <= (layer2_outputs(402)) and not (layer2_outputs(1099));
    layer3_outputs(1428) <= not((layer2_outputs(2498)) or (layer2_outputs(481)));
    layer3_outputs(1429) <= not(layer2_outputs(245));
    layer3_outputs(1430) <= not(layer2_outputs(2087));
    layer3_outputs(1431) <= layer2_outputs(315);
    layer3_outputs(1432) <= '1';
    layer3_outputs(1433) <= not(layer2_outputs(2114)) or (layer2_outputs(277));
    layer3_outputs(1434) <= (layer2_outputs(291)) or (layer2_outputs(1754));
    layer3_outputs(1435) <= not(layer2_outputs(427));
    layer3_outputs(1436) <= not(layer2_outputs(2268)) or (layer2_outputs(1859));
    layer3_outputs(1437) <= not((layer2_outputs(1315)) or (layer2_outputs(1292)));
    layer3_outputs(1438) <= not((layer2_outputs(1794)) and (layer2_outputs(104)));
    layer3_outputs(1439) <= (layer2_outputs(689)) and not (layer2_outputs(2237));
    layer3_outputs(1440) <= '0';
    layer3_outputs(1441) <= '0';
    layer3_outputs(1442) <= '0';
    layer3_outputs(1443) <= layer2_outputs(2238);
    layer3_outputs(1444) <= (layer2_outputs(843)) and not (layer2_outputs(1854));
    layer3_outputs(1445) <= (layer2_outputs(345)) and not (layer2_outputs(1000));
    layer3_outputs(1446) <= not(layer2_outputs(1972));
    layer3_outputs(1447) <= layer2_outputs(740);
    layer3_outputs(1448) <= (layer2_outputs(445)) and not (layer2_outputs(37));
    layer3_outputs(1449) <= layer2_outputs(490);
    layer3_outputs(1450) <= layer2_outputs(782);
    layer3_outputs(1451) <= '0';
    layer3_outputs(1452) <= not(layer2_outputs(846)) or (layer2_outputs(799));
    layer3_outputs(1453) <= not(layer2_outputs(188)) or (layer2_outputs(1495));
    layer3_outputs(1454) <= not(layer2_outputs(590));
    layer3_outputs(1455) <= (layer2_outputs(2461)) and not (layer2_outputs(498));
    layer3_outputs(1456) <= not((layer2_outputs(2365)) and (layer2_outputs(1339)));
    layer3_outputs(1457) <= layer2_outputs(1508);
    layer3_outputs(1458) <= not((layer2_outputs(1433)) and (layer2_outputs(2076)));
    layer3_outputs(1459) <= '1';
    layer3_outputs(1460) <= not(layer2_outputs(1798)) or (layer2_outputs(175));
    layer3_outputs(1461) <= not(layer2_outputs(1136));
    layer3_outputs(1462) <= not((layer2_outputs(1548)) and (layer2_outputs(1263)));
    layer3_outputs(1463) <= not(layer2_outputs(1640)) or (layer2_outputs(1246));
    layer3_outputs(1464) <= not((layer2_outputs(1682)) or (layer2_outputs(835)));
    layer3_outputs(1465) <= not((layer2_outputs(835)) or (layer2_outputs(1193)));
    layer3_outputs(1466) <= (layer2_outputs(862)) and not (layer2_outputs(2182));
    layer3_outputs(1467) <= (layer2_outputs(2486)) and (layer2_outputs(2558));
    layer3_outputs(1468) <= not((layer2_outputs(798)) xor (layer2_outputs(1971)));
    layer3_outputs(1469) <= not(layer2_outputs(40));
    layer3_outputs(1470) <= layer2_outputs(945);
    layer3_outputs(1471) <= (layer2_outputs(1728)) and (layer2_outputs(2549));
    layer3_outputs(1472) <= '1';
    layer3_outputs(1473) <= (layer2_outputs(2132)) and not (layer2_outputs(2351));
    layer3_outputs(1474) <= not(layer2_outputs(2209)) or (layer2_outputs(1144));
    layer3_outputs(1475) <= not(layer2_outputs(924)) or (layer2_outputs(833));
    layer3_outputs(1476) <= not(layer2_outputs(1869));
    layer3_outputs(1477) <= not(layer2_outputs(406)) or (layer2_outputs(172));
    layer3_outputs(1478) <= not((layer2_outputs(1030)) and (layer2_outputs(745)));
    layer3_outputs(1479) <= '1';
    layer3_outputs(1480) <= '0';
    layer3_outputs(1481) <= (layer2_outputs(988)) and not (layer2_outputs(1534));
    layer3_outputs(1482) <= layer2_outputs(1538);
    layer3_outputs(1483) <= not(layer2_outputs(804));
    layer3_outputs(1484) <= layer2_outputs(523);
    layer3_outputs(1485) <= '1';
    layer3_outputs(1486) <= not(layer2_outputs(486)) or (layer2_outputs(413));
    layer3_outputs(1487) <= not(layer2_outputs(277));
    layer3_outputs(1488) <= not((layer2_outputs(1762)) or (layer2_outputs(482)));
    layer3_outputs(1489) <= not((layer2_outputs(2559)) and (layer2_outputs(1775)));
    layer3_outputs(1490) <= layer2_outputs(463);
    layer3_outputs(1491) <= (layer2_outputs(2379)) xor (layer2_outputs(1515));
    layer3_outputs(1492) <= not(layer2_outputs(1384)) or (layer2_outputs(1249));
    layer3_outputs(1493) <= layer2_outputs(1735);
    layer3_outputs(1494) <= layer2_outputs(653);
    layer3_outputs(1495) <= (layer2_outputs(995)) or (layer2_outputs(1547));
    layer3_outputs(1496) <= not((layer2_outputs(1170)) or (layer2_outputs(917)));
    layer3_outputs(1497) <= not(layer2_outputs(1843));
    layer3_outputs(1498) <= not(layer2_outputs(381));
    layer3_outputs(1499) <= (layer2_outputs(496)) or (layer2_outputs(2090));
    layer3_outputs(1500) <= not(layer2_outputs(1833));
    layer3_outputs(1501) <= layer2_outputs(1040);
    layer3_outputs(1502) <= not((layer2_outputs(185)) or (layer2_outputs(2134)));
    layer3_outputs(1503) <= not(layer2_outputs(1058));
    layer3_outputs(1504) <= '0';
    layer3_outputs(1505) <= '0';
    layer3_outputs(1506) <= '1';
    layer3_outputs(1507) <= '0';
    layer3_outputs(1508) <= not(layer2_outputs(2452));
    layer3_outputs(1509) <= layer2_outputs(2186);
    layer3_outputs(1510) <= '1';
    layer3_outputs(1511) <= layer2_outputs(1753);
    layer3_outputs(1512) <= not((layer2_outputs(2318)) and (layer2_outputs(737)));
    layer3_outputs(1513) <= not((layer2_outputs(732)) and (layer2_outputs(695)));
    layer3_outputs(1514) <= not((layer2_outputs(1055)) xor (layer2_outputs(932)));
    layer3_outputs(1515) <= not(layer2_outputs(1167));
    layer3_outputs(1516) <= layer2_outputs(2291);
    layer3_outputs(1517) <= not(layer2_outputs(2082));
    layer3_outputs(1518) <= layer2_outputs(72);
    layer3_outputs(1519) <= layer2_outputs(306);
    layer3_outputs(1520) <= layer2_outputs(1772);
    layer3_outputs(1521) <= (layer2_outputs(549)) and not (layer2_outputs(1645));
    layer3_outputs(1522) <= layer2_outputs(2354);
    layer3_outputs(1523) <= not(layer2_outputs(187));
    layer3_outputs(1524) <= (layer2_outputs(694)) and not (layer2_outputs(1045));
    layer3_outputs(1525) <= (layer2_outputs(1540)) and not (layer2_outputs(866));
    layer3_outputs(1526) <= '0';
    layer3_outputs(1527) <= not((layer2_outputs(386)) xor (layer2_outputs(550)));
    layer3_outputs(1528) <= not(layer2_outputs(46));
    layer3_outputs(1529) <= not((layer2_outputs(440)) and (layer2_outputs(762)));
    layer3_outputs(1530) <= (layer2_outputs(371)) or (layer2_outputs(2253));
    layer3_outputs(1531) <= not((layer2_outputs(313)) and (layer2_outputs(1178)));
    layer3_outputs(1532) <= not((layer2_outputs(981)) or (layer2_outputs(1354)));
    layer3_outputs(1533) <= not(layer2_outputs(477));
    layer3_outputs(1534) <= (layer2_outputs(2270)) and not (layer2_outputs(2321));
    layer3_outputs(1535) <= not(layer2_outputs(2206));
    layer3_outputs(1536) <= not(layer2_outputs(808));
    layer3_outputs(1537) <= not((layer2_outputs(818)) or (layer2_outputs(1258)));
    layer3_outputs(1538) <= not(layer2_outputs(1017)) or (layer2_outputs(1727));
    layer3_outputs(1539) <= not(layer2_outputs(992));
    layer3_outputs(1540) <= (layer2_outputs(131)) and not (layer2_outputs(1685));
    layer3_outputs(1541) <= not(layer2_outputs(554)) or (layer2_outputs(1235));
    layer3_outputs(1542) <= layer2_outputs(1295);
    layer3_outputs(1543) <= (layer2_outputs(1923)) and not (layer2_outputs(2502));
    layer3_outputs(1544) <= not(layer2_outputs(89));
    layer3_outputs(1545) <= (layer2_outputs(1838)) and not (layer2_outputs(1578));
    layer3_outputs(1546) <= layer2_outputs(1132);
    layer3_outputs(1547) <= not(layer2_outputs(2497)) or (layer2_outputs(572));
    layer3_outputs(1548) <= not(layer2_outputs(2527)) or (layer2_outputs(1096));
    layer3_outputs(1549) <= '1';
    layer3_outputs(1550) <= not(layer2_outputs(2285)) or (layer2_outputs(882));
    layer3_outputs(1551) <= (layer2_outputs(1996)) and (layer2_outputs(1715));
    layer3_outputs(1552) <= (layer2_outputs(1260)) and not (layer2_outputs(759));
    layer3_outputs(1553) <= not((layer2_outputs(1698)) and (layer2_outputs(1001)));
    layer3_outputs(1554) <= '0';
    layer3_outputs(1555) <= '1';
    layer3_outputs(1556) <= not(layer2_outputs(863));
    layer3_outputs(1557) <= not((layer2_outputs(1725)) or (layer2_outputs(452)));
    layer3_outputs(1558) <= layer2_outputs(438);
    layer3_outputs(1559) <= not((layer2_outputs(2099)) or (layer2_outputs(1861)));
    layer3_outputs(1560) <= not(layer2_outputs(1485));
    layer3_outputs(1561) <= not(layer2_outputs(1325)) or (layer2_outputs(1296));
    layer3_outputs(1562) <= (layer2_outputs(815)) and (layer2_outputs(938));
    layer3_outputs(1563) <= (layer2_outputs(497)) and (layer2_outputs(1729));
    layer3_outputs(1564) <= not(layer2_outputs(2011)) or (layer2_outputs(2518));
    layer3_outputs(1565) <= (layer2_outputs(1429)) and (layer2_outputs(1406));
    layer3_outputs(1566) <= not(layer2_outputs(363));
    layer3_outputs(1567) <= layer2_outputs(1773);
    layer3_outputs(1568) <= not((layer2_outputs(687)) or (layer2_outputs(1195)));
    layer3_outputs(1569) <= (layer2_outputs(1830)) and not (layer2_outputs(1741));
    layer3_outputs(1570) <= layer2_outputs(184);
    layer3_outputs(1571) <= not(layer2_outputs(1182)) or (layer2_outputs(2207));
    layer3_outputs(1572) <= not((layer2_outputs(1561)) or (layer2_outputs(1207)));
    layer3_outputs(1573) <= layer2_outputs(643);
    layer3_outputs(1574) <= not(layer2_outputs(2202)) or (layer2_outputs(2102));
    layer3_outputs(1575) <= not((layer2_outputs(1536)) and (layer2_outputs(669)));
    layer3_outputs(1576) <= not(layer2_outputs(2174));
    layer3_outputs(1577) <= not((layer2_outputs(2050)) or (layer2_outputs(2198)));
    layer3_outputs(1578) <= (layer2_outputs(2073)) and not (layer2_outputs(257));
    layer3_outputs(1579) <= not(layer2_outputs(1772));
    layer3_outputs(1580) <= (layer2_outputs(875)) and not (layer2_outputs(1648));
    layer3_outputs(1581) <= (layer2_outputs(1553)) or (layer2_outputs(2234));
    layer3_outputs(1582) <= '0';
    layer3_outputs(1583) <= (layer2_outputs(1369)) and not (layer2_outputs(2489));
    layer3_outputs(1584) <= not(layer2_outputs(2413)) or (layer2_outputs(381));
    layer3_outputs(1585) <= layer2_outputs(1360);
    layer3_outputs(1586) <= not(layer2_outputs(793));
    layer3_outputs(1587) <= not(layer2_outputs(1119)) or (layer2_outputs(454));
    layer3_outputs(1588) <= not(layer2_outputs(1549)) or (layer2_outputs(1128));
    layer3_outputs(1589) <= layer2_outputs(1865);
    layer3_outputs(1590) <= not(layer2_outputs(1924)) or (layer2_outputs(354));
    layer3_outputs(1591) <= (layer2_outputs(721)) and not (layer2_outputs(1159));
    layer3_outputs(1592) <= layer2_outputs(1941);
    layer3_outputs(1593) <= (layer2_outputs(411)) and (layer2_outputs(1971));
    layer3_outputs(1594) <= not(layer2_outputs(939)) or (layer2_outputs(143));
    layer3_outputs(1595) <= layer2_outputs(720);
    layer3_outputs(1596) <= not(layer2_outputs(485)) or (layer2_outputs(2510));
    layer3_outputs(1597) <= '1';
    layer3_outputs(1598) <= (layer2_outputs(1853)) and (layer2_outputs(760));
    layer3_outputs(1599) <= '1';
    layer3_outputs(1600) <= '0';
    layer3_outputs(1601) <= (layer2_outputs(1188)) and (layer2_outputs(1745));
    layer3_outputs(1602) <= not((layer2_outputs(1795)) or (layer2_outputs(2386)));
    layer3_outputs(1603) <= (layer2_outputs(1089)) and not (layer2_outputs(805));
    layer3_outputs(1604) <= not(layer2_outputs(2499));
    layer3_outputs(1605) <= (layer2_outputs(1676)) and not (layer2_outputs(348));
    layer3_outputs(1606) <= layer2_outputs(1047);
    layer3_outputs(1607) <= (layer2_outputs(2433)) and not (layer2_outputs(2259));
    layer3_outputs(1608) <= not(layer2_outputs(182));
    layer3_outputs(1609) <= layer2_outputs(951);
    layer3_outputs(1610) <= '0';
    layer3_outputs(1611) <= (layer2_outputs(1600)) and not (layer2_outputs(2151));
    layer3_outputs(1612) <= '0';
    layer3_outputs(1613) <= (layer2_outputs(156)) or (layer2_outputs(102));
    layer3_outputs(1614) <= (layer2_outputs(2071)) and not (layer2_outputs(516));
    layer3_outputs(1615) <= not(layer2_outputs(859));
    layer3_outputs(1616) <= not(layer2_outputs(1438));
    layer3_outputs(1617) <= not((layer2_outputs(1230)) or (layer2_outputs(75)));
    layer3_outputs(1618) <= not(layer2_outputs(950));
    layer3_outputs(1619) <= layer2_outputs(1154);
    layer3_outputs(1620) <= (layer2_outputs(232)) or (layer2_outputs(2128));
    layer3_outputs(1621) <= (layer2_outputs(2523)) or (layer2_outputs(1326));
    layer3_outputs(1622) <= not(layer2_outputs(2289));
    layer3_outputs(1623) <= (layer2_outputs(1166)) and not (layer2_outputs(1002));
    layer3_outputs(1624) <= not(layer2_outputs(1700)) or (layer2_outputs(932));
    layer3_outputs(1625) <= (layer2_outputs(1063)) and (layer2_outputs(1217));
    layer3_outputs(1626) <= not(layer2_outputs(764));
    layer3_outputs(1627) <= (layer2_outputs(2093)) and not (layer2_outputs(2192));
    layer3_outputs(1628) <= layer2_outputs(1709);
    layer3_outputs(1629) <= layer2_outputs(1578);
    layer3_outputs(1630) <= not((layer2_outputs(159)) and (layer2_outputs(790)));
    layer3_outputs(1631) <= layer2_outputs(2302);
    layer3_outputs(1632) <= '0';
    layer3_outputs(1633) <= not((layer2_outputs(1507)) and (layer2_outputs(430)));
    layer3_outputs(1634) <= not(layer2_outputs(251));
    layer3_outputs(1635) <= (layer2_outputs(126)) and (layer2_outputs(703));
    layer3_outputs(1636) <= layer2_outputs(1339);
    layer3_outputs(1637) <= (layer2_outputs(1910)) or (layer2_outputs(1758));
    layer3_outputs(1638) <= not(layer2_outputs(2094));
    layer3_outputs(1639) <= not(layer2_outputs(1972));
    layer3_outputs(1640) <= not(layer2_outputs(920)) or (layer2_outputs(906));
    layer3_outputs(1641) <= layer2_outputs(2015);
    layer3_outputs(1642) <= not(layer2_outputs(771));
    layer3_outputs(1643) <= not((layer2_outputs(795)) or (layer2_outputs(124)));
    layer3_outputs(1644) <= not(layer2_outputs(1960)) or (layer2_outputs(2042));
    layer3_outputs(1645) <= not(layer2_outputs(678)) or (layer2_outputs(907));
    layer3_outputs(1646) <= not(layer2_outputs(450));
    layer3_outputs(1647) <= not((layer2_outputs(1124)) or (layer2_outputs(652)));
    layer3_outputs(1648) <= (layer2_outputs(1808)) and not (layer2_outputs(133));
    layer3_outputs(1649) <= not(layer2_outputs(10));
    layer3_outputs(1650) <= layer2_outputs(1328);
    layer3_outputs(1651) <= (layer2_outputs(1752)) or (layer2_outputs(2039));
    layer3_outputs(1652) <= (layer2_outputs(1752)) or (layer2_outputs(337));
    layer3_outputs(1653) <= not(layer2_outputs(2149));
    layer3_outputs(1654) <= layer2_outputs(2504);
    layer3_outputs(1655) <= (layer2_outputs(523)) and not (layer2_outputs(1672));
    layer3_outputs(1656) <= '1';
    layer3_outputs(1657) <= '1';
    layer3_outputs(1658) <= not(layer2_outputs(781)) or (layer2_outputs(167));
    layer3_outputs(1659) <= layer2_outputs(1167);
    layer3_outputs(1660) <= not(layer2_outputs(2275)) or (layer2_outputs(739));
    layer3_outputs(1661) <= not(layer2_outputs(2451)) or (layer2_outputs(1698));
    layer3_outputs(1662) <= '0';
    layer3_outputs(1663) <= (layer2_outputs(1087)) and not (layer2_outputs(1874));
    layer3_outputs(1664) <= (layer2_outputs(914)) and (layer2_outputs(1241));
    layer3_outputs(1665) <= layer2_outputs(1423);
    layer3_outputs(1666) <= (layer2_outputs(1992)) or (layer2_outputs(1649));
    layer3_outputs(1667) <= not((layer2_outputs(1945)) and (layer2_outputs(225)));
    layer3_outputs(1668) <= not(layer2_outputs(959));
    layer3_outputs(1669) <= not(layer2_outputs(413)) or (layer2_outputs(541));
    layer3_outputs(1670) <= (layer2_outputs(1844)) and not (layer2_outputs(2279));
    layer3_outputs(1671) <= (layer2_outputs(348)) and not (layer2_outputs(1607));
    layer3_outputs(1672) <= not((layer2_outputs(2488)) and (layer2_outputs(1612)));
    layer3_outputs(1673) <= layer2_outputs(335);
    layer3_outputs(1674) <= not(layer2_outputs(1106));
    layer3_outputs(1675) <= (layer2_outputs(1105)) and (layer2_outputs(1552));
    layer3_outputs(1676) <= (layer2_outputs(2028)) or (layer2_outputs(208));
    layer3_outputs(1677) <= layer2_outputs(1194);
    layer3_outputs(1678) <= not(layer2_outputs(1291));
    layer3_outputs(1679) <= (layer2_outputs(1503)) or (layer2_outputs(1654));
    layer3_outputs(1680) <= (layer2_outputs(879)) and not (layer2_outputs(1309));
    layer3_outputs(1681) <= not(layer2_outputs(2134));
    layer3_outputs(1682) <= not((layer2_outputs(1870)) or (layer2_outputs(136)));
    layer3_outputs(1683) <= not(layer2_outputs(1264)) or (layer2_outputs(1413));
    layer3_outputs(1684) <= (layer2_outputs(2537)) and (layer2_outputs(2526));
    layer3_outputs(1685) <= not(layer2_outputs(389));
    layer3_outputs(1686) <= (layer2_outputs(1481)) and (layer2_outputs(374));
    layer3_outputs(1687) <= not(layer2_outputs(1577)) or (layer2_outputs(766));
    layer3_outputs(1688) <= not(layer2_outputs(1056));
    layer3_outputs(1689) <= layer2_outputs(428);
    layer3_outputs(1690) <= (layer2_outputs(1335)) or (layer2_outputs(663));
    layer3_outputs(1691) <= '0';
    layer3_outputs(1692) <= layer2_outputs(292);
    layer3_outputs(1693) <= layer2_outputs(854);
    layer3_outputs(1694) <= not(layer2_outputs(1657));
    layer3_outputs(1695) <= '0';
    layer3_outputs(1696) <= not((layer2_outputs(987)) or (layer2_outputs(1579)));
    layer3_outputs(1697) <= not(layer2_outputs(2106));
    layer3_outputs(1698) <= (layer2_outputs(2072)) and not (layer2_outputs(1502));
    layer3_outputs(1699) <= not(layer2_outputs(2285));
    layer3_outputs(1700) <= (layer2_outputs(1650)) or (layer2_outputs(386));
    layer3_outputs(1701) <= '1';
    layer3_outputs(1702) <= layer2_outputs(2190);
    layer3_outputs(1703) <= layer2_outputs(727);
    layer3_outputs(1704) <= not((layer2_outputs(1329)) or (layer2_outputs(1597)));
    layer3_outputs(1705) <= not(layer2_outputs(884));
    layer3_outputs(1706) <= '1';
    layer3_outputs(1707) <= not((layer2_outputs(1750)) and (layer2_outputs(745)));
    layer3_outputs(1708) <= not(layer2_outputs(2219)) or (layer2_outputs(1460));
    layer3_outputs(1709) <= layer2_outputs(2178);
    layer3_outputs(1710) <= '0';
    layer3_outputs(1711) <= (layer2_outputs(1816)) and not (layer2_outputs(660));
    layer3_outputs(1712) <= not(layer2_outputs(1362)) or (layer2_outputs(2283));
    layer3_outputs(1713) <= layer2_outputs(1736);
    layer3_outputs(1714) <= not(layer2_outputs(2324)) or (layer2_outputs(1427));
    layer3_outputs(1715) <= (layer2_outputs(272)) or (layer2_outputs(1319));
    layer3_outputs(1716) <= not(layer2_outputs(117)) or (layer2_outputs(1304));
    layer3_outputs(1717) <= '1';
    layer3_outputs(1718) <= not(layer2_outputs(2557));
    layer3_outputs(1719) <= not(layer2_outputs(689));
    layer3_outputs(1720) <= (layer2_outputs(2476)) or (layer2_outputs(1520));
    layer3_outputs(1721) <= not(layer2_outputs(513));
    layer3_outputs(1722) <= (layer2_outputs(1710)) and (layer2_outputs(293));
    layer3_outputs(1723) <= not((layer2_outputs(106)) and (layer2_outputs(459)));
    layer3_outputs(1724) <= not(layer2_outputs(2164));
    layer3_outputs(1725) <= not(layer2_outputs(132));
    layer3_outputs(1726) <= not(layer2_outputs(2361)) or (layer2_outputs(375));
    layer3_outputs(1727) <= (layer2_outputs(1960)) and not (layer2_outputs(2253));
    layer3_outputs(1728) <= not(layer2_outputs(1042));
    layer3_outputs(1729) <= not(layer2_outputs(1515));
    layer3_outputs(1730) <= (layer2_outputs(2389)) xor (layer2_outputs(194));
    layer3_outputs(1731) <= layer2_outputs(2349);
    layer3_outputs(1732) <= (layer2_outputs(2324)) and not (layer2_outputs(1301));
    layer3_outputs(1733) <= layer2_outputs(1251);
    layer3_outputs(1734) <= not(layer2_outputs(1378));
    layer3_outputs(1735) <= not(layer2_outputs(1191));
    layer3_outputs(1736) <= not((layer2_outputs(2550)) and (layer2_outputs(1112)));
    layer3_outputs(1737) <= not((layer2_outputs(2079)) and (layer2_outputs(161)));
    layer3_outputs(1738) <= not((layer2_outputs(1373)) or (layer2_outputs(306)));
    layer3_outputs(1739) <= not(layer2_outputs(1911));
    layer3_outputs(1740) <= not(layer2_outputs(2120));
    layer3_outputs(1741) <= not(layer2_outputs(915)) or (layer2_outputs(2293));
    layer3_outputs(1742) <= not(layer2_outputs(615));
    layer3_outputs(1743) <= (layer2_outputs(1473)) or (layer2_outputs(1626));
    layer3_outputs(1744) <= not(layer2_outputs(509));
    layer3_outputs(1745) <= layer2_outputs(2334);
    layer3_outputs(1746) <= not(layer2_outputs(2531));
    layer3_outputs(1747) <= not(layer2_outputs(360));
    layer3_outputs(1748) <= '0';
    layer3_outputs(1749) <= (layer2_outputs(2244)) and not (layer2_outputs(60));
    layer3_outputs(1750) <= (layer2_outputs(584)) and not (layer2_outputs(129));
    layer3_outputs(1751) <= (layer2_outputs(1641)) and not (layer2_outputs(2327));
    layer3_outputs(1752) <= (layer2_outputs(1734)) or (layer2_outputs(18));
    layer3_outputs(1753) <= layer2_outputs(498);
    layer3_outputs(1754) <= not((layer2_outputs(2261)) and (layer2_outputs(1050)));
    layer3_outputs(1755) <= not(layer2_outputs(2364)) or (layer2_outputs(1285));
    layer3_outputs(1756) <= layer2_outputs(2410);
    layer3_outputs(1757) <= not((layer2_outputs(339)) and (layer2_outputs(165)));
    layer3_outputs(1758) <= not((layer2_outputs(416)) or (layer2_outputs(487)));
    layer3_outputs(1759) <= not(layer2_outputs(1568));
    layer3_outputs(1760) <= (layer2_outputs(1807)) and (layer2_outputs(1829));
    layer3_outputs(1761) <= '1';
    layer3_outputs(1762) <= '1';
    layer3_outputs(1763) <= '0';
    layer3_outputs(1764) <= layer2_outputs(1450);
    layer3_outputs(1765) <= not(layer2_outputs(2231));
    layer3_outputs(1766) <= not(layer2_outputs(2414));
    layer3_outputs(1767) <= not(layer2_outputs(1572)) or (layer2_outputs(2157));
    layer3_outputs(1768) <= not(layer2_outputs(2282));
    layer3_outputs(1769) <= (layer2_outputs(1838)) and (layer2_outputs(1271));
    layer3_outputs(1770) <= layer2_outputs(590);
    layer3_outputs(1771) <= (layer2_outputs(2088)) and (layer2_outputs(2544));
    layer3_outputs(1772) <= layer2_outputs(1506);
    layer3_outputs(1773) <= not(layer2_outputs(1067)) or (layer2_outputs(1800));
    layer3_outputs(1774) <= layer2_outputs(732);
    layer3_outputs(1775) <= '0';
    layer3_outputs(1776) <= layer2_outputs(806);
    layer3_outputs(1777) <= not(layer2_outputs(1174));
    layer3_outputs(1778) <= layer2_outputs(2091);
    layer3_outputs(1779) <= (layer2_outputs(674)) and not (layer2_outputs(1673));
    layer3_outputs(1780) <= not((layer2_outputs(298)) and (layer2_outputs(841)));
    layer3_outputs(1781) <= layer2_outputs(1399);
    layer3_outputs(1782) <= not(layer2_outputs(1836)) or (layer2_outputs(1880));
    layer3_outputs(1783) <= (layer2_outputs(2524)) and (layer2_outputs(31));
    layer3_outputs(1784) <= (layer2_outputs(1704)) and not (layer2_outputs(527));
    layer3_outputs(1785) <= not(layer2_outputs(2336)) or (layer2_outputs(1248));
    layer3_outputs(1786) <= layer2_outputs(1176);
    layer3_outputs(1787) <= (layer2_outputs(1182)) and not (layer2_outputs(538));
    layer3_outputs(1788) <= '0';
    layer3_outputs(1789) <= layer2_outputs(138);
    layer3_outputs(1790) <= not(layer2_outputs(1629));
    layer3_outputs(1791) <= not(layer2_outputs(1913));
    layer3_outputs(1792) <= (layer2_outputs(317)) or (layer2_outputs(622));
    layer3_outputs(1793) <= (layer2_outputs(1351)) and not (layer2_outputs(1604));
    layer3_outputs(1794) <= layer2_outputs(1554);
    layer3_outputs(1795) <= not(layer2_outputs(2379));
    layer3_outputs(1796) <= (layer2_outputs(1883)) and not (layer2_outputs(940));
    layer3_outputs(1797) <= not(layer2_outputs(2074)) or (layer2_outputs(2));
    layer3_outputs(1798) <= '0';
    layer3_outputs(1799) <= not(layer2_outputs(1426)) or (layer2_outputs(1070));
    layer3_outputs(1800) <= (layer2_outputs(1204)) and not (layer2_outputs(1088));
    layer3_outputs(1801) <= (layer2_outputs(2347)) or (layer2_outputs(1293));
    layer3_outputs(1802) <= layer2_outputs(1801);
    layer3_outputs(1803) <= '0';
    layer3_outputs(1804) <= (layer2_outputs(1015)) and not (layer2_outputs(542));
    layer3_outputs(1805) <= not((layer2_outputs(902)) or (layer2_outputs(45)));
    layer3_outputs(1806) <= not(layer2_outputs(2231)) or (layer2_outputs(1742));
    layer3_outputs(1807) <= (layer2_outputs(152)) and not (layer2_outputs(2302));
    layer3_outputs(1808) <= not((layer2_outputs(2325)) or (layer2_outputs(739)));
    layer3_outputs(1809) <= not(layer2_outputs(1786));
    layer3_outputs(1810) <= '1';
    layer3_outputs(1811) <= not(layer2_outputs(84)) or (layer2_outputs(2559));
    layer3_outputs(1812) <= layer2_outputs(2434);
    layer3_outputs(1813) <= not(layer2_outputs(834));
    layer3_outputs(1814) <= (layer2_outputs(1398)) or (layer2_outputs(2343));
    layer3_outputs(1815) <= layer2_outputs(1713);
    layer3_outputs(1816) <= layer2_outputs(2015);
    layer3_outputs(1817) <= (layer2_outputs(1579)) and not (layer2_outputs(1898));
    layer3_outputs(1818) <= '1';
    layer3_outputs(1819) <= not(layer2_outputs(130));
    layer3_outputs(1820) <= (layer2_outputs(2453)) and (layer2_outputs(1130));
    layer3_outputs(1821) <= layer2_outputs(1126);
    layer3_outputs(1822) <= not(layer2_outputs(1302));
    layer3_outputs(1823) <= (layer2_outputs(258)) and not (layer2_outputs(163));
    layer3_outputs(1824) <= not((layer2_outputs(1428)) and (layer2_outputs(43)));
    layer3_outputs(1825) <= (layer2_outputs(1914)) and (layer2_outputs(1770));
    layer3_outputs(1826) <= not((layer2_outputs(559)) xor (layer2_outputs(222)));
    layer3_outputs(1827) <= '0';
    layer3_outputs(1828) <= not(layer2_outputs(44));
    layer3_outputs(1829) <= not(layer2_outputs(503));
    layer3_outputs(1830) <= layer2_outputs(1241);
    layer3_outputs(1831) <= not(layer2_outputs(2204));
    layer3_outputs(1832) <= layer2_outputs(2201);
    layer3_outputs(1833) <= not(layer2_outputs(1072));
    layer3_outputs(1834) <= (layer2_outputs(1488)) or (layer2_outputs(826));
    layer3_outputs(1835) <= not((layer2_outputs(828)) and (layer2_outputs(1232)));
    layer3_outputs(1836) <= layer2_outputs(406);
    layer3_outputs(1837) <= (layer2_outputs(2174)) or (layer2_outputs(1980));
    layer3_outputs(1838) <= (layer2_outputs(1676)) or (layer2_outputs(708));
    layer3_outputs(1839) <= not(layer2_outputs(1782)) or (layer2_outputs(551));
    layer3_outputs(1840) <= layer2_outputs(814);
    layer3_outputs(1841) <= not(layer2_outputs(328));
    layer3_outputs(1842) <= layer2_outputs(1426);
    layer3_outputs(1843) <= layer2_outputs(567);
    layer3_outputs(1844) <= not(layer2_outputs(2429)) or (layer2_outputs(910));
    layer3_outputs(1845) <= '1';
    layer3_outputs(1846) <= not(layer2_outputs(488));
    layer3_outputs(1847) <= not(layer2_outputs(141));
    layer3_outputs(1848) <= layer2_outputs(1080);
    layer3_outputs(1849) <= layer2_outputs(536);
    layer3_outputs(1850) <= (layer2_outputs(1401)) and (layer2_outputs(955));
    layer3_outputs(1851) <= layer2_outputs(804);
    layer3_outputs(1852) <= not(layer2_outputs(190)) or (layer2_outputs(213));
    layer3_outputs(1853) <= (layer2_outputs(1163)) and not (layer2_outputs(1556));
    layer3_outputs(1854) <= (layer2_outputs(111)) or (layer2_outputs(479));
    layer3_outputs(1855) <= (layer2_outputs(1978)) xor (layer2_outputs(972));
    layer3_outputs(1856) <= '1';
    layer3_outputs(1857) <= not(layer2_outputs(627));
    layer3_outputs(1858) <= '0';
    layer3_outputs(1859) <= not((layer2_outputs(1629)) or (layer2_outputs(1542)));
    layer3_outputs(1860) <= layer2_outputs(840);
    layer3_outputs(1861) <= not(layer2_outputs(2075)) or (layer2_outputs(1630));
    layer3_outputs(1862) <= not(layer2_outputs(1770)) or (layer2_outputs(1731));
    layer3_outputs(1863) <= '0';
    layer3_outputs(1864) <= not((layer2_outputs(2256)) or (layer2_outputs(1153)));
    layer3_outputs(1865) <= not(layer2_outputs(49));
    layer3_outputs(1866) <= layer2_outputs(2520);
    layer3_outputs(1867) <= (layer2_outputs(1223)) and (layer2_outputs(2212));
    layer3_outputs(1868) <= (layer2_outputs(1199)) and not (layer2_outputs(2262));
    layer3_outputs(1869) <= (layer2_outputs(955)) and (layer2_outputs(473));
    layer3_outputs(1870) <= not((layer2_outputs(1877)) xor (layer2_outputs(1421)));
    layer3_outputs(1871) <= not(layer2_outputs(2159));
    layer3_outputs(1872) <= layer2_outputs(1987);
    layer3_outputs(1873) <= '0';
    layer3_outputs(1874) <= '1';
    layer3_outputs(1875) <= not(layer2_outputs(2131));
    layer3_outputs(1876) <= not(layer2_outputs(899));
    layer3_outputs(1877) <= not((layer2_outputs(2135)) or (layer2_outputs(393)));
    layer3_outputs(1878) <= not(layer2_outputs(1338));
    layer3_outputs(1879) <= (layer2_outputs(1160)) and not (layer2_outputs(2312));
    layer3_outputs(1880) <= not(layer2_outputs(1105)) or (layer2_outputs(1509));
    layer3_outputs(1881) <= not((layer2_outputs(2135)) or (layer2_outputs(315)));
    layer3_outputs(1882) <= layer2_outputs(959);
    layer3_outputs(1883) <= '0';
    layer3_outputs(1884) <= (layer2_outputs(2279)) and (layer2_outputs(443));
    layer3_outputs(1885) <= not(layer2_outputs(1617)) or (layer2_outputs(2355));
    layer3_outputs(1886) <= not((layer2_outputs(139)) or (layer2_outputs(2077)));
    layer3_outputs(1887) <= layer2_outputs(1664);
    layer3_outputs(1888) <= not(layer2_outputs(1899)) or (layer2_outputs(2322));
    layer3_outputs(1889) <= layer2_outputs(1557);
    layer3_outputs(1890) <= not((layer2_outputs(1209)) and (layer2_outputs(1993)));
    layer3_outputs(1891) <= (layer2_outputs(218)) or (layer2_outputs(1419));
    layer3_outputs(1892) <= (layer2_outputs(1593)) and (layer2_outputs(1179));
    layer3_outputs(1893) <= layer2_outputs(439);
    layer3_outputs(1894) <= not(layer2_outputs(1909)) or (layer2_outputs(2464));
    layer3_outputs(1895) <= not(layer2_outputs(1006)) or (layer2_outputs(805));
    layer3_outputs(1896) <= layer2_outputs(2232);
    layer3_outputs(1897) <= not(layer2_outputs(1292));
    layer3_outputs(1898) <= (layer2_outputs(726)) and (layer2_outputs(853));
    layer3_outputs(1899) <= layer2_outputs(2297);
    layer3_outputs(1900) <= not(layer2_outputs(2484));
    layer3_outputs(1901) <= not(layer2_outputs(96)) or (layer2_outputs(1005));
    layer3_outputs(1902) <= (layer2_outputs(822)) and not (layer2_outputs(30));
    layer3_outputs(1903) <= not(layer2_outputs(776));
    layer3_outputs(1904) <= not(layer2_outputs(2307)) or (layer2_outputs(2301));
    layer3_outputs(1905) <= (layer2_outputs(2382)) or (layer2_outputs(1647));
    layer3_outputs(1906) <= (layer2_outputs(430)) and (layer2_outputs(204));
    layer3_outputs(1907) <= '1';
    layer3_outputs(1908) <= not(layer2_outputs(729));
    layer3_outputs(1909) <= layer2_outputs(1600);
    layer3_outputs(1910) <= layer2_outputs(347);
    layer3_outputs(1911) <= (layer2_outputs(483)) and (layer2_outputs(1066));
    layer3_outputs(1912) <= (layer2_outputs(709)) and not (layer2_outputs(419));
    layer3_outputs(1913) <= '0';
    layer3_outputs(1914) <= not(layer2_outputs(535)) or (layer2_outputs(621));
    layer3_outputs(1915) <= (layer2_outputs(1705)) or (layer2_outputs(706));
    layer3_outputs(1916) <= layer2_outputs(1677);
    layer3_outputs(1917) <= layer2_outputs(1372);
    layer3_outputs(1918) <= '0';
    layer3_outputs(1919) <= layer2_outputs(519);
    layer3_outputs(1920) <= '0';
    layer3_outputs(1921) <= '1';
    layer3_outputs(1922) <= not((layer2_outputs(778)) and (layer2_outputs(2074)));
    layer3_outputs(1923) <= layer2_outputs(786);
    layer3_outputs(1924) <= (layer2_outputs(1570)) and not (layer2_outputs(1084));
    layer3_outputs(1925) <= '0';
    layer3_outputs(1926) <= layer2_outputs(143);
    layer3_outputs(1927) <= layer2_outputs(262);
    layer3_outputs(1928) <= layer2_outputs(1944);
    layer3_outputs(1929) <= layer2_outputs(1477);
    layer3_outputs(1930) <= layer2_outputs(2366);
    layer3_outputs(1931) <= layer2_outputs(217);
    layer3_outputs(1932) <= '1';
    layer3_outputs(1933) <= not(layer2_outputs(1921)) or (layer2_outputs(1000));
    layer3_outputs(1934) <= (layer2_outputs(1776)) and not (layer2_outputs(975));
    layer3_outputs(1935) <= (layer2_outputs(436)) and not (layer2_outputs(621));
    layer3_outputs(1936) <= (layer2_outputs(1100)) and (layer2_outputs(2073));
    layer3_outputs(1937) <= (layer2_outputs(2409)) and (layer2_outputs(1959));
    layer3_outputs(1938) <= not(layer2_outputs(1012));
    layer3_outputs(1939) <= not(layer2_outputs(1310));
    layer3_outputs(1940) <= not(layer2_outputs(1881)) or (layer2_outputs(2535));
    layer3_outputs(1941) <= not(layer2_outputs(761));
    layer3_outputs(1942) <= not(layer2_outputs(2388));
    layer3_outputs(1943) <= layer2_outputs(1932);
    layer3_outputs(1944) <= layer2_outputs(566);
    layer3_outputs(1945) <= (layer2_outputs(1200)) and (layer2_outputs(684));
    layer3_outputs(1946) <= not(layer2_outputs(1919));
    layer3_outputs(1947) <= not((layer2_outputs(1744)) and (layer2_outputs(331)));
    layer3_outputs(1948) <= (layer2_outputs(2528)) and not (layer2_outputs(939));
    layer3_outputs(1949) <= layer2_outputs(400);
    layer3_outputs(1950) <= (layer2_outputs(456)) and not (layer2_outputs(1761));
    layer3_outputs(1951) <= (layer2_outputs(1797)) and (layer2_outputs(120));
    layer3_outputs(1952) <= layer2_outputs(2518);
    layer3_outputs(1953) <= layer2_outputs(1453);
    layer3_outputs(1954) <= not(layer2_outputs(2453));
    layer3_outputs(1955) <= '1';
    layer3_outputs(1956) <= not((layer2_outputs(518)) xor (layer2_outputs(658)));
    layer3_outputs(1957) <= '1';
    layer3_outputs(1958) <= '0';
    layer3_outputs(1959) <= (layer2_outputs(1324)) and not (layer2_outputs(1122));
    layer3_outputs(1960) <= '0';
    layer3_outputs(1961) <= not((layer2_outputs(712)) and (layer2_outputs(219)));
    layer3_outputs(1962) <= not((layer2_outputs(2215)) or (layer2_outputs(1054)));
    layer3_outputs(1963) <= (layer2_outputs(2273)) and not (layer2_outputs(937));
    layer3_outputs(1964) <= not(layer2_outputs(2257)) or (layer2_outputs(56));
    layer3_outputs(1965) <= '0';
    layer3_outputs(1966) <= not((layer2_outputs(2054)) or (layer2_outputs(1638)));
    layer3_outputs(1967) <= not(layer2_outputs(1003));
    layer3_outputs(1968) <= (layer2_outputs(528)) and not (layer2_outputs(1334));
    layer3_outputs(1969) <= '0';
    layer3_outputs(1970) <= layer2_outputs(1577);
    layer3_outputs(1971) <= '1';
    layer3_outputs(1972) <= layer2_outputs(637);
    layer3_outputs(1973) <= (layer2_outputs(1374)) or (layer2_outputs(800));
    layer3_outputs(1974) <= not(layer2_outputs(1073)) or (layer2_outputs(598));
    layer3_outputs(1975) <= '0';
    layer3_outputs(1976) <= layer2_outputs(2255);
    layer3_outputs(1977) <= not((layer2_outputs(2085)) or (layer2_outputs(1382)));
    layer3_outputs(1978) <= not(layer2_outputs(2049));
    layer3_outputs(1979) <= layer2_outputs(389);
    layer3_outputs(1980) <= not((layer2_outputs(184)) and (layer2_outputs(21)));
    layer3_outputs(1981) <= not((layer2_outputs(2533)) and (layer2_outputs(1858)));
    layer3_outputs(1982) <= layer2_outputs(2351);
    layer3_outputs(1983) <= not(layer2_outputs(784));
    layer3_outputs(1984) <= '0';
    layer3_outputs(1985) <= not((layer2_outputs(1181)) or (layer2_outputs(758)));
    layer3_outputs(1986) <= (layer2_outputs(357)) and not (layer2_outputs(191));
    layer3_outputs(1987) <= '1';
    layer3_outputs(1988) <= not(layer2_outputs(79));
    layer3_outputs(1989) <= layer2_outputs(1557);
    layer3_outputs(1990) <= not(layer2_outputs(1456));
    layer3_outputs(1991) <= not((layer2_outputs(1402)) or (layer2_outputs(1131)));
    layer3_outputs(1992) <= not((layer2_outputs(2098)) or (layer2_outputs(741)));
    layer3_outputs(1993) <= not(layer2_outputs(484));
    layer3_outputs(1994) <= not(layer2_outputs(2450)) or (layer2_outputs(883));
    layer3_outputs(1995) <= not(layer2_outputs(894)) or (layer2_outputs(1484));
    layer3_outputs(1996) <= '1';
    layer3_outputs(1997) <= layer2_outputs(2195);
    layer3_outputs(1998) <= layer2_outputs(1860);
    layer3_outputs(1999) <= (layer2_outputs(503)) or (layer2_outputs(2298));
    layer3_outputs(2000) <= layer2_outputs(733);
    layer3_outputs(2001) <= not((layer2_outputs(1812)) or (layer2_outputs(1448)));
    layer3_outputs(2002) <= not(layer2_outputs(346));
    layer3_outputs(2003) <= '1';
    layer3_outputs(2004) <= '0';
    layer3_outputs(2005) <= (layer2_outputs(1107)) or (layer2_outputs(17));
    layer3_outputs(2006) <= not(layer2_outputs(109));
    layer3_outputs(2007) <= not((layer2_outputs(87)) and (layer2_outputs(2354)));
    layer3_outputs(2008) <= not(layer2_outputs(1659)) or (layer2_outputs(2454));
    layer3_outputs(2009) <= not((layer2_outputs(918)) or (layer2_outputs(2017)));
    layer3_outputs(2010) <= (layer2_outputs(1442)) and (layer2_outputs(114));
    layer3_outputs(2011) <= not(layer2_outputs(2539)) or (layer2_outputs(2305));
    layer3_outputs(2012) <= (layer2_outputs(340)) and not (layer2_outputs(5));
    layer3_outputs(2013) <= layer2_outputs(134);
    layer3_outputs(2014) <= (layer2_outputs(506)) and (layer2_outputs(2320));
    layer3_outputs(2015) <= layer2_outputs(2397);
    layer3_outputs(2016) <= not(layer2_outputs(1650));
    layer3_outputs(2017) <= (layer2_outputs(1321)) and not (layer2_outputs(2247));
    layer3_outputs(2018) <= (layer2_outputs(48)) and not (layer2_outputs(1196));
    layer3_outputs(2019) <= (layer2_outputs(2418)) and not (layer2_outputs(907));
    layer3_outputs(2020) <= not(layer2_outputs(2163));
    layer3_outputs(2021) <= layer2_outputs(852);
    layer3_outputs(2022) <= (layer2_outputs(1531)) and not (layer2_outputs(597));
    layer3_outputs(2023) <= not(layer2_outputs(1565)) or (layer2_outputs(415));
    layer3_outputs(2024) <= layer2_outputs(1326);
    layer3_outputs(2025) <= layer2_outputs(724);
    layer3_outputs(2026) <= (layer2_outputs(2526)) and not (layer2_outputs(1455));
    layer3_outputs(2027) <= not(layer2_outputs(1817));
    layer3_outputs(2028) <= not(layer2_outputs(2422)) or (layer2_outputs(860));
    layer3_outputs(2029) <= not(layer2_outputs(308));
    layer3_outputs(2030) <= layer2_outputs(2238);
    layer3_outputs(2031) <= not(layer2_outputs(536)) or (layer2_outputs(1634));
    layer3_outputs(2032) <= not(layer2_outputs(312));
    layer3_outputs(2033) <= (layer2_outputs(552)) or (layer2_outputs(1791));
    layer3_outputs(2034) <= not(layer2_outputs(1043)) or (layer2_outputs(1210));
    layer3_outputs(2035) <= not(layer2_outputs(573));
    layer3_outputs(2036) <= (layer2_outputs(1249)) and (layer2_outputs(2091));
    layer3_outputs(2037) <= not(layer2_outputs(301));
    layer3_outputs(2038) <= (layer2_outputs(2509)) and not (layer2_outputs(211));
    layer3_outputs(2039) <= '0';
    layer3_outputs(2040) <= (layer2_outputs(52)) and (layer2_outputs(825));
    layer3_outputs(2041) <= not(layer2_outputs(2133)) or (layer2_outputs(118));
    layer3_outputs(2042) <= not(layer2_outputs(2293));
    layer3_outputs(2043) <= not((layer2_outputs(1344)) or (layer2_outputs(1184)));
    layer3_outputs(2044) <= (layer2_outputs(421)) or (layer2_outputs(639));
    layer3_outputs(2045) <= (layer2_outputs(1857)) and not (layer2_outputs(2155));
    layer3_outputs(2046) <= (layer2_outputs(1030)) and not (layer2_outputs(1403));
    layer3_outputs(2047) <= (layer2_outputs(645)) or (layer2_outputs(479));
    layer3_outputs(2048) <= not(layer2_outputs(659));
    layer3_outputs(2049) <= not(layer2_outputs(1309));
    layer3_outputs(2050) <= layer2_outputs(577);
    layer3_outputs(2051) <= not(layer2_outputs(1492)) or (layer2_outputs(1826));
    layer3_outputs(2052) <= layer2_outputs(1510);
    layer3_outputs(2053) <= '1';
    layer3_outputs(2054) <= not(layer2_outputs(743)) or (layer2_outputs(1072));
    layer3_outputs(2055) <= layer2_outputs(1343);
    layer3_outputs(2056) <= not(layer2_outputs(2398));
    layer3_outputs(2057) <= '0';
    layer3_outputs(2058) <= not(layer2_outputs(492));
    layer3_outputs(2059) <= not(layer2_outputs(1035)) or (layer2_outputs(685));
    layer3_outputs(2060) <= '1';
    layer3_outputs(2061) <= layer2_outputs(1867);
    layer3_outputs(2062) <= not(layer2_outputs(1984));
    layer3_outputs(2063) <= not(layer2_outputs(1222)) or (layer2_outputs(1367));
    layer3_outputs(2064) <= not(layer2_outputs(428)) or (layer2_outputs(2141));
    layer3_outputs(2065) <= (layer2_outputs(1820)) or (layer2_outputs(1866));
    layer3_outputs(2066) <= (layer2_outputs(1583)) or (layer2_outputs(361));
    layer3_outputs(2067) <= (layer2_outputs(800)) and not (layer2_outputs(1839));
    layer3_outputs(2068) <= (layer2_outputs(2308)) or (layer2_outputs(718));
    layer3_outputs(2069) <= (layer2_outputs(1787)) and not (layer2_outputs(1768));
    layer3_outputs(2070) <= not(layer2_outputs(174));
    layer3_outputs(2071) <= layer2_outputs(1131);
    layer3_outputs(2072) <= (layer2_outputs(778)) xor (layer2_outputs(2111));
    layer3_outputs(2073) <= '0';
    layer3_outputs(2074) <= not(layer2_outputs(70)) or (layer2_outputs(644));
    layer3_outputs(2075) <= not(layer2_outputs(842));
    layer3_outputs(2076) <= '1';
    layer3_outputs(2077) <= not((layer2_outputs(1977)) and (layer2_outputs(2088)));
    layer3_outputs(2078) <= not(layer2_outputs(2305));
    layer3_outputs(2079) <= (layer2_outputs(52)) or (layer2_outputs(83));
    layer3_outputs(2080) <= (layer2_outputs(2333)) xor (layer2_outputs(3));
    layer3_outputs(2081) <= (layer2_outputs(373)) and (layer2_outputs(2505));
    layer3_outputs(2082) <= (layer2_outputs(2340)) and not (layer2_outputs(1049));
    layer3_outputs(2083) <= layer2_outputs(1031);
    layer3_outputs(2084) <= layer2_outputs(600);
    layer3_outputs(2085) <= (layer2_outputs(478)) or (layer2_outputs(1857));
    layer3_outputs(2086) <= layer2_outputs(2229);
    layer3_outputs(2087) <= '1';
    layer3_outputs(2088) <= (layer2_outputs(1320)) and not (layer2_outputs(1278));
    layer3_outputs(2089) <= layer2_outputs(1396);
    layer3_outputs(2090) <= not(layer2_outputs(1915)) or (layer2_outputs(937));
    layer3_outputs(2091) <= layer2_outputs(157);
    layer3_outputs(2092) <= (layer2_outputs(728)) and (layer2_outputs(2398));
    layer3_outputs(2093) <= layer2_outputs(191);
    layer3_outputs(2094) <= (layer2_outputs(279)) and not (layer2_outputs(1528));
    layer3_outputs(2095) <= not(layer2_outputs(1696));
    layer3_outputs(2096) <= not(layer2_outputs(1311));
    layer3_outputs(2097) <= not((layer2_outputs(1651)) and (layer2_outputs(565)));
    layer3_outputs(2098) <= not(layer2_outputs(2346));
    layer3_outputs(2099) <= not((layer2_outputs(1337)) and (layer2_outputs(2425)));
    layer3_outputs(2100) <= (layer2_outputs(2265)) and not (layer2_outputs(753));
    layer3_outputs(2101) <= layer2_outputs(646);
    layer3_outputs(2102) <= (layer2_outputs(656)) or (layer2_outputs(1240));
    layer3_outputs(2103) <= '1';
    layer3_outputs(2104) <= not(layer2_outputs(2499)) or (layer2_outputs(487));
    layer3_outputs(2105) <= (layer2_outputs(770)) or (layer2_outputs(2346));
    layer3_outputs(2106) <= not((layer2_outputs(1485)) or (layer2_outputs(285)));
    layer3_outputs(2107) <= layer2_outputs(2529);
    layer3_outputs(2108) <= layer2_outputs(5);
    layer3_outputs(2109) <= (layer2_outputs(1436)) or (layer2_outputs(2124));
    layer3_outputs(2110) <= not(layer2_outputs(2149));
    layer3_outputs(2111) <= not(layer2_outputs(1836));
    layer3_outputs(2112) <= (layer2_outputs(842)) and (layer2_outputs(1536));
    layer3_outputs(2113) <= not(layer2_outputs(1873));
    layer3_outputs(2114) <= not(layer2_outputs(1424));
    layer3_outputs(2115) <= not(layer2_outputs(382));
    layer3_outputs(2116) <= (layer2_outputs(1254)) and not (layer2_outputs(2169));
    layer3_outputs(2117) <= layer2_outputs(1425);
    layer3_outputs(2118) <= not((layer2_outputs(2057)) and (layer2_outputs(594)));
    layer3_outputs(2119) <= (layer2_outputs(2222)) and not (layer2_outputs(1180));
    layer3_outputs(2120) <= layer2_outputs(963);
    layer3_outputs(2121) <= layer2_outputs(1275);
    layer3_outputs(2122) <= (layer2_outputs(475)) and (layer2_outputs(1616));
    layer3_outputs(2123) <= layer2_outputs(744);
    layer3_outputs(2124) <= not(layer2_outputs(1533));
    layer3_outputs(2125) <= (layer2_outputs(1278)) and not (layer2_outputs(581));
    layer3_outputs(2126) <= not(layer2_outputs(116));
    layer3_outputs(2127) <= not(layer2_outputs(2347));
    layer3_outputs(2128) <= '1';
    layer3_outputs(2129) <= layer2_outputs(1034);
    layer3_outputs(2130) <= not((layer2_outputs(1471)) or (layer2_outputs(1361)));
    layer3_outputs(2131) <= (layer2_outputs(2245)) and not (layer2_outputs(227));
    layer3_outputs(2132) <= (layer2_outputs(641)) or (layer2_outputs(540));
    layer3_outputs(2133) <= not(layer2_outputs(2079)) or (layer2_outputs(971));
    layer3_outputs(2134) <= not((layer2_outputs(1666)) or (layer2_outputs(2516)));
    layer3_outputs(2135) <= layer2_outputs(365);
    layer3_outputs(2136) <= '1';
    layer3_outputs(2137) <= not((layer2_outputs(1655)) or (layer2_outputs(1560)));
    layer3_outputs(2138) <= layer2_outputs(2046);
    layer3_outputs(2139) <= layer2_outputs(85);
    layer3_outputs(2140) <= (layer2_outputs(2274)) and not (layer2_outputs(1790));
    layer3_outputs(2141) <= (layer2_outputs(1451)) and (layer2_outputs(1628));
    layer3_outputs(2142) <= not(layer2_outputs(2431));
    layer3_outputs(2143) <= not(layer2_outputs(1516));
    layer3_outputs(2144) <= (layer2_outputs(1417)) and (layer2_outputs(372));
    layer3_outputs(2145) <= (layer2_outputs(502)) and not (layer2_outputs(1231));
    layer3_outputs(2146) <= not((layer2_outputs(2481)) or (layer2_outputs(660)));
    layer3_outputs(2147) <= layer2_outputs(22);
    layer3_outputs(2148) <= not(layer2_outputs(1568));
    layer3_outputs(2149) <= not(layer2_outputs(1589));
    layer3_outputs(2150) <= not(layer2_outputs(1957));
    layer3_outputs(2151) <= not(layer2_outputs(654));
    layer3_outputs(2152) <= not((layer2_outputs(445)) and (layer2_outputs(180)));
    layer3_outputs(2153) <= not((layer2_outputs(456)) or (layer2_outputs(1702)));
    layer3_outputs(2154) <= layer2_outputs(1768);
    layer3_outputs(2155) <= not((layer2_outputs(1967)) and (layer2_outputs(1447)));
    layer3_outputs(2156) <= not(layer2_outputs(1039));
    layer3_outputs(2157) <= not(layer2_outputs(104)) or (layer2_outputs(668));
    layer3_outputs(2158) <= not(layer2_outputs(100));
    layer3_outputs(2159) <= not(layer2_outputs(763));
    layer3_outputs(2160) <= layer2_outputs(848);
    layer3_outputs(2161) <= not(layer2_outputs(1806));
    layer3_outputs(2162) <= not(layer2_outputs(493));
    layer3_outputs(2163) <= (layer2_outputs(120)) and (layer2_outputs(605));
    layer3_outputs(2164) <= (layer2_outputs(384)) or (layer2_outputs(1970));
    layer3_outputs(2165) <= not((layer2_outputs(1287)) and (layer2_outputs(1800)));
    layer3_outputs(2166) <= '0';
    layer3_outputs(2167) <= not(layer2_outputs(2108));
    layer3_outputs(2168) <= (layer2_outputs(1686)) and not (layer2_outputs(198));
    layer3_outputs(2169) <= '1';
    layer3_outputs(2170) <= layer2_outputs(748);
    layer3_outputs(2171) <= '0';
    layer3_outputs(2172) <= not((layer2_outputs(2521)) and (layer2_outputs(1417)));
    layer3_outputs(2173) <= (layer2_outputs(564)) and not (layer2_outputs(895));
    layer3_outputs(2174) <= not(layer2_outputs(1716));
    layer3_outputs(2175) <= (layer2_outputs(438)) and not (layer2_outputs(1864));
    layer3_outputs(2176) <= '1';
    layer3_outputs(2177) <= not(layer2_outputs(1837)) or (layer2_outputs(774));
    layer3_outputs(2178) <= '0';
    layer3_outputs(2179) <= (layer2_outputs(318)) and not (layer2_outputs(1980));
    layer3_outputs(2180) <= not((layer2_outputs(1804)) and (layer2_outputs(868)));
    layer3_outputs(2181) <= not((layer2_outputs(580)) or (layer2_outputs(1976)));
    layer3_outputs(2182) <= not(layer2_outputs(874));
    layer3_outputs(2183) <= (layer2_outputs(2129)) and not (layer2_outputs(557));
    layer3_outputs(2184) <= not(layer2_outputs(2236)) or (layer2_outputs(881));
    layer3_outputs(2185) <= not((layer2_outputs(284)) and (layer2_outputs(919)));
    layer3_outputs(2186) <= (layer2_outputs(1462)) xor (layer2_outputs(1522));
    layer3_outputs(2187) <= not((layer2_outputs(833)) and (layer2_outputs(1486)));
    layer3_outputs(2188) <= layer2_outputs(1625);
    layer3_outputs(2189) <= not(layer2_outputs(477));
    layer3_outputs(2190) <= not(layer2_outputs(1795));
    layer3_outputs(2191) <= '1';
    layer3_outputs(2192) <= (layer2_outputs(946)) and (layer2_outputs(1974));
    layer3_outputs(2193) <= layer2_outputs(359);
    layer3_outputs(2194) <= (layer2_outputs(1157)) and (layer2_outputs(2144));
    layer3_outputs(2195) <= (layer2_outputs(455)) and not (layer2_outputs(174));
    layer3_outputs(2196) <= not(layer2_outputs(759));
    layer3_outputs(2197) <= not(layer2_outputs(2474));
    layer3_outputs(2198) <= '1';
    layer3_outputs(2199) <= not((layer2_outputs(2528)) and (layer2_outputs(99)));
    layer3_outputs(2200) <= (layer2_outputs(2224)) xor (layer2_outputs(2385));
    layer3_outputs(2201) <= not(layer2_outputs(2543)) or (layer2_outputs(295));
    layer3_outputs(2202) <= layer2_outputs(2412);
    layer3_outputs(2203) <= not((layer2_outputs(1567)) or (layer2_outputs(2304)));
    layer3_outputs(2204) <= '0';
    layer3_outputs(2205) <= (layer2_outputs(1336)) and (layer2_outputs(1047));
    layer3_outputs(2206) <= not((layer2_outputs(2013)) or (layer2_outputs(1199)));
    layer3_outputs(2207) <= '0';
    layer3_outputs(2208) <= layer2_outputs(673);
    layer3_outputs(2209) <= not((layer2_outputs(1682)) and (layer2_outputs(511)));
    layer3_outputs(2210) <= (layer2_outputs(2377)) and (layer2_outputs(97));
    layer3_outputs(2211) <= not((layer2_outputs(2373)) and (layer2_outputs(1534)));
    layer3_outputs(2212) <= '1';
    layer3_outputs(2213) <= not(layer2_outputs(2370));
    layer3_outputs(2214) <= not(layer2_outputs(417));
    layer3_outputs(2215) <= not(layer2_outputs(623)) or (layer2_outputs(1615));
    layer3_outputs(2216) <= '1';
    layer3_outputs(2217) <= layer2_outputs(1952);
    layer3_outputs(2218) <= not((layer2_outputs(15)) and (layer2_outputs(2362)));
    layer3_outputs(2219) <= (layer2_outputs(1192)) and not (layer2_outputs(1497));
    layer3_outputs(2220) <= layer2_outputs(802);
    layer3_outputs(2221) <= '0';
    layer3_outputs(2222) <= (layer2_outputs(976)) and not (layer2_outputs(926));
    layer3_outputs(2223) <= layer2_outputs(1596);
    layer3_outputs(2224) <= layer2_outputs(830);
    layer3_outputs(2225) <= '1';
    layer3_outputs(2226) <= not(layer2_outputs(832)) or (layer2_outputs(1870));
    layer3_outputs(2227) <= '1';
    layer3_outputs(2228) <= layer2_outputs(68);
    layer3_outputs(2229) <= not((layer2_outputs(3)) or (layer2_outputs(2200)));
    layer3_outputs(2230) <= not(layer2_outputs(2010)) or (layer2_outputs(219));
    layer3_outputs(2231) <= not((layer2_outputs(1912)) or (layer2_outputs(1845)));
    layer3_outputs(2232) <= (layer2_outputs(1474)) and (layer2_outputs(1984));
    layer3_outputs(2233) <= layer2_outputs(78);
    layer3_outputs(2234) <= not((layer2_outputs(1851)) or (layer2_outputs(19)));
    layer3_outputs(2235) <= not(layer2_outputs(919));
    layer3_outputs(2236) <= (layer2_outputs(2278)) and not (layer2_outputs(210));
    layer3_outputs(2237) <= not(layer2_outputs(1383));
    layer3_outputs(2238) <= (layer2_outputs(1121)) and (layer2_outputs(1220));
    layer3_outputs(2239) <= layer2_outputs(533);
    layer3_outputs(2240) <= '0';
    layer3_outputs(2241) <= not(layer2_outputs(885));
    layer3_outputs(2242) <= not(layer2_outputs(1498));
    layer3_outputs(2243) <= '0';
    layer3_outputs(2244) <= not((layer2_outputs(1040)) or (layer2_outputs(1680)));
    layer3_outputs(2245) <= not(layer2_outputs(63)) or (layer2_outputs(2007));
    layer3_outputs(2246) <= (layer2_outputs(197)) or (layer2_outputs(1863));
    layer3_outputs(2247) <= layer2_outputs(175);
    layer3_outputs(2248) <= '0';
    layer3_outputs(2249) <= not(layer2_outputs(517));
    layer3_outputs(2250) <= '1';
    layer3_outputs(2251) <= (layer2_outputs(305)) or (layer2_outputs(499));
    layer3_outputs(2252) <= not(layer2_outputs(2416)) or (layer2_outputs(1458));
    layer3_outputs(2253) <= (layer2_outputs(80)) and not (layer2_outputs(2027));
    layer3_outputs(2254) <= '0';
    layer3_outputs(2255) <= not(layer2_outputs(2381));
    layer3_outputs(2256) <= layer2_outputs(1517);
    layer3_outputs(2257) <= not((layer2_outputs(631)) or (layer2_outputs(1139)));
    layer3_outputs(2258) <= (layer2_outputs(2558)) and (layer2_outputs(671));
    layer3_outputs(2259) <= '1';
    layer3_outputs(2260) <= not(layer2_outputs(16)) or (layer2_outputs(2008));
    layer3_outputs(2261) <= layer2_outputs(1591);
    layer3_outputs(2262) <= not(layer2_outputs(1117)) or (layer2_outputs(2000));
    layer3_outputs(2263) <= (layer2_outputs(453)) and (layer2_outputs(1571));
    layer3_outputs(2264) <= layer2_outputs(793);
    layer3_outputs(2265) <= not(layer2_outputs(563));
    layer3_outputs(2266) <= not(layer2_outputs(1587)) or (layer2_outputs(1713));
    layer3_outputs(2267) <= (layer2_outputs(1815)) and not (layer2_outputs(957));
    layer3_outputs(2268) <= layer2_outputs(1028);
    layer3_outputs(2269) <= not(layer2_outputs(2166));
    layer3_outputs(2270) <= layer2_outputs(930);
    layer3_outputs(2271) <= not(layer2_outputs(1717));
    layer3_outputs(2272) <= (layer2_outputs(1687)) or (layer2_outputs(933));
    layer3_outputs(2273) <= (layer2_outputs(59)) or (layer2_outputs(1832));
    layer3_outputs(2274) <= layer2_outputs(2220);
    layer3_outputs(2275) <= not(layer2_outputs(2553));
    layer3_outputs(2276) <= (layer2_outputs(1567)) and not (layer2_outputs(480));
    layer3_outputs(2277) <= (layer2_outputs(1123)) and (layer2_outputs(2374));
    layer3_outputs(2278) <= not((layer2_outputs(2059)) and (layer2_outputs(512)));
    layer3_outputs(2279) <= layer2_outputs(2241);
    layer3_outputs(2280) <= not(layer2_outputs(2009)) or (layer2_outputs(140));
    layer3_outputs(2281) <= not(layer2_outputs(2513));
    layer3_outputs(2282) <= not((layer2_outputs(108)) or (layer2_outputs(1720)));
    layer3_outputs(2283) <= (layer2_outputs(449)) and not (layer2_outputs(84));
    layer3_outputs(2284) <= not(layer2_outputs(323)) or (layer2_outputs(1511));
    layer3_outputs(2285) <= not(layer2_outputs(420));
    layer3_outputs(2286) <= not(layer2_outputs(270));
    layer3_outputs(2287) <= not(layer2_outputs(2075)) or (layer2_outputs(1166));
    layer3_outputs(2288) <= '0';
    layer3_outputs(2289) <= (layer2_outputs(1229)) and not (layer2_outputs(2537));
    layer3_outputs(2290) <= not((layer2_outputs(2055)) or (layer2_outputs(1165)));
    layer3_outputs(2291) <= '0';
    layer3_outputs(2292) <= layer2_outputs(985);
    layer3_outputs(2293) <= (layer2_outputs(555)) and (layer2_outputs(196));
    layer3_outputs(2294) <= (layer2_outputs(1885)) and not (layer2_outputs(151));
    layer3_outputs(2295) <= layer2_outputs(2173);
    layer3_outputs(2296) <= not((layer2_outputs(1675)) and (layer2_outputs(1489)));
    layer3_outputs(2297) <= not(layer2_outputs(1079));
    layer3_outputs(2298) <= not((layer2_outputs(1340)) and (layer2_outputs(796)));
    layer3_outputs(2299) <= '1';
    layer3_outputs(2300) <= (layer2_outputs(1824)) xor (layer2_outputs(2249));
    layer3_outputs(2301) <= not((layer2_outputs(387)) or (layer2_outputs(465)));
    layer3_outputs(2302) <= not((layer2_outputs(1939)) or (layer2_outputs(982)));
    layer3_outputs(2303) <= not(layer2_outputs(309)) or (layer2_outputs(2108));
    layer3_outputs(2304) <= (layer2_outputs(1253)) and not (layer2_outputs(101));
    layer3_outputs(2305) <= (layer2_outputs(2380)) and (layer2_outputs(1123));
    layer3_outputs(2306) <= not(layer2_outputs(157));
    layer3_outputs(2307) <= not(layer2_outputs(461));
    layer3_outputs(2308) <= not(layer2_outputs(949));
    layer3_outputs(2309) <= layer2_outputs(2389);
    layer3_outputs(2310) <= (layer2_outputs(1276)) or (layer2_outputs(2295));
    layer3_outputs(2311) <= layer2_outputs(2284);
    layer3_outputs(2312) <= layer2_outputs(1209);
    layer3_outputs(2313) <= not((layer2_outputs(1638)) and (layer2_outputs(1643)));
    layer3_outputs(2314) <= not(layer2_outputs(1562));
    layer3_outputs(2315) <= not(layer2_outputs(1622));
    layer3_outputs(2316) <= '0';
    layer3_outputs(2317) <= not((layer2_outputs(908)) or (layer2_outputs(1029)));
    layer3_outputs(2318) <= not(layer2_outputs(889));
    layer3_outputs(2319) <= not(layer2_outputs(840));
    layer3_outputs(2320) <= (layer2_outputs(426)) and not (layer2_outputs(2125));
    layer3_outputs(2321) <= not((layer2_outputs(1247)) or (layer2_outputs(586)));
    layer3_outputs(2322) <= (layer2_outputs(592)) or (layer2_outputs(2411));
    layer3_outputs(2323) <= '1';
    layer3_outputs(2324) <= not(layer2_outputs(2061)) or (layer2_outputs(1414));
    layer3_outputs(2325) <= '1';
    layer3_outputs(2326) <= layer2_outputs(2242);
    layer3_outputs(2327) <= (layer2_outputs(57)) or (layer2_outputs(1672));
    layer3_outputs(2328) <= (layer2_outputs(1294)) or (layer2_outputs(543));
    layer3_outputs(2329) <= not((layer2_outputs(111)) xor (layer2_outputs(1902)));
    layer3_outputs(2330) <= layer2_outputs(1260);
    layer3_outputs(2331) <= not((layer2_outputs(750)) and (layer2_outputs(1127)));
    layer3_outputs(2332) <= not(layer2_outputs(2130));
    layer3_outputs(2333) <= (layer2_outputs(1891)) and (layer2_outputs(1039));
    layer3_outputs(2334) <= layer2_outputs(1613);
    layer3_outputs(2335) <= not((layer2_outputs(1747)) or (layer2_outputs(2154)));
    layer3_outputs(2336) <= not(layer2_outputs(1932));
    layer3_outputs(2337) <= (layer2_outputs(67)) and not (layer2_outputs(1051));
    layer3_outputs(2338) <= '1';
    layer3_outputs(2339) <= not(layer2_outputs(2432)) or (layer2_outputs(1674));
    layer3_outputs(2340) <= not(layer2_outputs(2349)) or (layer2_outputs(2552));
    layer3_outputs(2341) <= (layer2_outputs(1374)) or (layer2_outputs(1764));
    layer3_outputs(2342) <= layer2_outputs(312);
    layer3_outputs(2343) <= not(layer2_outputs(290));
    layer3_outputs(2344) <= (layer2_outputs(1811)) and (layer2_outputs(2043));
    layer3_outputs(2345) <= '0';
    layer3_outputs(2346) <= (layer2_outputs(1711)) and not (layer2_outputs(796));
    layer3_outputs(2347) <= not(layer2_outputs(723));
    layer3_outputs(2348) <= not((layer2_outputs(1295)) xor (layer2_outputs(2182)));
    layer3_outputs(2349) <= not(layer2_outputs(1046)) or (layer2_outputs(905));
    layer3_outputs(2350) <= not(layer2_outputs(2367)) or (layer2_outputs(1759));
    layer3_outputs(2351) <= not(layer2_outputs(2066));
    layer3_outputs(2352) <= (layer2_outputs(1285)) and (layer2_outputs(1469));
    layer3_outputs(2353) <= (layer2_outputs(991)) and (layer2_outputs(1576));
    layer3_outputs(2354) <= not(layer2_outputs(522)) or (layer2_outputs(2081));
    layer3_outputs(2355) <= not((layer2_outputs(2243)) and (layer2_outputs(1397)));
    layer3_outputs(2356) <= not(layer2_outputs(2365));
    layer3_outputs(2357) <= layer2_outputs(2148);
    layer3_outputs(2358) <= (layer2_outputs(421)) and not (layer2_outputs(587));
    layer3_outputs(2359) <= not((layer2_outputs(2339)) and (layer2_outputs(1748)));
    layer3_outputs(2360) <= not(layer2_outputs(942));
    layer3_outputs(2361) <= layer2_outputs(1892);
    layer3_outputs(2362) <= (layer2_outputs(521)) or (layer2_outputs(1701));
    layer3_outputs(2363) <= (layer2_outputs(342)) xor (layer2_outputs(2168));
    layer3_outputs(2364) <= not((layer2_outputs(941)) and (layer2_outputs(1198)));
    layer3_outputs(2365) <= layer2_outputs(612);
    layer3_outputs(2366) <= (layer2_outputs(1008)) and not (layer2_outputs(1901));
    layer3_outputs(2367) <= '0';
    layer3_outputs(2368) <= not((layer2_outputs(1438)) and (layer2_outputs(2069)));
    layer3_outputs(2369) <= not((layer2_outputs(1622)) or (layer2_outputs(1891)));
    layer3_outputs(2370) <= not(layer2_outputs(1793));
    layer3_outputs(2371) <= (layer2_outputs(589)) and not (layer2_outputs(1202));
    layer3_outputs(2372) <= not(layer2_outputs(2320));
    layer3_outputs(2373) <= '0';
    layer3_outputs(2374) <= not(layer2_outputs(1962));
    layer3_outputs(2375) <= layer2_outputs(670);
    layer3_outputs(2376) <= (layer2_outputs(1868)) and not (layer2_outputs(405));
    layer3_outputs(2377) <= not((layer2_outputs(2025)) or (layer2_outputs(668)));
    layer3_outputs(2378) <= not(layer2_outputs(2403)) or (layer2_outputs(2335));
    layer3_outputs(2379) <= layer2_outputs(1751);
    layer3_outputs(2380) <= '0';
    layer3_outputs(2381) <= not(layer2_outputs(2109)) or (layer2_outputs(738));
    layer3_outputs(2382) <= layer2_outputs(1355);
    layer3_outputs(2383) <= (layer2_outputs(578)) and not (layer2_outputs(281));
    layer3_outputs(2384) <= layer2_outputs(2340);
    layer3_outputs(2385) <= (layer2_outputs(635)) and (layer2_outputs(2185));
    layer3_outputs(2386) <= not((layer2_outputs(521)) xor (layer2_outputs(1409)));
    layer3_outputs(2387) <= not((layer2_outputs(2281)) and (layer2_outputs(1604)));
    layer3_outputs(2388) <= layer2_outputs(987);
    layer3_outputs(2389) <= not(layer2_outputs(1262));
    layer3_outputs(2390) <= not(layer2_outputs(1454)) or (layer2_outputs(1783));
    layer3_outputs(2391) <= not((layer2_outputs(1222)) and (layer2_outputs(1667)));
    layer3_outputs(2392) <= '0';
    layer3_outputs(2393) <= layer2_outputs(1179);
    layer3_outputs(2394) <= not(layer2_outputs(525)) or (layer2_outputs(2029));
    layer3_outputs(2395) <= layer2_outputs(2326);
    layer3_outputs(2396) <= not((layer2_outputs(2254)) xor (layer2_outputs(492)));
    layer3_outputs(2397) <= layer2_outputs(253);
    layer3_outputs(2398) <= not(layer2_outputs(756));
    layer3_outputs(2399) <= '0';
    layer3_outputs(2400) <= not(layer2_outputs(1880));
    layer3_outputs(2401) <= not(layer2_outputs(755));
    layer3_outputs(2402) <= not(layer2_outputs(2186));
    layer3_outputs(2403) <= not(layer2_outputs(1273)) or (layer2_outputs(873));
    layer3_outputs(2404) <= layer2_outputs(1406);
    layer3_outputs(2405) <= not((layer2_outputs(2251)) and (layer2_outputs(1777)));
    layer3_outputs(2406) <= '1';
    layer3_outputs(2407) <= (layer2_outputs(1596)) and not (layer2_outputs(2491));
    layer3_outputs(2408) <= layer2_outputs(2031);
    layer3_outputs(2409) <= (layer2_outputs(294)) and (layer2_outputs(2278));
    layer3_outputs(2410) <= '0';
    layer3_outputs(2411) <= not((layer2_outputs(967)) or (layer2_outputs(127)));
    layer3_outputs(2412) <= not(layer2_outputs(229)) or (layer2_outputs(121));
    layer3_outputs(2413) <= not(layer2_outputs(617));
    layer3_outputs(2414) <= not((layer2_outputs(2404)) or (layer2_outputs(1617)));
    layer3_outputs(2415) <= layer2_outputs(1854);
    layer3_outputs(2416) <= not(layer2_outputs(566));
    layer3_outputs(2417) <= not(layer2_outputs(147));
    layer3_outputs(2418) <= not(layer2_outputs(11)) or (layer2_outputs(2260));
    layer3_outputs(2419) <= not(layer2_outputs(1178)) or (layer2_outputs(384));
    layer3_outputs(2420) <= (layer2_outputs(623)) and (layer2_outputs(1499));
    layer3_outputs(2421) <= not((layer2_outputs(626)) and (layer2_outputs(448)));
    layer3_outputs(2422) <= not(layer2_outputs(991)) or (layer2_outputs(2227));
    layer3_outputs(2423) <= not(layer2_outputs(1014));
    layer3_outputs(2424) <= '1';
    layer3_outputs(2425) <= not((layer2_outputs(592)) xor (layer2_outputs(146)));
    layer3_outputs(2426) <= (layer2_outputs(1750)) xor (layer2_outputs(2026));
    layer3_outputs(2427) <= (layer2_outputs(1494)) and not (layer2_outputs(2144));
    layer3_outputs(2428) <= (layer2_outputs(666)) and (layer2_outputs(2419));
    layer3_outputs(2429) <= layer2_outputs(1190);
    layer3_outputs(2430) <= (layer2_outputs(2297)) and not (layer2_outputs(1834));
    layer3_outputs(2431) <= (layer2_outputs(1519)) and not (layer2_outputs(2192));
    layer3_outputs(2432) <= '0';
    layer3_outputs(2433) <= '0';
    layer3_outputs(2434) <= '0';
    layer3_outputs(2435) <= layer2_outputs(717);
    layer3_outputs(2436) <= layer2_outputs(1236);
    layer3_outputs(2437) <= (layer2_outputs(266)) or (layer2_outputs(2463));
    layer3_outputs(2438) <= '1';
    layer3_outputs(2439) <= layer2_outputs(1572);
    layer3_outputs(2440) <= '0';
    layer3_outputs(2441) <= (layer2_outputs(88)) and not (layer2_outputs(2177));
    layer3_outputs(2442) <= (layer2_outputs(1626)) and (layer2_outputs(1273));
    layer3_outputs(2443) <= layer2_outputs(693);
    layer3_outputs(2444) <= (layer2_outputs(2115)) and not (layer2_outputs(2140));
    layer3_outputs(2445) <= layer2_outputs(1027);
    layer3_outputs(2446) <= not(layer2_outputs(2425));
    layer3_outputs(2447) <= not(layer2_outputs(2316)) or (layer2_outputs(1528));
    layer3_outputs(2448) <= layer2_outputs(44);
    layer3_outputs(2449) <= layer2_outputs(2219);
    layer3_outputs(2450) <= layer2_outputs(1120);
    layer3_outputs(2451) <= '1';
    layer3_outputs(2452) <= layer2_outputs(39);
    layer3_outputs(2453) <= '0';
    layer3_outputs(2454) <= '1';
    layer3_outputs(2455) <= (layer2_outputs(2205)) and not (layer2_outputs(1953));
    layer3_outputs(2456) <= not((layer2_outputs(93)) or (layer2_outputs(524)));
    layer3_outputs(2457) <= (layer2_outputs(1388)) or (layer2_outputs(1395));
    layer3_outputs(2458) <= not((layer2_outputs(4)) xor (layer2_outputs(332)));
    layer3_outputs(2459) <= not((layer2_outputs(269)) or (layer2_outputs(2283)));
    layer3_outputs(2460) <= not((layer2_outputs(488)) and (layer2_outputs(112)));
    layer3_outputs(2461) <= '1';
    layer3_outputs(2462) <= (layer2_outputs(595)) and not (layer2_outputs(2208));
    layer3_outputs(2463) <= not(layer2_outputs(1394));
    layer3_outputs(2464) <= '1';
    layer3_outputs(2465) <= '1';
    layer3_outputs(2466) <= (layer2_outputs(1257)) and (layer2_outputs(1696));
    layer3_outputs(2467) <= not((layer2_outputs(334)) xor (layer2_outputs(2040)));
    layer3_outputs(2468) <= (layer2_outputs(417)) and not (layer2_outputs(192));
    layer3_outputs(2469) <= not((layer2_outputs(544)) and (layer2_outputs(1281)));
    layer3_outputs(2470) <= (layer2_outputs(203)) and (layer2_outputs(34));
    layer3_outputs(2471) <= layer2_outputs(788);
    layer3_outputs(2472) <= not(layer2_outputs(1708));
    layer3_outputs(2473) <= (layer2_outputs(2007)) or (layer2_outputs(1156));
    layer3_outputs(2474) <= layer2_outputs(170);
    layer3_outputs(2475) <= (layer2_outputs(1268)) or (layer2_outputs(936));
    layer3_outputs(2476) <= not(layer2_outputs(390));
    layer3_outputs(2477) <= not(layer2_outputs(1532));
    layer3_outputs(2478) <= layer2_outputs(447);
    layer3_outputs(2479) <= layer2_outputs(577);
    layer3_outputs(2480) <= not((layer2_outputs(713)) and (layer2_outputs(1302)));
    layer3_outputs(2481) <= '1';
    layer3_outputs(2482) <= not(layer2_outputs(29));
    layer3_outputs(2483) <= (layer2_outputs(1397)) and not (layer2_outputs(1889));
    layer3_outputs(2484) <= (layer2_outputs(1548)) and not (layer2_outputs(2445));
    layer3_outputs(2485) <= layer2_outputs(1644);
    layer3_outputs(2486) <= layer2_outputs(2269);
    layer3_outputs(2487) <= '0';
    layer3_outputs(2488) <= not((layer2_outputs(918)) or (layer2_outputs(1322)));
    layer3_outputs(2489) <= (layer2_outputs(1479)) and not (layer2_outputs(2473));
    layer3_outputs(2490) <= '0';
    layer3_outputs(2491) <= not(layer2_outputs(168));
    layer3_outputs(2492) <= layer2_outputs(14);
    layer3_outputs(2493) <= not(layer2_outputs(2286));
    layer3_outputs(2494) <= not(layer2_outputs(502));
    layer3_outputs(2495) <= not(layer2_outputs(2064)) or (layer2_outputs(510));
    layer3_outputs(2496) <= (layer2_outputs(410)) and not (layer2_outputs(1879));
    layer3_outputs(2497) <= not(layer2_outputs(707));
    layer3_outputs(2498) <= (layer2_outputs(1296)) and not (layer2_outputs(1226));
    layer3_outputs(2499) <= (layer2_outputs(688)) and not (layer2_outputs(2138));
    layer3_outputs(2500) <= not(layer2_outputs(2184)) or (layer2_outputs(570));
    layer3_outputs(2501) <= not(layer2_outputs(1195));
    layer3_outputs(2502) <= (layer2_outputs(1476)) and (layer2_outputs(1862));
    layer3_outputs(2503) <= '0';
    layer3_outputs(2504) <= layer2_outputs(220);
    layer3_outputs(2505) <= (layer2_outputs(1953)) or (layer2_outputs(909));
    layer3_outputs(2506) <= layer2_outputs(379);
    layer3_outputs(2507) <= not(layer2_outputs(573));
    layer3_outputs(2508) <= layer2_outputs(2063);
    layer3_outputs(2509) <= '1';
    layer3_outputs(2510) <= '1';
    layer3_outputs(2511) <= '0';
    layer3_outputs(2512) <= layer2_outputs(457);
    layer3_outputs(2513) <= not((layer2_outputs(2353)) or (layer2_outputs(1725)));
    layer3_outputs(2514) <= layer2_outputs(142);
    layer3_outputs(2515) <= (layer2_outputs(576)) or (layer2_outputs(1886));
    layer3_outputs(2516) <= (layer2_outputs(1931)) or (layer2_outputs(2030));
    layer3_outputs(2517) <= not((layer2_outputs(0)) or (layer2_outputs(2242)));
    layer3_outputs(2518) <= '1';
    layer3_outputs(2519) <= (layer2_outputs(1411)) and not (layer2_outputs(2270));
    layer3_outputs(2520) <= not((layer2_outputs(1103)) and (layer2_outputs(393)));
    layer3_outputs(2521) <= layer2_outputs(2498);
    layer3_outputs(2522) <= (layer2_outputs(1648)) and not (layer2_outputs(1484));
    layer3_outputs(2523) <= (layer2_outputs(634)) and not (layer2_outputs(1867));
    layer3_outputs(2524) <= layer2_outputs(980);
    layer3_outputs(2525) <= (layer2_outputs(1202)) xor (layer2_outputs(1540));
    layer3_outputs(2526) <= layer2_outputs(1220);
    layer3_outputs(2527) <= not(layer2_outputs(378)) or (layer2_outputs(1716));
    layer3_outputs(2528) <= (layer2_outputs(2156)) and (layer2_outputs(1769));
    layer3_outputs(2529) <= layer2_outputs(1805);
    layer3_outputs(2530) <= not(layer2_outputs(1026));
    layer3_outputs(2531) <= layer2_outputs(517);
    layer3_outputs(2532) <= (layer2_outputs(2004)) and (layer2_outputs(524));
    layer3_outputs(2533) <= not(layer2_outputs(618)) or (layer2_outputs(850));
    layer3_outputs(2534) <= '0';
    layer3_outputs(2535) <= (layer2_outputs(2393)) and (layer2_outputs(2090));
    layer3_outputs(2536) <= (layer2_outputs(1998)) or (layer2_outputs(8));
    layer3_outputs(2537) <= (layer2_outputs(515)) and (layer2_outputs(1141));
    layer3_outputs(2538) <= not(layer2_outputs(68));
    layer3_outputs(2539) <= not((layer2_outputs(99)) and (layer2_outputs(1375)));
    layer3_outputs(2540) <= not(layer2_outputs(877));
    layer3_outputs(2541) <= (layer2_outputs(2065)) and not (layer2_outputs(534));
    layer3_outputs(2542) <= layer2_outputs(968);
    layer3_outputs(2543) <= (layer2_outputs(2188)) or (layer2_outputs(2101));
    layer3_outputs(2544) <= (layer2_outputs(790)) and not (layer2_outputs(1814));
    layer3_outputs(2545) <= (layer2_outputs(24)) and not (layer2_outputs(2292));
    layer3_outputs(2546) <= not(layer2_outputs(1677));
    layer3_outputs(2547) <= not((layer2_outputs(2227)) and (layer2_outputs(2359)));
    layer3_outputs(2548) <= not(layer2_outputs(319));
    layer3_outputs(2549) <= '0';
    layer3_outputs(2550) <= layer2_outputs(1032);
    layer3_outputs(2551) <= not((layer2_outputs(1227)) or (layer2_outputs(2006)));
    layer3_outputs(2552) <= (layer2_outputs(754)) and not (layer2_outputs(1610));
    layer3_outputs(2553) <= not(layer2_outputs(715));
    layer3_outputs(2554) <= layer2_outputs(1929);
    layer3_outputs(2555) <= not(layer2_outputs(1830));
    layer3_outputs(2556) <= layer2_outputs(2099);
    layer3_outputs(2557) <= (layer2_outputs(54)) and not (layer2_outputs(1384));
    layer3_outputs(2558) <= (layer2_outputs(236)) or (layer2_outputs(604));
    layer3_outputs(2559) <= not(layer2_outputs(1809)) or (layer2_outputs(1478));
    layer4_outputs(0) <= not(layer3_outputs(2542));
    layer4_outputs(1) <= not(layer3_outputs(2369)) or (layer3_outputs(357));
    layer4_outputs(2) <= layer3_outputs(888);
    layer4_outputs(3) <= layer3_outputs(2239);
    layer4_outputs(4) <= not((layer3_outputs(1786)) xor (layer3_outputs(189)));
    layer4_outputs(5) <= (layer3_outputs(1610)) and (layer3_outputs(452));
    layer4_outputs(6) <= (layer3_outputs(401)) or (layer3_outputs(182));
    layer4_outputs(7) <= '1';
    layer4_outputs(8) <= layer3_outputs(2276);
    layer4_outputs(9) <= (layer3_outputs(2518)) or (layer3_outputs(2464));
    layer4_outputs(10) <= not(layer3_outputs(493));
    layer4_outputs(11) <= not(layer3_outputs(2491));
    layer4_outputs(12) <= (layer3_outputs(2224)) and (layer3_outputs(1568));
    layer4_outputs(13) <= layer3_outputs(481);
    layer4_outputs(14) <= (layer3_outputs(2039)) and (layer3_outputs(2420));
    layer4_outputs(15) <= layer3_outputs(224);
    layer4_outputs(16) <= not(layer3_outputs(664));
    layer4_outputs(17) <= not(layer3_outputs(1898));
    layer4_outputs(18) <= layer3_outputs(2376);
    layer4_outputs(19) <= (layer3_outputs(411)) and not (layer3_outputs(38));
    layer4_outputs(20) <= not(layer3_outputs(487));
    layer4_outputs(21) <= not((layer3_outputs(662)) and (layer3_outputs(1455)));
    layer4_outputs(22) <= not(layer3_outputs(2352));
    layer4_outputs(23) <= not((layer3_outputs(1507)) and (layer3_outputs(2016)));
    layer4_outputs(24) <= not((layer3_outputs(223)) and (layer3_outputs(1853)));
    layer4_outputs(25) <= (layer3_outputs(249)) or (layer3_outputs(2117));
    layer4_outputs(26) <= not(layer3_outputs(1358)) or (layer3_outputs(72));
    layer4_outputs(27) <= (layer3_outputs(846)) and not (layer3_outputs(1308));
    layer4_outputs(28) <= not(layer3_outputs(367));
    layer4_outputs(29) <= layer3_outputs(376);
    layer4_outputs(30) <= (layer3_outputs(312)) and not (layer3_outputs(2437));
    layer4_outputs(31) <= not((layer3_outputs(2236)) xor (layer3_outputs(2021)));
    layer4_outputs(32) <= not(layer3_outputs(1546)) or (layer3_outputs(904));
    layer4_outputs(33) <= (layer3_outputs(868)) and (layer3_outputs(1516));
    layer4_outputs(34) <= not(layer3_outputs(932));
    layer4_outputs(35) <= (layer3_outputs(2150)) and not (layer3_outputs(1397));
    layer4_outputs(36) <= layer3_outputs(1313);
    layer4_outputs(37) <= (layer3_outputs(834)) and not (layer3_outputs(219));
    layer4_outputs(38) <= (layer3_outputs(2194)) or (layer3_outputs(381));
    layer4_outputs(39) <= not(layer3_outputs(1924));
    layer4_outputs(40) <= '0';
    layer4_outputs(41) <= not((layer3_outputs(1800)) or (layer3_outputs(737)));
    layer4_outputs(42) <= not(layer3_outputs(80)) or (layer3_outputs(177));
    layer4_outputs(43) <= layer3_outputs(1290);
    layer4_outputs(44) <= not(layer3_outputs(1987));
    layer4_outputs(45) <= layer3_outputs(432);
    layer4_outputs(46) <= (layer3_outputs(299)) and (layer3_outputs(1935));
    layer4_outputs(47) <= (layer3_outputs(1799)) xor (layer3_outputs(1334));
    layer4_outputs(48) <= not(layer3_outputs(144));
    layer4_outputs(49) <= not(layer3_outputs(708));
    layer4_outputs(50) <= (layer3_outputs(37)) and not (layer3_outputs(1121));
    layer4_outputs(51) <= not(layer3_outputs(612));
    layer4_outputs(52) <= not(layer3_outputs(700));
    layer4_outputs(53) <= (layer3_outputs(1606)) and not (layer3_outputs(141));
    layer4_outputs(54) <= (layer3_outputs(2257)) and (layer3_outputs(1396));
    layer4_outputs(55) <= not((layer3_outputs(2406)) xor (layer3_outputs(259)));
    layer4_outputs(56) <= (layer3_outputs(1725)) and (layer3_outputs(2127));
    layer4_outputs(57) <= not((layer3_outputs(614)) and (layer3_outputs(1061)));
    layer4_outputs(58) <= (layer3_outputs(981)) or (layer3_outputs(642));
    layer4_outputs(59) <= not((layer3_outputs(2180)) or (layer3_outputs(940)));
    layer4_outputs(60) <= (layer3_outputs(1885)) and not (layer3_outputs(1694));
    layer4_outputs(61) <= '0';
    layer4_outputs(62) <= not(layer3_outputs(2141));
    layer4_outputs(63) <= (layer3_outputs(627)) and not (layer3_outputs(777));
    layer4_outputs(64) <= (layer3_outputs(473)) and not (layer3_outputs(1014));
    layer4_outputs(65) <= (layer3_outputs(844)) or (layer3_outputs(2365));
    layer4_outputs(66) <= not((layer3_outputs(1874)) or (layer3_outputs(2509)));
    layer4_outputs(67) <= layer3_outputs(241);
    layer4_outputs(68) <= (layer3_outputs(1141)) and (layer3_outputs(64));
    layer4_outputs(69) <= layer3_outputs(1988);
    layer4_outputs(70) <= (layer3_outputs(1440)) and (layer3_outputs(1025));
    layer4_outputs(71) <= (layer3_outputs(1593)) and not (layer3_outputs(206));
    layer4_outputs(72) <= not(layer3_outputs(2307));
    layer4_outputs(73) <= not(layer3_outputs(2120));
    layer4_outputs(74) <= not((layer3_outputs(1336)) or (layer3_outputs(209)));
    layer4_outputs(75) <= not((layer3_outputs(1905)) and (layer3_outputs(1290)));
    layer4_outputs(76) <= (layer3_outputs(133)) or (layer3_outputs(1659));
    layer4_outputs(77) <= (layer3_outputs(1806)) and not (layer3_outputs(1703));
    layer4_outputs(78) <= not(layer3_outputs(1330));
    layer4_outputs(79) <= not(layer3_outputs(25));
    layer4_outputs(80) <= (layer3_outputs(212)) and not (layer3_outputs(1116));
    layer4_outputs(81) <= (layer3_outputs(763)) and (layer3_outputs(1441));
    layer4_outputs(82) <= not((layer3_outputs(327)) or (layer3_outputs(444)));
    layer4_outputs(83) <= not((layer3_outputs(2388)) or (layer3_outputs(682)));
    layer4_outputs(84) <= layer3_outputs(1762);
    layer4_outputs(85) <= not((layer3_outputs(2475)) and (layer3_outputs(732)));
    layer4_outputs(86) <= not((layer3_outputs(1128)) and (layer3_outputs(1716)));
    layer4_outputs(87) <= not(layer3_outputs(281));
    layer4_outputs(88) <= layer3_outputs(885);
    layer4_outputs(89) <= (layer3_outputs(343)) xor (layer3_outputs(2063));
    layer4_outputs(90) <= (layer3_outputs(1518)) xor (layer3_outputs(69));
    layer4_outputs(91) <= not((layer3_outputs(1758)) and (layer3_outputs(2393)));
    layer4_outputs(92) <= not(layer3_outputs(2090)) or (layer3_outputs(1581));
    layer4_outputs(93) <= layer3_outputs(1044);
    layer4_outputs(94) <= layer3_outputs(1134);
    layer4_outputs(95) <= not(layer3_outputs(33)) or (layer3_outputs(91));
    layer4_outputs(96) <= not(layer3_outputs(2305)) or (layer3_outputs(314));
    layer4_outputs(97) <= not(layer3_outputs(1674));
    layer4_outputs(98) <= not(layer3_outputs(1556)) or (layer3_outputs(600));
    layer4_outputs(99) <= not(layer3_outputs(869));
    layer4_outputs(100) <= layer3_outputs(852);
    layer4_outputs(101) <= layer3_outputs(287);
    layer4_outputs(102) <= (layer3_outputs(1785)) xor (layer3_outputs(488));
    layer4_outputs(103) <= not(layer3_outputs(1867)) or (layer3_outputs(1947));
    layer4_outputs(104) <= not((layer3_outputs(1863)) and (layer3_outputs(1218)));
    layer4_outputs(105) <= not((layer3_outputs(1994)) xor (layer3_outputs(362)));
    layer4_outputs(106) <= layer3_outputs(2431);
    layer4_outputs(107) <= not(layer3_outputs(2535));
    layer4_outputs(108) <= (layer3_outputs(2060)) xor (layer3_outputs(1056));
    layer4_outputs(109) <= '0';
    layer4_outputs(110) <= not((layer3_outputs(66)) or (layer3_outputs(1034)));
    layer4_outputs(111) <= not((layer3_outputs(1349)) xor (layer3_outputs(1106)));
    layer4_outputs(112) <= (layer3_outputs(2166)) and (layer3_outputs(2194));
    layer4_outputs(113) <= layer3_outputs(2073);
    layer4_outputs(114) <= not(layer3_outputs(1213)) or (layer3_outputs(777));
    layer4_outputs(115) <= not(layer3_outputs(2027));
    layer4_outputs(116) <= '0';
    layer4_outputs(117) <= not(layer3_outputs(2000));
    layer4_outputs(118) <= not(layer3_outputs(1563)) or (layer3_outputs(2202));
    layer4_outputs(119) <= layer3_outputs(2121);
    layer4_outputs(120) <= not(layer3_outputs(93)) or (layer3_outputs(1409));
    layer4_outputs(121) <= not((layer3_outputs(956)) and (layer3_outputs(393)));
    layer4_outputs(122) <= (layer3_outputs(344)) and not (layer3_outputs(992));
    layer4_outputs(123) <= (layer3_outputs(516)) or (layer3_outputs(976));
    layer4_outputs(124) <= not((layer3_outputs(44)) xor (layer3_outputs(2544)));
    layer4_outputs(125) <= not((layer3_outputs(1477)) or (layer3_outputs(2104)));
    layer4_outputs(126) <= not(layer3_outputs(1432));
    layer4_outputs(127) <= '0';
    layer4_outputs(128) <= not(layer3_outputs(1896));
    layer4_outputs(129) <= (layer3_outputs(2189)) and (layer3_outputs(2344));
    layer4_outputs(130) <= layer3_outputs(2526);
    layer4_outputs(131) <= not((layer3_outputs(2065)) or (layer3_outputs(1043)));
    layer4_outputs(132) <= (layer3_outputs(609)) and not (layer3_outputs(290));
    layer4_outputs(133) <= not(layer3_outputs(441)) or (layer3_outputs(718));
    layer4_outputs(134) <= not(layer3_outputs(1799));
    layer4_outputs(135) <= (layer3_outputs(1487)) or (layer3_outputs(2449));
    layer4_outputs(136) <= not(layer3_outputs(2435));
    layer4_outputs(137) <= layer3_outputs(1625);
    layer4_outputs(138) <= not(layer3_outputs(1692)) or (layer3_outputs(1363));
    layer4_outputs(139) <= not((layer3_outputs(2476)) or (layer3_outputs(1513)));
    layer4_outputs(140) <= not((layer3_outputs(541)) and (layer3_outputs(1312)));
    layer4_outputs(141) <= layer3_outputs(927);
    layer4_outputs(142) <= not(layer3_outputs(1999));
    layer4_outputs(143) <= layer3_outputs(2261);
    layer4_outputs(144) <= (layer3_outputs(2443)) and not (layer3_outputs(2143));
    layer4_outputs(145) <= layer3_outputs(678);
    layer4_outputs(146) <= not((layer3_outputs(284)) or (layer3_outputs(1288)));
    layer4_outputs(147) <= not(layer3_outputs(1474));
    layer4_outputs(148) <= (layer3_outputs(1247)) and (layer3_outputs(847));
    layer4_outputs(149) <= not(layer3_outputs(828));
    layer4_outputs(150) <= (layer3_outputs(135)) and not (layer3_outputs(1760));
    layer4_outputs(151) <= layer3_outputs(2096);
    layer4_outputs(152) <= (layer3_outputs(650)) and (layer3_outputs(1923));
    layer4_outputs(153) <= not(layer3_outputs(1265));
    layer4_outputs(154) <= (layer3_outputs(1089)) and (layer3_outputs(1214));
    layer4_outputs(155) <= not(layer3_outputs(1839));
    layer4_outputs(156) <= not(layer3_outputs(1815));
    layer4_outputs(157) <= layer3_outputs(1824);
    layer4_outputs(158) <= not(layer3_outputs(1957));
    layer4_outputs(159) <= not(layer3_outputs(72));
    layer4_outputs(160) <= (layer3_outputs(1609)) and (layer3_outputs(1638));
    layer4_outputs(161) <= not((layer3_outputs(2453)) and (layer3_outputs(808)));
    layer4_outputs(162) <= layer3_outputs(801);
    layer4_outputs(163) <= (layer3_outputs(2158)) and not (layer3_outputs(2322));
    layer4_outputs(164) <= (layer3_outputs(1152)) and (layer3_outputs(668));
    layer4_outputs(165) <= not(layer3_outputs(2040));
    layer4_outputs(166) <= not(layer3_outputs(710)) or (layer3_outputs(1400));
    layer4_outputs(167) <= layer3_outputs(1095);
    layer4_outputs(168) <= '1';
    layer4_outputs(169) <= not((layer3_outputs(2260)) and (layer3_outputs(870)));
    layer4_outputs(170) <= layer3_outputs(2042);
    layer4_outputs(171) <= (layer3_outputs(2195)) and not (layer3_outputs(1156));
    layer4_outputs(172) <= not((layer3_outputs(1112)) or (layer3_outputs(1584)));
    layer4_outputs(173) <= (layer3_outputs(1778)) and not (layer3_outputs(689));
    layer4_outputs(174) <= not(layer3_outputs(418)) or (layer3_outputs(629));
    layer4_outputs(175) <= '0';
    layer4_outputs(176) <= (layer3_outputs(107)) and (layer3_outputs(60));
    layer4_outputs(177) <= not(layer3_outputs(1623));
    layer4_outputs(178) <= (layer3_outputs(85)) xor (layer3_outputs(2057));
    layer4_outputs(179) <= (layer3_outputs(1500)) and not (layer3_outputs(623));
    layer4_outputs(180) <= (layer3_outputs(39)) xor (layer3_outputs(572));
    layer4_outputs(181) <= '0';
    layer4_outputs(182) <= '0';
    layer4_outputs(183) <= not(layer3_outputs(1927));
    layer4_outputs(184) <= (layer3_outputs(824)) xor (layer3_outputs(265));
    layer4_outputs(185) <= '1';
    layer4_outputs(186) <= '1';
    layer4_outputs(187) <= (layer3_outputs(1769)) and not (layer3_outputs(2214));
    layer4_outputs(188) <= not(layer3_outputs(804)) or (layer3_outputs(1318));
    layer4_outputs(189) <= not((layer3_outputs(975)) or (layer3_outputs(495)));
    layer4_outputs(190) <= not(layer3_outputs(394)) or (layer3_outputs(1395));
    layer4_outputs(191) <= layer3_outputs(1183);
    layer4_outputs(192) <= '0';
    layer4_outputs(193) <= layer3_outputs(1198);
    layer4_outputs(194) <= not(layer3_outputs(2249));
    layer4_outputs(195) <= layer3_outputs(749);
    layer4_outputs(196) <= (layer3_outputs(7)) and not (layer3_outputs(30));
    layer4_outputs(197) <= not(layer3_outputs(1514));
    layer4_outputs(198) <= (layer3_outputs(1159)) or (layer3_outputs(867));
    layer4_outputs(199) <= layer3_outputs(187);
    layer4_outputs(200) <= (layer3_outputs(795)) and not (layer3_outputs(1967));
    layer4_outputs(201) <= not((layer3_outputs(161)) or (layer3_outputs(1255)));
    layer4_outputs(202) <= not(layer3_outputs(1909));
    layer4_outputs(203) <= layer3_outputs(1602);
    layer4_outputs(204) <= not(layer3_outputs(2114));
    layer4_outputs(205) <= not(layer3_outputs(545));
    layer4_outputs(206) <= not((layer3_outputs(1929)) xor (layer3_outputs(651)));
    layer4_outputs(207) <= not((layer3_outputs(2235)) and (layer3_outputs(1101)));
    layer4_outputs(208) <= (layer3_outputs(416)) and not (layer3_outputs(487));
    layer4_outputs(209) <= layer3_outputs(486);
    layer4_outputs(210) <= '1';
    layer4_outputs(211) <= layer3_outputs(1618);
    layer4_outputs(212) <= (layer3_outputs(1809)) and not (layer3_outputs(196));
    layer4_outputs(213) <= not((layer3_outputs(1555)) or (layer3_outputs(1620)));
    layer4_outputs(214) <= '0';
    layer4_outputs(215) <= '0';
    layer4_outputs(216) <= layer3_outputs(149);
    layer4_outputs(217) <= layer3_outputs(82);
    layer4_outputs(218) <= not((layer3_outputs(1387)) xor (layer3_outputs(1820)));
    layer4_outputs(219) <= not(layer3_outputs(2274)) or (layer3_outputs(1061));
    layer4_outputs(220) <= layer3_outputs(0);
    layer4_outputs(221) <= (layer3_outputs(328)) and not (layer3_outputs(295));
    layer4_outputs(222) <= not(layer3_outputs(445));
    layer4_outputs(223) <= (layer3_outputs(1505)) and not (layer3_outputs(2213));
    layer4_outputs(224) <= layer3_outputs(2201);
    layer4_outputs(225) <= not(layer3_outputs(311));
    layer4_outputs(226) <= layer3_outputs(1586);
    layer4_outputs(227) <= not(layer3_outputs(1170));
    layer4_outputs(228) <= (layer3_outputs(406)) and (layer3_outputs(281));
    layer4_outputs(229) <= not((layer3_outputs(2428)) and (layer3_outputs(844)));
    layer4_outputs(230) <= '0';
    layer4_outputs(231) <= (layer3_outputs(550)) and not (layer3_outputs(385));
    layer4_outputs(232) <= layer3_outputs(1911);
    layer4_outputs(233) <= not((layer3_outputs(1077)) xor (layer3_outputs(2482)));
    layer4_outputs(234) <= not(layer3_outputs(2122)) or (layer3_outputs(1111));
    layer4_outputs(235) <= not((layer3_outputs(2446)) and (layer3_outputs(1787)));
    layer4_outputs(236) <= layer3_outputs(1398);
    layer4_outputs(237) <= not((layer3_outputs(317)) or (layer3_outputs(637)));
    layer4_outputs(238) <= not(layer3_outputs(2014));
    layer4_outputs(239) <= not(layer3_outputs(1012)) or (layer3_outputs(1902));
    layer4_outputs(240) <= layer3_outputs(1168);
    layer4_outputs(241) <= '0';
    layer4_outputs(242) <= (layer3_outputs(665)) or (layer3_outputs(863));
    layer4_outputs(243) <= '0';
    layer4_outputs(244) <= not((layer3_outputs(1757)) or (layer3_outputs(1456)));
    layer4_outputs(245) <= '1';
    layer4_outputs(246) <= not(layer3_outputs(2336));
    layer4_outputs(247) <= not(layer3_outputs(267)) or (layer3_outputs(1406));
    layer4_outputs(248) <= not((layer3_outputs(1732)) xor (layer3_outputs(820)));
    layer4_outputs(249) <= (layer3_outputs(1353)) xor (layer3_outputs(669));
    layer4_outputs(250) <= not((layer3_outputs(1435)) or (layer3_outputs(406)));
    layer4_outputs(251) <= not(layer3_outputs(103)) or (layer3_outputs(767));
    layer4_outputs(252) <= (layer3_outputs(290)) and (layer3_outputs(994));
    layer4_outputs(253) <= '0';
    layer4_outputs(254) <= (layer3_outputs(1567)) and (layer3_outputs(109));
    layer4_outputs(255) <= (layer3_outputs(2200)) or (layer3_outputs(556));
    layer4_outputs(256) <= layer3_outputs(1980);
    layer4_outputs(257) <= (layer3_outputs(440)) and (layer3_outputs(936));
    layer4_outputs(258) <= layer3_outputs(1400);
    layer4_outputs(259) <= not(layer3_outputs(991)) or (layer3_outputs(1645));
    layer4_outputs(260) <= (layer3_outputs(77)) and (layer3_outputs(436));
    layer4_outputs(261) <= not(layer3_outputs(304)) or (layer3_outputs(2474));
    layer4_outputs(262) <= not((layer3_outputs(2391)) or (layer3_outputs(2156)));
    layer4_outputs(263) <= '0';
    layer4_outputs(264) <= not(layer3_outputs(98));
    layer4_outputs(265) <= (layer3_outputs(1701)) or (layer3_outputs(1630));
    layer4_outputs(266) <= not(layer3_outputs(2444)) or (layer3_outputs(724));
    layer4_outputs(267) <= '0';
    layer4_outputs(268) <= '1';
    layer4_outputs(269) <= (layer3_outputs(1626)) and (layer3_outputs(7));
    layer4_outputs(270) <= (layer3_outputs(2409)) xor (layer3_outputs(2358));
    layer4_outputs(271) <= not(layer3_outputs(2122));
    layer4_outputs(272) <= not(layer3_outputs(1544));
    layer4_outputs(273) <= layer3_outputs(2255);
    layer4_outputs(274) <= not((layer3_outputs(2399)) and (layer3_outputs(1006)));
    layer4_outputs(275) <= layer3_outputs(1233);
    layer4_outputs(276) <= '0';
    layer4_outputs(277) <= layer3_outputs(875);
    layer4_outputs(278) <= (layer3_outputs(1463)) xor (layer3_outputs(478));
    layer4_outputs(279) <= not(layer3_outputs(2078));
    layer4_outputs(280) <= (layer3_outputs(977)) and not (layer3_outputs(779));
    layer4_outputs(281) <= '1';
    layer4_outputs(282) <= layer3_outputs(1291);
    layer4_outputs(283) <= not((layer3_outputs(112)) xor (layer3_outputs(1662)));
    layer4_outputs(284) <= not(layer3_outputs(943));
    layer4_outputs(285) <= not(layer3_outputs(263));
    layer4_outputs(286) <= (layer3_outputs(535)) or (layer3_outputs(232));
    layer4_outputs(287) <= layer3_outputs(273);
    layer4_outputs(288) <= not(layer3_outputs(1925)) or (layer3_outputs(2410));
    layer4_outputs(289) <= (layer3_outputs(195)) or (layer3_outputs(1521));
    layer4_outputs(290) <= (layer3_outputs(180)) and (layer3_outputs(1816));
    layer4_outputs(291) <= layer3_outputs(2142);
    layer4_outputs(292) <= (layer3_outputs(2268)) xor (layer3_outputs(957));
    layer4_outputs(293) <= not(layer3_outputs(1708));
    layer4_outputs(294) <= not((layer3_outputs(1730)) and (layer3_outputs(2032)));
    layer4_outputs(295) <= (layer3_outputs(446)) and not (layer3_outputs(17));
    layer4_outputs(296) <= not((layer3_outputs(1941)) and (layer3_outputs(2462)));
    layer4_outputs(297) <= not(layer3_outputs(611)) or (layer3_outputs(753));
    layer4_outputs(298) <= (layer3_outputs(849)) or (layer3_outputs(2133));
    layer4_outputs(299) <= not((layer3_outputs(278)) and (layer3_outputs(1632)));
    layer4_outputs(300) <= not((layer3_outputs(160)) or (layer3_outputs(291)));
    layer4_outputs(301) <= layer3_outputs(36);
    layer4_outputs(302) <= not(layer3_outputs(298)) or (layer3_outputs(1965));
    layer4_outputs(303) <= '1';
    layer4_outputs(304) <= (layer3_outputs(2340)) or (layer3_outputs(2493));
    layer4_outputs(305) <= '1';
    layer4_outputs(306) <= not((layer3_outputs(1642)) or (layer3_outputs(907)));
    layer4_outputs(307) <= not(layer3_outputs(2306));
    layer4_outputs(308) <= not(layer3_outputs(2052));
    layer4_outputs(309) <= layer3_outputs(2160);
    layer4_outputs(310) <= '1';
    layer4_outputs(311) <= not(layer3_outputs(1257));
    layer4_outputs(312) <= '0';
    layer4_outputs(313) <= not(layer3_outputs(1882)) or (layer3_outputs(194));
    layer4_outputs(314) <= not(layer3_outputs(2246));
    layer4_outputs(315) <= not(layer3_outputs(1427));
    layer4_outputs(316) <= not((layer3_outputs(1775)) or (layer3_outputs(46)));
    layer4_outputs(317) <= layer3_outputs(12);
    layer4_outputs(318) <= not(layer3_outputs(2362));
    layer4_outputs(319) <= (layer3_outputs(1553)) and not (layer3_outputs(1172));
    layer4_outputs(320) <= layer3_outputs(156);
    layer4_outputs(321) <= not(layer3_outputs(1936));
    layer4_outputs(322) <= layer3_outputs(2239);
    layer4_outputs(323) <= not(layer3_outputs(251));
    layer4_outputs(324) <= layer3_outputs(202);
    layer4_outputs(325) <= (layer3_outputs(1188)) and not (layer3_outputs(1666));
    layer4_outputs(326) <= not(layer3_outputs(84));
    layer4_outputs(327) <= layer3_outputs(1057);
    layer4_outputs(328) <= (layer3_outputs(391)) and not (layer3_outputs(1275));
    layer4_outputs(329) <= not((layer3_outputs(1038)) xor (layer3_outputs(1052)));
    layer4_outputs(330) <= not(layer3_outputs(2224));
    layer4_outputs(331) <= not(layer3_outputs(1256));
    layer4_outputs(332) <= (layer3_outputs(35)) and (layer3_outputs(2493));
    layer4_outputs(333) <= (layer3_outputs(382)) or (layer3_outputs(1928));
    layer4_outputs(334) <= not((layer3_outputs(83)) or (layer3_outputs(1851)));
    layer4_outputs(335) <= not(layer3_outputs(1792)) or (layer3_outputs(1132));
    layer4_outputs(336) <= not(layer3_outputs(1368)) or (layer3_outputs(2364));
    layer4_outputs(337) <= (layer3_outputs(246)) and (layer3_outputs(2397));
    layer4_outputs(338) <= not((layer3_outputs(1525)) or (layer3_outputs(366)));
    layer4_outputs(339) <= layer3_outputs(1993);
    layer4_outputs(340) <= layer3_outputs(156);
    layer4_outputs(341) <= (layer3_outputs(1776)) and (layer3_outputs(463));
    layer4_outputs(342) <= layer3_outputs(2031);
    layer4_outputs(343) <= layer3_outputs(949);
    layer4_outputs(344) <= not((layer3_outputs(569)) and (layer3_outputs(746)));
    layer4_outputs(345) <= not(layer3_outputs(2029));
    layer4_outputs(346) <= (layer3_outputs(345)) and not (layer3_outputs(717));
    layer4_outputs(347) <= not(layer3_outputs(282));
    layer4_outputs(348) <= not((layer3_outputs(1843)) and (layer3_outputs(1926)));
    layer4_outputs(349) <= not((layer3_outputs(94)) or (layer3_outputs(168)));
    layer4_outputs(350) <= not(layer3_outputs(423)) or (layer3_outputs(56));
    layer4_outputs(351) <= not((layer3_outputs(872)) or (layer3_outputs(1977)));
    layer4_outputs(352) <= layer3_outputs(2179);
    layer4_outputs(353) <= (layer3_outputs(525)) and not (layer3_outputs(1754));
    layer4_outputs(354) <= not(layer3_outputs(803)) or (layer3_outputs(2083));
    layer4_outputs(355) <= (layer3_outputs(1154)) or (layer3_outputs(43));
    layer4_outputs(356) <= not(layer3_outputs(1411));
    layer4_outputs(357) <= (layer3_outputs(559)) and (layer3_outputs(1251));
    layer4_outputs(358) <= (layer3_outputs(2218)) and not (layer3_outputs(1802));
    layer4_outputs(359) <= (layer3_outputs(2502)) and not (layer3_outputs(1835));
    layer4_outputs(360) <= '0';
    layer4_outputs(361) <= (layer3_outputs(1075)) and (layer3_outputs(1964));
    layer4_outputs(362) <= (layer3_outputs(1407)) and not (layer3_outputs(720));
    layer4_outputs(363) <= not(layer3_outputs(1981)) or (layer3_outputs(1502));
    layer4_outputs(364) <= (layer3_outputs(173)) and (layer3_outputs(533));
    layer4_outputs(365) <= not(layer3_outputs(350)) or (layer3_outputs(1874));
    layer4_outputs(366) <= (layer3_outputs(1767)) and not (layer3_outputs(986));
    layer4_outputs(367) <= (layer3_outputs(889)) or (layer3_outputs(1856));
    layer4_outputs(368) <= layer3_outputs(464);
    layer4_outputs(369) <= (layer3_outputs(518)) or (layer3_outputs(1316));
    layer4_outputs(370) <= not(layer3_outputs(1811));
    layer4_outputs(371) <= layer3_outputs(2467);
    layer4_outputs(372) <= not(layer3_outputs(1306));
    layer4_outputs(373) <= not(layer3_outputs(826)) or (layer3_outputs(857));
    layer4_outputs(374) <= (layer3_outputs(1264)) and (layer3_outputs(862));
    layer4_outputs(375) <= (layer3_outputs(114)) and not (layer3_outputs(1585));
    layer4_outputs(376) <= (layer3_outputs(649)) or (layer3_outputs(2049));
    layer4_outputs(377) <= (layer3_outputs(2126)) and (layer3_outputs(188));
    layer4_outputs(378) <= not((layer3_outputs(1771)) or (layer3_outputs(1452)));
    layer4_outputs(379) <= not((layer3_outputs(2319)) and (layer3_outputs(448)));
    layer4_outputs(380) <= not(layer3_outputs(543)) or (layer3_outputs(2262));
    layer4_outputs(381) <= not((layer3_outputs(1009)) and (layer3_outputs(1659)));
    layer4_outputs(382) <= not((layer3_outputs(2454)) or (layer3_outputs(1093)));
    layer4_outputs(383) <= '1';
    layer4_outputs(384) <= not(layer3_outputs(2068));
    layer4_outputs(385) <= '0';
    layer4_outputs(386) <= not(layer3_outputs(1257));
    layer4_outputs(387) <= not(layer3_outputs(2431));
    layer4_outputs(388) <= not(layer3_outputs(2412)) or (layer3_outputs(1423));
    layer4_outputs(389) <= layer3_outputs(2347);
    layer4_outputs(390) <= not((layer3_outputs(2219)) and (layer3_outputs(2105)));
    layer4_outputs(391) <= (layer3_outputs(1481)) and not (layer3_outputs(699));
    layer4_outputs(392) <= not(layer3_outputs(435));
    layer4_outputs(393) <= (layer3_outputs(531)) and (layer3_outputs(951));
    layer4_outputs(394) <= (layer3_outputs(2548)) or (layer3_outputs(394));
    layer4_outputs(395) <= layer3_outputs(638);
    layer4_outputs(396) <= '0';
    layer4_outputs(397) <= (layer3_outputs(2030)) and not (layer3_outputs(30));
    layer4_outputs(398) <= not(layer3_outputs(1499)) or (layer3_outputs(806));
    layer4_outputs(399) <= (layer3_outputs(264)) and (layer3_outputs(603));
    layer4_outputs(400) <= not((layer3_outputs(691)) or (layer3_outputs(1204)));
    layer4_outputs(401) <= not(layer3_outputs(2338));
    layer4_outputs(402) <= not((layer3_outputs(690)) and (layer3_outputs(1864)));
    layer4_outputs(403) <= not(layer3_outputs(789));
    layer4_outputs(404) <= not(layer3_outputs(1161));
    layer4_outputs(405) <= layer3_outputs(1928);
    layer4_outputs(406) <= not(layer3_outputs(2185));
    layer4_outputs(407) <= (layer3_outputs(723)) and not (layer3_outputs(132));
    layer4_outputs(408) <= not((layer3_outputs(840)) and (layer3_outputs(688)));
    layer4_outputs(409) <= '0';
    layer4_outputs(410) <= (layer3_outputs(108)) and (layer3_outputs(1757));
    layer4_outputs(411) <= not((layer3_outputs(209)) and (layer3_outputs(1860)));
    layer4_outputs(412) <= not(layer3_outputs(224));
    layer4_outputs(413) <= layer3_outputs(81);
    layer4_outputs(414) <= not((layer3_outputs(1888)) or (layer3_outputs(475)));
    layer4_outputs(415) <= '1';
    layer4_outputs(416) <= (layer3_outputs(2359)) and not (layer3_outputs(193));
    layer4_outputs(417) <= not(layer3_outputs(1575));
    layer4_outputs(418) <= layer3_outputs(1323);
    layer4_outputs(419) <= not(layer3_outputs(2209)) or (layer3_outputs(2430));
    layer4_outputs(420) <= '1';
    layer4_outputs(421) <= (layer3_outputs(2313)) and (layer3_outputs(27));
    layer4_outputs(422) <= (layer3_outputs(2465)) and not (layer3_outputs(105));
    layer4_outputs(423) <= not(layer3_outputs(2023));
    layer4_outputs(424) <= (layer3_outputs(333)) or (layer3_outputs(2251));
    layer4_outputs(425) <= '0';
    layer4_outputs(426) <= not((layer3_outputs(2146)) or (layer3_outputs(380)));
    layer4_outputs(427) <= not(layer3_outputs(2162));
    layer4_outputs(428) <= not(layer3_outputs(1092));
    layer4_outputs(429) <= (layer3_outputs(786)) and not (layer3_outputs(2135));
    layer4_outputs(430) <= not((layer3_outputs(1804)) or (layer3_outputs(2167)));
    layer4_outputs(431) <= not((layer3_outputs(828)) and (layer3_outputs(720)));
    layer4_outputs(432) <= layer3_outputs(2360);
    layer4_outputs(433) <= not(layer3_outputs(2097)) or (layer3_outputs(2308));
    layer4_outputs(434) <= (layer3_outputs(382)) and (layer3_outputs(2321));
    layer4_outputs(435) <= '0';
    layer4_outputs(436) <= layer3_outputs(58);
    layer4_outputs(437) <= layer3_outputs(311);
    layer4_outputs(438) <= not(layer3_outputs(438));
    layer4_outputs(439) <= (layer3_outputs(2159)) and not (layer3_outputs(990));
    layer4_outputs(440) <= not(layer3_outputs(139));
    layer4_outputs(441) <= (layer3_outputs(516)) or (layer3_outputs(2318));
    layer4_outputs(442) <= not(layer3_outputs(705));
    layer4_outputs(443) <= '0';
    layer4_outputs(444) <= not(layer3_outputs(2543));
    layer4_outputs(445) <= '0';
    layer4_outputs(446) <= layer3_outputs(1492);
    layer4_outputs(447) <= (layer3_outputs(2379)) and not (layer3_outputs(1405));
    layer4_outputs(448) <= not(layer3_outputs(1699));
    layer4_outputs(449) <= layer3_outputs(389);
    layer4_outputs(450) <= not(layer3_outputs(515)) or (layer3_outputs(956));
    layer4_outputs(451) <= layer3_outputs(2333);
    layer4_outputs(452) <= not(layer3_outputs(977));
    layer4_outputs(453) <= layer3_outputs(762);
    layer4_outputs(454) <= (layer3_outputs(1722)) and not (layer3_outputs(1968));
    layer4_outputs(455) <= not((layer3_outputs(2335)) and (layer3_outputs(1034)));
    layer4_outputs(456) <= layer3_outputs(146);
    layer4_outputs(457) <= not(layer3_outputs(650));
    layer4_outputs(458) <= layer3_outputs(1506);
    layer4_outputs(459) <= layer3_outputs(784);
    layer4_outputs(460) <= layer3_outputs(275);
    layer4_outputs(461) <= not(layer3_outputs(695));
    layer4_outputs(462) <= layer3_outputs(1681);
    layer4_outputs(463) <= (layer3_outputs(1712)) or (layer3_outputs(537));
    layer4_outputs(464) <= '1';
    layer4_outputs(465) <= (layer3_outputs(442)) and not (layer3_outputs(1493));
    layer4_outputs(466) <= not(layer3_outputs(1194));
    layer4_outputs(467) <= not(layer3_outputs(873)) or (layer3_outputs(968));
    layer4_outputs(468) <= not((layer3_outputs(387)) or (layer3_outputs(738)));
    layer4_outputs(469) <= (layer3_outputs(2333)) and (layer3_outputs(378));
    layer4_outputs(470) <= layer3_outputs(337);
    layer4_outputs(471) <= not(layer3_outputs(2211));
    layer4_outputs(472) <= '1';
    layer4_outputs(473) <= not(layer3_outputs(1071));
    layer4_outputs(474) <= not((layer3_outputs(1261)) and (layer3_outputs(1269)));
    layer4_outputs(475) <= not(layer3_outputs(208));
    layer4_outputs(476) <= '0';
    layer4_outputs(477) <= not(layer3_outputs(714)) or (layer3_outputs(519));
    layer4_outputs(478) <= (layer3_outputs(694)) and (layer3_outputs(841));
    layer4_outputs(479) <= (layer3_outputs(1696)) xor (layer3_outputs(1256));
    layer4_outputs(480) <= (layer3_outputs(1320)) or (layer3_outputs(395));
    layer4_outputs(481) <= not(layer3_outputs(2480));
    layer4_outputs(482) <= (layer3_outputs(2383)) and not (layer3_outputs(2372));
    layer4_outputs(483) <= '0';
    layer4_outputs(484) <= layer3_outputs(963);
    layer4_outputs(485) <= (layer3_outputs(1341)) and (layer3_outputs(1531));
    layer4_outputs(486) <= not(layer3_outputs(716));
    layer4_outputs(487) <= layer3_outputs(370);
    layer4_outputs(488) <= not(layer3_outputs(2208));
    layer4_outputs(489) <= layer3_outputs(1552);
    layer4_outputs(490) <= layer3_outputs(2147);
    layer4_outputs(491) <= not(layer3_outputs(1765));
    layer4_outputs(492) <= not((layer3_outputs(2235)) and (layer3_outputs(1554)));
    layer4_outputs(493) <= not((layer3_outputs(1347)) or (layer3_outputs(1952)));
    layer4_outputs(494) <= '1';
    layer4_outputs(495) <= (layer3_outputs(1212)) and (layer3_outputs(2270));
    layer4_outputs(496) <= layer3_outputs(544);
    layer4_outputs(497) <= layer3_outputs(578);
    layer4_outputs(498) <= not(layer3_outputs(2283)) or (layer3_outputs(312));
    layer4_outputs(499) <= not((layer3_outputs(1177)) xor (layer3_outputs(1852)));
    layer4_outputs(500) <= layer3_outputs(1553);
    layer4_outputs(501) <= not(layer3_outputs(1951));
    layer4_outputs(502) <= layer3_outputs(1106);
    layer4_outputs(503) <= '1';
    layer4_outputs(504) <= layer3_outputs(2461);
    layer4_outputs(505) <= (layer3_outputs(1022)) and not (layer3_outputs(1018));
    layer4_outputs(506) <= not(layer3_outputs(653));
    layer4_outputs(507) <= not((layer3_outputs(855)) and (layer3_outputs(1493)));
    layer4_outputs(508) <= not(layer3_outputs(1650)) or (layer3_outputs(2546));
    layer4_outputs(509) <= (layer3_outputs(1686)) and (layer3_outputs(493));
    layer4_outputs(510) <= not(layer3_outputs(371));
    layer4_outputs(511) <= not(layer3_outputs(1050));
    layer4_outputs(512) <= not((layer3_outputs(1074)) xor (layer3_outputs(827)));
    layer4_outputs(513) <= (layer3_outputs(1342)) and not (layer3_outputs(2498));
    layer4_outputs(514) <= not(layer3_outputs(2403)) or (layer3_outputs(1026));
    layer4_outputs(515) <= layer3_outputs(2489);
    layer4_outputs(516) <= (layer3_outputs(2442)) and not (layer3_outputs(1191));
    layer4_outputs(517) <= not(layer3_outputs(1896));
    layer4_outputs(518) <= '1';
    layer4_outputs(519) <= not(layer3_outputs(2105));
    layer4_outputs(520) <= not(layer3_outputs(428)) or (layer3_outputs(506));
    layer4_outputs(521) <= (layer3_outputs(739)) and not (layer3_outputs(321));
    layer4_outputs(522) <= not((layer3_outputs(421)) or (layer3_outputs(256)));
    layer4_outputs(523) <= not(layer3_outputs(1278)) or (layer3_outputs(1105));
    layer4_outputs(524) <= layer3_outputs(56);
    layer4_outputs(525) <= not(layer3_outputs(1058));
    layer4_outputs(526) <= layer3_outputs(2012);
    layer4_outputs(527) <= not(layer3_outputs(2476));
    layer4_outputs(528) <= (layer3_outputs(1525)) and not (layer3_outputs(1707));
    layer4_outputs(529) <= not(layer3_outputs(2061));
    layer4_outputs(530) <= not((layer3_outputs(2228)) and (layer3_outputs(2527)));
    layer4_outputs(531) <= layer3_outputs(1523);
    layer4_outputs(532) <= '1';
    layer4_outputs(533) <= (layer3_outputs(512)) and (layer3_outputs(2171));
    layer4_outputs(534) <= not((layer3_outputs(497)) or (layer3_outputs(1079)));
    layer4_outputs(535) <= layer3_outputs(2127);
    layer4_outputs(536) <= layer3_outputs(88);
    layer4_outputs(537) <= layer3_outputs(2494);
    layer4_outputs(538) <= layer3_outputs(1263);
    layer4_outputs(539) <= (layer3_outputs(829)) or (layer3_outputs(377));
    layer4_outputs(540) <= not(layer3_outputs(468)) or (layer3_outputs(2147));
    layer4_outputs(541) <= not(layer3_outputs(492));
    layer4_outputs(542) <= not(layer3_outputs(2470));
    layer4_outputs(543) <= layer3_outputs(1949);
    layer4_outputs(544) <= not(layer3_outputs(2272));
    layer4_outputs(545) <= not(layer3_outputs(1436));
    layer4_outputs(546) <= (layer3_outputs(886)) or (layer3_outputs(496));
    layer4_outputs(547) <= layer3_outputs(67);
    layer4_outputs(548) <= not(layer3_outputs(1125));
    layer4_outputs(549) <= (layer3_outputs(87)) xor (layer3_outputs(822));
    layer4_outputs(550) <= layer3_outputs(1355);
    layer4_outputs(551) <= (layer3_outputs(2478)) and not (layer3_outputs(2171));
    layer4_outputs(552) <= not(layer3_outputs(284));
    layer4_outputs(553) <= not((layer3_outputs(2373)) and (layer3_outputs(758)));
    layer4_outputs(554) <= layer3_outputs(33);
    layer4_outputs(555) <= layer3_outputs(2505);
    layer4_outputs(556) <= (layer3_outputs(1784)) or (layer3_outputs(1793));
    layer4_outputs(557) <= not((layer3_outputs(582)) and (layer3_outputs(1545)));
    layer4_outputs(558) <= not(layer3_outputs(1649));
    layer4_outputs(559) <= not((layer3_outputs(907)) xor (layer3_outputs(1954)));
    layer4_outputs(560) <= not((layer3_outputs(1003)) and (layer3_outputs(1346)));
    layer4_outputs(561) <= layer3_outputs(92);
    layer4_outputs(562) <= '1';
    layer4_outputs(563) <= (layer3_outputs(896)) and not (layer3_outputs(1921));
    layer4_outputs(564) <= '0';
    layer4_outputs(565) <= layer3_outputs(1989);
    layer4_outputs(566) <= (layer3_outputs(1042)) and not (layer3_outputs(1084));
    layer4_outputs(567) <= not((layer3_outputs(1689)) and (layer3_outputs(1496)));
    layer4_outputs(568) <= layer3_outputs(1388);
    layer4_outputs(569) <= not(layer3_outputs(980));
    layer4_outputs(570) <= not(layer3_outputs(1516));
    layer4_outputs(571) <= not(layer3_outputs(1420));
    layer4_outputs(572) <= (layer3_outputs(874)) and (layer3_outputs(1653));
    layer4_outputs(573) <= layer3_outputs(842);
    layer4_outputs(574) <= (layer3_outputs(1361)) and not (layer3_outputs(1790));
    layer4_outputs(575) <= not((layer3_outputs(1687)) or (layer3_outputs(654)));
    layer4_outputs(576) <= not(layer3_outputs(901));
    layer4_outputs(577) <= (layer3_outputs(1983)) and (layer3_outputs(2107));
    layer4_outputs(578) <= (layer3_outputs(1935)) and (layer3_outputs(566));
    layer4_outputs(579) <= layer3_outputs(797);
    layer4_outputs(580) <= not((layer3_outputs(42)) or (layer3_outputs(2501)));
    layer4_outputs(581) <= layer3_outputs(2193);
    layer4_outputs(582) <= '0';
    layer4_outputs(583) <= layer3_outputs(1202);
    layer4_outputs(584) <= (layer3_outputs(545)) and not (layer3_outputs(1945));
    layer4_outputs(585) <= '1';
    layer4_outputs(586) <= layer3_outputs(2371);
    layer4_outputs(587) <= '1';
    layer4_outputs(588) <= (layer3_outputs(2551)) and not (layer3_outputs(1094));
    layer4_outputs(589) <= not(layer3_outputs(2149)) or (layer3_outputs(59));
    layer4_outputs(590) <= not(layer3_outputs(1648)) or (layer3_outputs(1950));
    layer4_outputs(591) <= '0';
    layer4_outputs(592) <= (layer3_outputs(2322)) or (layer3_outputs(2045));
    layer4_outputs(593) <= (layer3_outputs(2524)) and not (layer3_outputs(1503));
    layer4_outputs(594) <= layer3_outputs(667);
    layer4_outputs(595) <= (layer3_outputs(1832)) xor (layer3_outputs(733));
    layer4_outputs(596) <= layer3_outputs(1800);
    layer4_outputs(597) <= not(layer3_outputs(317));
    layer4_outputs(598) <= layer3_outputs(221);
    layer4_outputs(599) <= not(layer3_outputs(1885));
    layer4_outputs(600) <= (layer3_outputs(116)) and (layer3_outputs(632));
    layer4_outputs(601) <= not(layer3_outputs(45));
    layer4_outputs(602) <= layer3_outputs(2482);
    layer4_outputs(603) <= layer3_outputs(1994);
    layer4_outputs(604) <= not((layer3_outputs(974)) and (layer3_outputs(2038)));
    layer4_outputs(605) <= layer3_outputs(559);
    layer4_outputs(606) <= (layer3_outputs(2422)) or (layer3_outputs(1973));
    layer4_outputs(607) <= (layer3_outputs(2126)) and not (layer3_outputs(386));
    layer4_outputs(608) <= (layer3_outputs(1521)) and not (layer3_outputs(1575));
    layer4_outputs(609) <= not((layer3_outputs(491)) and (layer3_outputs(1339)));
    layer4_outputs(610) <= not((layer3_outputs(5)) or (layer3_outputs(1230)));
    layer4_outputs(611) <= (layer3_outputs(191)) and not (layer3_outputs(1878));
    layer4_outputs(612) <= not((layer3_outputs(2225)) and (layer3_outputs(1586)));
    layer4_outputs(613) <= layer3_outputs(1533);
    layer4_outputs(614) <= layer3_outputs(617);
    layer4_outputs(615) <= not(layer3_outputs(760)) or (layer3_outputs(2220));
    layer4_outputs(616) <= not((layer3_outputs(485)) or (layer3_outputs(549)));
    layer4_outputs(617) <= (layer3_outputs(21)) and not (layer3_outputs(1470));
    layer4_outputs(618) <= not(layer3_outputs(2));
    layer4_outputs(619) <= layer3_outputs(170);
    layer4_outputs(620) <= not(layer3_outputs(1624));
    layer4_outputs(621) <= not(layer3_outputs(1588));
    layer4_outputs(622) <= not((layer3_outputs(1717)) and (layer3_outputs(1612)));
    layer4_outputs(623) <= not(layer3_outputs(597)) or (layer3_outputs(474));
    layer4_outputs(624) <= not(layer3_outputs(2528)) or (layer3_outputs(2056));
    layer4_outputs(625) <= (layer3_outputs(410)) and not (layer3_outputs(2534));
    layer4_outputs(626) <= layer3_outputs(2050);
    layer4_outputs(627) <= '0';
    layer4_outputs(628) <= '0';
    layer4_outputs(629) <= not(layer3_outputs(1732));
    layer4_outputs(630) <= not(layer3_outputs(2222));
    layer4_outputs(631) <= not(layer3_outputs(8));
    layer4_outputs(632) <= (layer3_outputs(2349)) or (layer3_outputs(1437));
    layer4_outputs(633) <= not(layer3_outputs(1263));
    layer4_outputs(634) <= (layer3_outputs(890)) and (layer3_outputs(459));
    layer4_outputs(635) <= (layer3_outputs(234)) and (layer3_outputs(2100));
    layer4_outputs(636) <= layer3_outputs(1423);
    layer4_outputs(637) <= not((layer3_outputs(2415)) or (layer3_outputs(2452)));
    layer4_outputs(638) <= not(layer3_outputs(875));
    layer4_outputs(639) <= layer3_outputs(1910);
    layer4_outputs(640) <= not(layer3_outputs(360));
    layer4_outputs(641) <= (layer3_outputs(2143)) and not (layer3_outputs(975));
    layer4_outputs(642) <= layer3_outputs(1526);
    layer4_outputs(643) <= not(layer3_outputs(2545));
    layer4_outputs(644) <= not(layer3_outputs(1226));
    layer4_outputs(645) <= '1';
    layer4_outputs(646) <= layer3_outputs(578);
    layer4_outputs(647) <= not(layer3_outputs(358)) or (layer3_outputs(2020));
    layer4_outputs(648) <= (layer3_outputs(484)) and (layer3_outputs(243));
    layer4_outputs(649) <= layer3_outputs(1363);
    layer4_outputs(650) <= (layer3_outputs(1025)) and (layer3_outputs(1070));
    layer4_outputs(651) <= (layer3_outputs(1333)) and not (layer3_outputs(515));
    layer4_outputs(652) <= not((layer3_outputs(2405)) xor (layer3_outputs(562)));
    layer4_outputs(653) <= '0';
    layer4_outputs(654) <= not((layer3_outputs(1917)) and (layer3_outputs(1962)));
    layer4_outputs(655) <= (layer3_outputs(272)) or (layer3_outputs(43));
    layer4_outputs(656) <= not(layer3_outputs(936)) or (layer3_outputs(41));
    layer4_outputs(657) <= layer3_outputs(1097);
    layer4_outputs(658) <= not(layer3_outputs(2360));
    layer4_outputs(659) <= not(layer3_outputs(2423));
    layer4_outputs(660) <= not(layer3_outputs(2402));
    layer4_outputs(661) <= layer3_outputs(1186);
    layer4_outputs(662) <= (layer3_outputs(1082)) and (layer3_outputs(233));
    layer4_outputs(663) <= (layer3_outputs(2411)) and not (layer3_outputs(2089));
    layer4_outputs(664) <= not(layer3_outputs(1020));
    layer4_outputs(665) <= (layer3_outputs(928)) xor (layer3_outputs(947));
    layer4_outputs(666) <= not((layer3_outputs(1680)) and (layer3_outputs(2532)));
    layer4_outputs(667) <= not(layer3_outputs(2472));
    layer4_outputs(668) <= not((layer3_outputs(792)) and (layer3_outputs(1592)));
    layer4_outputs(669) <= '1';
    layer4_outputs(670) <= '0';
    layer4_outputs(671) <= not((layer3_outputs(1569)) and (layer3_outputs(341)));
    layer4_outputs(672) <= layer3_outputs(1253);
    layer4_outputs(673) <= (layer3_outputs(216)) and not (layer3_outputs(701));
    layer4_outputs(674) <= not(layer3_outputs(47));
    layer4_outputs(675) <= not(layer3_outputs(750));
    layer4_outputs(676) <= layer3_outputs(1447);
    layer4_outputs(677) <= layer3_outputs(1857);
    layer4_outputs(678) <= '1';
    layer4_outputs(679) <= (layer3_outputs(772)) and not (layer3_outputs(734));
    layer4_outputs(680) <= layer3_outputs(1404);
    layer4_outputs(681) <= '1';
    layer4_outputs(682) <= (layer3_outputs(1171)) or (layer3_outputs(911));
    layer4_outputs(683) <= not(layer3_outputs(912));
    layer4_outputs(684) <= layer3_outputs(2309);
    layer4_outputs(685) <= not(layer3_outputs(2154)) or (layer3_outputs(2043));
    layer4_outputs(686) <= not(layer3_outputs(1227));
    layer4_outputs(687) <= not(layer3_outputs(625)) or (layer3_outputs(379));
    layer4_outputs(688) <= not(layer3_outputs(2456));
    layer4_outputs(689) <= not((layer3_outputs(1021)) xor (layer3_outputs(1463)));
    layer4_outputs(690) <= not(layer3_outputs(1000)) or (layer3_outputs(431));
    layer4_outputs(691) <= '0';
    layer4_outputs(692) <= (layer3_outputs(1072)) or (layer3_outputs(329));
    layer4_outputs(693) <= layer3_outputs(2159);
    layer4_outputs(694) <= (layer3_outputs(280)) and not (layer3_outputs(1289));
    layer4_outputs(695) <= not(layer3_outputs(468));
    layer4_outputs(696) <= not(layer3_outputs(1636));
    layer4_outputs(697) <= not(layer3_outputs(2005)) or (layer3_outputs(1197));
    layer4_outputs(698) <= layer3_outputs(1721);
    layer4_outputs(699) <= (layer3_outputs(2300)) or (layer3_outputs(1036));
    layer4_outputs(700) <= layer3_outputs(1622);
    layer4_outputs(701) <= (layer3_outputs(1270)) and not (layer3_outputs(358));
    layer4_outputs(702) <= not(layer3_outputs(483));
    layer4_outputs(703) <= not(layer3_outputs(1042));
    layer4_outputs(704) <= not(layer3_outputs(1522));
    layer4_outputs(705) <= not(layer3_outputs(2082));
    layer4_outputs(706) <= not((layer3_outputs(421)) and (layer3_outputs(1063)));
    layer4_outputs(707) <= (layer3_outputs(2175)) and not (layer3_outputs(1716));
    layer4_outputs(708) <= not(layer3_outputs(244));
    layer4_outputs(709) <= (layer3_outputs(229)) and (layer3_outputs(1764));
    layer4_outputs(710) <= not(layer3_outputs(201));
    layer4_outputs(711) <= not(layer3_outputs(2070));
    layer4_outputs(712) <= (layer3_outputs(1934)) and (layer3_outputs(1571));
    layer4_outputs(713) <= not((layer3_outputs(148)) or (layer3_outputs(1598)));
    layer4_outputs(714) <= not(layer3_outputs(621));
    layer4_outputs(715) <= (layer3_outputs(1889)) and not (layer3_outputs(1144));
    layer4_outputs(716) <= not(layer3_outputs(2123));
    layer4_outputs(717) <= layer3_outputs(706);
    layer4_outputs(718) <= '0';
    layer4_outputs(719) <= (layer3_outputs(2314)) and not (layer3_outputs(1579));
    layer4_outputs(720) <= (layer3_outputs(1747)) and not (layer3_outputs(1955));
    layer4_outputs(721) <= not(layer3_outputs(1774));
    layer4_outputs(722) <= not(layer3_outputs(2329));
    layer4_outputs(723) <= not(layer3_outputs(1153)) or (layer3_outputs(373));
    layer4_outputs(724) <= layer3_outputs(1426);
    layer4_outputs(725) <= not(layer3_outputs(1170));
    layer4_outputs(726) <= not(layer3_outputs(1734)) or (layer3_outputs(602));
    layer4_outputs(727) <= layer3_outputs(758);
    layer4_outputs(728) <= not((layer3_outputs(1772)) or (layer3_outputs(1544)));
    layer4_outputs(729) <= not(layer3_outputs(1518));
    layer4_outputs(730) <= not(layer3_outputs(957)) or (layer3_outputs(1274));
    layer4_outputs(731) <= (layer3_outputs(1645)) and not (layer3_outputs(2020));
    layer4_outputs(732) <= layer3_outputs(1347);
    layer4_outputs(733) <= (layer3_outputs(563)) and not (layer3_outputs(2047));
    layer4_outputs(734) <= not(layer3_outputs(949));
    layer4_outputs(735) <= layer3_outputs(1454);
    layer4_outputs(736) <= (layer3_outputs(2417)) and not (layer3_outputs(293));
    layer4_outputs(737) <= layer3_outputs(1233);
    layer4_outputs(738) <= not(layer3_outputs(1302));
    layer4_outputs(739) <= not(layer3_outputs(1685));
    layer4_outputs(740) <= not(layer3_outputs(2336));
    layer4_outputs(741) <= not(layer3_outputs(1010));
    layer4_outputs(742) <= layer3_outputs(1284);
    layer4_outputs(743) <= not((layer3_outputs(1724)) or (layer3_outputs(1357)));
    layer4_outputs(744) <= not(layer3_outputs(1802));
    layer4_outputs(745) <= (layer3_outputs(1578)) and (layer3_outputs(2018));
    layer4_outputs(746) <= (layer3_outputs(1968)) and not (layer3_outputs(652));
    layer4_outputs(747) <= (layer3_outputs(847)) and (layer3_outputs(2375));
    layer4_outputs(748) <= (layer3_outputs(2310)) or (layer3_outputs(1305));
    layer4_outputs(749) <= (layer3_outputs(2058)) or (layer3_outputs(1375));
    layer4_outputs(750) <= not((layer3_outputs(1227)) or (layer3_outputs(660)));
    layer4_outputs(751) <= (layer3_outputs(839)) and (layer3_outputs(2146));
    layer4_outputs(752) <= (layer3_outputs(2295)) or (layer3_outputs(1392));
    layer4_outputs(753) <= not(layer3_outputs(1346));
    layer4_outputs(754) <= layer3_outputs(2421);
    layer4_outputs(755) <= not(layer3_outputs(461));
    layer4_outputs(756) <= (layer3_outputs(1827)) and (layer3_outputs(101));
    layer4_outputs(757) <= layer3_outputs(1011);
    layer4_outputs(758) <= not(layer3_outputs(2243));
    layer4_outputs(759) <= (layer3_outputs(734)) xor (layer3_outputs(959));
    layer4_outputs(760) <= (layer3_outputs(655)) and (layer3_outputs(1647));
    layer4_outputs(761) <= not(layer3_outputs(90)) or (layer3_outputs(898));
    layer4_outputs(762) <= layer3_outputs(76);
    layer4_outputs(763) <= '1';
    layer4_outputs(764) <= not((layer3_outputs(465)) and (layer3_outputs(1331)));
    layer4_outputs(765) <= '0';
    layer4_outputs(766) <= not(layer3_outputs(2334));
    layer4_outputs(767) <= not(layer3_outputs(2238));
    layer4_outputs(768) <= not(layer3_outputs(2489));
    layer4_outputs(769) <= layer3_outputs(1895);
    layer4_outputs(770) <= not((layer3_outputs(348)) xor (layer3_outputs(668)));
    layer4_outputs(771) <= layer3_outputs(277);
    layer4_outputs(772) <= (layer3_outputs(631)) and not (layer3_outputs(1641));
    layer4_outputs(773) <= (layer3_outputs(1110)) and not (layer3_outputs(283));
    layer4_outputs(774) <= not((layer3_outputs(1035)) or (layer3_outputs(2148)));
    layer4_outputs(775) <= not(layer3_outputs(1307));
    layer4_outputs(776) <= (layer3_outputs(1908)) and not (layer3_outputs(239));
    layer4_outputs(777) <= layer3_outputs(61);
    layer4_outputs(778) <= not(layer3_outputs(964)) or (layer3_outputs(2230));
    layer4_outputs(779) <= '1';
    layer4_outputs(780) <= layer3_outputs(2553);
    layer4_outputs(781) <= (layer3_outputs(621)) and not (layer3_outputs(2441));
    layer4_outputs(782) <= not((layer3_outputs(1250)) and (layer3_outputs(517)));
    layer4_outputs(783) <= layer3_outputs(687);
    layer4_outputs(784) <= not(layer3_outputs(1284));
    layer4_outputs(785) <= not(layer3_outputs(218));
    layer4_outputs(786) <= not(layer3_outputs(1344));
    layer4_outputs(787) <= not(layer3_outputs(307));
    layer4_outputs(788) <= not(layer3_outputs(1501));
    layer4_outputs(789) <= (layer3_outputs(1880)) and not (layer3_outputs(507));
    layer4_outputs(790) <= not((layer3_outputs(917)) or (layer3_outputs(295)));
    layer4_outputs(791) <= not(layer3_outputs(997));
    layer4_outputs(792) <= not((layer3_outputs(1635)) and (layer3_outputs(950)));
    layer4_outputs(793) <= '1';
    layer4_outputs(794) <= not(layer3_outputs(862));
    layer4_outputs(795) <= not(layer3_outputs(1273));
    layer4_outputs(796) <= not(layer3_outputs(27));
    layer4_outputs(797) <= (layer3_outputs(1558)) and not (layer3_outputs(169));
    layer4_outputs(798) <= layer3_outputs(1234);
    layer4_outputs(799) <= layer3_outputs(1416);
    layer4_outputs(800) <= not(layer3_outputs(522));
    layer4_outputs(801) <= not(layer3_outputs(1774));
    layer4_outputs(802) <= (layer3_outputs(2180)) and not (layer3_outputs(1519));
    layer4_outputs(803) <= not(layer3_outputs(280));
    layer4_outputs(804) <= (layer3_outputs(23)) and not (layer3_outputs(1383));
    layer4_outputs(805) <= (layer3_outputs(316)) and (layer3_outputs(2093));
    layer4_outputs(806) <= '0';
    layer4_outputs(807) <= layer3_outputs(2196);
    layer4_outputs(808) <= (layer3_outputs(1538)) and not (layer3_outputs(1557));
    layer4_outputs(809) <= (layer3_outputs(1488)) or (layer3_outputs(1258));
    layer4_outputs(810) <= not(layer3_outputs(1096));
    layer4_outputs(811) <= not(layer3_outputs(1880));
    layer4_outputs(812) <= not((layer3_outputs(2429)) or (layer3_outputs(997)));
    layer4_outputs(813) <= not(layer3_outputs(157));
    layer4_outputs(814) <= (layer3_outputs(1796)) and not (layer3_outputs(1397));
    layer4_outputs(815) <= not(layer3_outputs(296));
    layer4_outputs(816) <= not(layer3_outputs(384));
    layer4_outputs(817) <= not(layer3_outputs(1494));
    layer4_outputs(818) <= (layer3_outputs(615)) and not (layer3_outputs(2342));
    layer4_outputs(819) <= not(layer3_outputs(2427)) or (layer3_outputs(1891));
    layer4_outputs(820) <= not(layer3_outputs(1543)) or (layer3_outputs(1761));
    layer4_outputs(821) <= layer3_outputs(652);
    layer4_outputs(822) <= layer3_outputs(476);
    layer4_outputs(823) <= not((layer3_outputs(1945)) and (layer3_outputs(1212)));
    layer4_outputs(824) <= (layer3_outputs(2181)) and not (layer3_outputs(646));
    layer4_outputs(825) <= (layer3_outputs(993)) and not (layer3_outputs(769));
    layer4_outputs(826) <= (layer3_outputs(155)) and not (layer3_outputs(1037));
    layer4_outputs(827) <= not(layer3_outputs(2076));
    layer4_outputs(828) <= not(layer3_outputs(1678)) or (layer3_outputs(2416));
    layer4_outputs(829) <= layer3_outputs(1939);
    layer4_outputs(830) <= not(layer3_outputs(1203)) or (layer3_outputs(1982));
    layer4_outputs(831) <= not((layer3_outputs(1606)) or (layer3_outputs(1101)));
    layer4_outputs(832) <= not(layer3_outputs(2038));
    layer4_outputs(833) <= layer3_outputs(1001);
    layer4_outputs(834) <= '0';
    layer4_outputs(835) <= (layer3_outputs(1952)) and not (layer3_outputs(2504));
    layer4_outputs(836) <= layer3_outputs(1859);
    layer4_outputs(837) <= not(layer3_outputs(1247));
    layer4_outputs(838) <= not(layer3_outputs(2381)) or (layer3_outputs(2516));
    layer4_outputs(839) <= (layer3_outputs(1309)) xor (layer3_outputs(1466));
    layer4_outputs(840) <= layer3_outputs(1147);
    layer4_outputs(841) <= not(layer3_outputs(1689));
    layer4_outputs(842) <= (layer3_outputs(2027)) and not (layer3_outputs(656));
    layer4_outputs(843) <= not(layer3_outputs(456));
    layer4_outputs(844) <= not(layer3_outputs(910));
    layer4_outputs(845) <= (layer3_outputs(659)) and not (layer3_outputs(497));
    layer4_outputs(846) <= not(layer3_outputs(1236)) or (layer3_outputs(1717));
    layer4_outputs(847) <= not((layer3_outputs(319)) or (layer3_outputs(500)));
    layer4_outputs(848) <= not((layer3_outputs(1711)) and (layer3_outputs(483)));
    layer4_outputs(849) <= (layer3_outputs(403)) and not (layer3_outputs(1414));
    layer4_outputs(850) <= '1';
    layer4_outputs(851) <= layer3_outputs(1675);
    layer4_outputs(852) <= (layer3_outputs(2039)) and (layer3_outputs(1278));
    layer4_outputs(853) <= not(layer3_outputs(2558));
    layer4_outputs(854) <= not(layer3_outputs(1959)) or (layer3_outputs(31));
    layer4_outputs(855) <= layer3_outputs(1843);
    layer4_outputs(856) <= layer3_outputs(178);
    layer4_outputs(857) <= not(layer3_outputs(2459)) or (layer3_outputs(2284));
    layer4_outputs(858) <= not(layer3_outputs(491));
    layer4_outputs(859) <= not((layer3_outputs(2264)) or (layer3_outputs(1848)));
    layer4_outputs(860) <= (layer3_outputs(585)) and not (layer3_outputs(1801));
    layer4_outputs(861) <= layer3_outputs(1446);
    layer4_outputs(862) <= not((layer3_outputs(2483)) and (layer3_outputs(2117)));
    layer4_outputs(863) <= (layer3_outputs(248)) and not (layer3_outputs(1356));
    layer4_outputs(864) <= layer3_outputs(1148);
    layer4_outputs(865) <= (layer3_outputs(1576)) and (layer3_outputs(2112));
    layer4_outputs(866) <= not(layer3_outputs(123));
    layer4_outputs(867) <= not(layer3_outputs(2142));
    layer4_outputs(868) <= '0';
    layer4_outputs(869) <= layer3_outputs(2186);
    layer4_outputs(870) <= not((layer3_outputs(554)) or (layer3_outputs(405)));
    layer4_outputs(871) <= not(layer3_outputs(1822));
    layer4_outputs(872) <= not(layer3_outputs(607)) or (layer3_outputs(1541));
    layer4_outputs(873) <= (layer3_outputs(764)) and (layer3_outputs(1051));
    layer4_outputs(874) <= (layer3_outputs(730)) or (layer3_outputs(1797));
    layer4_outputs(875) <= not(layer3_outputs(226));
    layer4_outputs(876) <= not(layer3_outputs(1742));
    layer4_outputs(877) <= not((layer3_outputs(182)) xor (layer3_outputs(364)));
    layer4_outputs(878) <= '1';
    layer4_outputs(879) <= (layer3_outputs(815)) or (layer3_outputs(2153));
    layer4_outputs(880) <= not(layer3_outputs(306)) or (layer3_outputs(120));
    layer4_outputs(881) <= not((layer3_outputs(2488)) xor (layer3_outputs(1552)));
    layer4_outputs(882) <= (layer3_outputs(1539)) and not (layer3_outputs(2400));
    layer4_outputs(883) <= not(layer3_outputs(590));
    layer4_outputs(884) <= not((layer3_outputs(612)) xor (layer3_outputs(1666)));
    layer4_outputs(885) <= '1';
    layer4_outputs(886) <= (layer3_outputs(2088)) and not (layer3_outputs(857));
    layer4_outputs(887) <= layer3_outputs(670);
    layer4_outputs(888) <= layer3_outputs(1202);
    layer4_outputs(889) <= layer3_outputs(1179);
    layer4_outputs(890) <= (layer3_outputs(1559)) and not (layer3_outputs(1287));
    layer4_outputs(891) <= layer3_outputs(1176);
    layer4_outputs(892) <= not(layer3_outputs(709));
    layer4_outputs(893) <= not(layer3_outputs(595)) or (layer3_outputs(575));
    layer4_outputs(894) <= layer3_outputs(1190);
    layer4_outputs(895) <= not((layer3_outputs(1668)) and (layer3_outputs(1973)));
    layer4_outputs(896) <= not(layer3_outputs(1324)) or (layer3_outputs(1821));
    layer4_outputs(897) <= '1';
    layer4_outputs(898) <= (layer3_outputs(1331)) and not (layer3_outputs(1846));
    layer4_outputs(899) <= layer3_outputs(2355);
    layer4_outputs(900) <= '0';
    layer4_outputs(901) <= not(layer3_outputs(261));
    layer4_outputs(902) <= layer3_outputs(1560);
    layer4_outputs(903) <= not(layer3_outputs(859));
    layer4_outputs(904) <= not((layer3_outputs(2269)) or (layer3_outputs(1744)));
    layer4_outputs(905) <= not((layer3_outputs(2320)) and (layer3_outputs(496)));
    layer4_outputs(906) <= not(layer3_outputs(2065));
    layer4_outputs(907) <= not(layer3_outputs(2189)) or (layer3_outputs(363));
    layer4_outputs(908) <= (layer3_outputs(28)) and (layer3_outputs(1217));
    layer4_outputs(909) <= not(layer3_outputs(1454));
    layer4_outputs(910) <= not(layer3_outputs(2361));
    layer4_outputs(911) <= (layer3_outputs(675)) or (layer3_outputs(2351));
    layer4_outputs(912) <= (layer3_outputs(640)) or (layer3_outputs(1828));
    layer4_outputs(913) <= not(layer3_outputs(891));
    layer4_outputs(914) <= not(layer3_outputs(1810));
    layer4_outputs(915) <= '1';
    layer4_outputs(916) <= not(layer3_outputs(704)) or (layer3_outputs(1698));
    layer4_outputs(917) <= not((layer3_outputs(785)) or (layer3_outputs(180)));
    layer4_outputs(918) <= (layer3_outputs(2001)) and not (layer3_outputs(760));
    layer4_outputs(919) <= not(layer3_outputs(1364));
    layer4_outputs(920) <= '1';
    layer4_outputs(921) <= (layer3_outputs(522)) and (layer3_outputs(2352));
    layer4_outputs(922) <= '1';
    layer4_outputs(923) <= layer3_outputs(1705);
    layer4_outputs(924) <= '1';
    layer4_outputs(925) <= layer3_outputs(1906);
    layer4_outputs(926) <= (layer3_outputs(670)) and (layer3_outputs(2317));
    layer4_outputs(927) <= not(layer3_outputs(2164));
    layer4_outputs(928) <= (layer3_outputs(2294)) xor (layer3_outputs(641));
    layer4_outputs(929) <= layer3_outputs(659);
    layer4_outputs(930) <= not(layer3_outputs(842));
    layer4_outputs(931) <= '1';
    layer4_outputs(932) <= not(layer3_outputs(1868));
    layer4_outputs(933) <= (layer3_outputs(1117)) and not (layer3_outputs(1617));
    layer4_outputs(934) <= not((layer3_outputs(447)) xor (layer3_outputs(419)));
    layer4_outputs(935) <= (layer3_outputs(77)) and (layer3_outputs(2198));
    layer4_outputs(936) <= not(layer3_outputs(2025)) or (layer3_outputs(1817));
    layer4_outputs(937) <= (layer3_outputs(1103)) and not (layer3_outputs(769));
    layer4_outputs(938) <= not(layer3_outputs(2228));
    layer4_outputs(939) <= not(layer3_outputs(1055));
    layer4_outputs(940) <= not((layer3_outputs(2492)) and (layer3_outputs(52)));
    layer4_outputs(941) <= (layer3_outputs(914)) and (layer3_outputs(1224));
    layer4_outputs(942) <= (layer3_outputs(1117)) and (layer3_outputs(1090));
    layer4_outputs(943) <= (layer3_outputs(1963)) and not (layer3_outputs(2034));
    layer4_outputs(944) <= not(layer3_outputs(588)) or (layer3_outputs(921));
    layer4_outputs(945) <= layer3_outputs(1919);
    layer4_outputs(946) <= layer3_outputs(1267);
    layer4_outputs(947) <= '1';
    layer4_outputs(948) <= not(layer3_outputs(2062));
    layer4_outputs(949) <= not(layer3_outputs(1208));
    layer4_outputs(950) <= (layer3_outputs(2241)) and not (layer3_outputs(682));
    layer4_outputs(951) <= (layer3_outputs(1947)) and not (layer3_outputs(1235));
    layer4_outputs(952) <= layer3_outputs(273);
    layer4_outputs(953) <= layer3_outputs(552);
    layer4_outputs(954) <= (layer3_outputs(579)) or (layer3_outputs(1215));
    layer4_outputs(955) <= (layer3_outputs(1498)) and not (layer3_outputs(2282));
    layer4_outputs(956) <= layer3_outputs(2374);
    layer4_outputs(957) <= not(layer3_outputs(1565)) or (layer3_outputs(2504));
    layer4_outputs(958) <= (layer3_outputs(1517)) or (layer3_outputs(1155));
    layer4_outputs(959) <= not(layer3_outputs(1546));
    layer4_outputs(960) <= not((layer3_outputs(2006)) and (layer3_outputs(594)));
    layer4_outputs(961) <= not(layer3_outputs(2116)) or (layer3_outputs(1676));
    layer4_outputs(962) <= not(layer3_outputs(1939)) or (layer3_outputs(353));
    layer4_outputs(963) <= (layer3_outputs(2484)) and (layer3_outputs(1760));
    layer4_outputs(964) <= not((layer3_outputs(2295)) and (layer3_outputs(1434)));
    layer4_outputs(965) <= not(layer3_outputs(92));
    layer4_outputs(966) <= (layer3_outputs(1663)) and (layer3_outputs(1446));
    layer4_outputs(967) <= (layer3_outputs(165)) and not (layer3_outputs(176));
    layer4_outputs(968) <= not(layer3_outputs(2395));
    layer4_outputs(969) <= not(layer3_outputs(843));
    layer4_outputs(970) <= layer3_outputs(1523);
    layer4_outputs(971) <= not((layer3_outputs(2533)) and (layer3_outputs(1852)));
    layer4_outputs(972) <= not(layer3_outputs(608));
    layer4_outputs(973) <= not((layer3_outputs(1985)) and (layer3_outputs(1867)));
    layer4_outputs(974) <= not(layer3_outputs(2551));
    layer4_outputs(975) <= layer3_outputs(1721);
    layer4_outputs(976) <= not(layer3_outputs(2427)) or (layer3_outputs(2402));
    layer4_outputs(977) <= '1';
    layer4_outputs(978) <= (layer3_outputs(1401)) and not (layer3_outputs(2031));
    layer4_outputs(979) <= not((layer3_outputs(1303)) and (layer3_outputs(1304)));
    layer4_outputs(980) <= '0';
    layer4_outputs(981) <= (layer3_outputs(1829)) xor (layer3_outputs(1150));
    layer4_outputs(982) <= layer3_outputs(320);
    layer4_outputs(983) <= layer3_outputs(1782);
    layer4_outputs(984) <= not((layer3_outputs(20)) xor (layer3_outputs(1086)));
    layer4_outputs(985) <= layer3_outputs(1582);
    layer4_outputs(986) <= not((layer3_outputs(2278)) or (layer3_outputs(1990)));
    layer4_outputs(987) <= (layer3_outputs(772)) and (layer3_outputs(429));
    layer4_outputs(988) <= (layer3_outputs(1429)) and not (layer3_outputs(1479));
    layer4_outputs(989) <= (layer3_outputs(586)) or (layer3_outputs(2380));
    layer4_outputs(990) <= (layer3_outputs(2507)) xor (layer3_outputs(26));
    layer4_outputs(991) <= layer3_outputs(2500);
    layer4_outputs(992) <= '1';
    layer4_outputs(993) <= (layer3_outputs(1555)) and not (layer3_outputs(2389));
    layer4_outputs(994) <= layer3_outputs(237);
    layer4_outputs(995) <= not(layer3_outputs(2369));
    layer4_outputs(996) <= not(layer3_outputs(897)) or (layer3_outputs(1932));
    layer4_outputs(997) <= layer3_outputs(749);
    layer4_outputs(998) <= layer3_outputs(473);
    layer4_outputs(999) <= not(layer3_outputs(938)) or (layer3_outputs(360));
    layer4_outputs(1000) <= not(layer3_outputs(796));
    layer4_outputs(1001) <= not((layer3_outputs(1181)) and (layer3_outputs(160)));
    layer4_outputs(1002) <= not(layer3_outputs(1983));
    layer4_outputs(1003) <= '1';
    layer4_outputs(1004) <= layer3_outputs(2348);
    layer4_outputs(1005) <= not(layer3_outputs(2304)) or (layer3_outputs(1577));
    layer4_outputs(1006) <= layer3_outputs(2071);
    layer4_outputs(1007) <= layer3_outputs(2485);
    layer4_outputs(1008) <= not(layer3_outputs(994));
    layer4_outputs(1009) <= not((layer3_outputs(1817)) xor (layer3_outputs(2340)));
    layer4_outputs(1010) <= not(layer3_outputs(361));
    layer4_outputs(1011) <= not(layer3_outputs(1426));
    layer4_outputs(1012) <= (layer3_outputs(908)) and not (layer3_outputs(1703));
    layer4_outputs(1013) <= layer3_outputs(434);
    layer4_outputs(1014) <= not(layer3_outputs(2124));
    layer4_outputs(1015) <= layer3_outputs(1437);
    layer4_outputs(1016) <= '1';
    layer4_outputs(1017) <= (layer3_outputs(518)) and (layer3_outputs(2523));
    layer4_outputs(1018) <= layer3_outputs(1870);
    layer4_outputs(1019) <= not(layer3_outputs(1959)) or (layer3_outputs(1634));
    layer4_outputs(1020) <= layer3_outputs(2530);
    layer4_outputs(1021) <= layer3_outputs(1142);
    layer4_outputs(1022) <= not(layer3_outputs(1814)) or (layer3_outputs(973));
    layer4_outputs(1023) <= not((layer3_outputs(617)) and (layer3_outputs(215)));
    layer4_outputs(1024) <= not(layer3_outputs(1770));
    layer4_outputs(1025) <= not((layer3_outputs(1032)) or (layer3_outputs(2096)));
    layer4_outputs(1026) <= layer3_outputs(1665);
    layer4_outputs(1027) <= (layer3_outputs(1030)) and (layer3_outputs(2302));
    layer4_outputs(1028) <= '1';
    layer4_outputs(1029) <= (layer3_outputs(1640)) or (layer3_outputs(1333));
    layer4_outputs(1030) <= not(layer3_outputs(1540));
    layer4_outputs(1031) <= not(layer3_outputs(1673));
    layer4_outputs(1032) <= not((layer3_outputs(2309)) or (layer3_outputs(1819)));
    layer4_outputs(1033) <= not(layer3_outputs(2321)) or (layer3_outputs(276));
    layer4_outputs(1034) <= layer3_outputs(770);
    layer4_outputs(1035) <= not(layer3_outputs(1930));
    layer4_outputs(1036) <= (layer3_outputs(664)) and not (layer3_outputs(1715));
    layer4_outputs(1037) <= layer3_outputs(658);
    layer4_outputs(1038) <= not((layer3_outputs(2013)) and (layer3_outputs(1771)));
    layer4_outputs(1039) <= (layer3_outputs(2354)) or (layer3_outputs(1711));
    layer4_outputs(1040) <= not(layer3_outputs(2190));
    layer4_outputs(1041) <= not(layer3_outputs(579));
    layer4_outputs(1042) <= layer3_outputs(1260);
    layer4_outputs(1043) <= '1';
    layer4_outputs(1044) <= not(layer3_outputs(2197));
    layer4_outputs(1045) <= layer3_outputs(213);
    layer4_outputs(1046) <= not(layer3_outputs(464));
    layer4_outputs(1047) <= not((layer3_outputs(2148)) and (layer3_outputs(1870)));
    layer4_outputs(1048) <= layer3_outputs(2061);
    layer4_outputs(1049) <= not((layer3_outputs(893)) or (layer3_outputs(243)));
    layer4_outputs(1050) <= not(layer3_outputs(943));
    layer4_outputs(1051) <= (layer3_outputs(2161)) and not (layer3_outputs(2080));
    layer4_outputs(1052) <= layer3_outputs(337);
    layer4_outputs(1053) <= '0';
    layer4_outputs(1054) <= (layer3_outputs(371)) and not (layer3_outputs(560));
    layer4_outputs(1055) <= layer3_outputs(1953);
    layer4_outputs(1056) <= layer3_outputs(1706);
    layer4_outputs(1057) <= not(layer3_outputs(470));
    layer4_outputs(1058) <= not(layer3_outputs(216)) or (layer3_outputs(1275));
    layer4_outputs(1059) <= not(layer3_outputs(402));
    layer4_outputs(1060) <= not((layer3_outputs(1425)) or (layer3_outputs(1357)));
    layer4_outputs(1061) <= not((layer3_outputs(620)) or (layer3_outputs(1113)));
    layer4_outputs(1062) <= not((layer3_outputs(570)) and (layer3_outputs(2511)));
    layer4_outputs(1063) <= not((layer3_outputs(2435)) and (layer3_outputs(2036)));
    layer4_outputs(1064) <= not(layer3_outputs(2197));
    layer4_outputs(1065) <= layer3_outputs(1998);
    layer4_outputs(1066) <= (layer3_outputs(1577)) and (layer3_outputs(1380));
    layer4_outputs(1067) <= not(layer3_outputs(1251));
    layer4_outputs(1068) <= not(layer3_outputs(179)) or (layer3_outputs(712));
    layer4_outputs(1069) <= (layer3_outputs(523)) or (layer3_outputs(1892));
    layer4_outputs(1070) <= layer3_outputs(2041);
    layer4_outputs(1071) <= not(layer3_outputs(118)) or (layer3_outputs(1780));
    layer4_outputs(1072) <= (layer3_outputs(1024)) and not (layer3_outputs(2259));
    layer4_outputs(1073) <= not(layer3_outputs(178));
    layer4_outputs(1074) <= layer3_outputs(1105);
    layer4_outputs(1075) <= not(layer3_outputs(541));
    layer4_outputs(1076) <= not(layer3_outputs(1)) or (layer3_outputs(1690));
    layer4_outputs(1077) <= not((layer3_outputs(965)) or (layer3_outputs(681)));
    layer4_outputs(1078) <= layer3_outputs(834);
    layer4_outputs(1079) <= layer3_outputs(2055);
    layer4_outputs(1080) <= (layer3_outputs(141)) or (layer3_outputs(960));
    layer4_outputs(1081) <= not(layer3_outputs(1990));
    layer4_outputs(1082) <= (layer3_outputs(1312)) or (layer3_outputs(2426));
    layer4_outputs(1083) <= not(layer3_outputs(1583));
    layer4_outputs(1084) <= not(layer3_outputs(1000));
    layer4_outputs(1085) <= layer3_outputs(60);
    layer4_outputs(1086) <= not(layer3_outputs(1325));
    layer4_outputs(1087) <= not(layer3_outputs(884)) or (layer3_outputs(1729));
    layer4_outputs(1088) <= layer3_outputs(2532);
    layer4_outputs(1089) <= (layer3_outputs(2446)) or (layer3_outputs(1673));
    layer4_outputs(1090) <= (layer3_outputs(230)) or (layer3_outputs(137));
    layer4_outputs(1091) <= layer3_outputs(1143);
    layer4_outputs(1092) <= not((layer3_outputs(1655)) xor (layer3_outputs(301)));
    layer4_outputs(1093) <= not(layer3_outputs(37));
    layer4_outputs(1094) <= not(layer3_outputs(159)) or (layer3_outputs(256));
    layer4_outputs(1095) <= not(layer3_outputs(1533));
    layer4_outputs(1096) <= layer3_outputs(183);
    layer4_outputs(1097) <= not(layer3_outputs(278)) or (layer3_outputs(2281));
    layer4_outputs(1098) <= not(layer3_outputs(1120)) or (layer3_outputs(1503));
    layer4_outputs(1099) <= not(layer3_outputs(731));
    layer4_outputs(1100) <= '0';
    layer4_outputs(1101) <= (layer3_outputs(1726)) or (layer3_outputs(488));
    layer4_outputs(1102) <= layer3_outputs(630);
    layer4_outputs(1103) <= not(layer3_outputs(2162)) or (layer3_outputs(2206));
    layer4_outputs(1104) <= layer3_outputs(510);
    layer4_outputs(1105) <= layer3_outputs(375);
    layer4_outputs(1106) <= layer3_outputs(384);
    layer4_outputs(1107) <= not(layer3_outputs(998));
    layer4_outputs(1108) <= (layer3_outputs(386)) or (layer3_outputs(2320));
    layer4_outputs(1109) <= layer3_outputs(1613);
    layer4_outputs(1110) <= not(layer3_outputs(1374));
    layer4_outputs(1111) <= not(layer3_outputs(2238));
    layer4_outputs(1112) <= (layer3_outputs(752)) and not (layer3_outputs(1637));
    layer4_outputs(1113) <= '1';
    layer4_outputs(1114) <= not(layer3_outputs(2506));
    layer4_outputs(1115) <= not((layer3_outputs(198)) or (layer3_outputs(1282)));
    layer4_outputs(1116) <= not((layer3_outputs(2384)) and (layer3_outputs(171)));
    layer4_outputs(1117) <= not(layer3_outputs(300));
    layer4_outputs(1118) <= layer3_outputs(86);
    layer4_outputs(1119) <= not((layer3_outputs(1211)) xor (layer3_outputs(1987)));
    layer4_outputs(1120) <= '1';
    layer4_outputs(1121) <= not(layer3_outputs(816)) or (layer3_outputs(1382));
    layer4_outputs(1122) <= layer3_outputs(97);
    layer4_outputs(1123) <= (layer3_outputs(968)) or (layer3_outputs(1168));
    layer4_outputs(1124) <= (layer3_outputs(654)) or (layer3_outputs(1584));
    layer4_outputs(1125) <= (layer3_outputs(2028)) xor (layer3_outputs(2033));
    layer4_outputs(1126) <= not((layer3_outputs(1081)) or (layer3_outputs(2443)));
    layer4_outputs(1127) <= not(layer3_outputs(566)) or (layer3_outputs(636));
    layer4_outputs(1128) <= '1';
    layer4_outputs(1129) <= not(layer3_outputs(135)) or (layer3_outputs(2508));
    layer4_outputs(1130) <= '0';
    layer4_outputs(1131) <= layer3_outputs(1588);
    layer4_outputs(1132) <= not(layer3_outputs(2357));
    layer4_outputs(1133) <= (layer3_outputs(1461)) or (layer3_outputs(1887));
    layer4_outputs(1134) <= (layer3_outputs(2380)) and not (layer3_outputs(24));
    layer4_outputs(1135) <= not(layer3_outputs(822));
    layer4_outputs(1136) <= (layer3_outputs(1883)) xor (layer3_outputs(1611));
    layer4_outputs(1137) <= not(layer3_outputs(193));
    layer4_outputs(1138) <= layer3_outputs(1904);
    layer4_outputs(1139) <= layer3_outputs(1104);
    layer4_outputs(1140) <= not(layer3_outputs(1136)) or (layer3_outputs(179));
    layer4_outputs(1141) <= '1';
    layer4_outputs(1142) <= (layer3_outputs(2182)) xor (layer3_outputs(908));
    layer4_outputs(1143) <= not(layer3_outputs(1342));
    layer4_outputs(1144) <= (layer3_outputs(2044)) xor (layer3_outputs(2013));
    layer4_outputs(1145) <= not(layer3_outputs(1982));
    layer4_outputs(1146) <= '1';
    layer4_outputs(1147) <= (layer3_outputs(643)) and not (layer3_outputs(1886));
    layer4_outputs(1148) <= layer3_outputs(583);
    layer4_outputs(1149) <= (layer3_outputs(1115)) and (layer3_outputs(1198));
    layer4_outputs(1150) <= (layer3_outputs(2485)) and (layer3_outputs(2245));
    layer4_outputs(1151) <= layer3_outputs(939);
    layer4_outputs(1152) <= not(layer3_outputs(2540));
    layer4_outputs(1153) <= not((layer3_outputs(2303)) and (layer3_outputs(2438)));
    layer4_outputs(1154) <= (layer3_outputs(2396)) and not (layer3_outputs(70));
    layer4_outputs(1155) <= (layer3_outputs(346)) and (layer3_outputs(1219));
    layer4_outputs(1156) <= '0';
    layer4_outputs(1157) <= not(layer3_outputs(2313));
    layer4_outputs(1158) <= (layer3_outputs(2001)) and not (layer3_outputs(1356));
    layer4_outputs(1159) <= layer3_outputs(2116);
    layer4_outputs(1160) <= not(layer3_outputs(1831));
    layer4_outputs(1161) <= not(layer3_outputs(2480));
    layer4_outputs(1162) <= not(layer3_outputs(1390));
    layer4_outputs(1163) <= not(layer3_outputs(771)) or (layer3_outputs(730));
    layer4_outputs(1164) <= (layer3_outputs(1809)) and (layer3_outputs(1998));
    layer4_outputs(1165) <= '0';
    layer4_outputs(1166) <= not(layer3_outputs(1362));
    layer4_outputs(1167) <= not((layer3_outputs(1216)) or (layer3_outputs(1778)));
    layer4_outputs(1168) <= not(layer3_outputs(674));
    layer4_outputs(1169) <= not(layer3_outputs(108)) or (layer3_outputs(164));
    layer4_outputs(1170) <= (layer3_outputs(1328)) and not (layer3_outputs(2111));
    layer4_outputs(1171) <= not(layer3_outputs(1073)) or (layer3_outputs(945));
    layer4_outputs(1172) <= not((layer3_outputs(989)) or (layer3_outputs(1834)));
    layer4_outputs(1173) <= not(layer3_outputs(660));
    layer4_outputs(1174) <= (layer3_outputs(1195)) or (layer3_outputs(1633));
    layer4_outputs(1175) <= layer3_outputs(1937);
    layer4_outputs(1176) <= layer3_outputs(413);
    layer4_outputs(1177) <= not((layer3_outputs(1729)) or (layer3_outputs(941)));
    layer4_outputs(1178) <= not(layer3_outputs(2131)) or (layer3_outputs(450));
    layer4_outputs(1179) <= layer3_outputs(2234);
    layer4_outputs(1180) <= layer3_outputs(1940);
    layer4_outputs(1181) <= (layer3_outputs(67)) and (layer3_outputs(2000));
    layer4_outputs(1182) <= (layer3_outputs(2408)) and (layer3_outputs(1727));
    layer4_outputs(1183) <= layer3_outputs(1846);
    layer4_outputs(1184) <= not((layer3_outputs(865)) or (layer3_outputs(2152)));
    layer4_outputs(1185) <= not(layer3_outputs(307));
    layer4_outputs(1186) <= '0';
    layer4_outputs(1187) <= not(layer3_outputs(1460));
    layer4_outputs(1188) <= not(layer3_outputs(437));
    layer4_outputs(1189) <= not(layer3_outputs(882));
    layer4_outputs(1190) <= layer3_outputs(2441);
    layer4_outputs(1191) <= (layer3_outputs(4)) or (layer3_outputs(1511));
    layer4_outputs(1192) <= not(layer3_outputs(32));
    layer4_outputs(1193) <= '0';
    layer4_outputs(1194) <= not(layer3_outputs(1008));
    layer4_outputs(1195) <= not(layer3_outputs(804)) or (layer3_outputs(1825));
    layer4_outputs(1196) <= (layer3_outputs(1390)) and not (layer3_outputs(1039));
    layer4_outputs(1197) <= (layer3_outputs(258)) and not (layer3_outputs(683));
    layer4_outputs(1198) <= not((layer3_outputs(97)) and (layer3_outputs(752)));
    layer4_outputs(1199) <= not(layer3_outputs(891)) or (layer3_outputs(2019));
    layer4_outputs(1200) <= layer3_outputs(1483);
    layer4_outputs(1201) <= not(layer3_outputs(1406));
    layer4_outputs(1202) <= not((layer3_outputs(1652)) or (layer3_outputs(1082)));
    layer4_outputs(1203) <= not(layer3_outputs(998));
    layer4_outputs(1204) <= not(layer3_outputs(438));
    layer4_outputs(1205) <= not(layer3_outputs(1223));
    layer4_outputs(1206) <= layer3_outputs(868);
    layer4_outputs(1207) <= (layer3_outputs(1069)) and (layer3_outputs(263));
    layer4_outputs(1208) <= (layer3_outputs(2343)) or (layer3_outputs(2182));
    layer4_outputs(1209) <= (layer3_outputs(399)) and (layer3_outputs(1214));
    layer4_outputs(1210) <= layer3_outputs(1860);
    layer4_outputs(1211) <= not((layer3_outputs(1380)) xor (layer3_outputs(2168)));
    layer4_outputs(1212) <= layer3_outputs(2331);
    layer4_outputs(1213) <= not(layer3_outputs(1745));
    layer4_outputs(1214) <= (layer3_outputs(16)) and not (layer3_outputs(1993));
    layer4_outputs(1215) <= not(layer3_outputs(792));
    layer4_outputs(1216) <= not((layer3_outputs(1806)) or (layer3_outputs(120)));
    layer4_outputs(1217) <= '1';
    layer4_outputs(1218) <= not(layer3_outputs(707));
    layer4_outputs(1219) <= not(layer3_outputs(498));
    layer4_outputs(1220) <= not(layer3_outputs(1833));
    layer4_outputs(1221) <= not(layer3_outputs(1408));
    layer4_outputs(1222) <= not(layer3_outputs(753));
    layer4_outputs(1223) <= not((layer3_outputs(2516)) or (layer3_outputs(553)));
    layer4_outputs(1224) <= (layer3_outputs(383)) and (layer3_outputs(1424));
    layer4_outputs(1225) <= not((layer3_outputs(1564)) and (layer3_outputs(2314)));
    layer4_outputs(1226) <= (layer3_outputs(51)) and (layer3_outputs(1243));
    layer4_outputs(1227) <= (layer3_outputs(729)) and (layer3_outputs(1022));
    layer4_outputs(1228) <= (layer3_outputs(448)) and not (layer3_outputs(1818));
    layer4_outputs(1229) <= (layer3_outputs(222)) and not (layer3_outputs(848));
    layer4_outputs(1230) <= not(layer3_outputs(2053));
    layer4_outputs(1231) <= not(layer3_outputs(1913));
    layer4_outputs(1232) <= layer3_outputs(1344);
    layer4_outputs(1233) <= not(layer3_outputs(2097));
    layer4_outputs(1234) <= not(layer3_outputs(1317));
    layer4_outputs(1235) <= '0';
    layer4_outputs(1236) <= (layer3_outputs(42)) and not (layer3_outputs(76));
    layer4_outputs(1237) <= not(layer3_outputs(2109)) or (layer3_outputs(463));
    layer4_outputs(1238) <= not(layer3_outputs(1049));
    layer4_outputs(1239) <= not((layer3_outputs(1914)) xor (layer3_outputs(18)));
    layer4_outputs(1240) <= (layer3_outputs(315)) and not (layer3_outputs(1601));
    layer4_outputs(1241) <= (layer3_outputs(1464)) and not (layer3_outputs(323));
    layer4_outputs(1242) <= (layer3_outputs(1749)) and not (layer3_outputs(955));
    layer4_outputs(1243) <= layer3_outputs(1068);
    layer4_outputs(1244) <= not(layer3_outputs(1766)) or (layer3_outputs(1323));
    layer4_outputs(1245) <= layer3_outputs(2404);
    layer4_outputs(1246) <= '0';
    layer4_outputs(1247) <= not(layer3_outputs(1098)) or (layer3_outputs(351));
    layer4_outputs(1248) <= '0';
    layer4_outputs(1249) <= (layer3_outputs(2249)) and not (layer3_outputs(2542));
    layer4_outputs(1250) <= not((layer3_outputs(1565)) or (layer3_outputs(1667)));
    layer4_outputs(1251) <= (layer3_outputs(73)) and not (layer3_outputs(1387));
    layer4_outputs(1252) <= layer3_outputs(1766);
    layer4_outputs(1253) <= (layer3_outputs(2201)) and not (layer3_outputs(54));
    layer4_outputs(1254) <= (layer3_outputs(620)) or (layer3_outputs(1977));
    layer4_outputs(1255) <= (layer3_outputs(338)) and not (layer3_outputs(154));
    layer4_outputs(1256) <= not(layer3_outputs(1861));
    layer4_outputs(1257) <= not(layer3_outputs(924)) or (layer3_outputs(2356));
    layer4_outputs(1258) <= not(layer3_outputs(961));
    layer4_outputs(1259) <= not(layer3_outputs(2203));
    layer4_outputs(1260) <= not(layer3_outputs(849)) or (layer3_outputs(1549));
    layer4_outputs(1261) <= not((layer3_outputs(732)) xor (layer3_outputs(669)));
    layer4_outputs(1262) <= layer3_outputs(309);
    layer4_outputs(1263) <= not(layer3_outputs(2048));
    layer4_outputs(1264) <= (layer3_outputs(2385)) and (layer3_outputs(308));
    layer4_outputs(1265) <= not(layer3_outputs(935));
    layer4_outputs(1266) <= (layer3_outputs(1899)) or (layer3_outputs(773));
    layer4_outputs(1267) <= (layer3_outputs(1794)) and not (layer3_outputs(2002));
    layer4_outputs(1268) <= (layer3_outputs(2259)) and not (layer3_outputs(561));
    layer4_outputs(1269) <= '0';
    layer4_outputs(1270) <= not(layer3_outputs(823));
    layer4_outputs(1271) <= (layer3_outputs(1396)) xor (layer3_outputs(1700));
    layer4_outputs(1272) <= (layer3_outputs(1276)) and (layer3_outputs(1276));
    layer4_outputs(1273) <= (layer3_outputs(606)) and not (layer3_outputs(900));
    layer4_outputs(1274) <= layer3_outputs(11);
    layer4_outputs(1275) <= (layer3_outputs(1961)) or (layer3_outputs(2308));
    layer4_outputs(1276) <= (layer3_outputs(1627)) and (layer3_outputs(286));
    layer4_outputs(1277) <= layer3_outputs(2457);
    layer4_outputs(1278) <= (layer3_outputs(214)) and (layer3_outputs(1884));
    layer4_outputs(1279) <= not(layer3_outputs(673)) or (layer3_outputs(336));
    layer4_outputs(1280) <= '1';
    layer4_outputs(1281) <= not(layer3_outputs(2008)) or (layer3_outputs(1650));
    layer4_outputs(1282) <= not((layer3_outputs(649)) xor (layer3_outputs(676)));
    layer4_outputs(1283) <= (layer3_outputs(490)) and not (layer3_outputs(1642));
    layer4_outputs(1284) <= layer3_outputs(1003);
    layer4_outputs(1285) <= '1';
    layer4_outputs(1286) <= '0';
    layer4_outputs(1287) <= (layer3_outputs(1395)) and not (layer3_outputs(462));
    layer4_outputs(1288) <= (layer3_outputs(1667)) or (layer3_outputs(751));
    layer4_outputs(1289) <= not((layer3_outputs(1248)) and (layer3_outputs(2305)));
    layer4_outputs(1290) <= not((layer3_outputs(1269)) and (layer3_outputs(63)));
    layer4_outputs(1291) <= layer3_outputs(814);
    layer4_outputs(1292) <= layer3_outputs(2024);
    layer4_outputs(1293) <= '0';
    layer4_outputs(1294) <= '1';
    layer4_outputs(1295) <= not(layer3_outputs(897)) or (layer3_outputs(1731));
    layer4_outputs(1296) <= layer3_outputs(1859);
    layer4_outputs(1297) <= not(layer3_outputs(314)) or (layer3_outputs(1098));
    layer4_outputs(1298) <= layer3_outputs(455);
    layer4_outputs(1299) <= not(layer3_outputs(2026));
    layer4_outputs(1300) <= not(layer3_outputs(1875)) or (layer3_outputs(228));
    layer4_outputs(1301) <= layer3_outputs(2549);
    layer4_outputs(1302) <= layer3_outputs(1897);
    layer4_outputs(1303) <= not((layer3_outputs(2373)) xor (layer3_outputs(2290)));
    layer4_outputs(1304) <= not(layer3_outputs(2468)) or (layer3_outputs(2338));
    layer4_outputs(1305) <= (layer3_outputs(1054)) xor (layer3_outputs(2463));
    layer4_outputs(1306) <= not(layer3_outputs(474));
    layer4_outputs(1307) <= (layer3_outputs(305)) and (layer3_outputs(1997));
    layer4_outputs(1308) <= layer3_outputs(1728);
    layer4_outputs(1309) <= not(layer3_outputs(1482));
    layer4_outputs(1310) <= layer3_outputs(1508);
    layer4_outputs(1311) <= layer3_outputs(1273);
    layer4_outputs(1312) <= not(layer3_outputs(2479));
    layer4_outputs(1313) <= layer3_outputs(1385);
    layer4_outputs(1314) <= layer3_outputs(169);
    layer4_outputs(1315) <= not(layer3_outputs(1100)) or (layer3_outputs(2444));
    layer4_outputs(1316) <= not((layer3_outputs(699)) or (layer3_outputs(2268)));
    layer4_outputs(1317) <= (layer3_outputs(1511)) or (layer3_outputs(2229));
    layer4_outputs(1318) <= not((layer3_outputs(2275)) or (layer3_outputs(1510)));
    layer4_outputs(1319) <= not(layer3_outputs(401));
    layer4_outputs(1320) <= (layer3_outputs(452)) and (layer3_outputs(1775));
    layer4_outputs(1321) <= not((layer3_outputs(486)) or (layer3_outputs(1453)));
    layer4_outputs(1322) <= (layer3_outputs(1232)) or (layer3_outputs(1792));
    layer4_outputs(1323) <= layer3_outputs(1786);
    layer4_outputs(1324) <= layer3_outputs(466);
    layer4_outputs(1325) <= '0';
    layer4_outputs(1326) <= (layer3_outputs(948)) and not (layer3_outputs(775));
    layer4_outputs(1327) <= layer3_outputs(177);
    layer4_outputs(1328) <= '0';
    layer4_outputs(1329) <= (layer3_outputs(1102)) and not (layer3_outputs(461));
    layer4_outputs(1330) <= not(layer3_outputs(1328));
    layer4_outputs(1331) <= layer3_outputs(2058);
    layer4_outputs(1332) <= not(layer3_outputs(205)) or (layer3_outputs(1015));
    layer4_outputs(1333) <= '1';
    layer4_outputs(1334) <= not(layer3_outputs(2271));
    layer4_outputs(1335) <= not(layer3_outputs(1886));
    layer4_outputs(1336) <= not(layer3_outputs(236));
    layer4_outputs(1337) <= layer3_outputs(568);
    layer4_outputs(1338) <= not((layer3_outputs(623)) and (layer3_outputs(2070)));
    layer4_outputs(1339) <= not(layer3_outputs(697)) or (layer3_outputs(1561));
    layer4_outputs(1340) <= layer3_outputs(333);
    layer4_outputs(1341) <= not(layer3_outputs(967));
    layer4_outputs(1342) <= not(layer3_outputs(873)) or (layer3_outputs(211));
    layer4_outputs(1343) <= not(layer3_outputs(2513));
    layer4_outputs(1344) <= not((layer3_outputs(2092)) or (layer3_outputs(2409)));
    layer4_outputs(1345) <= not(layer3_outputs(2212));
    layer4_outputs(1346) <= (layer3_outputs(9)) and not (layer3_outputs(2323));
    layer4_outputs(1347) <= (layer3_outputs(793)) xor (layer3_outputs(1899));
    layer4_outputs(1348) <= layer3_outputs(210);
    layer4_outputs(1349) <= '1';
    layer4_outputs(1350) <= '0';
    layer4_outputs(1351) <= layer3_outputs(1497);
    layer4_outputs(1352) <= not(layer3_outputs(554)) or (layer3_outputs(890));
    layer4_outputs(1353) <= not(layer3_outputs(1218)) or (layer3_outputs(1932));
    layer4_outputs(1354) <= (layer3_outputs(2392)) and not (layer3_outputs(865));
    layer4_outputs(1355) <= layer3_outputs(146);
    layer4_outputs(1356) <= not((layer3_outputs(598)) and (layer3_outputs(129)));
    layer4_outputs(1357) <= not(layer3_outputs(1359));
    layer4_outputs(1358) <= layer3_outputs(2537);
    layer4_outputs(1359) <= not(layer3_outputs(1238));
    layer4_outputs(1360) <= (layer3_outputs(2395)) and not (layer3_outputs(1855));
    layer4_outputs(1361) <= (layer3_outputs(441)) and not (layer3_outputs(1237));
    layer4_outputs(1362) <= (layer3_outputs(1391)) and not (layer3_outputs(1509));
    layer4_outputs(1363) <= not(layer3_outputs(667));
    layer4_outputs(1364) <= not((layer3_outputs(326)) or (layer3_outputs(1563)));
    layer4_outputs(1365) <= (layer3_outputs(1378)) and not (layer3_outputs(423));
    layer4_outputs(1366) <= not(layer3_outputs(2213));
    layer4_outputs(1367) <= layer3_outputs(1551);
    layer4_outputs(1368) <= not(layer3_outputs(1751)) or (layer3_outputs(2220));
    layer4_outputs(1369) <= '1';
    layer4_outputs(1370) <= not((layer3_outputs(2102)) or (layer3_outputs(2026)));
    layer4_outputs(1371) <= not((layer3_outputs(16)) or (layer3_outputs(1326)));
    layer4_outputs(1372) <= layer3_outputs(1833);
    layer4_outputs(1373) <= not(layer3_outputs(1628));
    layer4_outputs(1374) <= not(layer3_outputs(237));
    layer4_outputs(1375) <= not((layer3_outputs(1537)) or (layer3_outputs(1613)));
    layer4_outputs(1376) <= layer3_outputs(342);
    layer4_outputs(1377) <= not((layer3_outputs(2410)) and (layer3_outputs(1175)));
    layer4_outputs(1378) <= '1';
    layer4_outputs(1379) <= (layer3_outputs(2311)) or (layer3_outputs(324));
    layer4_outputs(1380) <= not((layer3_outputs(1601)) xor (layer3_outputs(535)));
    layer4_outputs(1381) <= not(layer3_outputs(356));
    layer4_outputs(1382) <= not((layer3_outputs(2286)) or (layer3_outputs(1739)));
    layer4_outputs(1383) <= (layer3_outputs(597)) and not (layer3_outputs(1513));
    layer4_outputs(1384) <= not(layer3_outputs(388));
    layer4_outputs(1385) <= not((layer3_outputs(1795)) or (layer3_outputs(142)));
    layer4_outputs(1386) <= not(layer3_outputs(443));
    layer4_outputs(1387) <= '0';
    layer4_outputs(1388) <= not(layer3_outputs(552));
    layer4_outputs(1389) <= '1';
    layer4_outputs(1390) <= (layer3_outputs(1442)) and (layer3_outputs(1205));
    layer4_outputs(1391) <= layer3_outputs(2386);
    layer4_outputs(1392) <= not(layer3_outputs(1449));
    layer4_outputs(1393) <= layer3_outputs(1199);
    layer4_outputs(1394) <= not((layer3_outputs(392)) and (layer3_outputs(1321)));
    layer4_outputs(1395) <= (layer3_outputs(1709)) and not (layer3_outputs(721));
    layer4_outputs(1396) <= (layer3_outputs(2078)) and (layer3_outputs(1637));
    layer4_outputs(1397) <= (layer3_outputs(2077)) or (layer3_outputs(674));
    layer4_outputs(1398) <= not(layer3_outputs(542)) or (layer3_outputs(1781));
    layer4_outputs(1399) <= layer3_outputs(2063);
    layer4_outputs(1400) <= layer3_outputs(932);
    layer4_outputs(1401) <= not(layer3_outputs(2240)) or (layer3_outputs(2252));
    layer4_outputs(1402) <= layer3_outputs(1753);
    layer4_outputs(1403) <= not(layer3_outputs(225));
    layer4_outputs(1404) <= (layer3_outputs(2170)) and (layer3_outputs(260));
    layer4_outputs(1405) <= (layer3_outputs(1530)) and not (layer3_outputs(2046));
    layer4_outputs(1406) <= (layer3_outputs(560)) and (layer3_outputs(232));
    layer4_outputs(1407) <= not((layer3_outputs(2386)) or (layer3_outputs(2193)));
    layer4_outputs(1408) <= (layer3_outputs(726)) and (layer3_outputs(1779));
    layer4_outputs(1409) <= not(layer3_outputs(531));
    layer4_outputs(1410) <= '1';
    layer4_outputs(1411) <= layer3_outputs(1335);
    layer4_outputs(1412) <= (layer3_outputs(1240)) and (layer3_outputs(2287));
    layer4_outputs(1413) <= layer3_outputs(715);
    layer4_outputs(1414) <= not(layer3_outputs(1345)) or (layer3_outputs(958));
    layer4_outputs(1415) <= layer3_outputs(2519);
    layer4_outputs(1416) <= layer3_outputs(378);
    layer4_outputs(1417) <= not((layer3_outputs(1261)) or (layer3_outputs(204)));
    layer4_outputs(1418) <= layer3_outputs(1340);
    layer4_outputs(1419) <= '0';
    layer4_outputs(1420) <= not(layer3_outputs(1311));
    layer4_outputs(1421) <= not(layer3_outputs(2315)) or (layer3_outputs(267));
    layer4_outputs(1422) <= (layer3_outputs(1719)) and not (layer3_outputs(469));
    layer4_outputs(1423) <= (layer3_outputs(563)) and not (layer3_outputs(1410));
    layer4_outputs(1424) <= not((layer3_outputs(2368)) xor (layer3_outputs(2404)));
    layer4_outputs(1425) <= not(layer3_outputs(253));
    layer4_outputs(1426) <= '1';
    layer4_outputs(1427) <= not((layer3_outputs(2304)) or (layer3_outputs(511)));
    layer4_outputs(1428) <= (layer3_outputs(1103)) and (layer3_outputs(1515));
    layer4_outputs(1429) <= not((layer3_outputs(1384)) and (layer3_outputs(1041)));
    layer4_outputs(1430) <= (layer3_outputs(2099)) or (layer3_outputs(987));
    layer4_outputs(1431) <= not(layer3_outputs(1457));
    layer4_outputs(1432) <= not(layer3_outputs(555));
    layer4_outputs(1433) <= not((layer3_outputs(2552)) and (layer3_outputs(117)));
    layer4_outputs(1434) <= layer3_outputs(837);
    layer4_outputs(1435) <= layer3_outputs(1704);
    layer4_outputs(1436) <= layer3_outputs(144);
    layer4_outputs(1437) <= '1';
    layer4_outputs(1438) <= (layer3_outputs(1244)) or (layer3_outputs(1984));
    layer4_outputs(1439) <= '0';
    layer4_outputs(1440) <= '0';
    layer4_outputs(1441) <= not(layer3_outputs(1592));
    layer4_outputs(1442) <= layer3_outputs(931);
    layer4_outputs(1443) <= '1';
    layer4_outputs(1444) <= layer3_outputs(996);
    layer4_outputs(1445) <= (layer3_outputs(538)) xor (layer3_outputs(596));
    layer4_outputs(1446) <= (layer3_outputs(152)) and (layer3_outputs(2387));
    layer4_outputs(1447) <= (layer3_outputs(121)) and not (layer3_outputs(158));
    layer4_outputs(1448) <= (layer3_outputs(598)) and not (layer3_outputs(1865));
    layer4_outputs(1449) <= (layer3_outputs(189)) and not (layer3_outputs(2327));
    layer4_outputs(1450) <= (layer3_outputs(2118)) and not (layer3_outputs(285));
    layer4_outputs(1451) <= layer3_outputs(1618);
    layer4_outputs(1452) <= layer3_outputs(544);
    layer4_outputs(1453) <= not(layer3_outputs(1274)) or (layer3_outputs(99));
    layer4_outputs(1454) <= not(layer3_outputs(344)) or (layer3_outputs(972));
    layer4_outputs(1455) <= not(layer3_outputs(123)) or (layer3_outputs(2136));
    layer4_outputs(1456) <= (layer3_outputs(331)) and not (layer3_outputs(800));
    layer4_outputs(1457) <= not(layer3_outputs(2074));
    layer4_outputs(1458) <= not(layer3_outputs(2192));
    layer4_outputs(1459) <= (layer3_outputs(1107)) or (layer3_outputs(1917));
    layer4_outputs(1460) <= not(layer3_outputs(195));
    layer4_outputs(1461) <= layer3_outputs(2028);
    layer4_outputs(1462) <= (layer3_outputs(2062)) or (layer3_outputs(2525));
    layer4_outputs(1463) <= not(layer3_outputs(1282)) or (layer3_outputs(799));
    layer4_outputs(1464) <= layer3_outputs(1460);
    layer4_outputs(1465) <= layer3_outputs(2179);
    layer4_outputs(1466) <= layer3_outputs(2362);
    layer4_outputs(1467) <= (layer3_outputs(1393)) or (layer3_outputs(812));
    layer4_outputs(1468) <= (layer3_outputs(2094)) and not (layer3_outputs(2253));
    layer4_outputs(1469) <= (layer3_outputs(1638)) or (layer3_outputs(1226));
    layer4_outputs(1470) <= not(layer3_outputs(2481));
    layer4_outputs(1471) <= (layer3_outputs(187)) and not (layer3_outputs(241));
    layer4_outputs(1472) <= layer3_outputs(2014);
    layer4_outputs(1473) <= '0';
    layer4_outputs(1474) <= (layer3_outputs(534)) and not (layer3_outputs(748));
    layer4_outputs(1475) <= layer3_outputs(638);
    layer4_outputs(1476) <= (layer3_outputs(2200)) and not (layer3_outputs(1023));
    layer4_outputs(1477) <= layer3_outputs(1895);
    layer4_outputs(1478) <= (layer3_outputs(1451)) and (layer3_outputs(1377));
    layer4_outputs(1479) <= layer3_outputs(1893);
    layer4_outputs(1480) <= not(layer3_outputs(701)) or (layer3_outputs(539));
    layer4_outputs(1481) <= '0';
    layer4_outputs(1482) <= (layer3_outputs(982)) xor (layer3_outputs(680));
    layer4_outputs(1483) <= (layer3_outputs(831)) and (layer3_outputs(429));
    layer4_outputs(1484) <= not((layer3_outputs(143)) or (layer3_outputs(1829)));
    layer4_outputs(1485) <= not(layer3_outputs(2521)) or (layer3_outputs(1182));
    layer4_outputs(1486) <= '0';
    layer4_outputs(1487) <= (layer3_outputs(1465)) and (layer3_outputs(489));
    layer4_outputs(1488) <= layer3_outputs(2512);
    layer4_outputs(1489) <= not(layer3_outputs(740));
    layer4_outputs(1490) <= not(layer3_outputs(2514));
    layer4_outputs(1491) <= '0';
    layer4_outputs(1492) <= '0';
    layer4_outputs(1493) <= (layer3_outputs(1876)) or (layer3_outputs(2378));
    layer4_outputs(1494) <= not(layer3_outputs(270));
    layer4_outputs(1495) <= (layer3_outputs(713)) and not (layer3_outputs(359));
    layer4_outputs(1496) <= not(layer3_outputs(99));
    layer4_outputs(1497) <= (layer3_outputs(1734)) xor (layer3_outputs(291));
    layer4_outputs(1498) <= (layer3_outputs(1187)) and (layer3_outputs(1072));
    layer4_outputs(1499) <= '1';
    layer4_outputs(1500) <= (layer3_outputs(397)) and not (layer3_outputs(250));
    layer4_outputs(1501) <= (layer3_outputs(1609)) and (layer3_outputs(931));
    layer4_outputs(1502) <= (layer3_outputs(1458)) or (layer3_outputs(778));
    layer4_outputs(1503) <= not((layer3_outputs(2066)) or (layer3_outputs(1597)));
    layer4_outputs(1504) <= not((layer3_outputs(347)) or (layer3_outputs(2160)));
    layer4_outputs(1505) <= not(layer3_outputs(1455));
    layer4_outputs(1506) <= layer3_outputs(1436);
    layer4_outputs(1507) <= (layer3_outputs(1779)) and not (layer3_outputs(446));
    layer4_outputs(1508) <= not(layer3_outputs(1134)) or (layer3_outputs(1023));
    layer4_outputs(1509) <= (layer3_outputs(1972)) and not (layer3_outputs(2426));
    layer4_outputs(1510) <= (layer3_outputs(192)) or (layer3_outputs(766));
    layer4_outputs(1511) <= '0';
    layer4_outputs(1512) <= '0';
    layer4_outputs(1513) <= not(layer3_outputs(1221)) or (layer3_outputs(600));
    layer4_outputs(1514) <= not((layer3_outputs(2508)) or (layer3_outputs(21)));
    layer4_outputs(1515) <= (layer3_outputs(2108)) and (layer3_outputs(1008));
    layer4_outputs(1516) <= '0';
    layer4_outputs(1517) <= (layer3_outputs(1372)) and not (layer3_outputs(705));
    layer4_outputs(1518) <= (layer3_outputs(2265)) and (layer3_outputs(574));
    layer4_outputs(1519) <= not(layer3_outputs(222)) or (layer3_outputs(1692));
    layer4_outputs(1520) <= (layer3_outputs(874)) xor (layer3_outputs(2358));
    layer4_outputs(1521) <= layer3_outputs(212);
    layer4_outputs(1522) <= not(layer3_outputs(511));
    layer4_outputs(1523) <= (layer3_outputs(2067)) and not (layer3_outputs(74));
    layer4_outputs(1524) <= (layer3_outputs(630)) or (layer3_outputs(163));
    layer4_outputs(1525) <= '1';
    layer4_outputs(1526) <= not(layer3_outputs(2176)) or (layer3_outputs(325));
    layer4_outputs(1527) <= '0';
    layer4_outputs(1528) <= (layer3_outputs(502)) and not (layer3_outputs(399));
    layer4_outputs(1529) <= not(layer3_outputs(942));
    layer4_outputs(1530) <= (layer3_outputs(952)) and (layer3_outputs(925));
    layer4_outputs(1531) <= (layer3_outputs(186)) and (layer3_outputs(1270));
    layer4_outputs(1532) <= not(layer3_outputs(449));
    layer4_outputs(1533) <= not(layer3_outputs(1184));
    layer4_outputs(1534) <= not(layer3_outputs(2223)) or (layer3_outputs(95));
    layer4_outputs(1535) <= not(layer3_outputs(1527)) or (layer3_outputs(1374));
    layer4_outputs(1536) <= not((layer3_outputs(1121)) and (layer3_outputs(1157)));
    layer4_outputs(1537) <= not(layer3_outputs(2134));
    layer4_outputs(1538) <= '0';
    layer4_outputs(1539) <= not((layer3_outputs(2125)) or (layer3_outputs(2245)));
    layer4_outputs(1540) <= layer3_outputs(2254);
    layer4_outputs(1541) <= not((layer3_outputs(1668)) or (layer3_outputs(2554)));
    layer4_outputs(1542) <= layer3_outputs(1199);
    layer4_outputs(1543) <= not(layer3_outputs(774));
    layer4_outputs(1544) <= '0';
    layer4_outputs(1545) <= not(layer3_outputs(905));
    layer4_outputs(1546) <= not(layer3_outputs(635));
    layer4_outputs(1547) <= not(layer3_outputs(374));
    layer4_outputs(1548) <= not((layer3_outputs(1068)) and (layer3_outputs(1722)));
    layer4_outputs(1549) <= not(layer3_outputs(1118));
    layer4_outputs(1550) <= not((layer3_outputs(2060)) xor (layer3_outputs(1039)));
    layer4_outputs(1551) <= '0';
    layer4_outputs(1552) <= not((layer3_outputs(2042)) and (layer3_outputs(2418)));
    layer4_outputs(1553) <= not(layer3_outputs(1920)) or (layer3_outputs(1064));
    layer4_outputs(1554) <= not((layer3_outputs(680)) or (layer3_outputs(1355)));
    layer4_outputs(1555) <= layer3_outputs(1912);
    layer4_outputs(1556) <= not(layer3_outputs(467)) or (layer3_outputs(1054));
    layer4_outputs(1557) <= '1';
    layer4_outputs(1558) <= not(layer3_outputs(2209));
    layer4_outputs(1559) <= not(layer3_outputs(2199)) or (layer3_outputs(1737));
    layer4_outputs(1560) <= (layer3_outputs(1178)) xor (layer3_outputs(1522));
    layer4_outputs(1561) <= (layer3_outputs(2346)) or (layer3_outputs(927));
    layer4_outputs(1562) <= (layer3_outputs(1102)) and (layer3_outputs(419));
    layer4_outputs(1563) <= (layer3_outputs(1100)) and not (layer3_outputs(1970));
    layer4_outputs(1564) <= not(layer3_outputs(188)) or (layer3_outputs(1017));
    layer4_outputs(1565) <= layer3_outputs(1128);
    layer4_outputs(1566) <= (layer3_outputs(914)) or (layer3_outputs(199));
    layer4_outputs(1567) <= not(layer3_outputs(823));
    layer4_outputs(1568) <= not((layer3_outputs(502)) xor (layer3_outputs(725)));
    layer4_outputs(1569) <= layer3_outputs(841);
    layer4_outputs(1570) <= (layer3_outputs(2473)) or (layer3_outputs(546));
    layer4_outputs(1571) <= layer3_outputs(2449);
    layer4_outputs(1572) <= (layer3_outputs(1540)) or (layer3_outputs(1245));
    layer4_outputs(1573) <= not((layer3_outputs(1143)) or (layer3_outputs(1583)));
    layer4_outputs(1574) <= layer3_outputs(735);
    layer4_outputs(1575) <= not((layer3_outputs(1595)) and (layer3_outputs(1536)));
    layer4_outputs(1576) <= not((layer3_outputs(1373)) or (layer3_outputs(794)));
    layer4_outputs(1577) <= not(layer3_outputs(2496)) or (layer3_outputs(2556));
    layer4_outputs(1578) <= (layer3_outputs(227)) and not (layer3_outputs(740));
    layer4_outputs(1579) <= not((layer3_outputs(1741)) or (layer3_outputs(1015)));
    layer4_outputs(1580) <= not(layer3_outputs(785));
    layer4_outputs(1581) <= layer3_outputs(181);
    layer4_outputs(1582) <= not(layer3_outputs(2375)) or (layer3_outputs(2072));
    layer4_outputs(1583) <= not((layer3_outputs(339)) or (layer3_outputs(945)));
    layer4_outputs(1584) <= not(layer3_outputs(2372));
    layer4_outputs(1585) <= layer3_outputs(437);
    layer4_outputs(1586) <= not(layer3_outputs(1006)) or (layer3_outputs(1296));
    layer4_outputs(1587) <= not((layer3_outputs(776)) and (layer3_outputs(1861)));
    layer4_outputs(1588) <= '1';
    layer4_outputs(1589) <= not((layer3_outputs(2271)) xor (layer3_outputs(941)));
    layer4_outputs(1590) <= (layer3_outputs(2064)) and (layer3_outputs(1259));
    layer4_outputs(1591) <= (layer3_outputs(1014)) or (layer3_outputs(926));
    layer4_outputs(1592) <= not(layer3_outputs(750));
    layer4_outputs(1593) <= not(layer3_outputs(1585));
    layer4_outputs(1594) <= (layer3_outputs(696)) or (layer3_outputs(1140));
    layer4_outputs(1595) <= layer3_outputs(1607);
    layer4_outputs(1596) <= layer3_outputs(1622);
    layer4_outputs(1597) <= layer3_outputs(161);
    layer4_outputs(1598) <= '0';
    layer4_outputs(1599) <= not(layer3_outputs(813));
    layer4_outputs(1600) <= layer3_outputs(2457);
    layer4_outputs(1601) <= layer3_outputs(2510);
    layer4_outputs(1602) <= not(layer3_outputs(1687));
    layer4_outputs(1603) <= (layer3_outputs(2144)) xor (layer3_outputs(933));
    layer4_outputs(1604) <= not(layer3_outputs(2294));
    layer4_outputs(1605) <= layer3_outputs(81);
    layer4_outputs(1606) <= (layer3_outputs(1804)) and not (layer3_outputs(2123));
    layer4_outputs(1607) <= layer3_outputs(251);
    layer4_outputs(1608) <= layer3_outputs(1232);
    layer4_outputs(1609) <= layer3_outputs(2152);
    layer4_outputs(1610) <= '0';
    layer4_outputs(1611) <= (layer3_outputs(79)) xor (layer3_outputs(2207));
    layer4_outputs(1612) <= not(layer3_outputs(477)) or (layer3_outputs(2266));
    layer4_outputs(1613) <= '0';
    layer4_outputs(1614) <= layer3_outputs(145);
    layer4_outputs(1615) <= layer3_outputs(661);
    layer4_outputs(1616) <= layer3_outputs(1095);
    layer4_outputs(1617) <= (layer3_outputs(802)) and not (layer3_outputs(2177));
    layer4_outputs(1618) <= not(layer3_outputs(1639));
    layer4_outputs(1619) <= not(layer3_outputs(632));
    layer4_outputs(1620) <= not(layer3_outputs(1217));
    layer4_outputs(1621) <= layer3_outputs(2455);
    layer4_outputs(1622) <= '0';
    layer4_outputs(1623) <= not(layer3_outputs(1394));
    layer4_outputs(1624) <= not(layer3_outputs(2415));
    layer4_outputs(1625) <= not(layer3_outputs(2081)) or (layer3_outputs(679));
    layer4_outputs(1626) <= '1';
    layer4_outputs(1627) <= not(layer3_outputs(2265)) or (layer3_outputs(1452));
    layer4_outputs(1628) <= '1';
    layer4_outputs(1629) <= not(layer3_outputs(422));
    layer4_outputs(1630) <= layer3_outputs(454);
    layer4_outputs(1631) <= (layer3_outputs(1165)) and not (layer3_outputs(115));
    layer4_outputs(1632) <= not(layer3_outputs(1755));
    layer4_outputs(1633) <= not(layer3_outputs(2137));
    layer4_outputs(1634) <= '0';
    layer4_outputs(1635) <= not(layer3_outputs(1830)) or (layer3_outputs(2165));
    layer4_outputs(1636) <= (layer3_outputs(887)) and not (layer3_outputs(1783));
    layer4_outputs(1637) <= not(layer3_outputs(1530));
    layer4_outputs(1638) <= not(layer3_outputs(258));
    layer4_outputs(1639) <= '1';
    layer4_outputs(1640) <= (layer3_outputs(1901)) and not (layer3_outputs(2109));
    layer4_outputs(1641) <= '0';
    layer4_outputs(1642) <= not(layer3_outputs(1158)) or (layer3_outputs(1173));
    layer4_outputs(1643) <= not(layer3_outputs(2285));
    layer4_outputs(1644) <= (layer3_outputs(1122)) or (layer3_outputs(2507));
    layer4_outputs(1645) <= layer3_outputs(892);
    layer4_outputs(1646) <= not(layer3_outputs(2533)) or (layer3_outputs(2066));
    layer4_outputs(1647) <= not(layer3_outputs(242)) or (layer3_outputs(798));
    layer4_outputs(1648) <= not((layer3_outputs(1184)) and (layer3_outputs(1781)));
    layer4_outputs(1649) <= layer3_outputs(629);
    layer4_outputs(1650) <= not(layer3_outputs(1850)) or (layer3_outputs(1209));
    layer4_outputs(1651) <= not((layer3_outputs(366)) and (layer3_outputs(2481)));
    layer4_outputs(1652) <= layer3_outputs(2524);
    layer4_outputs(1653) <= not((layer3_outputs(1836)) and (layer3_outputs(1756)));
    layer4_outputs(1654) <= (layer3_outputs(821)) and (layer3_outputs(1790));
    layer4_outputs(1655) <= (layer3_outputs(2326)) and (layer3_outputs(1087));
    layer4_outputs(1656) <= '0';
    layer4_outputs(1657) <= (layer3_outputs(1167)) or (layer3_outputs(217));
    layer4_outputs(1658) <= layer3_outputs(2514);
    layer4_outputs(1659) <= not(layer3_outputs(1894)) or (layer3_outputs(2129));
    layer4_outputs(1660) <= not(layer3_outputs(121));
    layer4_outputs(1661) <= not(layer3_outputs(2081));
    layer4_outputs(1662) <= not(layer3_outputs(999));
    layer4_outputs(1663) <= '1';
    layer4_outputs(1664) <= not(layer3_outputs(1756)) or (layer3_outputs(1696));
    layer4_outputs(1665) <= not(layer3_outputs(1021));
    layer4_outputs(1666) <= not((layer3_outputs(942)) or (layer3_outputs(104)));
    layer4_outputs(1667) <= not((layer3_outputs(2367)) and (layer3_outputs(385)));
    layer4_outputs(1668) <= not((layer3_outputs(2297)) or (layer3_outputs(2363)));
    layer4_outputs(1669) <= (layer3_outputs(938)) and not (layer3_outputs(506));
    layer4_outputs(1670) <= (layer3_outputs(1598)) and (layer3_outputs(1268));
    layer4_outputs(1671) <= layer3_outputs(2241);
    layer4_outputs(1672) <= not(layer3_outputs(381));
    layer4_outputs(1673) <= (layer3_outputs(1785)) or (layer3_outputs(363));
    layer4_outputs(1674) <= (layer3_outputs(1200)) and not (layer3_outputs(1417));
    layer4_outputs(1675) <= not(layer3_outputs(787)) or (layer3_outputs(365));
    layer4_outputs(1676) <= not(layer3_outputs(576));
    layer4_outputs(1677) <= (layer3_outputs(2140)) and not (layer3_outputs(410));
    layer4_outputs(1678) <= (layer3_outputs(111)) and (layer3_outputs(802));
    layer4_outputs(1679) <= (layer3_outputs(200)) or (layer3_outputs(415));
    layer4_outputs(1680) <= layer3_outputs(1336);
    layer4_outputs(1681) <= '1';
    layer4_outputs(1682) <= not(layer3_outputs(1604));
    layer4_outputs(1683) <= '1';
    layer4_outputs(1684) <= layer3_outputs(1580);
    layer4_outputs(1685) <= (layer3_outputs(2341)) or (layer3_outputs(2234));
    layer4_outputs(1686) <= not(layer3_outputs(2011));
    layer4_outputs(1687) <= not(layer3_outputs(861));
    layer4_outputs(1688) <= (layer3_outputs(1157)) and not (layer3_outputs(765));
    layer4_outputs(1689) <= (layer3_outputs(1548)) or (layer3_outputs(628));
    layer4_outputs(1690) <= layer3_outputs(915);
    layer4_outputs(1691) <= not(layer3_outputs(2541));
    layer4_outputs(1692) <= (layer3_outputs(1413)) xor (layer3_outputs(1088));
    layer4_outputs(1693) <= (layer3_outputs(2451)) or (layer3_outputs(1541));
    layer4_outputs(1694) <= (layer3_outputs(172)) or (layer3_outputs(1746));
    layer4_outputs(1695) <= (layer3_outputs(91)) and not (layer3_outputs(642));
    layer4_outputs(1696) <= layer3_outputs(444);
    layer4_outputs(1697) <= layer3_outputs(2416);
    layer4_outputs(1698) <= not(layer3_outputs(413));
    layer4_outputs(1699) <= (layer3_outputs(819)) xor (layer3_outputs(2157));
    layer4_outputs(1700) <= not(layer3_outputs(1723));
    layer4_outputs(1701) <= layer3_outputs(2445);
    layer4_outputs(1702) <= '0';
    layer4_outputs(1703) <= layer3_outputs(811);
    layer4_outputs(1704) <= layer3_outputs(2371);
    layer4_outputs(1705) <= not(layer3_outputs(101)) or (layer3_outputs(1281));
    layer4_outputs(1706) <= (layer3_outputs(2255)) or (layer3_outputs(1108));
    layer4_outputs(1707) <= not((layer3_outputs(1875)) and (layer3_outputs(1644)));
    layer4_outputs(1708) <= not(layer3_outputs(854));
    layer4_outputs(1709) <= not(layer3_outputs(2050));
    layer4_outputs(1710) <= '0';
    layer4_outputs(1711) <= not((layer3_outputs(1890)) and (layer3_outputs(322)));
    layer4_outputs(1712) <= not(layer3_outputs(2414));
    layer4_outputs(1713) <= layer3_outputs(2112);
    layer4_outputs(1714) <= not(layer3_outputs(925));
    layer4_outputs(1715) <= layer3_outputs(838);
    layer4_outputs(1716) <= (layer3_outputs(2470)) and (layer3_outputs(2383));
    layer4_outputs(1717) <= (layer3_outputs(492)) and not (layer3_outputs(1815));
    layer4_outputs(1718) <= '0';
    layer4_outputs(1719) <= '1';
    layer4_outputs(1720) <= not((layer3_outputs(848)) or (layer3_outputs(1845)));
    layer4_outputs(1721) <= not((layer3_outputs(1934)) xor (layer3_outputs(2011)));
    layer4_outputs(1722) <= layer3_outputs(1991);
    layer4_outputs(1723) <= not((layer3_outputs(1369)) or (layer3_outputs(1265)));
    layer4_outputs(1724) <= '1';
    layer4_outputs(1725) <= not(layer3_outputs(754));
    layer4_outputs(1726) <= (layer3_outputs(1910)) and not (layer3_outputs(2293));
    layer4_outputs(1727) <= layer3_outputs(233);
    layer4_outputs(1728) <= not(layer3_outputs(2335));
    layer4_outputs(1729) <= not(layer3_outputs(1119));
    layer4_outputs(1730) <= (layer3_outputs(2177)) or (layer3_outputs(1752));
    layer4_outputs(1731) <= (layer3_outputs(2347)) or (layer3_outputs(591));
    layer4_outputs(1732) <= not(layer3_outputs(1017));
    layer4_outputs(1733) <= (layer3_outputs(1574)) or (layer3_outputs(403));
    layer4_outputs(1734) <= not(layer3_outputs(1725));
    layer4_outputs(1735) <= layer3_outputs(2530);
    layer4_outputs(1736) <= (layer3_outputs(62)) and (layer3_outputs(2269));
    layer4_outputs(1737) <= not(layer3_outputs(854)) or (layer3_outputs(1643));
    layer4_outputs(1738) <= not(layer3_outputs(2183));
    layer4_outputs(1739) <= (layer3_outputs(587)) and not (layer3_outputs(1510));
    layer4_outputs(1740) <= (layer3_outputs(57)) and not (layer3_outputs(1365));
    layer4_outputs(1741) <= (layer3_outputs(851)) and (layer3_outputs(1849));
    layer4_outputs(1742) <= layer3_outputs(1979);
    layer4_outputs(1743) <= not(layer3_outputs(168)) or (layer3_outputs(1231));
    layer4_outputs(1744) <= not((layer3_outputs(2469)) and (layer3_outputs(1148)));
    layer4_outputs(1745) <= layer3_outputs(2377);
    layer4_outputs(1746) <= (layer3_outputs(481)) or (layer3_outputs(1748));
    layer4_outputs(1747) <= layer3_outputs(1508);
    layer4_outputs(1748) <= (layer3_outputs(901)) xor (layer3_outputs(1512));
    layer4_outputs(1749) <= '1';
    layer4_outputs(1750) <= layer3_outputs(1698);
    layer4_outputs(1751) <= layer3_outputs(29);
    layer4_outputs(1752) <= not(layer3_outputs(1868));
    layer4_outputs(1753) <= not(layer3_outputs(639)) or (layer3_outputs(2318));
    layer4_outputs(1754) <= not(layer3_outputs(679)) or (layer3_outputs(1517));
    layer4_outputs(1755) <= layer3_outputs(2266);
    layer4_outputs(1756) <= not(layer3_outputs(1491)) or (layer3_outputs(238));
    layer4_outputs(1757) <= (layer3_outputs(644)) or (layer3_outputs(2));
    layer4_outputs(1758) <= not(layer3_outputs(1719)) or (layer3_outputs(1825));
    layer4_outputs(1759) <= not(layer3_outputs(130)) or (layer3_outputs(325));
    layer4_outputs(1760) <= layer3_outputs(703);
    layer4_outputs(1761) <= not((layer3_outputs(2151)) or (layer3_outputs(1600)));
    layer4_outputs(1762) <= layer3_outputs(1309);
    layer4_outputs(1763) <= (layer3_outputs(845)) and not (layer3_outputs(1626));
    layer4_outputs(1764) <= (layer3_outputs(1573)) and (layer3_outputs(1720));
    layer4_outputs(1765) <= layer3_outputs(2237);
    layer4_outputs(1766) <= not(layer3_outputs(12)) or (layer3_outputs(1702));
    layer4_outputs(1767) <= (layer3_outputs(332)) and not (layer3_outputs(883));
    layer4_outputs(1768) <= layer3_outputs(820);
    layer4_outputs(1769) <= not(layer3_outputs(543)) or (layer3_outputs(1052));
    layer4_outputs(1770) <= not(layer3_outputs(1385));
    layer4_outputs(1771) <= layer3_outputs(2247);
    layer4_outputs(1772) <= (layer3_outputs(1933)) and not (layer3_outputs(2438));
    layer4_outputs(1773) <= layer3_outputs(274);
    layer4_outputs(1774) <= not((layer3_outputs(2456)) and (layer3_outputs(1468)));
    layer4_outputs(1775) <= (layer3_outputs(2328)) and not (layer3_outputs(1242));
    layer4_outputs(1776) <= layer3_outputs(2184);
    layer4_outputs(1777) <= layer3_outputs(126);
    layer4_outputs(1778) <= not(layer3_outputs(610)) or (layer3_outputs(78));
    layer4_outputs(1779) <= not(layer3_outputs(775));
    layer4_outputs(1780) <= (layer3_outputs(1616)) and not (layer3_outputs(299));
    layer4_outputs(1781) <= not(layer3_outputs(1469)) or (layer3_outputs(22));
    layer4_outputs(1782) <= (layer3_outputs(614)) and not (layer3_outputs(937));
    layer4_outputs(1783) <= layer3_outputs(1420);
    layer4_outputs(1784) <= '1';
    layer4_outputs(1785) <= not((layer3_outputs(500)) and (layer3_outputs(1051)));
    layer4_outputs(1786) <= not(layer3_outputs(1573)) or (layer3_outputs(529));
    layer4_outputs(1787) <= layer3_outputs(2250);
    layer4_outputs(1788) <= layer3_outputs(2163);
    layer4_outputs(1789) <= (layer3_outputs(2511)) xor (layer3_outputs(2114));
    layer4_outputs(1790) <= layer3_outputs(175);
    layer4_outputs(1791) <= not((layer3_outputs(1828)) or (layer3_outputs(48)));
    layer4_outputs(1792) <= (layer3_outputs(1131)) or (layer3_outputs(353));
    layer4_outputs(1793) <= (layer3_outputs(1164)) and (layer3_outputs(1862));
    layer4_outputs(1794) <= '0';
    layer4_outputs(1795) <= layer3_outputs(1365);
    layer4_outputs(1796) <= '1';
    layer4_outputs(1797) <= '1';
    layer4_outputs(1798) <= not(layer3_outputs(75)) or (layer3_outputs(2298));
    layer4_outputs(1799) <= not(layer3_outputs(1401));
    layer4_outputs(1800) <= not(layer3_outputs(1002));
    layer4_outputs(1801) <= not(layer3_outputs(2032));
    layer4_outputs(1802) <= not(layer3_outputs(1813));
    layer4_outputs(1803) <= '1';
    layer4_outputs(1804) <= not(layer3_outputs(1949));
    layer4_outputs(1805) <= layer3_outputs(3);
    layer4_outputs(1806) <= layer3_outputs(601);
    layer4_outputs(1807) <= not(layer3_outputs(744));
    layer4_outputs(1808) <= '0';
    layer4_outputs(1809) <= layer3_outputs(125);
    layer4_outputs(1810) <= (layer3_outputs(2471)) and not (layer3_outputs(1384));
    layer4_outputs(1811) <= layer3_outputs(807);
    layer4_outputs(1812) <= not((layer3_outputs(959)) or (layer3_outputs(306)));
    layer4_outputs(1813) <= (layer3_outputs(2495)) and not (layer3_outputs(269));
    layer4_outputs(1814) <= not(layer3_outputs(645));
    layer4_outputs(1815) <= not(layer3_outputs(1647));
    layer4_outputs(1816) <= not((layer3_outputs(1040)) and (layer3_outputs(247)));
    layer4_outputs(1817) <= (layer3_outputs(1743)) and (layer3_outputs(229));
    layer4_outputs(1818) <= (layer3_outputs(328)) and not (layer3_outputs(1408));
    layer4_outputs(1819) <= layer3_outputs(1755);
    layer4_outputs(1820) <= not((layer3_outputs(923)) or (layer3_outputs(415)));
    layer4_outputs(1821) <= (layer3_outputs(1441)) and (layer3_outputs(1600));
    layer4_outputs(1822) <= not(layer3_outputs(648)) or (layer3_outputs(124));
    layer4_outputs(1823) <= layer3_outputs(1254);
    layer4_outputs(1824) <= (layer3_outputs(2149)) and (layer3_outputs(715));
    layer4_outputs(1825) <= (layer3_outputs(1166)) or (layer3_outputs(766));
    layer4_outputs(1826) <= (layer3_outputs(2045)) and (layer3_outputs(75));
    layer4_outputs(1827) <= not(layer3_outputs(1281));
    layer4_outputs(1828) <= (layer3_outputs(80)) and (layer3_outputs(1139));
    layer4_outputs(1829) <= '1';
    layer4_outputs(1830) <= (layer3_outputs(1629)) and not (layer3_outputs(817));
    layer4_outputs(1831) <= not((layer3_outputs(1131)) and (layer3_outputs(1207)));
    layer4_outputs(1832) <= layer3_outputs(2007);
    layer4_outputs(1833) <= not((layer3_outputs(2217)) and (layer3_outputs(1572)));
    layer4_outputs(1834) <= not(layer3_outputs(783));
    layer4_outputs(1835) <= not(layer3_outputs(2289)) or (layer3_outputs(1596));
    layer4_outputs(1836) <= not(layer3_outputs(0));
    layer4_outputs(1837) <= layer3_outputs(727);
    layer4_outputs(1838) <= not(layer3_outputs(408)) or (layer3_outputs(964));
    layer4_outputs(1839) <= (layer3_outputs(1670)) and not (layer3_outputs(313));
    layer4_outputs(1840) <= not(layer3_outputs(1777)) or (layer3_outputs(1587));
    layer4_outputs(1841) <= (layer3_outputs(2165)) and (layer3_outputs(2048));
    layer4_outputs(1842) <= layer3_outputs(407);
    layer4_outputs(1843) <= not(layer3_outputs(2433)) or (layer3_outputs(1620));
    layer4_outputs(1844) <= '1';
    layer4_outputs(1845) <= layer3_outputs(784);
    layer4_outputs(1846) <= not(layer3_outputs(1438));
    layer4_outputs(1847) <= layer3_outputs(504);
    layer4_outputs(1848) <= layer3_outputs(1246);
    layer4_outputs(1849) <= not(layer3_outputs(976));
    layer4_outputs(1850) <= layer3_outputs(1326);
    layer4_outputs(1851) <= not((layer3_outputs(379)) and (layer3_outputs(590)));
    layer4_outputs(1852) <= not(layer3_outputs(467));
    layer4_outputs(1853) <= (layer3_outputs(1820)) and not (layer3_outputs(564));
    layer4_outputs(1854) <= not(layer3_outputs(909));
    layer4_outputs(1855) <= not(layer3_outputs(436));
    layer4_outputs(1856) <= not(layer3_outputs(618));
    layer4_outputs(1857) <= (layer3_outputs(2366)) and not (layer3_outputs(893));
    layer4_outputs(1858) <= layer3_outputs(2185);
    layer4_outputs(1859) <= not(layer3_outputs(355));
    layer4_outputs(1860) <= layer3_outputs(2370);
    layer4_outputs(1861) <= not((layer3_outputs(1329)) and (layer3_outputs(489)));
    layer4_outputs(1862) <= (layer3_outputs(2466)) and not (layer3_outputs(1834));
    layer4_outputs(1863) <= layer3_outputs(1697);
    layer4_outputs(1864) <= (layer3_outputs(2280)) and (layer3_outputs(805));
    layer4_outputs(1865) <= layer3_outputs(947);
    layer4_outputs(1866) <= not((layer3_outputs(558)) and (layer3_outputs(1096)));
    layer4_outputs(1867) <= not((layer3_outputs(738)) and (layer3_outputs(517)));
    layer4_outputs(1868) <= not(layer3_outputs(557));
    layer4_outputs(1869) <= layer3_outputs(747);
    layer4_outputs(1870) <= layer3_outputs(1443);
    layer4_outputs(1871) <= layer3_outputs(1900);
    layer4_outputs(1872) <= not(layer3_outputs(409)) or (layer3_outputs(1943));
    layer4_outputs(1873) <= (layer3_outputs(876)) and not (layer3_outputs(984));
    layer4_outputs(1874) <= not(layer3_outputs(1299));
    layer4_outputs(1875) <= not(layer3_outputs(824));
    layer4_outputs(1876) <= not(layer3_outputs(1569));
    layer4_outputs(1877) <= not((layer3_outputs(425)) or (layer3_outputs(1767)));
    layer4_outputs(1878) <= (layer3_outputs(1742)) and not (layer3_outputs(2188));
    layer4_outputs(1879) <= '0';
    layer4_outputs(1880) <= not(layer3_outputs(946));
    layer4_outputs(1881) <= not(layer3_outputs(2115)) or (layer3_outputs(915));
    layer4_outputs(1882) <= layer3_outputs(570);
    layer4_outputs(1883) <= (layer3_outputs(1057)) or (layer3_outputs(1996));
    layer4_outputs(1884) <= (layer3_outputs(1532)) and (layer3_outputs(1906));
    layer4_outputs(1885) <= not(layer3_outputs(274));
    layer4_outputs(1886) <= (layer3_outputs(902)) and not (layer3_outputs(944));
    layer4_outputs(1887) <= (layer3_outputs(53)) and (layer3_outputs(370));
    layer4_outputs(1888) <= not((layer3_outputs(1773)) or (layer3_outputs(702)));
    layer4_outputs(1889) <= layer3_outputs(1272);
    layer4_outputs(1890) <= not(layer3_outputs(1223)) or (layer3_outputs(376));
    layer4_outputs(1891) <= not((layer3_outputs(1129)) and (layer3_outputs(22)));
    layer4_outputs(1892) <= '0';
    layer4_outputs(1893) <= not(layer3_outputs(2108));
    layer4_outputs(1894) <= not(layer3_outputs(44));
    layer4_outputs(1895) <= (layer3_outputs(693)) and not (layer3_outputs(1697));
    layer4_outputs(1896) <= layer3_outputs(1723);
    layer4_outputs(1897) <= not((layer3_outputs(2303)) and (layer3_outputs(916)));
    layer4_outputs(1898) <= not(layer3_outputs(587)) or (layer3_outputs(1675));
    layer4_outputs(1899) <= (layer3_outputs(2172)) and not (layer3_outputs(1608));
    layer4_outputs(1900) <= not((layer3_outputs(2468)) and (layer3_outputs(1476)));
    layer4_outputs(1901) <= layer3_outputs(866);
    layer4_outputs(1902) <= not(layer3_outputs(151));
    layer4_outputs(1903) <= not(layer3_outputs(261));
    layer4_outputs(1904) <= layer3_outputs(818);
    layer4_outputs(1905) <= layer3_outputs(929);
    layer4_outputs(1906) <= layer3_outputs(2226);
    layer4_outputs(1907) <= not(layer3_outputs(972)) or (layer3_outputs(342));
    layer4_outputs(1908) <= (layer3_outputs(1206)) and not (layer3_outputs(1607));
    layer4_outputs(1909) <= (layer3_outputs(790)) and not (layer3_outputs(840));
    layer4_outputs(1910) <= layer3_outputs(851);
    layer4_outputs(1911) <= not(layer3_outputs(459));
    layer4_outputs(1912) <= not(layer3_outputs(1056));
    layer4_outputs(1913) <= layer3_outputs(550);
    layer4_outputs(1914) <= not((layer3_outputs(201)) and (layer3_outputs(137)));
    layer4_outputs(1915) <= not(layer3_outputs(1793)) or (layer3_outputs(1996));
    layer4_outputs(1916) <= layer3_outputs(1900);
    layer4_outputs(1917) <= not(layer3_outputs(191));
    layer4_outputs(1918) <= not(layer3_outputs(1603)) or (layer3_outputs(1193));
    layer4_outputs(1919) <= layer3_outputs(404);
    layer4_outputs(1920) <= not((layer3_outputs(1048)) and (layer3_outputs(1740)));
    layer4_outputs(1921) <= not((layer3_outputs(1590)) xor (layer3_outputs(2216)));
    layer4_outputs(1922) <= not((layer3_outputs(1803)) or (layer3_outputs(395)));
    layer4_outputs(1923) <= (layer3_outputs(1486)) and not (layer3_outputs(781));
    layer4_outputs(1924) <= not((layer3_outputs(260)) or (layer3_outputs(2388)));
    layer4_outputs(1925) <= not(layer3_outputs(647));
    layer4_outputs(1926) <= (layer3_outputs(551)) or (layer3_outputs(850));
    layer4_outputs(1927) <= not(layer3_outputs(501));
    layer4_outputs(1928) <= '1';
    layer4_outputs(1929) <= '1';
    layer4_outputs(1930) <= layer3_outputs(2111);
    layer4_outputs(1931) <= (layer3_outputs(472)) and not (layer3_outputs(1733));
    layer4_outputs(1932) <= not(layer3_outputs(2540));
    layer4_outputs(1933) <= (layer3_outputs(340)) and not (layer3_outputs(206));
    layer4_outputs(1934) <= (layer3_outputs(1085)) or (layer3_outputs(2125));
    layer4_outputs(1935) <= not(layer3_outputs(28));
    layer4_outputs(1936) <= not(layer3_outputs(793));
    layer4_outputs(1937) <= not(layer3_outputs(1413));
    layer4_outputs(1938) <= not((layer3_outputs(1908)) and (layer3_outputs(1435)));
    layer4_outputs(1939) <= layer3_outputs(1376);
    layer4_outputs(1940) <= (layer3_outputs(1950)) or (layer3_outputs(611));
    layer4_outputs(1941) <= (layer3_outputs(82)) and not (layer3_outputs(2450));
    layer4_outputs(1942) <= (layer3_outputs(130)) and (layer3_outputs(512));
    layer4_outputs(1943) <= layer3_outputs(879);
    layer4_outputs(1944) <= (layer3_outputs(154)) and not (layer3_outputs(2327));
    layer4_outputs(1945) <= not(layer3_outputs(149)) or (layer3_outputs(163));
    layer4_outputs(1946) <= layer3_outputs(442);
    layer4_outputs(1947) <= layer3_outputs(1140);
    layer4_outputs(1948) <= layer3_outputs(791);
    layer4_outputs(1949) <= not(layer3_outputs(69));
    layer4_outputs(1950) <= layer3_outputs(1919);
    layer4_outputs(1951) <= (layer3_outputs(2286)) or (layer3_outputs(2312));
    layer4_outputs(1952) <= (layer3_outputs(727)) and not (layer3_outputs(2417));
    layer4_outputs(1953) <= not((layer3_outputs(495)) or (layer3_outputs(2546)));
    layer4_outputs(1954) <= '1';
    layer4_outputs(1955) <= not(layer3_outputs(1310));
    layer4_outputs(1956) <= layer3_outputs(2425);
    layer4_outputs(1957) <= not((layer3_outputs(1926)) xor (layer3_outputs(2137)));
    layer4_outputs(1958) <= layer3_outputs(1362);
    layer4_outputs(1959) <= '0';
    layer4_outputs(1960) <= (layer3_outputs(2502)) and not (layer3_outputs(494));
    layer4_outputs(1961) <= not(layer3_outputs(244));
    layer4_outputs(1962) <= not(layer3_outputs(1348)) or (layer3_outputs(685));
    layer4_outputs(1963) <= (layer3_outputs(711)) xor (layer3_outputs(805));
    layer4_outputs(1964) <= not((layer3_outputs(2130)) xor (layer3_outputs(368)));
    layer4_outputs(1965) <= not(layer3_outputs(1976));
    layer4_outputs(1966) <= (layer3_outputs(104)) xor (layer3_outputs(1388));
    layer4_outputs(1967) <= not(layer3_outputs(794));
    layer4_outputs(1968) <= '0';
    layer4_outputs(1969) <= layer3_outputs(34);
    layer4_outputs(1970) <= layer3_outputs(2306);
    layer4_outputs(1971) <= (layer3_outputs(1183)) and (layer3_outputs(1059));
    layer4_outputs(1972) <= not(layer3_outputs(1693));
    layer4_outputs(1973) <= (layer3_outputs(1789)) and (layer3_outputs(2022));
    layer4_outputs(1974) <= not((layer3_outputs(803)) or (layer3_outputs(2216)));
    layer4_outputs(1975) <= not(layer3_outputs(1360));
    layer4_outputs(1976) <= not(layer3_outputs(1320));
    layer4_outputs(1977) <= (layer3_outputs(1651)) and not (layer3_outputs(1316));
    layer4_outputs(1978) <= not(layer3_outputs(47)) or (layer3_outputs(2198));
    layer4_outputs(1979) <= (layer3_outputs(2355)) and (layer3_outputs(1129));
    layer4_outputs(1980) <= not((layer3_outputs(589)) or (layer3_outputs(2384)));
    layer4_outputs(1981) <= '0';
    layer4_outputs(1982) <= not(layer3_outputs(435));
    layer4_outputs(1983) <= not(layer3_outputs(1882));
    layer4_outputs(1984) <= not(layer3_outputs(1262)) or (layer3_outputs(1773));
    layer4_outputs(1985) <= (layer3_outputs(953)) or (layer3_outputs(860));
    layer4_outputs(1986) <= '1';
    layer4_outputs(1987) <= '1';
    layer4_outputs(1988) <= not((layer3_outputs(1252)) and (layer3_outputs(1795)));
    layer4_outputs(1989) <= layer3_outputs(1791);
    layer4_outputs(1990) <= not(layer3_outputs(1988));
    layer4_outputs(1991) <= not(layer3_outputs(2436));
    layer4_outputs(1992) <= layer3_outputs(1416);
    layer4_outputs(1993) <= not(layer3_outputs(1484));
    layer4_outputs(1994) <= not(layer3_outputs(584));
    layer4_outputs(1995) <= '1';
    layer4_outputs(1996) <= (layer3_outputs(2500)) and (layer3_outputs(1616));
    layer4_outputs(1997) <= not(layer3_outputs(439)) or (layer3_outputs(1321));
    layer4_outputs(1998) <= layer3_outputs(1280);
    layer4_outputs(1999) <= not(layer3_outputs(974)) or (layer3_outputs(858));
    layer4_outputs(2000) <= layer3_outputs(2232);
    layer4_outputs(2001) <= '1';
    layer4_outputs(2002) <= (layer3_outputs(238)) and not (layer3_outputs(944));
    layer4_outputs(2003) <= layer3_outputs(1916);
    layer4_outputs(2004) <= not((layer3_outputs(741)) and (layer3_outputs(1376)));
    layer4_outputs(2005) <= not((layer3_outputs(2538)) or (layer3_outputs(1788)));
    layer4_outputs(2006) <= not((layer3_outputs(1635)) or (layer3_outputs(220)));
    layer4_outputs(2007) <= not((layer3_outputs(1461)) and (layer3_outputs(1496)));
    layer4_outputs(2008) <= not(layer3_outputs(1169));
    layer4_outputs(2009) <= (layer3_outputs(2254)) and not (layer3_outputs(2324));
    layer4_outputs(2010) <= not(layer3_outputs(334)) or (layer3_outputs(2377));
    layer4_outputs(2011) <= not(layer3_outputs(2520));
    layer4_outputs(2012) <= not((layer3_outputs(1450)) or (layer3_outputs(2037)));
    layer4_outputs(2013) <= not((layer3_outputs(2370)) xor (layer3_outputs(1662)));
    layer4_outputs(2014) <= '0';
    layer4_outputs(2015) <= layer3_outputs(2414);
    layer4_outputs(2016) <= not(layer3_outputs(2040)) or (layer3_outputs(877));
    layer4_outputs(2017) <= not(layer3_outputs(1948));
    layer4_outputs(2018) <= '1';
    layer4_outputs(2019) <= layer3_outputs(106);
    layer4_outputs(2020) <= not(layer3_outputs(929));
    layer4_outputs(2021) <= not(layer3_outputs(2002));
    layer4_outputs(2022) <= '0';
    layer4_outputs(2023) <= (layer3_outputs(504)) and not (layer3_outputs(1877));
    layer4_outputs(2024) <= not(layer3_outputs(2139));
    layer4_outputs(2025) <= layer3_outputs(2334);
    layer4_outputs(2026) <= (layer3_outputs(836)) and not (layer3_outputs(2292));
    layer4_outputs(2027) <= layer3_outputs(2397);
    layer4_outputs(2028) <= (layer3_outputs(220)) or (layer3_outputs(2501));
    layer4_outputs(2029) <= not(layer3_outputs(1231)) or (layer3_outputs(296));
    layer4_outputs(2030) <= '0';
    layer4_outputs(2031) <= not(layer3_outputs(1560));
    layer4_outputs(2032) <= not(layer3_outputs(1858));
    layer4_outputs(2033) <= (layer3_outputs(1494)) and (layer3_outputs(836));
    layer4_outputs(2034) <= layer3_outputs(1938);
    layer4_outputs(2035) <= layer3_outputs(2089);
    layer4_outputs(2036) <= '1';
    layer4_outputs(2037) <= layer3_outputs(2016);
    layer4_outputs(2038) <= '0';
    layer4_outputs(2039) <= '0';
    layer4_outputs(2040) <= not(layer3_outputs(1943));
    layer4_outputs(2041) <= (layer3_outputs(1431)) or (layer3_outputs(790));
    layer4_outputs(2042) <= layer3_outputs(797);
    layer4_outputs(2043) <= not(layer3_outputs(494));
    layer4_outputs(2044) <= not((layer3_outputs(2275)) or (layer3_outputs(105)));
    layer4_outputs(2045) <= '1';
    layer4_outputs(2046) <= (layer3_outputs(1515)) and (layer3_outputs(1862));
    layer4_outputs(2047) <= (layer3_outputs(134)) and not (layer3_outputs(318));
    layer4_outputs(2048) <= not(layer3_outputs(1382));
    layer4_outputs(2049) <= (layer3_outputs(270)) and not (layer3_outputs(140));
    layer4_outputs(2050) <= (layer3_outputs(986)) and not (layer3_outputs(427));
    layer4_outputs(2051) <= (layer3_outputs(2015)) and not (layer3_outputs(2473));
    layer4_outputs(2052) <= (layer3_outputs(1229)) and (layer3_outputs(202));
    layer4_outputs(2053) <= not(layer3_outputs(2300));
    layer4_outputs(2054) <= (layer3_outputs(594)) and not (layer3_outputs(833));
    layer4_outputs(2055) <= not(layer3_outputs(1529));
    layer4_outputs(2056) <= layer3_outputs(254);
    layer4_outputs(2057) <= (layer3_outputs(1142)) or (layer3_outputs(1488));
    layer4_outputs(2058) <= (layer3_outputs(747)) and not (layer3_outputs(336));
    layer4_outputs(2059) <= layer3_outputs(558);
    layer4_outputs(2060) <= not(layer3_outputs(1107)) or (layer3_outputs(1907));
    layer4_outputs(2061) <= not(layer3_outputs(1030)) or (layer3_outputs(881));
    layer4_outputs(2062) <= (layer3_outputs(1855)) and (layer3_outputs(1718));
    layer4_outputs(2063) <= (layer3_outputs(439)) or (layer3_outputs(2136));
    layer4_outputs(2064) <= (layer3_outputs(412)) and not (layer3_outputs(1624));
    layer4_outputs(2065) <= (layer3_outputs(761)) and (layer3_outputs(2550));
    layer4_outputs(2066) <= (layer3_outputs(1803)) and not (layer3_outputs(1301));
    layer4_outputs(2067) <= layer3_outputs(962);
    layer4_outputs(2068) <= not(layer3_outputs(1474));
    layer4_outputs(2069) <= (layer3_outputs(2226)) and not (layer3_outputs(2035));
    layer4_outputs(2070) <= not(layer3_outputs(171));
    layer4_outputs(2071) <= not(layer3_outputs(1872));
    layer4_outputs(2072) <= not(layer3_outputs(1944)) or (layer3_outputs(1891));
    layer4_outputs(2073) <= layer3_outputs(460);
    layer4_outputs(2074) <= layer3_outputs(1409);
    layer4_outputs(2075) <= not(layer3_outputs(859));
    layer4_outputs(2076) <= not((layer3_outputs(1617)) and (layer3_outputs(1534)));
    layer4_outputs(2077) <= not(layer3_outputs(2460)) or (layer3_outputs(2498));
    layer4_outputs(2078) <= layer3_outputs(639);
    layer4_outputs(2079) <= layer3_outputs(351);
    layer4_outputs(2080) <= (layer3_outputs(1078)) xor (layer3_outputs(498));
    layer4_outputs(2081) <= not(layer3_outputs(951)) or (layer3_outputs(1067));
    layer4_outputs(2082) <= not(layer3_outputs(2084)) or (layer3_outputs(456));
    layer4_outputs(2083) <= layer3_outputs(878);
    layer4_outputs(2084) <= (layer3_outputs(2559)) or (layer3_outputs(124));
    layer4_outputs(2085) <= (layer3_outputs(588)) and not (layer3_outputs(1780));
    layer4_outputs(2086) <= layer3_outputs(663);
    layer4_outputs(2087) <= not(layer3_outputs(1619));
    layer4_outputs(2088) <= layer3_outputs(1238);
    layer4_outputs(2089) <= (layer3_outputs(1109)) or (layer3_outputs(1787));
    layer4_outputs(2090) <= (layer3_outputs(718)) and not (layer3_outputs(2215));
    layer4_outputs(2091) <= '0';
    layer4_outputs(2092) <= not(layer3_outputs(272));
    layer4_outputs(2093) <= (layer3_outputs(1063)) and not (layer3_outputs(831));
    layer4_outputs(2094) <= not((layer3_outputs(1210)) and (layer3_outputs(869)));
    layer4_outputs(2095) <= (layer3_outputs(913)) and (layer3_outputs(1923));
    layer4_outputs(2096) <= (layer3_outputs(450)) and not (layer3_outputs(2101));
    layer4_outputs(2097) <= not(layer3_outputs(1661)) or (layer3_outputs(1884));
    layer4_outputs(2098) <= layer3_outputs(115);
    layer4_outputs(2099) <= (layer3_outputs(35)) or (layer3_outputs(1986));
    layer4_outputs(2100) <= (layer3_outputs(133)) xor (layer3_outputs(1062));
    layer4_outputs(2101) <= '1';
    layer4_outputs(2102) <= not(layer3_outputs(1174)) or (layer3_outputs(1453));
    layer4_outputs(2103) <= '0';
    layer4_outputs(2104) <= not(layer3_outputs(1614));
    layer4_outputs(2105) <= not(layer3_outputs(31)) or (layer3_outputs(2094));
    layer4_outputs(2106) <= (layer3_outputs(211)) and not (layer3_outputs(1873));
    layer4_outputs(2107) <= layer3_outputs(288);
    layer4_outputs(2108) <= layer3_outputs(644);
    layer4_outputs(2109) <= not((layer3_outputs(933)) xor (layer3_outputs(1605)));
    layer4_outputs(2110) <= layer3_outputs(1444);
    layer4_outputs(2111) <= '1';
    layer4_outputs(2112) <= (layer3_outputs(757)) and not (layer3_outputs(2091));
    layer4_outputs(2113) <= layer3_outputs(1845);
    layer4_outputs(2114) <= (layer3_outputs(1243)) and not (layer3_outputs(2368));
    layer4_outputs(2115) <= layer3_outputs(1844);
    layer4_outputs(2116) <= layer3_outputs(995);
    layer4_outputs(2117) <= not((layer3_outputs(809)) or (layer3_outputs(1136)));
    layer4_outputs(2118) <= (layer3_outputs(1940)) or (layer3_outputs(952));
    layer4_outputs(2119) <= not((layer3_outputs(1869)) and (layer3_outputs(1691)));
    layer4_outputs(2120) <= not((layer3_outputs(2513)) and (layer3_outputs(1163)));
    layer4_outputs(2121) <= (layer3_outputs(2301)) and not (layer3_outputs(1835));
    layer4_outputs(2122) <= (layer3_outputs(1180)) and not (layer3_outputs(484));
    layer4_outputs(2123) <= not((layer3_outputs(1422)) or (layer3_outputs(1255)));
    layer4_outputs(2124) <= (layer3_outputs(1332)) and not (layer3_outputs(2387));
    layer4_outputs(2125) <= not((layer3_outputs(855)) or (layer3_outputs(1242)));
    layer4_outputs(2126) <= layer3_outputs(369);
    layer4_outputs(2127) <= not(layer3_outputs(1317));
    layer4_outputs(2128) <= (layer3_outputs(2051)) xor (layer3_outputs(1220));
    layer4_outputs(2129) <= not((layer3_outputs(1691)) or (layer3_outputs(245)));
    layer4_outputs(2130) <= (layer3_outputs(832)) xor (layer3_outputs(1007));
    layer4_outputs(2131) <= layer3_outputs(2549);
    layer4_outputs(2132) <= (layer3_outputs(2128)) and not (layer3_outputs(826));
    layer4_outputs(2133) <= not(layer3_outputs(2264));
    layer4_outputs(2134) <= layer3_outputs(2010);
    layer4_outputs(2135) <= not(layer3_outputs(1641)) or (layer3_outputs(825));
    layer4_outputs(2136) <= not(layer3_outputs(1065)) or (layer3_outputs(2497));
    layer4_outputs(2137) <= not((layer3_outputs(1922)) and (layer3_outputs(2354)));
    layer4_outputs(2138) <= '1';
    layer4_outputs(2139) <= not(layer3_outputs(1682)) or (layer3_outputs(536));
    layer4_outputs(2140) <= not(layer3_outputs(1310));
    layer4_outputs(2141) <= layer3_outputs(1201);
    layer4_outputs(2142) <= (layer3_outputs(430)) and not (layer3_outputs(470));
    layer4_outputs(2143) <= not((layer3_outputs(152)) and (layer3_outputs(821)));
    layer4_outputs(2144) <= (layer3_outputs(2471)) and not (layer3_outputs(776));
    layer4_outputs(2145) <= not((layer3_outputs(1079)) xor (layer3_outputs(2083)));
    layer4_outputs(2146) <= layer3_outputs(110);
    layer4_outputs(2147) <= layer3_outputs(1822);
    layer4_outputs(2148) <= not(layer3_outputs(1046)) or (layer3_outputs(2168));
    layer4_outputs(2149) <= '1';
    layer4_outputs(2150) <= (layer3_outputs(375)) and (layer3_outputs(1904));
    layer4_outputs(2151) <= not(layer3_outputs(1869)) or (layer3_outputs(2547));
    layer4_outputs(2152) <= not(layer3_outputs(1330));
    layer4_outputs(2153) <= (layer3_outputs(549)) and (layer3_outputs(1664));
    layer4_outputs(2154) <= (layer3_outputs(1995)) and not (layer3_outputs(2467));
    layer4_outputs(2155) <= not(layer3_outputs(1367));
    layer4_outputs(2156) <= not((layer3_outputs(1375)) or (layer3_outputs(574)));
    layer4_outputs(2157) <= '1';
    layer4_outputs(2158) <= not(layer3_outputs(1048)) or (layer3_outputs(1029));
    layer4_outputs(2159) <= (layer3_outputs(68)) and not (layer3_outputs(2222));
    layer4_outputs(2160) <= (layer3_outputs(1091)) or (layer3_outputs(18));
    layer4_outputs(2161) <= not(layer3_outputs(482));
    layer4_outputs(2162) <= (layer3_outputs(2158)) and not (layer3_outputs(2053));
    layer4_outputs(2163) <= not(layer3_outputs(1660));
    layer4_outputs(2164) <= (layer3_outputs(398)) and (layer3_outputs(960));
    layer4_outputs(2165) <= layer3_outputs(271);
    layer4_outputs(2166) <= not(layer3_outputs(1986)) or (layer3_outputs(939));
    layer4_outputs(2167) <= (layer3_outputs(1579)) or (layer3_outputs(1295));
    layer4_outputs(2168) <= (layer3_outputs(582)) and (layer3_outputs(2337));
    layer4_outputs(2169) <= '0';
    layer4_outputs(2170) <= not(layer3_outputs(1283)) or (layer3_outputs(1920));
    layer4_outputs(2171) <= '1';
    layer4_outputs(2172) <= not((layer3_outputs(1907)) xor (layer3_outputs(2173)));
    layer4_outputs(2173) <= (layer3_outputs(1683)) and (layer3_outputs(1547));
    layer4_outputs(2174) <= (layer3_outputs(2548)) and (layer3_outputs(658));
    layer4_outputs(2175) <= (layer3_outputs(1459)) and not (layer3_outputs(1327));
    layer4_outputs(2176) <= (layer3_outputs(2247)) or (layer3_outputs(1179));
    layer4_outputs(2177) <= layer3_outputs(1604);
    layer4_outputs(2178) <= (layer3_outputs(530)) xor (layer3_outputs(1814));
    layer4_outputs(2179) <= not(layer3_outputs(671));
    layer4_outputs(2180) <= (layer3_outputs(1464)) and not (layer3_outputs(593));
    layer4_outputs(2181) <= not(layer3_outputs(700)) or (layer3_outputs(1319));
    layer4_outputs(2182) <= layer3_outputs(400);
    layer4_outputs(2183) <= not(layer3_outputs(2075)) or (layer3_outputs(2307));
    layer4_outputs(2184) <= layer3_outputs(1559);
    layer4_outputs(2185) <= not(layer3_outputs(1277)) or (layer3_outputs(184));
    layer4_outputs(2186) <= not(layer3_outputs(1669));
    layer4_outputs(2187) <= not((layer3_outputs(454)) xor (layer3_outputs(1646)));
    layer4_outputs(2188) <= (layer3_outputs(204)) and (layer3_outputs(573));
    layer4_outputs(2189) <= not(layer3_outputs(935)) or (layer3_outputs(368));
    layer4_outputs(2190) <= not(layer3_outputs(519));
    layer4_outputs(2191) <= layer3_outputs(2474);
    layer4_outputs(2192) <= (layer3_outputs(2447)) and not (layer3_outputs(613));
    layer4_outputs(2193) <= (layer3_outputs(89)) and not (layer3_outputs(721));
    layer4_outputs(2194) <= not(layer3_outputs(778)) or (layer3_outputs(2515));
    layer4_outputs(2195) <= not(layer3_outputs(605));
    layer4_outputs(2196) <= (layer3_outputs(2106)) and (layer3_outputs(905));
    layer4_outputs(2197) <= (layer3_outputs(1685)) and not (layer3_outputs(1213));
    layer4_outputs(2198) <= not(layer3_outputs(1631));
    layer4_outputs(2199) <= (layer3_outputs(1299)) or (layer3_outputs(2079));
    layer4_outputs(2200) <= not((layer3_outputs(1155)) and (layer3_outputs(1418)));
    layer4_outputs(2201) <= not(layer3_outputs(334));
    layer4_outputs(2202) <= layer3_outputs(1735);
    layer4_outputs(2203) <= not(layer3_outputs(2353));
    layer4_outputs(2204) <= (layer3_outputs(524)) and not (layer3_outputs(2330));
    layer4_outputs(2205) <= not(layer3_outputs(23));
    layer4_outputs(2206) <= not(layer3_outputs(106));
    layer4_outputs(2207) <= layer3_outputs(1163);
    layer4_outputs(2208) <= not(layer3_outputs(1053));
    layer4_outputs(2209) <= (layer3_outputs(1289)) xor (layer3_outputs(1027));
    layer4_outputs(2210) <= '0';
    layer4_outputs(2211) <= (layer3_outputs(894)) xor (layer3_outputs(126));
    layer4_outputs(2212) <= not(layer3_outputs(2153)) or (layer3_outputs(2422));
    layer4_outputs(2213) <= (layer3_outputs(787)) and not (layer3_outputs(2424));
    layer4_outputs(2214) <= (layer3_outputs(1124)) and (layer3_outputs(2051));
    layer4_outputs(2215) <= not(layer3_outputs(1658));
    layer4_outputs(2216) <= (layer3_outputs(1403)) or (layer3_outputs(1665));
    layer4_outputs(2217) <= not(layer3_outputs(761));
    layer4_outputs(2218) <= not(layer3_outputs(827)) or (layer3_outputs(1373));
    layer4_outputs(2219) <= layer3_outputs(934);
    layer4_outputs(2220) <= not(layer3_outputs(1942));
    layer4_outputs(2221) <= '1';
    layer4_outputs(2222) <= (layer3_outputs(990)) or (layer3_outputs(1053));
    layer4_outputs(2223) <= layer3_outputs(1561);
    layer4_outputs(2224) <= not(layer3_outputs(698));
    layer4_outputs(2225) <= (layer3_outputs(961)) and not (layer3_outputs(207));
    layer4_outputs(2226) <= (layer3_outputs(2544)) and (layer3_outputs(142));
    layer4_outputs(2227) <= not(layer3_outputs(1610));
    layer4_outputs(2228) <= '1';
    layer4_outputs(2229) <= (layer3_outputs(226)) xor (layer3_outputs(1501));
    layer4_outputs(2230) <= (layer3_outputs(902)) and not (layer3_outputs(1067));
    layer4_outputs(2231) <= not(layer3_outputs(17)) or (layer3_outputs(1759));
    layer4_outputs(2232) <= (layer3_outputs(2319)) and not (layer3_outputs(289));
    layer4_outputs(2233) <= layer3_outputs(980);
    layer4_outputs(2234) <= not(layer3_outputs(2227));
    layer4_outputs(2235) <= (layer3_outputs(2250)) xor (layer3_outputs(289));
    layer4_outputs(2236) <= layer3_outputs(818);
    layer4_outputs(2237) <= layer3_outputs(741);
    layer4_outputs(2238) <= layer3_outputs(318);
    layer4_outputs(2239) <= not(layer3_outputs(393));
    layer4_outputs(2240) <= not((layer3_outputs(838)) and (layer3_outputs(806)));
    layer4_outputs(2241) <= (layer3_outputs(965)) and (layer3_outputs(2356));
    layer4_outputs(2242) <= (layer3_outputs(661)) and (layer3_outputs(1657));
    layer4_outputs(2243) <= (layer3_outputs(1916)) and not (layer3_outputs(527));
    layer4_outputs(2244) <= '0';
    layer4_outputs(2245) <= (layer3_outputs(1467)) and (layer3_outputs(1164));
    layer4_outputs(2246) <= '1';
    layer4_outputs(2247) <= (layer3_outputs(2536)) xor (layer3_outputs(1369));
    layer4_outputs(2248) <= layer3_outputs(170);
    layer4_outputs(2249) <= layer3_outputs(1805);
    layer4_outputs(2250) <= (layer3_outputs(1816)) and (layer3_outputs(2214));
    layer4_outputs(2251) <= (layer3_outputs(1853)) and not (layer3_outputs(1189));
    layer4_outputs(2252) <= (layer3_outputs(1093)) or (layer3_outputs(262));
    layer4_outputs(2253) <= layer3_outputs(982);
    layer4_outputs(2254) <= not(layer3_outputs(199));
    layer4_outputs(2255) <= '0';
    layer4_outputs(2256) <= (layer3_outputs(388)) and not (layer3_outputs(748));
    layer4_outputs(2257) <= (layer3_outputs(1205)) and (layer3_outputs(1830));
    layer4_outputs(2258) <= not((layer3_outputs(2196)) or (layer3_outputs(1432)));
    layer4_outputs(2259) <= not(layer3_outputs(1931));
    layer4_outputs(2260) <= (layer3_outputs(2454)) xor (layer3_outputs(1724));
    layer4_outputs(2261) <= not((layer3_outputs(954)) and (layer3_outputs(555)));
    layer4_outputs(2262) <= (layer3_outputs(1627)) and (layer3_outputs(197));
    layer4_outputs(2263) <= '0';
    layer4_outputs(2264) <= not(layer3_outputs(432));
    layer4_outputs(2265) <= not(layer3_outputs(1999));
    layer4_outputs(2266) <= not((layer3_outputs(1679)) or (layer3_outputs(13)));
    layer4_outputs(2267) <= not(layer3_outputs(1439));
    layer4_outputs(2268) <= not(layer3_outputs(2522)) or (layer3_outputs(548));
    layer4_outputs(2269) <= layer3_outputs(2059);
    layer4_outputs(2270) <= layer3_outputs(2071);
    layer4_outputs(2271) <= not(layer3_outputs(1866)) or (layer3_outputs(1671));
    layer4_outputs(2272) <= layer3_outputs(1678);
    layer4_outputs(2273) <= not((layer3_outputs(1178)) xor (layer3_outputs(1654)));
    layer4_outputs(2274) <= not((layer3_outputs(756)) xor (layer3_outputs(1614)));
    layer4_outputs(2275) <= layer3_outputs(1681);
    layer4_outputs(2276) <= not(layer3_outputs(1837));
    layer4_outputs(2277) <= layer3_outputs(2497);
    layer4_outputs(2278) <= layer3_outputs(2357);
    layer4_outputs(2279) <= not(layer3_outputs(930));
    layer4_outputs(2280) <= layer3_outputs(2323);
    layer4_outputs(2281) <= layer3_outputs(2537);
    layer4_outputs(2282) <= not(layer3_outputs(2232));
    layer4_outputs(2283) <= (layer3_outputs(2242)) xor (layer3_outputs(2529));
    layer4_outputs(2284) <= not((layer3_outputs(1736)) or (layer3_outputs(96)));
    layer4_outputs(2285) <= not((layer3_outputs(870)) or (layer3_outputs(1345)));
    layer4_outputs(2286) <= (layer3_outputs(254)) and (layer3_outputs(1197));
    layer4_outputs(2287) <= not(layer3_outputs(118));
    layer4_outputs(2288) <= (layer3_outputs(2098)) and not (layer3_outputs(1871));
    layer4_outputs(2289) <= (layer3_outputs(357)) or (layer3_outputs(1980));
    layer4_outputs(2290) <= '1';
    layer4_outputs(2291) <= (layer3_outputs(2183)) and not (layer3_outputs(1459));
    layer4_outputs(2292) <= layer3_outputs(41);
    layer4_outputs(2293) <= not(layer3_outputs(839)) or (layer3_outputs(1300));
    layer4_outputs(2294) <= not((layer3_outputs(1808)) or (layer3_outputs(50)));
    layer4_outputs(2295) <= not((layer3_outputs(1108)) and (layer3_outputs(2339)));
    layer4_outputs(2296) <= layer3_outputs(1111);
    layer4_outputs(2297) <= not((layer3_outputs(1415)) and (layer3_outputs(1890)));
    layer4_outputs(2298) <= not(layer3_outputs(547));
    layer4_outputs(2299) <= layer3_outputs(485);
    layer4_outputs(2300) <= not(layer3_outputs(1350)) or (layer3_outputs(1174));
    layer4_outputs(2301) <= not(layer3_outputs(1770));
    layer4_outputs(2302) <= not(layer3_outputs(1348)) or (layer3_outputs(992));
    layer4_outputs(2303) <= not(layer3_outputs(1292)) or (layer3_outputs(513));
    layer4_outputs(2304) <= (layer3_outputs(1841)) and not (layer3_outputs(547));
    layer4_outputs(2305) <= (layer3_outputs(265)) xor (layer3_outputs(2288));
    layer4_outputs(2306) <= (layer3_outputs(1448)) or (layer3_outputs(2231));
    layer4_outputs(2307) <= layer3_outputs(508);
    layer4_outputs(2308) <= '1';
    layer4_outputs(2309) <= not(layer3_outputs(1482));
    layer4_outputs(2310) <= '0';
    layer4_outputs(2311) <= layer3_outputs(556);
    layer4_outputs(2312) <= not(layer3_outputs(1872));
    layer4_outputs(2313) <= not(layer3_outputs(525));
    layer4_outputs(2314) <= not(layer3_outputs(2035));
    layer4_outputs(2315) <= not(layer3_outputs(1946));
    layer4_outputs(2316) <= not(layer3_outputs(2401));
    layer4_outputs(2317) <= (layer3_outputs(139)) and not (layer3_outputs(979));
    layer4_outputs(2318) <= layer3_outputs(2408);
    layer4_outputs(2319) <= not(layer3_outputs(1044)) or (layer3_outputs(1499));
    layer4_outputs(2320) <= not((layer3_outputs(2341)) or (layer3_outputs(279)));
    layer4_outputs(2321) <= (layer3_outputs(1207)) xor (layer3_outputs(2099));
    layer4_outputs(2322) <= not(layer3_outputs(2312));
    layer4_outputs(2323) <= (layer3_outputs(2145)) xor (layer3_outputs(634));
    layer4_outputs(2324) <= (layer3_outputs(572)) and not (layer3_outputs(616));
    layer4_outputs(2325) <= not(layer3_outputs(305));
    layer4_outputs(2326) <= (layer3_outputs(2458)) and not (layer3_outputs(2054));
    layer4_outputs(2327) <= not(layer3_outputs(788)) or (layer3_outputs(1532));
    layer4_outputs(2328) <= layer3_outputs(239);
    layer4_outputs(2329) <= not(layer3_outputs(1471));
    layer4_outputs(2330) <= not(layer3_outputs(1137)) or (layer3_outputs(1838));
    layer4_outputs(2331) <= not(layer3_outputs(1761));
    layer4_outputs(2332) <= layer3_outputs(2186);
    layer4_outputs(2333) <= (layer3_outputs(1190)) and not (layer3_outputs(1036));
    layer4_outputs(2334) <= not(layer3_outputs(1283));
    layer4_outputs(2335) <= (layer3_outputs(1447)) and (layer3_outputs(2167));
    layer4_outputs(2336) <= '0';
    layer4_outputs(2337) <= not(layer3_outputs(1663));
    layer4_outputs(2338) <= layer3_outputs(1419);
    layer4_outputs(2339) <= not(layer3_outputs(1805)) or (layer3_outputs(292));
    layer4_outputs(2340) <= not(layer3_outputs(606)) or (layer3_outputs(1854));
    layer4_outputs(2341) <= not(layer3_outputs(151)) or (layer3_outputs(2174));
    layer4_outputs(2342) <= (layer3_outputs(896)) and (layer3_outputs(2512));
    layer4_outputs(2343) <= not(layer3_outputs(292));
    layer4_outputs(2344) <= (layer3_outputs(2337)) and not (layer3_outputs(666));
    layer4_outputs(2345) <= (layer3_outputs(1180)) and (layer3_outputs(1162));
    layer4_outputs(2346) <= layer3_outputs(2302);
    layer4_outputs(2347) <= layer3_outputs(759);
    layer4_outputs(2348) <= not((layer3_outputs(1196)) or (layer3_outputs(1810)));
    layer4_outputs(2349) <= (layer3_outputs(1076)) xor (layer3_outputs(1049));
    layer4_outputs(2350) <= (layer3_outputs(122)) and not (layer3_outputs(2074));
    layer4_outputs(2351) <= not(layer3_outputs(906));
    layer4_outputs(2352) <= not(layer3_outputs(1602)) or (layer3_outputs(131));
    layer4_outputs(2353) <= '1';
    layer4_outputs(2354) <= not(layer3_outputs(1909));
    layer4_outputs(2355) <= layer3_outputs(1700);
    layer4_outputs(2356) <= not(layer3_outputs(1300));
    layer4_outputs(2357) <= '0';
    layer4_outputs(2358) <= layer3_outputs(2539);
    layer4_outputs(2359) <= not((layer3_outputs(348)) xor (layer3_outputs(49)));
    layer4_outputs(2360) <= layer3_outputs(1639);
    layer4_outputs(2361) <= (layer3_outputs(283)) and not (layer3_outputs(1045));
    layer4_outputs(2362) <= (layer3_outputs(653)) or (layer3_outputs(1485));
    layer4_outputs(2363) <= (layer3_outputs(681)) and (layer3_outputs(1404));
    layer4_outputs(2364) <= layer3_outputs(159);
    layer4_outputs(2365) <= not(layer3_outputs(2499)) or (layer3_outputs(1509));
    layer4_outputs(2366) <= not(layer3_outputs(2055)) or (layer3_outputs(2376));
    layer4_outputs(2367) <= (layer3_outputs(1073)) and not (layer3_outputs(605));
    layer4_outputs(2368) <= layer3_outputs(346);
    layer4_outputs(2369) <= (layer3_outputs(249)) xor (layer3_outputs(946));
    layer4_outputs(2370) <= '1';
    layer4_outputs(2371) <= not((layer3_outputs(2003)) or (layer3_outputs(420)));
    layer4_outputs(2372) <= layer3_outputs(1119);
    layer4_outputs(2373) <= not(layer3_outputs(150));
    layer4_outputs(2374) <= layer3_outputs(657);
    layer4_outputs(2375) <= (layer3_outputs(297)) and (layer3_outputs(2113));
    layer4_outputs(2376) <= not(layer3_outputs(1772));
    layer4_outputs(2377) <= '0';
    layer4_outputs(2378) <= (layer3_outputs(1019)) and not (layer3_outputs(1354));
    layer4_outputs(2379) <= (layer3_outputs(2052)) or (layer3_outputs(1733));
    layer4_outputs(2380) <= not(layer3_outputs(817));
    layer4_outputs(2381) <= (layer3_outputs(1127)) and (layer3_outputs(754));
    layer4_outputs(2382) <= not(layer3_outputs(1903));
    layer4_outputs(2383) <= (layer3_outputs(1841)) and not (layer3_outputs(1695));
    layer4_outputs(2384) <= (layer3_outputs(1589)) or (layer3_outputs(214));
    layer4_outputs(2385) <= not((layer3_outputs(1699)) xor (layer3_outputs(1542)));
    layer4_outputs(2386) <= layer3_outputs(880);
    layer4_outputs(2387) <= layer3_outputs(595);
    layer4_outputs(2388) <= not((layer3_outputs(565)) or (layer3_outputs(1186)));
    layer4_outputs(2389) <= (layer3_outputs(2144)) and (layer3_outputs(1878));
    layer4_outputs(2390) <= (layer3_outputs(479)) and not (layer3_outputs(285));
    layer4_outputs(2391) <= layer3_outputs(2163);
    layer4_outputs(2392) <= not(layer3_outputs(2311));
    layer4_outputs(2393) <= not(layer3_outputs(695)) or (layer3_outputs(2412));
    layer4_outputs(2394) <= (layer3_outputs(102)) and not (layer3_outputs(162));
    layer4_outputs(2395) <= not(layer3_outputs(2161));
    layer4_outputs(2396) <= not(layer3_outputs(1964)) or (layer3_outputs(919));
    layer4_outputs(2397) <= (layer3_outputs(2503)) and not (layer3_outputs(71));
    layer4_outputs(2398) <= not((layer3_outputs(1657)) or (layer3_outputs(2363)));
    layer4_outputs(2399) <= not((layer3_outputs(2138)) and (layer3_outputs(1315)));
    layer4_outputs(2400) <= not((layer3_outputs(1201)) and (layer3_outputs(926)));
    layer4_outputs(2401) <= not(layer3_outputs(373)) or (layer3_outputs(520));
    layer4_outputs(2402) <= (layer3_outputs(1735)) or (layer3_outputs(979));
    layer4_outputs(2403) <= layer3_outputs(319);
    layer4_outputs(2404) <= (layer3_outputs(2400)) and not (layer3_outputs(843));
    layer4_outputs(2405) <= layer3_outputs(1246);
    layer4_outputs(2406) <= (layer3_outputs(655)) or (layer3_outputs(1506));
    layer4_outputs(2407) <= not(layer3_outputs(709));
    layer4_outputs(2408) <= layer3_outputs(25);
    layer4_outputs(2409) <= not(layer3_outputs(919));
    layer4_outputs(2410) <= layer3_outputs(303);
    layer4_outputs(2411) <= not((layer3_outputs(538)) and (layer3_outputs(1842)));
    layer4_outputs(2412) <= not(layer3_outputs(1975));
    layer4_outputs(2413) <= not(layer3_outputs(1424)) or (layer3_outputs(751));
    layer4_outputs(2414) <= not(layer3_outputs(640)) or (layer3_outputs(780));
    layer4_outputs(2415) <= not(layer3_outputs(1069)) or (layer3_outputs(1109));
    layer4_outputs(2416) <= layer3_outputs(608);
    layer4_outputs(2417) <= not(layer3_outputs(1956)) or (layer3_outputs(1957));
    layer4_outputs(2418) <= (layer3_outputs(708)) and not (layer3_outputs(789));
    layer4_outputs(2419) <= '1';
    layer4_outputs(2420) <= (layer3_outputs(2227)) or (layer3_outputs(2047));
    layer4_outputs(2421) <= not(layer3_outputs(298));
    layer4_outputs(2422) <= layer3_outputs(134);
    layer4_outputs(2423) <= (layer3_outputs(2156)) and not (layer3_outputs(1237));
    layer4_outputs(2424) <= layer3_outputs(1393);
    layer4_outputs(2425) <= not((layer3_outputs(2394)) and (layer3_outputs(2110)));
    layer4_outputs(2426) <= (layer3_outputs(2398)) and not (layer3_outputs(684));
    layer4_outputs(2427) <= not((layer3_outputs(1294)) or (layer3_outputs(1477)));
    layer4_outputs(2428) <= (layer3_outputs(1643)) and (layer3_outputs(2411));
    layer4_outputs(2429) <= not(layer3_outputs(1752));
    layer4_outputs(2430) <= not(layer3_outputs(1303)) or (layer3_outputs(1652));
    layer4_outputs(2431) <= not(layer3_outputs(1694));
    layer4_outputs(2432) <= (layer3_outputs(1252)) and (layer3_outputs(1361));
    layer4_outputs(2433) <= not(layer3_outputs(1656));
    layer4_outputs(2434) <= layer3_outputs(755);
    layer4_outputs(2435) <= not(layer3_outputs(1004)) or (layer3_outputs(1311));
    layer4_outputs(2436) <= layer3_outputs(427);
    layer4_outputs(2437) <= not((layer3_outputs(1386)) or (layer3_outputs(601)));
    layer4_outputs(2438) <= not(layer3_outputs(1893));
    layer4_outputs(2439) <= not(layer3_outputs(2394)) or (layer3_outputs(499));
    layer4_outputs(2440) <= '0';
    layer4_outputs(2441) <= '1';
    layer4_outputs(2442) <= not(layer3_outputs(1759));
    layer4_outputs(2443) <= not(layer3_outputs(1887)) or (layer3_outputs(1126));
    layer4_outputs(2444) <= (layer3_outputs(1670)) or (layer3_outputs(1185));
    layer4_outputs(2445) <= (layer3_outputs(1831)) or (layer3_outputs(2547));
    layer4_outputs(2446) <= not(layer3_outputs(1354));
    layer4_outputs(2447) <= (layer3_outputs(266)) and (layer3_outputs(1359));
    layer4_outputs(2448) <= (layer3_outputs(2459)) and (layer3_outputs(2017));
    layer4_outputs(2449) <= '0';
    layer4_outputs(2450) <= (layer3_outputs(1268)) and not (layer3_outputs(1535));
    layer4_outputs(2451) <= (layer3_outputs(1091)) and (layer3_outputs(1538));
    layer4_outputs(2452) <= (layer3_outputs(396)) and not (layer3_outputs(1562));
    layer4_outputs(2453) <= not(layer3_outputs(1291)) or (layer3_outputs(1808));
    layer4_outputs(2454) <= not(layer3_outputs(1087)) or (layer3_outputs(1220));
    layer4_outputs(2455) <= layer3_outputs(1318);
    layer4_outputs(2456) <= (layer3_outputs(2272)) and not (layer3_outputs(352));
    layer4_outputs(2457) <= (layer3_outputs(352)) and not (layer3_outputs(607));
    layer4_outputs(2458) <= not(layer3_outputs(1539));
    layer4_outputs(2459) <= (layer3_outputs(920)) and not (layer3_outputs(2207));
    layer4_outputs(2460) <= (layer3_outputs(928)) and not (layer3_outputs(1411));
    layer4_outputs(2461) <= layer3_outputs(96);
    layer4_outputs(2462) <= not(layer3_outputs(1288));
    layer4_outputs(2463) <= not((layer3_outputs(1842)) and (layer3_outputs(1764)));
    layer4_outputs(2464) <= layer3_outputs(1915);
    layer4_outputs(2465) <= not(layer3_outputs(1824));
    layer4_outputs(2466) <= (layer3_outputs(2157)) xor (layer3_outputs(397));
    layer4_outputs(2467) <= (layer3_outputs(1737)) and (layer3_outputs(807));
    layer4_outputs(2468) <= layer3_outputs(1114);
    layer4_outputs(2469) <= (layer3_outputs(2430)) and not (layer3_outputs(641));
    layer4_outputs(2470) <= '1';
    layer4_outputs(2471) <= (layer3_outputs(2538)) or (layer3_outputs(1644));
    layer4_outputs(2472) <= not(layer3_outputs(864)) or (layer3_outputs(2095));
    layer4_outputs(2473) <= '0';
    layer4_outputs(2474) <= not(layer3_outputs(2012));
    layer4_outputs(2475) <= not(layer3_outputs(210));
    layer4_outputs(2476) <= not(layer3_outputs(50)) or (layer3_outputs(592));
    layer4_outputs(2477) <= (layer3_outputs(2004)) xor (layer3_outputs(1942));
    layer4_outputs(2478) <= (layer3_outputs(340)) xor (layer3_outputs(275));
    layer4_outputs(2479) <= (layer3_outputs(1391)) and (layer3_outputs(2056));
    layer4_outputs(2480) <= not((layer3_outputs(757)) or (layer3_outputs(2154)));
    layer4_outputs(2481) <= not(layer3_outputs(1944));
    layer4_outputs(2482) <= not(layer3_outputs(2233));
    layer4_outputs(2483) <= not((layer3_outputs(1827)) and (layer3_outputs(1403)));
    layer4_outputs(2484) <= not((layer3_outputs(2187)) or (layer3_outputs(2119)));
    layer4_outputs(2485) <= not(layer3_outputs(308));
    layer4_outputs(2486) <= layer3_outputs(85);
    layer4_outputs(2487) <= not((layer3_outputs(810)) and (layer3_outputs(451)));
    layer4_outputs(2488) <= not((layer3_outputs(1567)) or (layer3_outputs(707)));
    layer4_outputs(2489) <= (layer3_outputs(2005)) or (layer3_outputs(744));
    layer4_outputs(2490) <= not(layer3_outputs(1076)) or (layer3_outputs(1433));
    layer4_outputs(2491) <= not(layer3_outputs(1191)) or (layer3_outputs(433));
    layer4_outputs(2492) <= not(layer3_outputs(703));
    layer4_outputs(2493) <= (layer3_outputs(999)) and (layer3_outputs(635));
    layer4_outputs(2494) <= (layer3_outputs(329)) and (layer3_outputs(1339));
    layer4_outputs(2495) <= not(layer3_outputs(119));
    layer4_outputs(2496) <= not(layer3_outputs(2492));
    layer4_outputs(2497) <= not(layer3_outputs(1615));
    layer4_outputs(2498) <= layer3_outputs(1071);
    layer4_outputs(2499) <= not(layer3_outputs(1550));
    layer4_outputs(2500) <= '1';
    layer4_outputs(2501) <= not(layer3_outputs(1394)) or (layer3_outputs(737));
    layer4_outputs(2502) <= (layer3_outputs(1248)) and not (layer3_outputs(1653));
    layer4_outputs(2503) <= not(layer3_outputs(1229));
    layer4_outputs(2504) <= (layer3_outputs(2448)) and not (layer3_outputs(2019));
    layer4_outputs(2505) <= layer3_outputs(1857);
    layer4_outputs(2506) <= (layer3_outputs(2405)) and (layer3_outputs(1007));
    layer4_outputs(2507) <= not((layer3_outputs(1632)) xor (layer3_outputs(150)));
    layer4_outputs(2508) <= not(layer3_outputs(1480));
    layer4_outputs(2509) <= not((layer3_outputs(2448)) xor (layer3_outputs(443)));
    layer4_outputs(2510) <= layer3_outputs(83);
    layer4_outputs(2511) <= '1';
    layer4_outputs(2512) <= layer3_outputs(768);
    layer4_outputs(2513) <= not(layer3_outputs(2535)) or (layer3_outputs(1832));
    layer4_outputs(2514) <= layer3_outputs(514);
    layer4_outputs(2515) <= (layer3_outputs(102)) xor (layer3_outputs(1296));
    layer4_outputs(2516) <= '1';
    layer4_outputs(2517) <= not(layer3_outputs(645));
    layer4_outputs(2518) <= not(layer3_outputs(1194));
    layer4_outputs(2519) <= (layer3_outputs(503)) and (layer3_outputs(1713));
    layer4_outputs(2520) <= not((layer3_outputs(1151)) and (layer3_outputs(646)));
    layer4_outputs(2521) <= (layer3_outputs(1135)) and (layer3_outputs(390));
    layer4_outputs(2522) <= (layer3_outputs(1478)) and not (layer3_outputs(1871));
    layer4_outputs(2523) <= not((layer3_outputs(1745)) or (layer3_outputs(1301)));
    layer4_outputs(2524) <= (layer3_outputs(1379)) and (layer3_outputs(1849));
    layer4_outputs(2525) <= not(layer3_outputs(2296)) or (layer3_outputs(1431));
    layer4_outputs(2526) <= not(layer3_outputs(780)) or (layer3_outputs(2382));
    layer4_outputs(2527) <= layer3_outputs(185);
    layer4_outputs(2528) <= not(layer3_outputs(2439)) or (layer3_outputs(1249));
    layer4_outputs(2529) <= not(layer3_outputs(1655)) or (layer3_outputs(702));
    layer4_outputs(2530) <= not(layer3_outputs(948));
    layer4_outputs(2531) <= not(layer3_outputs(1378));
    layer4_outputs(2532) <= (layer3_outputs(383)) or (layer3_outputs(2403));
    layer4_outputs(2533) <= not((layer3_outputs(551)) or (layer3_outputs(514)));
    layer4_outputs(2534) <= layer3_outputs(1654);
    layer4_outputs(2535) <= not(layer3_outputs(2101));
    layer4_outputs(2536) <= (layer3_outputs(879)) and not (layer3_outputs(2085));
    layer4_outputs(2537) <= (layer3_outputs(2093)) xor (layer3_outputs(316));
    layer4_outputs(2538) <= (layer3_outputs(1306)) and (layer3_outputs(1092));
    layer4_outputs(2539) <= layer3_outputs(2025);
    layer4_outputs(2540) <= layer3_outputs(1239);
    layer4_outputs(2541) <= not(layer3_outputs(571)) or (layer3_outputs(460));
    layer4_outputs(2542) <= (layer3_outputs(2439)) and not (layer3_outputs(1470));
    layer4_outputs(2543) <= not(layer3_outputs(633)) or (layer3_outputs(1930));
    layer4_outputs(2544) <= layer3_outputs(763);
    layer4_outputs(2545) <= (layer3_outputs(1962)) or (layer3_outputs(2007));
    layer4_outputs(2546) <= layer3_outputs(2270);
    layer4_outputs(2547) <= (layer3_outputs(59)) and not (layer3_outputs(15));
    layer4_outputs(2548) <= layer3_outputs(2155);
    layer4_outputs(2549) <= (layer3_outputs(53)) and not (layer3_outputs(245));
    layer4_outputs(2550) <= not(layer3_outputs(1040)) or (layer3_outputs(1171));
    layer4_outputs(2551) <= not(layer3_outputs(389)) or (layer3_outputs(1593));
    layer4_outputs(2552) <= not(layer3_outputs(2541));
    layer4_outputs(2553) <= (layer3_outputs(1628)) or (layer3_outputs(190));
    layer4_outputs(2554) <= layer3_outputs(116);
    layer4_outputs(2555) <= (layer3_outputs(1839)) and not (layer3_outputs(2351));
    layer4_outputs(2556) <= '0';
    layer4_outputs(2557) <= not(layer3_outputs(1658)) or (layer3_outputs(36));
    layer4_outputs(2558) <= not(layer3_outputs(1169));
    layer4_outputs(2559) <= '1';
    layer5_outputs(0) <= not(layer4_outputs(2017)) or (layer4_outputs(1133));
    layer5_outputs(1) <= layer4_outputs(1484);
    layer5_outputs(2) <= not((layer4_outputs(1817)) and (layer4_outputs(1911)));
    layer5_outputs(3) <= (layer4_outputs(2334)) and (layer4_outputs(182));
    layer5_outputs(4) <= layer4_outputs(50);
    layer5_outputs(5) <= (layer4_outputs(2019)) and (layer4_outputs(646));
    layer5_outputs(6) <= not(layer4_outputs(889));
    layer5_outputs(7) <= not((layer4_outputs(950)) and (layer4_outputs(1690)));
    layer5_outputs(8) <= not(layer4_outputs(1674));
    layer5_outputs(9) <= not(layer4_outputs(1625));
    layer5_outputs(10) <= not((layer4_outputs(1682)) xor (layer4_outputs(1883)));
    layer5_outputs(11) <= not((layer4_outputs(378)) xor (layer4_outputs(2087)));
    layer5_outputs(12) <= not(layer4_outputs(1701));
    layer5_outputs(13) <= not(layer4_outputs(450));
    layer5_outputs(14) <= layer4_outputs(967);
    layer5_outputs(15) <= layer4_outputs(1985);
    layer5_outputs(16) <= not(layer4_outputs(52));
    layer5_outputs(17) <= layer4_outputs(1947);
    layer5_outputs(18) <= not((layer4_outputs(892)) xor (layer4_outputs(2221)));
    layer5_outputs(19) <= layer4_outputs(2507);
    layer5_outputs(20) <= (layer4_outputs(1853)) and (layer4_outputs(64));
    layer5_outputs(21) <= layer4_outputs(2408);
    layer5_outputs(22) <= layer4_outputs(237);
    layer5_outputs(23) <= (layer4_outputs(1840)) and not (layer4_outputs(140));
    layer5_outputs(24) <= layer4_outputs(2067);
    layer5_outputs(25) <= not(layer4_outputs(2359));
    layer5_outputs(26) <= (layer4_outputs(1047)) and (layer4_outputs(2319));
    layer5_outputs(27) <= '0';
    layer5_outputs(28) <= not(layer4_outputs(2109));
    layer5_outputs(29) <= layer4_outputs(261);
    layer5_outputs(30) <= (layer4_outputs(2403)) xor (layer4_outputs(1995));
    layer5_outputs(31) <= not(layer4_outputs(451));
    layer5_outputs(32) <= (layer4_outputs(616)) and not (layer4_outputs(1279));
    layer5_outputs(33) <= (layer4_outputs(1127)) and (layer4_outputs(175));
    layer5_outputs(34) <= not(layer4_outputs(807));
    layer5_outputs(35) <= not(layer4_outputs(1730)) or (layer4_outputs(2445));
    layer5_outputs(36) <= not(layer4_outputs(325));
    layer5_outputs(37) <= layer4_outputs(2534);
    layer5_outputs(38) <= (layer4_outputs(2274)) and not (layer4_outputs(112));
    layer5_outputs(39) <= layer4_outputs(1526);
    layer5_outputs(40) <= not(layer4_outputs(1854));
    layer5_outputs(41) <= not(layer4_outputs(385)) or (layer4_outputs(185));
    layer5_outputs(42) <= (layer4_outputs(1616)) and not (layer4_outputs(591));
    layer5_outputs(43) <= not((layer4_outputs(943)) or (layer4_outputs(2154)));
    layer5_outputs(44) <= not((layer4_outputs(287)) and (layer4_outputs(1767)));
    layer5_outputs(45) <= (layer4_outputs(2492)) and (layer4_outputs(1052));
    layer5_outputs(46) <= not((layer4_outputs(2024)) xor (layer4_outputs(59)));
    layer5_outputs(47) <= layer4_outputs(228);
    layer5_outputs(48) <= not(layer4_outputs(2099));
    layer5_outputs(49) <= not((layer4_outputs(1192)) xor (layer4_outputs(2404)));
    layer5_outputs(50) <= (layer4_outputs(1733)) and not (layer4_outputs(356));
    layer5_outputs(51) <= (layer4_outputs(1367)) and not (layer4_outputs(945));
    layer5_outputs(52) <= not(layer4_outputs(1499));
    layer5_outputs(53) <= (layer4_outputs(1820)) and (layer4_outputs(588));
    layer5_outputs(54) <= not((layer4_outputs(707)) xor (layer4_outputs(2129)));
    layer5_outputs(55) <= not((layer4_outputs(1588)) and (layer4_outputs(634)));
    layer5_outputs(56) <= not(layer4_outputs(414));
    layer5_outputs(57) <= (layer4_outputs(888)) xor (layer4_outputs(1873));
    layer5_outputs(58) <= not(layer4_outputs(739));
    layer5_outputs(59) <= not(layer4_outputs(2474));
    layer5_outputs(60) <= (layer4_outputs(1408)) xor (layer4_outputs(552));
    layer5_outputs(61) <= not((layer4_outputs(746)) or (layer4_outputs(1671)));
    layer5_outputs(62) <= not(layer4_outputs(802));
    layer5_outputs(63) <= layer4_outputs(2069);
    layer5_outputs(64) <= not(layer4_outputs(817));
    layer5_outputs(65) <= layer4_outputs(1625);
    layer5_outputs(66) <= not(layer4_outputs(76));
    layer5_outputs(67) <= layer4_outputs(1680);
    layer5_outputs(68) <= not(layer4_outputs(1760));
    layer5_outputs(69) <= not((layer4_outputs(3)) xor (layer4_outputs(1590)));
    layer5_outputs(70) <= '1';
    layer5_outputs(71) <= layer4_outputs(405);
    layer5_outputs(72) <= layer4_outputs(2181);
    layer5_outputs(73) <= (layer4_outputs(2186)) and (layer4_outputs(1975));
    layer5_outputs(74) <= (layer4_outputs(1784)) xor (layer4_outputs(86));
    layer5_outputs(75) <= not((layer4_outputs(1019)) and (layer4_outputs(1825)));
    layer5_outputs(76) <= not(layer4_outputs(1896));
    layer5_outputs(77) <= layer4_outputs(1314);
    layer5_outputs(78) <= not(layer4_outputs(327));
    layer5_outputs(79) <= (layer4_outputs(1221)) or (layer4_outputs(1672));
    layer5_outputs(80) <= layer4_outputs(2045);
    layer5_outputs(81) <= not((layer4_outputs(2231)) or (layer4_outputs(1045)));
    layer5_outputs(82) <= '0';
    layer5_outputs(83) <= layer4_outputs(949);
    layer5_outputs(84) <= not(layer4_outputs(477));
    layer5_outputs(85) <= layer4_outputs(2094);
    layer5_outputs(86) <= not(layer4_outputs(2285));
    layer5_outputs(87) <= not(layer4_outputs(1178));
    layer5_outputs(88) <= layer4_outputs(2043);
    layer5_outputs(89) <= layer4_outputs(220);
    layer5_outputs(90) <= not((layer4_outputs(1575)) xor (layer4_outputs(2207)));
    layer5_outputs(91) <= not(layer4_outputs(222));
    layer5_outputs(92) <= (layer4_outputs(80)) or (layer4_outputs(1155));
    layer5_outputs(93) <= not(layer4_outputs(1371)) or (layer4_outputs(1689));
    layer5_outputs(94) <= layer4_outputs(1885);
    layer5_outputs(95) <= not(layer4_outputs(1095)) or (layer4_outputs(1318));
    layer5_outputs(96) <= not(layer4_outputs(1873)) or (layer4_outputs(1430));
    layer5_outputs(97) <= not(layer4_outputs(1878));
    layer5_outputs(98) <= not(layer4_outputs(1354)) or (layer4_outputs(1296));
    layer5_outputs(99) <= not(layer4_outputs(211));
    layer5_outputs(100) <= layer4_outputs(1547);
    layer5_outputs(101) <= layer4_outputs(2354);
    layer5_outputs(102) <= (layer4_outputs(629)) xor (layer4_outputs(1696));
    layer5_outputs(103) <= (layer4_outputs(676)) xor (layer4_outputs(2265));
    layer5_outputs(104) <= not((layer4_outputs(2221)) xor (layer4_outputs(1558)));
    layer5_outputs(105) <= layer4_outputs(517);
    layer5_outputs(106) <= not(layer4_outputs(353));
    layer5_outputs(107) <= '0';
    layer5_outputs(108) <= layer4_outputs(1260);
    layer5_outputs(109) <= not((layer4_outputs(437)) xor (layer4_outputs(1025)));
    layer5_outputs(110) <= '0';
    layer5_outputs(111) <= (layer4_outputs(2245)) and not (layer4_outputs(96));
    layer5_outputs(112) <= '1';
    layer5_outputs(113) <= not((layer4_outputs(1776)) and (layer4_outputs(767)));
    layer5_outputs(114) <= not(layer4_outputs(370));
    layer5_outputs(115) <= not((layer4_outputs(430)) and (layer4_outputs(1985)));
    layer5_outputs(116) <= (layer4_outputs(2549)) and (layer4_outputs(2208));
    layer5_outputs(117) <= not(layer4_outputs(1593));
    layer5_outputs(118) <= not(layer4_outputs(1012));
    layer5_outputs(119) <= (layer4_outputs(1223)) and not (layer4_outputs(1331));
    layer5_outputs(120) <= not(layer4_outputs(638));
    layer5_outputs(121) <= layer4_outputs(796);
    layer5_outputs(122) <= not((layer4_outputs(2108)) or (layer4_outputs(543)));
    layer5_outputs(123) <= (layer4_outputs(880)) and not (layer4_outputs(2463));
    layer5_outputs(124) <= not((layer4_outputs(203)) xor (layer4_outputs(1194)));
    layer5_outputs(125) <= (layer4_outputs(455)) and not (layer4_outputs(1700));
    layer5_outputs(126) <= not(layer4_outputs(623));
    layer5_outputs(127) <= (layer4_outputs(1816)) and not (layer4_outputs(1406));
    layer5_outputs(128) <= (layer4_outputs(1557)) and not (layer4_outputs(901));
    layer5_outputs(129) <= not(layer4_outputs(330)) or (layer4_outputs(600));
    layer5_outputs(130) <= not(layer4_outputs(2360));
    layer5_outputs(131) <= layer4_outputs(1841);
    layer5_outputs(132) <= layer4_outputs(753);
    layer5_outputs(133) <= layer4_outputs(577);
    layer5_outputs(134) <= (layer4_outputs(1423)) and not (layer4_outputs(1536));
    layer5_outputs(135) <= not((layer4_outputs(1366)) xor (layer4_outputs(1510)));
    layer5_outputs(136) <= layer4_outputs(434);
    layer5_outputs(137) <= not(layer4_outputs(1051));
    layer5_outputs(138) <= not((layer4_outputs(1167)) xor (layer4_outputs(967)));
    layer5_outputs(139) <= not((layer4_outputs(2121)) xor (layer4_outputs(2352)));
    layer5_outputs(140) <= '0';
    layer5_outputs(141) <= not(layer4_outputs(1805));
    layer5_outputs(142) <= not(layer4_outputs(680)) or (layer4_outputs(1236));
    layer5_outputs(143) <= not(layer4_outputs(1404));
    layer5_outputs(144) <= not(layer4_outputs(1559));
    layer5_outputs(145) <= layer4_outputs(2166);
    layer5_outputs(146) <= layer4_outputs(2355);
    layer5_outputs(147) <= (layer4_outputs(339)) xor (layer4_outputs(1900));
    layer5_outputs(148) <= layer4_outputs(142);
    layer5_outputs(149) <= layer4_outputs(256);
    layer5_outputs(150) <= layer4_outputs(1172);
    layer5_outputs(151) <= layer4_outputs(1336);
    layer5_outputs(152) <= not((layer4_outputs(1629)) or (layer4_outputs(255)));
    layer5_outputs(153) <= not(layer4_outputs(2103)) or (layer4_outputs(6));
    layer5_outputs(154) <= layer4_outputs(1081);
    layer5_outputs(155) <= not(layer4_outputs(744));
    layer5_outputs(156) <= not((layer4_outputs(1023)) or (layer4_outputs(2364)));
    layer5_outputs(157) <= (layer4_outputs(1872)) or (layer4_outputs(2151));
    layer5_outputs(158) <= not(layer4_outputs(2485));
    layer5_outputs(159) <= (layer4_outputs(1002)) and (layer4_outputs(1312));
    layer5_outputs(160) <= not(layer4_outputs(549)) or (layer4_outputs(364));
    layer5_outputs(161) <= (layer4_outputs(367)) or (layer4_outputs(305));
    layer5_outputs(162) <= '0';
    layer5_outputs(163) <= (layer4_outputs(889)) and not (layer4_outputs(540));
    layer5_outputs(164) <= (layer4_outputs(1274)) and (layer4_outputs(385));
    layer5_outputs(165) <= layer4_outputs(1783);
    layer5_outputs(166) <= (layer4_outputs(115)) and not (layer4_outputs(2025));
    layer5_outputs(167) <= not((layer4_outputs(1911)) and (layer4_outputs(1818)));
    layer5_outputs(168) <= layer4_outputs(1398);
    layer5_outputs(169) <= not((layer4_outputs(504)) xor (layer4_outputs(66)));
    layer5_outputs(170) <= not((layer4_outputs(2264)) or (layer4_outputs(2259)));
    layer5_outputs(171) <= not(layer4_outputs(2191)) or (layer4_outputs(117));
    layer5_outputs(172) <= not((layer4_outputs(929)) or (layer4_outputs(412)));
    layer5_outputs(173) <= layer4_outputs(1638);
    layer5_outputs(174) <= '1';
    layer5_outputs(175) <= layer4_outputs(569);
    layer5_outputs(176) <= not(layer4_outputs(2401));
    layer5_outputs(177) <= not((layer4_outputs(2502)) xor (layer4_outputs(446)));
    layer5_outputs(178) <= layer4_outputs(2546);
    layer5_outputs(179) <= (layer4_outputs(787)) and not (layer4_outputs(260));
    layer5_outputs(180) <= not(layer4_outputs(2473));
    layer5_outputs(181) <= (layer4_outputs(586)) or (layer4_outputs(481));
    layer5_outputs(182) <= not(layer4_outputs(1946));
    layer5_outputs(183) <= not((layer4_outputs(181)) xor (layer4_outputs(624)));
    layer5_outputs(184) <= layer4_outputs(2073);
    layer5_outputs(185) <= not(layer4_outputs(167));
    layer5_outputs(186) <= (layer4_outputs(894)) and (layer4_outputs(759));
    layer5_outputs(187) <= not(layer4_outputs(2197)) or (layer4_outputs(1602));
    layer5_outputs(188) <= not(layer4_outputs(316));
    layer5_outputs(189) <= not(layer4_outputs(1527)) or (layer4_outputs(779));
    layer5_outputs(190) <= not(layer4_outputs(219));
    layer5_outputs(191) <= layer4_outputs(1692);
    layer5_outputs(192) <= layer4_outputs(1102);
    layer5_outputs(193) <= (layer4_outputs(2327)) and (layer4_outputs(2558));
    layer5_outputs(194) <= not((layer4_outputs(1777)) xor (layer4_outputs(389)));
    layer5_outputs(195) <= not(layer4_outputs(2180)) or (layer4_outputs(535));
    layer5_outputs(196) <= (layer4_outputs(1448)) xor (layer4_outputs(1163));
    layer5_outputs(197) <= not(layer4_outputs(914));
    layer5_outputs(198) <= not(layer4_outputs(1967));
    layer5_outputs(199) <= layer4_outputs(346);
    layer5_outputs(200) <= (layer4_outputs(1093)) or (layer4_outputs(137));
    layer5_outputs(201) <= (layer4_outputs(203)) and (layer4_outputs(1961));
    layer5_outputs(202) <= not(layer4_outputs(488)) or (layer4_outputs(1327));
    layer5_outputs(203) <= '1';
    layer5_outputs(204) <= layer4_outputs(2296);
    layer5_outputs(205) <= layer4_outputs(459);
    layer5_outputs(206) <= layer4_outputs(1988);
    layer5_outputs(207) <= (layer4_outputs(82)) and not (layer4_outputs(355));
    layer5_outputs(208) <= not(layer4_outputs(2282));
    layer5_outputs(209) <= not(layer4_outputs(1698));
    layer5_outputs(210) <= layer4_outputs(2276);
    layer5_outputs(211) <= layer4_outputs(153);
    layer5_outputs(212) <= not(layer4_outputs(1847)) or (layer4_outputs(2013));
    layer5_outputs(213) <= not(layer4_outputs(1466));
    layer5_outputs(214) <= (layer4_outputs(2390)) and not (layer4_outputs(1833));
    layer5_outputs(215) <= not(layer4_outputs(474)) or (layer4_outputs(2150));
    layer5_outputs(216) <= layer4_outputs(2425);
    layer5_outputs(217) <= (layer4_outputs(2164)) or (layer4_outputs(908));
    layer5_outputs(218) <= not(layer4_outputs(2311)) or (layer4_outputs(70));
    layer5_outputs(219) <= not(layer4_outputs(709));
    layer5_outputs(220) <= not(layer4_outputs(1779));
    layer5_outputs(221) <= layer4_outputs(675);
    layer5_outputs(222) <= (layer4_outputs(2183)) xor (layer4_outputs(1997));
    layer5_outputs(223) <= not(layer4_outputs(1321)) or (layer4_outputs(1951));
    layer5_outputs(224) <= not(layer4_outputs(2456)) or (layer4_outputs(1029));
    layer5_outputs(225) <= not((layer4_outputs(1710)) and (layer4_outputs(963)));
    layer5_outputs(226) <= (layer4_outputs(1537)) and not (layer4_outputs(2476));
    layer5_outputs(227) <= not(layer4_outputs(1065));
    layer5_outputs(228) <= not(layer4_outputs(1555));
    layer5_outputs(229) <= not(layer4_outputs(2543));
    layer5_outputs(230) <= layer4_outputs(617);
    layer5_outputs(231) <= layer4_outputs(1652);
    layer5_outputs(232) <= '1';
    layer5_outputs(233) <= layer4_outputs(433);
    layer5_outputs(234) <= not((layer4_outputs(703)) or (layer4_outputs(799)));
    layer5_outputs(235) <= (layer4_outputs(2442)) xor (layer4_outputs(1149));
    layer5_outputs(236) <= not(layer4_outputs(2152));
    layer5_outputs(237) <= layer4_outputs(1814);
    layer5_outputs(238) <= not(layer4_outputs(2431)) or (layer4_outputs(719));
    layer5_outputs(239) <= layer4_outputs(136);
    layer5_outputs(240) <= (layer4_outputs(853)) and (layer4_outputs(1066));
    layer5_outputs(241) <= (layer4_outputs(1245)) and (layer4_outputs(1090));
    layer5_outputs(242) <= layer4_outputs(246);
    layer5_outputs(243) <= not(layer4_outputs(837)) or (layer4_outputs(2047));
    layer5_outputs(244) <= (layer4_outputs(1730)) and not (layer4_outputs(2533));
    layer5_outputs(245) <= layer4_outputs(750);
    layer5_outputs(246) <= not(layer4_outputs(2552)) or (layer4_outputs(1418));
    layer5_outputs(247) <= layer4_outputs(882);
    layer5_outputs(248) <= not(layer4_outputs(1254));
    layer5_outputs(249) <= layer4_outputs(1996);
    layer5_outputs(250) <= not(layer4_outputs(702)) or (layer4_outputs(353));
    layer5_outputs(251) <= (layer4_outputs(1027)) and (layer4_outputs(1743));
    layer5_outputs(252) <= (layer4_outputs(1424)) or (layer4_outputs(2321));
    layer5_outputs(253) <= not((layer4_outputs(2227)) or (layer4_outputs(186)));
    layer5_outputs(254) <= not((layer4_outputs(431)) or (layer4_outputs(465)));
    layer5_outputs(255) <= layer4_outputs(2015);
    layer5_outputs(256) <= not(layer4_outputs(2315));
    layer5_outputs(257) <= not(layer4_outputs(2392)) or (layer4_outputs(533));
    layer5_outputs(258) <= layer4_outputs(2548);
    layer5_outputs(259) <= (layer4_outputs(1192)) xor (layer4_outputs(1717));
    layer5_outputs(260) <= (layer4_outputs(1608)) xor (layer4_outputs(973));
    layer5_outputs(261) <= not(layer4_outputs(2164));
    layer5_outputs(262) <= layer4_outputs(1994);
    layer5_outputs(263) <= (layer4_outputs(1168)) and not (layer4_outputs(654));
    layer5_outputs(264) <= (layer4_outputs(837)) and not (layer4_outputs(1797));
    layer5_outputs(265) <= '1';
    layer5_outputs(266) <= not((layer4_outputs(50)) and (layer4_outputs(1653)));
    layer5_outputs(267) <= not((layer4_outputs(396)) xor (layer4_outputs(782)));
    layer5_outputs(268) <= (layer4_outputs(1272)) and (layer4_outputs(2279));
    layer5_outputs(269) <= layer4_outputs(1543);
    layer5_outputs(270) <= layer4_outputs(1957);
    layer5_outputs(271) <= layer4_outputs(909);
    layer5_outputs(272) <= '1';
    layer5_outputs(273) <= not(layer4_outputs(476));
    layer5_outputs(274) <= (layer4_outputs(1629)) and (layer4_outputs(257));
    layer5_outputs(275) <= not(layer4_outputs(971));
    layer5_outputs(276) <= not(layer4_outputs(1142));
    layer5_outputs(277) <= '0';
    layer5_outputs(278) <= '1';
    layer5_outputs(279) <= layer4_outputs(2198);
    layer5_outputs(280) <= not((layer4_outputs(2075)) or (layer4_outputs(2533)));
    layer5_outputs(281) <= layer4_outputs(301);
    layer5_outputs(282) <= layer4_outputs(953);
    layer5_outputs(283) <= (layer4_outputs(2098)) and not (layer4_outputs(2428));
    layer5_outputs(284) <= layer4_outputs(479);
    layer5_outputs(285) <= (layer4_outputs(1061)) xor (layer4_outputs(847));
    layer5_outputs(286) <= not(layer4_outputs(2205));
    layer5_outputs(287) <= layer4_outputs(1013);
    layer5_outputs(288) <= not(layer4_outputs(2008)) or (layer4_outputs(1631));
    layer5_outputs(289) <= layer4_outputs(2154);
    layer5_outputs(290) <= layer4_outputs(1816);
    layer5_outputs(291) <= layer4_outputs(1910);
    layer5_outputs(292) <= not(layer4_outputs(2363)) or (layer4_outputs(974));
    layer5_outputs(293) <= not(layer4_outputs(1188));
    layer5_outputs(294) <= not((layer4_outputs(202)) and (layer4_outputs(321)));
    layer5_outputs(295) <= (layer4_outputs(770)) and not (layer4_outputs(2281));
    layer5_outputs(296) <= not(layer4_outputs(621));
    layer5_outputs(297) <= (layer4_outputs(672)) xor (layer4_outputs(1487));
    layer5_outputs(298) <= (layer4_outputs(235)) and not (layer4_outputs(1377));
    layer5_outputs(299) <= layer4_outputs(2182);
    layer5_outputs(300) <= (layer4_outputs(805)) or (layer4_outputs(938));
    layer5_outputs(301) <= not(layer4_outputs(976)) or (layer4_outputs(1068));
    layer5_outputs(302) <= not((layer4_outputs(938)) and (layer4_outputs(1198)));
    layer5_outputs(303) <= not(layer4_outputs(1129)) or (layer4_outputs(1395));
    layer5_outputs(304) <= layer4_outputs(529);
    layer5_outputs(305) <= layer4_outputs(566);
    layer5_outputs(306) <= not(layer4_outputs(1050));
    layer5_outputs(307) <= layer4_outputs(1686);
    layer5_outputs(308) <= not(layer4_outputs(2133));
    layer5_outputs(309) <= layer4_outputs(67);
    layer5_outputs(310) <= (layer4_outputs(1341)) and not (layer4_outputs(2250));
    layer5_outputs(311) <= (layer4_outputs(442)) and (layer4_outputs(2401));
    layer5_outputs(312) <= '0';
    layer5_outputs(313) <= '0';
    layer5_outputs(314) <= not(layer4_outputs(1688)) or (layer4_outputs(43));
    layer5_outputs(315) <= '1';
    layer5_outputs(316) <= not(layer4_outputs(375)) or (layer4_outputs(123));
    layer5_outputs(317) <= not(layer4_outputs(1032));
    layer5_outputs(318) <= layer4_outputs(1407);
    layer5_outputs(319) <= not((layer4_outputs(257)) xor (layer4_outputs(1403)));
    layer5_outputs(320) <= layer4_outputs(313);
    layer5_outputs(321) <= (layer4_outputs(2444)) and not (layer4_outputs(2524));
    layer5_outputs(322) <= not(layer4_outputs(2101));
    layer5_outputs(323) <= layer4_outputs(33);
    layer5_outputs(324) <= not(layer4_outputs(788)) or (layer4_outputs(1008));
    layer5_outputs(325) <= not((layer4_outputs(1216)) or (layer4_outputs(2294)));
    layer5_outputs(326) <= (layer4_outputs(1650)) and not (layer4_outputs(1690));
    layer5_outputs(327) <= not((layer4_outputs(1108)) and (layer4_outputs(1632)));
    layer5_outputs(328) <= layer4_outputs(1265);
    layer5_outputs(329) <= layer4_outputs(2074);
    layer5_outputs(330) <= not((layer4_outputs(786)) or (layer4_outputs(1905)));
    layer5_outputs(331) <= layer4_outputs(1411);
    layer5_outputs(332) <= '0';
    layer5_outputs(333) <= layer4_outputs(220);
    layer5_outputs(334) <= not(layer4_outputs(224)) or (layer4_outputs(2375));
    layer5_outputs(335) <= not(layer4_outputs(822));
    layer5_outputs(336) <= layer4_outputs(1482);
    layer5_outputs(337) <= layer4_outputs(2305);
    layer5_outputs(338) <= layer4_outputs(2074);
    layer5_outputs(339) <= not(layer4_outputs(2387)) or (layer4_outputs(2041));
    layer5_outputs(340) <= '0';
    layer5_outputs(341) <= not((layer4_outputs(1584)) or (layer4_outputs(1387)));
    layer5_outputs(342) <= (layer4_outputs(885)) or (layer4_outputs(2471));
    layer5_outputs(343) <= not(layer4_outputs(640));
    layer5_outputs(344) <= layer4_outputs(945);
    layer5_outputs(345) <= (layer4_outputs(957)) and not (layer4_outputs(936));
    layer5_outputs(346) <= not(layer4_outputs(1275));
    layer5_outputs(347) <= not(layer4_outputs(1232));
    layer5_outputs(348) <= layer4_outputs(1034);
    layer5_outputs(349) <= layer4_outputs(821);
    layer5_outputs(350) <= layer4_outputs(243);
    layer5_outputs(351) <= (layer4_outputs(29)) and not (layer4_outputs(2330));
    layer5_outputs(352) <= (layer4_outputs(1020)) and (layer4_outputs(307));
    layer5_outputs(353) <= not(layer4_outputs(704));
    layer5_outputs(354) <= not((layer4_outputs(208)) or (layer4_outputs(183)));
    layer5_outputs(355) <= layer4_outputs(2165);
    layer5_outputs(356) <= (layer4_outputs(1301)) and not (layer4_outputs(492));
    layer5_outputs(357) <= (layer4_outputs(1823)) and not (layer4_outputs(1521));
    layer5_outputs(358) <= not(layer4_outputs(810)) or (layer4_outputs(2052));
    layer5_outputs(359) <= not(layer4_outputs(518)) or (layer4_outputs(1563));
    layer5_outputs(360) <= not((layer4_outputs(1812)) and (layer4_outputs(1018)));
    layer5_outputs(361) <= not((layer4_outputs(1002)) xor (layer4_outputs(1494)));
    layer5_outputs(362) <= not(layer4_outputs(1863)) or (layer4_outputs(1084));
    layer5_outputs(363) <= (layer4_outputs(1775)) or (layer4_outputs(1357));
    layer5_outputs(364) <= not(layer4_outputs(1752));
    layer5_outputs(365) <= not(layer4_outputs(735)) or (layer4_outputs(2186));
    layer5_outputs(366) <= not(layer4_outputs(973));
    layer5_outputs(367) <= layer4_outputs(722);
    layer5_outputs(368) <= not(layer4_outputs(2079));
    layer5_outputs(369) <= not((layer4_outputs(1612)) or (layer4_outputs(2520)));
    layer5_outputs(370) <= layer4_outputs(121);
    layer5_outputs(371) <= '0';
    layer5_outputs(372) <= not(layer4_outputs(296));
    layer5_outputs(373) <= not(layer4_outputs(509)) or (layer4_outputs(2334));
    layer5_outputs(374) <= not(layer4_outputs(254));
    layer5_outputs(375) <= not((layer4_outputs(2432)) and (layer4_outputs(493)));
    layer5_outputs(376) <= layer4_outputs(941);
    layer5_outputs(377) <= not(layer4_outputs(2079));
    layer5_outputs(378) <= not(layer4_outputs(1203));
    layer5_outputs(379) <= not((layer4_outputs(256)) or (layer4_outputs(222)));
    layer5_outputs(380) <= not(layer4_outputs(2158));
    layer5_outputs(381) <= (layer4_outputs(2282)) and not (layer4_outputs(1517));
    layer5_outputs(382) <= not(layer4_outputs(378));
    layer5_outputs(383) <= (layer4_outputs(524)) and not (layer4_outputs(854));
    layer5_outputs(384) <= not(layer4_outputs(553));
    layer5_outputs(385) <= not(layer4_outputs(2518));
    layer5_outputs(386) <= layer4_outputs(2215);
    layer5_outputs(387) <= (layer4_outputs(2402)) and (layer4_outputs(379));
    layer5_outputs(388) <= not(layer4_outputs(2505));
    layer5_outputs(389) <= (layer4_outputs(2028)) xor (layer4_outputs(274));
    layer5_outputs(390) <= (layer4_outputs(1127)) and not (layer4_outputs(1031));
    layer5_outputs(391) <= not(layer4_outputs(1574));
    layer5_outputs(392) <= not(layer4_outputs(841)) or (layer4_outputs(177));
    layer5_outputs(393) <= not(layer4_outputs(266));
    layer5_outputs(394) <= layer4_outputs(2489);
    layer5_outputs(395) <= not(layer4_outputs(421)) or (layer4_outputs(2225));
    layer5_outputs(396) <= layer4_outputs(1531);
    layer5_outputs(397) <= not((layer4_outputs(123)) xor (layer4_outputs(769)));
    layer5_outputs(398) <= not(layer4_outputs(1307)) or (layer4_outputs(2290));
    layer5_outputs(399) <= (layer4_outputs(440)) and not (layer4_outputs(601));
    layer5_outputs(400) <= not(layer4_outputs(531));
    layer5_outputs(401) <= not(layer4_outputs(891));
    layer5_outputs(402) <= not((layer4_outputs(1049)) xor (layer4_outputs(1684)));
    layer5_outputs(403) <= not(layer4_outputs(1431));
    layer5_outputs(404) <= (layer4_outputs(1287)) or (layer4_outputs(656));
    layer5_outputs(405) <= not((layer4_outputs(956)) or (layer4_outputs(1270)));
    layer5_outputs(406) <= layer4_outputs(1860);
    layer5_outputs(407) <= not(layer4_outputs(2035)) or (layer4_outputs(2391));
    layer5_outputs(408) <= (layer4_outputs(720)) and (layer4_outputs(1839));
    layer5_outputs(409) <= layer4_outputs(1245);
    layer5_outputs(410) <= layer4_outputs(250);
    layer5_outputs(411) <= (layer4_outputs(1970)) xor (layer4_outputs(1004));
    layer5_outputs(412) <= not(layer4_outputs(2068));
    layer5_outputs(413) <= layer4_outputs(2249);
    layer5_outputs(414) <= not(layer4_outputs(270));
    layer5_outputs(415) <= (layer4_outputs(1355)) or (layer4_outputs(62));
    layer5_outputs(416) <= not(layer4_outputs(1061));
    layer5_outputs(417) <= not(layer4_outputs(2498));
    layer5_outputs(418) <= not((layer4_outputs(2516)) and (layer4_outputs(491)));
    layer5_outputs(419) <= not(layer4_outputs(295)) or (layer4_outputs(1708));
    layer5_outputs(420) <= (layer4_outputs(1589)) xor (layer4_outputs(1749));
    layer5_outputs(421) <= (layer4_outputs(734)) and (layer4_outputs(844));
    layer5_outputs(422) <= layer4_outputs(901);
    layer5_outputs(423) <= not(layer4_outputs(1567)) or (layer4_outputs(2133));
    layer5_outputs(424) <= (layer4_outputs(1647)) and (layer4_outputs(1823));
    layer5_outputs(425) <= not(layer4_outputs(813));
    layer5_outputs(426) <= (layer4_outputs(776)) or (layer4_outputs(660));
    layer5_outputs(427) <= '0';
    layer5_outputs(428) <= not(layer4_outputs(1062));
    layer5_outputs(429) <= (layer4_outputs(1228)) and not (layer4_outputs(1356));
    layer5_outputs(430) <= not((layer4_outputs(1743)) or (layer4_outputs(171)));
    layer5_outputs(431) <= layer4_outputs(675);
    layer5_outputs(432) <= (layer4_outputs(1431)) and (layer4_outputs(1906));
    layer5_outputs(433) <= '1';
    layer5_outputs(434) <= not(layer4_outputs(2427));
    layer5_outputs(435) <= layer4_outputs(2436);
    layer5_outputs(436) <= (layer4_outputs(655)) xor (layer4_outputs(354));
    layer5_outputs(437) <= not(layer4_outputs(1728));
    layer5_outputs(438) <= (layer4_outputs(1258)) or (layer4_outputs(66));
    layer5_outputs(439) <= not(layer4_outputs(584));
    layer5_outputs(440) <= '1';
    layer5_outputs(441) <= layer4_outputs(2240);
    layer5_outputs(442) <= (layer4_outputs(1549)) and not (layer4_outputs(1442));
    layer5_outputs(443) <= not(layer4_outputs(1372));
    layer5_outputs(444) <= layer4_outputs(1094);
    layer5_outputs(445) <= '1';
    layer5_outputs(446) <= not((layer4_outputs(1216)) and (layer4_outputs(2398)));
    layer5_outputs(447) <= (layer4_outputs(1361)) and not (layer4_outputs(1224));
    layer5_outputs(448) <= not(layer4_outputs(871)) or (layer4_outputs(1394));
    layer5_outputs(449) <= layer4_outputs(768);
    layer5_outputs(450) <= '0';
    layer5_outputs(451) <= not(layer4_outputs(1360)) or (layer4_outputs(13));
    layer5_outputs(452) <= not(layer4_outputs(1862));
    layer5_outputs(453) <= layer4_outputs(1452);
    layer5_outputs(454) <= (layer4_outputs(1990)) and (layer4_outputs(1277));
    layer5_outputs(455) <= not(layer4_outputs(274));
    layer5_outputs(456) <= (layer4_outputs(492)) or (layer4_outputs(947));
    layer5_outputs(457) <= not(layer4_outputs(2240));
    layer5_outputs(458) <= not((layer4_outputs(2465)) xor (layer4_outputs(443)));
    layer5_outputs(459) <= not(layer4_outputs(910));
    layer5_outputs(460) <= not((layer4_outputs(93)) and (layer4_outputs(564)));
    layer5_outputs(461) <= (layer4_outputs(1385)) and not (layer4_outputs(2223));
    layer5_outputs(462) <= '0';
    layer5_outputs(463) <= layer4_outputs(1705);
    layer5_outputs(464) <= not(layer4_outputs(534));
    layer5_outputs(465) <= layer4_outputs(607);
    layer5_outputs(466) <= not(layer4_outputs(1939)) or (layer4_outputs(1175));
    layer5_outputs(467) <= layer4_outputs(1151);
    layer5_outputs(468) <= not((layer4_outputs(900)) and (layer4_outputs(2117)));
    layer5_outputs(469) <= not(layer4_outputs(884));
    layer5_outputs(470) <= not(layer4_outputs(463));
    layer5_outputs(471) <= not(layer4_outputs(318));
    layer5_outputs(472) <= not(layer4_outputs(438));
    layer5_outputs(473) <= not(layer4_outputs(1739));
    layer5_outputs(474) <= not((layer4_outputs(2345)) or (layer4_outputs(534)));
    layer5_outputs(475) <= not(layer4_outputs(2483));
    layer5_outputs(476) <= layer4_outputs(1043);
    layer5_outputs(477) <= not((layer4_outputs(1239)) or (layer4_outputs(33)));
    layer5_outputs(478) <= not(layer4_outputs(1750));
    layer5_outputs(479) <= not(layer4_outputs(919)) or (layer4_outputs(1038));
    layer5_outputs(480) <= (layer4_outputs(1290)) or (layer4_outputs(1822));
    layer5_outputs(481) <= (layer4_outputs(338)) or (layer4_outputs(457));
    layer5_outputs(482) <= (layer4_outputs(2472)) and not (layer4_outputs(2410));
    layer5_outputs(483) <= layer4_outputs(1501);
    layer5_outputs(484) <= layer4_outputs(297);
    layer5_outputs(485) <= layer4_outputs(2329);
    layer5_outputs(486) <= not(layer4_outputs(280)) or (layer4_outputs(395));
    layer5_outputs(487) <= (layer4_outputs(962)) and not (layer4_outputs(1197));
    layer5_outputs(488) <= not(layer4_outputs(1160)) or (layer4_outputs(2372));
    layer5_outputs(489) <= (layer4_outputs(1374)) xor (layer4_outputs(87));
    layer5_outputs(490) <= not((layer4_outputs(2167)) xor (layer4_outputs(483)));
    layer5_outputs(491) <= (layer4_outputs(1258)) or (layer4_outputs(1407));
    layer5_outputs(492) <= (layer4_outputs(119)) or (layer4_outputs(280));
    layer5_outputs(493) <= not(layer4_outputs(697));
    layer5_outputs(494) <= not((layer4_outputs(1626)) xor (layer4_outputs(133)));
    layer5_outputs(495) <= not(layer4_outputs(390));
    layer5_outputs(496) <= not(layer4_outputs(345));
    layer5_outputs(497) <= not(layer4_outputs(611));
    layer5_outputs(498) <= not(layer4_outputs(1508)) or (layer4_outputs(2518));
    layer5_outputs(499) <= not(layer4_outputs(902));
    layer5_outputs(500) <= not(layer4_outputs(1680));
    layer5_outputs(501) <= layer4_outputs(633);
    layer5_outputs(502) <= (layer4_outputs(2332)) or (layer4_outputs(1021));
    layer5_outputs(503) <= not(layer4_outputs(1937));
    layer5_outputs(504) <= (layer4_outputs(1056)) xor (layer4_outputs(1809));
    layer5_outputs(505) <= layer4_outputs(774);
    layer5_outputs(506) <= not(layer4_outputs(760));
    layer5_outputs(507) <= '1';
    layer5_outputs(508) <= not(layer4_outputs(1539));
    layer5_outputs(509) <= layer4_outputs(2021);
    layer5_outputs(510) <= (layer4_outputs(749)) and not (layer4_outputs(969));
    layer5_outputs(511) <= not(layer4_outputs(1897));
    layer5_outputs(512) <= not(layer4_outputs(2137)) or (layer4_outputs(864));
    layer5_outputs(513) <= not(layer4_outputs(1535));
    layer5_outputs(514) <= layer4_outputs(631);
    layer5_outputs(515) <= not((layer4_outputs(2343)) xor (layer4_outputs(1035)));
    layer5_outputs(516) <= layer4_outputs(2065);
    layer5_outputs(517) <= not((layer4_outputs(1089)) and (layer4_outputs(1602)));
    layer5_outputs(518) <= layer4_outputs(415);
    layer5_outputs(519) <= not((layer4_outputs(1801)) or (layer4_outputs(1711)));
    layer5_outputs(520) <= (layer4_outputs(1630)) xor (layer4_outputs(9));
    layer5_outputs(521) <= (layer4_outputs(1981)) and not (layer4_outputs(1097));
    layer5_outputs(522) <= (layer4_outputs(1311)) or (layer4_outputs(1902));
    layer5_outputs(523) <= not(layer4_outputs(1573));
    layer5_outputs(524) <= (layer4_outputs(1438)) and not (layer4_outputs(468));
    layer5_outputs(525) <= layer4_outputs(351);
    layer5_outputs(526) <= layer4_outputs(683);
    layer5_outputs(527) <= not(layer4_outputs(1963));
    layer5_outputs(528) <= layer4_outputs(550);
    layer5_outputs(529) <= not((layer4_outputs(1893)) or (layer4_outputs(1698)));
    layer5_outputs(530) <= layer4_outputs(581);
    layer5_outputs(531) <= (layer4_outputs(1786)) and (layer4_outputs(1917));
    layer5_outputs(532) <= not(layer4_outputs(366));
    layer5_outputs(533) <= (layer4_outputs(1913)) and (layer4_outputs(2056));
    layer5_outputs(534) <= not(layer4_outputs(2342));
    layer5_outputs(535) <= (layer4_outputs(1386)) and (layer4_outputs(737));
    layer5_outputs(536) <= (layer4_outputs(2550)) and not (layer4_outputs(2123));
    layer5_outputs(537) <= (layer4_outputs(190)) or (layer4_outputs(1274));
    layer5_outputs(538) <= not(layer4_outputs(246));
    layer5_outputs(539) <= layer4_outputs(2495);
    layer5_outputs(540) <= layer4_outputs(744);
    layer5_outputs(541) <= not(layer4_outputs(1264)) or (layer4_outputs(681));
    layer5_outputs(542) <= (layer4_outputs(76)) and not (layer4_outputs(496));
    layer5_outputs(543) <= layer4_outputs(526);
    layer5_outputs(544) <= (layer4_outputs(1488)) or (layer4_outputs(531));
    layer5_outputs(545) <= not((layer4_outputs(1859)) or (layer4_outputs(2012)));
    layer5_outputs(546) <= not((layer4_outputs(1482)) or (layer4_outputs(991)));
    layer5_outputs(547) <= layer4_outputs(1530);
    layer5_outputs(548) <= '0';
    layer5_outputs(549) <= (layer4_outputs(1195)) and not (layer4_outputs(283));
    layer5_outputs(550) <= not(layer4_outputs(1150));
    layer5_outputs(551) <= not(layer4_outputs(159)) or (layer4_outputs(918));
    layer5_outputs(552) <= layer4_outputs(2000);
    layer5_outputs(553) <= not(layer4_outputs(595));
    layer5_outputs(554) <= not((layer4_outputs(2552)) or (layer4_outputs(6)));
    layer5_outputs(555) <= not(layer4_outputs(2116));
    layer5_outputs(556) <= '0';
    layer5_outputs(557) <= not(layer4_outputs(968));
    layer5_outputs(558) <= not(layer4_outputs(1232));
    layer5_outputs(559) <= (layer4_outputs(1634)) xor (layer4_outputs(119));
    layer5_outputs(560) <= not(layer4_outputs(1417));
    layer5_outputs(561) <= (layer4_outputs(858)) xor (layer4_outputs(573));
    layer5_outputs(562) <= layer4_outputs(1802);
    layer5_outputs(563) <= layer4_outputs(2526);
    layer5_outputs(564) <= not(layer4_outputs(1951));
    layer5_outputs(565) <= not(layer4_outputs(1028));
    layer5_outputs(566) <= not(layer4_outputs(91));
    layer5_outputs(567) <= layer4_outputs(2486);
    layer5_outputs(568) <= not(layer4_outputs(2196)) or (layer4_outputs(1009));
    layer5_outputs(569) <= (layer4_outputs(176)) and (layer4_outputs(24));
    layer5_outputs(570) <= (layer4_outputs(2080)) and not (layer4_outputs(2202));
    layer5_outputs(571) <= layer4_outputs(1204);
    layer5_outputs(572) <= not(layer4_outputs(2335));
    layer5_outputs(573) <= not((layer4_outputs(1681)) xor (layer4_outputs(2234)));
    layer5_outputs(574) <= not((layer4_outputs(324)) and (layer4_outputs(2042)));
    layer5_outputs(575) <= layer4_outputs(2481);
    layer5_outputs(576) <= not(layer4_outputs(2273)) or (layer4_outputs(1826));
    layer5_outputs(577) <= not(layer4_outputs(1545));
    layer5_outputs(578) <= layer4_outputs(1500);
    layer5_outputs(579) <= (layer4_outputs(1646)) and (layer4_outputs(664));
    layer5_outputs(580) <= not(layer4_outputs(2214)) or (layer4_outputs(170));
    layer5_outputs(581) <= layer4_outputs(2479);
    layer5_outputs(582) <= '0';
    layer5_outputs(583) <= layer4_outputs(565);
    layer5_outputs(584) <= layer4_outputs(1382);
    layer5_outputs(585) <= (layer4_outputs(602)) and not (layer4_outputs(904));
    layer5_outputs(586) <= (layer4_outputs(2159)) and (layer4_outputs(1762));
    layer5_outputs(587) <= not(layer4_outputs(2386));
    layer5_outputs(588) <= not((layer4_outputs(1773)) and (layer4_outputs(1163)));
    layer5_outputs(589) <= layer4_outputs(1376);
    layer5_outputs(590) <= layer4_outputs(39);
    layer5_outputs(591) <= (layer4_outputs(1525)) xor (layer4_outputs(1452));
    layer5_outputs(592) <= '0';
    layer5_outputs(593) <= not(layer4_outputs(1875)) or (layer4_outputs(2292));
    layer5_outputs(594) <= not(layer4_outputs(2403));
    layer5_outputs(595) <= not(layer4_outputs(999)) or (layer4_outputs(2326));
    layer5_outputs(596) <= (layer4_outputs(1858)) and not (layer4_outputs(368));
    layer5_outputs(597) <= '0';
    layer5_outputs(598) <= (layer4_outputs(1445)) and not (layer4_outputs(657));
    layer5_outputs(599) <= layer4_outputs(1549);
    layer5_outputs(600) <= not(layer4_outputs(1665));
    layer5_outputs(601) <= not((layer4_outputs(1553)) xor (layer4_outputs(1726)));
    layer5_outputs(602) <= not(layer4_outputs(1157));
    layer5_outputs(603) <= (layer4_outputs(1478)) and (layer4_outputs(215));
    layer5_outputs(604) <= (layer4_outputs(38)) and not (layer4_outputs(1014));
    layer5_outputs(605) <= layer4_outputs(122);
    layer5_outputs(606) <= not((layer4_outputs(896)) and (layer4_outputs(579)));
    layer5_outputs(607) <= layer4_outputs(1599);
    layer5_outputs(608) <= not((layer4_outputs(2287)) and (layer4_outputs(1209)));
    layer5_outputs(609) <= not((layer4_outputs(477)) or (layer4_outputs(580)));
    layer5_outputs(610) <= '0';
    layer5_outputs(611) <= layer4_outputs(135);
    layer5_outputs(612) <= layer4_outputs(1131);
    layer5_outputs(613) <= not(layer4_outputs(34));
    layer5_outputs(614) <= not(layer4_outputs(986));
    layer5_outputs(615) <= layer4_outputs(1921);
    layer5_outputs(616) <= (layer4_outputs(2140)) or (layer4_outputs(436));
    layer5_outputs(617) <= not(layer4_outputs(791));
    layer5_outputs(618) <= not((layer4_outputs(920)) xor (layer4_outputs(1745)));
    layer5_outputs(619) <= layer4_outputs(1881);
    layer5_outputs(620) <= layer4_outputs(547);
    layer5_outputs(621) <= (layer4_outputs(1399)) and not (layer4_outputs(184));
    layer5_outputs(622) <= not(layer4_outputs(1017)) or (layer4_outputs(1445));
    layer5_outputs(623) <= (layer4_outputs(2506)) and not (layer4_outputs(2402));
    layer5_outputs(624) <= not(layer4_outputs(933));
    layer5_outputs(625) <= not(layer4_outputs(1242));
    layer5_outputs(626) <= not(layer4_outputs(1003));
    layer5_outputs(627) <= not((layer4_outputs(2090)) or (layer4_outputs(1559)));
    layer5_outputs(628) <= not((layer4_outputs(2135)) xor (layer4_outputs(150)));
    layer5_outputs(629) <= not((layer4_outputs(1409)) xor (layer4_outputs(336)));
    layer5_outputs(630) <= '1';
    layer5_outputs(631) <= not((layer4_outputs(71)) or (layer4_outputs(1520)));
    layer5_outputs(632) <= not(layer4_outputs(2118));
    layer5_outputs(633) <= not(layer4_outputs(948)) or (layer4_outputs(149));
    layer5_outputs(634) <= not(layer4_outputs(1781)) or (layer4_outputs(1097));
    layer5_outputs(635) <= (layer4_outputs(495)) and (layer4_outputs(1920));
    layer5_outputs(636) <= layer4_outputs(845);
    layer5_outputs(637) <= (layer4_outputs(1975)) and not (layer4_outputs(49));
    layer5_outputs(638) <= (layer4_outputs(35)) xor (layer4_outputs(1531));
    layer5_outputs(639) <= not((layer4_outputs(1266)) xor (layer4_outputs(578)));
    layer5_outputs(640) <= not(layer4_outputs(2447));
    layer5_outputs(641) <= layer4_outputs(1595);
    layer5_outputs(642) <= not(layer4_outputs(805));
    layer5_outputs(643) <= not(layer4_outputs(2232));
    layer5_outputs(644) <= '0';
    layer5_outputs(645) <= not(layer4_outputs(670)) or (layer4_outputs(1092));
    layer5_outputs(646) <= layer4_outputs(1576);
    layer5_outputs(647) <= (layer4_outputs(1268)) and (layer4_outputs(1558));
    layer5_outputs(648) <= not(layer4_outputs(72)) or (layer4_outputs(621));
    layer5_outputs(649) <= not(layer4_outputs(2146)) or (layer4_outputs(1294));
    layer5_outputs(650) <= not(layer4_outputs(2491)) or (layer4_outputs(1396));
    layer5_outputs(651) <= not(layer4_outputs(800)) or (layer4_outputs(1851));
    layer5_outputs(652) <= not(layer4_outputs(427));
    layer5_outputs(653) <= (layer4_outputs(298)) or (layer4_outputs(971));
    layer5_outputs(654) <= not((layer4_outputs(2544)) and (layer4_outputs(960)));
    layer5_outputs(655) <= not((layer4_outputs(194)) or (layer4_outputs(426)));
    layer5_outputs(656) <= not((layer4_outputs(2379)) or (layer4_outputs(472)));
    layer5_outputs(657) <= layer4_outputs(486);
    layer5_outputs(658) <= not(layer4_outputs(1360)) or (layer4_outputs(1372));
    layer5_outputs(659) <= layer4_outputs(99);
    layer5_outputs(660) <= layer4_outputs(1977);
    layer5_outputs(661) <= not((layer4_outputs(735)) or (layer4_outputs(1696)));
    layer5_outputs(662) <= not(layer4_outputs(1060));
    layer5_outputs(663) <= not(layer4_outputs(1760));
    layer5_outputs(664) <= not(layer4_outputs(313));
    layer5_outputs(665) <= not(layer4_outputs(2441));
    layer5_outputs(666) <= (layer4_outputs(2067)) and not (layer4_outputs(1511));
    layer5_outputs(667) <= layer4_outputs(1525);
    layer5_outputs(668) <= not(layer4_outputs(907));
    layer5_outputs(669) <= not((layer4_outputs(392)) or (layer4_outputs(2559)));
    layer5_outputs(670) <= not(layer4_outputs(984));
    layer5_outputs(671) <= not((layer4_outputs(862)) xor (layer4_outputs(14)));
    layer5_outputs(672) <= '1';
    layer5_outputs(673) <= not(layer4_outputs(2327));
    layer5_outputs(674) <= not(layer4_outputs(1196)) or (layer4_outputs(1010));
    layer5_outputs(675) <= not(layer4_outputs(2006));
    layer5_outputs(676) <= (layer4_outputs(838)) or (layer4_outputs(840));
    layer5_outputs(677) <= (layer4_outputs(2137)) and not (layer4_outputs(2135));
    layer5_outputs(678) <= (layer4_outputs(2362)) or (layer4_outputs(708));
    layer5_outputs(679) <= (layer4_outputs(1156)) and not (layer4_outputs(924));
    layer5_outputs(680) <= (layer4_outputs(976)) and not (layer4_outputs(2215));
    layer5_outputs(681) <= layer4_outputs(2114);
    layer5_outputs(682) <= (layer4_outputs(598)) xor (layer4_outputs(1883));
    layer5_outputs(683) <= not(layer4_outputs(1595)) or (layer4_outputs(1754));
    layer5_outputs(684) <= not(layer4_outputs(780));
    layer5_outputs(685) <= not((layer4_outputs(728)) or (layer4_outputs(1443)));
    layer5_outputs(686) <= not(layer4_outputs(2333)) or (layer4_outputs(1161));
    layer5_outputs(687) <= not((layer4_outputs(1660)) xor (layer4_outputs(244)));
    layer5_outputs(688) <= not(layer4_outputs(940)) or (layer4_outputs(859));
    layer5_outputs(689) <= layer4_outputs(2235);
    layer5_outputs(690) <= (layer4_outputs(18)) or (layer4_outputs(1922));
    layer5_outputs(691) <= not(layer4_outputs(2244));
    layer5_outputs(692) <= not(layer4_outputs(946));
    layer5_outputs(693) <= not((layer4_outputs(2224)) xor (layer4_outputs(719)));
    layer5_outputs(694) <= not(layer4_outputs(2422));
    layer5_outputs(695) <= layer4_outputs(2269);
    layer5_outputs(696) <= layer4_outputs(2172);
    layer5_outputs(697) <= '1';
    layer5_outputs(698) <= layer4_outputs(52);
    layer5_outputs(699) <= not(layer4_outputs(1998)) or (layer4_outputs(1858));
    layer5_outputs(700) <= (layer4_outputs(2047)) xor (layer4_outputs(2459));
    layer5_outputs(701) <= not(layer4_outputs(335));
    layer5_outputs(702) <= layer4_outputs(1176);
    layer5_outputs(703) <= not(layer4_outputs(1645));
    layer5_outputs(704) <= (layer4_outputs(1849)) or (layer4_outputs(836));
    layer5_outputs(705) <= (layer4_outputs(1441)) and not (layer4_outputs(503));
    layer5_outputs(706) <= layer4_outputs(776);
    layer5_outputs(707) <= layer4_outputs(1150);
    layer5_outputs(708) <= '0';
    layer5_outputs(709) <= (layer4_outputs(1065)) and not (layer4_outputs(2178));
    layer5_outputs(710) <= (layer4_outputs(1159)) and (layer4_outputs(264));
    layer5_outputs(711) <= not(layer4_outputs(941)) or (layer4_outputs(2209));
    layer5_outputs(712) <= layer4_outputs(168);
    layer5_outputs(713) <= layer4_outputs(1721);
    layer5_outputs(714) <= (layer4_outputs(2032)) and not (layer4_outputs(2256));
    layer5_outputs(715) <= not(layer4_outputs(634));
    layer5_outputs(716) <= layer4_outputs(1062);
    layer5_outputs(717) <= not((layer4_outputs(830)) or (layer4_outputs(2336)));
    layer5_outputs(718) <= layer4_outputs(1438);
    layer5_outputs(719) <= (layer4_outputs(2367)) and (layer4_outputs(1464));
    layer5_outputs(720) <= not(layer4_outputs(384));
    layer5_outputs(721) <= layer4_outputs(1457);
    layer5_outputs(722) <= (layer4_outputs(1194)) and not (layer4_outputs(2040));
    layer5_outputs(723) <= not((layer4_outputs(171)) xor (layer4_outputs(2080)));
    layer5_outputs(724) <= (layer4_outputs(2443)) and not (layer4_outputs(177));
    layer5_outputs(725) <= (layer4_outputs(400)) and (layer4_outputs(862));
    layer5_outputs(726) <= not(layer4_outputs(1210));
    layer5_outputs(727) <= not(layer4_outputs(1225)) or (layer4_outputs(1761));
    layer5_outputs(728) <= layer4_outputs(2487);
    layer5_outputs(729) <= layer4_outputs(501);
    layer5_outputs(730) <= (layer4_outputs(1904)) and not (layer4_outputs(245));
    layer5_outputs(731) <= not(layer4_outputs(1806));
    layer5_outputs(732) <= '1';
    layer5_outputs(733) <= layer4_outputs(2535);
    layer5_outputs(734) <= not((layer4_outputs(535)) and (layer4_outputs(1788)));
    layer5_outputs(735) <= (layer4_outputs(2464)) xor (layer4_outputs(565));
    layer5_outputs(736) <= (layer4_outputs(1987)) xor (layer4_outputs(1772));
    layer5_outputs(737) <= not(layer4_outputs(164)) or (layer4_outputs(122));
    layer5_outputs(738) <= (layer4_outputs(2040)) and not (layer4_outputs(438));
    layer5_outputs(739) <= (layer4_outputs(276)) and not (layer4_outputs(1275));
    layer5_outputs(740) <= not(layer4_outputs(1539)) or (layer4_outputs(2543));
    layer5_outputs(741) <= (layer4_outputs(694)) and not (layer4_outputs(218));
    layer5_outputs(742) <= (layer4_outputs(2509)) or (layer4_outputs(423));
    layer5_outputs(743) <= not(layer4_outputs(437));
    layer5_outputs(744) <= layer4_outputs(2010);
    layer5_outputs(745) <= not(layer4_outputs(710));
    layer5_outputs(746) <= not((layer4_outputs(2338)) or (layer4_outputs(1096)));
    layer5_outputs(747) <= layer4_outputs(1752);
    layer5_outputs(748) <= not(layer4_outputs(1885));
    layer5_outputs(749) <= not(layer4_outputs(2479)) or (layer4_outputs(1987));
    layer5_outputs(750) <= (layer4_outputs(165)) or (layer4_outputs(881));
    layer5_outputs(751) <= not((layer4_outputs(2085)) xor (layer4_outputs(212)));
    layer5_outputs(752) <= not(layer4_outputs(455));
    layer5_outputs(753) <= not(layer4_outputs(1656)) or (layer4_outputs(464));
    layer5_outputs(754) <= not(layer4_outputs(1654));
    layer5_outputs(755) <= not(layer4_outputs(2248));
    layer5_outputs(756) <= (layer4_outputs(1854)) or (layer4_outputs(465));
    layer5_outputs(757) <= layer4_outputs(1596);
    layer5_outputs(758) <= not(layer4_outputs(2290));
    layer5_outputs(759) <= not(layer4_outputs(1056));
    layer5_outputs(760) <= layer4_outputs(1278);
    layer5_outputs(761) <= layer4_outputs(1891);
    layer5_outputs(762) <= layer4_outputs(2152);
    layer5_outputs(763) <= layer4_outputs(65);
    layer5_outputs(764) <= not((layer4_outputs(2222)) xor (layer4_outputs(2525)));
    layer5_outputs(765) <= (layer4_outputs(902)) and not (layer4_outputs(551));
    layer5_outputs(766) <= (layer4_outputs(1337)) and (layer4_outputs(1042));
    layer5_outputs(767) <= layer4_outputs(2544);
    layer5_outputs(768) <= (layer4_outputs(1342)) or (layer4_outputs(1848));
    layer5_outputs(769) <= not(layer4_outputs(1657));
    layer5_outputs(770) <= not(layer4_outputs(1396));
    layer5_outputs(771) <= layer4_outputs(144);
    layer5_outputs(772) <= layer4_outputs(2309);
    layer5_outputs(773) <= not((layer4_outputs(884)) or (layer4_outputs(554)));
    layer5_outputs(774) <= layer4_outputs(2310);
    layer5_outputs(775) <= not(layer4_outputs(2256)) or (layer4_outputs(260));
    layer5_outputs(776) <= not(layer4_outputs(1429));
    layer5_outputs(777) <= not(layer4_outputs(1103));
    layer5_outputs(778) <= layer4_outputs(73);
    layer5_outputs(779) <= layer4_outputs(381);
    layer5_outputs(780) <= layer4_outputs(2262);
    layer5_outputs(781) <= (layer4_outputs(1660)) and not (layer4_outputs(1789));
    layer5_outputs(782) <= (layer4_outputs(2525)) and not (layer4_outputs(2119));
    layer5_outputs(783) <= not((layer4_outputs(2293)) xor (layer4_outputs(1607)));
    layer5_outputs(784) <= not(layer4_outputs(31));
    layer5_outputs(785) <= not((layer4_outputs(1029)) and (layer4_outputs(2071)));
    layer5_outputs(786) <= (layer4_outputs(1998)) and not (layer4_outputs(1878));
    layer5_outputs(787) <= '0';
    layer5_outputs(788) <= not(layer4_outputs(1469));
    layer5_outputs(789) <= layer4_outputs(551);
    layer5_outputs(790) <= layer4_outputs(2445);
    layer5_outputs(791) <= not(layer4_outputs(1263));
    layer5_outputs(792) <= layer4_outputs(1997);
    layer5_outputs(793) <= not(layer4_outputs(1180));
    layer5_outputs(794) <= not((layer4_outputs(870)) or (layer4_outputs(1352)));
    layer5_outputs(795) <= (layer4_outputs(1553)) xor (layer4_outputs(1132));
    layer5_outputs(796) <= not(layer4_outputs(765));
    layer5_outputs(797) <= layer4_outputs(933);
    layer5_outputs(798) <= (layer4_outputs(900)) and not (layer4_outputs(1124));
    layer5_outputs(799) <= (layer4_outputs(811)) and (layer4_outputs(1569));
    layer5_outputs(800) <= '1';
    layer5_outputs(801) <= not(layer4_outputs(2127));
    layer5_outputs(802) <= not(layer4_outputs(1319));
    layer5_outputs(803) <= not(layer4_outputs(1917));
    layer5_outputs(804) <= not(layer4_outputs(278)) or (layer4_outputs(1532));
    layer5_outputs(805) <= layer4_outputs(637);
    layer5_outputs(806) <= not(layer4_outputs(886));
    layer5_outputs(807) <= not(layer4_outputs(468));
    layer5_outputs(808) <= (layer4_outputs(25)) and not (layer4_outputs(1378));
    layer5_outputs(809) <= not(layer4_outputs(90)) or (layer4_outputs(2252));
    layer5_outputs(810) <= not(layer4_outputs(134)) or (layer4_outputs(340));
    layer5_outputs(811) <= layer4_outputs(2058);
    layer5_outputs(812) <= not(layer4_outputs(131));
    layer5_outputs(813) <= (layer4_outputs(78)) or (layer4_outputs(1449));
    layer5_outputs(814) <= not(layer4_outputs(502)) or (layer4_outputs(2083));
    layer5_outputs(815) <= layer4_outputs(2384);
    layer5_outputs(816) <= (layer4_outputs(654)) and (layer4_outputs(1765));
    layer5_outputs(817) <= (layer4_outputs(223)) and not (layer4_outputs(2376));
    layer5_outputs(818) <= (layer4_outputs(2261)) and (layer4_outputs(128));
    layer5_outputs(819) <= (layer4_outputs(1964)) and not (layer4_outputs(403));
    layer5_outputs(820) <= layer4_outputs(2550);
    layer5_outputs(821) <= (layer4_outputs(556)) and (layer4_outputs(724));
    layer5_outputs(822) <= layer4_outputs(964);
    layer5_outputs(823) <= layer4_outputs(304);
    layer5_outputs(824) <= (layer4_outputs(204)) and not (layer4_outputs(1588));
    layer5_outputs(825) <= not((layer4_outputs(754)) or (layer4_outputs(930)));
    layer5_outputs(826) <= not((layer4_outputs(28)) xor (layer4_outputs(1591)));
    layer5_outputs(827) <= not(layer4_outputs(373));
    layer5_outputs(828) <= not((layer4_outputs(1130)) xor (layer4_outputs(1716)));
    layer5_outputs(829) <= not((layer4_outputs(487)) and (layer4_outputs(522)));
    layer5_outputs(830) <= not((layer4_outputs(2348)) xor (layer4_outputs(1771)));
    layer5_outputs(831) <= not(layer4_outputs(1256));
    layer5_outputs(832) <= (layer4_outputs(878)) and (layer4_outputs(1370));
    layer5_outputs(833) <= not((layer4_outputs(2530)) and (layer4_outputs(979)));
    layer5_outputs(834) <= layer4_outputs(1716);
    layer5_outputs(835) <= (layer4_outputs(556)) and not (layer4_outputs(2380));
    layer5_outputs(836) <= layer4_outputs(2036);
    layer5_outputs(837) <= not(layer4_outputs(1234));
    layer5_outputs(838) <= layer4_outputs(786);
    layer5_outputs(839) <= (layer4_outputs(1603)) and not (layer4_outputs(532));
    layer5_outputs(840) <= (layer4_outputs(596)) and (layer4_outputs(1337));
    layer5_outputs(841) <= (layer4_outputs(24)) xor (layer4_outputs(2076));
    layer5_outputs(842) <= not(layer4_outputs(1281)) or (layer4_outputs(2558));
    layer5_outputs(843) <= (layer4_outputs(329)) and not (layer4_outputs(1852));
    layer5_outputs(844) <= layer4_outputs(2046);
    layer5_outputs(845) <= (layer4_outputs(1078)) and (layer4_outputs(1347));
    layer5_outputs(846) <= not(layer4_outputs(1727));
    layer5_outputs(847) <= '1';
    layer5_outputs(848) <= layer4_outputs(636);
    layer5_outputs(849) <= not(layer4_outputs(1953)) or (layer4_outputs(2340));
    layer5_outputs(850) <= (layer4_outputs(716)) and not (layer4_outputs(812));
    layer5_outputs(851) <= not(layer4_outputs(1836)) or (layer4_outputs(904));
    layer5_outputs(852) <= layer4_outputs(2145);
    layer5_outputs(853) <= (layer4_outputs(1908)) or (layer4_outputs(1021));
    layer5_outputs(854) <= not((layer4_outputs(1397)) or (layer4_outputs(2434)));
    layer5_outputs(855) <= layer4_outputs(1185);
    layer5_outputs(856) <= layer4_outputs(1694);
    layer5_outputs(857) <= (layer4_outputs(361)) and not (layer4_outputs(1587));
    layer5_outputs(858) <= (layer4_outputs(1791)) or (layer4_outputs(635));
    layer5_outputs(859) <= not(layer4_outputs(742));
    layer5_outputs(860) <= not(layer4_outputs(1299));
    layer5_outputs(861) <= not((layer4_outputs(2230)) xor (layer4_outputs(608)));
    layer5_outputs(862) <= layer4_outputs(1220);
    layer5_outputs(863) <= layer4_outputs(449);
    layer5_outputs(864) <= layer4_outputs(1076);
    layer5_outputs(865) <= '0';
    layer5_outputs(866) <= not((layer4_outputs(1115)) and (layer4_outputs(893)));
    layer5_outputs(867) <= not(layer4_outputs(1375));
    layer5_outputs(868) <= (layer4_outputs(1633)) xor (layer4_outputs(732));
    layer5_outputs(869) <= (layer4_outputs(992)) and not (layer4_outputs(847));
    layer5_outputs(870) <= (layer4_outputs(1691)) and (layer4_outputs(247));
    layer5_outputs(871) <= not((layer4_outputs(533)) xor (layer4_outputs(2011)));
    layer5_outputs(872) <= layer4_outputs(393);
    layer5_outputs(873) <= layer4_outputs(831);
    layer5_outputs(874) <= layer4_outputs(2314);
    layer5_outputs(875) <= not((layer4_outputs(2476)) xor (layer4_outputs(1579)));
    layer5_outputs(876) <= not(layer4_outputs(964));
    layer5_outputs(877) <= (layer4_outputs(2306)) and not (layer4_outputs(1186));
    layer5_outputs(878) <= (layer4_outputs(1110)) and not (layer4_outputs(145));
    layer5_outputs(879) <= not(layer4_outputs(242));
    layer5_outputs(880) <= not((layer4_outputs(575)) and (layer4_outputs(46)));
    layer5_outputs(881) <= not(layer4_outputs(1564));
    layer5_outputs(882) <= not(layer4_outputs(2354)) or (layer4_outputs(1637));
    layer5_outputs(883) <= not((layer4_outputs(2056)) and (layer4_outputs(1560)));
    layer5_outputs(884) <= layer4_outputs(1311);
    layer5_outputs(885) <= not((layer4_outputs(2380)) and (layer4_outputs(230)));
    layer5_outputs(886) <= not(layer4_outputs(2005)) or (layer4_outputs(108));
    layer5_outputs(887) <= layer4_outputs(323);
    layer5_outputs(888) <= layer4_outputs(860);
    layer5_outputs(889) <= (layer4_outputs(584)) and not (layer4_outputs(2147));
    layer5_outputs(890) <= not(layer4_outputs(1678));
    layer5_outputs(891) <= not(layer4_outputs(232));
    layer5_outputs(892) <= layer4_outputs(2454);
    layer5_outputs(893) <= not(layer4_outputs(1573));
    layer5_outputs(894) <= not(layer4_outputs(649));
    layer5_outputs(895) <= not((layer4_outputs(322)) or (layer4_outputs(53)));
    layer5_outputs(896) <= not(layer4_outputs(186)) or (layer4_outputs(1594));
    layer5_outputs(897) <= not((layer4_outputs(560)) and (layer4_outputs(1005)));
    layer5_outputs(898) <= not(layer4_outputs(2264));
    layer5_outputs(899) <= not(layer4_outputs(2366));
    layer5_outputs(900) <= (layer4_outputs(128)) or (layer4_outputs(2328));
    layer5_outputs(901) <= layer4_outputs(721);
    layer5_outputs(902) <= layer4_outputs(1344);
    layer5_outputs(903) <= layer4_outputs(508);
    layer5_outputs(904) <= (layer4_outputs(103)) and (layer4_outputs(1147));
    layer5_outputs(905) <= not(layer4_outputs(2134)) or (layer4_outputs(1518));
    layer5_outputs(906) <= layer4_outputs(1365);
    layer5_outputs(907) <= (layer4_outputs(126)) and (layer4_outputs(574));
    layer5_outputs(908) <= (layer4_outputs(1402)) and not (layer4_outputs(318));
    layer5_outputs(909) <= (layer4_outputs(491)) and (layer4_outputs(2493));
    layer5_outputs(910) <= (layer4_outputs(1166)) or (layer4_outputs(262));
    layer5_outputs(911) <= (layer4_outputs(1636)) and not (layer4_outputs(1310));
    layer5_outputs(912) <= layer4_outputs(22);
    layer5_outputs(913) <= (layer4_outputs(2180)) and not (layer4_outputs(758));
    layer5_outputs(914) <= not(layer4_outputs(225));
    layer5_outputs(915) <= not(layer4_outputs(549)) or (layer4_outputs(1894));
    layer5_outputs(916) <= not(layer4_outputs(833));
    layer5_outputs(917) <= layer4_outputs(2205);
    layer5_outputs(918) <= not(layer4_outputs(1608)) or (layer4_outputs(1570));
    layer5_outputs(919) <= (layer4_outputs(331)) xor (layer4_outputs(1748));
    layer5_outputs(920) <= not(layer4_outputs(1618)) or (layer4_outputs(243));
    layer5_outputs(921) <= layer4_outputs(1505);
    layer5_outputs(922) <= layer4_outputs(903);
    layer5_outputs(923) <= (layer4_outputs(1025)) xor (layer4_outputs(1845));
    layer5_outputs(924) <= (layer4_outputs(1907)) and not (layer4_outputs(1412));
    layer5_outputs(925) <= not((layer4_outputs(28)) xor (layer4_outputs(1974)));
    layer5_outputs(926) <= (layer4_outputs(407)) and not (layer4_outputs(103));
    layer5_outputs(927) <= not((layer4_outputs(1725)) xor (layer4_outputs(648)));
    layer5_outputs(928) <= not(layer4_outputs(1083));
    layer5_outputs(929) <= not((layer4_outputs(1243)) or (layer4_outputs(2346)));
    layer5_outputs(930) <= (layer4_outputs(1803)) and not (layer4_outputs(1661));
    layer5_outputs(931) <= not(layer4_outputs(88)) or (layer4_outputs(309));
    layer5_outputs(932) <= (layer4_outputs(970)) and (layer4_outputs(839));
    layer5_outputs(933) <= not(layer4_outputs(297)) or (layer4_outputs(1069));
    layer5_outputs(934) <= not(layer4_outputs(279));
    layer5_outputs(935) <= layer4_outputs(898);
    layer5_outputs(936) <= not(layer4_outputs(169));
    layer5_outputs(937) <= layer4_outputs(1484);
    layer5_outputs(938) <= not(layer4_outputs(442));
    layer5_outputs(939) <= (layer4_outputs(1428)) and not (layer4_outputs(1533));
    layer5_outputs(940) <= (layer4_outputs(539)) xor (layer4_outputs(1233));
    layer5_outputs(941) <= layer4_outputs(1033);
    layer5_outputs(942) <= layer4_outputs(15);
    layer5_outputs(943) <= layer4_outputs(1855);
    layer5_outputs(944) <= not(layer4_outputs(1373)) or (layer4_outputs(2306));
    layer5_outputs(945) <= not(layer4_outputs(1956));
    layer5_outputs(946) <= layer4_outputs(93);
    layer5_outputs(947) <= layer4_outputs(2092);
    layer5_outputs(948) <= layer4_outputs(2328);
    layer5_outputs(949) <= layer4_outputs(1632);
    layer5_outputs(950) <= (layer4_outputs(910)) or (layer4_outputs(2124));
    layer5_outputs(951) <= not((layer4_outputs(1963)) and (layer4_outputs(1562)));
    layer5_outputs(952) <= not(layer4_outputs(2083));
    layer5_outputs(953) <= not(layer4_outputs(2263));
    layer5_outputs(954) <= (layer4_outputs(2139)) xor (layer4_outputs(2523));
    layer5_outputs(955) <= (layer4_outputs(224)) and not (layer4_outputs(571));
    layer5_outputs(956) <= (layer4_outputs(2121)) and (layer4_outputs(2397));
    layer5_outputs(957) <= not(layer4_outputs(867));
    layer5_outputs(958) <= not((layer4_outputs(2002)) and (layer4_outputs(2095)));
    layer5_outputs(959) <= not((layer4_outputs(2251)) and (layer4_outputs(1140)));
    layer5_outputs(960) <= not(layer4_outputs(858));
    layer5_outputs(961) <= layer4_outputs(641);
    layer5_outputs(962) <= not(layer4_outputs(334));
    layer5_outputs(963) <= layer4_outputs(639);
    layer5_outputs(964) <= layer4_outputs(996);
    layer5_outputs(965) <= not(layer4_outputs(1189));
    layer5_outputs(966) <= layer4_outputs(876);
    layer5_outputs(967) <= layer4_outputs(2437);
    layer5_outputs(968) <= not(layer4_outputs(207));
    layer5_outputs(969) <= (layer4_outputs(174)) and (layer4_outputs(2325));
    layer5_outputs(970) <= layer4_outputs(2341);
    layer5_outputs(971) <= not((layer4_outputs(1957)) and (layer4_outputs(1624)));
    layer5_outputs(972) <= not(layer4_outputs(2424));
    layer5_outputs(973) <= layer4_outputs(2318);
    layer5_outputs(974) <= not(layer4_outputs(1738)) or (layer4_outputs(1299));
    layer5_outputs(975) <= not(layer4_outputs(153));
    layer5_outputs(976) <= not(layer4_outputs(676));
    layer5_outputs(977) <= '0';
    layer5_outputs(978) <= (layer4_outputs(2065)) and not (layer4_outputs(1830));
    layer5_outputs(979) <= not((layer4_outputs(832)) and (layer4_outputs(1654)));
    layer5_outputs(980) <= not(layer4_outputs(1093));
    layer5_outputs(981) <= (layer4_outputs(2455)) and (layer4_outputs(2390));
    layer5_outputs(982) <= not(layer4_outputs(577)) or (layer4_outputs(1831));
    layer5_outputs(983) <= not(layer4_outputs(2128));
    layer5_outputs(984) <= (layer4_outputs(630)) and not (layer4_outputs(139));
    layer5_outputs(985) <= (layer4_outputs(2298)) and not (layer4_outputs(1952));
    layer5_outputs(986) <= not(layer4_outputs(1795));
    layer5_outputs(987) <= (layer4_outputs(665)) or (layer4_outputs(830));
    layer5_outputs(988) <= not(layer4_outputs(1451));
    layer5_outputs(989) <= not(layer4_outputs(1316)) or (layer4_outputs(166));
    layer5_outputs(990) <= not(layer4_outputs(2494));
    layer5_outputs(991) <= not(layer4_outputs(1598)) or (layer4_outputs(1087));
    layer5_outputs(992) <= not(layer4_outputs(2200)) or (layer4_outputs(454));
    layer5_outputs(993) <= not((layer4_outputs(375)) xor (layer4_outputs(2236)));
    layer5_outputs(994) <= '1';
    layer5_outputs(995) <= not(layer4_outputs(1391));
    layer5_outputs(996) <= not((layer4_outputs(1546)) and (layer4_outputs(2365)));
    layer5_outputs(997) <= not(layer4_outputs(765));
    layer5_outputs(998) <= not((layer4_outputs(1139)) xor (layer4_outputs(1821)));
    layer5_outputs(999) <= not(layer4_outputs(1196));
    layer5_outputs(1000) <= not(layer4_outputs(1788));
    layer5_outputs(1001) <= (layer4_outputs(932)) or (layer4_outputs(1322));
    layer5_outputs(1002) <= not((layer4_outputs(1373)) xor (layer4_outputs(559)));
    layer5_outputs(1003) <= not(layer4_outputs(2293));
    layer5_outputs(1004) <= not(layer4_outputs(346));
    layer5_outputs(1005) <= not((layer4_outputs(1447)) and (layer4_outputs(179)));
    layer5_outputs(1006) <= not((layer4_outputs(957)) or (layer4_outputs(499)));
    layer5_outputs(1007) <= not(layer4_outputs(674));
    layer5_outputs(1008) <= not(layer4_outputs(433));
    layer5_outputs(1009) <= not((layer4_outputs(441)) and (layer4_outputs(1659)));
    layer5_outputs(1010) <= not(layer4_outputs(960));
    layer5_outputs(1011) <= layer4_outputs(824);
    layer5_outputs(1012) <= not(layer4_outputs(371));
    layer5_outputs(1013) <= not(layer4_outputs(1347));
    layer5_outputs(1014) <= layer4_outputs(362);
    layer5_outputs(1015) <= not((layer4_outputs(700)) xor (layer4_outputs(2278)));
    layer5_outputs(1016) <= not((layer4_outputs(2471)) xor (layer4_outputs(1976)));
    layer5_outputs(1017) <= not((layer4_outputs(2116)) or (layer4_outputs(2542)));
    layer5_outputs(1018) <= not((layer4_outputs(2312)) and (layer4_outputs(365)));
    layer5_outputs(1019) <= not((layer4_outputs(267)) xor (layer4_outputs(1249)));
    layer5_outputs(1020) <= (layer4_outputs(1711)) and not (layer4_outputs(1131));
    layer5_outputs(1021) <= not(layer4_outputs(1296)) or (layer4_outputs(2396));
    layer5_outputs(1022) <= not((layer4_outputs(1877)) xor (layer4_outputs(591)));
    layer5_outputs(1023) <= not(layer4_outputs(2376));
    layer5_outputs(1024) <= not(layer4_outputs(1335));
    layer5_outputs(1025) <= not(layer4_outputs(380)) or (layer4_outputs(890));
    layer5_outputs(1026) <= layer4_outputs(2126);
    layer5_outputs(1027) <= not((layer4_outputs(1099)) or (layer4_outputs(1767)));
    layer5_outputs(1028) <= not((layer4_outputs(544)) or (layer4_outputs(1869)));
    layer5_outputs(1029) <= not(layer4_outputs(500));
    layer5_outputs(1030) <= not((layer4_outputs(2475)) or (layer4_outputs(1300)));
    layer5_outputs(1031) <= (layer4_outputs(2510)) or (layer4_outputs(843));
    layer5_outputs(1032) <= not(layer4_outputs(1583));
    layer5_outputs(1033) <= not((layer4_outputs(2407)) xor (layer4_outputs(1943)));
    layer5_outputs(1034) <= layer4_outputs(636);
    layer5_outputs(1035) <= not(layer4_outputs(1617));
    layer5_outputs(1036) <= not(layer4_outputs(1916)) or (layer4_outputs(82));
    layer5_outputs(1037) <= (layer4_outputs(53)) and (layer4_outputs(2009));
    layer5_outputs(1038) <= (layer4_outputs(819)) xor (layer4_outputs(1817));
    layer5_outputs(1039) <= not((layer4_outputs(1292)) or (layer4_outputs(1784)));
    layer5_outputs(1040) <= not(layer4_outputs(1575));
    layer5_outputs(1041) <= layer4_outputs(1108);
    layer5_outputs(1042) <= not((layer4_outputs(710)) or (layer4_outputs(496)));
    layer5_outputs(1043) <= (layer4_outputs(1502)) and not (layer4_outputs(2184));
    layer5_outputs(1044) <= not(layer4_outputs(1121)) or (layer4_outputs(1577));
    layer5_outputs(1045) <= not(layer4_outputs(1317));
    layer5_outputs(1046) <= (layer4_outputs(1058)) and not (layer4_outputs(1842));
    layer5_outputs(1047) <= (layer4_outputs(2404)) and not (layer4_outputs(2513));
    layer5_outputs(1048) <= not(layer4_outputs(101)) or (layer4_outputs(147));
    layer5_outputs(1049) <= not(layer4_outputs(647));
    layer5_outputs(1050) <= not(layer4_outputs(2369));
    layer5_outputs(1051) <= not(layer4_outputs(1880));
    layer5_outputs(1052) <= not((layer4_outputs(425)) and (layer4_outputs(1147)));
    layer5_outputs(1053) <= layer4_outputs(867);
    layer5_outputs(1054) <= layer4_outputs(354);
    layer5_outputs(1055) <= (layer4_outputs(1007)) and not (layer4_outputs(422));
    layer5_outputs(1056) <= not((layer4_outputs(1506)) or (layer4_outputs(498)));
    layer5_outputs(1057) <= layer4_outputs(819);
    layer5_outputs(1058) <= not(layer4_outputs(1057));
    layer5_outputs(1059) <= (layer4_outputs(2387)) and not (layer4_outputs(1950));
    layer5_outputs(1060) <= layer4_outputs(984);
    layer5_outputs(1061) <= (layer4_outputs(1341)) and not (layer4_outputs(325));
    layer5_outputs(1062) <= not(layer4_outputs(2508)) or (layer4_outputs(2088));
    layer5_outputs(1063) <= layer4_outputs(2454);
    layer5_outputs(1064) <= (layer4_outputs(1089)) and not (layer4_outputs(645));
    layer5_outputs(1065) <= (layer4_outputs(877)) xor (layer4_outputs(1453));
    layer5_outputs(1066) <= not((layer4_outputs(196)) or (layer4_outputs(572)));
    layer5_outputs(1067) <= '1';
    layer5_outputs(1068) <= (layer4_outputs(180)) and (layer4_outputs(1134));
    layer5_outputs(1069) <= (layer4_outputs(2315)) and (layer4_outputs(161));
    layer5_outputs(1070) <= (layer4_outputs(1349)) and not (layer4_outputs(955));
    layer5_outputs(1071) <= not(layer4_outputs(2313));
    layer5_outputs(1072) <= (layer4_outputs(905)) or (layer4_outputs(2436));
    layer5_outputs(1073) <= layer4_outputs(2458);
    layer5_outputs(1074) <= (layer4_outputs(949)) and (layer4_outputs(970));
    layer5_outputs(1075) <= not(layer4_outputs(1420));
    layer5_outputs(1076) <= '1';
    layer5_outputs(1077) <= not(layer4_outputs(2159)) or (layer4_outputs(136));
    layer5_outputs(1078) <= not(layer4_outputs(598));
    layer5_outputs(1079) <= not((layer4_outputs(1356)) or (layer4_outputs(2541)));
    layer5_outputs(1080) <= (layer4_outputs(711)) or (layer4_outputs(1067));
    layer5_outputs(1081) <= (layer4_outputs(666)) and not (layer4_outputs(2498));
    layer5_outputs(1082) <= layer4_outputs(620);
    layer5_outputs(1083) <= not(layer4_outputs(86));
    layer5_outputs(1084) <= not(layer4_outputs(1909)) or (layer4_outputs(2106));
    layer5_outputs(1085) <= '0';
    layer5_outputs(1086) <= not((layer4_outputs(483)) xor (layer4_outputs(1368)));
    layer5_outputs(1087) <= (layer4_outputs(445)) and not (layer4_outputs(2072));
    layer5_outputs(1088) <= layer4_outputs(1766);
    layer5_outputs(1089) <= layer4_outputs(1930);
    layer5_outputs(1090) <= '0';
    layer5_outputs(1091) <= '1';
    layer5_outputs(1092) <= not((layer4_outputs(1385)) or (layer4_outputs(1265)));
    layer5_outputs(1093) <= not((layer4_outputs(1554)) or (layer4_outputs(2435)));
    layer5_outputs(1094) <= (layer4_outputs(1580)) and not (layer4_outputs(1167));
    layer5_outputs(1095) <= layer4_outputs(294);
    layer5_outputs(1096) <= not(layer4_outputs(255));
    layer5_outputs(1097) <= not(layer4_outputs(155)) or (layer4_outputs(1989));
    layer5_outputs(1098) <= not(layer4_outputs(1972));
    layer5_outputs(1099) <= not(layer4_outputs(1486));
    layer5_outputs(1100) <= (layer4_outputs(1032)) or (layer4_outputs(2141));
    layer5_outputs(1101) <= (layer4_outputs(195)) and not (layer4_outputs(530));
    layer5_outputs(1102) <= layer4_outputs(1503);
    layer5_outputs(1103) <= not((layer4_outputs(1336)) xor (layer4_outputs(248)));
    layer5_outputs(1104) <= (layer4_outputs(769)) or (layer4_outputs(1777));
    layer5_outputs(1105) <= not(layer4_outputs(1534));
    layer5_outputs(1106) <= (layer4_outputs(201)) and not (layer4_outputs(2006));
    layer5_outputs(1107) <= (layer4_outputs(2063)) and not (layer4_outputs(331));
    layer5_outputs(1108) <= not(layer4_outputs(2455));
    layer5_outputs(1109) <= not(layer4_outputs(1679));
    layer5_outputs(1110) <= (layer4_outputs(2462)) and not (layer4_outputs(2521));
    layer5_outputs(1111) <= not((layer4_outputs(2286)) and (layer4_outputs(2514)));
    layer5_outputs(1112) <= not(layer4_outputs(731)) or (layer4_outputs(1155));
    layer5_outputs(1113) <= not(layer4_outputs(181));
    layer5_outputs(1114) <= not(layer4_outputs(985)) or (layer4_outputs(1180));
    layer5_outputs(1115) <= not(layer4_outputs(1701));
    layer5_outputs(1116) <= not(layer4_outputs(2255)) or (layer4_outputs(2547));
    layer5_outputs(1117) <= not(layer4_outputs(738)) or (layer4_outputs(1070));
    layer5_outputs(1118) <= layer4_outputs(2172);
    layer5_outputs(1119) <= layer4_outputs(2322);
    layer5_outputs(1120) <= layer4_outputs(144);
    layer5_outputs(1121) <= not(layer4_outputs(2037));
    layer5_outputs(1122) <= layer4_outputs(1295);
    layer5_outputs(1123) <= (layer4_outputs(2059)) and not (layer4_outputs(2168));
    layer5_outputs(1124) <= layer4_outputs(1470);
    layer5_outputs(1125) <= not(layer4_outputs(2023));
    layer5_outputs(1126) <= not(layer4_outputs(79));
    layer5_outputs(1127) <= (layer4_outputs(264)) and not (layer4_outputs(471));
    layer5_outputs(1128) <= '0';
    layer5_outputs(1129) <= not((layer4_outputs(1958)) or (layer4_outputs(1605)));
    layer5_outputs(1130) <= layer4_outputs(2178);
    layer5_outputs(1131) <= '1';
    layer5_outputs(1132) <= not(layer4_outputs(238));
    layer5_outputs(1133) <= (layer4_outputs(672)) and not (layer4_outputs(2202));
    layer5_outputs(1134) <= layer4_outputs(341);
    layer5_outputs(1135) <= not(layer4_outputs(2457)) or (layer4_outputs(1071));
    layer5_outputs(1136) <= not((layer4_outputs(2277)) and (layer4_outputs(1190)));
    layer5_outputs(1137) <= (layer4_outputs(1874)) or (layer4_outputs(1485));
    layer5_outputs(1138) <= not((layer4_outputs(1304)) or (layer4_outputs(923)));
    layer5_outputs(1139) <= layer4_outputs(726);
    layer5_outputs(1140) <= (layer4_outputs(2163)) and not (layer4_outputs(324));
    layer5_outputs(1141) <= (layer4_outputs(985)) and (layer4_outputs(707));
    layer5_outputs(1142) <= layer4_outputs(700);
    layer5_outputs(1143) <= not(layer4_outputs(456));
    layer5_outputs(1144) <= (layer4_outputs(2038)) or (layer4_outputs(1712));
    layer5_outputs(1145) <= not(layer4_outputs(1313));
    layer5_outputs(1146) <= not(layer4_outputs(731)) or (layer4_outputs(593));
    layer5_outputs(1147) <= not(layer4_outputs(2208));
    layer5_outputs(1148) <= not(layer4_outputs(2333));
    layer5_outputs(1149) <= not((layer4_outputs(1732)) xor (layer4_outputs(730)));
    layer5_outputs(1150) <= layer4_outputs(139);
    layer5_outputs(1151) <= '0';
    layer5_outputs(1152) <= (layer4_outputs(1425)) and not (layer4_outputs(1269));
    layer5_outputs(1153) <= '0';
    layer5_outputs(1154) <= (layer4_outputs(163)) or (layer4_outputs(1145));
    layer5_outputs(1155) <= (layer4_outputs(1808)) or (layer4_outputs(238));
    layer5_outputs(1156) <= (layer4_outputs(2270)) and not (layer4_outputs(2519));
    layer5_outputs(1157) <= not(layer4_outputs(1475));
    layer5_outputs(1158) <= not(layer4_outputs(1673));
    layer5_outputs(1159) <= layer4_outputs(56);
    layer5_outputs(1160) <= not(layer4_outputs(190));
    layer5_outputs(1161) <= '0';
    layer5_outputs(1162) <= not((layer4_outputs(288)) xor (layer4_outputs(917)));
    layer5_outputs(1163) <= (layer4_outputs(1320)) xor (layer4_outputs(1355));
    layer5_outputs(1164) <= (layer4_outputs(266)) xor (layer4_outputs(7));
    layer5_outputs(1165) <= not(layer4_outputs(2482));
    layer5_outputs(1166) <= '1';
    layer5_outputs(1167) <= layer4_outputs(826);
    layer5_outputs(1168) <= (layer4_outputs(116)) xor (layer4_outputs(761));
    layer5_outputs(1169) <= not(layer4_outputs(1307)) or (layer4_outputs(2084));
    layer5_outputs(1170) <= layer4_outputs(229);
    layer5_outputs(1171) <= not((layer4_outputs(2323)) and (layer4_outputs(816)));
    layer5_outputs(1172) <= not((layer4_outputs(1287)) xor (layer4_outputs(896)));
    layer5_outputs(1173) <= layer4_outputs(851);
    layer5_outputs(1174) <= layer4_outputs(777);
    layer5_outputs(1175) <= layer4_outputs(218);
    layer5_outputs(1176) <= (layer4_outputs(469)) and not (layer4_outputs(580));
    layer5_outputs(1177) <= (layer4_outputs(2489)) xor (layer4_outputs(367));
    layer5_outputs(1178) <= layer4_outputs(806);
    layer5_outputs(1179) <= (layer4_outputs(803)) and (layer4_outputs(755));
    layer5_outputs(1180) <= not((layer4_outputs(1479)) and (layer4_outputs(730)));
    layer5_outputs(1181) <= layer4_outputs(2230);
    layer5_outputs(1182) <= (layer4_outputs(1529)) and not (layer4_outputs(1114));
    layer5_outputs(1183) <= not((layer4_outputs(1398)) and (layer4_outputs(1138)));
    layer5_outputs(1184) <= not(layer4_outputs(2347));
    layer5_outputs(1185) <= not(layer4_outputs(721));
    layer5_outputs(1186) <= '0';
    layer5_outputs(1187) <= (layer4_outputs(1687)) and not (layer4_outputs(783));
    layer5_outputs(1188) <= layer4_outputs(1190);
    layer5_outputs(1189) <= (layer4_outputs(610)) and (layer4_outputs(2291));
    layer5_outputs(1190) <= not(layer4_outputs(1284));
    layer5_outputs(1191) <= not(layer4_outputs(2251));
    layer5_outputs(1192) <= (layer4_outputs(129)) and (layer4_outputs(834));
    layer5_outputs(1193) <= layer4_outputs(2528);
    layer5_outputs(1194) <= layer4_outputs(1566);
    layer5_outputs(1195) <= layer4_outputs(1876);
    layer5_outputs(1196) <= not(layer4_outputs(271));
    layer5_outputs(1197) <= not(layer4_outputs(1379));
    layer5_outputs(1198) <= layer4_outputs(2385);
    layer5_outputs(1199) <= not((layer4_outputs(1383)) xor (layer4_outputs(2546)));
    layer5_outputs(1200) <= (layer4_outputs(2426)) xor (layer4_outputs(1740));
    layer5_outputs(1201) <= layer4_outputs(1807);
    layer5_outputs(1202) <= layer4_outputs(395);
    layer5_outputs(1203) <= (layer4_outputs(851)) or (layer4_outputs(485));
    layer5_outputs(1204) <= not(layer4_outputs(117));
    layer5_outputs(1205) <= not((layer4_outputs(37)) xor (layer4_outputs(2532)));
    layer5_outputs(1206) <= (layer4_outputs(1432)) and not (layer4_outputs(1074));
    layer5_outputs(1207) <= (layer4_outputs(608)) and not (layer4_outputs(1846));
    layer5_outputs(1208) <= (layer4_outputs(1259)) and (layer4_outputs(661));
    layer5_outputs(1209) <= not(layer4_outputs(1584));
    layer5_outputs(1210) <= layer4_outputs(204);
    layer5_outputs(1211) <= (layer4_outputs(555)) xor (layer4_outputs(673));
    layer5_outputs(1212) <= '1';
    layer5_outputs(1213) <= not((layer4_outputs(774)) or (layer4_outputs(982)));
    layer5_outputs(1214) <= layer4_outputs(1422);
    layer5_outputs(1215) <= not(layer4_outputs(2176)) or (layer4_outputs(2472));
    layer5_outputs(1216) <= not(layer4_outputs(1313)) or (layer4_outputs(809));
    layer5_outputs(1217) <= (layer4_outputs(1827)) and not (layer4_outputs(590));
    layer5_outputs(1218) <= not(layer4_outputs(157));
    layer5_outputs(1219) <= not(layer4_outputs(11));
    layer5_outputs(1220) <= (layer4_outputs(1077)) xor (layer4_outputs(170));
    layer5_outputs(1221) <= layer4_outputs(249);
    layer5_outputs(1222) <= not((layer4_outputs(614)) xor (layer4_outputs(1900)));
    layer5_outputs(1223) <= (layer4_outputs(2277)) and not (layer4_outputs(2530));
    layer5_outputs(1224) <= not(layer4_outputs(2204));
    layer5_outputs(1225) <= layer4_outputs(2418);
    layer5_outputs(1226) <= (layer4_outputs(480)) and not (layer4_outputs(814));
    layer5_outputs(1227) <= not((layer4_outputs(1861)) xor (layer4_outputs(352)));
    layer5_outputs(1228) <= layer4_outputs(2481);
    layer5_outputs(1229) <= layer4_outputs(2393);
    layer5_outputs(1230) <= not((layer4_outputs(1240)) or (layer4_outputs(801)));
    layer5_outputs(1231) <= not(layer4_outputs(195));
    layer5_outputs(1232) <= not(layer4_outputs(2359)) or (layer4_outputs(1932));
    layer5_outputs(1233) <= not((layer4_outputs(2502)) xor (layer4_outputs(859)));
    layer5_outputs(1234) <= not((layer4_outputs(863)) or (layer4_outputs(714)));
    layer5_outputs(1235) <= layer4_outputs(2448);
    layer5_outputs(1236) <= layer4_outputs(687);
    layer5_outputs(1237) <= not(layer4_outputs(1527));
    layer5_outputs(1238) <= not(layer4_outputs(279)) or (layer4_outputs(475));
    layer5_outputs(1239) <= not((layer4_outputs(2049)) or (layer4_outputs(633)));
    layer5_outputs(1240) <= not(layer4_outputs(1641)) or (layer4_outputs(1332));
    layer5_outputs(1241) <= (layer4_outputs(1888)) and (layer4_outputs(2179));
    layer5_outputs(1242) <= (layer4_outputs(1751)) and not (layer4_outputs(1175));
    layer5_outputs(1243) <= not(layer4_outputs(2175));
    layer5_outputs(1244) <= layer4_outputs(1684);
    layer5_outputs(1245) <= not(layer4_outputs(1415)) or (layer4_outputs(94));
    layer5_outputs(1246) <= not(layer4_outputs(497));
    layer5_outputs(1247) <= layer4_outputs(432);
    layer5_outputs(1248) <= layer4_outputs(2260);
    layer5_outputs(1249) <= not(layer4_outputs(990)) or (layer4_outputs(800));
    layer5_outputs(1250) <= (layer4_outputs(2136)) or (layer4_outputs(764));
    layer5_outputs(1251) <= '1';
    layer5_outputs(1252) <= not(layer4_outputs(1792));
    layer5_outputs(1253) <= not(layer4_outputs(2557)) or (layer4_outputs(1572));
    layer5_outputs(1254) <= '0';
    layer5_outputs(1255) <= not(layer4_outputs(2266));
    layer5_outputs(1256) <= (layer4_outputs(1571)) and not (layer4_outputs(632));
    layer5_outputs(1257) <= not(layer4_outputs(1867)) or (layer4_outputs(2002));
    layer5_outputs(1258) <= not(layer4_outputs(2233));
    layer5_outputs(1259) <= layer4_outputs(2082);
    layer5_outputs(1260) <= (layer4_outputs(1208)) or (layer4_outputs(1304));
    layer5_outputs(1261) <= not((layer4_outputs(448)) and (layer4_outputs(272)));
    layer5_outputs(1262) <= not(layer4_outputs(2430));
    layer5_outputs(1263) <= not(layer4_outputs(1022));
    layer5_outputs(1264) <= layer4_outputs(2350);
    layer5_outputs(1265) <= '1';
    layer5_outputs(1266) <= not(layer4_outputs(79));
    layer5_outputs(1267) <= not(layer4_outputs(2112));
    layer5_outputs(1268) <= (layer4_outputs(332)) and not (layer4_outputs(1742));
    layer5_outputs(1269) <= (layer4_outputs(60)) and not (layer4_outputs(1522));
    layer5_outputs(1270) <= (layer4_outputs(734)) and not (layer4_outputs(343));
    layer5_outputs(1271) <= layer4_outputs(2213);
    layer5_outputs(1272) <= layer4_outputs(2499);
    layer5_outputs(1273) <= (layer4_outputs(891)) and (layer4_outputs(1327));
    layer5_outputs(1274) <= (layer4_outputs(1682)) and not (layer4_outputs(2283));
    layer5_outputs(1275) <= (layer4_outputs(1019)) and not (layer4_outputs(1548));
    layer5_outputs(1276) <= layer4_outputs(1901);
    layer5_outputs(1277) <= not(layer4_outputs(1736));
    layer5_outputs(1278) <= not(layer4_outputs(20));
    layer5_outputs(1279) <= (layer4_outputs(1969)) xor (layer4_outputs(1984));
    layer5_outputs(1280) <= '1';
    layer5_outputs(1281) <= (layer4_outputs(54)) xor (layer4_outputs(698));
    layer5_outputs(1282) <= not((layer4_outputs(1746)) or (layer4_outputs(1364)));
    layer5_outputs(1283) <= not(layer4_outputs(102)) or (layer4_outputs(1923));
    layer5_outputs(1284) <= (layer4_outputs(2480)) or (layer4_outputs(2477));
    layer5_outputs(1285) <= not(layer4_outputs(1747));
    layer5_outputs(1286) <= not(layer4_outputs(0));
    layer5_outputs(1287) <= not(layer4_outputs(355));
    layer5_outputs(1288) <= not(layer4_outputs(2437));
    layer5_outputs(1289) <= layer4_outputs(951);
    layer5_outputs(1290) <= (layer4_outputs(290)) xor (layer4_outputs(2406));
    layer5_outputs(1291) <= (layer4_outputs(1361)) and (layer4_outputs(376));
    layer5_outputs(1292) <= not(layer4_outputs(652)) or (layer4_outputs(74));
    layer5_outputs(1293) <= layer4_outputs(130);
    layer5_outputs(1294) <= not(layer4_outputs(2194));
    layer5_outputs(1295) <= layer4_outputs(1126);
    layer5_outputs(1296) <= layer4_outputs(1143);
    layer5_outputs(1297) <= layer4_outputs(1252);
    layer5_outputs(1298) <= not(layer4_outputs(1414)) or (layer4_outputs(148));
    layer5_outputs(1299) <= not(layer4_outputs(1470)) or (layer4_outputs(2442));
    layer5_outputs(1300) <= not(layer4_outputs(1794));
    layer5_outputs(1301) <= (layer4_outputs(2259)) xor (layer4_outputs(1498));
    layer5_outputs(1302) <= (layer4_outputs(922)) and not (layer4_outputs(390));
    layer5_outputs(1303) <= layer4_outputs(1393);
    layer5_outputs(1304) <= layer4_outputs(2512);
    layer5_outputs(1305) <= (layer4_outputs(1881)) and (layer4_outputs(240));
    layer5_outputs(1306) <= layer4_outputs(1416);
    layer5_outputs(1307) <= not((layer4_outputs(2548)) xor (layer4_outputs(2415)));
    layer5_outputs(1308) <= not(layer4_outputs(1538));
    layer5_outputs(1309) <= not(layer4_outputs(2196));
    layer5_outputs(1310) <= not(layer4_outputs(772));
    layer5_outputs(1311) <= layer4_outputs(209);
    layer5_outputs(1312) <= not(layer4_outputs(1210));
    layer5_outputs(1313) <= not(layer4_outputs(311));
    layer5_outputs(1314) <= not(layer4_outputs(109)) or (layer4_outputs(1288));
    layer5_outputs(1315) <= not((layer4_outputs(874)) xor (layer4_outputs(1633)));
    layer5_outputs(1316) <= not(layer4_outputs(1764)) or (layer4_outputs(2171));
    layer5_outputs(1317) <= not(layer4_outputs(1863)) or (layer4_outputs(1300));
    layer5_outputs(1318) <= layer4_outputs(2465);
    layer5_outputs(1319) <= (layer4_outputs(2167)) or (layer4_outputs(678));
    layer5_outputs(1320) <= (layer4_outputs(1879)) and (layer4_outputs(291));
    layer5_outputs(1321) <= '0';
    layer5_outputs(1322) <= layer4_outputs(1956);
    layer5_outputs(1323) <= not(layer4_outputs(1400)) or (layer4_outputs(709));
    layer5_outputs(1324) <= not((layer4_outputs(341)) xor (layer4_outputs(1847)));
    layer5_outputs(1325) <= not(layer4_outputs(225));
    layer5_outputs(1326) <= not(layer4_outputs(1220)) or (layer4_outputs(1169));
    layer5_outputs(1327) <= not(layer4_outputs(2399)) or (layer4_outputs(2521));
    layer5_outputs(1328) <= (layer4_outputs(1456)) and not (layer4_outputs(405));
    layer5_outputs(1329) <= not(layer4_outputs(1349)) or (layer4_outputs(1850));
    layer5_outputs(1330) <= not(layer4_outputs(461));
    layer5_outputs(1331) <= layer4_outputs(1826);
    layer5_outputs(1332) <= not((layer4_outputs(770)) and (layer4_outputs(205)));
    layer5_outputs(1333) <= (layer4_outputs(1766)) and not (layer4_outputs(2233));
    layer5_outputs(1334) <= not((layer4_outputs(217)) xor (layer4_outputs(1815)));
    layer5_outputs(1335) <= not(layer4_outputs(977));
    layer5_outputs(1336) <= (layer4_outputs(665)) and (layer4_outputs(981));
    layer5_outputs(1337) <= (layer4_outputs(1733)) and not (layer4_outputs(762));
    layer5_outputs(1338) <= layer4_outputs(440);
    layer5_outputs(1339) <= layer4_outputs(1886);
    layer5_outputs(1340) <= not(layer4_outputs(928));
    layer5_outputs(1341) <= not(layer4_outputs(466));
    layer5_outputs(1342) <= layer4_outputs(2484);
    layer5_outputs(1343) <= not(layer4_outputs(1779));
    layer5_outputs(1344) <= (layer4_outputs(1648)) and not (layer4_outputs(1563));
    layer5_outputs(1345) <= layer4_outputs(2084);
    layer5_outputs(1346) <= (layer4_outputs(1729)) and (layer4_outputs(2266));
    layer5_outputs(1347) <= not(layer4_outputs(506));
    layer5_outputs(1348) <= not(layer4_outputs(2307));
    layer5_outputs(1349) <= layer4_outputs(1199);
    layer5_outputs(1350) <= layer4_outputs(510);
    layer5_outputs(1351) <= not(layer4_outputs(1254));
    layer5_outputs(1352) <= not((layer4_outputs(2351)) and (layer4_outputs(2499)));
    layer5_outputs(1353) <= (layer4_outputs(1521)) and (layer4_outputs(1515));
    layer5_outputs(1354) <= not((layer4_outputs(659)) and (layer4_outputs(1772)));
    layer5_outputs(1355) <= not(layer4_outputs(2104)) or (layer4_outputs(2361));
    layer5_outputs(1356) <= (layer4_outputs(1013)) or (layer4_outputs(1329));
    layer5_outputs(1357) <= layer4_outputs(2036);
    layer5_outputs(1358) <= not(layer4_outputs(382)) or (layer4_outputs(550));
    layer5_outputs(1359) <= (layer4_outputs(846)) or (layer4_outputs(1955));
    layer5_outputs(1360) <= layer4_outputs(470);
    layer5_outputs(1361) <= not(layer4_outputs(335));
    layer5_outputs(1362) <= not(layer4_outputs(1755));
    layer5_outputs(1363) <= not(layer4_outputs(1392)) or (layer4_outputs(1895));
    layer5_outputs(1364) <= layer4_outputs(1524);
    layer5_outputs(1365) <= layer4_outputs(1435);
    layer5_outputs(1366) <= not(layer4_outputs(2303));
    layer5_outputs(1367) <= layer4_outputs(370);
    layer5_outputs(1368) <= (layer4_outputs(742)) xor (layer4_outputs(589));
    layer5_outputs(1369) <= layer4_outputs(586);
    layer5_outputs(1370) <= (layer4_outputs(528)) and not (layer4_outputs(2411));
    layer5_outputs(1371) <= not((layer4_outputs(2515)) or (layer4_outputs(1638)));
    layer5_outputs(1372) <= layer4_outputs(2275);
    layer5_outputs(1373) <= not(layer4_outputs(959));
    layer5_outputs(1374) <= not(layer4_outputs(1063));
    layer5_outputs(1375) <= not(layer4_outputs(868)) or (layer4_outputs(2035));
    layer5_outputs(1376) <= layer4_outputs(845);
    layer5_outputs(1377) <= layer4_outputs(1468);
    layer5_outputs(1378) <= (layer4_outputs(981)) and not (layer4_outputs(2389));
    layer5_outputs(1379) <= layer4_outputs(1790);
    layer5_outputs(1380) <= layer4_outputs(821);
    layer5_outputs(1381) <= not(layer4_outputs(200));
    layer5_outputs(1382) <= (layer4_outputs(963)) and (layer4_outputs(2285));
    layer5_outputs(1383) <= not((layer4_outputs(1182)) xor (layer4_outputs(557)));
    layer5_outputs(1384) <= not(layer4_outputs(2405));
    layer5_outputs(1385) <= not(layer4_outputs(146)) or (layer4_outputs(942));
    layer5_outputs(1386) <= not((layer4_outputs(2364)) and (layer4_outputs(501)));
    layer5_outputs(1387) <= (layer4_outputs(1244)) and not (layer4_outputs(2484));
    layer5_outputs(1388) <= layer4_outputs(416);
    layer5_outputs(1389) <= not(layer4_outputs(2275)) or (layer4_outputs(1801));
    layer5_outputs(1390) <= not(layer4_outputs(394));
    layer5_outputs(1391) <= (layer4_outputs(1554)) and not (layer4_outputs(317));
    layer5_outputs(1392) <= not(layer4_outputs(921));
    layer5_outputs(1393) <= not((layer4_outputs(2341)) xor (layer4_outputs(462)));
    layer5_outputs(1394) <= (layer4_outputs(63)) and not (layer4_outputs(1030));
    layer5_outputs(1395) <= (layer4_outputs(829)) and not (layer4_outputs(486));
    layer5_outputs(1396) <= (layer4_outputs(404)) xor (layer4_outputs(982));
    layer5_outputs(1397) <= layer4_outputs(861);
    layer5_outputs(1398) <= (layer4_outputs(397)) and not (layer4_outputs(236));
    layer5_outputs(1399) <= layer4_outputs(1250);
    layer5_outputs(1400) <= not(layer4_outputs(618));
    layer5_outputs(1401) <= layer4_outputs(1162);
    layer5_outputs(1402) <= not(layer4_outputs(250));
    layer5_outputs(1403) <= layer4_outputs(1064);
    layer5_outputs(1404) <= (layer4_outputs(724)) xor (layer4_outputs(606));
    layer5_outputs(1405) <= (layer4_outputs(2490)) and (layer4_outputs(2156));
    layer5_outputs(1406) <= layer4_outputs(2120);
    layer5_outputs(1407) <= (layer4_outputs(883)) and not (layer4_outputs(512));
    layer5_outputs(1408) <= not((layer4_outputs(1084)) xor (layer4_outputs(747)));
    layer5_outputs(1409) <= not((layer4_outputs(1444)) xor (layer4_outputs(1088)));
    layer5_outputs(1410) <= '1';
    layer5_outputs(1411) <= not(layer4_outputs(1565));
    layer5_outputs(1412) <= not((layer4_outputs(576)) xor (layer4_outputs(1782)));
    layer5_outputs(1413) <= not((layer4_outputs(1201)) xor (layer4_outputs(516)));
    layer5_outputs(1414) <= not(layer4_outputs(47));
    layer5_outputs(1415) <= (layer4_outputs(399)) and (layer4_outputs(792));
    layer5_outputs(1416) <= layer4_outputs(1619);
    layer5_outputs(1417) <= not(layer4_outputs(1427));
    layer5_outputs(1418) <= not((layer4_outputs(2066)) or (layer4_outputs(2214)));
    layer5_outputs(1419) <= layer4_outputs(2203);
    layer5_outputs(1420) <= (layer4_outputs(1463)) and (layer4_outputs(2145));
    layer5_outputs(1421) <= layer4_outputs(2265);
    layer5_outputs(1422) <= not(layer4_outputs(1188)) or (layer4_outputs(457));
    layer5_outputs(1423) <= not((layer4_outputs(558)) and (layer4_outputs(85)));
    layer5_outputs(1424) <= layer4_outputs(113);
    layer5_outputs(1425) <= not(layer4_outputs(453));
    layer5_outputs(1426) <= (layer4_outputs(1513)) and not (layer4_outputs(1493));
    layer5_outputs(1427) <= layer4_outputs(358);
    layer5_outputs(1428) <= not(layer4_outputs(282)) or (layer4_outputs(978));
    layer5_outputs(1429) <= layer4_outputs(2382);
    layer5_outputs(1430) <= not(layer4_outputs(1798)) or (layer4_outputs(1090));
    layer5_outputs(1431) <= not((layer4_outputs(16)) or (layer4_outputs(1640)));
    layer5_outputs(1432) <= layer4_outputs(348);
    layer5_outputs(1433) <= layer4_outputs(25);
    layer5_outputs(1434) <= '0';
    layer5_outputs(1435) <= not(layer4_outputs(308)) or (layer4_outputs(1593));
    layer5_outputs(1436) <= layer4_outputs(1117);
    layer5_outputs(1437) <= (layer4_outputs(1122)) and not (layer4_outputs(1152));
    layer5_outputs(1438) <= not(layer4_outputs(1516));
    layer5_outputs(1439) <= (layer4_outputs(1583)) and (layer4_outputs(160));
    layer5_outputs(1440) <= not(layer4_outputs(1362));
    layer5_outputs(1441) <= (layer4_outputs(1673)) or (layer4_outputs(2089));
    layer5_outputs(1442) <= not(layer4_outputs(2427)) or (layer4_outputs(708));
    layer5_outputs(1443) <= not((layer4_outputs(1044)) or (layer4_outputs(1868)));
    layer5_outputs(1444) <= not((layer4_outputs(263)) and (layer4_outputs(582)));
    layer5_outputs(1445) <= layer4_outputs(946);
    layer5_outputs(1446) <= layer4_outputs(1862);
    layer5_outputs(1447) <= layer4_outputs(948);
    layer5_outputs(1448) <= not((layer4_outputs(1879)) xor (layer4_outputs(1867)));
    layer5_outputs(1449) <= not(layer4_outputs(38));
    layer5_outputs(1450) <= layer4_outputs(747);
    layer5_outputs(1451) <= '1';
    layer5_outputs(1452) <= (layer4_outputs(44)) and (layer4_outputs(886));
    layer5_outputs(1453) <= not(layer4_outputs(2272)) or (layer4_outputs(1011));
    layer5_outputs(1454) <= layer4_outputs(1278);
    layer5_outputs(1455) <= layer4_outputs(935);
    layer5_outputs(1456) <= (layer4_outputs(723)) and not (layer4_outputs(2400));
    layer5_outputs(1457) <= layer4_outputs(60);
    layer5_outputs(1458) <= not(layer4_outputs(1709)) or (layer4_outputs(2168));
    layer5_outputs(1459) <= '1';
    layer5_outputs(1460) <= (layer4_outputs(51)) xor (layer4_outputs(1737));
    layer5_outputs(1461) <= '0';
    layer5_outputs(1462) <= layer4_outputs(2467);
    layer5_outputs(1463) <= '1';
    layer5_outputs(1464) <= not(layer4_outputs(1582)) or (layer4_outputs(226));
    layer5_outputs(1465) <= not(layer4_outputs(2424)) or (layer4_outputs(2057));
    layer5_outputs(1466) <= not(layer4_outputs(1091));
    layer5_outputs(1467) <= layer4_outputs(568);
    layer5_outputs(1468) <= (layer4_outputs(0)) and (layer4_outputs(2201));
    layer5_outputs(1469) <= (layer4_outputs(1303)) and (layer4_outputs(529));
    layer5_outputs(1470) <= not((layer4_outputs(935)) and (layer4_outputs(987)));
    layer5_outputs(1471) <= not((layer4_outputs(977)) or (layer4_outputs(2554)));
    layer5_outputs(1472) <= not(layer4_outputs(1734));
    layer5_outputs(1473) <= not(layer4_outputs(372));
    layer5_outputs(1474) <= not(layer4_outputs(292));
    layer5_outputs(1475) <= '1';
    layer5_outputs(1476) <= not(layer4_outputs(1463)) or (layer4_outputs(2034));
    layer5_outputs(1477) <= layer4_outputs(538);
    layer5_outputs(1478) <= not((layer4_outputs(1723)) xor (layer4_outputs(2226)));
    layer5_outputs(1479) <= '1';
    layer5_outputs(1480) <= layer4_outputs(1496);
    layer5_outputs(1481) <= layer4_outputs(2217);
    layer5_outputs(1482) <= not((layer4_outputs(239)) xor (layer4_outputs(1207)));
    layer5_outputs(1483) <= not((layer4_outputs(1318)) and (layer4_outputs(439)));
    layer5_outputs(1484) <= (layer4_outputs(1238)) or (layer4_outputs(921));
    layer5_outputs(1485) <= not((layer4_outputs(2358)) and (layer4_outputs(1283)));
    layer5_outputs(1486) <= not(layer4_outputs(197)) or (layer4_outputs(223));
    layer5_outputs(1487) <= (layer4_outputs(1466)) and (layer4_outputs(2319));
    layer5_outputs(1488) <= not(layer4_outputs(2261));
    layer5_outputs(1489) <= (layer4_outputs(2469)) or (layer4_outputs(1179));
    layer5_outputs(1490) <= not(layer4_outputs(2110)) or (layer4_outputs(470));
    layer5_outputs(1491) <= layer4_outputs(1379);
    layer5_outputs(1492) <= (layer4_outputs(55)) and (layer4_outputs(706));
    layer5_outputs(1493) <= (layer4_outputs(2391)) and not (layer4_outputs(2440));
    layer5_outputs(1494) <= not(layer4_outputs(1119)) or (layer4_outputs(2374));
    layer5_outputs(1495) <= not(layer4_outputs(1364));
    layer5_outputs(1496) <= (layer4_outputs(286)) and (layer4_outputs(563));
    layer5_outputs(1497) <= (layer4_outputs(359)) xor (layer4_outputs(124));
    layer5_outputs(1498) <= not((layer4_outputs(1309)) or (layer4_outputs(1489)));
    layer5_outputs(1499) <= (layer4_outputs(1542)) and (layer4_outputs(760));
    layer5_outputs(1500) <= not(layer4_outputs(2453));
    layer5_outputs(1501) <= (layer4_outputs(1433)) and not (layer4_outputs(1852));
    layer5_outputs(1502) <= layer4_outputs(2150);
    layer5_outputs(1503) <= layer4_outputs(2466);
    layer5_outputs(1504) <= (layer4_outputs(1149)) or (layer4_outputs(140));
    layer5_outputs(1505) <= (layer4_outputs(241)) and (layer4_outputs(926));
    layer5_outputs(1506) <= not(layer4_outputs(1753));
    layer5_outputs(1507) <= layer4_outputs(478);
    layer5_outputs(1508) <= layer4_outputs(1782);
    layer5_outputs(1509) <= not(layer4_outputs(1992)) or (layer4_outputs(1251));
    layer5_outputs(1510) <= not((layer4_outputs(1944)) or (layer4_outputs(818)));
    layer5_outputs(1511) <= (layer4_outputs(546)) or (layer4_outputs(187));
    layer5_outputs(1512) <= not((layer4_outputs(1635)) xor (layer4_outputs(926)));
    layer5_outputs(1513) <= layer4_outputs(677);
    layer5_outputs(1514) <= layer4_outputs(2075);
    layer5_outputs(1515) <= layer4_outputs(895);
    layer5_outputs(1516) <= not(layer4_outputs(2399));
    layer5_outputs(1517) <= (layer4_outputs(1367)) and (layer4_outputs(2193));
    layer5_outputs(1518) <= layer4_outputs(953);
    layer5_outputs(1519) <= (layer4_outputs(1628)) xor (layer4_outputs(1015));
    layer5_outputs(1520) <= (layer4_outputs(702)) xor (layer4_outputs(1999));
    layer5_outputs(1521) <= layer4_outputs(2003);
    layer5_outputs(1522) <= not((layer4_outputs(1822)) xor (layer4_outputs(2421)));
    layer5_outputs(1523) <= (layer4_outputs(1938)) xor (layer4_outputs(1450));
    layer5_outputs(1524) <= (layer4_outputs(1261)) or (layer4_outputs(2200));
    layer5_outputs(1525) <= layer4_outputs(391);
    layer5_outputs(1526) <= not((layer4_outputs(65)) or (layer4_outputs(2536)));
    layer5_outputs(1527) <= (layer4_outputs(1498)) or (layer4_outputs(2407));
    layer5_outputs(1528) <= not(layer4_outputs(2052)) or (layer4_outputs(1949));
    layer5_outputs(1529) <= not(layer4_outputs(1011));
    layer5_outputs(1530) <= '1';
    layer5_outputs(1531) <= (layer4_outputs(2260)) and not (layer4_outputs(725));
    layer5_outputs(1532) <= layer4_outputs(2016);
    layer5_outputs(1533) <= not(layer4_outputs(659));
    layer5_outputs(1534) <= not(layer4_outputs(1468)) or (layer4_outputs(2496));
    layer5_outputs(1535) <= not((layer4_outputs(15)) or (layer4_outputs(1530)));
    layer5_outputs(1536) <= not(layer4_outputs(2144));
    layer5_outputs(1537) <= (layer4_outputs(301)) and not (layer4_outputs(1006));
    layer5_outputs(1538) <= not((layer4_outputs(1556)) and (layer4_outputs(1399)));
    layer5_outputs(1539) <= layer4_outputs(1248);
    layer5_outputs(1540) <= not(layer4_outputs(1802));
    layer5_outputs(1541) <= layer4_outputs(130);
    layer5_outputs(1542) <= '1';
    layer5_outputs(1543) <= (layer4_outputs(1756)) or (layer4_outputs(1982));
    layer5_outputs(1544) <= not(layer4_outputs(1164)) or (layer4_outputs(1754));
    layer5_outputs(1545) <= layer4_outputs(798);
    layer5_outputs(1546) <= '1';
    layer5_outputs(1547) <= not(layer4_outputs(1818)) or (layer4_outputs(602));
    layer5_outputs(1548) <= not(layer4_outputs(1991));
    layer5_outputs(1549) <= layer4_outputs(231);
    layer5_outputs(1550) <= (layer4_outputs(1722)) xor (layer4_outputs(1204));
    layer5_outputs(1551) <= not(layer4_outputs(614)) or (layer4_outputs(1966));
    layer5_outputs(1552) <= (layer4_outputs(775)) and not (layer4_outputs(2073));
    layer5_outputs(1553) <= not(layer4_outputs(326));
    layer5_outputs(1554) <= not(layer4_outputs(174));
    layer5_outputs(1555) <= (layer4_outputs(836)) and not (layer4_outputs(1902));
    layer5_outputs(1556) <= not(layer4_outputs(693));
    layer5_outputs(1557) <= not(layer4_outputs(1137));
    layer5_outputs(1558) <= not(layer4_outputs(45));
    layer5_outputs(1559) <= not((layer4_outputs(1476)) or (layer4_outputs(515)));
    layer5_outputs(1560) <= '1';
    layer5_outputs(1561) <= not(layer4_outputs(2551)) or (layer4_outputs(404));
    layer5_outputs(1562) <= layer4_outputs(1510);
    layer5_outputs(1563) <= (layer4_outputs(952)) and not (layer4_outputs(1388));
    layer5_outputs(1564) <= layer4_outputs(2216);
    layer5_outputs(1565) <= '0';
    layer5_outputs(1566) <= (layer4_outputs(1507)) and (layer4_outputs(469));
    layer5_outputs(1567) <= layer4_outputs(927);
    layer5_outputs(1568) <= (layer4_outputs(803)) and (layer4_outputs(684));
    layer5_outputs(1569) <= not(layer4_outputs(2410));
    layer5_outputs(1570) <= not(layer4_outputs(666));
    layer5_outputs(1571) <= not(layer4_outputs(293));
    layer5_outputs(1572) <= '0';
    layer5_outputs(1573) <= not(layer4_outputs(151));
    layer5_outputs(1574) <= (layer4_outputs(369)) xor (layer4_outputs(1323));
    layer5_outputs(1575) <= layer4_outputs(699);
    layer5_outputs(1576) <= (layer4_outputs(1722)) and not (layer4_outputs(1829));
    layer5_outputs(1577) <= layer4_outputs(2504);
    layer5_outputs(1578) <= not(layer4_outputs(21)) or (layer4_outputs(311));
    layer5_outputs(1579) <= not(layer4_outputs(1940));
    layer5_outputs(1580) <= (layer4_outputs(34)) and not (layer4_outputs(1384));
    layer5_outputs(1581) <= layer4_outputs(2128);
    layer5_outputs(1582) <= not(layer4_outputs(1535));
    layer5_outputs(1583) <= (layer4_outputs(254)) and not (layer4_outputs(1615));
    layer5_outputs(1584) <= (layer4_outputs(2532)) and not (layer4_outputs(988));
    layer5_outputs(1585) <= layer4_outputs(1475);
    layer5_outputs(1586) <= layer4_outputs(1135);
    layer5_outputs(1587) <= (layer4_outputs(2395)) and not (layer4_outputs(780));
    layer5_outputs(1588) <= '1';
    layer5_outputs(1589) <= not(layer4_outputs(1621));
    layer5_outputs(1590) <= layer4_outputs(252);
    layer5_outputs(1591) <= layer4_outputs(1541);
    layer5_outputs(1592) <= not((layer4_outputs(1314)) or (layer4_outputs(692)));
    layer5_outputs(1593) <= not(layer4_outputs(1119));
    layer5_outputs(1594) <= not((layer4_outputs(962)) and (layer4_outputs(555)));
    layer5_outputs(1595) <= not(layer4_outputs(1178));
    layer5_outputs(1596) <= not(layer4_outputs(2189));
    layer5_outputs(1597) <= (layer4_outputs(2044)) and (layer4_outputs(2234));
    layer5_outputs(1598) <= not(layer4_outputs(1741));
    layer5_outputs(1599) <= (layer4_outputs(1334)) xor (layer4_outputs(1257));
    layer5_outputs(1600) <= not(layer4_outputs(513)) or (layer4_outputs(696));
    layer5_outputs(1601) <= (layer4_outputs(2281)) and not (layer4_outputs(518));
    layer5_outputs(1602) <= not(layer4_outputs(1704)) or (layer4_outputs(1864));
    layer5_outputs(1603) <= not(layer4_outputs(740));
    layer5_outputs(1604) <= not((layer4_outputs(999)) xor (layer4_outputs(1773)));
    layer5_outputs(1605) <= (layer4_outputs(1483)) and not (layer4_outputs(605));
    layer5_outputs(1606) <= not(layer4_outputs(430));
    layer5_outputs(1607) <= layer4_outputs(662);
    layer5_outputs(1608) <= not(layer4_outputs(1446)) or (layer4_outputs(183));
    layer5_outputs(1609) <= not(layer4_outputs(402));
    layer5_outputs(1610) <= (layer4_outputs(330)) and not (layer4_outputs(825));
    layer5_outputs(1611) <= not((layer4_outputs(1667)) xor (layer4_outputs(137)));
    layer5_outputs(1612) <= (layer4_outputs(1643)) or (layer4_outputs(1101));
    layer5_outputs(1613) <= not(layer4_outputs(392)) or (layer4_outputs(1765));
    layer5_outputs(1614) <= (layer4_outputs(736)) and not (layer4_outputs(1503));
    layer5_outputs(1615) <= '0';
    layer5_outputs(1616) <= not(layer4_outputs(519));
    layer5_outputs(1617) <= not(layer4_outputs(2355));
    layer5_outputs(1618) <= (layer4_outputs(2024)) xor (layer4_outputs(944));
    layer5_outputs(1619) <= layer4_outputs(127);
    layer5_outputs(1620) <= not(layer4_outputs(570));
    layer5_outputs(1621) <= not((layer4_outputs(337)) xor (layer4_outputs(1170)));
    layer5_outputs(1622) <= (layer4_outputs(2173)) and not (layer4_outputs(1620));
    layer5_outputs(1623) <= (layer4_outputs(1436)) and (layer4_outputs(613));
    layer5_outputs(1624) <= (layer4_outputs(107)) and not (layer4_outputs(284));
    layer5_outputs(1625) <= layer4_outputs(1133);
    layer5_outputs(1626) <= layer4_outputs(1824);
    layer5_outputs(1627) <= layer4_outputs(2027);
    layer5_outputs(1628) <= '1';
    layer5_outputs(1629) <= not((layer4_outputs(688)) and (layer4_outputs(41)));
    layer5_outputs(1630) <= not(layer4_outputs(1001)) or (layer4_outputs(398));
    layer5_outputs(1631) <= (layer4_outputs(1454)) and not (layer4_outputs(980));
    layer5_outputs(1632) <= layer4_outputs(1729);
    layer5_outputs(1633) <= (layer4_outputs(689)) and not (layer4_outputs(568));
    layer5_outputs(1634) <= (layer4_outputs(2077)) xor (layer4_outputs(1290));
    layer5_outputs(1635) <= (layer4_outputs(1342)) or (layer4_outputs(1358));
    layer5_outputs(1636) <= layer4_outputs(1255);
    layer5_outputs(1637) <= (layer4_outputs(1243)) and (layer4_outputs(2393));
    layer5_outputs(1638) <= not((layer4_outputs(1871)) or (layer4_outputs(1868)));
    layer5_outputs(1639) <= not(layer4_outputs(1735));
    layer5_outputs(1640) <= not(layer4_outputs(2236));
    layer5_outputs(1641) <= '1';
    layer5_outputs(1642) <= not(layer4_outputs(932)) or (layer4_outputs(569));
    layer5_outputs(1643) <= layer4_outputs(1391);
    layer5_outputs(1644) <= (layer4_outputs(987)) and (layer4_outputs(1656));
    layer5_outputs(1645) <= (layer4_outputs(1058)) and not (layer4_outputs(750));
    layer5_outputs(1646) <= not((layer4_outputs(1033)) or (layer4_outputs(2522)));
    layer5_outputs(1647) <= not(layer4_outputs(799));
    layer5_outputs(1648) <= layer4_outputs(1490);
    layer5_outputs(1649) <= layer4_outputs(1087);
    layer5_outputs(1650) <= (layer4_outputs(2388)) and not (layer4_outputs(1040));
    layer5_outputs(1651) <= (layer4_outputs(1659)) and not (layer4_outputs(2100));
    layer5_outputs(1652) <= (layer4_outputs(2352)) or (layer4_outputs(907));
    layer5_outputs(1653) <= layer4_outputs(1613);
    layer5_outputs(1654) <= (layer4_outputs(613)) or (layer4_outputs(2174));
    layer5_outputs(1655) <= (layer4_outputs(1838)) and not (layer4_outputs(2070));
    layer5_outputs(1656) <= not(layer4_outputs(1579));
    layer5_outputs(1657) <= (layer4_outputs(2017)) and not (layer4_outputs(2192));
    layer5_outputs(1658) <= layer4_outputs(2381);
    layer5_outputs(1659) <= layer4_outputs(1721);
    layer5_outputs(1660) <= not(layer4_outputs(1151));
    layer5_outputs(1661) <= (layer4_outputs(57)) or (layer4_outputs(2108));
    layer5_outputs(1662) <= not((layer4_outputs(2115)) and (layer4_outputs(201)));
    layer5_outputs(1663) <= not(layer4_outputs(73));
    layer5_outputs(1664) <= not(layer4_outputs(523)) or (layer4_outputs(1871));
    layer5_outputs(1665) <= (layer4_outputs(1465)) and not (layer4_outputs(1611));
    layer5_outputs(1666) <= not(layer4_outputs(2081));
    layer5_outputs(1667) <= layer4_outputs(1572);
    layer5_outputs(1668) <= not((layer4_outputs(519)) xor (layer4_outputs(2549)));
    layer5_outputs(1669) <= not(layer4_outputs(767));
    layer5_outputs(1670) <= not(layer4_outputs(1880)) or (layer4_outputs(377));
    layer5_outputs(1671) <= not(layer4_outputs(685));
    layer5_outputs(1672) <= (layer4_outputs(869)) or (layer4_outputs(1650));
    layer5_outputs(1673) <= (layer4_outputs(1714)) and (layer4_outputs(247));
    layer5_outputs(1674) <= layer4_outputs(2415);
    layer5_outputs(1675) <= (layer4_outputs(655)) xor (layer4_outputs(1742));
    layer5_outputs(1676) <= layer4_outputs(1983);
    layer5_outputs(1677) <= (layer4_outputs(2501)) and not (layer4_outputs(1605));
    layer5_outputs(1678) <= not((layer4_outputs(1692)) xor (layer4_outputs(1668)));
    layer5_outputs(1679) <= not(layer4_outputs(489));
    layer5_outputs(1680) <= not(layer4_outputs(478));
    layer5_outputs(1681) <= (layer4_outputs(1481)) and (layer4_outputs(1112));
    layer5_outputs(1682) <= layer4_outputs(648);
    layer5_outputs(1683) <= not(layer4_outputs(2335));
    layer5_outputs(1684) <= not(layer4_outputs(306));
    layer5_outputs(1685) <= (layer4_outputs(1552)) and not (layer4_outputs(2037));
    layer5_outputs(1686) <= layer4_outputs(160);
    layer5_outputs(1687) <= (layer4_outputs(1424)) and not (layer4_outputs(80));
    layer5_outputs(1688) <= not((layer4_outputs(146)) or (layer4_outputs(1661)));
    layer5_outputs(1689) <= layer4_outputs(1518);
    layer5_outputs(1690) <= not(layer4_outputs(2187));
    layer5_outputs(1691) <= layer4_outputs(1298);
    layer5_outputs(1692) <= not(layer4_outputs(1267));
    layer5_outputs(1693) <= layer4_outputs(1667);
    layer5_outputs(1694) <= not(layer4_outputs(1905));
    layer5_outputs(1695) <= (layer4_outputs(2276)) and not (layer4_outputs(1418));
    layer5_outputs(1696) <= '0';
    layer5_outputs(1697) <= not((layer4_outputs(1326)) and (layer4_outputs(1117)));
    layer5_outputs(1698) <= not(layer4_outputs(2267));
    layer5_outputs(1699) <= '1';
    layer5_outputs(1700) <= not(layer4_outputs(560));
    layer5_outputs(1701) <= not(layer4_outputs(494)) or (layer4_outputs(2237));
    layer5_outputs(1702) <= not(layer4_outputs(490));
    layer5_outputs(1703) <= '1';
    layer5_outputs(1704) <= not((layer4_outputs(319)) or (layer4_outputs(816)));
    layer5_outputs(1705) <= not((layer4_outputs(951)) or (layer4_outputs(2086)));
    layer5_outputs(1706) <= not((layer4_outputs(2310)) and (layer4_outputs(736)));
    layer5_outputs(1707) <= layer4_outputs(111);
    layer5_outputs(1708) <= (layer4_outputs(1293)) xor (layer4_outputs(2309));
    layer5_outputs(1709) <= not((layer4_outputs(1154)) or (layer4_outputs(2432)));
    layer5_outputs(1710) <= (layer4_outputs(1420)) and not (layer4_outputs(217));
    layer5_outputs(1711) <= not(layer4_outputs(2141)) or (layer4_outputs(661));
    layer5_outputs(1712) <= (layer4_outputs(2122)) and not (layer4_outputs(1612));
    layer5_outputs(1713) <= not((layer4_outputs(1515)) and (layer4_outputs(1325)));
    layer5_outputs(1714) <= not((layer4_outputs(180)) and (layer4_outputs(214)));
    layer5_outputs(1715) <= not(layer4_outputs(1710)) or (layer4_outputs(104));
    layer5_outputs(1716) <= not(layer4_outputs(426));
    layer5_outputs(1717) <= layer4_outputs(1376);
    layer5_outputs(1718) <= (layer4_outputs(1174)) and (layer4_outputs(2371));
    layer5_outputs(1719) <= not(layer4_outputs(2430));
    layer5_outputs(1720) <= not((layer4_outputs(1982)) and (layer4_outputs(358)));
    layer5_outputs(1721) <= '0';
    layer5_outputs(1722) <= (layer4_outputs(2300)) and (layer4_outputs(609));
    layer5_outputs(1723) <= (layer4_outputs(2014)) and not (layer4_outputs(1082));
    layer5_outputs(1724) <= (layer4_outputs(944)) or (layer4_outputs(1244));
    layer5_outputs(1725) <= not((layer4_outputs(1853)) and (layer4_outputs(1111)));
    layer5_outputs(1726) <= (layer4_outputs(1546)) or (layer4_outputs(1821));
    layer5_outputs(1727) <= layer4_outputs(1339);
    layer5_outputs(1728) <= not(layer4_outputs(162)) or (layer4_outputs(1055));
    layer5_outputs(1729) <= not(layer4_outputs(595));
    layer5_outputs(1730) <= not(layer4_outputs(284)) or (layer4_outputs(8));
    layer5_outputs(1731) <= not(layer4_outputs(1461));
    layer5_outputs(1732) <= not(layer4_outputs(1340)) or (layer4_outputs(1173));
    layer5_outputs(1733) <= not((layer4_outputs(1049)) or (layer4_outputs(1292)));
    layer5_outputs(1734) <= (layer4_outputs(881)) xor (layer4_outputs(2497));
    layer5_outputs(1735) <= '1';
    layer5_outputs(1736) <= layer4_outputs(1577);
    layer5_outputs(1737) <= not(layer4_outputs(1977));
    layer5_outputs(1738) <= layer4_outputs(2258);
    layer5_outputs(1739) <= layer4_outputs(2122);
    layer5_outputs(1740) <= not((layer4_outputs(2284)) xor (layer4_outputs(651)));
    layer5_outputs(1741) <= not((layer4_outputs(1789)) xor (layer4_outputs(849)));
    layer5_outputs(1742) <= layer4_outputs(2392);
    layer5_outputs(1743) <= layer4_outputs(1919);
    layer5_outputs(1744) <= layer4_outputs(2501);
    layer5_outputs(1745) <= not(layer4_outputs(2041));
    layer5_outputs(1746) <= not(layer4_outputs(2535));
    layer5_outputs(1747) <= layer4_outputs(2372);
    layer5_outputs(1748) <= '0';
    layer5_outputs(1749) <= layer4_outputs(1857);
    layer5_outputs(1750) <= layer4_outputs(570);
    layer5_outputs(1751) <= (layer4_outputs(1686)) and (layer4_outputs(298));
    layer5_outputs(1752) <= layer4_outputs(548);
    layer5_outputs(1753) <= not(layer4_outputs(2517));
    layer5_outputs(1754) <= (layer4_outputs(1860)) and not (layer4_outputs(590));
    layer5_outputs(1755) <= not((layer4_outputs(2478)) or (layer4_outputs(216)));
    layer5_outputs(1756) <= (layer4_outputs(30)) or (layer4_outputs(1442));
    layer5_outputs(1757) <= (layer4_outputs(92)) or (layer4_outputs(954));
    layer5_outputs(1758) <= not(layer4_outputs(1859));
    layer5_outputs(1759) <= not(layer4_outputs(753));
    layer5_outputs(1760) <= '1';
    layer5_outputs(1761) <= layer4_outputs(2129);
    layer5_outputs(1762) <= layer4_outputs(1344);
    layer5_outputs(1763) <= '1';
    layer5_outputs(1764) <= (layer4_outputs(2192)) and (layer4_outputs(679));
    layer5_outputs(1765) <= not(layer4_outputs(1707)) or (layer4_outputs(200));
    layer5_outputs(1766) <= not(layer4_outputs(943));
    layer5_outputs(1767) <= layer4_outputs(2262);
    layer5_outputs(1768) <= (layer4_outputs(1835)) and not (layer4_outputs(373));
    layer5_outputs(1769) <= not(layer4_outputs(632));
    layer5_outputs(1770) <= layer4_outputs(56);
    layer5_outputs(1771) <= layer4_outputs(1359);
    layer5_outputs(1772) <= not(layer4_outputs(1825));
    layer5_outputs(1773) <= (layer4_outputs(336)) and not (layer4_outputs(2496));
    layer5_outputs(1774) <= layer4_outputs(2286);
    layer5_outputs(1775) <= layer4_outputs(1930);
    layer5_outputs(1776) <= not((layer4_outputs(1709)) and (layer4_outputs(1297)));
    layer5_outputs(1777) <= layer4_outputs(285);
    layer5_outputs(1778) <= (layer4_outputs(592)) or (layer4_outputs(1409));
    layer5_outputs(1779) <= not(layer4_outputs(8));
    layer5_outputs(1780) <= not(layer4_outputs(1109)) or (layer4_outputs(2307));
    layer5_outputs(1781) <= not(layer4_outputs(2312));
    layer5_outputs(1782) <= layer4_outputs(1166);
    layer5_outputs(1783) <= layer4_outputs(2127);
    layer5_outputs(1784) <= '1';
    layer5_outputs(1785) <= not((layer4_outputs(567)) and (layer4_outputs(2468)));
    layer5_outputs(1786) <= not((layer4_outputs(1948)) and (layer4_outputs(356)));
    layer5_outputs(1787) <= not(layer4_outputs(544));
    layer5_outputs(1788) <= not(layer4_outputs(855));
    layer5_outputs(1789) <= (layer4_outputs(213)) and (layer4_outputs(127));
    layer5_outputs(1790) <= not((layer4_outputs(1809)) or (layer4_outputs(1811)));
    layer5_outputs(1791) <= not(layer4_outputs(939));
    layer5_outputs(1792) <= layer4_outputs(312);
    layer5_outputs(1793) <= not((layer4_outputs(623)) or (layer4_outputs(2031)));
    layer5_outputs(1794) <= not(layer4_outputs(1897));
    layer5_outputs(1795) <= layer4_outputs(954);
    layer5_outputs(1796) <= layer4_outputs(2131);
    layer5_outputs(1797) <= (layer4_outputs(2409)) and (layer4_outputs(2431));
    layer5_outputs(1798) <= not(layer4_outputs(522)) or (layer4_outputs(441));
    layer5_outputs(1799) <= layer4_outputs(1397);
    layer5_outputs(1800) <= layer4_outputs(887);
    layer5_outputs(1801) <= not(layer4_outputs(626));
    layer5_outputs(1802) <= not(layer4_outputs(138));
    layer5_outputs(1803) <= not(layer4_outputs(1814)) or (layer4_outputs(1075));
    layer5_outputs(1804) <= not((layer4_outputs(1323)) and (layer4_outputs(7)));
    layer5_outputs(1805) <= not(layer4_outputs(2111)) or (layer4_outputs(4));
    layer5_outputs(1806) <= (layer4_outputs(990)) or (layer4_outputs(41));
    layer5_outputs(1807) <= layer4_outputs(1717);
    layer5_outputs(1808) <= not(layer4_outputs(323));
    layer5_outputs(1809) <= not((layer4_outputs(713)) or (layer4_outputs(1202)));
    layer5_outputs(1810) <= (layer4_outputs(484)) and not (layer4_outputs(112));
    layer5_outputs(1811) <= layer4_outputs(1280);
    layer5_outputs(1812) <= layer4_outputs(1493);
    layer5_outputs(1813) <= (layer4_outputs(2429)) xor (layer4_outputs(1471));
    layer5_outputs(1814) <= not(layer4_outputs(2071)) or (layer4_outputs(583));
    layer5_outputs(1815) <= not(layer4_outputs(460));
    layer5_outputs(1816) <= not((layer4_outputs(2434)) and (layer4_outputs(429)));
    layer5_outputs(1817) <= (layer4_outputs(1105)) and not (layer4_outputs(1266));
    layer5_outputs(1818) <= not(layer4_outputs(1707));
    layer5_outputs(1819) <= (layer4_outputs(2143)) xor (layer4_outputs(2190));
    layer5_outputs(1820) <= not(layer4_outputs(2438));
    layer5_outputs(1821) <= not((layer4_outputs(1294)) or (layer4_outputs(228)));
    layer5_outputs(1822) <= layer4_outputs(2439);
    layer5_outputs(1823) <= not(layer4_outputs(1280)) or (layer4_outputs(2217));
    layer5_outputs(1824) <= layer4_outputs(869);
    layer5_outputs(1825) <= not((layer4_outputs(856)) and (layer4_outputs(299)));
    layer5_outputs(1826) <= not(layer4_outputs(2468));
    layer5_outputs(1827) <= not(layer4_outputs(1289));
    layer5_outputs(1828) <= not(layer4_outputs(1925)) or (layer4_outputs(2450));
    layer5_outputs(1829) <= not(layer4_outputs(1132)) or (layer4_outputs(1456));
    layer5_outputs(1830) <= (layer4_outputs(2374)) and (layer4_outputs(227));
    layer5_outputs(1831) <= (layer4_outputs(795)) and (layer4_outputs(211));
    layer5_outputs(1832) <= not((layer4_outputs(810)) or (layer4_outputs(814)));
    layer5_outputs(1833) <= not(layer4_outputs(1543)) or (layer4_outputs(1200));
    layer5_outputs(1834) <= layer4_outputs(693);
    layer5_outputs(1835) <= (layer4_outputs(511)) or (layer4_outputs(2324));
    layer5_outputs(1836) <= not((layer4_outputs(420)) or (layer4_outputs(2148)));
    layer5_outputs(1837) <= layer4_outputs(1974);
    layer5_outputs(1838) <= not((layer4_outputs(2086)) and (layer4_outputs(880)));
    layer5_outputs(1839) <= (layer4_outputs(466)) and not (layer4_outputs(1931));
    layer5_outputs(1840) <= not(layer4_outputs(1306));
    layer5_outputs(1841) <= layer4_outputs(1035);
    layer5_outputs(1842) <= '0';
    layer5_outputs(1843) <= layer4_outputs(2365);
    layer5_outputs(1844) <= '0';
    layer5_outputs(1845) <= layer4_outputs(419);
    layer5_outputs(1846) <= not(layer4_outputs(852)) or (layer4_outputs(1870));
    layer5_outputs(1847) <= layer4_outputs(2255);
    layer5_outputs(1848) <= not(layer4_outputs(138));
    layer5_outputs(1849) <= not((layer4_outputs(1125)) xor (layer4_outputs(545)));
    layer5_outputs(1850) <= layer4_outputs(283);
    layer5_outputs(1851) <= not(layer4_outputs(794));
    layer5_outputs(1852) <= '0';
    layer5_outputs(1853) <= layer4_outputs(489);
    layer5_outputs(1854) <= not(layer4_outputs(1615));
    layer5_outputs(1855) <= layer4_outputs(259);
    layer5_outputs(1856) <= layer4_outputs(1935);
    layer5_outputs(1857) <= layer4_outputs(1316);
    layer5_outputs(1858) <= (layer4_outputs(875)) and not (layer4_outputs(1644));
    layer5_outputs(1859) <= '1';
    layer5_outputs(1860) <= layer4_outputs(2278);
    layer5_outputs(1861) <= not((layer4_outputs(1622)) xor (layer4_outputs(1037)));
    layer5_outputs(1862) <= '0';
    layer5_outputs(1863) <= (layer4_outputs(2130)) and not (layer4_outputs(1524));
    layer5_outputs(1864) <= (layer4_outputs(1628)) and not (layer4_outputs(1942));
    layer5_outputs(1865) <= layer4_outputs(2292);
    layer5_outputs(1866) <= not((layer4_outputs(386)) or (layer4_outputs(74)));
    layer5_outputs(1867) <= (layer4_outputs(59)) and (layer4_outputs(788));
    layer5_outputs(1868) <= not(layer4_outputs(1464));
    layer5_outputs(1869) <= not(layer4_outputs(604));
    layer5_outputs(1870) <= not((layer4_outputs(1643)) and (layer4_outputs(512)));
    layer5_outputs(1871) <= layer4_outputs(1526);
    layer5_outputs(1872) <= not(layer4_outputs(406)) or (layer4_outputs(879));
    layer5_outputs(1873) <= not((layer4_outputs(1158)) xor (layer4_outputs(741)));
    layer5_outputs(1874) <= (layer4_outputs(1317)) or (layer4_outputs(1645));
    layer5_outputs(1875) <= (layer4_outputs(1320)) and not (layer4_outputs(958));
    layer5_outputs(1876) <= (layer4_outputs(2459)) and not (layer4_outputs(2153));
    layer5_outputs(1877) <= not(layer4_outputs(1623));
    layer5_outputs(1878) <= (layer4_outputs(808)) and not (layer4_outputs(1989));
    layer5_outputs(1879) <= (layer4_outputs(2416)) and not (layer4_outputs(30));
    layer5_outputs(1880) <= layer4_outputs(790);
    layer5_outputs(1881) <= not(layer4_outputs(2438));
    layer5_outputs(1882) <= layer4_outputs(2460);
    layer5_outputs(1883) <= not(layer4_outputs(785));
    layer5_outputs(1884) <= (layer4_outputs(2004)) and (layer4_outputs(1106));
    layer5_outputs(1885) <= layer4_outputs(1606);
    layer5_outputs(1886) <= layer4_outputs(1522);
    layer5_outputs(1887) <= not(layer4_outputs(965));
    layer5_outputs(1888) <= not(layer4_outputs(90));
    layer5_outputs(1889) <= not((layer4_outputs(1228)) and (layer4_outputs(887)));
    layer5_outputs(1890) <= not(layer4_outputs(950)) or (layer4_outputs(2433));
    layer5_outputs(1891) <= (layer4_outputs(2408)) or (layer4_outputs(625));
    layer5_outputs(1892) <= not(layer4_outputs(2503));
    layer5_outputs(1893) <= (layer4_outputs(2)) xor (layer4_outputs(2330));
    layer5_outputs(1894) <= not(layer4_outputs(616));
    layer5_outputs(1895) <= '1';
    layer5_outputs(1896) <= '1';
    layer5_outputs(1897) <= not(layer4_outputs(2301));
    layer5_outputs(1898) <= (layer4_outputs(334)) xor (layer4_outputs(515));
    layer5_outputs(1899) <= '0';
    layer5_outputs(1900) <= layer4_outputs(1926);
    layer5_outputs(1901) <= not(layer4_outputs(111));
    layer5_outputs(1902) <= not(layer4_outputs(2245));
    layer5_outputs(1903) <= '0';
    layer5_outputs(1904) <= not(layer4_outputs(1923));
    layer5_outputs(1905) <= (layer4_outputs(2343)) and not (layer4_outputs(2048));
    layer5_outputs(1906) <= (layer4_outputs(1380)) and not (layer4_outputs(1649));
    layer5_outputs(1907) <= not(layer4_outputs(1874));
    layer5_outputs(1908) <= layer4_outputs(1663);
    layer5_outputs(1909) <= layer4_outputs(1651);
    layer5_outputs(1910) <= not(layer4_outputs(1966));
    layer5_outputs(1911) <= (layer4_outputs(2033)) and (layer4_outputs(603));
    layer5_outputs(1912) <= not(layer4_outputs(1365));
    layer5_outputs(1913) <= not(layer4_outputs(828)) or (layer4_outputs(804));
    layer5_outputs(1914) <= not(layer4_outputs(2242));
    layer5_outputs(1915) <= not(layer4_outputs(796));
    layer5_outputs(1916) <= not((layer4_outputs(1125)) and (layer4_outputs(975)));
    layer5_outputs(1917) <= '1';
    layer5_outputs(1918) <= layer4_outputs(17);
    layer5_outputs(1919) <= not(layer4_outputs(1338)) or (layer4_outputs(934));
    layer5_outputs(1920) <= layer4_outputs(1350);
    layer5_outputs(1921) <= not((layer4_outputs(316)) and (layer4_outputs(2219)));
    layer5_outputs(1922) <= not((layer4_outputs(2018)) xor (layer4_outputs(125)));
    layer5_outputs(1923) <= not(layer4_outputs(727)) or (layer4_outputs(2247));
    layer5_outputs(1924) <= (layer4_outputs(1565)) and not (layer4_outputs(1770));
    layer5_outputs(1925) <= not(layer4_outputs(1533));
    layer5_outputs(1926) <= (layer4_outputs(115)) and not (layer4_outputs(338));
    layer5_outputs(1927) <= not((layer4_outputs(101)) xor (layer4_outputs(409)));
    layer5_outputs(1928) <= layer4_outputs(1940);
    layer5_outputs(1929) <= (layer4_outputs(371)) xor (layer4_outputs(428));
    layer5_outputs(1930) <= not(layer4_outputs(1725));
    layer5_outputs(1931) <= layer4_outputs(2046);
    layer5_outputs(1932) <= layer4_outputs(812);
    layer5_outputs(1933) <= not(layer4_outputs(2486));
    layer5_outputs(1934) <= not(layer4_outputs(1964)) or (layer4_outputs(552));
    layer5_outputs(1935) <= (layer4_outputs(712)) xor (layer4_outputs(2448));
    layer5_outputs(1936) <= '1';
    layer5_outputs(1937) <= layer4_outputs(2197);
    layer5_outputs(1938) <= not((layer4_outputs(1719)) xor (layer4_outputs(1655)));
    layer5_outputs(1939) <= layer4_outputs(1000);
    layer5_outputs(1940) <= (layer4_outputs(2377)) and not (layer4_outputs(1043));
    layer5_outputs(1941) <= (layer4_outputs(1542)) and not (layer4_outputs(662));
    layer5_outputs(1942) <= not(layer4_outputs(713)) or (layer4_outputs(955));
    layer5_outputs(1943) <= '0';
    layer5_outputs(1944) <= (layer4_outputs(1544)) xor (layer4_outputs(236));
    layer5_outputs(1945) <= not(layer4_outputs(646));
    layer5_outputs(1946) <= not(layer4_outputs(282));
    layer5_outputs(1947) <= not(layer4_outputs(1189));
    layer5_outputs(1948) <= (layer4_outputs(915)) or (layer4_outputs(2406));
    layer5_outputs(1949) <= not((layer4_outputs(1041)) and (layer4_outputs(1111)));
    layer5_outputs(1950) <= layer4_outputs(1237);
    layer5_outputs(1951) <= not(layer4_outputs(683));
    layer5_outputs(1952) <= not((layer4_outputs(300)) xor (layer4_outputs(1165)));
    layer5_outputs(1953) <= not((layer4_outputs(2490)) xor (layer4_outputs(189)));
    layer5_outputs(1954) <= layer4_outputs(1338);
    layer5_outputs(1955) <= (layer4_outputs(2105)) and (layer4_outputs(852));
    layer5_outputs(1956) <= '1';
    layer5_outputs(1957) <= layer4_outputs(379);
    layer5_outputs(1958) <= (layer4_outputs(699)) and not (layer4_outputs(1113));
    layer5_outputs(1959) <= layer4_outputs(1474);
    layer5_outputs(1960) <= (layer4_outputs(1181)) xor (layer4_outputs(1703));
    layer5_outputs(1961) <= not(layer4_outputs(172));
    layer5_outputs(1962) <= not(layer4_outputs(781));
    layer5_outputs(1963) <= layer4_outputs(453);
    layer5_outputs(1964) <= layer4_outputs(2185);
    layer5_outputs(1965) <= layer4_outputs(846);
    layer5_outputs(1966) <= not(layer4_outputs(643));
    layer5_outputs(1967) <= not((layer4_outputs(303)) xor (layer4_outputs(1910)));
    layer5_outputs(1968) <= layer4_outputs(1618);
    layer5_outputs(1969) <= layer4_outputs(432);
    layer5_outputs(1970) <= not(layer4_outputs(1519)) or (layer4_outputs(2295));
    layer5_outputs(1971) <= not((layer4_outputs(2091)) or (layer4_outputs(449)));
    layer5_outputs(1972) <= (layer4_outputs(1321)) and not (layer4_outputs(1184));
    layer5_outputs(1973) <= (layer4_outputs(653)) or (layer4_outputs(1561));
    layer5_outputs(1974) <= not(layer4_outputs(680));
    layer5_outputs(1975) <= not((layer4_outputs(474)) or (layer4_outputs(1724)));
    layer5_outputs(1976) <= '1';
    layer5_outputs(1977) <= not((layer4_outputs(768)) and (layer4_outputs(2458)));
    layer5_outputs(1978) <= not((layer4_outputs(344)) and (layer4_outputs(1848)));
    layer5_outputs(1979) <= not(layer4_outputs(1748));
    layer5_outputs(1980) <= not((layer4_outputs(1590)) and (layer4_outputs(159)));
    layer5_outputs(1981) <= (layer4_outputs(825)) and (layer4_outputs(2516));
    layer5_outputs(1982) <= layer4_outputs(132);
    layer5_outputs(1983) <= not(layer4_outputs(2177));
    layer5_outputs(1984) <= not(layer4_outputs(2531));
    layer5_outputs(1985) <= (layer4_outputs(1903)) and not (layer4_outputs(717));
    layer5_outputs(1986) <= not(layer4_outputs(1501));
    layer5_outputs(1987) <= not(layer4_outputs(2254));
    layer5_outputs(1988) <= (layer4_outputs(873)) and (layer4_outputs(1098));
    layer5_outputs(1989) <= layer4_outputs(269);
    layer5_outputs(1990) <= not(layer4_outputs(667));
    layer5_outputs(1991) <= not(layer4_outputs(704)) or (layer4_outputs(1256));
    layer5_outputs(1992) <= (layer4_outputs(2095)) and not (layer4_outputs(1702));
    layer5_outputs(1993) <= (layer4_outputs(539)) and not (layer4_outputs(514));
    layer5_outputs(1994) <= not((layer4_outputs(997)) and (layer4_outputs(1238)));
    layer5_outputs(1995) <= not(layer4_outputs(1159));
    layer5_outputs(1996) <= not(layer4_outputs(2243)) or (layer4_outputs(1458));
    layer5_outputs(1997) <= (layer4_outputs(1285)) or (layer4_outputs(173));
    layer5_outputs(1998) <= (layer4_outputs(1102)) or (layer4_outputs(899));
    layer5_outputs(1999) <= not(layer4_outputs(1462)) or (layer4_outputs(1623));
    layer5_outputs(2000) <= layer4_outputs(1988);
    layer5_outputs(2001) <= not((layer4_outputs(302)) xor (layer4_outputs(1764)));
    layer5_outputs(2002) <= (layer4_outputs(307)) and not (layer4_outputs(2409));
    layer5_outputs(2003) <= layer4_outputs(322);
    layer5_outputs(2004) <= '1';
    layer5_outputs(2005) <= (layer4_outputs(194)) or (layer4_outputs(2051));
    layer5_outputs(2006) <= (layer4_outputs(892)) and not (layer4_outputs(913));
    layer5_outputs(2007) <= layer4_outputs(1467);
    layer5_outputs(2008) <= not((layer4_outputs(77)) xor (layer4_outputs(841)));
    layer5_outputs(2009) <= '0';
    layer5_outputs(2010) <= not((layer4_outputs(2497)) xor (layer4_outputs(1619)));
    layer5_outputs(2011) <= layer4_outputs(314);
    layer5_outputs(2012) <= not(layer4_outputs(1143));
    layer5_outputs(2013) <= layer4_outputs(513);
    layer5_outputs(2014) <= not(layer4_outputs(2369));
    layer5_outputs(2015) <= '0';
    layer5_outputs(2016) <= layer4_outputs(1432);
    layer5_outputs(2017) <= layer4_outputs(2144);
    layer5_outputs(2018) <= (layer4_outputs(752)) and (layer4_outputs(1285));
    layer5_outputs(2019) <= layer4_outputs(1890);
    layer5_outputs(2020) <= not(layer4_outputs(1529));
    layer5_outputs(2021) <= (layer4_outputs(1642)) and not (layer4_outputs(1172));
    layer5_outputs(2022) <= not((layer4_outputs(42)) and (layer4_outputs(2185)));
    layer5_outputs(2023) <= (layer4_outputs(471)) and not (layer4_outputs(1086));
    layer5_outputs(2024) <= layer4_outputs(1700);
    layer5_outputs(2025) <= layer4_outputs(688);
    layer5_outputs(2026) <= not(layer4_outputs(1877));
    layer5_outputs(2027) <= layer4_outputs(607);
    layer5_outputs(2028) <= (layer4_outputs(1774)) xor (layer4_outputs(462));
    layer5_outputs(2029) <= not(layer4_outputs(1555));
    layer5_outputs(2030) <= not(layer4_outputs(843));
    layer5_outputs(2031) <= not(layer4_outputs(3)) or (layer4_outputs(537));
    layer5_outputs(2032) <= (layer4_outputs(2394)) and (layer4_outputs(473));
    layer5_outputs(2033) <= not(layer4_outputs(1933)) or (layer4_outputs(1142));
    layer5_outputs(2034) <= (layer4_outputs(1948)) and not (layer4_outputs(1796));
    layer5_outputs(2035) <= not(layer4_outputs(1912));
    layer5_outputs(2036) <= layer4_outputs(1305);
    layer5_outputs(2037) <= (layer4_outputs(1844)) or (layer4_outputs(2362));
    layer5_outputs(2038) <= layer4_outputs(2023);
    layer5_outputs(2039) <= layer4_outputs(1621);
    layer5_outputs(2040) <= not(layer4_outputs(773)) or (layer4_outputs(558));
    layer5_outputs(2041) <= layer4_outputs(890);
    layer5_outputs(2042) <= (layer4_outputs(1803)) or (layer4_outputs(2151));
    layer5_outputs(2043) <= layer4_outputs(2081);
    layer5_outputs(2044) <= layer4_outputs(622);
    layer5_outputs(2045) <= not((layer4_outputs(548)) xor (layer4_outputs(2494)));
    layer5_outputs(2046) <= layer4_outputs(975);
    layer5_outputs(2047) <= (layer4_outputs(147)) or (layer4_outputs(1981));
    layer5_outputs(2048) <= not((layer4_outputs(1810)) and (layer4_outputs(1203)));
    layer5_outputs(2049) <= not(layer4_outputs(578));
    layer5_outputs(2050) <= layer4_outputs(583);
    layer5_outputs(2051) <= not((layer4_outputs(2470)) or (layer4_outputs(488)));
    layer5_outputs(2052) <= not((layer4_outputs(1842)) or (layer4_outputs(527)));
    layer5_outputs(2053) <= not(layer4_outputs(1218));
    layer5_outputs(2054) <= not((layer4_outputs(540)) and (layer4_outputs(612)));
    layer5_outputs(2055) <= not((layer4_outputs(2524)) or (layer4_outputs(2051)));
    layer5_outputs(2056) <= not(layer4_outputs(2201));
    layer5_outputs(2057) <= layer4_outputs(1509);
    layer5_outputs(2058) <= not((layer4_outputs(275)) xor (layer4_outputs(1568)));
    layer5_outputs(2059) <= not(layer4_outputs(2096)) or (layer4_outputs(2279));
    layer5_outputs(2060) <= not(layer4_outputs(1807));
    layer5_outputs(2061) <= not(layer4_outputs(1734));
    layer5_outputs(2062) <= (layer4_outputs(2440)) or (layer4_outputs(2239));
    layer5_outputs(2063) <= (layer4_outputs(658)) xor (layer4_outputs(1500));
    layer5_outputs(2064) <= (layer4_outputs(328)) and not (layer4_outputs(507));
    layer5_outputs(2065) <= (layer4_outputs(2034)) or (layer4_outputs(2527));
    layer5_outputs(2066) <= not(layer4_outputs(617));
    layer5_outputs(2067) <= layer4_outputs(911);
    layer5_outputs(2068) <= layer4_outputs(1020);
    layer5_outputs(2069) <= (layer4_outputs(1411)) or (layer4_outputs(1370));
    layer5_outputs(2070) <= not((layer4_outputs(801)) and (layer4_outputs(1614)));
    layer5_outputs(2071) <= not(layer4_outputs(1514));
    layer5_outputs(2072) <= (layer4_outputs(2300)) and (layer4_outputs(877));
    layer5_outputs(2073) <= layer4_outputs(1576);
    layer5_outputs(2074) <= not(layer4_outputs(1435));
    layer5_outputs(2075) <= layer4_outputs(2147);
    layer5_outputs(2076) <= not(layer4_outputs(1264)) or (layer4_outputs(532));
    layer5_outputs(2077) <= not(layer4_outputs(163)) or (layer4_outputs(705));
    layer5_outputs(2078) <= not((layer4_outputs(1676)) and (layer4_outputs(615)));
    layer5_outputs(2079) <= '1';
    layer5_outputs(2080) <= '1';
    layer5_outputs(2081) <= layer4_outputs(1688);
    layer5_outputs(2082) <= (layer4_outputs(26)) and (layer4_outputs(1291));
    layer5_outputs(2083) <= not((layer4_outputs(494)) and (layer4_outputs(273)));
    layer5_outputs(2084) <= (layer4_outputs(156)) or (layer4_outputs(418));
    layer5_outputs(2085) <= not((layer4_outputs(966)) xor (layer4_outputs(1578)));
    layer5_outputs(2086) <= (layer4_outputs(364)) and not (layer4_outputs(872));
    layer5_outputs(2087) <= (layer4_outputs(2384)) and not (layer4_outputs(31));
    layer5_outputs(2088) <= (layer4_outputs(1206)) or (layer4_outputs(2289));
    layer5_outputs(2089) <= not(layer4_outputs(2060));
    layer5_outputs(2090) <= (layer4_outputs(2134)) and (layer4_outputs(1509));
    layer5_outputs(2091) <= not(layer4_outputs(511));
    layer5_outputs(2092) <= layer4_outputs(1813);
    layer5_outputs(2093) <= layer4_outputs(1106);
    layer5_outputs(2094) <= (layer4_outputs(108)) and not (layer4_outputs(227));
    layer5_outputs(2095) <= not((layer4_outputs(989)) and (layer4_outputs(1414)));
    layer5_outputs(2096) <= not(layer4_outputs(1516));
    layer5_outputs(2097) <= layer4_outputs(1247);
    layer5_outputs(2098) <= layer4_outputs(1164);
    layer5_outputs(2099) <= (layer4_outputs(1)) and not (layer4_outputs(1253));
    layer5_outputs(2100) <= layer4_outputs(729);
    layer5_outputs(2101) <= layer4_outputs(2379);
    layer5_outputs(2102) <= not(layer4_outputs(226));
    layer5_outputs(2103) <= layer4_outputs(554);
    layer5_outputs(2104) <= layer4_outputs(1187);
    layer5_outputs(2105) <= '0';
    layer5_outputs(2106) <= layer4_outputs(1939);
    layer5_outputs(2107) <= not(layer4_outputs(2010));
    layer5_outputs(2108) <= not((layer4_outputs(2020)) or (layer4_outputs(572)));
    layer5_outputs(2109) <= not(layer4_outputs(844));
    layer5_outputs(2110) <= not(layer4_outputs(620));
    layer5_outputs(2111) <= (layer4_outputs(386)) xor (layer4_outputs(1888));
    layer5_outputs(2112) <= not(layer4_outputs(2206));
    layer5_outputs(2113) <= not(layer4_outputs(2473)) or (layer4_outputs(1978));
    layer5_outputs(2114) <= (layer4_outputs(1556)) and not (layer4_outputs(2039));
    layer5_outputs(2115) <= (layer4_outputs(2026)) or (layer4_outputs(883));
    layer5_outputs(2116) <= not(layer4_outputs(1302));
    layer5_outputs(2117) <= '1';
    layer5_outputs(2118) <= not(layer4_outputs(357)) or (layer4_outputs(2213));
    layer5_outputs(2119) <= layer4_outputs(2229);
    layer5_outputs(2120) <= not((layer4_outputs(272)) or (layer4_outputs(1865)));
    layer5_outputs(2121) <= layer4_outputs(1731);
    layer5_outputs(2122) <= not((layer4_outputs(1366)) or (layer4_outputs(134)));
    layer5_outputs(2123) <= layer4_outputs(1586);
    layer5_outputs(2124) <= (layer4_outputs(917)) and (layer4_outputs(920));
    layer5_outputs(2125) <= not((layer4_outputs(1829)) or (layer4_outputs(645)));
    layer5_outputs(2126) <= not(layer4_outputs(1745)) or (layer4_outputs(1934));
    layer5_outputs(2127) <= (layer4_outputs(1984)) and (layer4_outputs(740));
    layer5_outputs(2128) <= layer4_outputs(2545);
    layer5_outputs(2129) <= not((layer4_outputs(2308)) xor (layer4_outputs(22)));
    layer5_outputs(2130) <= layer4_outputs(1139);
    layer5_outputs(2131) <= not(layer4_outputs(2447));
    layer5_outputs(2132) <= layer4_outputs(1697);
    layer5_outputs(2133) <= not(layer4_outputs(289));
    layer5_outputs(2134) <= not(layer4_outputs(1046));
    layer5_outputs(2135) <= not(layer4_outputs(361));
    layer5_outputs(2136) <= not(layer4_outputs(1755));
    layer5_outputs(2137) <= layer4_outputs(2218);
    layer5_outputs(2138) <= layer4_outputs(48);
    layer5_outputs(2139) <= (layer4_outputs(1875)) and not (layer4_outputs(1567));
    layer5_outputs(2140) <= not(layer4_outputs(452)) or (layer4_outputs(979));
    layer5_outputs(2141) <= not((layer4_outputs(2349)) and (layer4_outputs(1267)));
    layer5_outputs(2142) <= not(layer4_outputs(1351)) or (layer4_outputs(939));
    layer5_outputs(2143) <= not(layer4_outputs(315));
    layer5_outputs(2144) <= not(layer4_outputs(1812)) or (layer4_outputs(2149));
    layer5_outputs(2145) <= layer4_outputs(972);
    layer5_outputs(2146) <= layer4_outputs(1672);
    layer5_outputs(2147) <= '1';
    layer5_outputs(2148) <= layer4_outputs(1843);
    layer5_outputs(2149) <= '0';
    layer5_outputs(2150) <= (layer4_outputs(1929)) and not (layer4_outputs(2181));
    layer5_outputs(2151) <= not(layer4_outputs(467));
    layer5_outputs(2152) <= (layer4_outputs(929)) and (layer4_outputs(1664));
    layer5_outputs(2153) <= layer4_outputs(273);
    layer5_outputs(2154) <= layer4_outputs(1609);
    layer5_outputs(2155) <= not(layer4_outputs(1421));
    layer5_outputs(2156) <= (layer4_outputs(88)) and not (layer4_outputs(113));
    layer5_outputs(2157) <= (layer4_outputs(333)) and not (layer4_outputs(351));
    layer5_outputs(2158) <= (layer4_outputs(2174)) and (layer4_outputs(401));
    layer5_outputs(2159) <= (layer4_outputs(993)) xor (layer4_outputs(143));
    layer5_outputs(2160) <= layer4_outputs(262);
    layer5_outputs(2161) <= '0';
    layer5_outputs(2162) <= (layer4_outputs(1281)) or (layer4_outputs(2482));
    layer5_outputs(2163) <= (layer4_outputs(2353)) and not (layer4_outputs(1129));
    layer5_outputs(2164) <= '1';
    layer5_outputs(2165) <= not((layer4_outputs(1610)) and (layer4_outputs(1472)));
    layer5_outputs(2166) <= (layer4_outputs(1523)) and (layer4_outputs(1177));
    layer5_outputs(2167) <= not(layer4_outputs(1775));
    layer5_outputs(2168) <= layer4_outputs(2250);
    layer5_outputs(2169) <= not(layer4_outputs(435));
    layer5_outputs(2170) <= (layer4_outputs(2093)) and not (layer4_outputs(1014));
    layer5_outputs(2171) <= not((layer4_outputs(1451)) or (layer4_outputs(1793)));
    layer5_outputs(2172) <= not(layer4_outputs(2161));
    layer5_outputs(2173) <= not(layer4_outputs(561)) or (layer4_outputs(2271));
    layer5_outputs(2174) <= layer4_outputs(2461);
    layer5_outputs(2175) <= layer4_outputs(1222);
    layer5_outputs(2176) <= layer4_outputs(2049);
    layer5_outputs(2177) <= not((layer4_outputs(848)) xor (layer4_outputs(1353)));
    layer5_outputs(2178) <= not(layer4_outputs(597)) or (layer4_outputs(1537));
    layer5_outputs(2179) <= (layer4_outputs(1072)) and not (layer4_outputs(1251));
    layer5_outputs(2180) <= layer4_outputs(807);
    layer5_outputs(2181) <= (layer4_outputs(2477)) xor (layer4_outputs(2488));
    layer5_outputs(2182) <= not(layer4_outputs(1804));
    layer5_outputs(2183) <= '0';
    layer5_outputs(2184) <= not(layer4_outputs(2538));
    layer5_outputs(2185) <= not(layer4_outputs(1804));
    layer5_outputs(2186) <= not(layer4_outputs(1889));
    layer5_outputs(2187) <= not(layer4_outputs(1980));
    layer5_outputs(2188) <= not(layer4_outputs(57)) or (layer4_outputs(1024));
    layer5_outputs(2189) <= layer4_outputs(1218);
    layer5_outputs(2190) <= '0';
    layer5_outputs(2191) <= not(layer4_outputs(679));
    layer5_outputs(2192) <= (layer4_outputs(1792)) xor (layer4_outputs(423));
    layer5_outputs(2193) <= layer4_outputs(2383);
    layer5_outputs(2194) <= (layer4_outputs(2087)) and (layer4_outputs(2348));
    layer5_outputs(2195) <= layer4_outputs(2299);
    layer5_outputs(2196) <= layer4_outputs(1965);
    layer5_outputs(2197) <= not((layer4_outputs(1663)) and (layer4_outputs(2506)));
    layer5_outputs(2198) <= not(layer4_outputs(1066));
    layer5_outputs(2199) <= not(layer4_outputs(167));
    layer5_outputs(2200) <= layer4_outputs(715);
    layer5_outputs(2201) <= (layer4_outputs(1219)) and (layer4_outputs(493));
    layer5_outputs(2202) <= layer4_outputs(940);
    layer5_outputs(2203) <= layer4_outputs(1866);
    layer5_outputs(2204) <= (layer4_outputs(923)) or (layer4_outputs(1778));
    layer5_outputs(2205) <= (layer4_outputs(2474)) and (layer4_outputs(561));
    layer5_outputs(2206) <= (layer4_outputs(717)) and not (layer4_outputs(1750));
    layer5_outputs(2207) <= not(layer4_outputs(2232));
    layer5_outputs(2208) <= (layer4_outputs(27)) and (layer4_outputs(798));
    layer5_outputs(2209) <= not(layer4_outputs(2237));
    layer5_outputs(2210) <= not((layer4_outputs(1291)) or (layer4_outputs(1651)));
    layer5_outputs(2211) <= not(layer4_outputs(2244));
    layer5_outputs(2212) <= not(layer4_outputs(745)) or (layer4_outputs(1954));
    layer5_outputs(2213) <= not(layer4_outputs(524));
    layer5_outputs(2214) <= (layer4_outputs(1820)) or (layer4_outputs(368));
    layer5_outputs(2215) <= not(layer4_outputs(1031)) or (layer4_outputs(1229));
    layer5_outputs(2216) <= not(layer4_outputs(191));
    layer5_outputs(2217) <= layer4_outputs(1581);
    layer5_outputs(2218) <= layer4_outputs(1335);
    layer5_outputs(2219) <= not(layer4_outputs(589));
    layer5_outputs(2220) <= (layer4_outputs(1269)) and (layer4_outputs(2210));
    layer5_outputs(2221) <= layer4_outputs(1237);
    layer5_outputs(2222) <= not(layer4_outputs(1968));
    layer5_outputs(2223) <= (layer4_outputs(686)) or (layer4_outputs(1434));
    layer5_outputs(2224) <= '0';
    layer5_outputs(2225) <= layer4_outputs(2220);
    layer5_outputs(2226) <= (layer4_outputs(1677)) and not (layer4_outputs(823));
    layer5_outputs(2227) <= not(layer4_outputs(237));
    layer5_outputs(2228) <= not(layer4_outputs(1226));
    layer5_outputs(2229) <= layer4_outputs(208);
    layer5_outputs(2230) <= '1';
    layer5_outputs(2231) <= (layer4_outputs(994)) and not (layer4_outputs(2412));
    layer5_outputs(2232) <= not(layer4_outputs(1412)) or (layer4_outputs(135));
    layer5_outputs(2233) <= not(layer4_outputs(309)) or (layer4_outputs(1105));
    layer5_outputs(2234) <= not((layer4_outputs(164)) or (layer4_outputs(1811)));
    layer5_outputs(2235) <= not((layer4_outputs(1262)) and (layer4_outputs(435)));
    layer5_outputs(2236) <= layer4_outputs(388);
    layer5_outputs(2237) <= not((layer4_outputs(972)) or (layer4_outputs(499)));
    layer5_outputs(2238) <= not(layer4_outputs(97));
    layer5_outputs(2239) <= not(layer4_outputs(2107)) or (layer4_outputs(475));
    layer5_outputs(2240) <= not(layer4_outputs(705)) or (layer4_outputs(1580));
    layer5_outputs(2241) <= layer4_outputs(2466);
    layer5_outputs(2242) <= not(layer4_outputs(1958));
    layer5_outputs(2243) <= not(layer4_outputs(2425)) or (layer4_outputs(911));
    layer5_outputs(2244) <= (layer4_outputs(1085)) and not (layer4_outputs(1000));
    layer5_outputs(2245) <= not(layer4_outputs(1460));
    layer5_outputs(2246) <= not(layer4_outputs(2054)) or (layer4_outputs(1746));
    layer5_outputs(2247) <= (layer4_outputs(1592)) and (layer4_outputs(1359));
    layer5_outputs(2248) <= layer4_outputs(1662);
    layer5_outputs(2249) <= not((layer4_outputs(919)) and (layer4_outputs(992)));
    layer5_outputs(2250) <= (layer4_outputs(2487)) and not (layer4_outputs(36));
    layer5_outputs(2251) <= not(layer4_outputs(363));
    layer5_outputs(2252) <= not(layer4_outputs(781));
    layer5_outputs(2253) <= not(layer4_outputs(1079));
    layer5_outputs(2254) <= not(layer4_outputs(2289));
    layer5_outputs(2255) <= not(layer4_outputs(1215));
    layer5_outputs(2256) <= layer4_outputs(1912);
    layer5_outputs(2257) <= (layer4_outputs(1363)) and (layer4_outputs(1776));
    layer5_outputs(2258) <= not(layer4_outputs(563)) or (layer4_outputs(1201));
    layer5_outputs(2259) <= '0';
    layer5_outputs(2260) <= '0';
    layer5_outputs(2261) <= layer4_outputs(1276);
    layer5_outputs(2262) <= not((layer4_outputs(116)) and (layer4_outputs(1687)));
    layer5_outputs(2263) <= not(layer4_outputs(417));
    layer5_outputs(2264) <= not(layer4_outputs(1454)) or (layer4_outputs(1199));
    layer5_outputs(2265) <= layer4_outputs(2540);
    layer5_outputs(2266) <= (layer4_outputs(2539)) and (layer4_outputs(1850));
    layer5_outputs(2267) <= (layer4_outputs(1737)) or (layer4_outputs(947));
    layer5_outputs(2268) <= not(layer4_outputs(2395));
    layer5_outputs(2269) <= not(layer4_outputs(1592));
    layer5_outputs(2270) <= (layer4_outputs(1467)) and (layer4_outputs(871));
    layer5_outputs(2271) <= not(layer4_outputs(2491));
    layer5_outputs(2272) <= layer4_outputs(2195);
    layer5_outputs(2273) <= layer4_outputs(2338);
    layer5_outputs(2274) <= layer4_outputs(2509);
    layer5_outputs(2275) <= layer4_outputs(712);
    layer5_outputs(2276) <= layer4_outputs(2418);
    layer5_outputs(2277) <= layer4_outputs(1893);
    layer5_outputs(2278) <= not(layer4_outputs(366));
    layer5_outputs(2279) <= not(layer4_outputs(232));
    layer5_outputs(2280) <= layer4_outputs(875);
    layer5_outputs(2281) <= not((layer4_outputs(785)) or (layer4_outputs(627)));
    layer5_outputs(2282) <= not(layer4_outputs(1641));
    layer5_outputs(2283) <= not(layer4_outputs(1473));
    layer5_outputs(2284) <= not(layer4_outputs(658));
    layer5_outputs(2285) <= not((layer4_outputs(1810)) or (layer4_outputs(764)));
    layer5_outputs(2286) <= not(layer4_outputs(467));
    layer5_outputs(2287) <= (layer4_outputs(2475)) and not (layer4_outputs(347));
    layer5_outputs(2288) <= not(layer4_outputs(2423));
    layer5_outputs(2289) <= not(layer4_outputs(300)) or (layer4_outputs(110));
    layer5_outputs(2290) <= not((layer4_outputs(1386)) or (layer4_outputs(277)));
    layer5_outputs(2291) <= not(layer4_outputs(1261));
    layer5_outputs(2292) <= not(layer4_outputs(538));
    layer5_outputs(2293) <= layer4_outputs(2272);
    layer5_outputs(2294) <= not(layer4_outputs(1215));
    layer5_outputs(2295) <= not((layer4_outputs(1207)) or (layer4_outputs(1209)));
    layer5_outputs(2296) <= '0';
    layer5_outputs(2297) <= not((layer4_outputs(682)) and (layer4_outputs(2268)));
    layer5_outputs(2298) <= not(layer4_outputs(669)) or (layer4_outputs(1284));
    layer5_outputs(2299) <= layer4_outputs(89);
    layer5_outputs(2300) <= layer4_outputs(1907);
    layer5_outputs(2301) <= (layer4_outputs(1604)) and (layer4_outputs(480));
    layer5_outputs(2302) <= not((layer4_outputs(557)) or (layer4_outputs(2031)));
    layer5_outputs(2303) <= (layer4_outputs(543)) and not (layer4_outputs(1747));
    layer5_outputs(2304) <= layer4_outputs(751);
    layer5_outputs(2305) <= (layer4_outputs(1073)) and (layer4_outputs(815));
    layer5_outputs(2306) <= '0';
    layer5_outputs(2307) <= not(layer4_outputs(1298)) or (layer4_outputs(497));
    layer5_outputs(2308) <= not(layer4_outputs(502));
    layer5_outputs(2309) <= not(layer4_outputs(517));
    layer5_outputs(2310) <= '0';
    layer5_outputs(2311) <= (layer4_outputs(91)) and not (layer4_outputs(2545));
    layer5_outputs(2312) <= (layer4_outputs(1781)) and not (layer4_outputs(2356));
    layer5_outputs(2313) <= (layer4_outputs(1986)) and not (layer4_outputs(357));
    layer5_outputs(2314) <= layer4_outputs(906);
    layer5_outputs(2315) <= not(layer4_outputs(2538));
    layer5_outputs(2316) <= not(layer4_outputs(898));
    layer5_outputs(2317) <= (layer4_outputs(714)) and not (layer4_outputs(1504));
    layer5_outputs(2318) <= not(layer4_outputs(1960));
    layer5_outputs(2319) <= not(layer4_outputs(1128));
    layer5_outputs(2320) <= layer4_outputs(221);
    layer5_outputs(2321) <= not((layer4_outputs(2085)) xor (layer4_outputs(418)));
    layer5_outputs(2322) <= not(layer4_outputs(143));
    layer5_outputs(2323) <= layer4_outputs(1233);
    layer5_outputs(2324) <= layer4_outputs(528);
    layer5_outputs(2325) <= not(layer4_outputs(2160)) or (layer4_outputs(118));
    layer5_outputs(2326) <= not(layer4_outputs(599));
    layer5_outputs(2327) <= layer4_outputs(1564);
    layer5_outputs(2328) <= not((layer4_outputs(928)) and (layer4_outputs(1685)));
    layer5_outputs(2329) <= (layer4_outputs(2297)) xor (layer4_outputs(2553));
    layer5_outputs(2330) <= (layer4_outputs(1213)) and (layer4_outputs(1352));
    layer5_outputs(2331) <= layer4_outputs(98);
    layer5_outputs(2332) <= not((layer4_outputs(790)) and (layer4_outputs(1959)));
    layer5_outputs(2333) <= (layer4_outputs(778)) and not (layer4_outputs(784));
    layer5_outputs(2334) <= '0';
    layer5_outputs(2335) <= not(layer4_outputs(1330)) or (layer4_outputs(1732));
    layer5_outputs(2336) <= (layer4_outputs(187)) or (layer4_outputs(1315));
    layer5_outputs(2337) <= layer4_outputs(81);
    layer5_outputs(2338) <= layer4_outputs(1305);
    layer5_outputs(2339) <= not(layer4_outputs(2113)) or (layer4_outputs(631));
    layer5_outputs(2340) <= not(layer4_outputs(2175)) or (layer4_outputs(1669));
    layer5_outputs(2341) <= '0';
    layer5_outputs(2342) <= (layer4_outputs(978)) and not (layer4_outputs(2536));
    layer5_outputs(2343) <= not(layer4_outputs(1173));
    layer5_outputs(2344) <= (layer4_outputs(1944)) and (layer4_outputs(2539));
    layer5_outputs(2345) <= (layer4_outputs(1026)) or (layer4_outputs(2050));
    layer5_outputs(2346) <= not((layer4_outputs(1042)) xor (layer4_outputs(773)));
    layer5_outputs(2347) <= layer4_outputs(1658);
    layer5_outputs(2348) <= (layer4_outputs(154)) and (layer4_outputs(1736));
    layer5_outputs(2349) <= (layer4_outputs(1695)) and not (layer4_outputs(445));
    layer5_outputs(2350) <= layer4_outputs(1205);
    layer5_outputs(2351) <= (layer4_outputs(1310)) or (layer4_outputs(1938));
    layer5_outputs(2352) <= layer4_outputs(106);
    layer5_outputs(2353) <= '1';
    layer5_outputs(2354) <= not(layer4_outputs(2451));
    layer5_outputs(2355) <= not(layer4_outputs(1845)) or (layer4_outputs(1441));
    layer5_outputs(2356) <= '0';
    layer5_outputs(2357) <= layer4_outputs(1488);
    layer5_outputs(2358) <= not(layer4_outputs(756)) or (layer4_outputs(507));
    layer5_outputs(2359) <= layer4_outputs(1921);
    layer5_outputs(2360) <= not(layer4_outputs(2216));
    layer5_outputs(2361) <= (layer4_outputs(1695)) and not (layer4_outputs(995));
    layer5_outputs(2362) <= layer4_outputs(1227);
    layer5_outputs(2363) <= (layer4_outputs(299)) and not (layer4_outputs(1324));
    layer5_outputs(2364) <= layer4_outputs(2189);
    layer5_outputs(2365) <= not(layer4_outputs(1222));
    layer5_outputs(2366) <= not((layer4_outputs(450)) or (layer4_outputs(2547)));
    layer5_outputs(2367) <= not(layer4_outputs(1148));
    layer5_outputs(2368) <= '0';
    layer5_outputs(2369) <= (layer4_outputs(261)) and not (layer4_outputs(2304));
    layer5_outputs(2370) <= not(layer4_outputs(2452));
    layer5_outputs(2371) <= not(layer4_outputs(2195));
    layer5_outputs(2372) <= layer4_outputs(43);
    layer5_outputs(2373) <= not(layer4_outputs(1666));
    layer5_outputs(2374) <= (layer4_outputs(1113)) and (layer4_outputs(741));
    layer5_outputs(2375) <= '1';
    layer5_outputs(2376) <= (layer4_outputs(1363)) xor (layer4_outputs(265));
    layer5_outputs(2377) <= not(layer4_outputs(2346)) or (layer4_outputs(1152));
    layer5_outputs(2378) <= not(layer4_outputs(2043));
    layer5_outputs(2379) <= not(layer4_outputs(365)) or (layer4_outputs(1334));
    layer5_outputs(2380) <= (layer4_outputs(1384)) or (layer4_outputs(1272));
    layer5_outputs(2381) <= not((layer4_outputs(895)) and (layer4_outputs(2097)));
    layer5_outputs(2382) <= layer4_outputs(937);
    layer5_outputs(2383) <= (layer4_outputs(1918)) and (layer4_outputs(1890));
    layer5_outputs(2384) <= not(layer4_outputs(823));
    layer5_outputs(2385) <= layer4_outputs(21);
    layer5_outputs(2386) <= (layer4_outputs(1309)) and not (layer4_outputs(2258));
    layer5_outputs(2387) <= not(layer4_outputs(2368));
    layer5_outputs(2388) <= not((layer4_outputs(1405)) xor (layer4_outputs(2022)));
    layer5_outputs(2389) <= not((layer4_outputs(579)) and (layer4_outputs(885)));
    layer5_outputs(2390) <= (layer4_outputs(510)) and not (layer4_outputs(342));
    layer5_outputs(2391) <= (layer4_outputs(983)) and not (layer4_outputs(863));
    layer5_outputs(2392) <= not((layer4_outputs(54)) or (layer4_outputs(78)));
    layer5_outputs(2393) <= not(layer4_outputs(1712));
    layer5_outputs(2394) <= not(layer4_outputs(1308)) or (layer4_outputs(428));
    layer5_outputs(2395) <= (layer4_outputs(99)) or (layer4_outputs(436));
    layer5_outputs(2396) <= (layer4_outputs(2351)) and not (layer4_outputs(1184));
    layer5_outputs(2397) <= layer4_outputs(1109);
    layer5_outputs(2398) <= (layer4_outputs(644)) or (layer4_outputs(1993));
    layer5_outputs(2399) <= (layer4_outputs(530)) or (layer4_outputs(828));
    layer5_outputs(2400) <= layer4_outputs(1704);
    layer5_outputs(2401) <= (layer4_outputs(596)) and (layer4_outputs(1074));
    layer5_outputs(2402) <= not(layer4_outputs(2057));
    layer5_outputs(2403) <= (layer4_outputs(411)) and not (layer4_outputs(1154));
    layer5_outputs(2404) <= not(layer4_outputs(48));
    layer5_outputs(2405) <= not(layer4_outputs(695));
    layer5_outputs(2406) <= not(layer4_outputs(795));
    layer5_outputs(2407) <= not((layer4_outputs(2077)) and (layer4_outputs(408)));
    layer5_outputs(2408) <= (layer4_outputs(1889)) or (layer4_outputs(1153));
    layer5_outputs(2409) <= not(layer4_outputs(13));
    layer5_outputs(2410) <= not(layer4_outputs(746));
    layer5_outputs(2411) <= (layer4_outputs(413)) and not (layer4_outputs(1362));
    layer5_outputs(2412) <= not(layer4_outputs(1289)) or (layer4_outputs(1293));
    layer5_outputs(2413) <= layer4_outputs(874);
    layer5_outputs(2414) <= layer4_outputs(419);
    layer5_outputs(2415) <= not(layer4_outputs(69));
    layer5_outputs(2416) <= layer4_outputs(2000);
    layer5_outputs(2417) <= not((layer4_outputs(1426)) xor (layer4_outputs(2542)));
    layer5_outputs(2418) <= (layer4_outputs(75)) and (layer4_outputs(1460));
    layer5_outputs(2419) <= (layer4_outputs(989)) and not (layer4_outputs(1972));
    layer5_outputs(2420) <= (layer4_outputs(1494)) xor (layer4_outputs(1249));
    layer5_outputs(2421) <= (layer4_outputs(359)) or (layer4_outputs(1263));
    layer5_outputs(2422) <= not(layer4_outputs(141));
    layer5_outputs(2423) <= (layer4_outputs(328)) or (layer4_outputs(2241));
    layer5_outputs(2424) <= '0';
    layer5_outputs(2425) <= layer4_outputs(2143);
    layer5_outputs(2426) <= not(layer4_outputs(1864));
    layer5_outputs(2427) <= not((layer4_outputs(209)) and (layer4_outputs(2078)));
    layer5_outputs(2428) <= (layer4_outputs(172)) xor (layer4_outputs(1227));
    layer5_outputs(2429) <= (layer4_outputs(2198)) and (layer4_outputs(1552));
    layer5_outputs(2430) <= not(layer4_outputs(1727));
    layer5_outputs(2431) <= not(layer4_outputs(2453)) or (layer4_outputs(295));
    layer5_outputs(2432) <= (layer4_outputs(2165)) and (layer4_outputs(783));
    layer5_outputs(2433) <= (layer4_outputs(2187)) or (layer4_outputs(1758));
    layer5_outputs(2434) <= (layer4_outputs(1697)) and not (layer4_outputs(235));
    layer5_outputs(2435) <= not(layer4_outputs(188));
    layer5_outputs(2436) <= '1';
    layer5_outputs(2437) <= not(layer4_outputs(1906));
    layer5_outputs(2438) <= '1';
    layer5_outputs(2439) <= layer4_outputs(444);
    layer5_outputs(2440) <= (layer4_outputs(1202)) xor (layer4_outputs(11));
    layer5_outputs(2441) <= layer4_outputs(387);
    layer5_outputs(2442) <= not(layer4_outputs(1135)) or (layer4_outputs(1052));
    layer5_outputs(2443) <= not((layer4_outputs(132)) or (layer4_outputs(2177)));
    layer5_outputs(2444) <= not(layer4_outputs(873));
    layer5_outputs(2445) <= '1';
    layer5_outputs(2446) <= not(layer4_outputs(348)) or (layer4_outputs(594));
    layer5_outputs(2447) <= (layer4_outputs(102)) and (layer4_outputs(766));
    layer5_outputs(2448) <= not(layer4_outputs(1348));
    layer5_outputs(2449) <= not(layer4_outputs(626));
    layer5_outputs(2450) <= not(layer4_outputs(1480));
    layer5_outputs(2451) <= layer4_outputs(2301);
    layer5_outputs(2452) <= (layer4_outputs(2323)) and not (layer4_outputs(2062));
    layer5_outputs(2453) <= (layer4_outputs(1620)) and (layer4_outputs(677));
    layer5_outputs(2454) <= layer4_outputs(815);
    layer5_outputs(2455) <= not((layer4_outputs(1107)) or (layer4_outputs(387)));
    layer5_outputs(2456) <= not((layer4_outputs(1916)) or (layer4_outputs(1094)));
    layer5_outputs(2457) <= (layer4_outputs(2382)) and not (layer4_outputs(1986));
    layer5_outputs(2458) <= not((layer4_outputs(1308)) or (layer4_outputs(1731)));
    layer5_outputs(2459) <= (layer4_outputs(2428)) and (layer4_outputs(1055));
    layer5_outputs(2460) <= not((layer4_outputs(1208)) or (layer4_outputs(1247)));
    layer5_outputs(2461) <= not(layer4_outputs(337));
    layer5_outputs(2462) <= not((layer4_outputs(2050)) or (layer4_outputs(1644)));
    layer5_outputs(2463) <= layer4_outputs(2528);
    layer5_outputs(2464) <= (layer4_outputs(2254)) or (layer4_outputs(2303));
    layer5_outputs(2465) <= (layer4_outputs(756)) xor (layer4_outputs(2033));
    layer5_outputs(2466) <= (layer4_outputs(2203)) and (layer4_outputs(1507));
    layer5_outputs(2467) <= layer4_outputs(1099);
    layer5_outputs(2468) <= not(layer4_outputs(1328)) or (layer4_outputs(248));
    layer5_outputs(2469) <= layer4_outputs(1471);
    layer5_outputs(2470) <= (layer4_outputs(2131)) xor (layer4_outputs(2492));
    layer5_outputs(2471) <= (layer4_outputs(1702)) and not (layer4_outputs(905));
    layer5_outputs(2472) <= (layer4_outputs(1815)) and not (layer4_outputs(1647));
    layer5_outputs(2473) <= layer4_outputs(1790);
    layer5_outputs(2474) <= (layer4_outputs(61)) or (layer4_outputs(1331));
    layer5_outputs(2475) <= not(layer4_outputs(888)) or (layer4_outputs(748));
    layer5_outputs(2476) <= not(layer4_outputs(2512)) or (layer4_outputs(131));
    layer5_outputs(2477) <= not(layer4_outputs(339));
    layer5_outputs(2478) <= not(layer4_outputs(1720)) or (layer4_outputs(2160));
    layer5_outputs(2479) <= not(layer4_outputs(1262));
    layer5_outputs(2480) <= layer4_outputs(1486);
    layer5_outputs(2481) <= not(layer4_outputs(1609)) or (layer4_outputs(775));
    layer5_outputs(2482) <= (layer4_outputs(2162)) and not (layer4_outputs(1639));
    layer5_outputs(2483) <= (layer4_outputs(1408)) or (layer4_outputs(759));
    layer5_outputs(2484) <= not(layer4_outputs(545)) or (layer4_outputs(1630));
    layer5_outputs(2485) <= layer4_outputs(118);
    layer5_outputs(2486) <= '0';
    layer5_outputs(2487) <= not((layer4_outputs(1101)) xor (layer4_outputs(1606)));
    layer5_outputs(2488) <= (layer4_outputs(1453)) and not (layer4_outputs(1081));
    layer5_outputs(2489) <= not(layer4_outputs(400)) or (layer4_outputs(251));
    layer5_outputs(2490) <= layer4_outputs(2161);
    layer5_outputs(2491) <= not((layer4_outputs(1181)) or (layer4_outputs(771)));
    layer5_outputs(2492) <= layer4_outputs(2414);
    layer5_outputs(2493) <= (layer4_outputs(866)) xor (layer4_outputs(424));
    layer5_outputs(2494) <= '0';
    layer5_outputs(2495) <= layer4_outputs(2026);
    layer5_outputs(2496) <= layer4_outputs(1479);
    layer5_outputs(2497) <= not(layer4_outputs(1751));
    layer5_outputs(2498) <= (layer4_outputs(1869)) and not (layer4_outputs(1570));
    layer5_outputs(2499) <= layer4_outputs(1544);
    layer5_outputs(2500) <= not((layer4_outputs(120)) and (layer4_outputs(2526)));
    layer5_outputs(2501) <= layer4_outputs(1953);
    layer5_outputs(2502) <= not(layer4_outputs(997)) or (layer4_outputs(1485));
    layer5_outputs(2503) <= not(layer4_outputs(1763));
    layer5_outputs(2504) <= layer4_outputs(1666);
    layer5_outputs(2505) <= not(layer4_outputs(315));
    layer5_outputs(2506) <= '0';
    layer5_outputs(2507) <= '0';
    layer5_outputs(2508) <= '0';
    layer5_outputs(2509) <= not((layer4_outputs(2166)) and (layer4_outputs(1036)));
    layer5_outputs(2510) <= not(layer4_outputs(2218));
    layer5_outputs(2511) <= not((layer4_outputs(2375)) xor (layer4_outputs(1165)));
    layer5_outputs(2512) <= layer4_outputs(380);
    layer5_outputs(2513) <= layer4_outputs(2029);
    layer5_outputs(2514) <= not((layer4_outputs(485)) and (layer4_outputs(2107)));
    layer5_outputs(2515) <= not(layer4_outputs(993)) or (layer4_outputs(1171));
    layer5_outputs(2516) <= layer4_outputs(258);
    layer5_outputs(2517) <= layer4_outputs(619);
    layer5_outputs(2518) <= not(layer4_outputs(2248));
    layer5_outputs(2519) <= layer4_outputs(39);
    layer5_outputs(2520) <= layer4_outputs(913);
    layer5_outputs(2521) <= '1';
    layer5_outputs(2522) <= (layer4_outputs(1144)) and not (layer4_outputs(2267));
    layer5_outputs(2523) <= layer4_outputs(1474);
    layer5_outputs(2524) <= (layer4_outputs(752)) or (layer4_outputs(1120));
    layer5_outputs(2525) <= (layer4_outputs(2183)) xor (layer4_outputs(456));
    layer5_outputs(2526) <= layer4_outputs(1426);
    layer5_outputs(2527) <= layer4_outputs(1295);
    layer5_outputs(2528) <= layer4_outputs(630);
    layer5_outputs(2529) <= (layer4_outputs(1104)) xor (layer4_outputs(1279));
    layer5_outputs(2530) <= (layer4_outputs(2027)) and not (layer4_outputs(2339));
    layer5_outputs(2531) <= not(layer4_outputs(2066));
    layer5_outputs(2532) <= not(layer4_outputs(1846)) or (layer4_outputs(2018));
    layer5_outputs(2533) <= (layer4_outputs(213)) and (layer4_outputs(349));
    layer5_outputs(2534) <= not(layer4_outputs(849));
    layer5_outputs(2535) <= not(layer4_outputs(1800));
    layer5_outputs(2536) <= not(layer4_outputs(100)) or (layer4_outputs(2551));
    layer5_outputs(2537) <= not((layer4_outputs(1770)) or (layer4_outputs(876)));
    layer5_outputs(2538) <= not(layer4_outputs(1080));
    layer5_outputs(2539) <= layer4_outputs(1472);
    layer5_outputs(2540) <= (layer4_outputs(1253)) and not (layer4_outputs(2461));
    layer5_outputs(2541) <= not((layer4_outputs(2096)) or (layer4_outputs(2246)));
    layer5_outputs(2542) <= (layer4_outputs(506)) and not (layer4_outputs(1920));
    layer5_outputs(2543) <= not(layer4_outputs(1597)) or (layer4_outputs(149));
    layer5_outputs(2544) <= layer4_outputs(1662);
    layer5_outputs(2545) <= layer4_outputs(1995);
    layer5_outputs(2546) <= (layer4_outputs(1677)) and not (layer4_outputs(1950));
    layer5_outputs(2547) <= (layer4_outputs(2069)) and not (layer4_outputs(1671));
    layer5_outputs(2548) <= not((layer4_outputs(2329)) or (layer4_outputs(1904)));
    layer5_outputs(2549) <= not(layer4_outputs(81)) or (layer4_outputs(2503));
    layer5_outputs(2550) <= (layer4_outputs(2063)) and not (layer4_outputs(909));
    layer5_outputs(2551) <= not(layer4_outputs(2225)) or (layer4_outputs(1114));
    layer5_outputs(2552) <= layer4_outputs(2385);
    layer5_outputs(2553) <= (layer4_outputs(1914)) and (layer4_outputs(1693));
    layer5_outputs(2554) <= not((layer4_outputs(178)) and (layer4_outputs(1655)));
    layer5_outputs(2555) <= not(layer4_outputs(2394));
    layer5_outputs(2556) <= (layer4_outputs(1603)) xor (layer4_outputs(619));
    layer5_outputs(2557) <= not(layer4_outputs(1351));
    layer5_outputs(2558) <= (layer4_outputs(2053)) or (layer4_outputs(2048));
    layer5_outputs(2559) <= not(layer4_outputs(415)) or (layer4_outputs(1738));
    layer6_outputs(0) <= layer5_outputs(1842);
    layer6_outputs(1) <= not((layer5_outputs(1511)) xor (layer5_outputs(1068)));
    layer6_outputs(2) <= not(layer5_outputs(2555)) or (layer5_outputs(1162));
    layer6_outputs(3) <= not(layer5_outputs(1671));
    layer6_outputs(4) <= not((layer5_outputs(2495)) xor (layer5_outputs(282)));
    layer6_outputs(5) <= (layer5_outputs(1955)) and not (layer5_outputs(2282));
    layer6_outputs(6) <= layer5_outputs(870);
    layer6_outputs(7) <= layer5_outputs(556);
    layer6_outputs(8) <= layer5_outputs(25);
    layer6_outputs(9) <= layer5_outputs(233);
    layer6_outputs(10) <= not(layer5_outputs(2222)) or (layer5_outputs(2343));
    layer6_outputs(11) <= not(layer5_outputs(1020));
    layer6_outputs(12) <= layer5_outputs(2028);
    layer6_outputs(13) <= (layer5_outputs(692)) and not (layer5_outputs(1842));
    layer6_outputs(14) <= not((layer5_outputs(973)) and (layer5_outputs(372)));
    layer6_outputs(15) <= not(layer5_outputs(2046));
    layer6_outputs(16) <= layer5_outputs(1187);
    layer6_outputs(17) <= not(layer5_outputs(558)) or (layer5_outputs(519));
    layer6_outputs(18) <= (layer5_outputs(801)) xor (layer5_outputs(517));
    layer6_outputs(19) <= not(layer5_outputs(2195));
    layer6_outputs(20) <= not(layer5_outputs(1503));
    layer6_outputs(21) <= (layer5_outputs(531)) xor (layer5_outputs(1867));
    layer6_outputs(22) <= (layer5_outputs(928)) xor (layer5_outputs(696));
    layer6_outputs(23) <= layer5_outputs(1805);
    layer6_outputs(24) <= not(layer5_outputs(797)) or (layer5_outputs(2211));
    layer6_outputs(25) <= layer5_outputs(2503);
    layer6_outputs(26) <= (layer5_outputs(1201)) and not (layer5_outputs(1985));
    layer6_outputs(27) <= (layer5_outputs(1224)) or (layer5_outputs(1598));
    layer6_outputs(28) <= (layer5_outputs(160)) or (layer5_outputs(1930));
    layer6_outputs(29) <= layer5_outputs(755);
    layer6_outputs(30) <= (layer5_outputs(1311)) xor (layer5_outputs(1668));
    layer6_outputs(31) <= not(layer5_outputs(2178));
    layer6_outputs(32) <= not((layer5_outputs(979)) and (layer5_outputs(1045)));
    layer6_outputs(33) <= not(layer5_outputs(1124)) or (layer5_outputs(856));
    layer6_outputs(34) <= layer5_outputs(1112);
    layer6_outputs(35) <= layer5_outputs(1563);
    layer6_outputs(36) <= not(layer5_outputs(802));
    layer6_outputs(37) <= not((layer5_outputs(682)) and (layer5_outputs(1551)));
    layer6_outputs(38) <= '0';
    layer6_outputs(39) <= layer5_outputs(1527);
    layer6_outputs(40) <= (layer5_outputs(2248)) and (layer5_outputs(1592));
    layer6_outputs(41) <= not(layer5_outputs(553));
    layer6_outputs(42) <= (layer5_outputs(44)) and (layer5_outputs(793));
    layer6_outputs(43) <= layer5_outputs(2253);
    layer6_outputs(44) <= not((layer5_outputs(474)) or (layer5_outputs(2090)));
    layer6_outputs(45) <= (layer5_outputs(498)) and (layer5_outputs(2071));
    layer6_outputs(46) <= not(layer5_outputs(2415)) or (layer5_outputs(820));
    layer6_outputs(47) <= not(layer5_outputs(2284));
    layer6_outputs(48) <= (layer5_outputs(117)) and not (layer5_outputs(1682));
    layer6_outputs(49) <= layer5_outputs(2236);
    layer6_outputs(50) <= not(layer5_outputs(1701)) or (layer5_outputs(1202));
    layer6_outputs(51) <= not(layer5_outputs(1354)) or (layer5_outputs(2058));
    layer6_outputs(52) <= layer5_outputs(1738);
    layer6_outputs(53) <= (layer5_outputs(770)) xor (layer5_outputs(2230));
    layer6_outputs(54) <= layer5_outputs(1698);
    layer6_outputs(55) <= layer5_outputs(2113);
    layer6_outputs(56) <= not(layer5_outputs(2239));
    layer6_outputs(57) <= layer5_outputs(46);
    layer6_outputs(58) <= not(layer5_outputs(731));
    layer6_outputs(59) <= not(layer5_outputs(2213)) or (layer5_outputs(1173));
    layer6_outputs(60) <= layer5_outputs(1642);
    layer6_outputs(61) <= layer5_outputs(2360);
    layer6_outputs(62) <= layer5_outputs(1508);
    layer6_outputs(63) <= (layer5_outputs(641)) and not (layer5_outputs(1972));
    layer6_outputs(64) <= (layer5_outputs(1413)) xor (layer5_outputs(557));
    layer6_outputs(65) <= not(layer5_outputs(2248));
    layer6_outputs(66) <= layer5_outputs(1552);
    layer6_outputs(67) <= not((layer5_outputs(2364)) xor (layer5_outputs(189)));
    layer6_outputs(68) <= not(layer5_outputs(1433));
    layer6_outputs(69) <= layer5_outputs(402);
    layer6_outputs(70) <= '0';
    layer6_outputs(71) <= not(layer5_outputs(367)) or (layer5_outputs(1992));
    layer6_outputs(72) <= not((layer5_outputs(945)) xor (layer5_outputs(812)));
    layer6_outputs(73) <= not(layer5_outputs(115));
    layer6_outputs(74) <= not((layer5_outputs(1724)) xor (layer5_outputs(2129)));
    layer6_outputs(75) <= not(layer5_outputs(2025)) or (layer5_outputs(227));
    layer6_outputs(76) <= (layer5_outputs(2477)) and (layer5_outputs(1515));
    layer6_outputs(77) <= (layer5_outputs(18)) and not (layer5_outputs(519));
    layer6_outputs(78) <= not(layer5_outputs(1648)) or (layer5_outputs(1439));
    layer6_outputs(79) <= not(layer5_outputs(2254));
    layer6_outputs(80) <= not((layer5_outputs(1807)) or (layer5_outputs(644)));
    layer6_outputs(81) <= layer5_outputs(1179);
    layer6_outputs(82) <= (layer5_outputs(29)) and (layer5_outputs(1464));
    layer6_outputs(83) <= layer5_outputs(329);
    layer6_outputs(84) <= not(layer5_outputs(1611));
    layer6_outputs(85) <= not(layer5_outputs(1356)) or (layer5_outputs(1401));
    layer6_outputs(86) <= not(layer5_outputs(1421)) or (layer5_outputs(1824));
    layer6_outputs(87) <= layer5_outputs(1590);
    layer6_outputs(88) <= layer5_outputs(1464);
    layer6_outputs(89) <= not((layer5_outputs(1348)) or (layer5_outputs(1200)));
    layer6_outputs(90) <= not(layer5_outputs(1507));
    layer6_outputs(91) <= layer5_outputs(2383);
    layer6_outputs(92) <= not(layer5_outputs(652));
    layer6_outputs(93) <= not((layer5_outputs(704)) and (layer5_outputs(726)));
    layer6_outputs(94) <= (layer5_outputs(880)) xor (layer5_outputs(385));
    layer6_outputs(95) <= not((layer5_outputs(1435)) or (layer5_outputs(258)));
    layer6_outputs(96) <= not(layer5_outputs(1266));
    layer6_outputs(97) <= not(layer5_outputs(2075));
    layer6_outputs(98) <= not((layer5_outputs(1028)) xor (layer5_outputs(446)));
    layer6_outputs(99) <= layer5_outputs(889);
    layer6_outputs(100) <= layer5_outputs(2151);
    layer6_outputs(101) <= (layer5_outputs(1569)) and not (layer5_outputs(1342));
    layer6_outputs(102) <= layer5_outputs(752);
    layer6_outputs(103) <= not(layer5_outputs(130)) or (layer5_outputs(1289));
    layer6_outputs(104) <= not(layer5_outputs(839));
    layer6_outputs(105) <= layer5_outputs(1617);
    layer6_outputs(106) <= layer5_outputs(1202);
    layer6_outputs(107) <= (layer5_outputs(449)) and not (layer5_outputs(2465));
    layer6_outputs(108) <= not(layer5_outputs(1449));
    layer6_outputs(109) <= layer5_outputs(836);
    layer6_outputs(110) <= not(layer5_outputs(1801));
    layer6_outputs(111) <= (layer5_outputs(187)) and (layer5_outputs(1859));
    layer6_outputs(112) <= layer5_outputs(1906);
    layer6_outputs(113) <= (layer5_outputs(548)) xor (layer5_outputs(1772));
    layer6_outputs(114) <= not((layer5_outputs(2013)) and (layer5_outputs(992)));
    layer6_outputs(115) <= layer5_outputs(2357);
    layer6_outputs(116) <= not(layer5_outputs(2205));
    layer6_outputs(117) <= not((layer5_outputs(1897)) xor (layer5_outputs(1836)));
    layer6_outputs(118) <= not(layer5_outputs(38));
    layer6_outputs(119) <= '1';
    layer6_outputs(120) <= (layer5_outputs(1935)) xor (layer5_outputs(1033));
    layer6_outputs(121) <= (layer5_outputs(1292)) and not (layer5_outputs(144));
    layer6_outputs(122) <= not((layer5_outputs(1492)) or (layer5_outputs(555)));
    layer6_outputs(123) <= not((layer5_outputs(439)) or (layer5_outputs(1716)));
    layer6_outputs(124) <= (layer5_outputs(382)) and not (layer5_outputs(1132));
    layer6_outputs(125) <= not(layer5_outputs(699)) or (layer5_outputs(1210));
    layer6_outputs(126) <= not(layer5_outputs(1408)) or (layer5_outputs(2421));
    layer6_outputs(127) <= not(layer5_outputs(272));
    layer6_outputs(128) <= (layer5_outputs(2509)) and (layer5_outputs(1142));
    layer6_outputs(129) <= not(layer5_outputs(2327));
    layer6_outputs(130) <= not(layer5_outputs(1698));
    layer6_outputs(131) <= not(layer5_outputs(981));
    layer6_outputs(132) <= layer5_outputs(47);
    layer6_outputs(133) <= not(layer5_outputs(1785));
    layer6_outputs(134) <= layer5_outputs(1183);
    layer6_outputs(135) <= not((layer5_outputs(1944)) or (layer5_outputs(1487)));
    layer6_outputs(136) <= (layer5_outputs(112)) or (layer5_outputs(1954));
    layer6_outputs(137) <= not(layer5_outputs(353));
    layer6_outputs(138) <= layer5_outputs(1648);
    layer6_outputs(139) <= (layer5_outputs(771)) or (layer5_outputs(376));
    layer6_outputs(140) <= (layer5_outputs(2377)) xor (layer5_outputs(529));
    layer6_outputs(141) <= not(layer5_outputs(1929));
    layer6_outputs(142) <= not(layer5_outputs(1230));
    layer6_outputs(143) <= not(layer5_outputs(1408));
    layer6_outputs(144) <= layer5_outputs(296);
    layer6_outputs(145) <= not(layer5_outputs(2077)) or (layer5_outputs(1298));
    layer6_outputs(146) <= not((layer5_outputs(1989)) xor (layer5_outputs(2550)));
    layer6_outputs(147) <= not((layer5_outputs(1157)) and (layer5_outputs(1930)));
    layer6_outputs(148) <= layer5_outputs(1569);
    layer6_outputs(149) <= (layer5_outputs(2370)) xor (layer5_outputs(1091));
    layer6_outputs(150) <= layer5_outputs(331);
    layer6_outputs(151) <= layer5_outputs(8);
    layer6_outputs(152) <= not(layer5_outputs(1783));
    layer6_outputs(153) <= (layer5_outputs(274)) xor (layer5_outputs(243));
    layer6_outputs(154) <= not((layer5_outputs(1896)) xor (layer5_outputs(181)));
    layer6_outputs(155) <= not(layer5_outputs(901));
    layer6_outputs(156) <= not((layer5_outputs(2348)) xor (layer5_outputs(1733)));
    layer6_outputs(157) <= (layer5_outputs(2234)) xor (layer5_outputs(2009));
    layer6_outputs(158) <= not(layer5_outputs(96));
    layer6_outputs(159) <= not(layer5_outputs(1557));
    layer6_outputs(160) <= not((layer5_outputs(1015)) and (layer5_outputs(2060)));
    layer6_outputs(161) <= not(layer5_outputs(1415));
    layer6_outputs(162) <= (layer5_outputs(2188)) xor (layer5_outputs(1038));
    layer6_outputs(163) <= (layer5_outputs(1960)) xor (layer5_outputs(731));
    layer6_outputs(164) <= (layer5_outputs(1786)) and (layer5_outputs(545));
    layer6_outputs(165) <= layer5_outputs(409);
    layer6_outputs(166) <= not((layer5_outputs(1463)) xor (layer5_outputs(2128)));
    layer6_outputs(167) <= not((layer5_outputs(2255)) xor (layer5_outputs(401)));
    layer6_outputs(168) <= layer5_outputs(1380);
    layer6_outputs(169) <= not(layer5_outputs(243));
    layer6_outputs(170) <= not((layer5_outputs(1659)) and (layer5_outputs(2000)));
    layer6_outputs(171) <= not((layer5_outputs(1394)) and (layer5_outputs(2452)));
    layer6_outputs(172) <= (layer5_outputs(596)) and (layer5_outputs(1966));
    layer6_outputs(173) <= layer5_outputs(748);
    layer6_outputs(174) <= layer5_outputs(466);
    layer6_outputs(175) <= (layer5_outputs(1963)) and not (layer5_outputs(708));
    layer6_outputs(176) <= not((layer5_outputs(2524)) xor (layer5_outputs(511)));
    layer6_outputs(177) <= (layer5_outputs(476)) and (layer5_outputs(567));
    layer6_outputs(178) <= layer5_outputs(1597);
    layer6_outputs(179) <= not((layer5_outputs(140)) xor (layer5_outputs(533)));
    layer6_outputs(180) <= (layer5_outputs(840)) xor (layer5_outputs(2449));
    layer6_outputs(181) <= not(layer5_outputs(859));
    layer6_outputs(182) <= layer5_outputs(586);
    layer6_outputs(183) <= (layer5_outputs(886)) or (layer5_outputs(694));
    layer6_outputs(184) <= layer5_outputs(101);
    layer6_outputs(185) <= not((layer5_outputs(1011)) xor (layer5_outputs(877)));
    layer6_outputs(186) <= (layer5_outputs(1888)) and not (layer5_outputs(831));
    layer6_outputs(187) <= not(layer5_outputs(1706)) or (layer5_outputs(2035));
    layer6_outputs(188) <= (layer5_outputs(297)) xor (layer5_outputs(382));
    layer6_outputs(189) <= (layer5_outputs(2201)) or (layer5_outputs(43));
    layer6_outputs(190) <= not((layer5_outputs(636)) or (layer5_outputs(1461)));
    layer6_outputs(191) <= (layer5_outputs(950)) and (layer5_outputs(180));
    layer6_outputs(192) <= layer5_outputs(2340);
    layer6_outputs(193) <= not((layer5_outputs(2370)) and (layer5_outputs(158)));
    layer6_outputs(194) <= not(layer5_outputs(2069));
    layer6_outputs(195) <= (layer5_outputs(1593)) or (layer5_outputs(1732));
    layer6_outputs(196) <= layer5_outputs(2496);
    layer6_outputs(197) <= layer5_outputs(2448);
    layer6_outputs(198) <= not(layer5_outputs(2186));
    layer6_outputs(199) <= not(layer5_outputs(487));
    layer6_outputs(200) <= (layer5_outputs(341)) and not (layer5_outputs(380));
    layer6_outputs(201) <= not(layer5_outputs(1414));
    layer6_outputs(202) <= layer5_outputs(1708);
    layer6_outputs(203) <= layer5_outputs(1411);
    layer6_outputs(204) <= (layer5_outputs(47)) or (layer5_outputs(158));
    layer6_outputs(205) <= not(layer5_outputs(1615)) or (layer5_outputs(1265));
    layer6_outputs(206) <= layer5_outputs(1563);
    layer6_outputs(207) <= not(layer5_outputs(1748));
    layer6_outputs(208) <= not((layer5_outputs(874)) or (layer5_outputs(504)));
    layer6_outputs(209) <= not(layer5_outputs(452));
    layer6_outputs(210) <= layer5_outputs(824);
    layer6_outputs(211) <= not((layer5_outputs(1757)) xor (layer5_outputs(520)));
    layer6_outputs(212) <= not((layer5_outputs(398)) and (layer5_outputs(1167)));
    layer6_outputs(213) <= not(layer5_outputs(768));
    layer6_outputs(214) <= layer5_outputs(898);
    layer6_outputs(215) <= layer5_outputs(2216);
    layer6_outputs(216) <= layer5_outputs(2138);
    layer6_outputs(217) <= not(layer5_outputs(1333));
    layer6_outputs(218) <= layer5_outputs(644);
    layer6_outputs(219) <= not((layer5_outputs(138)) or (layer5_outputs(1415)));
    layer6_outputs(220) <= not(layer5_outputs(388)) or (layer5_outputs(2053));
    layer6_outputs(221) <= not(layer5_outputs(724));
    layer6_outputs(222) <= (layer5_outputs(1196)) and (layer5_outputs(1730));
    layer6_outputs(223) <= not((layer5_outputs(2468)) or (layer5_outputs(1844)));
    layer6_outputs(224) <= (layer5_outputs(913)) and not (layer5_outputs(1641));
    layer6_outputs(225) <= not(layer5_outputs(414));
    layer6_outputs(226) <= not((layer5_outputs(122)) xor (layer5_outputs(2004)));
    layer6_outputs(227) <= not((layer5_outputs(1154)) xor (layer5_outputs(443)));
    layer6_outputs(228) <= not((layer5_outputs(525)) and (layer5_outputs(1670)));
    layer6_outputs(229) <= layer5_outputs(1056);
    layer6_outputs(230) <= not((layer5_outputs(1875)) or (layer5_outputs(2462)));
    layer6_outputs(231) <= layer5_outputs(1018);
    layer6_outputs(232) <= not(layer5_outputs(2054));
    layer6_outputs(233) <= layer5_outputs(1281);
    layer6_outputs(234) <= layer5_outputs(1392);
    layer6_outputs(235) <= (layer5_outputs(632)) or (layer5_outputs(211));
    layer6_outputs(236) <= layer5_outputs(540);
    layer6_outputs(237) <= (layer5_outputs(2475)) xor (layer5_outputs(2274));
    layer6_outputs(238) <= not(layer5_outputs(575));
    layer6_outputs(239) <= not(layer5_outputs(2069));
    layer6_outputs(240) <= layer5_outputs(2398);
    layer6_outputs(241) <= layer5_outputs(855);
    layer6_outputs(242) <= not(layer5_outputs(245)) or (layer5_outputs(1852));
    layer6_outputs(243) <= not(layer5_outputs(2109));
    layer6_outputs(244) <= layer5_outputs(24);
    layer6_outputs(245) <= not((layer5_outputs(1554)) xor (layer5_outputs(517)));
    layer6_outputs(246) <= not(layer5_outputs(1974));
    layer6_outputs(247) <= not((layer5_outputs(439)) or (layer5_outputs(2542)));
    layer6_outputs(248) <= not(layer5_outputs(1453));
    layer6_outputs(249) <= not(layer5_outputs(1051));
    layer6_outputs(250) <= not((layer5_outputs(1693)) or (layer5_outputs(658)));
    layer6_outputs(251) <= (layer5_outputs(1231)) or (layer5_outputs(1689));
    layer6_outputs(252) <= not((layer5_outputs(1104)) and (layer5_outputs(2408)));
    layer6_outputs(253) <= (layer5_outputs(190)) or (layer5_outputs(16));
    layer6_outputs(254) <= (layer5_outputs(1396)) xor (layer5_outputs(898));
    layer6_outputs(255) <= (layer5_outputs(2367)) xor (layer5_outputs(1719));
    layer6_outputs(256) <= (layer5_outputs(1489)) and not (layer5_outputs(2504));
    layer6_outputs(257) <= (layer5_outputs(1886)) or (layer5_outputs(1726));
    layer6_outputs(258) <= (layer5_outputs(2479)) xor (layer5_outputs(1402));
    layer6_outputs(259) <= not(layer5_outputs(1494));
    layer6_outputs(260) <= layer5_outputs(360);
    layer6_outputs(261) <= (layer5_outputs(2290)) and (layer5_outputs(63));
    layer6_outputs(262) <= '0';
    layer6_outputs(263) <= not(layer5_outputs(2089));
    layer6_outputs(264) <= not(layer5_outputs(501)) or (layer5_outputs(841));
    layer6_outputs(265) <= not((layer5_outputs(2114)) xor (layer5_outputs(225)));
    layer6_outputs(266) <= layer5_outputs(591);
    layer6_outputs(267) <= layer5_outputs(2315);
    layer6_outputs(268) <= layer5_outputs(565);
    layer6_outputs(269) <= not(layer5_outputs(946));
    layer6_outputs(270) <= not(layer5_outputs(1999));
    layer6_outputs(271) <= not(layer5_outputs(2326)) or (layer5_outputs(2292));
    layer6_outputs(272) <= not(layer5_outputs(550));
    layer6_outputs(273) <= not(layer5_outputs(1208));
    layer6_outputs(274) <= not(layer5_outputs(160));
    layer6_outputs(275) <= not(layer5_outputs(1826));
    layer6_outputs(276) <= not(layer5_outputs(2147));
    layer6_outputs(277) <= layer5_outputs(2297);
    layer6_outputs(278) <= layer5_outputs(512);
    layer6_outputs(279) <= (layer5_outputs(1322)) or (layer5_outputs(779));
    layer6_outputs(280) <= layer5_outputs(1558);
    layer6_outputs(281) <= not(layer5_outputs(709));
    layer6_outputs(282) <= not(layer5_outputs(989));
    layer6_outputs(283) <= (layer5_outputs(812)) xor (layer5_outputs(1420));
    layer6_outputs(284) <= layer5_outputs(562);
    layer6_outputs(285) <= not(layer5_outputs(2534));
    layer6_outputs(286) <= layer5_outputs(1642);
    layer6_outputs(287) <= not(layer5_outputs(1369));
    layer6_outputs(288) <= not(layer5_outputs(726)) or (layer5_outputs(1779));
    layer6_outputs(289) <= layer5_outputs(70);
    layer6_outputs(290) <= layer5_outputs(1636);
    layer6_outputs(291) <= not(layer5_outputs(48));
    layer6_outputs(292) <= not((layer5_outputs(1696)) xor (layer5_outputs(1232)));
    layer6_outputs(293) <= (layer5_outputs(1427)) and not (layer5_outputs(268));
    layer6_outputs(294) <= layer5_outputs(970);
    layer6_outputs(295) <= not(layer5_outputs(2309));
    layer6_outputs(296) <= (layer5_outputs(1827)) xor (layer5_outputs(723));
    layer6_outputs(297) <= not(layer5_outputs(1876));
    layer6_outputs(298) <= (layer5_outputs(753)) and (layer5_outputs(1250));
    layer6_outputs(299) <= not(layer5_outputs(677));
    layer6_outputs(300) <= not(layer5_outputs(2331)) or (layer5_outputs(1970));
    layer6_outputs(301) <= layer5_outputs(225);
    layer6_outputs(302) <= not(layer5_outputs(1949));
    layer6_outputs(303) <= (layer5_outputs(1106)) and not (layer5_outputs(1715));
    layer6_outputs(304) <= (layer5_outputs(696)) and (layer5_outputs(2345));
    layer6_outputs(305) <= not(layer5_outputs(2093));
    layer6_outputs(306) <= (layer5_outputs(294)) and not (layer5_outputs(497));
    layer6_outputs(307) <= not((layer5_outputs(969)) or (layer5_outputs(1270)));
    layer6_outputs(308) <= not(layer5_outputs(581));
    layer6_outputs(309) <= layer5_outputs(1908);
    layer6_outputs(310) <= not((layer5_outputs(121)) xor (layer5_outputs(356)));
    layer6_outputs(311) <= (layer5_outputs(1246)) or (layer5_outputs(1554));
    layer6_outputs(312) <= layer5_outputs(2392);
    layer6_outputs(313) <= not(layer5_outputs(1950));
    layer6_outputs(314) <= (layer5_outputs(1575)) and not (layer5_outputs(1407));
    layer6_outputs(315) <= '1';
    layer6_outputs(316) <= not(layer5_outputs(50));
    layer6_outputs(317) <= not(layer5_outputs(2045)) or (layer5_outputs(2140));
    layer6_outputs(318) <= layer5_outputs(1100);
    layer6_outputs(319) <= not(layer5_outputs(105));
    layer6_outputs(320) <= not(layer5_outputs(1049));
    layer6_outputs(321) <= not(layer5_outputs(987)) or (layer5_outputs(1799));
    layer6_outputs(322) <= not(layer5_outputs(92));
    layer6_outputs(323) <= layer5_outputs(2085);
    layer6_outputs(324) <= not(layer5_outputs(1326));
    layer6_outputs(325) <= not(layer5_outputs(690)) or (layer5_outputs(2378));
    layer6_outputs(326) <= not(layer5_outputs(1573)) or (layer5_outputs(434));
    layer6_outputs(327) <= layer5_outputs(584);
    layer6_outputs(328) <= not(layer5_outputs(248));
    layer6_outputs(329) <= not((layer5_outputs(951)) xor (layer5_outputs(6)));
    layer6_outputs(330) <= not(layer5_outputs(1705));
    layer6_outputs(331) <= not(layer5_outputs(88));
    layer6_outputs(332) <= not(layer5_outputs(666));
    layer6_outputs(333) <= not(layer5_outputs(944));
    layer6_outputs(334) <= layer5_outputs(235);
    layer6_outputs(335) <= (layer5_outputs(1846)) and (layer5_outputs(128));
    layer6_outputs(336) <= not((layer5_outputs(35)) xor (layer5_outputs(1095)));
    layer6_outputs(337) <= not(layer5_outputs(1053));
    layer6_outputs(338) <= not((layer5_outputs(1442)) xor (layer5_outputs(2124)));
    layer6_outputs(339) <= not((layer5_outputs(1146)) or (layer5_outputs(2500)));
    layer6_outputs(340) <= layer5_outputs(763);
    layer6_outputs(341) <= layer5_outputs(1007);
    layer6_outputs(342) <= not(layer5_outputs(652));
    layer6_outputs(343) <= layer5_outputs(2316);
    layer6_outputs(344) <= (layer5_outputs(1334)) or (layer5_outputs(600));
    layer6_outputs(345) <= not(layer5_outputs(923)) or (layer5_outputs(1462));
    layer6_outputs(346) <= (layer5_outputs(1883)) and (layer5_outputs(971));
    layer6_outputs(347) <= not((layer5_outputs(2273)) and (layer5_outputs(1247)));
    layer6_outputs(348) <= layer5_outputs(2378);
    layer6_outputs(349) <= layer5_outputs(2441);
    layer6_outputs(350) <= not(layer5_outputs(66));
    layer6_outputs(351) <= (layer5_outputs(1522)) xor (layer5_outputs(156));
    layer6_outputs(352) <= not(layer5_outputs(377));
    layer6_outputs(353) <= not(layer5_outputs(933)) or (layer5_outputs(791));
    layer6_outputs(354) <= (layer5_outputs(435)) xor (layer5_outputs(93));
    layer6_outputs(355) <= layer5_outputs(491);
    layer6_outputs(356) <= not(layer5_outputs(1059));
    layer6_outputs(357) <= not((layer5_outputs(2112)) xor (layer5_outputs(396)));
    layer6_outputs(358) <= layer5_outputs(1239);
    layer6_outputs(359) <= not(layer5_outputs(1759));
    layer6_outputs(360) <= '0';
    layer6_outputs(361) <= layer5_outputs(1262);
    layer6_outputs(362) <= not(layer5_outputs(657));
    layer6_outputs(363) <= not(layer5_outputs(814)) or (layer5_outputs(505));
    layer6_outputs(364) <= not((layer5_outputs(2506)) xor (layer5_outputs(1387)));
    layer6_outputs(365) <= (layer5_outputs(1370)) xor (layer5_outputs(1738));
    layer6_outputs(366) <= layer5_outputs(421);
    layer6_outputs(367) <= not((layer5_outputs(956)) xor (layer5_outputs(2407)));
    layer6_outputs(368) <= layer5_outputs(1362);
    layer6_outputs(369) <= not(layer5_outputs(1389));
    layer6_outputs(370) <= not(layer5_outputs(223));
    layer6_outputs(371) <= not(layer5_outputs(1443));
    layer6_outputs(372) <= not(layer5_outputs(694)) or (layer5_outputs(1784));
    layer6_outputs(373) <= layer5_outputs(1491);
    layer6_outputs(374) <= not((layer5_outputs(206)) and (layer5_outputs(729)));
    layer6_outputs(375) <= not((layer5_outputs(2539)) xor (layer5_outputs(2515)));
    layer6_outputs(376) <= not((layer5_outputs(1860)) and (layer5_outputs(2431)));
    layer6_outputs(377) <= layer5_outputs(792);
    layer6_outputs(378) <= (layer5_outputs(699)) and not (layer5_outputs(1545));
    layer6_outputs(379) <= not(layer5_outputs(743));
    layer6_outputs(380) <= (layer5_outputs(2416)) xor (layer5_outputs(613));
    layer6_outputs(381) <= (layer5_outputs(1440)) xor (layer5_outputs(2299));
    layer6_outputs(382) <= not(layer5_outputs(168));
    layer6_outputs(383) <= not(layer5_outputs(2489));
    layer6_outputs(384) <= layer5_outputs(729);
    layer6_outputs(385) <= '1';
    layer6_outputs(386) <= not(layer5_outputs(1431));
    layer6_outputs(387) <= (layer5_outputs(306)) or (layer5_outputs(2181));
    layer6_outputs(388) <= not(layer5_outputs(1925));
    layer6_outputs(389) <= (layer5_outputs(578)) xor (layer5_outputs(548));
    layer6_outputs(390) <= not((layer5_outputs(772)) or (layer5_outputs(1711)));
    layer6_outputs(391) <= layer5_outputs(2536);
    layer6_outputs(392) <= layer5_outputs(2020);
    layer6_outputs(393) <= layer5_outputs(1306);
    layer6_outputs(394) <= not((layer5_outputs(470)) and (layer5_outputs(1242)));
    layer6_outputs(395) <= (layer5_outputs(2333)) xor (layer5_outputs(413));
    layer6_outputs(396) <= not(layer5_outputs(1)) or (layer5_outputs(715));
    layer6_outputs(397) <= (layer5_outputs(114)) and not (layer5_outputs(23));
    layer6_outputs(398) <= layer5_outputs(451);
    layer6_outputs(399) <= not((layer5_outputs(2079)) or (layer5_outputs(1888)));
    layer6_outputs(400) <= not(layer5_outputs(1260)) or (layer5_outputs(1458));
    layer6_outputs(401) <= (layer5_outputs(648)) and (layer5_outputs(835));
    layer6_outputs(402) <= not((layer5_outputs(2516)) or (layer5_outputs(170)));
    layer6_outputs(403) <= layer5_outputs(10);
    layer6_outputs(404) <= not((layer5_outputs(1245)) or (layer5_outputs(1995)));
    layer6_outputs(405) <= not(layer5_outputs(1849));
    layer6_outputs(406) <= '0';
    layer6_outputs(407) <= not(layer5_outputs(1395));
    layer6_outputs(408) <= (layer5_outputs(1622)) xor (layer5_outputs(1695));
    layer6_outputs(409) <= (layer5_outputs(1666)) xor (layer5_outputs(541));
    layer6_outputs(410) <= (layer5_outputs(2101)) and not (layer5_outputs(2433));
    layer6_outputs(411) <= not((layer5_outputs(1055)) xor (layer5_outputs(1005)));
    layer6_outputs(412) <= layer5_outputs(687);
    layer6_outputs(413) <= not(layer5_outputs(775));
    layer6_outputs(414) <= not(layer5_outputs(807));
    layer6_outputs(415) <= not(layer5_outputs(1541)) or (layer5_outputs(917));
    layer6_outputs(416) <= (layer5_outputs(1979)) and not (layer5_outputs(1854));
    layer6_outputs(417) <= (layer5_outputs(1853)) xor (layer5_outputs(2428));
    layer6_outputs(418) <= not((layer5_outputs(394)) xor (layer5_outputs(2217)));
    layer6_outputs(419) <= (layer5_outputs(257)) and (layer5_outputs(1240));
    layer6_outputs(420) <= (layer5_outputs(1275)) or (layer5_outputs(821));
    layer6_outputs(421) <= not(layer5_outputs(815));
    layer6_outputs(422) <= layer5_outputs(1311);
    layer6_outputs(423) <= layer5_outputs(1332);
    layer6_outputs(424) <= not(layer5_outputs(1697));
    layer6_outputs(425) <= not(layer5_outputs(2124));
    layer6_outputs(426) <= layer5_outputs(1426);
    layer6_outputs(427) <= (layer5_outputs(1257)) and (layer5_outputs(2068));
    layer6_outputs(428) <= layer5_outputs(403);
    layer6_outputs(429) <= (layer5_outputs(515)) and not (layer5_outputs(1770));
    layer6_outputs(430) <= layer5_outputs(414);
    layer6_outputs(431) <= (layer5_outputs(1633)) and not (layer5_outputs(1700));
    layer6_outputs(432) <= not(layer5_outputs(192));
    layer6_outputs(433) <= (layer5_outputs(123)) or (layer5_outputs(612));
    layer6_outputs(434) <= layer5_outputs(1536);
    layer6_outputs(435) <= not(layer5_outputs(1906));
    layer6_outputs(436) <= (layer5_outputs(365)) and (layer5_outputs(1684));
    layer6_outputs(437) <= (layer5_outputs(338)) xor (layer5_outputs(327));
    layer6_outputs(438) <= not(layer5_outputs(200));
    layer6_outputs(439) <= not((layer5_outputs(437)) and (layer5_outputs(166)));
    layer6_outputs(440) <= not(layer5_outputs(1677)) or (layer5_outputs(1689));
    layer6_outputs(441) <= '0';
    layer6_outputs(442) <= not(layer5_outputs(2084));
    layer6_outputs(443) <= layer5_outputs(1081);
    layer6_outputs(444) <= layer5_outputs(2172);
    layer6_outputs(445) <= not((layer5_outputs(918)) and (layer5_outputs(1138)));
    layer6_outputs(446) <= layer5_outputs(125);
    layer6_outputs(447) <= layer5_outputs(1558);
    layer6_outputs(448) <= not(layer5_outputs(1174));
    layer6_outputs(449) <= not((layer5_outputs(221)) or (layer5_outputs(739)));
    layer6_outputs(450) <= layer5_outputs(1121);
    layer6_outputs(451) <= not(layer5_outputs(679));
    layer6_outputs(452) <= not(layer5_outputs(941));
    layer6_outputs(453) <= (layer5_outputs(1761)) and not (layer5_outputs(1403));
    layer6_outputs(454) <= layer5_outputs(1716);
    layer6_outputs(455) <= (layer5_outputs(2003)) and not (layer5_outputs(1761));
    layer6_outputs(456) <= (layer5_outputs(2335)) and (layer5_outputs(846));
    layer6_outputs(457) <= not((layer5_outputs(714)) and (layer5_outputs(142)));
    layer6_outputs(458) <= not((layer5_outputs(1871)) or (layer5_outputs(163)));
    layer6_outputs(459) <= layer5_outputs(1600);
    layer6_outputs(460) <= layer5_outputs(1269);
    layer6_outputs(461) <= layer5_outputs(1167);
    layer6_outputs(462) <= layer5_outputs(2386);
    layer6_outputs(463) <= layer5_outputs(1074);
    layer6_outputs(464) <= (layer5_outputs(844)) xor (layer5_outputs(566));
    layer6_outputs(465) <= not(layer5_outputs(1523)) or (layer5_outputs(36));
    layer6_outputs(466) <= (layer5_outputs(95)) and not (layer5_outputs(1796));
    layer6_outputs(467) <= layer5_outputs(1290);
    layer6_outputs(468) <= not(layer5_outputs(1940)) or (layer5_outputs(656));
    layer6_outputs(469) <= not(layer5_outputs(378)) or (layer5_outputs(1535));
    layer6_outputs(470) <= not(layer5_outputs(1199));
    layer6_outputs(471) <= not((layer5_outputs(2513)) xor (layer5_outputs(2543)));
    layer6_outputs(472) <= not((layer5_outputs(81)) xor (layer5_outputs(13)));
    layer6_outputs(473) <= layer5_outputs(1687);
    layer6_outputs(474) <= (layer5_outputs(1804)) or (layer5_outputs(234));
    layer6_outputs(475) <= layer5_outputs(387);
    layer6_outputs(476) <= (layer5_outputs(462)) or (layer5_outputs(1816));
    layer6_outputs(477) <= (layer5_outputs(320)) and not (layer5_outputs(2200));
    layer6_outputs(478) <= not(layer5_outputs(1264));
    layer6_outputs(479) <= not(layer5_outputs(1603));
    layer6_outputs(480) <= (layer5_outputs(549)) xor (layer5_outputs(1521));
    layer6_outputs(481) <= not((layer5_outputs(1369)) and (layer5_outputs(2182)));
    layer6_outputs(482) <= not(layer5_outputs(1305));
    layer6_outputs(483) <= not(layer5_outputs(1634));
    layer6_outputs(484) <= not(layer5_outputs(2132));
    layer6_outputs(485) <= not((layer5_outputs(312)) and (layer5_outputs(2412)));
    layer6_outputs(486) <= layer5_outputs(1570);
    layer6_outputs(487) <= not(layer5_outputs(68));
    layer6_outputs(488) <= (layer5_outputs(1272)) xor (layer5_outputs(2123));
    layer6_outputs(489) <= not(layer5_outputs(422));
    layer6_outputs(490) <= not(layer5_outputs(803));
    layer6_outputs(491) <= not((layer5_outputs(704)) or (layer5_outputs(179)));
    layer6_outputs(492) <= not(layer5_outputs(2326));
    layer6_outputs(493) <= not(layer5_outputs(499));
    layer6_outputs(494) <= layer5_outputs(2210);
    layer6_outputs(495) <= not(layer5_outputs(2011)) or (layer5_outputs(299));
    layer6_outputs(496) <= (layer5_outputs(1845)) xor (layer5_outputs(111));
    layer6_outputs(497) <= (layer5_outputs(1378)) and not (layer5_outputs(1986));
    layer6_outputs(498) <= (layer5_outputs(1001)) or (layer5_outputs(541));
    layer6_outputs(499) <= not(layer5_outputs(2226)) or (layer5_outputs(363));
    layer6_outputs(500) <= (layer5_outputs(1172)) and (layer5_outputs(1571));
    layer6_outputs(501) <= not(layer5_outputs(2508));
    layer6_outputs(502) <= layer5_outputs(1291);
    layer6_outputs(503) <= layer5_outputs(2162);
    layer6_outputs(504) <= not((layer5_outputs(765)) or (layer5_outputs(1165)));
    layer6_outputs(505) <= not(layer5_outputs(1286));
    layer6_outputs(506) <= (layer5_outputs(872)) and not (layer5_outputs(2100));
    layer6_outputs(507) <= not(layer5_outputs(2167)) or (layer5_outputs(133));
    layer6_outputs(508) <= (layer5_outputs(2313)) and (layer5_outputs(2274));
    layer6_outputs(509) <= layer5_outputs(101);
    layer6_outputs(510) <= not((layer5_outputs(5)) or (layer5_outputs(2065)));
    layer6_outputs(511) <= not((layer5_outputs(1739)) and (layer5_outputs(259)));
    layer6_outputs(512) <= layer5_outputs(349);
    layer6_outputs(513) <= layer5_outputs(1339);
    layer6_outputs(514) <= layer5_outputs(407);
    layer6_outputs(515) <= not(layer5_outputs(2143)) or (layer5_outputs(1008));
    layer6_outputs(516) <= layer5_outputs(741);
    layer6_outputs(517) <= not(layer5_outputs(737));
    layer6_outputs(518) <= (layer5_outputs(378)) or (layer5_outputs(2227));
    layer6_outputs(519) <= not(layer5_outputs(1881));
    layer6_outputs(520) <= not(layer5_outputs(1173));
    layer6_outputs(521) <= not(layer5_outputs(1165));
    layer6_outputs(522) <= not((layer5_outputs(792)) or (layer5_outputs(1647)));
    layer6_outputs(523) <= layer5_outputs(1901);
    layer6_outputs(524) <= layer5_outputs(2028);
    layer6_outputs(525) <= (layer5_outputs(2098)) and (layer5_outputs(750));
    layer6_outputs(526) <= (layer5_outputs(1650)) and not (layer5_outputs(187));
    layer6_outputs(527) <= layer5_outputs(908);
    layer6_outputs(528) <= layer5_outputs(2418);
    layer6_outputs(529) <= not(layer5_outputs(178));
    layer6_outputs(530) <= not(layer5_outputs(1814));
    layer6_outputs(531) <= not((layer5_outputs(1652)) xor (layer5_outputs(597)));
    layer6_outputs(532) <= layer5_outputs(2191);
    layer6_outputs(533) <= not((layer5_outputs(2072)) or (layer5_outputs(531)));
    layer6_outputs(534) <= not(layer5_outputs(1850));
    layer6_outputs(535) <= (layer5_outputs(2514)) and (layer5_outputs(2355));
    layer6_outputs(536) <= not(layer5_outputs(2091));
    layer6_outputs(537) <= not((layer5_outputs(2504)) xor (layer5_outputs(434)));
    layer6_outputs(538) <= '0';
    layer6_outputs(539) <= (layer5_outputs(1972)) and not (layer5_outputs(633));
    layer6_outputs(540) <= (layer5_outputs(734)) or (layer5_outputs(1768));
    layer6_outputs(541) <= not(layer5_outputs(720));
    layer6_outputs(542) <= layer5_outputs(397);
    layer6_outputs(543) <= layer5_outputs(246);
    layer6_outputs(544) <= (layer5_outputs(1409)) and (layer5_outputs(75));
    layer6_outputs(545) <= layer5_outputs(716);
    layer6_outputs(546) <= not(layer5_outputs(1465));
    layer6_outputs(547) <= not(layer5_outputs(309));
    layer6_outputs(548) <= not((layer5_outputs(1098)) xor (layer5_outputs(1882)));
    layer6_outputs(549) <= (layer5_outputs(1741)) and (layer5_outputs(210));
    layer6_outputs(550) <= layer5_outputs(364);
    layer6_outputs(551) <= (layer5_outputs(1354)) and (layer5_outputs(1999));
    layer6_outputs(552) <= '1';
    layer6_outputs(553) <= not(layer5_outputs(1757)) or (layer5_outputs(1540));
    layer6_outputs(554) <= not(layer5_outputs(452));
    layer6_outputs(555) <= not(layer5_outputs(983)) or (layer5_outputs(13));
    layer6_outputs(556) <= not(layer5_outputs(2548));
    layer6_outputs(557) <= not(layer5_outputs(1594)) or (layer5_outputs(1037));
    layer6_outputs(558) <= layer5_outputs(1462);
    layer6_outputs(559) <= not((layer5_outputs(718)) and (layer5_outputs(2389)));
    layer6_outputs(560) <= layer5_outputs(483);
    layer6_outputs(561) <= layer5_outputs(394);
    layer6_outputs(562) <= not(layer5_outputs(1364)) or (layer5_outputs(838));
    layer6_outputs(563) <= not(layer5_outputs(1877)) or (layer5_outputs(1448));
    layer6_outputs(564) <= not((layer5_outputs(2059)) and (layer5_outputs(129)));
    layer6_outputs(565) <= not(layer5_outputs(1052));
    layer6_outputs(566) <= (layer5_outputs(360)) and (layer5_outputs(1840));
    layer6_outputs(567) <= not(layer5_outputs(1117)) or (layer5_outputs(586));
    layer6_outputs(568) <= layer5_outputs(1288);
    layer6_outputs(569) <= not((layer5_outputs(2454)) and (layer5_outputs(1543)));
    layer6_outputs(570) <= not(layer5_outputs(1466));
    layer6_outputs(571) <= not((layer5_outputs(181)) and (layer5_outputs(1115)));
    layer6_outputs(572) <= (layer5_outputs(115)) and not (layer5_outputs(1566));
    layer6_outputs(573) <= not((layer5_outputs(606)) and (layer5_outputs(1009)));
    layer6_outputs(574) <= not(layer5_outputs(893));
    layer6_outputs(575) <= layer5_outputs(1893);
    layer6_outputs(576) <= not(layer5_outputs(148)) or (layer5_outputs(1870));
    layer6_outputs(577) <= layer5_outputs(1582);
    layer6_outputs(578) <= (layer5_outputs(354)) and (layer5_outputs(1230));
    layer6_outputs(579) <= (layer5_outputs(2220)) xor (layer5_outputs(1443));
    layer6_outputs(580) <= layer5_outputs(2547);
    layer6_outputs(581) <= (layer5_outputs(1214)) xor (layer5_outputs(1885));
    layer6_outputs(582) <= not((layer5_outputs(405)) or (layer5_outputs(1832)));
    layer6_outputs(583) <= not((layer5_outputs(265)) xor (layer5_outputs(1221)));
    layer6_outputs(584) <= not((layer5_outputs(131)) xor (layer5_outputs(1452)));
    layer6_outputs(585) <= not((layer5_outputs(1388)) or (layer5_outputs(2097)));
    layer6_outputs(586) <= layer5_outputs(775);
    layer6_outputs(587) <= layer5_outputs(1968);
    layer6_outputs(588) <= '1';
    layer6_outputs(589) <= (layer5_outputs(1123)) and not (layer5_outputs(2424));
    layer6_outputs(590) <= (layer5_outputs(871)) and not (layer5_outputs(2056));
    layer6_outputs(591) <= (layer5_outputs(889)) or (layer5_outputs(233));
    layer6_outputs(592) <= not(layer5_outputs(292)) or (layer5_outputs(543));
    layer6_outputs(593) <= not(layer5_outputs(1159));
    layer6_outputs(594) <= '1';
    layer6_outputs(595) <= not(layer5_outputs(633)) or (layer5_outputs(1953));
    layer6_outputs(596) <= not((layer5_outputs(1280)) and (layer5_outputs(1937)));
    layer6_outputs(597) <= not(layer5_outputs(827));
    layer6_outputs(598) <= layer5_outputs(261);
    layer6_outputs(599) <= (layer5_outputs(803)) xor (layer5_outputs(1601));
    layer6_outputs(600) <= layer5_outputs(2380);
    layer6_outputs(601) <= (layer5_outputs(1328)) or (layer5_outputs(884));
    layer6_outputs(602) <= layer5_outputs(2115);
    layer6_outputs(603) <= not(layer5_outputs(2265));
    layer6_outputs(604) <= not(layer5_outputs(1273));
    layer6_outputs(605) <= not(layer5_outputs(2155)) or (layer5_outputs(2102));
    layer6_outputs(606) <= layer5_outputs(1133);
    layer6_outputs(607) <= not((layer5_outputs(99)) or (layer5_outputs(2008)));
    layer6_outputs(608) <= not(layer5_outputs(570)) or (layer5_outputs(805));
    layer6_outputs(609) <= layer5_outputs(1180);
    layer6_outputs(610) <= not((layer5_outputs(1378)) and (layer5_outputs(1071)));
    layer6_outputs(611) <= not(layer5_outputs(1769));
    layer6_outputs(612) <= (layer5_outputs(935)) xor (layer5_outputs(635));
    layer6_outputs(613) <= not(layer5_outputs(1706)) or (layer5_outputs(1087));
    layer6_outputs(614) <= '1';
    layer6_outputs(615) <= layer5_outputs(793);
    layer6_outputs(616) <= layer5_outputs(1145);
    layer6_outputs(617) <= (layer5_outputs(975)) and not (layer5_outputs(328));
    layer6_outputs(618) <= not(layer5_outputs(1199));
    layer6_outputs(619) <= not(layer5_outputs(1909));
    layer6_outputs(620) <= not(layer5_outputs(2163)) or (layer5_outputs(2257));
    layer6_outputs(621) <= not((layer5_outputs(242)) xor (layer5_outputs(468)));
    layer6_outputs(622) <= not((layer5_outputs(249)) and (layer5_outputs(248)));
    layer6_outputs(623) <= not(layer5_outputs(2540));
    layer6_outputs(624) <= (layer5_outputs(1848)) or (layer5_outputs(698));
    layer6_outputs(625) <= not(layer5_outputs(977));
    layer6_outputs(626) <= (layer5_outputs(1074)) and not (layer5_outputs(1657));
    layer6_outputs(627) <= (layer5_outputs(2150)) or (layer5_outputs(1042));
    layer6_outputs(628) <= (layer5_outputs(128)) and not (layer5_outputs(1532));
    layer6_outputs(629) <= not(layer5_outputs(348));
    layer6_outputs(630) <= layer5_outputs(2091);
    layer6_outputs(631) <= layer5_outputs(83);
    layer6_outputs(632) <= layer5_outputs(1782);
    layer6_outputs(633) <= not(layer5_outputs(1107));
    layer6_outputs(634) <= (layer5_outputs(2116)) and not (layer5_outputs(1490));
    layer6_outputs(635) <= not(layer5_outputs(1117));
    layer6_outputs(636) <= '1';
    layer6_outputs(637) <= (layer5_outputs(1992)) xor (layer5_outputs(2331));
    layer6_outputs(638) <= not(layer5_outputs(1075));
    layer6_outputs(639) <= (layer5_outputs(2341)) and not (layer5_outputs(849));
    layer6_outputs(640) <= '0';
    layer6_outputs(641) <= (layer5_outputs(2413)) and not (layer5_outputs(1843));
    layer6_outputs(642) <= not((layer5_outputs(897)) and (layer5_outputs(1381)));
    layer6_outputs(643) <= layer5_outputs(489);
    layer6_outputs(644) <= layer5_outputs(1590);
    layer6_outputs(645) <= layer5_outputs(1160);
    layer6_outputs(646) <= layer5_outputs(1629);
    layer6_outputs(647) <= not(layer5_outputs(2519)) or (layer5_outputs(2034));
    layer6_outputs(648) <= (layer5_outputs(2033)) xor (layer5_outputs(617));
    layer6_outputs(649) <= not(layer5_outputs(1608)) or (layer5_outputs(500));
    layer6_outputs(650) <= not(layer5_outputs(2001));
    layer6_outputs(651) <= (layer5_outputs(742)) and not (layer5_outputs(1733));
    layer6_outputs(652) <= (layer5_outputs(1833)) and (layer5_outputs(994));
    layer6_outputs(653) <= (layer5_outputs(1714)) and not (layer5_outputs(2297));
    layer6_outputs(654) <= (layer5_outputs(219)) and not (layer5_outputs(789));
    layer6_outputs(655) <= not((layer5_outputs(685)) xor (layer5_outputs(2008)));
    layer6_outputs(656) <= layer5_outputs(724);
    layer6_outputs(657) <= not(layer5_outputs(594));
    layer6_outputs(658) <= not(layer5_outputs(927));
    layer6_outputs(659) <= not(layer5_outputs(2065));
    layer6_outputs(660) <= (layer5_outputs(1051)) and not (layer5_outputs(1452));
    layer6_outputs(661) <= layer5_outputs(684);
    layer6_outputs(662) <= not((layer5_outputs(924)) or (layer5_outputs(2311)));
    layer6_outputs(663) <= layer5_outputs(2427);
    layer6_outputs(664) <= (layer5_outputs(1574)) or (layer5_outputs(2384));
    layer6_outputs(665) <= layer5_outputs(1893);
    layer6_outputs(666) <= layer5_outputs(1256);
    layer6_outputs(667) <= not(layer5_outputs(150));
    layer6_outputs(668) <= not((layer5_outputs(1802)) xor (layer5_outputs(896)));
    layer6_outputs(669) <= not(layer5_outputs(2010));
    layer6_outputs(670) <= (layer5_outputs(2482)) xor (layer5_outputs(2430));
    layer6_outputs(671) <= (layer5_outputs(2)) xor (layer5_outputs(2402));
    layer6_outputs(672) <= not(layer5_outputs(2110)) or (layer5_outputs(1566));
    layer6_outputs(673) <= (layer5_outputs(882)) and not (layer5_outputs(1688));
    layer6_outputs(674) <= (layer5_outputs(1046)) or (layer5_outputs(776));
    layer6_outputs(675) <= (layer5_outputs(1033)) and (layer5_outputs(1310));
    layer6_outputs(676) <= layer5_outputs(1457);
    layer6_outputs(677) <= not(layer5_outputs(1887)) or (layer5_outputs(1513));
    layer6_outputs(678) <= not(layer5_outputs(1478));
    layer6_outputs(679) <= not((layer5_outputs(679)) xor (layer5_outputs(1704)));
    layer6_outputs(680) <= (layer5_outputs(2557)) and not (layer5_outputs(1210));
    layer6_outputs(681) <= layer5_outputs(720);
    layer6_outputs(682) <= not(layer5_outputs(2352));
    layer6_outputs(683) <= not((layer5_outputs(1855)) and (layer5_outputs(2286)));
    layer6_outputs(684) <= (layer5_outputs(1122)) xor (layer5_outputs(141));
    layer6_outputs(685) <= not(layer5_outputs(122)) or (layer5_outputs(336));
    layer6_outputs(686) <= not(layer5_outputs(2181)) or (layer5_outputs(2219));
    layer6_outputs(687) <= layer5_outputs(1484);
    layer6_outputs(688) <= (layer5_outputs(997)) and not (layer5_outputs(102));
    layer6_outputs(689) <= (layer5_outputs(1156)) xor (layer5_outputs(393));
    layer6_outputs(690) <= not((layer5_outputs(77)) or (layer5_outputs(2064)));
    layer6_outputs(691) <= not(layer5_outputs(895));
    layer6_outputs(692) <= layer5_outputs(935);
    layer6_outputs(693) <= not(layer5_outputs(2492)) or (layer5_outputs(2024));
    layer6_outputs(694) <= (layer5_outputs(599)) xor (layer5_outputs(2166));
    layer6_outputs(695) <= not(layer5_outputs(579));
    layer6_outputs(696) <= layer5_outputs(1206);
    layer6_outputs(697) <= layer5_outputs(2014);
    layer6_outputs(698) <= (layer5_outputs(1901)) xor (layer5_outputs(1846));
    layer6_outputs(699) <= not((layer5_outputs(344)) xor (layer5_outputs(1025)));
    layer6_outputs(700) <= layer5_outputs(1451);
    layer6_outputs(701) <= not(layer5_outputs(410));
    layer6_outputs(702) <= layer5_outputs(2516);
    layer6_outputs(703) <= not((layer5_outputs(2111)) xor (layer5_outputs(1868)));
    layer6_outputs(704) <= layer5_outputs(1010);
    layer6_outputs(705) <= (layer5_outputs(2039)) or (layer5_outputs(2195));
    layer6_outputs(706) <= not(layer5_outputs(454));
    layer6_outputs(707) <= (layer5_outputs(1495)) or (layer5_outputs(1891));
    layer6_outputs(708) <= not((layer5_outputs(444)) xor (layer5_outputs(962)));
    layer6_outputs(709) <= (layer5_outputs(1860)) and (layer5_outputs(357));
    layer6_outputs(710) <= not(layer5_outputs(279)) or (layer5_outputs(853));
    layer6_outputs(711) <= layer5_outputs(400);
    layer6_outputs(712) <= (layer5_outputs(411)) and (layer5_outputs(1547));
    layer6_outputs(713) <= not(layer5_outputs(165));
    layer6_outputs(714) <= (layer5_outputs(1459)) xor (layer5_outputs(2115));
    layer6_outputs(715) <= layer5_outputs(1500);
    layer6_outputs(716) <= layer5_outputs(1384);
    layer6_outputs(717) <= not(layer5_outputs(255));
    layer6_outputs(718) <= (layer5_outputs(939)) xor (layer5_outputs(1454));
    layer6_outputs(719) <= layer5_outputs(147);
    layer6_outputs(720) <= layer5_outputs(310);
    layer6_outputs(721) <= not((layer5_outputs(1395)) or (layer5_outputs(2047)));
    layer6_outputs(722) <= not(layer5_outputs(1446)) or (layer5_outputs(2073));
    layer6_outputs(723) <= not((layer5_outputs(1106)) and (layer5_outputs(2453)));
    layer6_outputs(724) <= not((layer5_outputs(1659)) and (layer5_outputs(273)));
    layer6_outputs(725) <= not(layer5_outputs(1604));
    layer6_outputs(726) <= (layer5_outputs(1368)) or (layer5_outputs(1623));
    layer6_outputs(727) <= layer5_outputs(900);
    layer6_outputs(728) <= layer5_outputs(202);
    layer6_outputs(729) <= (layer5_outputs(1626)) or (layer5_outputs(2074));
    layer6_outputs(730) <= (layer5_outputs(1728)) xor (layer5_outputs(593));
    layer6_outputs(731) <= (layer5_outputs(107)) xor (layer5_outputs(1029));
    layer6_outputs(732) <= layer5_outputs(598);
    layer6_outputs(733) <= layer5_outputs(536);
    layer6_outputs(734) <= not(layer5_outputs(1050));
    layer6_outputs(735) <= (layer5_outputs(1521)) and (layer5_outputs(764));
    layer6_outputs(736) <= not(layer5_outputs(582)) or (layer5_outputs(1746));
    layer6_outputs(737) <= layer5_outputs(915);
    layer6_outputs(738) <= layer5_outputs(2317);
    layer6_outputs(739) <= not((layer5_outputs(1875)) xor (layer5_outputs(1385)));
    layer6_outputs(740) <= not(layer5_outputs(1487));
    layer6_outputs(741) <= not((layer5_outputs(2071)) xor (layer5_outputs(1307)));
    layer6_outputs(742) <= not(layer5_outputs(1916));
    layer6_outputs(743) <= (layer5_outputs(453)) xor (layer5_outputs(1020));
    layer6_outputs(744) <= (layer5_outputs(2057)) and (layer5_outputs(974));
    layer6_outputs(745) <= not(layer5_outputs(484));
    layer6_outputs(746) <= not(layer5_outputs(500));
    layer6_outputs(747) <= not(layer5_outputs(530));
    layer6_outputs(748) <= not(layer5_outputs(588)) or (layer5_outputs(639));
    layer6_outputs(749) <= not(layer5_outputs(747));
    layer6_outputs(750) <= (layer5_outputs(1453)) and (layer5_outputs(358));
    layer6_outputs(751) <= not(layer5_outputs(2501));
    layer6_outputs(752) <= (layer5_outputs(175)) and not (layer5_outputs(828));
    layer6_outputs(753) <= layer5_outputs(1833);
    layer6_outputs(754) <= not(layer5_outputs(1691));
    layer6_outputs(755) <= (layer5_outputs(2269)) and (layer5_outputs(524));
    layer6_outputs(756) <= not(layer5_outputs(1510));
    layer6_outputs(757) <= not(layer5_outputs(1287));
    layer6_outputs(758) <= not(layer5_outputs(976));
    layer6_outputs(759) <= layer5_outputs(2277);
    layer6_outputs(760) <= (layer5_outputs(894)) and (layer5_outputs(2397));
    layer6_outputs(761) <= (layer5_outputs(2336)) and (layer5_outputs(668));
    layer6_outputs(762) <= not(layer5_outputs(2456));
    layer6_outputs(763) <= layer5_outputs(2130);
    layer6_outputs(764) <= not(layer5_outputs(799)) or (layer5_outputs(180));
    layer6_outputs(765) <= layer5_outputs(2187);
    layer6_outputs(766) <= not(layer5_outputs(215));
    layer6_outputs(767) <= layer5_outputs(1128);
    layer6_outputs(768) <= not((layer5_outputs(1099)) or (layer5_outputs(608)));
    layer6_outputs(769) <= layer5_outputs(779);
    layer6_outputs(770) <= layer5_outputs(1958);
    layer6_outputs(771) <= '1';
    layer6_outputs(772) <= layer5_outputs(872);
    layer6_outputs(773) <= not(layer5_outputs(1190));
    layer6_outputs(774) <= not((layer5_outputs(1007)) or (layer5_outputs(352)));
    layer6_outputs(775) <= not((layer5_outputs(2107)) and (layer5_outputs(1629)));
    layer6_outputs(776) <= not(layer5_outputs(108));
    layer6_outputs(777) <= (layer5_outputs(2296)) and not (layer5_outputs(1528));
    layer6_outputs(778) <= not((layer5_outputs(776)) and (layer5_outputs(22)));
    layer6_outputs(779) <= not(layer5_outputs(1313));
    layer6_outputs(780) <= (layer5_outputs(911)) and (layer5_outputs(2426));
    layer6_outputs(781) <= (layer5_outputs(1258)) and not (layer5_outputs(55));
    layer6_outputs(782) <= not(layer5_outputs(1506));
    layer6_outputs(783) <= layer5_outputs(1163);
    layer6_outputs(784) <= layer5_outputs(92);
    layer6_outputs(785) <= not(layer5_outputs(617));
    layer6_outputs(786) <= not(layer5_outputs(2344));
    layer6_outputs(787) <= not((layer5_outputs(240)) xor (layer5_outputs(686)));
    layer6_outputs(788) <= not(layer5_outputs(77));
    layer6_outputs(789) <= '0';
    layer6_outputs(790) <= not(layer5_outputs(2108)) or (layer5_outputs(680));
    layer6_outputs(791) <= not(layer5_outputs(1219));
    layer6_outputs(792) <= layer5_outputs(1058);
    layer6_outputs(793) <= (layer5_outputs(267)) and not (layer5_outputs(1468));
    layer6_outputs(794) <= not(layer5_outputs(818));
    layer6_outputs(795) <= not(layer5_outputs(2446));
    layer6_outputs(796) <= (layer5_outputs(858)) and not (layer5_outputs(1321));
    layer6_outputs(797) <= layer5_outputs(2221);
    layer6_outputs(798) <= layer5_outputs(203);
    layer6_outputs(799) <= not((layer5_outputs(2373)) and (layer5_outputs(589)));
    layer6_outputs(800) <= layer5_outputs(2256);
    layer6_outputs(801) <= not(layer5_outputs(906)) or (layer5_outputs(1261));
    layer6_outputs(802) <= layer5_outputs(505);
    layer6_outputs(803) <= not(layer5_outputs(900));
    layer6_outputs(804) <= not(layer5_outputs(1774)) or (layer5_outputs(2376));
    layer6_outputs(805) <= (layer5_outputs(2229)) and not (layer5_outputs(2320));
    layer6_outputs(806) <= (layer5_outputs(30)) xor (layer5_outputs(1221));
    layer6_outputs(807) <= layer5_outputs(1585);
    layer6_outputs(808) <= layer5_outputs(2204);
    layer6_outputs(809) <= (layer5_outputs(1704)) and (layer5_outputs(1612));
    layer6_outputs(810) <= (layer5_outputs(643)) and not (layer5_outputs(962));
    layer6_outputs(811) <= not(layer5_outputs(658)) or (layer5_outputs(2109));
    layer6_outputs(812) <= not(layer5_outputs(2285));
    layer6_outputs(813) <= not((layer5_outputs(339)) and (layer5_outputs(1730)));
    layer6_outputs(814) <= not(layer5_outputs(1483)) or (layer5_outputs(1432));
    layer6_outputs(815) <= not((layer5_outputs(1084)) and (layer5_outputs(2016)));
    layer6_outputs(816) <= not((layer5_outputs(1977)) or (layer5_outputs(756)));
    layer6_outputs(817) <= not((layer5_outputs(2502)) xor (layer5_outputs(569)));
    layer6_outputs(818) <= layer5_outputs(1324);
    layer6_outputs(819) <= layer5_outputs(931);
    layer6_outputs(820) <= not((layer5_outputs(1735)) or (layer5_outputs(98)));
    layer6_outputs(821) <= not(layer5_outputs(1910));
    layer6_outputs(822) <= not(layer5_outputs(1044)) or (layer5_outputs(42));
    layer6_outputs(823) <= not(layer5_outputs(1373));
    layer6_outputs(824) <= (layer5_outputs(1938)) and not (layer5_outputs(2108));
    layer6_outputs(825) <= layer5_outputs(2190);
    layer6_outputs(826) <= layer5_outputs(2341);
    layer6_outputs(827) <= (layer5_outputs(2535)) or (layer5_outputs(425));
    layer6_outputs(828) <= not(layer5_outputs(2125)) or (layer5_outputs(34));
    layer6_outputs(829) <= not((layer5_outputs(2216)) and (layer5_outputs(875)));
    layer6_outputs(830) <= not(layer5_outputs(259));
    layer6_outputs(831) <= not((layer5_outputs(1470)) xor (layer5_outputs(1533)));
    layer6_outputs(832) <= not(layer5_outputs(156));
    layer6_outputs(833) <= layer5_outputs(1089);
    layer6_outputs(834) <= layer5_outputs(8);
    layer6_outputs(835) <= not(layer5_outputs(2410));
    layer6_outputs(836) <= not(layer5_outputs(2206));
    layer6_outputs(837) <= (layer5_outputs(760)) and not (layer5_outputs(2287));
    layer6_outputs(838) <= not((layer5_outputs(1880)) xor (layer5_outputs(2237)));
    layer6_outputs(839) <= not(layer5_outputs(2536));
    layer6_outputs(840) <= layer5_outputs(796);
    layer6_outputs(841) <= layer5_outputs(996);
    layer6_outputs(842) <= layer5_outputs(1680);
    layer6_outputs(843) <= (layer5_outputs(801)) and (layer5_outputs(1678));
    layer6_outputs(844) <= layer5_outputs(2523);
    layer6_outputs(845) <= (layer5_outputs(381)) and (layer5_outputs(1780));
    layer6_outputs(846) <= not(layer5_outputs(1073));
    layer6_outputs(847) <= not((layer5_outputs(910)) xor (layer5_outputs(964)));
    layer6_outputs(848) <= not((layer5_outputs(1286)) xor (layer5_outputs(327)));
    layer6_outputs(849) <= not(layer5_outputs(1657)) or (layer5_outputs(1609));
    layer6_outputs(850) <= not(layer5_outputs(1347));
    layer6_outputs(851) <= not(layer5_outputs(62));
    layer6_outputs(852) <= not(layer5_outputs(861));
    layer6_outputs(853) <= not((layer5_outputs(2183)) xor (layer5_outputs(301)));
    layer6_outputs(854) <= not((layer5_outputs(1016)) or (layer5_outputs(1264)));
    layer6_outputs(855) <= not(layer5_outputs(1752));
    layer6_outputs(856) <= not((layer5_outputs(1862)) and (layer5_outputs(983)));
    layer6_outputs(857) <= layer5_outputs(2457);
    layer6_outputs(858) <= not(layer5_outputs(448));
    layer6_outputs(859) <= not(layer5_outputs(1482));
    layer6_outputs(860) <= layer5_outputs(2490);
    layer6_outputs(861) <= not((layer5_outputs(616)) and (layer5_outputs(837)));
    layer6_outputs(862) <= layer5_outputs(2173);
    layer6_outputs(863) <= (layer5_outputs(886)) xor (layer5_outputs(1002));
    layer6_outputs(864) <= (layer5_outputs(72)) and not (layer5_outputs(2484));
    layer6_outputs(865) <= not(layer5_outputs(2001)) or (layer5_outputs(27));
    layer6_outputs(866) <= not((layer5_outputs(484)) or (layer5_outputs(1115)));
    layer6_outputs(867) <= not((layer5_outputs(1486)) or (layer5_outputs(461)));
    layer6_outputs(868) <= not(layer5_outputs(404));
    layer6_outputs(869) <= not(layer5_outputs(561)) or (layer5_outputs(1283));
    layer6_outputs(870) <= layer5_outputs(1012);
    layer6_outputs(871) <= not(layer5_outputs(1278)) or (layer5_outputs(788));
    layer6_outputs(872) <= (layer5_outputs(1266)) and not (layer5_outputs(1391));
    layer6_outputs(873) <= not(layer5_outputs(2056));
    layer6_outputs(874) <= not(layer5_outputs(2012));
    layer6_outputs(875) <= layer5_outputs(1663);
    layer6_outputs(876) <= layer5_outputs(1309);
    layer6_outputs(877) <= layer5_outputs(1392);
    layer6_outputs(878) <= not((layer5_outputs(2316)) xor (layer5_outputs(1771)));
    layer6_outputs(879) <= layer5_outputs(1514);
    layer6_outputs(880) <= not(layer5_outputs(1785));
    layer6_outputs(881) <= layer5_outputs(44);
    layer6_outputs(882) <= (layer5_outputs(236)) xor (layer5_outputs(2049));
    layer6_outputs(883) <= (layer5_outputs(713)) and not (layer5_outputs(1669));
    layer6_outputs(884) <= not((layer5_outputs(745)) and (layer5_outputs(1157)));
    layer6_outputs(885) <= (layer5_outputs(1836)) and not (layer5_outputs(1598));
    layer6_outputs(886) <= (layer5_outputs(1773)) xor (layer5_outputs(2006));
    layer6_outputs(887) <= not((layer5_outputs(1871)) and (layer5_outputs(829)));
    layer6_outputs(888) <= layer5_outputs(1987);
    layer6_outputs(889) <= (layer5_outputs(37)) or (layer5_outputs(1410));
    layer6_outputs(890) <= (layer5_outputs(1847)) and not (layer5_outputs(1902));
    layer6_outputs(891) <= not(layer5_outputs(1272));
    layer6_outputs(892) <= not(layer5_outputs(878));
    layer6_outputs(893) <= not((layer5_outputs(1170)) and (layer5_outputs(1856)));
    layer6_outputs(894) <= layer5_outputs(1145);
    layer6_outputs(895) <= not(layer5_outputs(1416));
    layer6_outputs(896) <= '0';
    layer6_outputs(897) <= (layer5_outputs(2425)) xor (layer5_outputs(2095));
    layer6_outputs(898) <= (layer5_outputs(2024)) xor (layer5_outputs(1138));
    layer6_outputs(899) <= not(layer5_outputs(1125));
    layer6_outputs(900) <= layer5_outputs(1676);
    layer6_outputs(901) <= not(layer5_outputs(2520));
    layer6_outputs(902) <= not(layer5_outputs(515));
    layer6_outputs(903) <= layer5_outputs(1125);
    layer6_outputs(904) <= (layer5_outputs(2358)) xor (layer5_outputs(1291));
    layer6_outputs(905) <= (layer5_outputs(1722)) and not (layer5_outputs(411));
    layer6_outputs(906) <= not(layer5_outputs(1812));
    layer6_outputs(907) <= not(layer5_outputs(1904)) or (layer5_outputs(818));
    layer6_outputs(908) <= not((layer5_outputs(2385)) and (layer5_outputs(228)));
    layer6_outputs(909) <= layer5_outputs(437);
    layer6_outputs(910) <= not(layer5_outputs(1570)) or (layer5_outputs(2268));
    layer6_outputs(911) <= not(layer5_outputs(1488));
    layer6_outputs(912) <= not((layer5_outputs(1223)) or (layer5_outputs(413)));
    layer6_outputs(913) <= layer5_outputs(1372);
    layer6_outputs(914) <= not((layer5_outputs(1774)) or (layer5_outputs(750)));
    layer6_outputs(915) <= layer5_outputs(94);
    layer6_outputs(916) <= not(layer5_outputs(536));
    layer6_outputs(917) <= layer5_outputs(1374);
    layer6_outputs(918) <= layer5_outputs(1431);
    layer6_outputs(919) <= not(layer5_outputs(1257));
    layer6_outputs(920) <= layer5_outputs(307);
    layer6_outputs(921) <= (layer5_outputs(1914)) and not (layer5_outputs(953));
    layer6_outputs(922) <= layer5_outputs(362);
    layer6_outputs(923) <= layer5_outputs(2365);
    layer6_outputs(924) <= layer5_outputs(527);
    layer6_outputs(925) <= (layer5_outputs(363)) and (layer5_outputs(117));
    layer6_outputs(926) <= not(layer5_outputs(453));
    layer6_outputs(927) <= (layer5_outputs(919)) xor (layer5_outputs(207));
    layer6_outputs(928) <= not(layer5_outputs(2480)) or (layer5_outputs(1325));
    layer6_outputs(929) <= not((layer5_outputs(1222)) xor (layer5_outputs(1456)));
    layer6_outputs(930) <= not(layer5_outputs(894)) or (layer5_outputs(1263));
    layer6_outputs(931) <= not(layer5_outputs(2436));
    layer6_outputs(932) <= layer5_outputs(2070);
    layer6_outputs(933) <= layer5_outputs(1729);
    layer6_outputs(934) <= (layer5_outputs(2517)) or (layer5_outputs(105));
    layer6_outputs(935) <= not(layer5_outputs(705));
    layer6_outputs(936) <= layer5_outputs(1720);
    layer6_outputs(937) <= not((layer5_outputs(2288)) xor (layer5_outputs(618)));
    layer6_outputs(938) <= layer5_outputs(62);
    layer6_outputs(939) <= not((layer5_outputs(1835)) xor (layer5_outputs(932)));
    layer6_outputs(940) <= not(layer5_outputs(2496));
    layer6_outputs(941) <= not((layer5_outputs(1236)) xor (layer5_outputs(1779)));
    layer6_outputs(942) <= (layer5_outputs(11)) xor (layer5_outputs(33));
    layer6_outputs(943) <= not((layer5_outputs(1946)) or (layer5_outputs(910)));
    layer6_outputs(944) <= layer5_outputs(127);
    layer6_outputs(945) <= not(layer5_outputs(934)) or (layer5_outputs(2497));
    layer6_outputs(946) <= not(layer5_outputs(354));
    layer6_outputs(947) <= layer5_outputs(594);
    layer6_outputs(948) <= not(layer5_outputs(1894));
    layer6_outputs(949) <= not(layer5_outputs(1867));
    layer6_outputs(950) <= (layer5_outputs(1263)) or (layer5_outputs(1988));
    layer6_outputs(951) <= layer5_outputs(2007);
    layer6_outputs(952) <= (layer5_outputs(1297)) and not (layer5_outputs(1492));
    layer6_outputs(953) <= (layer5_outputs(2396)) xor (layer5_outputs(2342));
    layer6_outputs(954) <= not(layer5_outputs(2162));
    layer6_outputs(955) <= (layer5_outputs(1919)) and not (layer5_outputs(639));
    layer6_outputs(956) <= (layer5_outputs(1245)) or (layer5_outputs(1004));
    layer6_outputs(957) <= layer5_outputs(2420);
    layer6_outputs(958) <= not(layer5_outputs(1668));
    layer6_outputs(959) <= not(layer5_outputs(427));
    layer6_outputs(960) <= (layer5_outputs(1250)) and not (layer5_outputs(2057));
    layer6_outputs(961) <= layer5_outputs(307);
    layer6_outputs(962) <= not(layer5_outputs(840));
    layer6_outputs(963) <= (layer5_outputs(376)) or (layer5_outputs(478));
    layer6_outputs(964) <= not(layer5_outputs(2255));
    layer6_outputs(965) <= not((layer5_outputs(2483)) xor (layer5_outputs(2210)));
    layer6_outputs(966) <= not(layer5_outputs(2253));
    layer6_outputs(967) <= (layer5_outputs(1665)) xor (layer5_outputs(868));
    layer6_outputs(968) <= (layer5_outputs(735)) xor (layer5_outputs(1087));
    layer6_outputs(969) <= (layer5_outputs(538)) and not (layer5_outputs(1123));
    layer6_outputs(970) <= (layer5_outputs(397)) and (layer5_outputs(1758));
    layer6_outputs(971) <= (layer5_outputs(2404)) and not (layer5_outputs(1876));
    layer6_outputs(972) <= not(layer5_outputs(1874));
    layer6_outputs(973) <= not(layer5_outputs(97));
    layer6_outputs(974) <= (layer5_outputs(71)) and not (layer5_outputs(1341));
    layer6_outputs(975) <= not(layer5_outputs(1194));
    layer6_outputs(976) <= not((layer5_outputs(1147)) or (layer5_outputs(1177)));
    layer6_outputs(977) <= not((layer5_outputs(1878)) xor (layer5_outputs(2194)));
    layer6_outputs(978) <= not(layer5_outputs(920));
    layer6_outputs(979) <= not(layer5_outputs(2417));
    layer6_outputs(980) <= not((layer5_outputs(190)) and (layer5_outputs(251)));
    layer6_outputs(981) <= layer5_outputs(1447);
    layer6_outputs(982) <= (layer5_outputs(1568)) and (layer5_outputs(2112));
    layer6_outputs(983) <= not((layer5_outputs(1710)) or (layer5_outputs(1416)));
    layer6_outputs(984) <= not((layer5_outputs(2123)) xor (layer5_outputs(2414)));
    layer6_outputs(985) <= not((layer5_outputs(2150)) or (layer5_outputs(1883)));
    layer6_outputs(986) <= (layer5_outputs(583)) and (layer5_outputs(1577));
    layer6_outputs(987) <= not(layer5_outputs(1163));
    layer6_outputs(988) <= layer5_outputs(646);
    layer6_outputs(989) <= not(layer5_outputs(1707));
    layer6_outputs(990) <= layer5_outputs(65);
    layer6_outputs(991) <= (layer5_outputs(706)) and not (layer5_outputs(318));
    layer6_outputs(992) <= layer5_outputs(493);
    layer6_outputs(993) <= (layer5_outputs(1339)) and not (layer5_outputs(1961));
    layer6_outputs(994) <= (layer5_outputs(1664)) and not (layer5_outputs(1957));
    layer6_outputs(995) <= layer5_outputs(1745);
    layer6_outputs(996) <= layer5_outputs(299);
    layer6_outputs(997) <= layer5_outputs(172);
    layer6_outputs(998) <= not((layer5_outputs(2039)) or (layer5_outputs(1372)));
    layer6_outputs(999) <= not(layer5_outputs(1077));
    layer6_outputs(1000) <= not(layer5_outputs(1361));
    layer6_outputs(1001) <= (layer5_outputs(705)) or (layer5_outputs(860));
    layer6_outputs(1002) <= (layer5_outputs(384)) and not (layer5_outputs(637));
    layer6_outputs(1003) <= layer5_outputs(1548);
    layer6_outputs(1004) <= (layer5_outputs(1329)) and (layer5_outputs(275));
    layer6_outputs(1005) <= not(layer5_outputs(857));
    layer6_outputs(1006) <= (layer5_outputs(1304)) and (layer5_outputs(2196));
    layer6_outputs(1007) <= not((layer5_outputs(1197)) or (layer5_outputs(1627)));
    layer6_outputs(1008) <= (layer5_outputs(1148)) and not (layer5_outputs(2553));
    layer6_outputs(1009) <= not(layer5_outputs(2301));
    layer6_outputs(1010) <= not(layer5_outputs(1918));
    layer6_outputs(1011) <= not(layer5_outputs(2050));
    layer6_outputs(1012) <= not(layer5_outputs(2250));
    layer6_outputs(1013) <= not(layer5_outputs(2400));
    layer6_outputs(1014) <= layer5_outputs(1962);
    layer6_outputs(1015) <= layer5_outputs(867);
    layer6_outputs(1016) <= (layer5_outputs(939)) and (layer5_outputs(224));
    layer6_outputs(1017) <= '0';
    layer6_outputs(1018) <= layer5_outputs(2214);
    layer6_outputs(1019) <= not(layer5_outputs(1610)) or (layer5_outputs(574));
    layer6_outputs(1020) <= (layer5_outputs(1624)) or (layer5_outputs(1350));
    layer6_outputs(1021) <= layer5_outputs(1193);
    layer6_outputs(1022) <= layer5_outputs(1166);
    layer6_outputs(1023) <= (layer5_outputs(2289)) or (layer5_outputs(31));
    layer6_outputs(1024) <= (layer5_outputs(1054)) and not (layer5_outputs(309));
    layer6_outputs(1025) <= (layer5_outputs(585)) and not (layer5_outputs(1618));
    layer6_outputs(1026) <= not((layer5_outputs(2202)) xor (layer5_outputs(650)));
    layer6_outputs(1027) <= (layer5_outputs(1242)) xor (layer5_outputs(25));
    layer6_outputs(1028) <= (layer5_outputs(12)) and not (layer5_outputs(283));
    layer6_outputs(1029) <= not((layer5_outputs(1491)) or (layer5_outputs(290)));
    layer6_outputs(1030) <= not(layer5_outputs(110)) or (layer5_outputs(445));
    layer6_outputs(1031) <= not((layer5_outputs(2538)) xor (layer5_outputs(1062)));
    layer6_outputs(1032) <= layer5_outputs(1078);
    layer6_outputs(1033) <= not((layer5_outputs(942)) or (layer5_outputs(1891)));
    layer6_outputs(1034) <= not((layer5_outputs(2467)) or (layer5_outputs(202)));
    layer6_outputs(1035) <= not((layer5_outputs(1812)) or (layer5_outputs(2094)));
    layer6_outputs(1036) <= layer5_outputs(1111);
    layer6_outputs(1037) <= not(layer5_outputs(2419)) or (layer5_outputs(257));
    layer6_outputs(1038) <= not(layer5_outputs(2371));
    layer6_outputs(1039) <= (layer5_outputs(1614)) xor (layer5_outputs(2557));
    layer6_outputs(1040) <= not((layer5_outputs(68)) or (layer5_outputs(800)));
    layer6_outputs(1041) <= (layer5_outputs(147)) and (layer5_outputs(2419));
    layer6_outputs(1042) <= layer5_outputs(1810);
    layer6_outputs(1043) <= not(layer5_outputs(1204)) or (layer5_outputs(148));
    layer6_outputs(1044) <= not((layer5_outputs(406)) and (layer5_outputs(1823)));
    layer6_outputs(1045) <= not(layer5_outputs(1599));
    layer6_outputs(1046) <= layer5_outputs(998);
    layer6_outputs(1047) <= not(layer5_outputs(2249));
    layer6_outputs(1048) <= not(layer5_outputs(2177)) or (layer5_outputs(745));
    layer6_outputs(1049) <= not(layer5_outputs(2098));
    layer6_outputs(1050) <= '0';
    layer6_outputs(1051) <= layer5_outputs(1476);
    layer6_outputs(1052) <= not((layer5_outputs(959)) and (layer5_outputs(1024)));
    layer6_outputs(1053) <= (layer5_outputs(73)) and not (layer5_outputs(2137));
    layer6_outputs(1054) <= not(layer5_outputs(2128));
    layer6_outputs(1055) <= (layer5_outputs(2023)) and not (layer5_outputs(403));
    layer6_outputs(1056) <= layer5_outputs(1578);
    layer6_outputs(1057) <= not((layer5_outputs(1076)) or (layer5_outputs(1663)));
    layer6_outputs(1058) <= (layer5_outputs(698)) or (layer5_outputs(349));
    layer6_outputs(1059) <= layer5_outputs(152);
    layer6_outputs(1060) <= not(layer5_outputs(908));
    layer6_outputs(1061) <= not((layer5_outputs(881)) xor (layer5_outputs(1519)));
    layer6_outputs(1062) <= not((layer5_outputs(764)) or (layer5_outputs(194)));
    layer6_outputs(1063) <= layer5_outputs(2345);
    layer6_outputs(1064) <= (layer5_outputs(102)) and (layer5_outputs(1031));
    layer6_outputs(1065) <= not(layer5_outputs(264));
    layer6_outputs(1066) <= layer5_outputs(58);
    layer6_outputs(1067) <= not(layer5_outputs(2099));
    layer6_outputs(1068) <= (layer5_outputs(2461)) xor (layer5_outputs(6));
    layer6_outputs(1069) <= (layer5_outputs(2443)) and not (layer5_outputs(2361));
    layer6_outputs(1070) <= layer5_outputs(86);
    layer6_outputs(1071) <= not(layer5_outputs(1941)) or (layer5_outputs(0));
    layer6_outputs(1072) <= (layer5_outputs(1995)) xor (layer5_outputs(2022));
    layer6_outputs(1073) <= not(layer5_outputs(1341));
    layer6_outputs(1074) <= not(layer5_outputs(1841));
    layer6_outputs(1075) <= layer5_outputs(1177);
    layer6_outputs(1076) <= not(layer5_outputs(510));
    layer6_outputs(1077) <= layer5_outputs(675);
    layer6_outputs(1078) <= not(layer5_outputs(2241));
    layer6_outputs(1079) <= layer5_outputs(571);
    layer6_outputs(1080) <= layer5_outputs(559);
    layer6_outputs(1081) <= layer5_outputs(542);
    layer6_outputs(1082) <= not(layer5_outputs(346));
    layer6_outputs(1083) <= not(layer5_outputs(2531)) or (layer5_outputs(857));
    layer6_outputs(1084) <= not((layer5_outputs(1105)) and (layer5_outputs(1018)));
    layer6_outputs(1085) <= not(layer5_outputs(1379)) or (layer5_outputs(214));
    layer6_outputs(1086) <= (layer5_outputs(1081)) or (layer5_outputs(435));
    layer6_outputs(1087) <= not(layer5_outputs(651));
    layer6_outputs(1088) <= layer5_outputs(502);
    layer6_outputs(1089) <= layer5_outputs(1297);
    layer6_outputs(1090) <= not(layer5_outputs(2505)) or (layer5_outputs(1755));
    layer6_outputs(1091) <= layer5_outputs(954);
    layer6_outputs(1092) <= (layer5_outputs(1865)) and (layer5_outputs(2192));
    layer6_outputs(1093) <= layer5_outputs(2301);
    layer6_outputs(1094) <= (layer5_outputs(1781)) xor (layer5_outputs(1130));
    layer6_outputs(1095) <= not(layer5_outputs(2019));
    layer6_outputs(1096) <= not(layer5_outputs(2360));
    layer6_outputs(1097) <= layer5_outputs(1303);
    layer6_outputs(1098) <= not((layer5_outputs(2187)) or (layer5_outputs(1094)));
    layer6_outputs(1099) <= (layer5_outputs(1080)) and not (layer5_outputs(1019));
    layer6_outputs(1100) <= not(layer5_outputs(832));
    layer6_outputs(1101) <= not((layer5_outputs(692)) and (layer5_outputs(1612)));
    layer6_outputs(1102) <= (layer5_outputs(404)) xor (layer5_outputs(1306));
    layer6_outputs(1103) <= not(layer5_outputs(2168)) or (layer5_outputs(236));
    layer6_outputs(1104) <= (layer5_outputs(1589)) and not (layer5_outputs(1155));
    layer6_outputs(1105) <= not(layer5_outputs(711)) or (layer5_outputs(334));
    layer6_outputs(1106) <= not((layer5_outputs(1720)) and (layer5_outputs(308)));
    layer6_outputs(1107) <= layer5_outputs(1555);
    layer6_outputs(1108) <= (layer5_outputs(2144)) and not (layer5_outputs(79));
    layer6_outputs(1109) <= (layer5_outputs(783)) and (layer5_outputs(1252));
    layer6_outputs(1110) <= not(layer5_outputs(1153));
    layer6_outputs(1111) <= not(layer5_outputs(605));
    layer6_outputs(1112) <= layer5_outputs(331);
    layer6_outputs(1113) <= not(layer5_outputs(2221));
    layer6_outputs(1114) <= layer5_outputs(2185);
    layer6_outputs(1115) <= not(layer5_outputs(277));
    layer6_outputs(1116) <= not(layer5_outputs(420));
    layer6_outputs(1117) <= layer5_outputs(1244);
    layer6_outputs(1118) <= not(layer5_outputs(2354));
    layer6_outputs(1119) <= not(layer5_outputs(1234));
    layer6_outputs(1120) <= not(layer5_outputs(454));
    layer6_outputs(1121) <= not(layer5_outputs(154));
    layer6_outputs(1122) <= (layer5_outputs(1222)) and not (layer5_outputs(2021));
    layer6_outputs(1123) <= not((layer5_outputs(2406)) or (layer5_outputs(605)));
    layer6_outputs(1124) <= layer5_outputs(1469);
    layer6_outputs(1125) <= not(layer5_outputs(1538));
    layer6_outputs(1126) <= (layer5_outputs(957)) and (layer5_outputs(237));
    layer6_outputs(1127) <= (layer5_outputs(2228)) and (layer5_outputs(1673));
    layer6_outputs(1128) <= (layer5_outputs(1531)) xor (layer5_outputs(1798));
    layer6_outputs(1129) <= not(layer5_outputs(1747));
    layer6_outputs(1130) <= not(layer5_outputs(1654));
    layer6_outputs(1131) <= layer5_outputs(2180);
    layer6_outputs(1132) <= layer5_outputs(756);
    layer6_outputs(1133) <= (layer5_outputs(581)) and not (layer5_outputs(1837));
    layer6_outputs(1134) <= (layer5_outputs(325)) and (layer5_outputs(1496));
    layer6_outputs(1135) <= not(layer5_outputs(2271));
    layer6_outputs(1136) <= not((layer5_outputs(892)) xor (layer5_outputs(507)));
    layer6_outputs(1137) <= not((layer5_outputs(67)) or (layer5_outputs(1361)));
    layer6_outputs(1138) <= not(layer5_outputs(2414));
    layer6_outputs(1139) <= layer5_outputs(351);
    layer6_outputs(1140) <= not(layer5_outputs(178));
    layer6_outputs(1141) <= not(layer5_outputs(2436));
    layer6_outputs(1142) <= not((layer5_outputs(1312)) xor (layer5_outputs(121)));
    layer6_outputs(1143) <= not(layer5_outputs(1350));
    layer6_outputs(1144) <= not((layer5_outputs(2066)) xor (layer5_outputs(2165)));
    layer6_outputs(1145) <= not(layer5_outputs(1929));
    layer6_outputs(1146) <= not(layer5_outputs(1477)) or (layer5_outputs(1234));
    layer6_outputs(1147) <= not(layer5_outputs(966));
    layer6_outputs(1148) <= not((layer5_outputs(960)) and (layer5_outputs(2240)));
    layer6_outputs(1149) <= (layer5_outputs(1300)) xor (layer5_outputs(369));
    layer6_outputs(1150) <= layer5_outputs(1485);
    layer6_outputs(1151) <= (layer5_outputs(2377)) and not (layer5_outputs(1803));
    layer6_outputs(1152) <= '0';
    layer6_outputs(1153) <= not(layer5_outputs(2520));
    layer6_outputs(1154) <= not(layer5_outputs(811)) or (layer5_outputs(72));
    layer6_outputs(1155) <= layer5_outputs(143);
    layer6_outputs(1156) <= not((layer5_outputs(2272)) xor (layer5_outputs(2085)));
    layer6_outputs(1157) <= (layer5_outputs(1861)) xor (layer5_outputs(862));
    layer6_outputs(1158) <= layer5_outputs(914);
    layer6_outputs(1159) <= not(layer5_outputs(702));
    layer6_outputs(1160) <= layer5_outputs(1120);
    layer6_outputs(1161) <= not(layer5_outputs(213));
    layer6_outputs(1162) <= layer5_outputs(629);
    layer6_outputs(1163) <= (layer5_outputs(2030)) or (layer5_outputs(1283));
    layer6_outputs(1164) <= (layer5_outputs(2322)) xor (layer5_outputs(971));
    layer6_outputs(1165) <= (layer5_outputs(1188)) and (layer5_outputs(20));
    layer6_outputs(1166) <= (layer5_outputs(1473)) and not (layer5_outputs(1641));
    layer6_outputs(1167) <= not((layer5_outputs(456)) xor (layer5_outputs(1458)));
    layer6_outputs(1168) <= layer5_outputs(1065);
    layer6_outputs(1169) <= layer5_outputs(842);
    layer6_outputs(1170) <= layer5_outputs(544);
    layer6_outputs(1171) <= layer5_outputs(881);
    layer6_outputs(1172) <= layer5_outputs(2052);
    layer6_outputs(1173) <= not(layer5_outputs(2032)) or (layer5_outputs(554));
    layer6_outputs(1174) <= (layer5_outputs(960)) and not (layer5_outputs(2141));
    layer6_outputs(1175) <= not(layer5_outputs(1564));
    layer6_outputs(1176) <= not((layer5_outputs(1637)) or (layer5_outputs(1066)));
    layer6_outputs(1177) <= (layer5_outputs(1895)) xor (layer5_outputs(1268));
    layer6_outputs(1178) <= layer5_outputs(2529);
    layer6_outputs(1179) <= layer5_outputs(84);
    layer6_outputs(1180) <= layer5_outputs(850);
    layer6_outputs(1181) <= not(layer5_outputs(1446)) or (layer5_outputs(1398));
    layer6_outputs(1182) <= not(layer5_outputs(660)) or (layer5_outputs(141));
    layer6_outputs(1183) <= layer5_outputs(621);
    layer6_outputs(1184) <= not((layer5_outputs(855)) and (layer5_outputs(2421)));
    layer6_outputs(1185) <= not(layer5_outputs(751));
    layer6_outputs(1186) <= layer5_outputs(2470);
    layer6_outputs(1187) <= not(layer5_outputs(1067));
    layer6_outputs(1188) <= not(layer5_outputs(200));
    layer6_outputs(1189) <= '0';
    layer6_outputs(1190) <= (layer5_outputs(1412)) and not (layer5_outputs(323));
    layer6_outputs(1191) <= not((layer5_outputs(1213)) xor (layer5_outputs(1695)));
    layer6_outputs(1192) <= not(layer5_outputs(1474));
    layer6_outputs(1193) <= layer5_outputs(1313);
    layer6_outputs(1194) <= not((layer5_outputs(244)) and (layer5_outputs(2430)));
    layer6_outputs(1195) <= not(layer5_outputs(2207));
    layer6_outputs(1196) <= (layer5_outputs(968)) xor (layer5_outputs(276));
    layer6_outputs(1197) <= not(layer5_outputs(1149)) or (layer5_outputs(2305));
    layer6_outputs(1198) <= (layer5_outputs(2329)) and not (layer5_outputs(1367));
    layer6_outputs(1199) <= layer5_outputs(254);
    layer6_outputs(1200) <= not((layer5_outputs(676)) xor (layer5_outputs(2214)));
    layer6_outputs(1201) <= (layer5_outputs(2170)) xor (layer5_outputs(2304));
    layer6_outputs(1202) <= layer5_outputs(1766);
    layer6_outputs(1203) <= layer5_outputs(769);
    layer6_outputs(1204) <= not(layer5_outputs(298));
    layer6_outputs(1205) <= (layer5_outputs(748)) xor (layer5_outputs(419));
    layer6_outputs(1206) <= layer5_outputs(1857);
    layer6_outputs(1207) <= not(layer5_outputs(157));
    layer6_outputs(1208) <= (layer5_outputs(2129)) xor (layer5_outputs(1128));
    layer6_outputs(1209) <= not(layer5_outputs(2500)) or (layer5_outputs(1512));
    layer6_outputs(1210) <= (layer5_outputs(2223)) and not (layer5_outputs(933));
    layer6_outputs(1211) <= not(layer5_outputs(2016));
    layer6_outputs(1212) <= not(layer5_outputs(332)) or (layer5_outputs(2121));
    layer6_outputs(1213) <= not(layer5_outputs(1243));
    layer6_outputs(1214) <= (layer5_outputs(2116)) and not (layer5_outputs(572));
    layer6_outputs(1215) <= not((layer5_outputs(1060)) xor (layer5_outputs(595)));
    layer6_outputs(1216) <= not(layer5_outputs(1583));
    layer6_outputs(1217) <= (layer5_outputs(600)) and not (layer5_outputs(996));
    layer6_outputs(1218) <= not(layer5_outputs(373));
    layer6_outputs(1219) <= (layer5_outputs(921)) or (layer5_outputs(1276));
    layer6_outputs(1220) <= not((layer5_outputs(390)) or (layer5_outputs(820)));
    layer6_outputs(1221) <= not((layer5_outputs(1732)) and (layer5_outputs(1686)));
    layer6_outputs(1222) <= (layer5_outputs(938)) xor (layer5_outputs(2359));
    layer6_outputs(1223) <= not(layer5_outputs(1036)) or (layer5_outputs(407));
    layer6_outputs(1224) <= (layer5_outputs(2131)) and (layer5_outputs(2363));
    layer6_outputs(1225) <= not(layer5_outputs(324)) or (layer5_outputs(1803));
    layer6_outputs(1226) <= layer5_outputs(424);
    layer6_outputs(1227) <= layer5_outputs(816);
    layer6_outputs(1228) <= (layer5_outputs(119)) xor (layer5_outputs(40));
    layer6_outputs(1229) <= not(layer5_outputs(2070));
    layer6_outputs(1230) <= (layer5_outputs(501)) and not (layer5_outputs(502));
    layer6_outputs(1231) <= (layer5_outputs(485)) or (layer5_outputs(1102));
    layer6_outputs(1232) <= not((layer5_outputs(2143)) or (layer5_outputs(2506)));
    layer6_outputs(1233) <= (layer5_outputs(987)) and not (layer5_outputs(482));
    layer6_outputs(1234) <= not((layer5_outputs(1514)) and (layer5_outputs(825)));
    layer6_outputs(1235) <= not((layer5_outputs(1586)) xor (layer5_outputs(1116)));
    layer6_outputs(1236) <= (layer5_outputs(1636)) xor (layer5_outputs(602));
    layer6_outputs(1237) <= layer5_outputs(304);
    layer6_outputs(1238) <= (layer5_outputs(289)) or (layer5_outputs(2203));
    layer6_outputs(1239) <= (layer5_outputs(52)) and not (layer5_outputs(1108));
    layer6_outputs(1240) <= (layer5_outputs(716)) and not (layer5_outputs(1201));
    layer6_outputs(1241) <= not((layer5_outputs(319)) or (layer5_outputs(2017)));
    layer6_outputs(1242) <= '0';
    layer6_outputs(1243) <= layer5_outputs(664);
    layer6_outputs(1244) <= not(layer5_outputs(1071));
    layer6_outputs(1245) <= (layer5_outputs(848)) and not (layer5_outputs(400));
    layer6_outputs(1246) <= (layer5_outputs(43)) and not (layer5_outputs(2242));
    layer6_outputs(1247) <= (layer5_outputs(1834)) and not (layer5_outputs(2380));
    layer6_outputs(1248) <= not(layer5_outputs(459)) or (layer5_outputs(940));
    layer6_outputs(1249) <= not(layer5_outputs(1948));
    layer6_outputs(1250) <= (layer5_outputs(2498)) and (layer5_outputs(1069));
    layer6_outputs(1251) <= not((layer5_outputs(1279)) and (layer5_outputs(1271)));
    layer6_outputs(1252) <= (layer5_outputs(214)) xor (layer5_outputs(199));
    layer6_outputs(1253) <= not(layer5_outputs(417));
    layer6_outputs(1254) <= not(layer5_outputs(2448));
    layer6_outputs(1255) <= (layer5_outputs(1472)) and (layer5_outputs(2096));
    layer6_outputs(1256) <= layer5_outputs(2383);
    layer6_outputs(1257) <= not(layer5_outputs(2442)) or (layer5_outputs(1402));
    layer6_outputs(1258) <= not(layer5_outputs(2415));
    layer6_outputs(1259) <= '1';
    layer6_outputs(1260) <= (layer5_outputs(661)) and not (layer5_outputs(1581));
    layer6_outputs(1261) <= not(layer5_outputs(544)) or (layer5_outputs(733));
    layer6_outputs(1262) <= not(layer5_outputs(1526));
    layer6_outputs(1263) <= not(layer5_outputs(222)) or (layer5_outputs(1118));
    layer6_outputs(1264) <= not(layer5_outputs(1407)) or (layer5_outputs(1976));
    layer6_outputs(1265) <= layer5_outputs(40);
    layer6_outputs(1266) <= layer5_outputs(270);
    layer6_outputs(1267) <= not(layer5_outputs(482));
    layer6_outputs(1268) <= (layer5_outputs(473)) and (layer5_outputs(2537));
    layer6_outputs(1269) <= not(layer5_outputs(1246));
    layer6_outputs(1270) <= not(layer5_outputs(2082)) or (layer5_outputs(1782));
    layer6_outputs(1271) <= layer5_outputs(806);
    layer6_outputs(1272) <= layer5_outputs(1083);
    layer6_outputs(1273) <= layer5_outputs(60);
    layer6_outputs(1274) <= layer5_outputs(1923);
    layer6_outputs(1275) <= not(layer5_outputs(1666)) or (layer5_outputs(995));
    layer6_outputs(1276) <= not(layer5_outputs(2351));
    layer6_outputs(1277) <= not((layer5_outputs(921)) and (layer5_outputs(267)));
    layer6_outputs(1278) <= (layer5_outputs(891)) xor (layer5_outputs(321));
    layer6_outputs(1279) <= not((layer5_outputs(979)) xor (layer5_outputs(74)));
    layer6_outputs(1280) <= not(layer5_outputs(417));
    layer6_outputs(1281) <= (layer5_outputs(1358)) xor (layer5_outputs(513));
    layer6_outputs(1282) <= (layer5_outputs(1748)) and (layer5_outputs(1186));
    layer6_outputs(1283) <= layer5_outputs(296);
    layer6_outputs(1284) <= not(layer5_outputs(985)) or (layer5_outputs(2485));
    layer6_outputs(1285) <= (layer5_outputs(2371)) and not (layer5_outputs(2422));
    layer6_outputs(1286) <= not(layer5_outputs(443));
    layer6_outputs(1287) <= not(layer5_outputs(1915));
    layer6_outputs(1288) <= not(layer5_outputs(1371));
    layer6_outputs(1289) <= not(layer5_outputs(883));
    layer6_outputs(1290) <= (layer5_outputs(612)) and (layer5_outputs(182));
    layer6_outputs(1291) <= not(layer5_outputs(350)) or (layer5_outputs(483));
    layer6_outputs(1292) <= (layer5_outputs(640)) and not (layer5_outputs(2554));
    layer6_outputs(1293) <= layer5_outputs(980);
    layer6_outputs(1294) <= layer5_outputs(1159);
    layer6_outputs(1295) <= not((layer5_outputs(2453)) xor (layer5_outputs(140)));
    layer6_outputs(1296) <= not((layer5_outputs(2325)) and (layer5_outputs(733)));
    layer6_outputs(1297) <= not(layer5_outputs(1838)) or (layer5_outputs(1632));
    layer6_outputs(1298) <= not((layer5_outputs(10)) xor (layer5_outputs(2482)));
    layer6_outputs(1299) <= layer5_outputs(2100);
    layer6_outputs(1300) <= layer5_outputs(1602);
    layer6_outputs(1301) <= layer5_outputs(2106);
    layer6_outputs(1302) <= not((layer5_outputs(2026)) xor (layer5_outputs(2310)));
    layer6_outputs(1303) <= not(layer5_outputs(835));
    layer6_outputs(1304) <= not(layer5_outputs(2518));
    layer6_outputs(1305) <= (layer5_outputs(1651)) xor (layer5_outputs(1005));
    layer6_outputs(1306) <= layer5_outputs(993);
    layer6_outputs(1307) <= not((layer5_outputs(1463)) xor (layer5_outputs(76)));
    layer6_outputs(1308) <= layer5_outputs(28);
    layer6_outputs(1309) <= (layer5_outputs(1318)) or (layer5_outputs(1788));
    layer6_outputs(1310) <= layer5_outputs(2455);
    layer6_outputs(1311) <= '0';
    layer6_outputs(1312) <= not(layer5_outputs(606));
    layer6_outputs(1313) <= not(layer5_outputs(2350));
    layer6_outputs(1314) <= (layer5_outputs(1445)) and not (layer5_outputs(2051));
    layer6_outputs(1315) <= layer5_outputs(2136);
    layer6_outputs(1316) <= not((layer5_outputs(1268)) and (layer5_outputs(35)));
    layer6_outputs(1317) <= not((layer5_outputs(2204)) and (layer5_outputs(26)));
    layer6_outputs(1318) <= not(layer5_outputs(1942));
    layer6_outputs(1319) <= layer5_outputs(1048);
    layer6_outputs(1320) <= not(layer5_outputs(1707));
    layer6_outputs(1321) <= not(layer5_outputs(218));
    layer6_outputs(1322) <= not(layer5_outputs(1905)) or (layer5_outputs(530));
    layer6_outputs(1323) <= not(layer5_outputs(984)) or (layer5_outputs(1187));
    layer6_outputs(1324) <= (layer5_outputs(1783)) and (layer5_outputs(1195));
    layer6_outputs(1325) <= (layer5_outputs(2055)) and not (layer5_outputs(1212));
    layer6_outputs(1326) <= (layer5_outputs(508)) and not (layer5_outputs(2106));
    layer6_outputs(1327) <= layer5_outputs(1006);
    layer6_outputs(1328) <= not((layer5_outputs(2512)) xor (layer5_outputs(2556)));
    layer6_outputs(1329) <= not((layer5_outputs(870)) xor (layer5_outputs(1038)));
    layer6_outputs(1330) <= (layer5_outputs(41)) and (layer5_outputs(1197));
    layer6_outputs(1331) <= not((layer5_outputs(75)) and (layer5_outputs(1327)));
    layer6_outputs(1332) <= (layer5_outputs(2348)) xor (layer5_outputs(78));
    layer6_outputs(1333) <= (layer5_outputs(1423)) and not (layer5_outputs(609));
    layer6_outputs(1334) <= not(layer5_outputs(2463));
    layer6_outputs(1335) <= (layer5_outputs(118)) xor (layer5_outputs(1776));
    layer6_outputs(1336) <= not(layer5_outputs(2060));
    layer6_outputs(1337) <= not((layer5_outputs(472)) and (layer5_outputs(740)));
    layer6_outputs(1338) <= not(layer5_outputs(136));
    layer6_outputs(1339) <= layer5_outputs(1806);
    layer6_outputs(1340) <= (layer5_outputs(884)) and not (layer5_outputs(2238));
    layer6_outputs(1341) <= not(layer5_outputs(398));
    layer6_outputs(1342) <= not(layer5_outputs(1678));
    layer6_outputs(1343) <= (layer5_outputs(2334)) and not (layer5_outputs(1614));
    layer6_outputs(1344) <= layer5_outputs(599);
    layer6_outputs(1345) <= not((layer5_outputs(676)) xor (layer5_outputs(1584)));
    layer6_outputs(1346) <= '0';
    layer6_outputs(1347) <= layer5_outputs(547);
    layer6_outputs(1348) <= layer5_outputs(1253);
    layer6_outputs(1349) <= (layer5_outputs(2303)) and not (layer5_outputs(701));
    layer6_outputs(1350) <= layer5_outputs(851);
    layer6_outputs(1351) <= (layer5_outputs(1601)) and (layer5_outputs(1717));
    layer6_outputs(1352) <= layer5_outputs(682);
    layer6_outputs(1353) <= not(layer5_outputs(1649));
    layer6_outputs(1354) <= layer5_outputs(1401);
    layer6_outputs(1355) <= not(layer5_outputs(2444));
    layer6_outputs(1356) <= not(layer5_outputs(261)) or (layer5_outputs(832));
    layer6_outputs(1357) <= not(layer5_outputs(1075));
    layer6_outputs(1358) <= (layer5_outputs(1691)) and not (layer5_outputs(2188));
    layer6_outputs(1359) <= not(layer5_outputs(317)) or (layer5_outputs(937));
    layer6_outputs(1360) <= not(layer5_outputs(999));
    layer6_outputs(1361) <= layer5_outputs(1454);
    layer6_outputs(1362) <= '0';
    layer6_outputs(1363) <= layer5_outputs(2167);
    layer6_outputs(1364) <= not(layer5_outputs(1646));
    layer6_outputs(1365) <= layer5_outputs(2061);
    layer6_outputs(1366) <= '1';
    layer6_outputs(1367) <= (layer5_outputs(1905)) and not (layer5_outputs(549));
    layer6_outputs(1368) <= not(layer5_outputs(905));
    layer6_outputs(1369) <= layer5_outputs(208);
    layer6_outputs(1370) <= not((layer5_outputs(1971)) xor (layer5_outputs(1404)));
    layer6_outputs(1371) <= (layer5_outputs(1764)) xor (layer5_outputs(2357));
    layer6_outputs(1372) <= not(layer5_outputs(1544)) or (layer5_outputs(1289));
    layer6_outputs(1373) <= layer5_outputs(2172);
    layer6_outputs(1374) <= layer5_outputs(794);
    layer6_outputs(1375) <= not(layer5_outputs(2549));
    layer6_outputs(1376) <= not(layer5_outputs(2134)) or (layer5_outputs(406));
    layer6_outputs(1377) <= not(layer5_outputs(2059));
    layer6_outputs(1378) <= not(layer5_outputs(2265));
    layer6_outputs(1379) <= (layer5_outputs(1872)) and not (layer5_outputs(2027));
    layer6_outputs(1380) <= layer5_outputs(432);
    layer6_outputs(1381) <= layer5_outputs(1682);
    layer6_outputs(1382) <= not(layer5_outputs(655));
    layer6_outputs(1383) <= not(layer5_outputs(791));
    layer6_outputs(1384) <= layer5_outputs(314);
    layer6_outputs(1385) <= (layer5_outputs(287)) and not (layer5_outputs(1134));
    layer6_outputs(1386) <= not((layer5_outputs(2364)) and (layer5_outputs(212)));
    layer6_outputs(1387) <= not(layer5_outputs(813));
    layer6_outputs(1388) <= layer5_outputs(1604);
    layer6_outputs(1389) <= not((layer5_outputs(286)) and (layer5_outputs(389)));
    layer6_outputs(1390) <= not(layer5_outputs(1206));
    layer6_outputs(1391) <= (layer5_outputs(2369)) xor (layer5_outputs(817));
    layer6_outputs(1392) <= not(layer5_outputs(491));
    layer6_outputs(1393) <= not(layer5_outputs(385));
    layer6_outputs(1394) <= layer5_outputs(1349);
    layer6_outputs(1395) <= not((layer5_outputs(1232)) xor (layer5_outputs(23)));
    layer6_outputs(1396) <= not(layer5_outputs(2532));
    layer6_outputs(1397) <= (layer5_outputs(497)) and not (layer5_outputs(2458));
    layer6_outputs(1398) <= layer5_outputs(1532);
    layer6_outputs(1399) <= (layer5_outputs(326)) and not (layer5_outputs(2170));
    layer6_outputs(1400) <= (layer5_outputs(732)) xor (layer5_outputs(1675));
    layer6_outputs(1401) <= layer5_outputs(167);
    layer6_outputs(1402) <= layer5_outputs(120);
    layer6_outputs(1403) <= layer5_outputs(2522);
    layer6_outputs(1404) <= (layer5_outputs(1683)) and (layer5_outputs(1996));
    layer6_outputs(1405) <= (layer5_outputs(1143)) or (layer5_outputs(1775));
    layer6_outputs(1406) <= not((layer5_outputs(804)) xor (layer5_outputs(1397)));
    layer6_outputs(1407) <= not((layer5_outputs(2182)) xor (layer5_outputs(2023)));
    layer6_outputs(1408) <= not(layer5_outputs(902));
    layer6_outputs(1409) <= (layer5_outputs(2176)) and (layer5_outputs(2293));
    layer6_outputs(1410) <= (layer5_outputs(528)) and not (layer5_outputs(1063));
    layer6_outputs(1411) <= not((layer5_outputs(1015)) xor (layer5_outputs(85)));
    layer6_outputs(1412) <= layer5_outputs(1151);
    layer6_outputs(1413) <= not(layer5_outputs(2155));
    layer6_outputs(1414) <= not(layer5_outputs(197)) or (layer5_outputs(890));
    layer6_outputs(1415) <= not(layer5_outputs(899));
    layer6_outputs(1416) <= (layer5_outputs(678)) xor (layer5_outputs(631));
    layer6_outputs(1417) <= (layer5_outputs(1061)) or (layer5_outputs(1127));
    layer6_outputs(1418) <= not(layer5_outputs(1938));
    layer6_outputs(1419) <= (layer5_outputs(1498)) xor (layer5_outputs(2459));
    layer6_outputs(1420) <= (layer5_outputs(1219)) or (layer5_outputs(54));
    layer6_outputs(1421) <= layer5_outputs(1804);
    layer6_outputs(1422) <= not(layer5_outputs(1039)) or (layer5_outputs(2286));
    layer6_outputs(1423) <= not((layer5_outputs(168)) xor (layer5_outputs(1665)));
    layer6_outputs(1424) <= (layer5_outputs(481)) and not (layer5_outputs(1166));
    layer6_outputs(1425) <= (layer5_outputs(1429)) and not (layer5_outputs(1031));
    layer6_outputs(1426) <= layer5_outputs(1746);
    layer6_outputs(1427) <= not(layer5_outputs(773));
    layer6_outputs(1428) <= (layer5_outputs(1447)) or (layer5_outputs(24));
    layer6_outputs(1429) <= not((layer5_outputs(833)) and (layer5_outputs(1041)));
    layer6_outputs(1430) <= (layer5_outputs(2374)) or (layer5_outputs(1879));
    layer6_outputs(1431) <= not((layer5_outputs(1533)) xor (layer5_outputs(1990)));
    layer6_outputs(1432) <= layer5_outputs(2465);
    layer6_outputs(1433) <= layer5_outputs(2243);
    layer6_outputs(1434) <= layer5_outputs(681);
    layer6_outputs(1435) <= not(layer5_outputs(2350));
    layer6_outputs(1436) <= layer5_outputs(428);
    layer6_outputs(1437) <= layer5_outputs(370);
    layer6_outputs(1438) <= (layer5_outputs(2461)) and not (layer5_outputs(1535));
    layer6_outputs(1439) <= not((layer5_outputs(2174)) or (layer5_outputs(205)));
    layer6_outputs(1440) <= (layer5_outputs(99)) xor (layer5_outputs(1091));
    layer6_outputs(1441) <= not(layer5_outputs(1898));
    layer6_outputs(1442) <= layer5_outputs(670);
    layer6_outputs(1443) <= (layer5_outputs(59)) or (layer5_outputs(1717));
    layer6_outputs(1444) <= not((layer5_outputs(2325)) xor (layer5_outputs(206)));
    layer6_outputs(1445) <= layer5_outputs(546);
    layer6_outputs(1446) <= not(layer5_outputs(2239));
    layer6_outputs(1447) <= layer5_outputs(1684);
    layer6_outputs(1448) <= layer5_outputs(1994);
    layer6_outputs(1449) <= not(layer5_outputs(2369));
    layer6_outputs(1450) <= (layer5_outputs(1978)) or (layer5_outputs(2470));
    layer6_outputs(1451) <= not(layer5_outputs(1826));
    layer6_outputs(1452) <= '1';
    layer6_outputs(1453) <= not(layer5_outputs(1565));
    layer6_outputs(1454) <= layer5_outputs(942);
    layer6_outputs(1455) <= (layer5_outputs(1134)) or (layer5_outputs(1825));
    layer6_outputs(1456) <= layer5_outputs(374);
    layer6_outputs(1457) <= layer5_outputs(887);
    layer6_outputs(1458) <= not(layer5_outputs(2544));
    layer6_outputs(1459) <= not(layer5_outputs(1982));
    layer6_outputs(1460) <= not(layer5_outputs(1253));
    layer6_outputs(1461) <= not(layer5_outputs(1228));
    layer6_outputs(1462) <= (layer5_outputs(1921)) xor (layer5_outputs(1506));
    layer6_outputs(1463) <= not((layer5_outputs(535)) or (layer5_outputs(2279)));
    layer6_outputs(1464) <= (layer5_outputs(237)) and not (layer5_outputs(1161));
    layer6_outputs(1465) <= not(layer5_outputs(2554));
    layer6_outputs(1466) <= layer5_outputs(193);
    layer6_outputs(1467) <= not(layer5_outputs(1700));
    layer6_outputs(1468) <= not((layer5_outputs(1388)) or (layer5_outputs(1772)));
    layer6_outputs(1469) <= not(layer5_outputs(1300)) or (layer5_outputs(176));
    layer6_outputs(1470) <= (layer5_outputs(1390)) and not (layer5_outputs(1225));
    layer6_outputs(1471) <= (layer5_outputs(1438)) xor (layer5_outputs(1270));
    layer6_outputs(1472) <= not(layer5_outputs(1751));
    layer6_outputs(1473) <= not((layer5_outputs(784)) and (layer5_outputs(2385)));
    layer6_outputs(1474) <= layer5_outputs(715);
    layer6_outputs(1475) <= layer5_outputs(205);
    layer6_outputs(1476) <= not((layer5_outputs(1342)) xor (layer5_outputs(695)));
    layer6_outputs(1477) <= not((layer5_outputs(1420)) xor (layer5_outputs(2054)));
    layer6_outputs(1478) <= (layer5_outputs(978)) and not (layer5_outputs(66));
    layer6_outputs(1479) <= not(layer5_outputs(2236));
    layer6_outputs(1480) <= not(layer5_outputs(1295));
    layer6_outputs(1481) <= (layer5_outputs(744)) and not (layer5_outputs(325));
    layer6_outputs(1482) <= layer5_outputs(1822);
    layer6_outputs(1483) <= layer5_outputs(1022);
    layer6_outputs(1484) <= not(layer5_outputs(1818));
    layer6_outputs(1485) <= not(layer5_outputs(2372));
    layer6_outputs(1486) <= layer5_outputs(189);
    layer6_outputs(1487) <= not((layer5_outputs(1393)) and (layer5_outputs(1154)));
    layer6_outputs(1488) <= layer5_outputs(270);
    layer6_outputs(1489) <= (layer5_outputs(2142)) and (layer5_outputs(146));
    layer6_outputs(1490) <= layer5_outputs(253);
    layer6_outputs(1491) <= (layer5_outputs(807)) and (layer5_outputs(427));
    layer6_outputs(1492) <= (layer5_outputs(664)) and not (layer5_outputs(988));
    layer6_outputs(1493) <= layer5_outputs(1343);
    layer6_outputs(1494) <= layer5_outputs(2083);
    layer6_outputs(1495) <= layer5_outputs(1749);
    layer6_outputs(1496) <= not(layer5_outputs(446));
    layer6_outputs(1497) <= not(layer5_outputs(2339));
    layer6_outputs(1498) <= (layer5_outputs(1470)) xor (layer5_outputs(1674));
    layer6_outputs(1499) <= layer5_outputs(1191);
    layer6_outputs(1500) <= layer5_outputs(208);
    layer6_outputs(1501) <= layer5_outputs(338);
    layer6_outputs(1502) <= not(layer5_outputs(1957));
    layer6_outputs(1503) <= '1';
    layer6_outputs(1504) <= layer5_outputs(1140);
    layer6_outputs(1505) <= not((layer5_outputs(765)) or (layer5_outputs(1545)));
    layer6_outputs(1506) <= not(layer5_outputs(2344));
    layer6_outputs(1507) <= (layer5_outputs(495)) and not (layer5_outputs(948));
    layer6_outputs(1508) <= not(layer5_outputs(1174)) or (layer5_outputs(1096));
    layer6_outputs(1509) <= layer5_outputs(2041);
    layer6_outputs(1510) <= not(layer5_outputs(1607));
    layer6_outputs(1511) <= not(layer5_outputs(492));
    layer6_outputs(1512) <= not(layer5_outputs(2455));
    layer6_outputs(1513) <= (layer5_outputs(648)) and (layer5_outputs(2223));
    layer6_outputs(1514) <= not(layer5_outputs(1575)) or (layer5_outputs(276));
    layer6_outputs(1515) <= layer5_outputs(1866);
    layer6_outputs(1516) <= not((layer5_outputs(455)) xor (layer5_outputs(622)));
    layer6_outputs(1517) <= not((layer5_outputs(1169)) and (layer5_outputs(198)));
    layer6_outputs(1518) <= not((layer5_outputs(342)) or (layer5_outputs(1425)));
    layer6_outputs(1519) <= not(layer5_outputs(2107));
    layer6_outputs(1520) <= not(layer5_outputs(1323));
    layer6_outputs(1521) <= not(layer5_outputs(2478));
    layer6_outputs(1522) <= layer5_outputs(1791);
    layer6_outputs(1523) <= not((layer5_outputs(1022)) or (layer5_outputs(2163)));
    layer6_outputs(1524) <= (layer5_outputs(2241)) xor (layer5_outputs(335));
    layer6_outputs(1525) <= (layer5_outputs(2025)) and (layer5_outputs(1690));
    layer6_outputs(1526) <= layer5_outputs(149);
    layer6_outputs(1527) <= not(layer5_outputs(1428));
    layer6_outputs(1528) <= layer5_outputs(1809);
    layer6_outputs(1529) <= (layer5_outputs(805)) or (layer5_outputs(1249));
    layer6_outputs(1530) <= (layer5_outputs(1832)) and not (layer5_outputs(57));
    layer6_outputs(1531) <= not(layer5_outputs(2443));
    layer6_outputs(1532) <= (layer5_outputs(2328)) xor (layer5_outputs(209));
    layer6_outputs(1533) <= (layer5_outputs(51)) xor (layer5_outputs(2235));
    layer6_outputs(1534) <= (layer5_outputs(543)) and not (layer5_outputs(2156));
    layer6_outputs(1535) <= not(layer5_outputs(2199));
    layer6_outputs(1536) <= not(layer5_outputs(923));
    layer6_outputs(1537) <= not((layer5_outputs(1950)) xor (layer5_outputs(32)));
    layer6_outputs(1538) <= not(layer5_outputs(969));
    layer6_outputs(1539) <= not(layer5_outputs(1784)) or (layer5_outputs(2447));
    layer6_outputs(1540) <= not(layer5_outputs(1571));
    layer6_outputs(1541) <= layer5_outputs(1274);
    layer6_outputs(1542) <= not(layer5_outputs(1680));
    layer6_outputs(1543) <= (layer5_outputs(135)) and (layer5_outputs(1998));
    layer6_outputs(1544) <= not((layer5_outputs(145)) or (layer5_outputs(253)));
    layer6_outputs(1545) <= not(layer5_outputs(222)) or (layer5_outputs(1442));
    layer6_outputs(1546) <= (layer5_outputs(488)) or (layer5_outputs(451));
    layer6_outputs(1547) <= layer5_outputs(503);
    layer6_outputs(1548) <= layer5_outputs(171);
    layer6_outputs(1549) <= (layer5_outputs(1923)) or (layer5_outputs(1486));
    layer6_outputs(1550) <= (layer5_outputs(2330)) and not (layer5_outputs(2474));
    layer6_outputs(1551) <= not(layer5_outputs(250));
    layer6_outputs(1552) <= '0';
    layer6_outputs(1553) <= not(layer5_outputs(1043));
    layer6_outputs(1554) <= (layer5_outputs(926)) and not (layer5_outputs(598));
    layer6_outputs(1555) <= not((layer5_outputs(221)) xor (layer5_outputs(396)));
    layer6_outputs(1556) <= (layer5_outputs(2298)) and (layer5_outputs(2473));
    layer6_outputs(1557) <= (layer5_outputs(1620)) or (layer5_outputs(1434));
    layer6_outputs(1558) <= (layer5_outputs(1667)) xor (layer5_outputs(2467));
    layer6_outputs(1559) <= not((layer5_outputs(981)) and (layer5_outputs(39)));
    layer6_outputs(1560) <= (layer5_outputs(1885)) and not (layer5_outputs(316));
    layer6_outputs(1561) <= layer5_outputs(33);
    layer6_outputs(1562) <= layer5_outputs(90);
    layer6_outputs(1563) <= (layer5_outputs(368)) and not (layer5_outputs(1696));
    layer6_outputs(1564) <= (layer5_outputs(282)) or (layer5_outputs(2122));
    layer6_outputs(1565) <= (layer5_outputs(395)) xor (layer5_outputs(1217));
    layer6_outputs(1566) <= (layer5_outputs(2437)) and not (layer5_outputs(514));
    layer6_outputs(1567) <= (layer5_outputs(2505)) and not (layer5_outputs(263));
    layer6_outputs(1568) <= layer5_outputs(1976);
    layer6_outputs(1569) <= (layer5_outputs(1502)) or (layer5_outputs(133));
    layer6_outputs(1570) <= not((layer5_outputs(2501)) xor (layer5_outputs(1820)));
    layer6_outputs(1571) <= not(layer5_outputs(1934));
    layer6_outputs(1572) <= not((layer5_outputs(1360)) xor (layer5_outputs(2201)));
    layer6_outputs(1573) <= (layer5_outputs(36)) or (layer5_outputs(709));
    layer6_outputs(1574) <= not(layer5_outputs(56));
    layer6_outputs(1575) <= not(layer5_outputs(2300));
    layer6_outputs(1576) <= layer5_outputs(1807);
    layer6_outputs(1577) <= (layer5_outputs(580)) and (layer5_outputs(401));
    layer6_outputs(1578) <= not(layer5_outputs(410));
    layer6_outputs(1579) <= not(layer5_outputs(54));
    layer6_outputs(1580) <= not((layer5_outputs(1945)) or (layer5_outputs(162)));
    layer6_outputs(1581) <= not(layer5_outputs(1477)) or (layer5_outputs(1731));
    layer6_outputs(1582) <= not((layer5_outputs(1056)) and (layer5_outputs(2233)));
    layer6_outputs(1583) <= not(layer5_outputs(1729));
    layer6_outputs(1584) <= not(layer5_outputs(1853));
    layer6_outputs(1585) <= layer5_outputs(238);
    layer6_outputs(1586) <= not(layer5_outputs(1568));
    layer6_outputs(1587) <= not(layer5_outputs(1343)) or (layer5_outputs(646));
    layer6_outputs(1588) <= not(layer5_outputs(347));
    layer6_outputs(1589) <= layer5_outputs(306);
    layer6_outputs(1590) <= layer5_outputs(61);
    layer6_outputs(1591) <= not(layer5_outputs(854));
    layer6_outputs(1592) <= (layer5_outputs(1725)) or (layer5_outputs(1082));
    layer6_outputs(1593) <= not(layer5_outputs(1551));
    layer6_outputs(1594) <= (layer5_outputs(294)) and not (layer5_outputs(492));
    layer6_outputs(1595) <= not(layer5_outputs(333));
    layer6_outputs(1596) <= (layer5_outputs(1925)) and not (layer5_outputs(2072));
    layer6_outputs(1597) <= (layer5_outputs(418)) and not (layer5_outputs(1061));
    layer6_outputs(1598) <= (layer5_outputs(1797)) and not (layer5_outputs(359));
    layer6_outputs(1599) <= (layer5_outputs(300)) and not (layer5_outputs(2469));
    layer6_outputs(1600) <= not(layer5_outputs(671));
    layer6_outputs(1601) <= layer5_outputs(513);
    layer6_outputs(1602) <= layer5_outputs(1653);
    layer6_outputs(1603) <= (layer5_outputs(1067)) or (layer5_outputs(518));
    layer6_outputs(1604) <= layer5_outputs(931);
    layer6_outputs(1605) <= not(layer5_outputs(18)) or (layer5_outputs(902));
    layer6_outputs(1606) <= layer5_outputs(1337);
    layer6_outputs(1607) <= (layer5_outputs(37)) or (layer5_outputs(1736));
    layer6_outputs(1608) <= not(layer5_outputs(2545));
    layer6_outputs(1609) <= not((layer5_outputs(247)) xor (layer5_outputs(1068)));
    layer6_outputs(1610) <= (layer5_outputs(481)) and not (layer5_outputs(2196));
    layer6_outputs(1611) <= layer5_outputs(1907);
    layer6_outputs(1612) <= not(layer5_outputs(1605));
    layer6_outputs(1613) <= not(layer5_outputs(636));
    layer6_outputs(1614) <= not(layer5_outputs(2209));
    layer6_outputs(1615) <= not(layer5_outputs(213));
    layer6_outputs(1616) <= not(layer5_outputs(659));
    layer6_outputs(1617) <= not(layer5_outputs(2405));
    layer6_outputs(1618) <= not((layer5_outputs(1445)) xor (layer5_outputs(2499)));
    layer6_outputs(1619) <= layer5_outputs(2032);
    layer6_outputs(1620) <= layer5_outputs(126);
    layer6_outputs(1621) <= not(layer5_outputs(945));
    layer6_outputs(1622) <= not(layer5_outputs(104));
    layer6_outputs(1623) <= not(layer5_outputs(1660));
    layer6_outputs(1624) <= layer5_outputs(305);
    layer6_outputs(1625) <= not((layer5_outputs(1686)) xor (layer5_outputs(2111)));
    layer6_outputs(1626) <= not(layer5_outputs(736));
    layer6_outputs(1627) <= layer5_outputs(395);
    layer6_outputs(1628) <= (layer5_outputs(1973)) and not (layer5_outputs(1964));
    layer6_outputs(1629) <= layer5_outputs(1643);
    layer6_outputs(1630) <= layer5_outputs(684);
    layer6_outputs(1631) <= (layer5_outputs(2323)) and (layer5_outputs(2528));
    layer6_outputs(1632) <= (layer5_outputs(1703)) and not (layer5_outputs(538));
    layer6_outputs(1633) <= not(layer5_outputs(1017));
    layer6_outputs(1634) <= not(layer5_outputs(2447));
    layer6_outputs(1635) <= not(layer5_outputs(2053));
    layer6_outputs(1636) <= not(layer5_outputs(1679));
    layer6_outputs(1637) <= not((layer5_outputs(2153)) and (layer5_outputs(1136)));
    layer6_outputs(1638) <= (layer5_outputs(2515)) xor (layer5_outputs(1436));
    layer6_outputs(1639) <= not(layer5_outputs(466));
    layer6_outputs(1640) <= not((layer5_outputs(509)) xor (layer5_outputs(1381)));
    layer6_outputs(1641) <= not(layer5_outputs(408));
    layer6_outputs(1642) <= (layer5_outputs(229)) and not (layer5_outputs(2324));
    layer6_outputs(1643) <= layer5_outputs(869);
    layer6_outputs(1644) <= not(layer5_outputs(1110)) or (layer5_outputs(986));
    layer6_outputs(1645) <= not((layer5_outputs(1911)) xor (layer5_outputs(795)));
    layer6_outputs(1646) <= (layer5_outputs(1628)) and not (layer5_outputs(1325));
    layer6_outputs(1647) <= layer5_outputs(179);
    layer6_outputs(1648) <= not(layer5_outputs(2262));
    layer6_outputs(1649) <= layer5_outputs(2555);
    layer6_outputs(1650) <= not(layer5_outputs(1613));
    layer6_outputs(1651) <= not((layer5_outputs(766)) xor (layer5_outputs(2479)));
    layer6_outputs(1652) <= layer5_outputs(2437);
    layer6_outputs(1653) <= layer5_outputs(2381);
    layer6_outputs(1654) <= layer5_outputs(405);
    layer6_outputs(1655) <= not(layer5_outputs(1884));
    layer6_outputs(1656) <= not((layer5_outputs(48)) or (layer5_outputs(654)));
    layer6_outputs(1657) <= not(layer5_outputs(1450));
    layer6_outputs(1658) <= not(layer5_outputs(1198));
    layer6_outputs(1659) <= (layer5_outputs(64)) and (layer5_outputs(241));
    layer6_outputs(1660) <= not(layer5_outputs(1980)) or (layer5_outputs(1866));
    layer6_outputs(1661) <= not(layer5_outputs(1829)) or (layer5_outputs(220));
    layer6_outputs(1662) <= layer5_outputs(621);
    layer6_outputs(1663) <= layer5_outputs(29);
    layer6_outputs(1664) <= not((layer5_outputs(2451)) and (layer5_outputs(1886)));
    layer6_outputs(1665) <= not(layer5_outputs(1550));
    layer6_outputs(1666) <= not(layer5_outputs(813));
    layer6_outputs(1667) <= (layer5_outputs(1155)) and not (layer5_outputs(1422));
    layer6_outputs(1668) <= layer5_outputs(554);
    layer6_outputs(1669) <= (layer5_outputs(741)) and not (layer5_outputs(280));
    layer6_outputs(1670) <= not(layer5_outputs(1259));
    layer6_outputs(1671) <= layer5_outputs(328);
    layer6_outputs(1672) <= not(layer5_outputs(880));
    layer6_outputs(1673) <= not((layer5_outputs(1499)) and (layer5_outputs(15)));
    layer6_outputs(1674) <= '0';
    layer6_outputs(1675) <= '0';
    layer6_outputs(1676) <= layer5_outputs(744);
    layer6_outputs(1677) <= (layer5_outputs(2351)) and (layer5_outputs(0));
    layer6_outputs(1678) <= not(layer5_outputs(1337));
    layer6_outputs(1679) <= layer5_outputs(532);
    layer6_outputs(1680) <= (layer5_outputs(1060)) xor (layer5_outputs(665));
    layer6_outputs(1681) <= (layer5_outputs(1837)) and (layer5_outputs(1539));
    layer6_outputs(1682) <= not(layer5_outputs(825));
    layer6_outputs(1683) <= layer5_outputs(275);
    layer6_outputs(1684) <= (layer5_outputs(2422)) or (layer5_outputs(184));
    layer6_outputs(1685) <= layer5_outputs(1964);
    layer6_outputs(1686) <= not(layer5_outputs(1276)) or (layer5_outputs(1302));
    layer6_outputs(1687) <= (layer5_outputs(782)) xor (layer5_outputs(288));
    layer6_outputs(1688) <= not(layer5_outputs(1913)) or (layer5_outputs(504));
    layer6_outputs(1689) <= not(layer5_outputs(1239));
    layer6_outputs(1690) <= layer5_outputs(126);
    layer6_outputs(1691) <= (layer5_outputs(1066)) and not (layer5_outputs(2257));
    layer6_outputs(1692) <= not((layer5_outputs(154)) and (layer5_outputs(2205)));
    layer6_outputs(1693) <= (layer5_outputs(560)) and not (layer5_outputs(662));
    layer6_outputs(1694) <= (layer5_outputs(1861)) and (layer5_outputs(545));
    layer6_outputs(1695) <= (layer5_outputs(1101)) and not (layer5_outputs(856));
    layer6_outputs(1696) <= not(layer5_outputs(1814));
    layer6_outputs(1697) <= layer5_outputs(2184);
    layer6_outputs(1698) <= not(layer5_outputs(1520));
    layer6_outputs(1699) <= layer5_outputs(1787);
    layer6_outputs(1700) <= layer5_outputs(627);
    layer6_outputs(1701) <= '1';
    layer6_outputs(1702) <= not(layer5_outputs(1872));
    layer6_outputs(1703) <= layer5_outputs(659);
    layer6_outputs(1704) <= layer5_outputs(2037);
    layer6_outputs(1705) <= not(layer5_outputs(2047));
    layer6_outputs(1706) <= not(layer5_outputs(2273)) or (layer5_outputs(1639));
    layer6_outputs(1707) <= (layer5_outputs(38)) or (layer5_outputs(2400));
    layer6_outputs(1708) <= not(layer5_outputs(1393));
    layer6_outputs(1709) <= not(layer5_outputs(125));
    layer6_outputs(1710) <= (layer5_outputs(2537)) xor (layer5_outputs(1141));
    layer6_outputs(1711) <= (layer5_outputs(1329)) xor (layer5_outputs(2462));
    layer6_outputs(1712) <= layer5_outputs(262);
    layer6_outputs(1713) <= (layer5_outputs(2510)) and not (layer5_outputs(2530));
    layer6_outputs(1714) <= (layer5_outputs(474)) or (layer5_outputs(846));
    layer6_outputs(1715) <= not(layer5_outputs(388));
    layer6_outputs(1716) <= layer5_outputs(2177);
    layer6_outputs(1717) <= not(layer5_outputs(2502));
    layer6_outputs(1718) <= layer5_outputs(1593);
    layer6_outputs(1719) <= layer5_outputs(2429);
    layer6_outputs(1720) <= not(layer5_outputs(2481));
    layer6_outputs(1721) <= (layer5_outputs(767)) and not (layer5_outputs(9));
    layer6_outputs(1722) <= not(layer5_outputs(2135));
    layer6_outputs(1723) <= layer5_outputs(569);
    layer6_outputs(1724) <= not(layer5_outputs(1119));
    layer6_outputs(1725) <= not(layer5_outputs(1775));
    layer6_outputs(1726) <= not(layer5_outputs(1654));
    layer6_outputs(1727) <= not(layer5_outputs(1368));
    layer6_outputs(1728) <= (layer5_outputs(863)) xor (layer5_outputs(203));
    layer6_outputs(1729) <= not(layer5_outputs(1621));
    layer6_outputs(1730) <= (layer5_outputs(810)) and (layer5_outputs(2452));
    layer6_outputs(1731) <= layer5_outputs(1);
    layer6_outputs(1732) <= not(layer5_outputs(193));
    layer6_outputs(1733) <= not(layer5_outputs(2176));
    layer6_outputs(1734) <= (layer5_outputs(63)) and not (layer5_outputs(2514));
    layer6_outputs(1735) <= not(layer5_outputs(1850)) or (layer5_outputs(727));
    layer6_outputs(1736) <= (layer5_outputs(2487)) and not (layer5_outputs(2229));
    layer6_outputs(1737) <= not((layer5_outputs(2208)) or (layer5_outputs(707)));
    layer6_outputs(1738) <= not(layer5_outputs(1667));
    layer6_outputs(1739) <= (layer5_outputs(97)) and not (layer5_outputs(701));
    layer6_outputs(1740) <= layer5_outputs(1334);
    layer6_outputs(1741) <= not(layer5_outputs(1993));
    layer6_outputs(1742) <= not((layer5_outputs(1863)) and (layer5_outputs(1522)));
    layer6_outputs(1743) <= layer5_outputs(975);
    layer6_outputs(1744) <= layer5_outputs(1634);
    layer6_outputs(1745) <= (layer5_outputs(1756)) xor (layer5_outputs(119));
    layer6_outputs(1746) <= not((layer5_outputs(109)) xor (layer5_outputs(2212)));
    layer6_outputs(1747) <= layer5_outputs(290);
    layer6_outputs(1748) <= not((layer5_outputs(1421)) or (layer5_outputs(271)));
    layer6_outputs(1749) <= (layer5_outputs(1596)) and not (layer5_outputs(2411));
    layer6_outputs(1750) <= not(layer5_outputs(1137)) or (layer5_outputs(988));
    layer6_outputs(1751) <= layer5_outputs(888);
    layer6_outputs(1752) <= (layer5_outputs(138)) xor (layer5_outputs(2198));
    layer6_outputs(1753) <= layer5_outputs(2518);
    layer6_outputs(1754) <= (layer5_outputs(603)) xor (layer5_outputs(113));
    layer6_outputs(1755) <= (layer5_outputs(293)) and not (layer5_outputs(770));
    layer6_outputs(1756) <= (layer5_outputs(2362)) and not (layer5_outputs(145));
    layer6_outputs(1757) <= not(layer5_outputs(350));
    layer6_outputs(1758) <= not(layer5_outputs(763));
    layer6_outputs(1759) <= '0';
    layer6_outputs(1760) <= layer5_outputs(1750);
    layer6_outputs(1761) <= layer5_outputs(1878);
    layer6_outputs(1762) <= (layer5_outputs(391)) and not (layer5_outputs(1026));
    layer6_outputs(1763) <= layer5_outputs(1913);
    layer6_outputs(1764) <= not(layer5_outputs(2092));
    layer6_outputs(1765) <= layer5_outputs(1441);
    layer6_outputs(1766) <= not(layer5_outputs(2324)) or (layer5_outputs(1555));
    layer6_outputs(1767) <= not(layer5_outputs(1721)) or (layer5_outputs(2206));
    layer6_outputs(1768) <= (layer5_outputs(642)) and not (layer5_outputs(1338));
    layer6_outputs(1769) <= not(layer5_outputs(1468));
    layer6_outputs(1770) <= not((layer5_outputs(1815)) xor (layer5_outputs(853)));
    layer6_outputs(1771) <= not(layer5_outputs(1000));
    layer6_outputs(1772) <= (layer5_outputs(1233)) and not (layer5_outputs(2246));
    layer6_outputs(1773) <= layer5_outputs(503);
    layer6_outputs(1774) <= layer5_outputs(2075);
    layer6_outputs(1775) <= not((layer5_outputs(1688)) and (layer5_outputs(1432)));
    layer6_outputs(1776) <= layer5_outputs(2294);
    layer6_outputs(1777) <= not(layer5_outputs(1528));
    layer6_outputs(1778) <= not(layer5_outputs(2160));
    layer6_outputs(1779) <= not((layer5_outputs(1192)) and (layer5_outputs(1086)));
    layer6_outputs(1780) <= layer5_outputs(1030);
    layer6_outputs(1781) <= not((layer5_outputs(2006)) or (layer5_outputs(155)));
    layer6_outputs(1782) <= not(layer5_outputs(1536)) or (layer5_outputs(2132));
    layer6_outputs(1783) <= not((layer5_outputs(1741)) and (layer5_outputs(2527)));
    layer6_outputs(1784) <= not((layer5_outputs(2078)) xor (layer5_outputs(118)));
    layer6_outputs(1785) <= layer5_outputs(1969);
    layer6_outputs(1786) <= layer5_outputs(175);
    layer6_outputs(1787) <= not(layer5_outputs(1928));
    layer6_outputs(1788) <= (layer5_outputs(2035)) xor (layer5_outputs(2356));
    layer6_outputs(1789) <= (layer5_outputs(564)) and not (layer5_outputs(1247));
    layer6_outputs(1790) <= not((layer5_outputs(2260)) and (layer5_outputs(2310)));
    layer6_outputs(1791) <= layer5_outputs(1977);
    layer6_outputs(1792) <= not(layer5_outputs(69)) or (layer5_outputs(952));
    layer6_outputs(1793) <= not(layer5_outputs(1660));
    layer6_outputs(1794) <= layer5_outputs(1753);
    layer6_outputs(1795) <= not(layer5_outputs(516));
    layer6_outputs(1796) <= (layer5_outputs(997)) and not (layer5_outputs(2432));
    layer6_outputs(1797) <= not(layer5_outputs(116)) or (layer5_outputs(2266));
    layer6_outputs(1798) <= (layer5_outputs(2308)) and (layer5_outputs(2332));
    layer6_outputs(1799) <= not(layer5_outputs(625));
    layer6_outputs(1800) <= layer5_outputs(587);
    layer6_outputs(1801) <= layer5_outputs(1500);
    layer6_outputs(1802) <= not(layer5_outputs(1744)) or (layer5_outputs(480));
    layer6_outputs(1803) <= (layer5_outputs(1229)) xor (layer5_outputs(2379));
    layer6_outputs(1804) <= not(layer5_outputs(2251)) or (layer5_outputs(1411));
    layer6_outputs(1805) <= not(layer5_outputs(1143));
    layer6_outputs(1806) <= not(layer5_outputs(245));
    layer6_outputs(1807) <= not((layer5_outputs(2485)) xor (layer5_outputs(1303)));
    layer6_outputs(1808) <= (layer5_outputs(2463)) xor (layer5_outputs(1271));
    layer6_outputs(1809) <= layer5_outputs(1540);
    layer6_outputs(1810) <= not(layer5_outputs(965));
    layer6_outputs(1811) <= layer5_outputs(1926);
    layer6_outputs(1812) <= layer5_outputs(1021);
    layer6_outputs(1813) <= not(layer5_outputs(1248));
    layer6_outputs(1814) <= not(layer5_outputs(164)) or (layer5_outputs(2405));
    layer6_outputs(1815) <= (layer5_outputs(909)) xor (layer5_outputs(890));
    layer6_outputs(1816) <= not((layer5_outputs(478)) xor (layer5_outputs(2356)));
    layer6_outputs(1817) <= layer5_outputs(2218);
    layer6_outputs(1818) <= layer5_outputs(1121);
    layer6_outputs(1819) <= layer5_outputs(677);
    layer6_outputs(1820) <= (layer5_outputs(1382)) and not (layer5_outputs(1178));
    layer6_outputs(1821) <= (layer5_outputs(1899)) xor (layer5_outputs(1800));
    layer6_outputs(1822) <= layer5_outputs(1417);
    layer6_outputs(1823) <= not(layer5_outputs(576));
    layer6_outputs(1824) <= not(layer5_outputs(1095));
    layer6_outputs(1825) <= not(layer5_outputs(1517)) or (layer5_outputs(2433));
    layer6_outputs(1826) <= (layer5_outputs(1040)) xor (layer5_outputs(1579));
    layer6_outputs(1827) <= not((layer5_outputs(1808)) or (layer5_outputs(622)));
    layer6_outputs(1828) <= '0';
    layer6_outputs(1829) <= not(layer5_outputs(797)) or (layer5_outputs(258));
    layer6_outputs(1830) <= (layer5_outputs(1553)) and (layer5_outputs(1189));
    layer6_outputs(1831) <= not(layer5_outputs(1277)) or (layer5_outputs(882));
    layer6_outputs(1832) <= layer5_outputs(615);
    layer6_outputs(1833) <= layer5_outputs(1762);
    layer6_outputs(1834) <= (layer5_outputs(2416)) or (layer5_outputs(1651));
    layer6_outputs(1835) <= (layer5_outputs(2475)) xor (layer5_outputs(604));
    layer6_outputs(1836) <= not(layer5_outputs(712));
    layer6_outputs(1837) <= not(layer5_outputs(1983)) or (layer5_outputs(1937));
    layer6_outputs(1838) <= not((layer5_outputs(976)) and (layer5_outputs(1501)));
    layer6_outputs(1839) <= (layer5_outputs(1063)) or (layer5_outputs(2287));
    layer6_outputs(1840) <= not(layer5_outputs(1932));
    layer6_outputs(1841) <= '0';
    layer6_outputs(1842) <= not(layer5_outputs(412));
    layer6_outputs(1843) <= layer5_outputs(2519);
    layer6_outputs(1844) <= layer5_outputs(711);
    layer6_outputs(1845) <= (layer5_outputs(1735)) and (layer5_outputs(2392));
    layer6_outputs(1846) <= (layer5_outputs(1050)) or (layer5_outputs(436));
    layer6_outputs(1847) <= not(layer5_outputs(380));
    layer6_outputs(1848) <= layer5_outputs(1743);
    layer6_outputs(1849) <= not(layer5_outputs(479));
    layer6_outputs(1850) <= not(layer5_outputs(329));
    layer6_outputs(1851) <= not((layer5_outputs(1653)) xor (layer5_outputs(1915)));
    layer6_outputs(1852) <= not((layer5_outputs(1620)) and (layer5_outputs(1747)));
    layer6_outputs(1853) <= (layer5_outputs(34)) or (layer5_outputs(1448));
    layer6_outputs(1854) <= not(layer5_outputs(2003));
    layer6_outputs(1855) <= not((layer5_outputs(17)) xor (layer5_outputs(509)));
    layer6_outputs(1856) <= not(layer5_outputs(169));
    layer6_outputs(1857) <= not((layer5_outputs(1899)) xor (layer5_outputs(1444)));
    layer6_outputs(1858) <= not(layer5_outputs(1574));
    layer6_outputs(1859) <= not(layer5_outputs(224));
    layer6_outputs(1860) <= layer5_outputs(2120);
    layer6_outputs(1861) <= layer5_outputs(634);
    layer6_outputs(1862) <= layer5_outputs(1924);
    layer6_outputs(1863) <= layer5_outputs(2484);
    layer6_outputs(1864) <= layer5_outputs(670);
    layer6_outputs(1865) <= not(layer5_outputs(1480)) or (layer5_outputs(1703));
    layer6_outputs(1866) <= layer5_outputs(1984);
    layer6_outputs(1867) <= (layer5_outputs(563)) and not (layer5_outputs(1797));
    layer6_outputs(1868) <= layer5_outputs(1685);
    layer6_outputs(1869) <= not((layer5_outputs(1819)) or (layer5_outputs(231)));
    layer6_outputs(1870) <= layer5_outputs(2525);
    layer6_outputs(1871) <= (layer5_outputs(249)) and not (layer5_outputs(256));
    layer6_outputs(1872) <= not(layer5_outputs(954)) or (layer5_outputs(2156));
    layer6_outputs(1873) <= (layer5_outputs(1207)) xor (layer5_outputs(1302));
    layer6_outputs(1874) <= not(layer5_outputs(74));
    layer6_outputs(1875) <= not(layer5_outputs(291));
    layer6_outputs(1876) <= (layer5_outputs(1970)) and not (layer5_outputs(1855));
    layer6_outputs(1877) <= not((layer5_outputs(1763)) or (layer5_outputs(182)));
    layer6_outputs(1878) <= layer5_outputs(1255);
    layer6_outputs(1879) <= layer5_outputs(2218);
    layer6_outputs(1880) <= layer5_outputs(1335);
    layer6_outputs(1881) <= layer5_outputs(814);
    layer6_outputs(1882) <= (layer5_outputs(45)) and not (layer5_outputs(337));
    layer6_outputs(1883) <= layer5_outputs(831);
    layer6_outputs(1884) <= layer5_outputs(1092);
    layer6_outputs(1885) <= not((layer5_outputs(1912)) xor (layer5_outputs(781)));
    layer6_outputs(1886) <= not(layer5_outputs(2476));
    layer6_outputs(1887) <= (layer5_outputs(1037)) and (layer5_outputs(462));
    layer6_outputs(1888) <= not(layer5_outputs(1086)) or (layer5_outputs(2471));
    layer6_outputs(1889) <= not((layer5_outputs(690)) or (layer5_outputs(2045)));
    layer6_outputs(1890) <= (layer5_outputs(210)) and not (layer5_outputs(2232));
    layer6_outputs(1891) <= not(layer5_outputs(1220));
    layer6_outputs(1892) <= (layer5_outputs(571)) and (layer5_outputs(2141));
    layer6_outputs(1893) <= not((layer5_outputs(2396)) and (layer5_outputs(871)));
    layer6_outputs(1894) <= not(layer5_outputs(82));
    layer6_outputs(1895) <= layer5_outputs(1150);
    layer6_outputs(1896) <= not(layer5_outputs(912));
    layer6_outputs(1897) <= not(layer5_outputs(1630));
    layer6_outputs(1898) <= not(layer5_outputs(370));
    layer6_outputs(1899) <= not(layer5_outputs(601));
    layer6_outputs(1900) <= (layer5_outputs(2534)) and not (layer5_outputs(1781));
    layer6_outputs(1901) <= not(layer5_outputs(2149));
    layer6_outputs(1902) <= not((layer5_outputs(738)) xor (layer5_outputs(1887)));
    layer6_outputs(1903) <= not(layer5_outputs(284));
    layer6_outputs(1904) <= not((layer5_outputs(322)) xor (layer5_outputs(1681)));
    layer6_outputs(1905) <= layer5_outputs(1435);
    layer6_outputs(1906) <= not(layer5_outputs(1968));
    layer6_outputs(1907) <= (layer5_outputs(1736)) or (layer5_outputs(2005));
    layer6_outputs(1908) <= layer5_outputs(1529);
    layer6_outputs(1909) <= not(layer5_outputs(69));
    layer6_outputs(1910) <= (layer5_outputs(157)) or (layer5_outputs(582));
    layer6_outputs(1911) <= not((layer5_outputs(821)) or (layer5_outputs(2018)));
    layer6_outputs(1912) <= not(layer5_outputs(1482));
    layer6_outputs(1913) <= (layer5_outputs(1059)) xor (layer5_outputs(632));
    layer6_outputs(1914) <= not(layer5_outputs(526));
    layer6_outputs(1915) <= '0';
    layer6_outputs(1916) <= not(layer5_outputs(323));
    layer6_outputs(1917) <= not(layer5_outputs(506));
    layer6_outputs(1918) <= (layer5_outputs(1410)) and not (layer5_outputs(995));
    layer6_outputs(1919) <= layer5_outputs(929);
    layer6_outputs(1920) <= layer5_outputs(688);
    layer6_outputs(1921) <= layer5_outputs(1001);
    layer6_outputs(1922) <= not(layer5_outputs(1586)) or (layer5_outputs(266));
    layer6_outputs(1923) <= (layer5_outputs(289)) or (layer5_outputs(2480));
    layer6_outputs(1924) <= (layer5_outputs(1485)) and not (layer5_outputs(330));
    layer6_outputs(1925) <= not(layer5_outputs(227));
    layer6_outputs(1926) <= not((layer5_outputs(777)) and (layer5_outputs(2332)));
    layer6_outputs(1927) <= (layer5_outputs(204)) xor (layer5_outputs(1169));
    layer6_outputs(1928) <= not(layer5_outputs(2317));
    layer6_outputs(1929) <= layer5_outputs(1218);
    layer6_outputs(1930) <= not((layer5_outputs(1631)) or (layer5_outputs(1070)));
    layer6_outputs(1931) <= layer5_outputs(1216);
    layer6_outputs(1932) <= not(layer5_outputs(377)) or (layer5_outputs(580));
    layer6_outputs(1933) <= layer5_outputs(1692);
    layer6_outputs(1934) <= not((layer5_outputs(2290)) xor (layer5_outputs(2118)));
    layer6_outputs(1935) <= (layer5_outputs(201)) and not (layer5_outputs(1991));
    layer6_outputs(1936) <= not(layer5_outputs(1578)) or (layer5_outputs(318));
    layer6_outputs(1937) <= not(layer5_outputs(471));
    layer6_outputs(1938) <= not(layer5_outputs(1591)) or (layer5_outputs(708));
    layer6_outputs(1939) <= (layer5_outputs(2478)) xor (layer5_outputs(936));
    layer6_outputs(1940) <= (layer5_outputs(759)) and not (layer5_outputs(1584));
    layer6_outputs(1941) <= (layer5_outputs(59)) and (layer5_outputs(649));
    layer6_outputs(1942) <= not(layer5_outputs(2152)) or (layer5_outputs(1326));
    layer6_outputs(1943) <= layer5_outputs(16);
    layer6_outputs(1944) <= (layer5_outputs(1765)) and not (layer5_outputs(2131));
    layer6_outputs(1945) <= layer5_outputs(2040);
    layer6_outputs(1946) <= not((layer5_outputs(1808)) xor (layer5_outputs(1386)));
    layer6_outputs(1947) <= (layer5_outputs(1961)) xor (layer5_outputs(2391));
    layer6_outputs(1948) <= not(layer5_outputs(1771)) or (layer5_outputs(1079));
    layer6_outputs(1949) <= not(layer5_outputs(1045));
    layer6_outputs(1950) <= layer5_outputs(1120);
    layer6_outputs(1951) <= (layer5_outputs(2259)) and not (layer5_outputs(1035));
    layer6_outputs(1952) <= (layer5_outputs(2252)) and not (layer5_outputs(2291));
    layer6_outputs(1953) <= not((layer5_outputs(355)) and (layer5_outputs(447)));
    layer6_outputs(1954) <= layer5_outputs(936);
    layer6_outputs(1955) <= not((layer5_outputs(195)) xor (layer5_outputs(1966)));
    layer6_outputs(1956) <= not((layer5_outputs(2208)) and (layer5_outputs(2151)));
    layer6_outputs(1957) <= not(layer5_outputs(607));
    layer6_outputs(1958) <= not(layer5_outputs(728));
    layer6_outputs(1959) <= not(layer5_outputs(963));
    layer6_outputs(1960) <= layer5_outputs(2278);
    layer6_outputs(1961) <= layer5_outputs(2043);
    layer6_outputs(1962) <= layer5_outputs(433);
    layer6_outputs(1963) <= (layer5_outputs(356)) xor (layer5_outputs(2450));
    layer6_outputs(1964) <= not(layer5_outputs(50));
    layer6_outputs(1965) <= layer5_outputs(1892);
    layer6_outputs(1966) <= not(layer5_outputs(1196));
    layer6_outputs(1967) <= not(layer5_outputs(28)) or (layer5_outputs(389));
    layer6_outputs(1968) <= not(layer5_outputs(2012));
    layer6_outputs(1969) <= not((layer5_outputs(1549)) and (layer5_outputs(1449)));
    layer6_outputs(1970) <= layer5_outputs(2449);
    layer6_outputs(1971) <= (layer5_outputs(106)) or (layer5_outputs(826));
    layer6_outputs(1972) <= (layer5_outputs(89)) and not (layer5_outputs(1638));
    layer6_outputs(1973) <= not(layer5_outputs(2234)) or (layer5_outputs(1321));
    layer6_outputs(1974) <= layer5_outputs(1028);
    layer6_outputs(1975) <= (layer5_outputs(1560)) xor (layer5_outputs(106));
    layer6_outputs(1976) <= layer5_outputs(1843);
    layer6_outputs(1977) <= (layer5_outputs(486)) and not (layer5_outputs(2446));
    layer6_outputs(1978) <= not(layer5_outputs(722));
    layer6_outputs(1979) <= (layer5_outputs(843)) xor (layer5_outputs(672));
    layer6_outputs(1980) <= layer5_outputs(673);
    layer6_outputs(1981) <= not(layer5_outputs(619));
    layer6_outputs(1982) <= (layer5_outputs(426)) and not (layer5_outputs(1243));
    layer6_outputs(1983) <= layer5_outputs(1734);
    layer6_outputs(1984) <= layer5_outputs(869);
    layer6_outputs(1985) <= not(layer5_outputs(2099));
    layer6_outputs(1986) <= layer5_outputs(1926);
    layer6_outputs(1987) <= (layer5_outputs(550)) and not (layer5_outputs(860));
    layer6_outputs(1988) <= layer5_outputs(1556);
    layer6_outputs(1989) <= layer5_outputs(2466);
    layer6_outputs(1990) <= (layer5_outputs(879)) xor (layer5_outputs(1595));
    layer6_outputs(1991) <= (layer5_outputs(1513)) and not (layer5_outputs(171));
    layer6_outputs(1992) <= layer5_outputs(1530);
    layer6_outputs(1993) <= (layer5_outputs(1390)) or (layer5_outputs(358));
    layer6_outputs(1994) <= not((layer5_outputs(2386)) or (layer5_outputs(1959)));
    layer6_outputs(1995) <= not(layer5_outputs(1419)) or (layer5_outputs(494));
    layer6_outputs(1996) <= not(layer5_outputs(827));
    layer6_outputs(1997) <= layer5_outputs(1422);
    layer6_outputs(1998) <= (layer5_outputs(1580)) and not (layer5_outputs(2381));
    layer6_outputs(1999) <= layer5_outputs(1525);
    layer6_outputs(2000) <= (layer5_outputs(1076)) and not (layer5_outputs(19));
    layer6_outputs(2001) <= not(layer5_outputs(1600)) or (layer5_outputs(2094));
    layer6_outputs(2002) <= not(layer5_outputs(703));
    layer6_outputs(2003) <= layer5_outputs(539);
    layer6_outputs(2004) <= not(layer5_outputs(326));
    layer6_outputs(2005) <= layer5_outputs(1982);
    layer6_outputs(2006) <= not(layer5_outputs(1331));
    layer6_outputs(2007) <= not(layer5_outputs(897)) or (layer5_outputs(1949));
    layer6_outputs(2008) <= not((layer5_outputs(967)) and (layer5_outputs(2101)));
    layer6_outputs(2009) <= not(layer5_outputs(1008));
    layer6_outputs(2010) <= layer5_outputs(1795);
    layer6_outputs(2011) <= not((layer5_outputs(577)) and (layer5_outputs(2529)));
    layer6_outputs(2012) <= not(layer5_outputs(1909));
    layer6_outputs(2013) <= not(layer5_outputs(1288));
    layer6_outputs(2014) <= not(layer5_outputs(1132));
    layer6_outputs(2015) <= layer5_outputs(1591);
    layer6_outputs(2016) <= layer5_outputs(467);
    layer6_outputs(2017) <= not(layer5_outputs(552));
    layer6_outputs(2018) <= not((layer5_outputs(1317)) xor (layer5_outputs(834)));
    layer6_outputs(2019) <= (layer5_outputs(1244)) and (layer5_outputs(1191));
    layer6_outputs(2020) <= not(layer5_outputs(285)) or (layer5_outputs(1939));
    layer6_outputs(2021) <= not(layer5_outputs(1557));
    layer6_outputs(2022) <= (layer5_outputs(1895)) and not (layer5_outputs(561));
    layer6_outputs(2023) <= (layer5_outputs(2347)) or (layer5_outputs(941));
    layer6_outputs(2024) <= (layer5_outputs(1677)) and not (layer5_outputs(2245));
    layer6_outputs(2025) <= (layer5_outputs(172)) and (layer5_outputs(577));
    layer6_outputs(2026) <= not((layer5_outputs(1508)) or (layer5_outputs(457)));
    layer6_outputs(2027) <= (layer5_outputs(2145)) and (layer5_outputs(2280));
    layer6_outputs(2028) <= layer5_outputs(2095);
    layer6_outputs(2029) <= layer5_outputs(2251);
    layer6_outputs(2030) <= not(layer5_outputs(1017));
    layer6_outputs(2031) <= not(layer5_outputs(1127));
    layer6_outputs(2032) <= (layer5_outputs(1572)) and not (layer5_outputs(1956));
    layer6_outputs(2033) <= not(layer5_outputs(2363));
    layer6_outputs(2034) <= not(layer5_outputs(896)) or (layer5_outputs(663));
    layer6_outputs(2035) <= not(layer5_outputs(713));
    layer6_outputs(2036) <= not(layer5_outputs(1182));
    layer6_outputs(2037) <= layer5_outputs(675);
    layer6_outputs(2038) <= layer5_outputs(613);
    layer6_outputs(2039) <= layer5_outputs(1226);
    layer6_outputs(2040) <= not(layer5_outputs(1034));
    layer6_outputs(2041) <= not(layer5_outputs(1494));
    layer6_outputs(2042) <= (layer5_outputs(1744)) and (layer5_outputs(295));
    layer6_outputs(2043) <= not((layer5_outputs(1595)) xor (layer5_outputs(2149)));
    layer6_outputs(2044) <= not(layer5_outputs(1441)) or (layer5_outputs(1013));
    layer6_outputs(2045) <= not(layer5_outputs(2121)) or (layer5_outputs(1296));
    layer6_outputs(2046) <= not((layer5_outputs(2338)) or (layer5_outputs(2435)));
    layer6_outputs(2047) <= not((layer5_outputs(1635)) and (layer5_outputs(1726)));
    layer6_outputs(2048) <= not(layer5_outputs(2352)) or (layer5_outputs(2193));
    layer6_outputs(2049) <= (layer5_outputs(1552)) and (layer5_outputs(1273));
    layer6_outputs(2050) <= not(layer5_outputs(2270));
    layer6_outputs(2051) <= not(layer5_outputs(1516));
    layer6_outputs(2052) <= not(layer5_outputs(1697)) or (layer5_outputs(1611));
    layer6_outputs(2053) <= (layer5_outputs(293)) and not (layer5_outputs(2403));
    layer6_outputs(2054) <= not(layer5_outputs(2087));
    layer6_outputs(2055) <= not(layer5_outputs(845)) or (layer5_outputs(794));
    layer6_outputs(2056) <= not((layer5_outputs(551)) and (layer5_outputs(256)));
    layer6_outputs(2057) <= not((layer5_outputs(2013)) and (layer5_outputs(2007)));
    layer6_outputs(2058) <= layer5_outputs(2140);
    layer6_outputs(2059) <= not((layer5_outputs(1399)) xor (layer5_outputs(1802)));
    layer6_outputs(2060) <= (layer5_outputs(1048)) or (layer5_outputs(667));
    layer6_outputs(2061) <= not((layer5_outputs(2412)) and (layer5_outputs(345)));
    layer6_outputs(2062) <= (layer5_outputs(984)) and not (layer5_outputs(1518));
    layer6_outputs(2063) <= layer5_outputs(1742);
    layer6_outputs(2064) <= not(layer5_outputs(1838));
    layer6_outputs(2065) <= (layer5_outputs(909)) and (layer5_outputs(766));
    layer6_outputs(2066) <= not(layer5_outputs(2440));
    layer6_outputs(2067) <= not((layer5_outputs(575)) xor (layer5_outputs(2460)));
    layer6_outputs(2068) <= not(layer5_outputs(912));
    layer6_outputs(2069) <= layer5_outputs(1758);
    layer6_outputs(2070) <= layer5_outputs(1565);
    layer6_outputs(2071) <= layer5_outputs(238);
    layer6_outputs(2072) <= (layer5_outputs(1637)) and not (layer5_outputs(722));
    layer6_outputs(2073) <= not(layer5_outputs(1897));
    layer6_outputs(2074) <= layer5_outputs(1370);
    layer6_outputs(2075) <= not(layer5_outputs(1589));
    layer6_outputs(2076) <= layer5_outputs(1498);
    layer6_outputs(2077) <= (layer5_outputs(727)) and (layer5_outputs(2198));
    layer6_outputs(2078) <= not(layer5_outputs(2552));
    layer6_outputs(2079) <= layer5_outputs(1742);
    layer6_outputs(2080) <= not((layer5_outputs(2544)) xor (layer5_outputs(1451)));
    layer6_outputs(2081) <= layer5_outputs(673);
    layer6_outputs(2082) <= (layer5_outputs(87)) and not (layer5_outputs(1436));
    layer6_outputs(2083) <= not((layer5_outputs(2302)) or (layer5_outputs(1345)));
    layer6_outputs(2084) <= (layer5_outputs(1148)) and not (layer5_outputs(2103));
    layer6_outputs(2085) <= (layer5_outputs(2061)) xor (layer5_outputs(1122));
    layer6_outputs(2086) <= '1';
    layer6_outputs(2087) <= (layer5_outputs(477)) xor (layer5_outputs(2038));
    layer6_outputs(2088) <= (layer5_outputs(2389)) and not (layer5_outputs(1529));
    layer6_outputs(2089) <= not((layer5_outputs(641)) or (layer5_outputs(1495)));
    layer6_outputs(2090) <= not((layer5_outputs(21)) xor (layer5_outputs(1985)));
    layer6_outputs(2091) <= (layer5_outputs(89)) and not (layer5_outputs(2026));
    layer6_outputs(2092) <= not((layer5_outputs(1265)) and (layer5_outputs(1531)));
    layer6_outputs(2093) <= (layer5_outputs(1376)) and (layer5_outputs(1581));
    layer6_outputs(2094) <= not(layer5_outputs(2247));
    layer6_outputs(2095) <= not(layer5_outputs(1940)) or (layer5_outputs(892));
    layer6_outputs(2096) <= '1';
    layer6_outputs(2097) <= not((layer5_outputs(2498)) xor (layer5_outputs(1147)));
    layer6_outputs(2098) <= not(layer5_outputs(1396)) or (layer5_outputs(1467));
    layer6_outputs(2099) <= layer5_outputs(2390);
    layer6_outputs(2100) <= (layer5_outputs(2469)) or (layer5_outputs(1504));
    layer6_outputs(2101) <= not(layer5_outputs(2464)) or (layer5_outputs(689));
    layer6_outputs(2102) <= '1';
    layer6_outputs(2103) <= not((layer5_outputs(1959)) and (layer5_outputs(124)));
    layer6_outputs(2104) <= not(layer5_outputs(185));
    layer6_outputs(2105) <= (layer5_outputs(1080)) and (layer5_outputs(1124));
    layer6_outputs(2106) <= not(layer5_outputs(572)) or (layer5_outputs(304));
    layer6_outputs(2107) <= layer5_outputs(1503);
    layer6_outputs(2108) <= (layer5_outputs(1713)) or (layer5_outputs(1437));
    layer6_outputs(2109) <= (layer5_outputs(2142)) or (layer5_outputs(1456));
    layer6_outputs(2110) <= layer5_outputs(590);
    layer6_outputs(2111) <= (layer5_outputs(601)) and not (layer5_outputs(961));
    layer6_outputs(2112) <= (layer5_outputs(1019)) and not (layer5_outputs(819));
    layer6_outputs(2113) <= layer5_outputs(1579);
    layer6_outputs(2114) <= not((layer5_outputs(2104)) and (layer5_outputs(2019)));
    layer6_outputs(2115) <= not((layer5_outputs(628)) and (layer5_outputs(2073)));
    layer6_outputs(2116) <= layer5_outputs(2559);
    layer6_outputs(2117) <= not(layer5_outputs(784));
    layer6_outputs(2118) <= layer5_outputs(2135);
    layer6_outputs(2119) <= layer5_outputs(88);
    layer6_outputs(2120) <= not((layer5_outputs(1823)) xor (layer5_outputs(2042)));
    layer6_outputs(2121) <= not(layer5_outputs(144));
    layer6_outputs(2122) <= (layer5_outputs(1258)) and not (layer5_outputs(163));
    layer6_outputs(2123) <= (layer5_outputs(523)) and (layer5_outputs(2055));
    layer6_outputs(2124) <= (layer5_outputs(139)) and not (layer5_outputs(1386));
    layer6_outputs(2125) <= (layer5_outputs(611)) and (layer5_outputs(1974));
    layer6_outputs(2126) <= (layer5_outputs(432)) or (layer5_outputs(472));
    layer6_outputs(2127) <= not((layer5_outputs(2361)) or (layer5_outputs(1384)));
    layer6_outputs(2128) <= not(layer5_outputs(620));
    layer6_outputs(2129) <= (layer5_outputs(2034)) and (layer5_outputs(1064));
    layer6_outputs(2130) <= not((layer5_outputs(153)) xor (layer5_outputs(826)));
    layer6_outputs(2131) <= not(layer5_outputs(1928));
    layer6_outputs(2132) <= not(layer5_outputs(2036)) or (layer5_outputs(1427));
    layer6_outputs(2133) <= not((layer5_outputs(610)) and (layer5_outputs(298)));
    layer6_outputs(2134) <= not((layer5_outputs(899)) xor (layer5_outputs(1953)));
    layer6_outputs(2135) <= layer5_outputs(1233);
    layer6_outputs(2136) <= layer5_outputs(1650);
    layer6_outputs(2137) <= not(layer5_outputs(2225));
    layer6_outputs(2138) <= not((layer5_outputs(1670)) xor (layer5_outputs(1192)));
    layer6_outputs(2139) <= not(layer5_outputs(1399)) or (layer5_outputs(1786));
    layer6_outputs(2140) <= not(layer5_outputs(978));
    layer6_outputs(2141) <= not(layer5_outputs(1156));
    layer6_outputs(2142) <= not((layer5_outputs(1983)) xor (layer5_outputs(1675)));
    layer6_outputs(2143) <= layer5_outputs(2481);
    layer6_outputs(2144) <= (layer5_outputs(31)) xor (layer5_outputs(2220));
    layer6_outputs(2145) <= not(layer5_outputs(771));
    layer6_outputs(2146) <= layer5_outputs(2300);
    layer6_outputs(2147) <= not(layer5_outputs(1813));
    layer6_outputs(2148) <= layer5_outputs(1722);
    layer6_outputs(2149) <= not(layer5_outputs(151));
    layer6_outputs(2150) <= not(layer5_outputs(1702));
    layer6_outputs(2151) <= layer5_outputs(2404);
    layer6_outputs(2152) <= not(layer5_outputs(1728)) or (layer5_outputs(1204));
    layer6_outputs(2153) <= not(layer5_outputs(2473)) or (layer5_outputs(1911));
    layer6_outputs(2154) <= not(layer5_outputs(2442));
    layer6_outputs(2155) <= not(layer5_outputs(2030));
    layer6_outputs(2156) <= layer5_outputs(1021);
    layer6_outputs(2157) <= (layer5_outputs(1859)) xor (layer5_outputs(2410));
    layer6_outputs(2158) <= not((layer5_outputs(1365)) and (layer5_outputs(295)));
    layer6_outputs(2159) <= layer5_outputs(838);
    layer6_outputs(2160) <= (layer5_outputs(1962)) xor (layer5_outputs(1397));
    layer6_outputs(2161) <= not(layer5_outputs(2263));
    layer6_outputs(2162) <= not(layer5_outputs(1839));
    layer6_outputs(2163) <= not((layer5_outputs(2367)) or (layer5_outputs(919)));
    layer6_outputs(2164) <= not(layer5_outputs(76));
    layer6_outputs(2165) <= not(layer5_outputs(2209));
    layer6_outputs(2166) <= not(layer5_outputs(1073));
    layer6_outputs(2167) <= layer5_outputs(1818);
    layer6_outputs(2168) <= not(layer5_outputs(83)) or (layer5_outputs(2238));
    layer6_outputs(2169) <= not((layer5_outputs(688)) or (layer5_outputs(1673)));
    layer6_outputs(2170) <= '0';
    layer6_outputs(2171) <= (layer5_outputs(1626)) xor (layer5_outputs(851));
    layer6_outputs(2172) <= not((layer5_outputs(262)) and (layer5_outputs(2312)));
    layer6_outputs(2173) <= not(layer5_outputs(2088)) or (layer5_outputs(2493));
    layer6_outputs(2174) <= not(layer5_outputs(1760));
    layer6_outputs(2175) <= not(layer5_outputs(1009));
    layer6_outputs(2176) <= not((layer5_outputs(219)) xor (layer5_outputs(242)));
    layer6_outputs(2177) <= not(layer5_outputs(700));
    layer6_outputs(2178) <= layer5_outputs(392);
    layer6_outputs(2179) <= (layer5_outputs(507)) xor (layer5_outputs(2219));
    layer6_outputs(2180) <= not(layer5_outputs(1831));
    layer6_outputs(2181) <= not((layer5_outputs(239)) xor (layer5_outputs(2077)));
    layer6_outputs(2182) <= layer5_outputs(1308);
    layer6_outputs(2183) <= not((layer5_outputs(161)) xor (layer5_outputs(686)));
    layer6_outputs(2184) <= (layer5_outputs(2491)) or (layer5_outputs(972));
    layer6_outputs(2185) <= not(layer5_outputs(2417));
    layer6_outputs(2186) <= not((layer5_outputs(1455)) and (layer5_outputs(1032)));
    layer6_outputs(2187) <= not((layer5_outputs(2440)) and (layer5_outputs(1543)));
    layer6_outputs(2188) <= layer5_outputs(2488);
    layer6_outputs(2189) <= (layer5_outputs(650)) and not (layer5_outputs(629));
    layer6_outputs(2190) <= layer5_outputs(2531);
    layer6_outputs(2191) <= not(layer5_outputs(2513));
    layer6_outputs(2192) <= layer5_outputs(1314);
    layer6_outputs(2193) <= not(layer5_outputs(1351));
    layer6_outputs(2194) <= (layer5_outputs(1054)) and not (layer5_outputs(2511));
    layer6_outputs(2195) <= '1';
    layer6_outputs(2196) <= not(layer5_outputs(746));
    layer6_outputs(2197) <= '1';
    layer6_outputs(2198) <= layer5_outputs(2014);
    layer6_outputs(2199) <= not(layer5_outputs(520));
    layer6_outputs(2200) <= (layer5_outputs(2503)) and not (layer5_outputs(1550));
    layer6_outputs(2201) <= layer5_outputs(1560);
    layer6_outputs(2202) <= layer5_outputs(655);
    layer6_outputs(2203) <= layer5_outputs(320);
    layer6_outputs(2204) <= not(layer5_outputs(2281));
    layer6_outputs(2205) <= not(layer5_outputs(1119));
    layer6_outputs(2206) <= not(layer5_outputs(421));
    layer6_outputs(2207) <= layer5_outputs(333);
    layer6_outputs(2208) <= not(layer5_outputs(1844));
    layer6_outputs(2209) <= layer5_outputs(1281);
    layer6_outputs(2210) <= not(layer5_outputs(79));
    layer6_outputs(2211) <= layer5_outputs(458);
    layer6_outputs(2212) <= layer5_outputs(1030);
    layer6_outputs(2213) <= not(layer5_outputs(91));
    layer6_outputs(2214) <= not(layer5_outputs(1267)) or (layer5_outputs(1089));
    layer6_outputs(2215) <= (layer5_outputs(1986)) and (layer5_outputs(1509));
    layer6_outputs(2216) <= layer5_outputs(146);
    layer6_outputs(2217) <= (layer5_outputs(551)) and not (layer5_outputs(1013));
    layer6_outputs(2218) <= (layer5_outputs(286)) or (layer5_outputs(782));
    layer6_outputs(2219) <= not(layer5_outputs(1737)) or (layer5_outputs(303));
    layer6_outputs(2220) <= not(layer5_outputs(244));
    layer6_outputs(2221) <= (layer5_outputs(631)) and (layer5_outputs(663));
    layer6_outputs(2222) <= not(layer5_outputs(867)) or (layer5_outputs(1363));
    layer6_outputs(2223) <= (layer5_outputs(645)) and (layer5_outputs(2134));
    layer6_outputs(2224) <= layer5_outputs(2553);
    layer6_outputs(2225) <= not(layer5_outputs(850)) or (layer5_outputs(1815));
    layer6_outputs(2226) <= layer5_outputs(1139);
    layer6_outputs(2227) <= layer5_outputs(1919);
    layer6_outputs(2228) <= not((layer5_outputs(553)) and (layer5_outputs(1100)));
    layer6_outputs(2229) <= (layer5_outputs(1481)) and (layer5_outputs(625));
    layer6_outputs(2230) <= not(layer5_outputs(1900));
    layer6_outputs(2231) <= not(layer5_outputs(2395)) or (layer5_outputs(150));
    layer6_outputs(2232) <= (layer5_outputs(1346)) and not (layer5_outputs(96));
    layer6_outputs(2233) <= layer5_outputs(2368);
    layer6_outputs(2234) <= not(layer5_outputs(1093));
    layer6_outputs(2235) <= not(layer5_outputs(2148));
    layer6_outputs(2236) <= not((layer5_outputs(990)) or (layer5_outputs(2011)));
    layer6_outputs(2237) <= not(layer5_outputs(124));
    layer6_outputs(2238) <= not(layer5_outputs(2164));
    layer6_outputs(2239) <= not(layer5_outputs(1355));
    layer6_outputs(2240) <= not((layer5_outputs(1817)) or (layer5_outputs(2064)));
    layer6_outputs(2241) <= not(layer5_outputs(567));
    layer6_outputs(2242) <= (layer5_outputs(1737)) xor (layer5_outputs(830));
    layer6_outputs(2243) <= not((layer5_outputs(1318)) and (layer5_outputs(1990)));
    layer6_outputs(2244) <= not(layer5_outputs(1269));
    layer6_outputs(2245) <= not(layer5_outputs(308));
    layer6_outputs(2246) <= not((layer5_outputs(747)) and (layer5_outputs(1820)));
    layer6_outputs(2247) <= not(layer5_outputs(2154));
    layer6_outputs(2248) <= (layer5_outputs(767)) or (layer5_outputs(647));
    layer6_outputs(2249) <= '1';
    layer6_outputs(2250) <= (layer5_outputs(1077)) and (layer5_outputs(1998));
    layer6_outputs(2251) <= layer5_outputs(2087);
    layer6_outputs(2252) <= not(layer5_outputs(934));
    layer6_outputs(2253) <= not((layer5_outputs(1501)) and (layer5_outputs(1211)));
    layer6_outputs(2254) <= (layer5_outputs(1366)) and not (layer5_outputs(1144));
    layer6_outputs(2255) <= not(layer5_outputs(916));
    layer6_outputs(2256) <= not((layer5_outputs(2511)) and (layer5_outputs(188)));
    layer6_outputs(2257) <= (layer5_outputs(1900)) xor (layer5_outputs(2015));
    layer6_outputs(2258) <= layer5_outputs(1078);
    layer6_outputs(2259) <= not((layer5_outputs(854)) and (layer5_outputs(1171)));
    layer6_outputs(2260) <= not(layer5_outputs(1284));
    layer6_outputs(2261) <= layer5_outputs(514);
    layer6_outputs(2262) <= layer5_outputs(129);
    layer6_outputs(2263) <= (layer5_outputs(660)) or (layer5_outputs(2199));
    layer6_outputs(2264) <= layer5_outputs(4);
    layer6_outputs(2265) <= layer5_outputs(1227);
    layer6_outputs(2266) <= layer5_outputs(493);
    layer6_outputs(2267) <= not(layer5_outputs(1027));
    layer6_outputs(2268) <= layer5_outputs(230);
    layer6_outputs(2269) <= layer5_outputs(2429);
    layer6_outputs(2270) <= not(layer5_outputs(32));
    layer6_outputs(2271) <= layer5_outputs(1103);
    layer6_outputs(2272) <= not(layer5_outputs(1181)) or (layer5_outputs(932));
    layer6_outputs(2273) <= not(layer5_outputs(1335));
    layer6_outputs(2274) <= (layer5_outputs(136)) xor (layer5_outputs(1101));
    layer6_outputs(2275) <= not(layer5_outputs(883)) or (layer5_outputs(2215));
    layer6_outputs(2276) <= not((layer5_outputs(311)) and (layer5_outputs(70)));
    layer6_outputs(2277) <= not((layer5_outputs(1430)) xor (layer5_outputs(1171)));
    layer6_outputs(2278) <= (layer5_outputs(2434)) or (layer5_outputs(386));
    layer6_outputs(2279) <= not(layer5_outputs(137));
    layer6_outputs(2280) <= not(layer5_outputs(564));
    layer6_outputs(2281) <= '0';
    layer6_outputs(2282) <= not((layer5_outputs(2398)) and (layer5_outputs(1140)));
    layer6_outputs(2283) <= not(layer5_outputs(212));
    layer6_outputs(2284) <= (layer5_outputs(263)) xor (layer5_outputs(1340));
    layer6_outputs(2285) <= (layer5_outputs(778)) and not (layer5_outputs(961));
    layer6_outputs(2286) <= (layer5_outputs(95)) and (layer5_outputs(64));
    layer6_outputs(2287) <= layer5_outputs(228);
    layer6_outputs(2288) <= layer5_outputs(1947);
    layer6_outputs(2289) <= not((layer5_outputs(522)) xor (layer5_outputs(2166)));
    layer6_outputs(2290) <= (layer5_outputs(139)) xor (layer5_outputs(60));
    layer6_outputs(2291) <= not(layer5_outputs(2427));
    layer6_outputs(2292) <= not((layer5_outputs(893)) and (layer5_outputs(1754)));
    layer6_outputs(2293) <= (layer5_outputs(1472)) xor (layer5_outputs(774));
    layer6_outputs(2294) <= not(layer5_outputs(1538));
    layer6_outputs(2295) <= layer5_outputs(1084);
    layer6_outputs(2296) <= not((layer5_outputs(2037)) xor (layer5_outputs(2074)));
    layer6_outputs(2297) <= not(layer5_outputs(904)) or (layer5_outputs(2490));
    layer6_outputs(2298) <= not((layer5_outputs(84)) or (layer5_outputs(1502)));
    layer6_outputs(2299) <= not(layer5_outputs(2343));
    layer6_outputs(2300) <= layer5_outputs(211);
    layer6_outputs(2301) <= not((layer5_outputs(1364)) xor (layer5_outputs(2320)));
    layer6_outputs(2302) <= layer5_outputs(2441);
    layer6_outputs(2303) <= layer5_outputs(21);
    layer6_outputs(2304) <= (layer5_outputs(1798)) xor (layer5_outputs(1927));
    layer6_outputs(2305) <= not(layer5_outputs(1363)) or (layer5_outputs(1987));
    layer6_outputs(2306) <= layer5_outputs(837);
    layer6_outputs(2307) <= layer5_outputs(425);
    layer6_outputs(2308) <= not(layer5_outputs(1767));
    layer6_outputs(2309) <= layer5_outputs(736);
    layer6_outputs(2310) <= layer5_outputs(1296);
    layer6_outputs(2311) <= not(layer5_outputs(1559));
    layer6_outputs(2312) <= (layer5_outputs(2539)) xor (layer5_outputs(1424));
    layer6_outputs(2313) <= not(layer5_outputs(2264));
    layer6_outputs(2314) <= layer5_outputs(1112);
    layer6_outputs(2315) <= not((layer5_outputs(2458)) and (layer5_outputs(743)));
    layer6_outputs(2316) <= (layer5_outputs(2203)) and (layer5_outputs(1625));
    layer6_outputs(2317) <= (layer5_outputs(12)) and not (layer5_outputs(1497));
    layer6_outputs(2318) <= (layer5_outputs(78)) and not (layer5_outputs(1489));
    layer6_outputs(2319) <= not((layer5_outputs(465)) and (layer5_outputs(1960)));
    layer6_outputs(2320) <= '0';
    layer6_outputs(2321) <= (layer5_outputs(1621)) and not (layer5_outputs(1367));
    layer6_outputs(2322) <= (layer5_outputs(86)) and not (layer5_outputs(937));
    layer6_outputs(2323) <= not(layer5_outputs(430));
    layer6_outputs(2324) <= not(layer5_outputs(1931)) or (layer5_outputs(816));
    layer6_outputs(2325) <= not(layer5_outputs(2133));
    layer6_outputs(2326) <= not(layer5_outputs(2178));
    layer6_outputs(2327) <= layer5_outputs(2340);
    layer6_outputs(2328) <= (layer5_outputs(862)) and (layer5_outputs(217));
    layer6_outputs(2329) <= layer5_outputs(1488);
    layer6_outputs(2330) <= (layer5_outputs(1357)) xor (layer5_outputs(2076));
    layer6_outputs(2331) <= not((layer5_outputs(2270)) or (layer5_outputs(337)));
    layer6_outputs(2332) <= not(layer5_outputs(2127));
    layer6_outputs(2333) <= (layer5_outputs(1548)) or (layer5_outputs(231));
    layer6_outputs(2334) <= not(layer5_outputs(866)) or (layer5_outputs(216));
    layer6_outputs(2335) <= not(layer5_outputs(347));
    layer6_outputs(2336) <= (layer5_outputs(26)) and not (layer5_outputs(1922));
    layer6_outputs(2337) <= not(layer5_outputs(315));
    layer6_outputs(2338) <= not((layer5_outputs(2120)) xor (layer5_outputs(1394)));
    layer6_outputs(2339) <= not(layer5_outputs(2476));
    layer6_outputs(2340) <= not(layer5_outputs(1810));
    layer6_outputs(2341) <= layer5_outputs(419);
    layer6_outputs(2342) <= not(layer5_outputs(2267));
    layer6_outputs(2343) <= not(layer5_outputs(1770));
    layer6_outputs(2344) <= layer5_outputs(1207);
    layer6_outputs(2345) <= not((layer5_outputs(2068)) and (layer5_outputs(1179)));
    layer6_outputs(2346) <= (layer5_outputs(790)) and (layer5_outputs(643));
    layer6_outputs(2347) <= (layer5_outputs(2379)) xor (layer5_outputs(1793));
    layer6_outputs(2348) <= '1';
    layer6_outputs(2349) <= layer5_outputs(1918);
    layer6_outputs(2350) <= layer5_outputs(132);
    layer6_outputs(2351) <= not((layer5_outputs(1072)) xor (layer5_outputs(471)));
    layer6_outputs(2352) <= not(layer5_outputs(100));
    layer6_outputs(2353) <= not((layer5_outputs(2318)) and (layer5_outputs(2200)));
    layer6_outputs(2354) <= (layer5_outputs(833)) and not (layer5_outputs(757));
    layer6_outputs(2355) <= (layer5_outputs(1355)) and (layer5_outputs(977));
    layer6_outputs(2356) <= layer5_outputs(788);
    layer6_outputs(2357) <= not(layer5_outputs(1828));
    layer6_outputs(2358) <= not(layer5_outputs(657));
    layer6_outputs(2359) <= not((layer5_outputs(110)) or (layer5_outputs(1969)));
    layer6_outputs(2360) <= (layer5_outputs(1671)) and not (layer5_outputs(2027));
    layer6_outputs(2361) <= not(layer5_outputs(1609));
    layer6_outputs(2362) <= layer5_outputs(2376);
    layer6_outputs(2363) <= not((layer5_outputs(714)) or (layer5_outputs(1750)));
    layer6_outputs(2364) <= layer5_outputs(1515);
    layer6_outputs(2365) <= not(layer5_outputs(2278));
    layer6_outputs(2366) <= not(layer5_outputs(1645));
    layer6_outputs(2367) <= not(layer5_outputs(2168)) or (layer5_outputs(1607));
    layer6_outputs(2368) <= layer5_outputs(159);
    layer6_outputs(2369) <= not(layer5_outputs(1344));
    layer6_outputs(2370) <= not(layer5_outputs(234));
    layer6_outputs(2371) <= (layer5_outputs(2559)) xor (layer5_outputs(2512));
    layer6_outputs(2372) <= layer5_outputs(480);
    layer6_outputs(2373) <= not(layer5_outputs(1745));
    layer6_outputs(2374) <= not((layer5_outputs(762)) and (layer5_outputs(1111)));
    layer6_outputs(2375) <= '1';
    layer6_outputs(2376) <= layer5_outputs(1715);
    layer6_outputs(2377) <= (layer5_outputs(1133)) and (layer5_outputs(449));
    layer6_outputs(2378) <= not(layer5_outputs(1580)) or (layer5_outputs(438));
    layer6_outputs(2379) <= not((layer5_outputs(111)) xor (layer5_outputs(2233)));
    layer6_outputs(2380) <= layer5_outputs(420);
    layer6_outputs(2381) <= not((layer5_outputs(2050)) or (layer5_outputs(1946)));
    layer6_outputs(2382) <= (layer5_outputs(352)) and (layer5_outputs(2418));
    layer6_outputs(2383) <= not((layer5_outputs(2021)) or (layer5_outputs(1052)));
    layer6_outputs(2384) <= layer5_outputs(448);
    layer6_outputs(2385) <= not(layer5_outputs(2413));
    layer6_outputs(2386) <= (layer5_outputs(1430)) and (layer5_outputs(738));
    layer6_outputs(2387) <= not(layer5_outputs(1817));
    layer6_outputs(2388) <= not(layer5_outputs(534));
    layer6_outputs(2389) <= layer5_outputs(155);
    layer6_outputs(2390) <= not(layer5_outputs(2426)) or (layer5_outputs(393));
    layer6_outputs(2391) <= (layer5_outputs(2242)) xor (layer5_outputs(153));
    layer6_outputs(2392) <= (layer5_outputs(710)) and (layer5_outputs(1505));
    layer6_outputs(2393) <= not(layer5_outputs(1226));
    layer6_outputs(2394) <= not(layer5_outputs(845));
    layer6_outputs(2395) <= (layer5_outputs(2497)) xor (layer5_outputs(1409));
    layer6_outputs(2396) <= layer5_outputs(1248);
    layer6_outputs(2397) <= not((layer5_outputs(1249)) or (layer5_outputs(1530)));
    layer6_outputs(2398) <= (layer5_outputs(1389)) or (layer5_outputs(1200));
    layer6_outputs(2399) <= not((layer5_outputs(685)) and (layer5_outputs(1920)));
    layer6_outputs(2400) <= not(layer5_outputs(589)) or (layer5_outputs(368));
    layer6_outputs(2401) <= '1';
    layer6_outputs(2402) <= (layer5_outputs(359)) or (layer5_outputs(2250));
    layer6_outputs(2403) <= (layer5_outputs(381)) and not (layer5_outputs(730));
    layer6_outputs(2404) <= '0';
    layer6_outputs(2405) <= layer5_outputs(2202);
    layer6_outputs(2406) <= not(layer5_outputs(1858));
    layer6_outputs(2407) <= layer5_outputs(2382);
    layer6_outputs(2408) <= not(layer5_outputs(1150));
    layer6_outputs(2409) <= (layer5_outputs(926)) xor (layer5_outputs(1845));
    layer6_outputs(2410) <= layer5_outputs(861);
    layer6_outputs(2411) <= layer5_outputs(2406);
    layer6_outputs(2412) <= layer5_outputs(1788);
    layer6_outputs(2413) <= not(layer5_outputs(1190));
    layer6_outputs(2414) <= not((layer5_outputs(2217)) or (layer5_outputs(465)));
    layer6_outputs(2415) <= layer5_outputs(524);
    layer6_outputs(2416) <= layer5_outputs(2052);
    layer6_outputs(2417) <= (layer5_outputs(1466)) and (layer5_outputs(2358));
    layer6_outputs(2418) <= layer5_outputs(526);
    layer6_outputs(2419) <= (layer5_outputs(957)) and (layer5_outputs(751));
    layer6_outputs(2420) <= '1';
    layer6_outputs(2421) <= layer5_outputs(416);
    layer6_outputs(2422) <= not((layer5_outputs(1723)) xor (layer5_outputs(671)));
    layer6_outputs(2423) <= (layer5_outputs(288)) and (layer5_outputs(1711));
    layer6_outputs(2424) <= layer5_outputs(1419);
    layer6_outputs(2425) <= not(layer5_outputs(344));
    layer6_outputs(2426) <= (layer5_outputs(781)) xor (layer5_outputs(2393));
    layer6_outputs(2427) <= layer5_outputs(1162);
    layer6_outputs(2428) <= (layer5_outputs(1952)) and not (layer5_outputs(1618));
    layer6_outputs(2429) <= not(layer5_outputs(2231));
    layer6_outputs(2430) <= not((layer5_outputs(2526)) xor (layer5_outputs(516)));
    layer6_outputs(2431) <= layer5_outputs(2207);
    layer6_outputs(2432) <= (layer5_outputs(1014)) or (layer5_outputs(1324));
    layer6_outputs(2433) <= not(layer5_outputs(1687));
    layer6_outputs(2434) <= not(layer5_outputs(67));
    layer6_outputs(2435) <= not(layer5_outputs(2029));
    layer6_outputs(2436) <= (layer5_outputs(2311)) and not (layer5_outputs(1317));
    layer6_outputs(2437) <= (layer5_outputs(195)) and (layer5_outputs(1605));
    layer6_outputs(2438) <= (layer5_outputs(1692)) and not (layer5_outputs(235));
    layer6_outputs(2439) <= not(layer5_outputs(1158));
    layer6_outputs(2440) <= not(layer5_outputs(532)) or (layer5_outputs(2119));
    layer6_outputs(2441) <= not(layer5_outputs(1556));
    layer6_outputs(2442) <= not(layer5_outputs(2042));
    layer6_outputs(2443) <= not(layer5_outputs(963)) or (layer5_outputs(1304));
    layer6_outputs(2444) <= not((layer5_outputs(1164)) xor (layer5_outputs(1205)));
    layer6_outputs(2445) <= layer5_outputs(2263);
    layer6_outputs(2446) <= layer5_outputs(785);
    layer6_outputs(2447) <= layer5_outputs(907);
    layer6_outputs(2448) <= not((layer5_outputs(1093)) and (layer5_outputs(2492)));
    layer6_outputs(2449) <= not((layer5_outputs(737)) and (layer5_outputs(841)));
    layer6_outputs(2450) <= not(layer5_outputs(1417)) or (layer5_outputs(1405));
    layer6_outputs(2451) <= not(layer5_outputs(459)) or (layer5_outputs(968));
    layer6_outputs(2452) <= layer5_outputs(1831);
    layer6_outputs(2453) <= layer5_outputs(1602);
    layer6_outputs(2454) <= not(layer5_outputs(1377)) or (layer5_outputs(173));
    layer6_outputs(2455) <= layer5_outputs(1282);
    layer6_outputs(2456) <= not(layer5_outputs(58));
    layer6_outputs(2457) <= '0';
    layer6_outputs(2458) <= not(layer5_outputs(2393)) or (layer5_outputs(1583));
    layer6_outputs(2459) <= (layer5_outputs(1114)) or (layer5_outputs(2164));
    layer6_outputs(2460) <= layer5_outputs(2153);
    layer6_outputs(2461) <= not((layer5_outputs(55)) xor (layer5_outputs(2318)));
    layer6_outputs(2462) <= layer5_outputs(1238);
    layer6_outputs(2463) <= layer5_outputs(1152);
    layer6_outputs(2464) <= not((layer5_outputs(2083)) and (layer5_outputs(1175)));
    layer6_outputs(2465) <= not(layer5_outputs(2261));
    layer6_outputs(2466) <= layer5_outputs(39);
    layer6_outputs(2467) <= not((layer5_outputs(1126)) or (layer5_outputs(104)));
    layer6_outputs(2468) <= layer5_outputs(2403);
    layer6_outputs(2469) <= (layer5_outputs(1373)) and (layer5_outputs(1336));
    layer6_outputs(2470) <= (layer5_outputs(1592)) xor (layer5_outputs(537));
    layer6_outputs(2471) <= not(layer5_outputs(346));
    layer6_outputs(2472) <= not((layer5_outputs(123)) xor (layer5_outputs(760)));
    layer6_outputs(2473) <= layer5_outputs(2306);
    layer6_outputs(2474) <= not(layer5_outputs(786));
    layer6_outputs(2475) <= (layer5_outputs(1662)) xor (layer5_outputs(903));
    layer6_outputs(2476) <= not(layer5_outputs(2139)) or (layer5_outputs(992));
    layer6_outputs(2477) <= layer5_outputs(1016);
    layer6_outputs(2478) <= layer5_outputs(1524);
    layer6_outputs(2479) <= layer5_outputs(2031);
    layer6_outputs(2480) <= not(layer5_outputs(1505));
    layer6_outputs(2481) <= not(layer5_outputs(2526));
    layer6_outputs(2482) <= not(layer5_outputs(1694));
    layer6_outputs(2483) <= (layer5_outputs(341)) or (layer5_outputs(1499));
    layer6_outputs(2484) <= layer5_outputs(583);
    layer6_outputs(2485) <= layer5_outputs(488);
    layer6_outputs(2486) <= not(layer5_outputs(1975));
    layer6_outputs(2487) <= (layer5_outputs(431)) xor (layer5_outputs(371));
    layer6_outputs(2488) <= layer5_outputs(927);
    layer6_outputs(2489) <= not(layer5_outputs(229));
    layer6_outputs(2490) <= not(layer5_outputs(2362));
    layer6_outputs(2491) <= (layer5_outputs(2086)) xor (layer5_outputs(1129));
    layer6_outputs(2492) <= layer5_outputs(2291);
    layer6_outputs(2493) <= not(layer5_outputs(2423)) or (layer5_outputs(2102));
    layer6_outputs(2494) <= not(layer5_outputs(1594));
    layer6_outputs(2495) <= not(layer5_outputs(1638)) or (layer5_outputs(264));
    layer6_outputs(2496) <= not(layer5_outputs(2139)) or (layer5_outputs(1991));
    layer6_outputs(2497) <= '1';
    layer6_outputs(2498) <= (layer5_outputs(342)) and not (layer5_outputs(1044));
    layer6_outputs(2499) <= (layer5_outputs(2046)) and not (layer5_outputs(680));
    layer6_outputs(2500) <= not(layer5_outputs(42));
    layer6_outputs(2501) <= not(layer5_outputs(2252));
    layer6_outputs(2502) <= layer5_outputs(321);
    layer6_outputs(2503) <= layer5_outputs(2394);
    layer6_outputs(2504) <= (layer5_outputs(1635)) and not (layer5_outputs(2533));
    layer6_outputs(2505) <= not(layer5_outputs(1186));
    layer6_outputs(2506) <= not(layer5_outputs(518));
    layer6_outputs(2507) <= layer5_outputs(185);
    layer6_outputs(2508) <= not((layer5_outputs(925)) xor (layer5_outputs(1816)));
    layer6_outputs(2509) <= layer5_outputs(260);
    layer6_outputs(2510) <= layer5_outputs(1617);
    layer6_outputs(2511) <= not((layer5_outputs(2138)) and (layer5_outputs(73)));
    layer6_outputs(2512) <= (layer5_outputs(302)) and not (layer5_outputs(858));
    layer6_outputs(2513) <= not(layer5_outputs(2472)) or (layer5_outputs(955));
    layer6_outputs(2514) <= not(layer5_outputs(2294));
    layer6_outputs(2515) <= not(layer5_outputs(223));
    layer6_outputs(2516) <= (layer5_outputs(2246)) and not (layer5_outputs(1801));
    layer6_outputs(2517) <= not(layer5_outputs(1647));
    layer6_outputs(2518) <= not(layer5_outputs(423));
    layer6_outputs(2519) <= not(layer5_outputs(239));
    layer6_outputs(2520) <= (layer5_outputs(1767)) and not (layer5_outputs(1144));
    layer6_outputs(2521) <= layer5_outputs(1790);
    layer6_outputs(2522) <= not(layer5_outputs(2049));
    layer6_outputs(2523) <= (layer5_outputs(651)) and not (layer5_outputs(1710));
    layer6_outputs(2524) <= not(layer5_outputs(2307));
    layer6_outputs(2525) <= not(layer5_outputs(762)) or (layer5_outputs(2302));
    layer6_outputs(2526) <= not(layer5_outputs(1541)) or (layer5_outputs(1870));
    layer6_outputs(2527) <= (layer5_outputs(2322)) or (layer5_outputs(412));
    layer6_outputs(2528) <= not((layer5_outputs(574)) or (layer5_outputs(661)));
    layer6_outputs(2529) <= (layer5_outputs(1366)) and not (layer5_outputs(2493));
    layer6_outputs(2530) <= not(layer5_outputs(778));
    layer6_outputs(2531) <= not(layer5_outputs(1639));
    layer6_outputs(2532) <= not(layer5_outputs(1476));
    layer6_outputs(2533) <= layer5_outputs(186);
    layer6_outputs(2534) <= not(layer5_outputs(525));
    layer6_outputs(2535) <= layer5_outputs(1333);
    layer6_outputs(2536) <= not((layer5_outputs(1428)) xor (layer5_outputs(1104)));
    layer6_outputs(2537) <= not((layer5_outputs(1029)) xor (layer5_outputs(929)));
    layer6_outputs(2538) <= (layer5_outputs(952)) or (layer5_outputs(1141));
    layer6_outputs(2539) <= not(layer5_outputs(982));
    layer6_outputs(2540) <= not((layer5_outputs(780)) or (layer5_outputs(170)));
    layer6_outputs(2541) <= not(layer5_outputs(591));
    layer6_outputs(2542) <= layer5_outputs(2225);
    layer6_outputs(2543) <= (layer5_outputs(2002)) or (layer5_outputs(1979));
    layer6_outputs(2544) <= not(layer5_outputs(1910));
    layer6_outputs(2545) <= not(layer5_outputs(441));
    layer6_outputs(2546) <= not((layer5_outputs(749)) or (layer5_outputs(2387)));
    layer6_outputs(2547) <= (layer5_outputs(1493)) and not (layer5_outputs(1213));
    layer6_outputs(2548) <= not(layer5_outputs(1587)) or (layer5_outputs(1069));
    layer6_outputs(2549) <= not((layer5_outputs(1438)) and (layer5_outputs(441)));
    layer6_outputs(2550) <= not(layer5_outputs(1208));
    layer6_outputs(2551) <= not(layer5_outputs(283));
    layer6_outputs(2552) <= (layer5_outputs(1828)) and (layer5_outputs(1942));
    layer6_outputs(2553) <= not((layer5_outputs(510)) xor (layer5_outputs(1616)));
    layer6_outputs(2554) <= not(layer5_outputs(2439));
    layer6_outputs(2555) <= layer5_outputs(1520);
    layer6_outputs(2556) <= not(layer5_outputs(330));
    layer6_outputs(2557) <= layer5_outputs(303);
    layer6_outputs(2558) <= layer5_outputs(2247);
    layer6_outputs(2559) <= not(layer5_outputs(2185)) or (layer5_outputs(950));
    outputs(0) <= not(layer6_outputs(105));
    outputs(1) <= (layer6_outputs(1595)) and not (layer6_outputs(2403));
    outputs(2) <= (layer6_outputs(443)) and not (layer6_outputs(2523));
    outputs(3) <= not(layer6_outputs(2));
    outputs(4) <= layer6_outputs(1903);
    outputs(5) <= (layer6_outputs(1614)) xor (layer6_outputs(1549));
    outputs(6) <= not(layer6_outputs(2462));
    outputs(7) <= not(layer6_outputs(1447));
    outputs(8) <= not(layer6_outputs(165));
    outputs(9) <= not(layer6_outputs(312)) or (layer6_outputs(2392));
    outputs(10) <= (layer6_outputs(1534)) or (layer6_outputs(42));
    outputs(11) <= not(layer6_outputs(1696));
    outputs(12) <= layer6_outputs(1190);
    outputs(13) <= (layer6_outputs(696)) and (layer6_outputs(1354));
    outputs(14) <= not(layer6_outputs(1268));
    outputs(15) <= not((layer6_outputs(2093)) or (layer6_outputs(464)));
    outputs(16) <= not((layer6_outputs(550)) or (layer6_outputs(236)));
    outputs(17) <= (layer6_outputs(1180)) and not (layer6_outputs(2041));
    outputs(18) <= layer6_outputs(638);
    outputs(19) <= not((layer6_outputs(1292)) or (layer6_outputs(803)));
    outputs(20) <= (layer6_outputs(1201)) and not (layer6_outputs(265));
    outputs(21) <= not(layer6_outputs(2282)) or (layer6_outputs(1056));
    outputs(22) <= (layer6_outputs(2280)) and (layer6_outputs(72));
    outputs(23) <= not((layer6_outputs(145)) xor (layer6_outputs(1526)));
    outputs(24) <= layer6_outputs(2356);
    outputs(25) <= not(layer6_outputs(2468));
    outputs(26) <= (layer6_outputs(1508)) xor (layer6_outputs(2496));
    outputs(27) <= not((layer6_outputs(1133)) or (layer6_outputs(224)));
    outputs(28) <= layer6_outputs(161);
    outputs(29) <= layer6_outputs(940);
    outputs(30) <= (layer6_outputs(869)) and not (layer6_outputs(1668));
    outputs(31) <= not((layer6_outputs(1663)) or (layer6_outputs(662)));
    outputs(32) <= (layer6_outputs(1958)) xor (layer6_outputs(2338));
    outputs(33) <= (layer6_outputs(750)) and not (layer6_outputs(2219));
    outputs(34) <= not(layer6_outputs(567));
    outputs(35) <= layer6_outputs(2224);
    outputs(36) <= not(layer6_outputs(2017)) or (layer6_outputs(921));
    outputs(37) <= (layer6_outputs(1632)) and not (layer6_outputs(686));
    outputs(38) <= layer6_outputs(1670);
    outputs(39) <= layer6_outputs(295);
    outputs(40) <= not(layer6_outputs(460));
    outputs(41) <= not(layer6_outputs(1392));
    outputs(42) <= not((layer6_outputs(2006)) or (layer6_outputs(1502)));
    outputs(43) <= not(layer6_outputs(534));
    outputs(44) <= not(layer6_outputs(238));
    outputs(45) <= layer6_outputs(73);
    outputs(46) <= layer6_outputs(1818);
    outputs(47) <= (layer6_outputs(2483)) and not (layer6_outputs(1138));
    outputs(48) <= not(layer6_outputs(1686));
    outputs(49) <= layer6_outputs(1039);
    outputs(50) <= not(layer6_outputs(1043));
    outputs(51) <= (layer6_outputs(600)) and (layer6_outputs(2181));
    outputs(52) <= not(layer6_outputs(286));
    outputs(53) <= (layer6_outputs(930)) and not (layer6_outputs(2358));
    outputs(54) <= not((layer6_outputs(2482)) or (layer6_outputs(490)));
    outputs(55) <= not(layer6_outputs(1686));
    outputs(56) <= (layer6_outputs(571)) and (layer6_outputs(1295));
    outputs(57) <= not(layer6_outputs(1121));
    outputs(58) <= not(layer6_outputs(875));
    outputs(59) <= not(layer6_outputs(1480)) or (layer6_outputs(1208));
    outputs(60) <= layer6_outputs(1957);
    outputs(61) <= not(layer6_outputs(1694));
    outputs(62) <= layer6_outputs(2018);
    outputs(63) <= not(layer6_outputs(729));
    outputs(64) <= not(layer6_outputs(1092));
    outputs(65) <= layer6_outputs(48);
    outputs(66) <= not(layer6_outputs(2079));
    outputs(67) <= (layer6_outputs(1374)) and not (layer6_outputs(1864));
    outputs(68) <= not(layer6_outputs(653));
    outputs(69) <= not(layer6_outputs(2408));
    outputs(70) <= layer6_outputs(2410);
    outputs(71) <= not(layer6_outputs(362));
    outputs(72) <= not((layer6_outputs(1397)) or (layer6_outputs(1646)));
    outputs(73) <= (layer6_outputs(67)) and not (layer6_outputs(1827));
    outputs(74) <= not((layer6_outputs(1768)) or (layer6_outputs(2000)));
    outputs(75) <= not(layer6_outputs(1430)) or (layer6_outputs(1940));
    outputs(76) <= layer6_outputs(63);
    outputs(77) <= not(layer6_outputs(32));
    outputs(78) <= (layer6_outputs(1755)) xor (layer6_outputs(2230));
    outputs(79) <= not(layer6_outputs(1924));
    outputs(80) <= not(layer6_outputs(24)) or (layer6_outputs(1142));
    outputs(81) <= layer6_outputs(647);
    outputs(82) <= not(layer6_outputs(1044));
    outputs(83) <= layer6_outputs(558);
    outputs(84) <= not(layer6_outputs(1467));
    outputs(85) <= not(layer6_outputs(1747));
    outputs(86) <= (layer6_outputs(5)) xor (layer6_outputs(2453));
    outputs(87) <= not(layer6_outputs(1851));
    outputs(88) <= not((layer6_outputs(1784)) or (layer6_outputs(402)));
    outputs(89) <= not(layer6_outputs(1457));
    outputs(90) <= (layer6_outputs(792)) xor (layer6_outputs(2515));
    outputs(91) <= not(layer6_outputs(1967));
    outputs(92) <= (layer6_outputs(2466)) xor (layer6_outputs(1207));
    outputs(93) <= not(layer6_outputs(112));
    outputs(94) <= layer6_outputs(1882);
    outputs(95) <= layer6_outputs(930);
    outputs(96) <= (layer6_outputs(2367)) and not (layer6_outputs(1322));
    outputs(97) <= not(layer6_outputs(2343));
    outputs(98) <= (layer6_outputs(2457)) xor (layer6_outputs(1256));
    outputs(99) <= (layer6_outputs(308)) and (layer6_outputs(773));
    outputs(100) <= layer6_outputs(2537);
    outputs(101) <= not((layer6_outputs(511)) or (layer6_outputs(2066)));
    outputs(102) <= not(layer6_outputs(706));
    outputs(103) <= layer6_outputs(1987);
    outputs(104) <= (layer6_outputs(1200)) and not (layer6_outputs(1403));
    outputs(105) <= layer6_outputs(1129);
    outputs(106) <= not(layer6_outputs(9));
    outputs(107) <= (layer6_outputs(2232)) xor (layer6_outputs(1365));
    outputs(108) <= not(layer6_outputs(2460));
    outputs(109) <= not(layer6_outputs(527));
    outputs(110) <= (layer6_outputs(1109)) or (layer6_outputs(1358));
    outputs(111) <= not(layer6_outputs(982));
    outputs(112) <= not(layer6_outputs(922));
    outputs(113) <= not(layer6_outputs(897));
    outputs(114) <= (layer6_outputs(984)) and not (layer6_outputs(1289));
    outputs(115) <= layer6_outputs(2446);
    outputs(116) <= (layer6_outputs(1417)) and not (layer6_outputs(53));
    outputs(117) <= (layer6_outputs(1825)) and not (layer6_outputs(1531));
    outputs(118) <= layer6_outputs(491);
    outputs(119) <= layer6_outputs(2137);
    outputs(120) <= layer6_outputs(2470);
    outputs(121) <= (layer6_outputs(1580)) xor (layer6_outputs(162));
    outputs(122) <= (layer6_outputs(992)) and (layer6_outputs(537));
    outputs(123) <= not((layer6_outputs(1443)) xor (layer6_outputs(1847)));
    outputs(124) <= not(layer6_outputs(216));
    outputs(125) <= not(layer6_outputs(530));
    outputs(126) <= (layer6_outputs(1779)) and (layer6_outputs(1255));
    outputs(127) <= not(layer6_outputs(337));
    outputs(128) <= not(layer6_outputs(1922));
    outputs(129) <= not((layer6_outputs(1742)) xor (layer6_outputs(2220)));
    outputs(130) <= (layer6_outputs(433)) xor (layer6_outputs(1917));
    outputs(131) <= (layer6_outputs(1937)) and (layer6_outputs(720));
    outputs(132) <= (layer6_outputs(2559)) and not (layer6_outputs(1835));
    outputs(133) <= not(layer6_outputs(956));
    outputs(134) <= layer6_outputs(1500);
    outputs(135) <= not(layer6_outputs(117));
    outputs(136) <= (layer6_outputs(206)) xor (layer6_outputs(1878));
    outputs(137) <= layer6_outputs(1488);
    outputs(138) <= not(layer6_outputs(1193));
    outputs(139) <= (layer6_outputs(1613)) and (layer6_outputs(819));
    outputs(140) <= layer6_outputs(2223);
    outputs(141) <= not(layer6_outputs(587));
    outputs(142) <= not(layer6_outputs(1267));
    outputs(143) <= (layer6_outputs(750)) and not (layer6_outputs(555));
    outputs(144) <= layer6_outputs(2279);
    outputs(145) <= layer6_outputs(1089);
    outputs(146) <= layer6_outputs(173);
    outputs(147) <= (layer6_outputs(738)) and not (layer6_outputs(77));
    outputs(148) <= (layer6_outputs(2167)) and (layer6_outputs(1512));
    outputs(149) <= not(layer6_outputs(2183));
    outputs(150) <= layer6_outputs(2417);
    outputs(151) <= layer6_outputs(1423);
    outputs(152) <= not(layer6_outputs(1991)) or (layer6_outputs(538));
    outputs(153) <= (layer6_outputs(2413)) and (layer6_outputs(911));
    outputs(154) <= not((layer6_outputs(1168)) xor (layer6_outputs(1239)));
    outputs(155) <= layer6_outputs(219);
    outputs(156) <= not((layer6_outputs(1666)) or (layer6_outputs(2523)));
    outputs(157) <= layer6_outputs(1636);
    outputs(158) <= (layer6_outputs(1157)) xor (layer6_outputs(2397));
    outputs(159) <= not(layer6_outputs(1216));
    outputs(160) <= layer6_outputs(2004);
    outputs(161) <= (layer6_outputs(1488)) and not (layer6_outputs(1970));
    outputs(162) <= layer6_outputs(536);
    outputs(163) <= layer6_outputs(860);
    outputs(164) <= not(layer6_outputs(1185));
    outputs(165) <= (layer6_outputs(1209)) and not (layer6_outputs(1336));
    outputs(166) <= layer6_outputs(1359);
    outputs(167) <= not(layer6_outputs(912));
    outputs(168) <= not(layer6_outputs(313));
    outputs(169) <= layer6_outputs(74);
    outputs(170) <= not(layer6_outputs(2312));
    outputs(171) <= not(layer6_outputs(1437));
    outputs(172) <= not((layer6_outputs(2496)) xor (layer6_outputs(894)));
    outputs(173) <= layer6_outputs(1569);
    outputs(174) <= layer6_outputs(505);
    outputs(175) <= (layer6_outputs(2331)) and not (layer6_outputs(2188));
    outputs(176) <= (layer6_outputs(1068)) and (layer6_outputs(2484));
    outputs(177) <= not((layer6_outputs(2110)) or (layer6_outputs(694)));
    outputs(178) <= not(layer6_outputs(1838));
    outputs(179) <= not(layer6_outputs(279));
    outputs(180) <= not(layer6_outputs(1710));
    outputs(181) <= layer6_outputs(2524);
    outputs(182) <= layer6_outputs(342);
    outputs(183) <= not((layer6_outputs(959)) xor (layer6_outputs(1941)));
    outputs(184) <= not(layer6_outputs(2262));
    outputs(185) <= not(layer6_outputs(1499)) or (layer6_outputs(890));
    outputs(186) <= layer6_outputs(176);
    outputs(187) <= (layer6_outputs(111)) and not (layer6_outputs(1600));
    outputs(188) <= (layer6_outputs(1294)) and not (layer6_outputs(142));
    outputs(189) <= not((layer6_outputs(169)) or (layer6_outputs(550)));
    outputs(190) <= layer6_outputs(633);
    outputs(191) <= layer6_outputs(1192);
    outputs(192) <= not(layer6_outputs(831));
    outputs(193) <= not(layer6_outputs(1084)) or (layer6_outputs(275));
    outputs(194) <= not(layer6_outputs(1627));
    outputs(195) <= not(layer6_outputs(1333));
    outputs(196) <= (layer6_outputs(1378)) and (layer6_outputs(1840));
    outputs(197) <= layer6_outputs(1658);
    outputs(198) <= layer6_outputs(1007);
    outputs(199) <= (layer6_outputs(2314)) and not (layer6_outputs(2283));
    outputs(200) <= (layer6_outputs(2055)) and (layer6_outputs(2543));
    outputs(201) <= not((layer6_outputs(2238)) xor (layer6_outputs(1764)));
    outputs(202) <= not(layer6_outputs(1446));
    outputs(203) <= not(layer6_outputs(2127));
    outputs(204) <= layer6_outputs(1752);
    outputs(205) <= layer6_outputs(61);
    outputs(206) <= layer6_outputs(590);
    outputs(207) <= not(layer6_outputs(55)) or (layer6_outputs(1682));
    outputs(208) <= (layer6_outputs(2444)) and not (layer6_outputs(428));
    outputs(209) <= not(layer6_outputs(1918));
    outputs(210) <= not(layer6_outputs(1662));
    outputs(211) <= layer6_outputs(891);
    outputs(212) <= not((layer6_outputs(1764)) or (layer6_outputs(2552)));
    outputs(213) <= not(layer6_outputs(322));
    outputs(214) <= not(layer6_outputs(591));
    outputs(215) <= layer6_outputs(1494);
    outputs(216) <= not(layer6_outputs(1045));
    outputs(217) <= (layer6_outputs(355)) and not (layer6_outputs(846));
    outputs(218) <= (layer6_outputs(1731)) and not (layer6_outputs(1104));
    outputs(219) <= layer6_outputs(2064);
    outputs(220) <= layer6_outputs(1952);
    outputs(221) <= (layer6_outputs(46)) xor (layer6_outputs(829));
    outputs(222) <= (layer6_outputs(119)) xor (layer6_outputs(1390));
    outputs(223) <= not((layer6_outputs(2340)) xor (layer6_outputs(1362)));
    outputs(224) <= not(layer6_outputs(1583));
    outputs(225) <= (layer6_outputs(1795)) and (layer6_outputs(1602));
    outputs(226) <= layer6_outputs(2331);
    outputs(227) <= not(layer6_outputs(1280));
    outputs(228) <= not(layer6_outputs(2228));
    outputs(229) <= (layer6_outputs(1971)) xor (layer6_outputs(1992));
    outputs(230) <= not((layer6_outputs(1047)) or (layer6_outputs(2106)));
    outputs(231) <= not(layer6_outputs(788));
    outputs(232) <= layer6_outputs(626);
    outputs(233) <= not(layer6_outputs(1527));
    outputs(234) <= layer6_outputs(1895);
    outputs(235) <= layer6_outputs(997);
    outputs(236) <= (layer6_outputs(2348)) and not (layer6_outputs(1261));
    outputs(237) <= layer6_outputs(1677);
    outputs(238) <= layer6_outputs(1705);
    outputs(239) <= layer6_outputs(2302);
    outputs(240) <= not(layer6_outputs(2350));
    outputs(241) <= layer6_outputs(938);
    outputs(242) <= layer6_outputs(795);
    outputs(243) <= not(layer6_outputs(1113));
    outputs(244) <= (layer6_outputs(2180)) and (layer6_outputs(125));
    outputs(245) <= not(layer6_outputs(1456));
    outputs(246) <= not(layer6_outputs(1015));
    outputs(247) <= not((layer6_outputs(154)) xor (layer6_outputs(735)));
    outputs(248) <= not(layer6_outputs(1223));
    outputs(249) <= layer6_outputs(2028);
    outputs(250) <= not(layer6_outputs(794));
    outputs(251) <= (layer6_outputs(1573)) and not (layer6_outputs(448));
    outputs(252) <= layer6_outputs(1340);
    outputs(253) <= not(layer6_outputs(413));
    outputs(254) <= not(layer6_outputs(1738));
    outputs(255) <= not(layer6_outputs(1769));
    outputs(256) <= not(layer6_outputs(611));
    outputs(257) <= layer6_outputs(2475);
    outputs(258) <= layer6_outputs(1230);
    outputs(259) <= not(layer6_outputs(1331));
    outputs(260) <= not((layer6_outputs(298)) xor (layer6_outputs(1930)));
    outputs(261) <= not(layer6_outputs(2103));
    outputs(262) <= not(layer6_outputs(235));
    outputs(263) <= layer6_outputs(2026);
    outputs(264) <= layer6_outputs(1850);
    outputs(265) <= not(layer6_outputs(1969));
    outputs(266) <= not(layer6_outputs(870));
    outputs(267) <= (layer6_outputs(2114)) and not (layer6_outputs(1054));
    outputs(268) <= layer6_outputs(1328);
    outputs(269) <= not((layer6_outputs(2489)) or (layer6_outputs(1534)));
    outputs(270) <= not(layer6_outputs(862));
    outputs(271) <= layer6_outputs(985);
    outputs(272) <= not(layer6_outputs(1803));
    outputs(273) <= (layer6_outputs(382)) and not (layer6_outputs(295));
    outputs(274) <= (layer6_outputs(2286)) and not (layer6_outputs(1188));
    outputs(275) <= not((layer6_outputs(1772)) xor (layer6_outputs(2028)));
    outputs(276) <= layer6_outputs(1246);
    outputs(277) <= (layer6_outputs(560)) and not (layer6_outputs(2266));
    outputs(278) <= not((layer6_outputs(619)) or (layer6_outputs(2252)));
    outputs(279) <= not((layer6_outputs(376)) xor (layer6_outputs(201)));
    outputs(280) <= not(layer6_outputs(28));
    outputs(281) <= (layer6_outputs(473)) and not (layer6_outputs(797));
    outputs(282) <= (layer6_outputs(462)) and not (layer6_outputs(616));
    outputs(283) <= not(layer6_outputs(1098));
    outputs(284) <= (layer6_outputs(357)) xor (layer6_outputs(1150));
    outputs(285) <= (layer6_outputs(2059)) and not (layer6_outputs(2513));
    outputs(286) <= (layer6_outputs(2091)) and (layer6_outputs(1853));
    outputs(287) <= not(layer6_outputs(702));
    outputs(288) <= (layer6_outputs(1540)) and not (layer6_outputs(2454));
    outputs(289) <= layer6_outputs(401);
    outputs(290) <= (layer6_outputs(1614)) and not (layer6_outputs(1003));
    outputs(291) <= (layer6_outputs(1083)) and (layer6_outputs(242));
    outputs(292) <= not(layer6_outputs(1071));
    outputs(293) <= layer6_outputs(2024);
    outputs(294) <= layer6_outputs(2317);
    outputs(295) <= layer6_outputs(972);
    outputs(296) <= (layer6_outputs(1282)) xor (layer6_outputs(1761));
    outputs(297) <= (layer6_outputs(177)) and not (layer6_outputs(252));
    outputs(298) <= not(layer6_outputs(1753));
    outputs(299) <= (layer6_outputs(1182)) and (layer6_outputs(12));
    outputs(300) <= (layer6_outputs(763)) xor (layer6_outputs(1076));
    outputs(301) <= not(layer6_outputs(707));
    outputs(302) <= (layer6_outputs(1678)) and not (layer6_outputs(1090));
    outputs(303) <= layer6_outputs(1510);
    outputs(304) <= layer6_outputs(2430);
    outputs(305) <= (layer6_outputs(480)) and not (layer6_outputs(1010));
    outputs(306) <= not(layer6_outputs(1993));
    outputs(307) <= not(layer6_outputs(515));
    outputs(308) <= not((layer6_outputs(170)) or (layer6_outputs(2109)));
    outputs(309) <= not(layer6_outputs(784));
    outputs(310) <= (layer6_outputs(2548)) and not (layer6_outputs(1599));
    outputs(311) <= not(layer6_outputs(1140));
    outputs(312) <= (layer6_outputs(915)) and not (layer6_outputs(1139));
    outputs(313) <= (layer6_outputs(617)) or (layer6_outputs(1141));
    outputs(314) <= (layer6_outputs(1496)) or (layer6_outputs(2200));
    outputs(315) <= layer6_outputs(239);
    outputs(316) <= (layer6_outputs(381)) and not (layer6_outputs(1990));
    outputs(317) <= (layer6_outputs(1788)) and not (layer6_outputs(417));
    outputs(318) <= layer6_outputs(2089);
    outputs(319) <= not(layer6_outputs(2484));
    outputs(320) <= (layer6_outputs(754)) and not (layer6_outputs(2120));
    outputs(321) <= not(layer6_outputs(1005));
    outputs(322) <= layer6_outputs(370);
    outputs(323) <= layer6_outputs(1360);
    outputs(324) <= layer6_outputs(1033);
    outputs(325) <= not((layer6_outputs(946)) or (layer6_outputs(2118)));
    outputs(326) <= not(layer6_outputs(2541));
    outputs(327) <= layer6_outputs(2386);
    outputs(328) <= not(layer6_outputs(1655));
    outputs(329) <= (layer6_outputs(160)) and not (layer6_outputs(1293));
    outputs(330) <= (layer6_outputs(675)) and not (layer6_outputs(283));
    outputs(331) <= not(layer6_outputs(2190)) or (layer6_outputs(239));
    outputs(332) <= (layer6_outputs(168)) and not (layer6_outputs(2365));
    outputs(333) <= layer6_outputs(2248);
    outputs(334) <= (layer6_outputs(1349)) and not (layer6_outputs(1371));
    outputs(335) <= not((layer6_outputs(1717)) xor (layer6_outputs(1267)));
    outputs(336) <= not(layer6_outputs(1021));
    outputs(337) <= layer6_outputs(2142);
    outputs(338) <= (layer6_outputs(382)) and not (layer6_outputs(699));
    outputs(339) <= (layer6_outputs(1948)) and (layer6_outputs(2512));
    outputs(340) <= layer6_outputs(1862);
    outputs(341) <= not((layer6_outputs(2386)) xor (layer6_outputs(2196)));
    outputs(342) <= (layer6_outputs(2209)) and not (layer6_outputs(1796));
    outputs(343) <= not((layer6_outputs(1323)) xor (layer6_outputs(2546)));
    outputs(344) <= (layer6_outputs(978)) and (layer6_outputs(227));
    outputs(345) <= (layer6_outputs(2089)) and not (layer6_outputs(2418));
    outputs(346) <= layer6_outputs(1061);
    outputs(347) <= not(layer6_outputs(707));
    outputs(348) <= not(layer6_outputs(415));
    outputs(349) <= not(layer6_outputs(1684));
    outputs(350) <= not(layer6_outputs(1116));
    outputs(351) <= (layer6_outputs(1961)) xor (layer6_outputs(592));
    outputs(352) <= not(layer6_outputs(1023));
    outputs(353) <= not(layer6_outputs(1184));
    outputs(354) <= layer6_outputs(1292);
    outputs(355) <= not(layer6_outputs(317));
    outputs(356) <= not((layer6_outputs(1012)) xor (layer6_outputs(2260)));
    outputs(357) <= layer6_outputs(546);
    outputs(358) <= not(layer6_outputs(2514));
    outputs(359) <= (layer6_outputs(1101)) and (layer6_outputs(2530));
    outputs(360) <= (layer6_outputs(439)) xor (layer6_outputs(1545));
    outputs(361) <= layer6_outputs(1465);
    outputs(362) <= layer6_outputs(880);
    outputs(363) <= (layer6_outputs(838)) and not (layer6_outputs(782));
    outputs(364) <= not(layer6_outputs(1074));
    outputs(365) <= (layer6_outputs(470)) xor (layer6_outputs(1672));
    outputs(366) <= (layer6_outputs(163)) and not (layer6_outputs(1867));
    outputs(367) <= not(layer6_outputs(799));
    outputs(368) <= not(layer6_outputs(1009));
    outputs(369) <= layer6_outputs(2515);
    outputs(370) <= (layer6_outputs(429)) and not (layer6_outputs(2547));
    outputs(371) <= not((layer6_outputs(441)) xor (layer6_outputs(67)));
    outputs(372) <= (layer6_outputs(1688)) xor (layer6_outputs(2057));
    outputs(373) <= not((layer6_outputs(1944)) or (layer6_outputs(1090)));
    outputs(374) <= not(layer6_outputs(85));
    outputs(375) <= layer6_outputs(1199);
    outputs(376) <= not(layer6_outputs(574));
    outputs(377) <= layer6_outputs(582);
    outputs(378) <= (layer6_outputs(2107)) and not (layer6_outputs(929));
    outputs(379) <= (layer6_outputs(1651)) xor (layer6_outputs(1572));
    outputs(380) <= layer6_outputs(2512);
    outputs(381) <= layer6_outputs(672);
    outputs(382) <= layer6_outputs(1972);
    outputs(383) <= (layer6_outputs(1536)) and not (layer6_outputs(892));
    outputs(384) <= (layer6_outputs(80)) and not (layer6_outputs(380));
    outputs(385) <= not(layer6_outputs(573));
    outputs(386) <= not(layer6_outputs(2308));
    outputs(387) <= not(layer6_outputs(1388));
    outputs(388) <= not(layer6_outputs(503));
    outputs(389) <= layer6_outputs(2390);
    outputs(390) <= (layer6_outputs(1205)) xor (layer6_outputs(1165));
    outputs(391) <= (layer6_outputs(954)) and not (layer6_outputs(221));
    outputs(392) <= not(layer6_outputs(1545)) or (layer6_outputs(1643));
    outputs(393) <= (layer6_outputs(723)) xor (layer6_outputs(1526));
    outputs(394) <= (layer6_outputs(444)) and not (layer6_outputs(1529));
    outputs(395) <= not((layer6_outputs(995)) xor (layer6_outputs(465)));
    outputs(396) <= (layer6_outputs(1451)) and not (layer6_outputs(1321));
    outputs(397) <= (layer6_outputs(1646)) and not (layer6_outputs(2394));
    outputs(398) <= (layer6_outputs(378)) and not (layer6_outputs(2212));
    outputs(399) <= layer6_outputs(2453);
    outputs(400) <= not(layer6_outputs(373));
    outputs(401) <= (layer6_outputs(1813)) and not (layer6_outputs(139));
    outputs(402) <= (layer6_outputs(1768)) and (layer6_outputs(1900));
    outputs(403) <= not(layer6_outputs(1389)) or (layer6_outputs(19));
    outputs(404) <= not(layer6_outputs(2477));
    outputs(405) <= not(layer6_outputs(671));
    outputs(406) <= not((layer6_outputs(1844)) xor (layer6_outputs(456)));
    outputs(407) <= layer6_outputs(1198);
    outputs(408) <= layer6_outputs(1523);
    outputs(409) <= layer6_outputs(66);
    outputs(410) <= not(layer6_outputs(1005));
    outputs(411) <= (layer6_outputs(620)) and not (layer6_outputs(76));
    outputs(412) <= (layer6_outputs(1345)) and (layer6_outputs(2074));
    outputs(413) <= layer6_outputs(2125);
    outputs(414) <= not(layer6_outputs(2140));
    outputs(415) <= layer6_outputs(107);
    outputs(416) <= not(layer6_outputs(1795));
    outputs(417) <= (layer6_outputs(1615)) and not (layer6_outputs(2559));
    outputs(418) <= not(layer6_outputs(1868));
    outputs(419) <= (layer6_outputs(1370)) and (layer6_outputs(2452));
    outputs(420) <= (layer6_outputs(255)) and (layer6_outputs(627));
    outputs(421) <= (layer6_outputs(1400)) and (layer6_outputs(1730));
    outputs(422) <= (layer6_outputs(237)) and not (layer6_outputs(1906));
    outputs(423) <= layer6_outputs(1224);
    outputs(424) <= layer6_outputs(1583);
    outputs(425) <= layer6_outputs(925);
    outputs(426) <= not((layer6_outputs(407)) or (layer6_outputs(2178)));
    outputs(427) <= (layer6_outputs(1708)) and not (layer6_outputs(1419));
    outputs(428) <= (layer6_outputs(858)) and not (layer6_outputs(1319));
    outputs(429) <= layer6_outputs(1846);
    outputs(430) <= layer6_outputs(1539);
    outputs(431) <= (layer6_outputs(693)) and (layer6_outputs(148));
    outputs(432) <= (layer6_outputs(1745)) and not (layer6_outputs(1977));
    outputs(433) <= (layer6_outputs(2090)) and (layer6_outputs(698));
    outputs(434) <= (layer6_outputs(1179)) xor (layer6_outputs(1282));
    outputs(435) <= (layer6_outputs(1142)) and (layer6_outputs(687));
    outputs(436) <= layer6_outputs(1822);
    outputs(437) <= not(layer6_outputs(571));
    outputs(438) <= not(layer6_outputs(679));
    outputs(439) <= not(layer6_outputs(877));
    outputs(440) <= (layer6_outputs(954)) and not (layer6_outputs(93));
    outputs(441) <= (layer6_outputs(968)) or (layer6_outputs(52));
    outputs(442) <= layer6_outputs(924);
    outputs(443) <= layer6_outputs(1897);
    outputs(444) <= not((layer6_outputs(481)) or (layer6_outputs(1419)));
    outputs(445) <= layer6_outputs(1989);
    outputs(446) <= (layer6_outputs(1171)) and (layer6_outputs(420));
    outputs(447) <= (layer6_outputs(360)) or (layer6_outputs(1272));
    outputs(448) <= not(layer6_outputs(86));
    outputs(449) <= layer6_outputs(745);
    outputs(450) <= layer6_outputs(2091);
    outputs(451) <= layer6_outputs(1214);
    outputs(452) <= not((layer6_outputs(1966)) xor (layer6_outputs(406)));
    outputs(453) <= (layer6_outputs(1328)) and not (layer6_outputs(1108));
    outputs(454) <= (layer6_outputs(2087)) and not (layer6_outputs(882));
    outputs(455) <= (layer6_outputs(1601)) and not (layer6_outputs(542));
    outputs(456) <= (layer6_outputs(1513)) and (layer6_outputs(1237));
    outputs(457) <= not((layer6_outputs(1484)) xor (layer6_outputs(394)));
    outputs(458) <= not(layer6_outputs(1458));
    outputs(459) <= not(layer6_outputs(2051));
    outputs(460) <= not((layer6_outputs(1112)) and (layer6_outputs(1873)));
    outputs(461) <= (layer6_outputs(1423)) and not (layer6_outputs(221));
    outputs(462) <= layer6_outputs(1114);
    outputs(463) <= layer6_outputs(2284);
    outputs(464) <= (layer6_outputs(1117)) and not (layer6_outputs(358));
    outputs(465) <= not(layer6_outputs(479));
    outputs(466) <= (layer6_outputs(1735)) and not (layer6_outputs(2458));
    outputs(467) <= not(layer6_outputs(2545));
    outputs(468) <= not(layer6_outputs(661));
    outputs(469) <= not(layer6_outputs(737)) or (layer6_outputs(52));
    outputs(470) <= (layer6_outputs(2383)) xor (layer6_outputs(10));
    outputs(471) <= not(layer6_outputs(1555));
    outputs(472) <= not((layer6_outputs(2100)) or (layer6_outputs(191)));
    outputs(473) <= (layer6_outputs(412)) and (layer6_outputs(412));
    outputs(474) <= (layer6_outputs(1100)) xor (layer6_outputs(523));
    outputs(475) <= not((layer6_outputs(1320)) or (layer6_outputs(1791)));
    outputs(476) <= (layer6_outputs(393)) and not (layer6_outputs(1359));
    outputs(477) <= (layer6_outputs(54)) and not (layer6_outputs(388));
    outputs(478) <= (layer6_outputs(1268)) and not (layer6_outputs(496));
    outputs(479) <= layer6_outputs(282);
    outputs(480) <= layer6_outputs(1386);
    outputs(481) <= not(layer6_outputs(1950));
    outputs(482) <= layer6_outputs(1244);
    outputs(483) <= (layer6_outputs(1093)) and not (layer6_outputs(539));
    outputs(484) <= layer6_outputs(2363);
    outputs(485) <= (layer6_outputs(666)) and (layer6_outputs(1234));
    outputs(486) <= not((layer6_outputs(2480)) xor (layer6_outputs(98)));
    outputs(487) <= not((layer6_outputs(573)) or (layer6_outputs(81)));
    outputs(488) <= not(layer6_outputs(1542));
    outputs(489) <= layer6_outputs(1001);
    outputs(490) <= not(layer6_outputs(2325));
    outputs(491) <= (layer6_outputs(236)) and not (layer6_outputs(2433));
    outputs(492) <= (layer6_outputs(905)) and not (layer6_outputs(966));
    outputs(493) <= (layer6_outputs(570)) or (layer6_outputs(854));
    outputs(494) <= not((layer6_outputs(1579)) or (layer6_outputs(2357)));
    outputs(495) <= not(layer6_outputs(1018));
    outputs(496) <= not(layer6_outputs(814)) or (layer6_outputs(998));
    outputs(497) <= (layer6_outputs(2530)) and (layer6_outputs(2202));
    outputs(498) <= layer6_outputs(101);
    outputs(499) <= (layer6_outputs(1434)) xor (layer6_outputs(1935));
    outputs(500) <= not(layer6_outputs(631));
    outputs(501) <= (layer6_outputs(770)) or (layer6_outputs(807));
    outputs(502) <= not(layer6_outputs(430));
    outputs(503) <= not(layer6_outputs(2213));
    outputs(504) <= layer6_outputs(2046);
    outputs(505) <= not(layer6_outputs(893));
    outputs(506) <= (layer6_outputs(1334)) and not (layer6_outputs(1905));
    outputs(507) <= layer6_outputs(275);
    outputs(508) <= not(layer6_outputs(2055));
    outputs(509) <= layer6_outputs(497);
    outputs(510) <= not((layer6_outputs(1532)) or (layer6_outputs(232)));
    outputs(511) <= (layer6_outputs(1106)) and not (layer6_outputs(511));
    outputs(512) <= not(layer6_outputs(320));
    outputs(513) <= layer6_outputs(1826);
    outputs(514) <= (layer6_outputs(2020)) and not (layer6_outputs(942));
    outputs(515) <= (layer6_outputs(2325)) and (layer6_outputs(174));
    outputs(516) <= not((layer6_outputs(1994)) xor (layer6_outputs(1033)));
    outputs(517) <= not((layer6_outputs(1880)) xor (layer6_outputs(2115)));
    outputs(518) <= layer6_outputs(204);
    outputs(519) <= (layer6_outputs(941)) and not (layer6_outputs(1471));
    outputs(520) <= layer6_outputs(1541);
    outputs(521) <= layer6_outputs(961);
    outputs(522) <= layer6_outputs(138);
    outputs(523) <= layer6_outputs(2350);
    outputs(524) <= (layer6_outputs(2543)) and not (layer6_outputs(2078));
    outputs(525) <= not(layer6_outputs(753)) or (layer6_outputs(1519));
    outputs(526) <= (layer6_outputs(1881)) and not (layer6_outputs(102));
    outputs(527) <= not((layer6_outputs(1778)) xor (layer6_outputs(911)));
    outputs(528) <= layer6_outputs(386);
    outputs(529) <= not(layer6_outputs(166));
    outputs(530) <= not(layer6_outputs(697));
    outputs(531) <= not(layer6_outputs(2197)) or (layer6_outputs(1874));
    outputs(532) <= not((layer6_outputs(309)) and (layer6_outputs(1140)));
    outputs(533) <= not(layer6_outputs(2545));
    outputs(534) <= not(layer6_outputs(2069));
    outputs(535) <= not(layer6_outputs(452)) or (layer6_outputs(1674));
    outputs(536) <= layer6_outputs(1785);
    outputs(537) <= layer6_outputs(159);
    outputs(538) <= layer6_outputs(2145);
    outputs(539) <= (layer6_outputs(1198)) xor (layer6_outputs(1880));
    outputs(540) <= (layer6_outputs(1487)) xor (layer6_outputs(497));
    outputs(541) <= (layer6_outputs(1604)) and not (layer6_outputs(1650));
    outputs(542) <= layer6_outputs(1079);
    outputs(543) <= layer6_outputs(605);
    outputs(544) <= (layer6_outputs(1557)) and not (layer6_outputs(2269));
    outputs(545) <= layer6_outputs(1470);
    outputs(546) <= (layer6_outputs(711)) and not (layer6_outputs(2359));
    outputs(547) <= not(layer6_outputs(129));
    outputs(548) <= not((layer6_outputs(1213)) or (layer6_outputs(88)));
    outputs(549) <= layer6_outputs(1643);
    outputs(550) <= not(layer6_outputs(1309)) or (layer6_outputs(1342));
    outputs(551) <= (layer6_outputs(907)) xor (layer6_outputs(1777));
    outputs(552) <= not((layer6_outputs(218)) xor (layer6_outputs(859)));
    outputs(553) <= not(layer6_outputs(2264));
    outputs(554) <= not(layer6_outputs(901));
    outputs(555) <= not(layer6_outputs(1129));
    outputs(556) <= not(layer6_outputs(2553));
    outputs(557) <= not((layer6_outputs(273)) xor (layer6_outputs(1305)));
    outputs(558) <= not((layer6_outputs(229)) xor (layer6_outputs(30)));
    outputs(559) <= (layer6_outputs(384)) and not (layer6_outputs(787));
    outputs(560) <= layer6_outputs(610);
    outputs(561) <= not(layer6_outputs(638));
    outputs(562) <= not(layer6_outputs(115));
    outputs(563) <= (layer6_outputs(116)) xor (layer6_outputs(1644));
    outputs(564) <= not(layer6_outputs(1835));
    outputs(565) <= (layer6_outputs(1283)) or (layer6_outputs(1882));
    outputs(566) <= (layer6_outputs(1195)) xor (layer6_outputs(1239));
    outputs(567) <= not(layer6_outputs(1610));
    outputs(568) <= (layer6_outputs(1896)) and not (layer6_outputs(266));
    outputs(569) <= (layer6_outputs(2550)) xor (layer6_outputs(1410));
    outputs(570) <= not(layer6_outputs(2387)) or (layer6_outputs(1562));
    outputs(571) <= not(layer6_outputs(1472));
    outputs(572) <= layer6_outputs(1542);
    outputs(573) <= not(layer6_outputs(1964)) or (layer6_outputs(2236));
    outputs(574) <= not((layer6_outputs(1003)) xor (layer6_outputs(2550)));
    outputs(575) <= not(layer6_outputs(2272));
    outputs(576) <= not(layer6_outputs(1155));
    outputs(577) <= not(layer6_outputs(588)) or (layer6_outputs(1653));
    outputs(578) <= not(layer6_outputs(2184));
    outputs(579) <= not(layer6_outputs(1584));
    outputs(580) <= layer6_outputs(1957);
    outputs(581) <= (layer6_outputs(1372)) xor (layer6_outputs(1756));
    outputs(582) <= not(layer6_outputs(2274));
    outputs(583) <= layer6_outputs(632);
    outputs(584) <= not((layer6_outputs(175)) xor (layer6_outputs(1432)));
    outputs(585) <= layer6_outputs(1054);
    outputs(586) <= not(layer6_outputs(791));
    outputs(587) <= not(layer6_outputs(1363));
    outputs(588) <= (layer6_outputs(1702)) xor (layer6_outputs(1145));
    outputs(589) <= (layer6_outputs(401)) xor (layer6_outputs(1938));
    outputs(590) <= not((layer6_outputs(1248)) xor (layer6_outputs(201)));
    outputs(591) <= layer6_outputs(2210);
    outputs(592) <= not(layer6_outputs(48));
    outputs(593) <= (layer6_outputs(1353)) xor (layer6_outputs(465));
    outputs(594) <= not((layer6_outputs(2022)) xor (layer6_outputs(1641)));
    outputs(595) <= layer6_outputs(1395);
    outputs(596) <= layer6_outputs(186);
    outputs(597) <= layer6_outputs(100);
    outputs(598) <= (layer6_outputs(2193)) and not (layer6_outputs(1242));
    outputs(599) <= not(layer6_outputs(915));
    outputs(600) <= (layer6_outputs(1667)) and not (layer6_outputs(635));
    outputs(601) <= not((layer6_outputs(2228)) and (layer6_outputs(2208)));
    outputs(602) <= not(layer6_outputs(2389));
    outputs(603) <= layer6_outputs(919);
    outputs(604) <= not(layer6_outputs(1004));
    outputs(605) <= not(layer6_outputs(419));
    outputs(606) <= layer6_outputs(1131);
    outputs(607) <= (layer6_outputs(785)) xor (layer6_outputs(1819));
    outputs(608) <= (layer6_outputs(1438)) and not (layer6_outputs(2508));
    outputs(609) <= not(layer6_outputs(1621));
    outputs(610) <= (layer6_outputs(2079)) or (layer6_outputs(1016));
    outputs(611) <= not(layer6_outputs(519));
    outputs(612) <= not((layer6_outputs(2455)) xor (layer6_outputs(2400)));
    outputs(613) <= layer6_outputs(314);
    outputs(614) <= not(layer6_outputs(1293));
    outputs(615) <= not(layer6_outputs(806));
    outputs(616) <= not(layer6_outputs(2297)) or (layer6_outputs(1842));
    outputs(617) <= not(layer6_outputs(1382));
    outputs(618) <= (layer6_outputs(1318)) and not (layer6_outputs(2381));
    outputs(619) <= not((layer6_outputs(1127)) xor (layer6_outputs(474)));
    outputs(620) <= (layer6_outputs(2474)) and not (layer6_outputs(789));
    outputs(621) <= not(layer6_outputs(1739));
    outputs(622) <= (layer6_outputs(1270)) and not (layer6_outputs(388));
    outputs(623) <= layer6_outputs(989);
    outputs(624) <= not((layer6_outputs(1757)) xor (layer6_outputs(648)));
    outputs(625) <= not(layer6_outputs(1885));
    outputs(626) <= (layer6_outputs(1673)) xor (layer6_outputs(2385));
    outputs(627) <= not((layer6_outputs(1559)) xor (layer6_outputs(1098)));
    outputs(628) <= layer6_outputs(21);
    outputs(629) <= not(layer6_outputs(984));
    outputs(630) <= not((layer6_outputs(2540)) xor (layer6_outputs(581)));
    outputs(631) <= layer6_outputs(2321);
    outputs(632) <= not((layer6_outputs(423)) xor (layer6_outputs(545)));
    outputs(633) <= layer6_outputs(1403);
    outputs(634) <= not((layer6_outputs(2368)) or (layer6_outputs(641)));
    outputs(635) <= not((layer6_outputs(903)) xor (layer6_outputs(1934)));
    outputs(636) <= (layer6_outputs(1933)) and not (layer6_outputs(426));
    outputs(637) <= not(layer6_outputs(2556)) or (layer6_outputs(232));
    outputs(638) <= not((layer6_outputs(1664)) or (layer6_outputs(554)));
    outputs(639) <= not(layer6_outputs(2045));
    outputs(640) <= (layer6_outputs(1719)) xor (layer6_outputs(1905));
    outputs(641) <= layer6_outputs(2250);
    outputs(642) <= not((layer6_outputs(1027)) or (layer6_outputs(1211)));
    outputs(643) <= layer6_outputs(2189);
    outputs(644) <= not((layer6_outputs(1424)) xor (layer6_outputs(1297)));
    outputs(645) <= not(layer6_outputs(407));
    outputs(646) <= (layer6_outputs(1564)) and (layer6_outputs(2066));
    outputs(647) <= layer6_outputs(1860);
    outputs(648) <= layer6_outputs(575);
    outputs(649) <= not((layer6_outputs(2420)) and (layer6_outputs(1929)));
    outputs(650) <= not(layer6_outputs(1706)) or (layer6_outputs(729));
    outputs(651) <= (layer6_outputs(1479)) and not (layer6_outputs(285));
    outputs(652) <= not((layer6_outputs(225)) or (layer6_outputs(234)));
    outputs(653) <= layer6_outputs(213);
    outputs(654) <= not((layer6_outputs(1057)) xor (layer6_outputs(1407)));
    outputs(655) <= layer6_outputs(1617);
    outputs(656) <= layer6_outputs(2284);
    outputs(657) <= layer6_outputs(813);
    outputs(658) <= (layer6_outputs(359)) xor (layer6_outputs(1050));
    outputs(659) <= layer6_outputs(772);
    outputs(660) <= (layer6_outputs(689)) and not (layer6_outputs(324));
    outputs(661) <= not(layer6_outputs(943));
    outputs(662) <= not(layer6_outputs(2087)) or (layer6_outputs(2082));
    outputs(663) <= (layer6_outputs(916)) and not (layer6_outputs(47));
    outputs(664) <= (layer6_outputs(1844)) xor (layer6_outputs(519));
    outputs(665) <= (layer6_outputs(1031)) and not (layer6_outputs(189));
    outputs(666) <= not((layer6_outputs(208)) xor (layer6_outputs(1489)));
    outputs(667) <= layer6_outputs(1899);
    outputs(668) <= not((layer6_outputs(65)) xor (layer6_outputs(1478)));
    outputs(669) <= layer6_outputs(900);
    outputs(670) <= not((layer6_outputs(194)) xor (layer6_outputs(2464)));
    outputs(671) <= not((layer6_outputs(2243)) xor (layer6_outputs(215)));
    outputs(672) <= layer6_outputs(458);
    outputs(673) <= layer6_outputs(2498);
    outputs(674) <= not(layer6_outputs(1754));
    outputs(675) <= (layer6_outputs(1069)) and not (layer6_outputs(712));
    outputs(676) <= (layer6_outputs(703)) and not (layer6_outputs(467));
    outputs(677) <= layer6_outputs(328);
    outputs(678) <= not((layer6_outputs(890)) xor (layer6_outputs(650)));
    outputs(679) <= layer6_outputs(21);
    outputs(680) <= (layer6_outputs(2164)) and (layer6_outputs(748));
    outputs(681) <= not((layer6_outputs(2092)) xor (layer6_outputs(1980)));
    outputs(682) <= (layer6_outputs(2136)) xor (layer6_outputs(492));
    outputs(683) <= (layer6_outputs(166)) xor (layer6_outputs(2197));
    outputs(684) <= (layer6_outputs(1338)) and (layer6_outputs(2376));
    outputs(685) <= not(layer6_outputs(1739));
    outputs(686) <= layer6_outputs(1147);
    outputs(687) <= not((layer6_outputs(1221)) xor (layer6_outputs(1634)));
    outputs(688) <= layer6_outputs(476);
    outputs(689) <= not(layer6_outputs(886));
    outputs(690) <= layer6_outputs(893);
    outputs(691) <= layer6_outputs(659);
    outputs(692) <= (layer6_outputs(1938)) and not (layer6_outputs(1699));
    outputs(693) <= (layer6_outputs(2186)) and (layer6_outputs(1318));
    outputs(694) <= layer6_outputs(1306);
    outputs(695) <= (layer6_outputs(1019)) xor (layer6_outputs(185));
    outputs(696) <= not(layer6_outputs(1912));
    outputs(697) <= layer6_outputs(730);
    outputs(698) <= not(layer6_outputs(1522));
    outputs(699) <= not(layer6_outputs(942));
    outputs(700) <= layer6_outputs(1748);
    outputs(701) <= not(layer6_outputs(2527));
    outputs(702) <= layer6_outputs(2370);
    outputs(703) <= layer6_outputs(2040);
    outputs(704) <= not(layer6_outputs(2495));
    outputs(705) <= layer6_outputs(2520);
    outputs(706) <= not(layer6_outputs(193)) or (layer6_outputs(941));
    outputs(707) <= (layer6_outputs(2332)) xor (layer6_outputs(25));
    outputs(708) <= layer6_outputs(124);
    outputs(709) <= layer6_outputs(1395);
    outputs(710) <= not((layer6_outputs(1689)) xor (layer6_outputs(1756)));
    outputs(711) <= (layer6_outputs(1884)) and (layer6_outputs(2073));
    outputs(712) <= not(layer6_outputs(155));
    outputs(713) <= not(layer6_outputs(2246));
    outputs(714) <= layer6_outputs(72);
    outputs(715) <= (layer6_outputs(2106)) and not (layer6_outputs(1670));
    outputs(716) <= not((layer6_outputs(1046)) xor (layer6_outputs(1134)));
    outputs(717) <= (layer6_outputs(2154)) or (layer6_outputs(1653));
    outputs(718) <= (layer6_outputs(1746)) and (layer6_outputs(2243));
    outputs(719) <= layer6_outputs(976);
    outputs(720) <= not(layer6_outputs(180));
    outputs(721) <= not((layer6_outputs(1947)) xor (layer6_outputs(1381)));
    outputs(722) <= layer6_outputs(500);
    outputs(723) <= not(layer6_outputs(2507));
    outputs(724) <= layer6_outputs(1811);
    outputs(725) <= (layer6_outputs(342)) xor (layer6_outputs(1926));
    outputs(726) <= not(layer6_outputs(1514));
    outputs(727) <= layer6_outputs(1099);
    outputs(728) <= not(layer6_outputs(426));
    outputs(729) <= not((layer6_outputs(971)) or (layer6_outputs(140)));
    outputs(730) <= not((layer6_outputs(990)) xor (layer6_outputs(2065)));
    outputs(731) <= (layer6_outputs(2542)) and (layer6_outputs(2432));
    outputs(732) <= not((layer6_outputs(1444)) xor (layer6_outputs(1541)));
    outputs(733) <= layer6_outputs(446);
    outputs(734) <= layer6_outputs(2071);
    outputs(735) <= layer6_outputs(1726);
    outputs(736) <= layer6_outputs(1010);
    outputs(737) <= not((layer6_outputs(2060)) and (layer6_outputs(2374)));
    outputs(738) <= (layer6_outputs(1680)) or (layer6_outputs(916));
    outputs(739) <= layer6_outputs(784);
    outputs(740) <= not(layer6_outputs(2295)) or (layer6_outputs(1308));
    outputs(741) <= layer6_outputs(600);
    outputs(742) <= not(layer6_outputs(765));
    outputs(743) <= layer6_outputs(1227);
    outputs(744) <= not(layer6_outputs(599));
    outputs(745) <= layer6_outputs(619);
    outputs(746) <= not(layer6_outputs(469));
    outputs(747) <= (layer6_outputs(257)) and not (layer6_outputs(1378));
    outputs(748) <= (layer6_outputs(1866)) xor (layer6_outputs(1912));
    outputs(749) <= layer6_outputs(869);
    outputs(750) <= (layer6_outputs(94)) xor (layer6_outputs(345));
    outputs(751) <= not((layer6_outputs(655)) xor (layer6_outputs(1832)));
    outputs(752) <= (layer6_outputs(2123)) xor (layer6_outputs(738));
    outputs(753) <= layer6_outputs(822);
    outputs(754) <= layer6_outputs(54);
    outputs(755) <= layer6_outputs(1360);
    outputs(756) <= layer6_outputs(1773);
    outputs(757) <= not(layer6_outputs(2423));
    outputs(758) <= not(layer6_outputs(1834));
    outputs(759) <= not(layer6_outputs(668));
    outputs(760) <= not(layer6_outputs(1570));
    outputs(761) <= not(layer6_outputs(584));
    outputs(762) <= (layer6_outputs(1859)) xor (layer6_outputs(507));
    outputs(763) <= not((layer6_outputs(109)) xor (layer6_outputs(1072)));
    outputs(764) <= (layer6_outputs(1808)) and (layer6_outputs(922));
    outputs(765) <= layer6_outputs(173);
    outputs(766) <= not((layer6_outputs(2407)) xor (layer6_outputs(1231)));
    outputs(767) <= not((layer6_outputs(32)) xor (layer6_outputs(393)));
    outputs(768) <= not(layer6_outputs(1464));
    outputs(769) <= layer6_outputs(438);
    outputs(770) <= (layer6_outputs(1982)) xor (layer6_outputs(103));
    outputs(771) <= layer6_outputs(1173);
    outputs(772) <= not(layer6_outputs(1193)) or (layer6_outputs(852));
    outputs(773) <= not(layer6_outputs(1665));
    outputs(774) <= not(layer6_outputs(473));
    outputs(775) <= (layer6_outputs(1358)) and (layer6_outputs(1609));
    outputs(776) <= layer6_outputs(2364);
    outputs(777) <= not(layer6_outputs(710));
    outputs(778) <= not((layer6_outputs(2320)) xor (layer6_outputs(2440)));
    outputs(779) <= layer6_outputs(1128);
    outputs(780) <= layer6_outputs(2064);
    outputs(781) <= (layer6_outputs(815)) and not (layer6_outputs(697));
    outputs(782) <= layer6_outputs(823);
    outputs(783) <= not((layer6_outputs(1873)) xor (layer6_outputs(1690)));
    outputs(784) <= layer6_outputs(1096);
    outputs(785) <= not(layer6_outputs(807));
    outputs(786) <= not((layer6_outputs(296)) and (layer6_outputs(14)));
    outputs(787) <= (layer6_outputs(567)) and (layer6_outputs(2048));
    outputs(788) <= not((layer6_outputs(856)) and (layer6_outputs(648)));
    outputs(789) <= layer6_outputs(1260);
    outputs(790) <= layer6_outputs(319);
    outputs(791) <= (layer6_outputs(1593)) and not (layer6_outputs(1120));
    outputs(792) <= not(layer6_outputs(2237));
    outputs(793) <= (layer6_outputs(2191)) or (layer6_outputs(463));
    outputs(794) <= (layer6_outputs(705)) and not (layer6_outputs(395));
    outputs(795) <= (layer6_outputs(2095)) and not (layer6_outputs(1219));
    outputs(796) <= not(layer6_outputs(2424));
    outputs(797) <= (layer6_outputs(872)) and (layer6_outputs(300));
    outputs(798) <= not(layer6_outputs(396)) or (layer6_outputs(42));
    outputs(799) <= not((layer6_outputs(1350)) or (layer6_outputs(234)));
    outputs(800) <= not((layer6_outputs(635)) xor (layer6_outputs(1713)));
    outputs(801) <= (layer6_outputs(387)) and (layer6_outputs(1435));
    outputs(802) <= not(layer6_outputs(1474));
    outputs(803) <= (layer6_outputs(2391)) and not (layer6_outputs(448));
    outputs(804) <= not(layer6_outputs(2220)) or (layer6_outputs(1805));
    outputs(805) <= (layer6_outputs(1433)) xor (layer6_outputs(1303));
    outputs(806) <= layer6_outputs(1886);
    outputs(807) <= not((layer6_outputs(617)) or (layer6_outputs(2387)));
    outputs(808) <= layer6_outputs(543);
    outputs(809) <= not((layer6_outputs(1556)) or (layer6_outputs(844)));
    outputs(810) <= not((layer6_outputs(885)) xor (layer6_outputs(996)));
    outputs(811) <= not(layer6_outputs(821));
    outputs(812) <= layer6_outputs(1246);
    outputs(813) <= not(layer6_outputs(563));
    outputs(814) <= layer6_outputs(244);
    outputs(815) <= layer6_outputs(1266);
    outputs(816) <= not(layer6_outputs(2234));
    outputs(817) <= not(layer6_outputs(1167));
    outputs(818) <= (layer6_outputs(816)) and not (layer6_outputs(2393));
    outputs(819) <= not(layer6_outputs(2116));
    outputs(820) <= (layer6_outputs(1170)) and not (layer6_outputs(782));
    outputs(821) <= (layer6_outputs(433)) xor (layer6_outputs(1087));
    outputs(822) <= not(layer6_outputs(2001));
    outputs(823) <= not(layer6_outputs(2200));
    outputs(824) <= (layer6_outputs(2203)) xor (layer6_outputs(2406));
    outputs(825) <= not(layer6_outputs(2229));
    outputs(826) <= layer6_outputs(115);
    outputs(827) <= layer6_outputs(2382);
    outputs(828) <= not((layer6_outputs(2222)) xor (layer6_outputs(2531)));
    outputs(829) <= not((layer6_outputs(1202)) xor (layer6_outputs(2119)));
    outputs(830) <= (layer6_outputs(768)) xor (layer6_outputs(1188));
    outputs(831) <= (layer6_outputs(614)) and not (layer6_outputs(1186));
    outputs(832) <= not((layer6_outputs(1486)) xor (layer6_outputs(2547)));
    outputs(833) <= layer6_outputs(1884);
    outputs(834) <= (layer6_outputs(2319)) and (layer6_outputs(1578));
    outputs(835) <= (layer6_outputs(1197)) and not (layer6_outputs(827));
    outputs(836) <= not((layer6_outputs(333)) or (layer6_outputs(8)));
    outputs(837) <= not((layer6_outputs(683)) or (layer6_outputs(1791)));
    outputs(838) <= not(layer6_outputs(521));
    outputs(839) <= (layer6_outputs(654)) and not (layer6_outputs(1418));
    outputs(840) <= not(layer6_outputs(624));
    outputs(841) <= not(layer6_outputs(1175));
    outputs(842) <= layer6_outputs(53);
    outputs(843) <= layer6_outputs(436);
    outputs(844) <= not(layer6_outputs(2012));
    outputs(845) <= layer6_outputs(1063);
    outputs(846) <= (layer6_outputs(2368)) and not (layer6_outputs(332));
    outputs(847) <= (layer6_outputs(447)) and not (layer6_outputs(688));
    outputs(848) <= not((layer6_outputs(544)) xor (layer6_outputs(1194)));
    outputs(849) <= not(layer6_outputs(120));
    outputs(850) <= (layer6_outputs(758)) and not (layer6_outputs(1941));
    outputs(851) <= (layer6_outputs(1453)) xor (layer6_outputs(1460));
    outputs(852) <= not((layer6_outputs(2448)) or (layer6_outputs(2438)));
    outputs(853) <= (layer6_outputs(1771)) and not (layer6_outputs(2306));
    outputs(854) <= layer6_outputs(898);
    outputs(855) <= (layer6_outputs(1690)) xor (layer6_outputs(1174));
    outputs(856) <= layer6_outputs(1029);
    outputs(857) <= (layer6_outputs(676)) and not (layer6_outputs(1155));
    outputs(858) <= not(layer6_outputs(1037));
    outputs(859) <= not(layer6_outputs(1113));
    outputs(860) <= not(layer6_outputs(1061));
    outputs(861) <= layer6_outputs(1302);
    outputs(862) <= (layer6_outputs(2053)) xor (layer6_outputs(2384));
    outputs(863) <= not((layer6_outputs(1858)) and (layer6_outputs(1621)));
    outputs(864) <= (layer6_outputs(923)) and not (layer6_outputs(489));
    outputs(865) <= layer6_outputs(796);
    outputs(866) <= not(layer6_outputs(1677));
    outputs(867) <= layer6_outputs(802);
    outputs(868) <= (layer6_outputs(1563)) xor (layer6_outputs(226));
    outputs(869) <= (layer6_outputs(2376)) xor (layer6_outputs(609));
    outputs(870) <= not(layer6_outputs(1404));
    outputs(871) <= (layer6_outputs(321)) and not (layer6_outputs(209));
    outputs(872) <= (layer6_outputs(2270)) xor (layer6_outputs(1376));
    outputs(873) <= layer6_outputs(1868);
    outputs(874) <= layer6_outputs(1567);
    outputs(875) <= not((layer6_outputs(963)) xor (layer6_outputs(1602)));
    outputs(876) <= not((layer6_outputs(57)) or (layer6_outputs(2305)));
    outputs(877) <= (layer6_outputs(2288)) and not (layer6_outputs(403));
    outputs(878) <= not(layer6_outputs(1624));
    outputs(879) <= layer6_outputs(1520);
    outputs(880) <= not((layer6_outputs(773)) or (layer6_outputs(1656)));
    outputs(881) <= not(layer6_outputs(1481));
    outputs(882) <= not(layer6_outputs(2349));
    outputs(883) <= not(layer6_outputs(1073));
    outputs(884) <= layer6_outputs(1013);
    outputs(885) <= layer6_outputs(1191);
    outputs(886) <= layer6_outputs(1183);
    outputs(887) <= (layer6_outputs(636)) xor (layer6_outputs(305));
    outputs(888) <= not(layer6_outputs(2333));
    outputs(889) <= layer6_outputs(909);
    outputs(890) <= (layer6_outputs(449)) or (layer6_outputs(1759));
    outputs(891) <= (layer6_outputs(2548)) xor (layer6_outputs(2043));
    outputs(892) <= not(layer6_outputs(1080));
    outputs(893) <= layer6_outputs(860);
    outputs(894) <= not((layer6_outputs(2153)) xor (layer6_outputs(1401)));
    outputs(895) <= (layer6_outputs(160)) and (layer6_outputs(2373));
    outputs(896) <= not((layer6_outputs(2008)) xor (layer6_outputs(70)));
    outputs(897) <= layer6_outputs(2300);
    outputs(898) <= not(layer6_outputs(1413));
    outputs(899) <= not(layer6_outputs(2003));
    outputs(900) <= not((layer6_outputs(1779)) xor (layer6_outputs(898)));
    outputs(901) <= not(layer6_outputs(2519)) or (layer6_outputs(1915));
    outputs(902) <= not(layer6_outputs(683));
    outputs(903) <= not(layer6_outputs(1420));
    outputs(904) <= not(layer6_outputs(979));
    outputs(905) <= layer6_outputs(2443);
    outputs(906) <= layer6_outputs(1599);
    outputs(907) <= not(layer6_outputs(597));
    outputs(908) <= layer6_outputs(1214);
    outputs(909) <= not((layer6_outputs(2229)) and (layer6_outputs(1281)));
    outputs(910) <= (layer6_outputs(1828)) or (layer6_outputs(1798));
    outputs(911) <= layer6_outputs(2371);
    outputs(912) <= layer6_outputs(293);
    outputs(913) <= (layer6_outputs(630)) and (layer6_outputs(1781));
    outputs(914) <= not((layer6_outputs(1298)) xor (layer6_outputs(3)));
    outputs(915) <= not(layer6_outputs(1622)) or (layer6_outputs(1594));
    outputs(916) <= not((layer6_outputs(1750)) or (layer6_outputs(509)));
    outputs(917) <= not(layer6_outputs(1220));
    outputs(918) <= not(layer6_outputs(2353));
    outputs(919) <= not(layer6_outputs(2023));
    outputs(920) <= (layer6_outputs(796)) and not (layer6_outputs(1194));
    outputs(921) <= not(layer6_outputs(2536));
    outputs(922) <= (layer6_outputs(1601)) and not (layer6_outputs(2185));
    outputs(923) <= (layer6_outputs(1641)) and (layer6_outputs(833));
    outputs(924) <= (layer6_outputs(1229)) and not (layer6_outputs(1540));
    outputs(925) <= (layer6_outputs(2218)) and (layer6_outputs(1787));
    outputs(926) <= not(layer6_outputs(569));
    outputs(927) <= layer6_outputs(1320);
    outputs(928) <= not(layer6_outputs(2396));
    outputs(929) <= not((layer6_outputs(2143)) or (layer6_outputs(1944)));
    outputs(930) <= not(layer6_outputs(1213));
    outputs(931) <= layer6_outputs(1801);
    outputs(932) <= (layer6_outputs(1854)) and (layer6_outputs(2117));
    outputs(933) <= not((layer6_outputs(1369)) xor (layer6_outputs(1498)));
    outputs(934) <= layer6_outputs(872);
    outputs(935) <= not(layer6_outputs(987));
    outputs(936) <= layer6_outputs(513);
    outputs(937) <= not((layer6_outputs(1351)) xor (layer6_outputs(194)));
    outputs(938) <= layer6_outputs(1114);
    outputs(939) <= (layer6_outputs(203)) and not (layer6_outputs(91));
    outputs(940) <= (layer6_outputs(386)) and (layer6_outputs(2030));
    outputs(941) <= layer6_outputs(60);
    outputs(942) <= (layer6_outputs(334)) and (layer6_outputs(2162));
    outputs(943) <= layer6_outputs(2377);
    outputs(944) <= not((layer6_outputs(1094)) xor (layer6_outputs(321)));
    outputs(945) <= not(layer6_outputs(2052));
    outputs(946) <= layer6_outputs(456);
    outputs(947) <= not(layer6_outputs(384));
    outputs(948) <= not(layer6_outputs(96));
    outputs(949) <= not((layer6_outputs(1816)) xor (layer6_outputs(1790)));
    outputs(950) <= (layer6_outputs(835)) and not (layer6_outputs(749));
    outputs(951) <= not((layer6_outputs(99)) or (layer6_outputs(277)));
    outputs(952) <= (layer6_outputs(364)) and (layer6_outputs(2398));
    outputs(953) <= not(layer6_outputs(1767)) or (layer6_outputs(2013));
    outputs(954) <= not((layer6_outputs(1347)) and (layer6_outputs(311)));
    outputs(955) <= (layer6_outputs(1302)) and not (layer6_outputs(1659));
    outputs(956) <= not(layer6_outputs(2314));
    outputs(957) <= not(layer6_outputs(1058));
    outputs(958) <= not(layer6_outputs(78));
    outputs(959) <= layer6_outputs(2153);
    outputs(960) <= layer6_outputs(576);
    outputs(961) <= layer6_outputs(182);
    outputs(962) <= layer6_outputs(2347);
    outputs(963) <= layer6_outputs(2378);
    outputs(964) <= layer6_outputs(1516);
    outputs(965) <= layer6_outputs(604);
    outputs(966) <= (layer6_outputs(216)) and (layer6_outputs(1094));
    outputs(967) <= not((layer6_outputs(1551)) or (layer6_outputs(83)));
    outputs(968) <= not(layer6_outputs(2234));
    outputs(969) <= not(layer6_outputs(2051));
    outputs(970) <= not(layer6_outputs(1147));
    outputs(971) <= (layer6_outputs(2080)) and not (layer6_outputs(1464));
    outputs(972) <= not((layer6_outputs(2053)) xor (layer6_outputs(279)));
    outputs(973) <= not(layer6_outputs(2461));
    outputs(974) <= not(layer6_outputs(936));
    outputs(975) <= not(layer6_outputs(1462));
    outputs(976) <= not(layer6_outputs(1501));
    outputs(977) <= (layer6_outputs(2422)) and not (layer6_outputs(303));
    outputs(978) <= (layer6_outputs(958)) and not (layer6_outputs(434));
    outputs(979) <= layer6_outputs(834);
    outputs(980) <= not(layer6_outputs(1119));
    outputs(981) <= (layer6_outputs(1105)) and (layer6_outputs(353));
    outputs(982) <= not((layer6_outputs(126)) or (layer6_outputs(1088)));
    outputs(983) <= not(layer6_outputs(2307));
    outputs(984) <= (layer6_outputs(989)) and (layer6_outputs(1125));
    outputs(985) <= layer6_outputs(1095);
    outputs(986) <= not((layer6_outputs(2187)) or (layer6_outputs(390)));
    outputs(987) <= not((layer6_outputs(1047)) or (layer6_outputs(493)));
    outputs(988) <= not((layer6_outputs(603)) or (layer6_outputs(1725)));
    outputs(989) <= layer6_outputs(1168);
    outputs(990) <= not(layer6_outputs(249));
    outputs(991) <= (layer6_outputs(1714)) and (layer6_outputs(1576));
    outputs(992) <= not((layer6_outputs(133)) or (layer6_outputs(2120)));
    outputs(993) <= (layer6_outputs(861)) xor (layer6_outputs(2457));
    outputs(994) <= not((layer6_outputs(217)) and (layer6_outputs(1366)));
    outputs(995) <= (layer6_outputs(1185)) and not (layer6_outputs(130));
    outputs(996) <= not(layer6_outputs(2278));
    outputs(997) <= layer6_outputs(783);
    outputs(998) <= layer6_outputs(2492);
    outputs(999) <= not(layer6_outputs(1810));
    outputs(1000) <= not(layer6_outputs(1538));
    outputs(1001) <= (layer6_outputs(1634)) xor (layer6_outputs(1702));
    outputs(1002) <= layer6_outputs(1709);
    outputs(1003) <= not(layer6_outputs(1388));
    outputs(1004) <= layer6_outputs(2029);
    outputs(1005) <= (layer6_outputs(475)) and not (layer6_outputs(446));
    outputs(1006) <= not(layer6_outputs(2549));
    outputs(1007) <= not((layer6_outputs(203)) xor (layer6_outputs(2085)));
    outputs(1008) <= layer6_outputs(1397);
    outputs(1009) <= layer6_outputs(1112);
    outputs(1010) <= layer6_outputs(2398);
    outputs(1011) <= not(layer6_outputs(663));
    outputs(1012) <= (layer6_outputs(1103)) xor (layer6_outputs(540));
    outputs(1013) <= layer6_outputs(744);
    outputs(1014) <= not((layer6_outputs(346)) xor (layer6_outputs(128)));
    outputs(1015) <= not((layer6_outputs(379)) xor (layer6_outputs(1948)));
    outputs(1016) <= layer6_outputs(1557);
    outputs(1017) <= not(layer6_outputs(775));
    outputs(1018) <= (layer6_outputs(1865)) and not (layer6_outputs(77));
    outputs(1019) <= not(layer6_outputs(965));
    outputs(1020) <= not(layer6_outputs(997));
    outputs(1021) <= not((layer6_outputs(2397)) xor (layer6_outputs(934)));
    outputs(1022) <= not(layer6_outputs(926));
    outputs(1023) <= not(layer6_outputs(147));
    outputs(1024) <= layer6_outputs(2503);
    outputs(1025) <= (layer6_outputs(354)) xor (layer6_outputs(840));
    outputs(1026) <= layer6_outputs(1379);
    outputs(1027) <= not(layer6_outputs(1244));
    outputs(1028) <= layer6_outputs(953);
    outputs(1029) <= not(layer6_outputs(1633));
    outputs(1030) <= not((layer6_outputs(1695)) xor (layer6_outputs(1782)));
    outputs(1031) <= layer6_outputs(1776);
    outputs(1032) <= (layer6_outputs(472)) xor (layer6_outputs(629));
    outputs(1033) <= layer6_outputs(548);
    outputs(1034) <= layer6_outputs(2304);
    outputs(1035) <= not(layer6_outputs(2172));
    outputs(1036) <= (layer6_outputs(1280)) and not (layer6_outputs(387));
    outputs(1037) <= layer6_outputs(1385);
    outputs(1038) <= layer6_outputs(879);
    outputs(1039) <= not(layer6_outputs(151));
    outputs(1040) <= not(layer6_outputs(1502));
    outputs(1041) <= not(layer6_outputs(871)) or (layer6_outputs(1518));
    outputs(1042) <= not(layer6_outputs(1654));
    outputs(1043) <= (layer6_outputs(349)) xor (layer6_outputs(1343));
    outputs(1044) <= not(layer6_outputs(190));
    outputs(1045) <= not((layer6_outputs(1603)) xor (layer6_outputs(1501)));
    outputs(1046) <= not(layer6_outputs(1474));
    outputs(1047) <= layer6_outputs(1689);
    outputs(1048) <= layer6_outputs(1954);
    outputs(1049) <= not((layer6_outputs(2399)) xor (layer6_outputs(682)));
    outputs(1050) <= layer6_outputs(1483);
    outputs(1051) <= layer6_outputs(1104);
    outputs(1052) <= (layer6_outputs(1722)) and not (layer6_outputs(2491));
    outputs(1053) <= (layer6_outputs(1696)) xor (layer6_outputs(606));
    outputs(1054) <= not(layer6_outputs(257));
    outputs(1055) <= not(layer6_outputs(1683));
    outputs(1056) <= not(layer6_outputs(1312));
    outputs(1057) <= not(layer6_outputs(1170));
    outputs(1058) <= (layer6_outputs(2542)) and not (layer6_outputs(1028));
    outputs(1059) <= (layer6_outputs(1622)) xor (layer6_outputs(209));
    outputs(1060) <= (layer6_outputs(912)) and not (layer6_outputs(1196));
    outputs(1061) <= not(layer6_outputs(2022));
    outputs(1062) <= not((layer6_outputs(1383)) or (layer6_outputs(660)));
    outputs(1063) <= layer6_outputs(553);
    outputs(1064) <= layer6_outputs(60);
    outputs(1065) <= not(layer6_outputs(1148));
    outputs(1066) <= layer6_outputs(283);
    outputs(1067) <= not(layer6_outputs(899));
    outputs(1068) <= not(layer6_outputs(2165));
    outputs(1069) <= (layer6_outputs(2365)) and not (layer6_outputs(1290));
    outputs(1070) <= layer6_outputs(424);
    outputs(1071) <= layer6_outputs(780);
    outputs(1072) <= (layer6_outputs(895)) xor (layer6_outputs(1221));
    outputs(1073) <= not(layer6_outputs(2021));
    outputs(1074) <= (layer6_outputs(722)) and not (layer6_outputs(994));
    outputs(1075) <= (layer6_outputs(1287)) and not (layer6_outputs(2159));
    outputs(1076) <= layer6_outputs(2151);
    outputs(1077) <= not(layer6_outputs(2339));
    outputs(1078) <= not(layer6_outputs(627));
    outputs(1079) <= not(layer6_outputs(447)) or (layer6_outputs(123));
    outputs(1080) <= not(layer6_outputs(1473));
    outputs(1081) <= not((layer6_outputs(406)) xor (layer6_outputs(264)));
    outputs(1082) <= not(layer6_outputs(2369));
    outputs(1083) <= (layer6_outputs(793)) and (layer6_outputs(1233));
    outputs(1084) <= layer6_outputs(1627);
    outputs(1085) <= (layer6_outputs(1943)) xor (layer6_outputs(2201));
    outputs(1086) <= not(layer6_outputs(613));
    outputs(1087) <= not(layer6_outputs(2054));
    outputs(1088) <= (layer6_outputs(599)) and (layer6_outputs(2414));
    outputs(1089) <= not((layer6_outputs(1755)) xor (layer6_outputs(2216)));
    outputs(1090) <= (layer6_outputs(2248)) and (layer6_outputs(1738));
    outputs(1091) <= layer6_outputs(2076);
    outputs(1092) <= not(layer6_outputs(727));
    outputs(1093) <= layer6_outputs(1744);
    outputs(1094) <= not(layer6_outputs(367));
    outputs(1095) <= not((layer6_outputs(187)) and (layer6_outputs(2343)));
    outputs(1096) <= not((layer6_outputs(789)) xor (layer6_outputs(235)));
    outputs(1097) <= not(layer6_outputs(2204));
    outputs(1098) <= not(layer6_outputs(2094));
    outputs(1099) <= layer6_outputs(2414);
    outputs(1100) <= layer6_outputs(467);
    outputs(1101) <= not(layer6_outputs(1348));
    outputs(1102) <= (layer6_outputs(1387)) and not (layer6_outputs(100));
    outputs(1103) <= not(layer6_outputs(1492));
    outputs(1104) <= not((layer6_outputs(2244)) xor (layer6_outputs(2518)));
    outputs(1105) <= (layer6_outputs(1146)) and not (layer6_outputs(1939));
    outputs(1106) <= layer6_outputs(2487);
    outputs(1107) <= (layer6_outputs(1893)) xor (layer6_outputs(1866));
    outputs(1108) <= layer6_outputs(1729);
    outputs(1109) <= not(layer6_outputs(1937));
    outputs(1110) <= not(layer6_outputs(1609));
    outputs(1111) <= not((layer6_outputs(1011)) xor (layer6_outputs(2347)));
    outputs(1112) <= not((layer6_outputs(2324)) xor (layer6_outputs(2539)));
    outputs(1113) <= not(layer6_outputs(29));
    outputs(1114) <= (layer6_outputs(824)) xor (layer6_outputs(168));
    outputs(1115) <= layer6_outputs(2006);
    outputs(1116) <= layer6_outputs(1285);
    outputs(1117) <= (layer6_outputs(884)) and not (layer6_outputs(1342));
    outputs(1118) <= not((layer6_outputs(2077)) or (layer6_outputs(925)));
    outputs(1119) <= not((layer6_outputs(1982)) xor (layer6_outputs(289)));
    outputs(1120) <= layer6_outputs(2538);
    outputs(1121) <= (layer6_outputs(1344)) and not (layer6_outputs(200));
    outputs(1122) <= layer6_outputs(733);
    outputs(1123) <= not(layer6_outputs(1132)) or (layer6_outputs(631));
    outputs(1124) <= layer6_outputs(174);
    outputs(1125) <= not((layer6_outputs(2323)) xor (layer6_outputs(1778)));
    outputs(1126) <= not((layer6_outputs(414)) or (layer6_outputs(1869)));
    outputs(1127) <= layer6_outputs(47);
    outputs(1128) <= (layer6_outputs(1845)) and not (layer6_outputs(1367));
    outputs(1129) <= (layer6_outputs(749)) and (layer6_outputs(466));
    outputs(1130) <= (layer6_outputs(245)) and (layer6_outputs(1000));
    outputs(1131) <= (layer6_outputs(1203)) and not (layer6_outputs(1305));
    outputs(1132) <= layer6_outputs(1304);
    outputs(1133) <= (layer6_outputs(1507)) and not (layer6_outputs(510));
    outputs(1134) <= layer6_outputs(2456);
    outputs(1135) <= (layer6_outputs(2029)) xor (layer6_outputs(470));
    outputs(1136) <= layer6_outputs(1920);
    outputs(1137) <= not((layer6_outputs(805)) or (layer6_outputs(1330)));
    outputs(1138) <= not(layer6_outputs(845));
    outputs(1139) <= not(layer6_outputs(2058));
    outputs(1140) <= (layer6_outputs(2322)) and not (layer6_outputs(11));
    outputs(1141) <= layer6_outputs(152);
    outputs(1142) <= not(layer6_outputs(975));
    outputs(1143) <= not((layer6_outputs(1366)) xor (layer6_outputs(1304)));
    outputs(1144) <= not((layer6_outputs(1354)) xor (layer6_outputs(931)));
    outputs(1145) <= not(layer6_outputs(2135));
    outputs(1146) <= not(layer6_outputs(1319));
    outputs(1147) <= not((layer6_outputs(378)) xor (layer6_outputs(1038)));
    outputs(1148) <= (layer6_outputs(225)) and (layer6_outputs(1721));
    outputs(1149) <= not(layer6_outputs(59));
    outputs(1150) <= not(layer6_outputs(1840));
    outputs(1151) <= layer6_outputs(1916);
    outputs(1152) <= not(layer6_outputs(1976));
    outputs(1153) <= (layer6_outputs(15)) xor (layer6_outputs(1806));
    outputs(1154) <= layer6_outputs(1399);
    outputs(1155) <= (layer6_outputs(1769)) and not (layer6_outputs(2137));
    outputs(1156) <= layer6_outputs(2313);
    outputs(1157) <= (layer6_outputs(288)) and not (layer6_outputs(1639));
    outputs(1158) <= not(layer6_outputs(2276));
    outputs(1159) <= layer6_outputs(44);
    outputs(1160) <= layer6_outputs(1871);
    outputs(1161) <= layer6_outputs(901);
    outputs(1162) <= not(layer6_outputs(425));
    outputs(1163) <= (layer6_outputs(2245)) and not (layer6_outputs(1299));
    outputs(1164) <= not((layer6_outputs(1749)) or (layer6_outputs(2411)));
    outputs(1165) <= not((layer6_outputs(1034)) or (layer6_outputs(2116)));
    outputs(1166) <= layer6_outputs(1858);
    outputs(1167) <= layer6_outputs(2179);
    outputs(1168) <= not((layer6_outputs(1533)) and (layer6_outputs(1348)));
    outputs(1169) <= layer6_outputs(1500);
    outputs(1170) <= not(layer6_outputs(2526));
    outputs(1171) <= layer6_outputs(547);
    outputs(1172) <= not(layer6_outputs(1182)) or (layer6_outputs(981));
    outputs(1173) <= not(layer6_outputs(2400));
    outputs(1174) <= layer6_outputs(1809);
    outputs(1175) <= (layer6_outputs(2549)) xor (layer6_outputs(1050));
    outputs(1176) <= layer6_outputs(1051);
    outputs(1177) <= (layer6_outputs(692)) and not (layer6_outputs(914));
    outputs(1178) <= (layer6_outputs(2374)) and not (layer6_outputs(2534));
    outputs(1179) <= layer6_outputs(2206);
    outputs(1180) <= not((layer6_outputs(435)) xor (layer6_outputs(826)));
    outputs(1181) <= not(layer6_outputs(449));
    outputs(1182) <= not(layer6_outputs(2054));
    outputs(1183) <= not(layer6_outputs(740));
    outputs(1184) <= not(layer6_outputs(1547));
    outputs(1185) <= (layer6_outputs(527)) and (layer6_outputs(2144));
    outputs(1186) <= not(layer6_outputs(1854));
    outputs(1187) <= not(layer6_outputs(2063));
    outputs(1188) <= not(layer6_outputs(1881));
    outputs(1189) <= (layer6_outputs(1060)) xor (layer6_outputs(532));
    outputs(1190) <= layer6_outputs(2308);
    outputs(1191) <= layer6_outputs(290);
    outputs(1192) <= not((layer6_outputs(1577)) xor (layer6_outputs(1076)));
    outputs(1193) <= layer6_outputs(1253);
    outputs(1194) <= layer6_outputs(991);
    outputs(1195) <= layer6_outputs(2499);
    outputs(1196) <= not(layer6_outputs(280));
    outputs(1197) <= not(layer6_outputs(1099));
    outputs(1198) <= not((layer6_outputs(825)) xor (layer6_outputs(1277)));
    outputs(1199) <= not((layer6_outputs(207)) and (layer6_outputs(23)));
    outputs(1200) <= not((layer6_outputs(1992)) xor (layer6_outputs(2206)));
    outputs(1201) <= not(layer6_outputs(716));
    outputs(1202) <= (layer6_outputs(555)) and not (layer6_outputs(1523));
    outputs(1203) <= layer6_outputs(846);
    outputs(1204) <= (layer6_outputs(2519)) and not (layer6_outputs(2524));
    outputs(1205) <= layer6_outputs(185);
    outputs(1206) <= layer6_outputs(766);
    outputs(1207) <= not((layer6_outputs(1364)) xor (layer6_outputs(657)));
    outputs(1208) <= not(layer6_outputs(1921));
    outputs(1209) <= (layer6_outputs(2256)) xor (layer6_outputs(786));
    outputs(1210) <= not((layer6_outputs(525)) xor (layer6_outputs(1202)));
    outputs(1211) <= not((layer6_outputs(1783)) xor (layer6_outputs(2173)));
    outputs(1212) <= not((layer6_outputs(117)) or (layer6_outputs(121)));
    outputs(1213) <= not(layer6_outputs(2324));
    outputs(1214) <= (layer6_outputs(334)) xor (layer6_outputs(289));
    outputs(1215) <= not(layer6_outputs(541));
    outputs(1216) <= layer6_outputs(184);
    outputs(1217) <= not(layer6_outputs(639));
    outputs(1218) <= (layer6_outputs(75)) xor (layer6_outputs(1865));
    outputs(1219) <= not(layer6_outputs(2276));
    outputs(1220) <= (layer6_outputs(1707)) and not (layer6_outputs(1726));
    outputs(1221) <= not(layer6_outputs(1896));
    outputs(1222) <= layer6_outputs(1176);
    outputs(1223) <= layer6_outputs(524);
    outputs(1224) <= layer6_outputs(759);
    outputs(1225) <= layer6_outputs(307);
    outputs(1226) <= layer6_outputs(149);
    outputs(1227) <= layer6_outputs(1460);
    outputs(1228) <= layer6_outputs(113);
    outputs(1229) <= layer6_outputs(1698);
    outputs(1230) <= not((layer6_outputs(2190)) xor (layer6_outputs(1628)));
    outputs(1231) <= layer6_outputs(2558);
    outputs(1232) <= layer6_outputs(2127);
    outputs(1233) <= (layer6_outputs(2435)) xor (layer6_outputs(1252));
    outputs(1234) <= not(layer6_outputs(1119));
    outputs(1235) <= layer6_outputs(1226);
    outputs(1236) <= not(layer6_outputs(85));
    outputs(1237) <= (layer6_outputs(2146)) and not (layer6_outputs(969));
    outputs(1238) <= not(layer6_outputs(2017));
    outputs(1239) <= layer6_outputs(1949);
    outputs(1240) <= not(layer6_outputs(253));
    outputs(1241) <= not(layer6_outputs(202));
    outputs(1242) <= not(layer6_outputs(964));
    outputs(1243) <= not(layer6_outputs(1679)) or (layer6_outputs(1208));
    outputs(1244) <= not(layer6_outputs(1493));
    outputs(1245) <= layer6_outputs(504);
    outputs(1246) <= not(layer6_outputs(2253));
    outputs(1247) <= layer6_outputs(19);
    outputs(1248) <= layer6_outputs(111);
    outputs(1249) <= layer6_outputs(2242);
    outputs(1250) <= not(layer6_outputs(1048));
    outputs(1251) <= (layer6_outputs(717)) and not (layer6_outputs(2003));
    outputs(1252) <= not(layer6_outputs(417));
    outputs(1253) <= not((layer6_outputs(645)) xor (layer6_outputs(2502)));
    outputs(1254) <= not(layer6_outputs(693));
    outputs(1255) <= layer6_outputs(1927);
    outputs(1256) <= not(layer6_outputs(644));
    outputs(1257) <= not(layer6_outputs(2033));
    outputs(1258) <= not((layer6_outputs(1995)) xor (layer6_outputs(250)));
    outputs(1259) <= not(layer6_outputs(1831)) or (layer6_outputs(1864));
    outputs(1260) <= (layer6_outputs(1212)) xor (layer6_outputs(1733));
    outputs(1261) <= (layer6_outputs(39)) and (layer6_outputs(1446));
    outputs(1262) <= (layer6_outputs(2036)) and not (layer6_outputs(302));
    outputs(1263) <= layer6_outputs(832);
    outputs(1264) <= (layer6_outputs(2423)) xor (layer6_outputs(1134));
    outputs(1265) <= (layer6_outputs(249)) and (layer6_outputs(2527));
    outputs(1266) <= (layer6_outputs(1931)) and (layer6_outputs(375));
    outputs(1267) <= not((layer6_outputs(1953)) and (layer6_outputs(1307)));
    outputs(1268) <= not((layer6_outputs(2098)) or (layer6_outputs(1223)));
    outputs(1269) <= not(layer6_outputs(145));
    outputs(1270) <= layer6_outputs(2258);
    outputs(1271) <= layer6_outputs(580);
    outputs(1272) <= (layer6_outputs(2345)) and not (layer6_outputs(1563));
    outputs(1273) <= layer6_outputs(323);
    outputs(1274) <= not(layer6_outputs(1899));
    outputs(1275) <= (layer6_outputs(849)) and not (layer6_outputs(250));
    outputs(1276) <= (layer6_outputs(2479)) xor (layer6_outputs(1030));
    outputs(1277) <= (layer6_outputs(1851)) and not (layer6_outputs(1685));
    outputs(1278) <= not(layer6_outputs(1049));
    outputs(1279) <= (layer6_outputs(1415)) and (layer6_outputs(1390));
    outputs(1280) <= layer6_outputs(2477);
    outputs(1281) <= layer6_outputs(35);
    outputs(1282) <= not(layer6_outputs(1224));
    outputs(1283) <= not((layer6_outputs(2382)) xor (layer6_outputs(1671)));
    outputs(1284) <= not(layer6_outputs(871));
    outputs(1285) <= not(layer6_outputs(769));
    outputs(1286) <= layer6_outputs(2471);
    outputs(1287) <= (layer6_outputs(2245)) and not (layer6_outputs(641));
    outputs(1288) <= layer6_outputs(1357);
    outputs(1289) <= layer6_outputs(409);
    outputs(1290) <= layer6_outputs(2255);
    outputs(1291) <= (layer6_outputs(118)) or (layer6_outputs(1626));
    outputs(1292) <= (layer6_outputs(608)) xor (layer6_outputs(390));
    outputs(1293) <= not((layer6_outputs(1252)) xor (layer6_outputs(1807)));
    outputs(1294) <= (layer6_outputs(2401)) and not (layer6_outputs(2544));
    outputs(1295) <= layer6_outputs(1528);
    outputs(1296) <= layer6_outputs(1771);
    outputs(1297) <= not((layer6_outputs(335)) xor (layer6_outputs(40)));
    outputs(1298) <= not(layer6_outputs(2488));
    outputs(1299) <= (layer6_outputs(597)) xor (layer6_outputs(2433));
    outputs(1300) <= (layer6_outputs(1284)) and not (layer6_outputs(1990));
    outputs(1301) <= (layer6_outputs(471)) xor (layer6_outputs(1091));
    outputs(1302) <= not(layer6_outputs(484));
    outputs(1303) <= not(layer6_outputs(611)) or (layer6_outputs(1032));
    outputs(1304) <= not((layer6_outputs(883)) xor (layer6_outputs(2286)));
    outputs(1305) <= (layer6_outputs(2149)) xor (layer6_outputs(1369));
    outputs(1306) <= not(layer6_outputs(2126));
    outputs(1307) <= not((layer6_outputs(1000)) and (layer6_outputs(842)));
    outputs(1308) <= layer6_outputs(1383);
    outputs(1309) <= layer6_outputs(82);
    outputs(1310) <= (layer6_outputs(786)) and not (layer6_outputs(623));
    outputs(1311) <= not(layer6_outputs(1018));
    outputs(1312) <= layer6_outputs(1515);
    outputs(1313) <= layer6_outputs(2322);
    outputs(1314) <= (layer6_outputs(2111)) and not (layer6_outputs(902));
    outputs(1315) <= not((layer6_outputs(2451)) xor (layer6_outputs(2227)));
    outputs(1316) <= (layer6_outputs(1039)) and not (layer6_outputs(1491));
    outputs(1317) <= layer6_outputs(2269);
    outputs(1318) <= (layer6_outputs(2016)) xor (layer6_outputs(1647));
    outputs(1319) <= not((layer6_outputs(2312)) or (layer6_outputs(607)));
    outputs(1320) <= layer6_outputs(654);
    outputs(1321) <= layer6_outputs(82);
    outputs(1322) <= layer6_outputs(1898);
    outputs(1323) <= (layer6_outputs(453)) and not (layer6_outputs(1138));
    outputs(1324) <= not(layer6_outputs(2379));
    outputs(1325) <= not(layer6_outputs(1431));
    outputs(1326) <= (layer6_outputs(2450)) and not (layer6_outputs(176));
    outputs(1327) <= (layer6_outputs(2058)) xor (layer6_outputs(377));
    outputs(1328) <= not((layer6_outputs(1434)) xor (layer6_outputs(1730)));
    outputs(1329) <= not(layer6_outputs(1616));
    outputs(1330) <= not(layer6_outputs(1173));
    outputs(1331) <= (layer6_outputs(2553)) xor (layer6_outputs(1776));
    outputs(1332) <= not(layer6_outputs(1737));
    outputs(1333) <= not((layer6_outputs(931)) xor (layer6_outputs(2366)));
    outputs(1334) <= not((layer6_outputs(970)) xor (layer6_outputs(1831)));
    outputs(1335) <= layer6_outputs(365);
    outputs(1336) <= not((layer6_outputs(2525)) and (layer6_outputs(906)));
    outputs(1337) <= not((layer6_outputs(2326)) or (layer6_outputs(437)));
    outputs(1338) <= not((layer6_outputs(2146)) xor (layer6_outputs(1126)));
    outputs(1339) <= (layer6_outputs(2111)) or (layer6_outputs(175));
    outputs(1340) <= layer6_outputs(1428);
    outputs(1341) <= (layer6_outputs(1640)) and not (layer6_outputs(245));
    outputs(1342) <= not((layer6_outputs(593)) xor (layer6_outputs(2505)));
    outputs(1343) <= layer6_outputs(1004);
    outputs(1344) <= not((layer6_outputs(196)) xor (layer6_outputs(365)));
    outputs(1345) <= (layer6_outputs(2043)) xor (layer6_outputs(2504));
    outputs(1346) <= not((layer6_outputs(95)) xor (layer6_outputs(1089)));
    outputs(1347) <= layer6_outputs(504);
    outputs(1348) <= layer6_outputs(1676);
    outputs(1349) <= layer6_outputs(2050);
    outputs(1350) <= not(layer6_outputs(946));
    outputs(1351) <= (layer6_outputs(752)) xor (layer6_outputs(189));
    outputs(1352) <= layer6_outputs(2332);
    outputs(1353) <= layer6_outputs(2085);
    outputs(1354) <= not(layer6_outputs(1617));
    outputs(1355) <= not(layer6_outputs(1797));
    outputs(1356) <= (layer6_outputs(674)) and not (layer6_outputs(2123));
    outputs(1357) <= (layer6_outputs(620)) and (layer6_outputs(888));
    outputs(1358) <= not(layer6_outputs(1793));
    outputs(1359) <= layer6_outputs(505);
    outputs(1360) <= not((layer6_outputs(1723)) xor (layer6_outputs(50)));
    outputs(1361) <= (layer6_outputs(1967)) and not (layer6_outputs(1373));
    outputs(1362) <= layer6_outputs(126);
    outputs(1363) <= not((layer6_outputs(973)) xor (layer6_outputs(564)));
    outputs(1364) <= not(layer6_outputs(1949));
    outputs(1365) <= (layer6_outputs(2334)) xor (layer6_outputs(58));
    outputs(1366) <= not(layer6_outputs(2251));
    outputs(1367) <= not((layer6_outputs(331)) xor (layer6_outputs(1457)));
    outputs(1368) <= (layer6_outputs(1988)) and not (layer6_outputs(2247));
    outputs(1369) <= not(layer6_outputs(2067));
    outputs(1370) <= not((layer6_outputs(1752)) xor (layer6_outputs(319)));
    outputs(1371) <= not(layer6_outputs(1287));
    outputs(1372) <= not(layer6_outputs(838)) or (layer6_outputs(1260));
    outputs(1373) <= (layer6_outputs(2202)) xor (layer6_outputs(1251));
    outputs(1374) <= (layer6_outputs(91)) and not (layer6_outputs(16));
    outputs(1375) <= (layer6_outputs(803)) xor (layer6_outputs(959));
    outputs(1376) <= not(layer6_outputs(2026));
    outputs(1377) <= not(layer6_outputs(623));
    outputs(1378) <= not(layer6_outputs(2356));
    outputs(1379) <= not((layer6_outputs(2164)) xor (layer6_outputs(2482)));
    outputs(1380) <= layer6_outputs(487);
    outputs(1381) <= layer6_outputs(45);
    outputs(1382) <= not(layer6_outputs(1604)) or (layer6_outputs(526));
    outputs(1383) <= layer6_outputs(1914);
    outputs(1384) <= layer6_outputs(1889);
    outputs(1385) <= layer6_outputs(503);
    outputs(1386) <= not(layer6_outputs(1399));
    outputs(1387) <= (layer6_outputs(851)) and (layer6_outputs(1783));
    outputs(1388) <= layer6_outputs(1991);
    outputs(1389) <= not((layer6_outputs(478)) xor (layer6_outputs(188)));
    outputs(1390) <= layer6_outputs(1724);
    outputs(1391) <= not((layer6_outputs(1654)) xor (layer6_outputs(1525)));
    outputs(1392) <= (layer6_outputs(18)) and not (layer6_outputs(1398));
    outputs(1393) <= layer6_outputs(169);
    outputs(1394) <= not((layer6_outputs(589)) or (layer6_outputs(1657)));
    outputs(1395) <= (layer6_outputs(776)) xor (layer6_outputs(1079));
    outputs(1396) <= layer6_outputs(88);
    outputs(1397) <= (layer6_outputs(2015)) and (layer6_outputs(241));
    outputs(1398) <= not((layer6_outputs(1326)) and (layer6_outputs(2372)));
    outputs(1399) <= (layer6_outputs(713)) and not (layer6_outputs(110));
    outputs(1400) <= not(layer6_outputs(621));
    outputs(1401) <= layer6_outputs(1650);
    outputs(1402) <= not(layer6_outputs(1381));
    outputs(1403) <= not(layer6_outputs(1932));
    outputs(1404) <= not((layer6_outputs(517)) xor (layer6_outputs(1410)));
    outputs(1405) <= not((layer6_outputs(2011)) xor (layer6_outputs(713)));
    outputs(1406) <= not(layer6_outputs(1257));
    outputs(1407) <= layer6_outputs(419);
    outputs(1408) <= (layer6_outputs(702)) xor (layer6_outputs(677));
    outputs(1409) <= not(layer6_outputs(1598));
    outputs(1410) <= layer6_outputs(1711);
    outputs(1411) <= (layer6_outputs(1828)) xor (layer6_outputs(724));
    outputs(1412) <= layer6_outputs(1630);
    outputs(1413) <= layer6_outputs(156);
    outputs(1414) <= not(layer6_outputs(1741));
    outputs(1415) <= not(layer6_outputs(2062)) or (layer6_outputs(1040));
    outputs(1416) <= not((layer6_outputs(431)) or (layer6_outputs(1435)));
    outputs(1417) <= not(layer6_outputs(728));
    outputs(1418) <= layer6_outputs(680);
    outputs(1419) <= (layer6_outputs(508)) and not (layer6_outputs(1977));
    outputs(1420) <= not((layer6_outputs(2447)) or (layer6_outputs(863)));
    outputs(1421) <= (layer6_outputs(357)) and not (layer6_outputs(392));
    outputs(1422) <= (layer6_outputs(291)) and (layer6_outputs(2044));
    outputs(1423) <= not((layer6_outputs(821)) and (layer6_outputs(1506)));
    outputs(1424) <= not((layer6_outputs(581)) or (layer6_outputs(718)));
    outputs(1425) <= layer6_outputs(2160);
    outputs(1426) <= not((layer6_outputs(2501)) or (layer6_outputs(2463)));
    outputs(1427) <= layer6_outputs(741);
    outputs(1428) <= not((layer6_outputs(1748)) or (layer6_outputs(1959)));
    outputs(1429) <= layer6_outputs(1439);
    outputs(1430) <= not(layer6_outputs(1728));
    outputs(1431) <= layer6_outputs(422);
    outputs(1432) <= not((layer6_outputs(298)) xor (layer6_outputs(526)));
    outputs(1433) <= not(layer6_outputs(1157));
    outputs(1434) <= (layer6_outputs(2215)) and not (layer6_outputs(1649));
    outputs(1435) <= (layer6_outputs(1171)) and not (layer6_outputs(259));
    outputs(1436) <= not((layer6_outputs(228)) xor (layer6_outputs(579)));
    outputs(1437) <= (layer6_outputs(1259)) xor (layer6_outputs(790));
    outputs(1438) <= layer6_outputs(2419);
    outputs(1439) <= not((layer6_outputs(2201)) xor (layer6_outputs(1945)));
    outputs(1440) <= (layer6_outputs(510)) xor (layer6_outputs(486));
    outputs(1441) <= layer6_outputs(1706);
    outputs(1442) <= layer6_outputs(421);
    outputs(1443) <= layer6_outputs(562);
    outputs(1444) <= layer6_outputs(2175);
    outputs(1445) <= not(layer6_outputs(880)) or (layer6_outputs(2151));
    outputs(1446) <= layer6_outputs(186);
    outputs(1447) <= layer6_outputs(1199);
    outputs(1448) <= (layer6_outputs(1600)) xor (layer6_outputs(691));
    outputs(1449) <= not((layer6_outputs(462)) xor (layer6_outputs(1705)));
    outputs(1450) <= not(layer6_outputs(1103));
    outputs(1451) <= not(layer6_outputs(840)) or (layer6_outputs(2177));
    outputs(1452) <= not(layer6_outputs(1709));
    outputs(1453) <= layer6_outputs(2004);
    outputs(1454) <= not(layer6_outputs(2166));
    outputs(1455) <= layer6_outputs(1042);
    outputs(1456) <= not((layer6_outputs(1100)) xor (layer6_outputs(867)));
    outputs(1457) <= (layer6_outputs(1703)) and (layer6_outputs(1715));
    outputs(1458) <= not(layer6_outputs(2431));
    outputs(1459) <= not(layer6_outputs(507));
    outputs(1460) <= (layer6_outputs(1536)) xor (layer6_outputs(1999));
    outputs(1461) <= not((layer6_outputs(1297)) xor (layer6_outputs(1036)));
    outputs(1462) <= (layer6_outputs(136)) xor (layer6_outputs(570));
    outputs(1463) <= layer6_outputs(1101);
    outputs(1464) <= layer6_outputs(986);
    outputs(1465) <= layer6_outputs(2301);
    outputs(1466) <= (layer6_outputs(2167)) and (layer6_outputs(679));
    outputs(1467) <= (layer6_outputs(533)) xor (layer6_outputs(307));
    outputs(1468) <= not((layer6_outputs(1644)) xor (layer6_outputs(2107)));
    outputs(1469) <= layer6_outputs(1954);
    outputs(1470) <= (layer6_outputs(2215)) and (layer6_outputs(587));
    outputs(1471) <= not(layer6_outputs(905));
    outputs(1472) <= layer6_outputs(1658);
    outputs(1473) <= not((layer6_outputs(1786)) xor (layer6_outputs(1983)));
    outputs(1474) <= not((layer6_outputs(1232)) or (layer6_outputs(2290)));
    outputs(1475) <= (layer6_outputs(227)) and (layer6_outputs(140));
    outputs(1476) <= not(layer6_outputs(2148));
    outputs(1477) <= not((layer6_outputs(1338)) or (layer6_outputs(884)));
    outputs(1478) <= not(layer6_outputs(369));
    outputs(1479) <= layer6_outputs(2537);
    outputs(1480) <= not(layer6_outputs(1222));
    outputs(1481) <= layer6_outputs(953);
    outputs(1482) <= not((layer6_outputs(1528)) xor (layer6_outputs(828)));
    outputs(1483) <= not(layer6_outputs(534));
    outputs(1484) <= (layer6_outputs(135)) or (layer6_outputs(977));
    outputs(1485) <= not(layer6_outputs(701));
    outputs(1486) <= layer6_outputs(1158);
    outputs(1487) <= not((layer6_outputs(812)) xor (layer6_outputs(121)));
    outputs(1488) <= not((layer6_outputs(1242)) xor (layer6_outputs(1059)));
    outputs(1489) <= layer6_outputs(2013);
    outputs(1490) <= not((layer6_outputs(2402)) xor (layer6_outputs(1753)));
    outputs(1491) <= layer6_outputs(1595);
    outputs(1492) <= layer6_outputs(137);
    outputs(1493) <= layer6_outputs(2155);
    outputs(1494) <= not(layer6_outputs(2456));
    outputs(1495) <= not(layer6_outputs(2209));
    outputs(1496) <= (layer6_outputs(460)) xor (layer6_outputs(2319));
    outputs(1497) <= (layer6_outputs(1477)) and not (layer6_outputs(709));
    outputs(1498) <= not(layer6_outputs(1981));
    outputs(1499) <= layer6_outputs(566);
    outputs(1500) <= not((layer6_outputs(316)) xor (layer6_outputs(657)));
    outputs(1501) <= not((layer6_outputs(2090)) xor (layer6_outputs(1308)));
    outputs(1502) <= not(layer6_outputs(2544));
    outputs(1503) <= not(layer6_outputs(728)) or (layer6_outputs(1081));
    outputs(1504) <= (layer6_outputs(1625)) xor (layer6_outputs(1981));
    outputs(1505) <= layer6_outputs(1519);
    outputs(1506) <= not(layer6_outputs(1203));
    outputs(1507) <= layer6_outputs(674);
    outputs(1508) <= not(layer6_outputs(920));
    outputs(1509) <= layer6_outputs(1725);
    outputs(1510) <= not(layer6_outputs(255));
    outputs(1511) <= not(layer6_outputs(1461));
    outputs(1512) <= (layer6_outputs(303)) xor (layer6_outputs(35));
    outputs(1513) <= not((layer6_outputs(1947)) or (layer6_outputs(725)));
    outputs(1514) <= layer6_outputs(2018);
    outputs(1515) <= not((layer6_outputs(381)) or (layer6_outputs(2351)));
    outputs(1516) <= (layer6_outputs(1505)) xor (layer6_outputs(1891));
    outputs(1517) <= not((layer6_outputs(1062)) and (layer6_outputs(2391)));
    outputs(1518) <= not(layer6_outputs(1394));
    outputs(1519) <= (layer6_outputs(873)) and not (layer6_outputs(199));
    outputs(1520) <= not(layer6_outputs(22));
    outputs(1521) <= (layer6_outputs(537)) xor (layer6_outputs(1809));
    outputs(1522) <= layer6_outputs(1195);
    outputs(1523) <= not(layer6_outputs(1456));
    outputs(1524) <= layer6_outputs(290);
    outputs(1525) <= not(layer6_outputs(416));
    outputs(1526) <= layer6_outputs(1428);
    outputs(1527) <= layer6_outputs(411);
    outputs(1528) <= not((layer6_outputs(1102)) xor (layer6_outputs(1843)));
    outputs(1529) <= not((layer6_outputs(1298)) or (layer6_outputs(678)));
    outputs(1530) <= not(layer6_outputs(819));
    outputs(1531) <= not(layer6_outputs(1330));
    outputs(1532) <= (layer6_outputs(1339)) xor (layer6_outputs(1215));
    outputs(1533) <= (layer6_outputs(2434)) and not (layer6_outputs(1394));
    outputs(1534) <= layer6_outputs(1950);
    outputs(1535) <= not(layer6_outputs(340));
    outputs(1536) <= not((layer6_outputs(756)) xor (layer6_outputs(897)));
    outputs(1537) <= layer6_outputs(1964);
    outputs(1538) <= (layer6_outputs(215)) and (layer6_outputs(2416));
    outputs(1539) <= layer6_outputs(1347);
    outputs(1540) <= not((layer6_outputs(1591)) xor (layer6_outputs(1476)));
    outputs(1541) <= layer6_outputs(1994);
    outputs(1542) <= not(layer6_outputs(1437));
    outputs(1543) <= layer6_outputs(2283);
    outputs(1544) <= layer6_outputs(2335);
    outputs(1545) <= not((layer6_outputs(2354)) or (layer6_outputs(2425)));
    outputs(1546) <= not(layer6_outputs(1537));
    outputs(1547) <= layer6_outputs(2528);
    outputs(1548) <= (layer6_outputs(2555)) and not (layer6_outputs(2005));
    outputs(1549) <= not(layer6_outputs(1124));
    outputs(1550) <= layer6_outputs(1691);
    outputs(1551) <= layer6_outputs(1069);
    outputs(1552) <= (layer6_outputs(2303)) and (layer6_outputs(495));
    outputs(1553) <= not(layer6_outputs(1473)) or (layer6_outputs(695));
    outputs(1554) <= not(layer6_outputs(646));
    outputs(1555) <= not(layer6_outputs(1846));
    outputs(1556) <= layer6_outputs(1968);
    outputs(1557) <= (layer6_outputs(2188)) and (layer6_outputs(861));
    outputs(1558) <= layer6_outputs(1220);
    outputs(1559) <= not(layer6_outputs(818));
    outputs(1560) <= (layer6_outputs(790)) and not (layer6_outputs(1801));
    outputs(1561) <= layer6_outputs(2075);
    outputs(1562) <= not(layer6_outputs(1228));
    outputs(1563) <= layer6_outputs(2410);
    outputs(1564) <= layer6_outputs(746);
    outputs(1565) <= (layer6_outputs(440)) and not (layer6_outputs(781));
    outputs(1566) <= not((layer6_outputs(1984)) or (layer6_outputs(602)));
    outputs(1567) <= layer6_outputs(464);
    outputs(1568) <= layer6_outputs(179);
    outputs(1569) <= (layer6_outputs(34)) and not (layer6_outputs(703));
    outputs(1570) <= (layer6_outputs(251)) and not (layer6_outputs(1449));
    outputs(1571) <= layer6_outputs(416);
    outputs(1572) <= (layer6_outputs(348)) and (layer6_outputs(2132));
    outputs(1573) <= not(layer6_outputs(436));
    outputs(1574) <= (layer6_outputs(2221)) and not (layer6_outputs(755));
    outputs(1575) <= layer6_outputs(2529);
    outputs(1576) <= not(layer6_outputs(1907));
    outputs(1577) <= (layer6_outputs(482)) and not (layer6_outputs(211));
    outputs(1578) <= (layer6_outputs(1740)) and (layer6_outputs(1257));
    outputs(1579) <= (layer6_outputs(1482)) and (layer6_outputs(665));
    outputs(1580) <= layer6_outputs(1870);
    outputs(1581) <= (layer6_outputs(2504)) and not (layer6_outputs(192));
    outputs(1582) <= not((layer6_outputs(1775)) or (layer6_outputs(1445)));
    outputs(1583) <= (layer6_outputs(892)) and not (layer6_outputs(1151));
    outputs(1584) <= layer6_outputs(2483);
    outputs(1585) <= not(layer6_outputs(187));
    outputs(1586) <= not(layer6_outputs(1082));
    outputs(1587) <= (layer6_outputs(2156)) and not (layer6_outputs(343));
    outputs(1588) <= not((layer6_outputs(1549)) xor (layer6_outputs(1290)));
    outputs(1589) <= (layer6_outputs(1566)) and not (layer6_outputs(591));
    outputs(1590) <= layer6_outputs(1312);
    outputs(1591) <= layer6_outputs(369);
    outputs(1592) <= not(layer6_outputs(1607)) or (layer6_outputs(466));
    outputs(1593) <= layer6_outputs(1556);
    outputs(1594) <= layer6_outputs(689);
    outputs(1595) <= not((layer6_outputs(1301)) or (layer6_outputs(1183)));
    outputs(1596) <= not((layer6_outputs(1806)) xor (layer6_outputs(1209)));
    outputs(1597) <= not(layer6_outputs(371));
    outputs(1598) <= layer6_outputs(1373);
    outputs(1599) <= not((layer6_outputs(385)) xor (layer6_outputs(2303)));
    outputs(1600) <= (layer6_outputs(734)) and not (layer6_outputs(690));
    outputs(1601) <= not(layer6_outputs(990)) or (layer6_outputs(1571));
    outputs(1602) <= not((layer6_outputs(391)) or (layer6_outputs(1853)));
    outputs(1603) <= layer6_outputs(695);
    outputs(1604) <= layer6_outputs(1628);
    outputs(1605) <= layer6_outputs(23);
    outputs(1606) <= layer6_outputs(2041);
    outputs(1607) <= not(layer6_outputs(151));
    outputs(1608) <= not((layer6_outputs(1574)) xor (layer6_outputs(1984)));
    outputs(1609) <= not(layer6_outputs(2131));
    outputs(1610) <= not(layer6_outputs(1137));
    outputs(1611) <= layer6_outputs(488);
    outputs(1612) <= (layer6_outputs(1449)) xor (layer6_outputs(2459));
    outputs(1613) <= not(layer6_outputs(514));
    outputs(1614) <= not(layer6_outputs(2371));
    outputs(1615) <= not(layer6_outputs(621));
    outputs(1616) <= layer6_outputs(1980);
    outputs(1617) <= (layer6_outputs(624)) and not (layer6_outputs(563));
    outputs(1618) <= (layer6_outputs(1484)) or (layer6_outputs(578));
    outputs(1619) <= (layer6_outputs(69)) and not (layer6_outputs(1475));
    outputs(1620) <= layer6_outputs(1649);
    outputs(1621) <= layer6_outputs(1225);
    outputs(1622) <= (layer6_outputs(811)) and (layer6_outputs(242));
    outputs(1623) <= not(layer6_outputs(1531));
    outputs(1624) <= not(layer6_outputs(2278));
    outputs(1625) <= not(layer6_outputs(350));
    outputs(1626) <= (layer6_outputs(1021)) and (layer6_outputs(341));
    outputs(1627) <= layer6_outputs(1900);
    outputs(1628) <= layer6_outputs(2199);
    outputs(1629) <= layer6_outputs(914);
    outputs(1630) <= layer6_outputs(2529);
    outputs(1631) <= not(layer6_outputs(1664));
    outputs(1632) <= not(layer6_outputs(2275));
    outputs(1633) <= not((layer6_outputs(1317)) or (layer6_outputs(2514)));
    outputs(1634) <= not(layer6_outputs(2351));
    outputs(1635) <= not(layer6_outputs(1382));
    outputs(1636) <= (layer6_outputs(1510)) xor (layer6_outputs(2144));
    outputs(1637) <= not((layer6_outputs(395)) xor (layer6_outputs(1560)));
    outputs(1638) <= not(layer6_outputs(1596));
    outputs(1639) <= layer6_outputs(1430);
    outputs(1640) <= layer6_outputs(347);
    outputs(1641) <= not((layer6_outputs(13)) or (layer6_outputs(195)));
    outputs(1642) <= not((layer6_outputs(2088)) or (layer6_outputs(352)));
    outputs(1643) <= layer6_outputs(853);
    outputs(1644) <= not(layer6_outputs(785));
    outputs(1645) <= layer6_outputs(957);
    outputs(1646) <= not(layer6_outputs(518));
    outputs(1647) <= not((layer6_outputs(79)) xor (layer6_outputs(2056)));
    outputs(1648) <= not((layer6_outputs(1466)) xor (layer6_outputs(1890)));
    outputs(1649) <= not(layer6_outputs(452));
    outputs(1650) <= (layer6_outputs(1876)) or (layer6_outputs(1288));
    outputs(1651) <= layer6_outputs(568);
    outputs(1652) <= layer6_outputs(806);
    outputs(1653) <= (layer6_outputs(1637)) and (layer6_outputs(1663));
    outputs(1654) <= not(layer6_outputs(163));
    outputs(1655) <= not((layer6_outputs(1567)) or (layer6_outputs(58)));
    outputs(1656) <= (layer6_outputs(1136)) and not (layer6_outputs(1340));
    outputs(1657) <= not((layer6_outputs(2122)) or (layer6_outputs(2299)));
    outputs(1658) <= not(layer6_outputs(162));
    outputs(1659) <= (layer6_outputs(694)) xor (layer6_outputs(1053));
    outputs(1660) <= (layer6_outputs(2046)) and not (layer6_outputs(2241));
    outputs(1661) <= not(layer6_outputs(1265));
    outputs(1662) <= (layer6_outputs(190)) and (layer6_outputs(668));
    outputs(1663) <= not((layer6_outputs(1158)) or (layer6_outputs(2491)));
    outputs(1664) <= layer6_outputs(240);
    outputs(1665) <= not((layer6_outputs(1787)) or (layer6_outputs(2255)));
    outputs(1666) <= not((layer6_outputs(192)) or (layer6_outputs(368)));
    outputs(1667) <= layer6_outputs(1794);
    outputs(1668) <= (layer6_outputs(2000)) or (layer6_outputs(908));
    outputs(1669) <= (layer6_outputs(1679)) and (layer6_outputs(422));
    outputs(1670) <= (layer6_outputs(423)) and not (layer6_outputs(1176));
    outputs(1671) <= not(layer6_outputs(1052));
    outputs(1672) <= not(layer6_outputs(1939));
    outputs(1673) <= layer6_outputs(1961);
    outputs(1674) <= not(layer6_outputs(2323));
    outputs(1675) <= not(layer6_outputs(375));
    outputs(1676) <= (layer6_outputs(2472)) and (layer6_outputs(1878));
    outputs(1677) <= (layer6_outputs(2407)) or (layer6_outputs(1636));
    outputs(1678) <= (layer6_outputs(1016)) xor (layer6_outputs(756));
    outputs(1679) <= layer6_outputs(1386);
    outputs(1680) <= not((layer6_outputs(1146)) or (layer6_outputs(1426)));
    outputs(1681) <= not(layer6_outputs(152));
    outputs(1682) <= not(layer6_outputs(1718));
    outputs(1683) <= (layer6_outputs(1096)) xor (layer6_outputs(1102));
    outputs(1684) <= layer6_outputs(364);
    outputs(1685) <= layer6_outputs(206);
    outputs(1686) <= not((layer6_outputs(1814)) and (layer6_outputs(1661)));
    outputs(1687) <= layer6_outputs(204);
    outputs(1688) <= (layer6_outputs(1960)) and (layer6_outputs(605));
    outputs(1689) <= (layer6_outputs(851)) and not (layer6_outputs(285));
    outputs(1690) <= not((layer6_outputs(1139)) xor (layer6_outputs(1026)));
    outputs(1691) <= not(layer6_outputs(1837));
    outputs(1692) <= layer6_outputs(280);
    outputs(1693) <= not((layer6_outputs(4)) xor (layer6_outputs(2534)));
    outputs(1694) <= (layer6_outputs(962)) xor (layer6_outputs(1548));
    outputs(1695) <= layer6_outputs(2311);
    outputs(1696) <= (layer6_outputs(800)) and (layer6_outputs(928));
    outputs(1697) <= layer6_outputs(259);
    outputs(1698) <= not((layer6_outputs(177)) xor (layer6_outputs(532)));
    outputs(1699) <= layer6_outputs(1952);
    outputs(1700) <= not(layer6_outputs(1106));
    outputs(1701) <= layer6_outputs(1588);
    outputs(1702) <= (layer6_outputs(2156)) and (layer6_outputs(603));
    outputs(1703) <= not(layer6_outputs(1671));
    outputs(1704) <= layer6_outputs(420);
    outputs(1705) <= layer6_outputs(2435);
    outputs(1706) <= (layer6_outputs(1131)) and (layer6_outputs(1300));
    outputs(1707) <= not(layer6_outputs(2114));
    outputs(1708) <= layer6_outputs(1482);
    outputs(1709) <= not((layer6_outputs(2207)) xor (layer6_outputs(263)));
    outputs(1710) <= layer6_outputs(489);
    outputs(1711) <= layer6_outputs(913);
    outputs(1712) <= not((layer6_outputs(881)) and (layer6_outputs(1928)));
    outputs(1713) <= layer6_outputs(512);
    outputs(1714) <= (layer6_outputs(1625)) and not (layer6_outputs(1093));
    outputs(1715) <= layer6_outputs(590);
    outputs(1716) <= (layer6_outputs(1832)) and not (layer6_outputs(556));
    outputs(1717) <= not((layer6_outputs(731)) xor (layer6_outputs(1130)));
    outputs(1718) <= layer6_outputs(1393);
    outputs(1719) <= layer6_outputs(2451);
    outputs(1720) <= (layer6_outputs(2165)) and (layer6_outputs(474));
    outputs(1721) <= not((layer6_outputs(1161)) or (layer6_outputs(1780)));
    outputs(1722) <= not(layer6_outputs(1315));
    outputs(1723) <= not((layer6_outputs(783)) or (layer6_outputs(2138)));
    outputs(1724) <= (layer6_outputs(1652)) and not (layer6_outputs(198));
    outputs(1725) <= layer6_outputs(2557);
    outputs(1726) <= not((layer6_outputs(1582)) xor (layer6_outputs(2295)));
    outputs(1727) <= layer6_outputs(517);
    outputs(1728) <= not((layer6_outputs(1757)) xor (layer6_outputs(730)));
    outputs(1729) <= layer6_outputs(2187);
    outputs(1730) <= (layer6_outputs(2057)) and not (layer6_outputs(154));
    outputs(1731) <= not(layer6_outputs(2162));
    outputs(1732) <= layer6_outputs(1892);
    outputs(1733) <= (layer6_outputs(2104)) xor (layer6_outputs(38));
    outputs(1734) <= (layer6_outputs(2494)) xor (layer6_outputs(1848));
    outputs(1735) <= not(layer6_outputs(2501));
    outputs(1736) <= not(layer6_outputs(1255));
    outputs(1737) <= layer6_outputs(477);
    outputs(1738) <= layer6_outputs(1660);
    outputs(1739) <= layer6_outputs(1109);
    outputs(1740) <= layer6_outputs(839);
    outputs(1741) <= not(layer6_outputs(1200));
    outputs(1742) <= not(layer6_outputs(556));
    outputs(1743) <= (layer6_outputs(1372)) and (layer6_outputs(1015));
    outputs(1744) <= layer6_outputs(1774);
    outputs(1745) <= not((layer6_outputs(106)) xor (layer6_outputs(2060)));
    outputs(1746) <= not(layer6_outputs(182));
    outputs(1747) <= (layer6_outputs(2459)) xor (layer6_outputs(214));
    outputs(1748) <= (layer6_outputs(252)) xor (layer6_outputs(2342));
    outputs(1749) <= not(layer6_outputs(286));
    outputs(1750) <= layer6_outputs(628);
    outputs(1751) <= not(layer6_outputs(1716)) or (layer6_outputs(1789));
    outputs(1752) <= (layer6_outputs(1824)) xor (layer6_outputs(1887));
    outputs(1753) <= not((layer6_outputs(1576)) or (layer6_outputs(1727)));
    outputs(1754) <= (layer6_outputs(947)) and not (layer6_outputs(1618));
    outputs(1755) <= layer6_outputs(1867);
    outputs(1756) <= layer6_outputs(1743);
    outputs(1757) <= not((layer6_outputs(1978)) xor (layer6_outputs(2259)));
    outputs(1758) <= layer6_outputs(1566);
    outputs(1759) <= not((layer6_outputs(1924)) or (layer6_outputs(211)));
    outputs(1760) <= not((layer6_outputs(265)) or (layer6_outputs(520)));
    outputs(1761) <= (layer6_outputs(299)) and (layer6_outputs(251));
    outputs(1762) <= (layer6_outputs(1535)) and (layer6_outputs(1172));
    outputs(1763) <= not(layer6_outputs(457));
    outputs(1764) <= not(layer6_outputs(2507));
    outputs(1765) <= (layer6_outputs(1429)) xor (layer6_outputs(506));
    outputs(1766) <= layer6_outputs(1623);
    outputs(1767) <= layer6_outputs(969);
    outputs(1768) <= not(layer6_outputs(2009));
    outputs(1769) <= not(layer6_outputs(2381));
    outputs(1770) <= not(layer6_outputs(2432));
    outputs(1771) <= not(layer6_outputs(918));
    outputs(1772) <= (layer6_outputs(408)) xor (layer6_outputs(814));
    outputs(1773) <= not(layer6_outputs(1775));
    outputs(1774) <= (layer6_outputs(696)) and (layer6_outputs(1316));
    outputs(1775) <= not(layer6_outputs(1243));
    outputs(1776) <= (layer6_outputs(717)) and not (layer6_outputs(181));
    outputs(1777) <= not(layer6_outputs(6));
    outputs(1778) <= not(layer6_outputs(1673));
    outputs(1779) <= not((layer6_outputs(1310)) or (layer6_outputs(1974)));
    outputs(1780) <= layer6_outputs(1586);
    outputs(1781) <= not((layer6_outputs(1362)) xor (layer6_outputs(484)));
    outputs(1782) <= not(layer6_outputs(9));
    outputs(1783) <= layer6_outputs(428);
    outputs(1784) <= not((layer6_outputs(2294)) or (layer6_outputs(622)));
    outputs(1785) <= (layer6_outputs(950)) and not (layer6_outputs(752));
    outputs(1786) <= not(layer6_outputs(2280));
    outputs(1787) <= layer6_outputs(968);
    outputs(1788) <= (layer6_outputs(144)) and (layer6_outputs(2475));
    outputs(1789) <= not((layer6_outputs(1546)) xor (layer6_outputs(2428)));
    outputs(1790) <= not(layer6_outputs(2141));
    outputs(1791) <= layer6_outputs(1587);
    outputs(1792) <= layer6_outputs(233);
    outputs(1793) <= not(layer6_outputs(2532));
    outputs(1794) <= not(layer6_outputs(1605)) or (layer6_outputs(742));
    outputs(1795) <= layer6_outputs(1380);
    outputs(1796) <= layer6_outputs(1544);
    outputs(1797) <= (layer6_outputs(2222)) and not (layer6_outputs(2221));
    outputs(1798) <= not(layer6_outputs(2444));
    outputs(1799) <= (layer6_outputs(1325)) xor (layer6_outputs(1056));
    outputs(1800) <= (layer6_outputs(2176)) and not (layer6_outputs(1611));
    outputs(1801) <= layer6_outputs(848);
    outputs(1802) <= layer6_outputs(339);
    outputs(1803) <= layer6_outputs(6);
    outputs(1804) <= not(layer6_outputs(976));
    outputs(1805) <= layer6_outputs(939);
    outputs(1806) <= (layer6_outputs(322)) and not (layer6_outputs(90));
    outputs(1807) <= (layer6_outputs(2370)) and (layer6_outputs(2240));
    outputs(1808) <= not(layer6_outputs(1454));
    outputs(1809) <= (layer6_outputs(2327)) and (layer6_outputs(1803));
    outputs(1810) <= (layer6_outputs(1772)) xor (layer6_outputs(1059));
    outputs(1811) <= (layer6_outputs(531)) xor (layer6_outputs(137));
    outputs(1812) <= (layer6_outputs(2063)) and not (layer6_outputs(1240));
    outputs(1813) <= not(layer6_outputs(1275)) or (layer6_outputs(2149));
    outputs(1814) <= layer6_outputs(479);
    outputs(1815) <= not(layer6_outputs(414));
    outputs(1816) <= not(layer6_outputs(134));
    outputs(1817) <= layer6_outputs(2088);
    outputs(1818) <= not(layer6_outputs(1046));
    outputs(1819) <= (layer6_outputs(1715)) and (layer6_outputs(1606));
    outputs(1820) <= not(layer6_outputs(2489));
    outputs(1821) <= (layer6_outputs(1953)) and (layer6_outputs(2293));
    outputs(1822) <= not(layer6_outputs(1979));
    outputs(1823) <= (layer6_outputs(1452)) xor (layer6_outputs(453));
    outputs(1824) <= layer6_outputs(939);
    outputs(1825) <= layer6_outputs(1788);
    outputs(1826) <= not(layer6_outputs(424));
    outputs(1827) <= not(layer6_outputs(1391));
    outputs(1828) <= layer6_outputs(1398);
    outputs(1829) <= (layer6_outputs(1629)) and (layer6_outputs(1842));
    outputs(1830) <= layer6_outputs(2265);
    outputs(1831) <= (layer6_outputs(330)) xor (layer6_outputs(1875));
    outputs(1832) <= not((layer6_outputs(272)) or (layer6_outputs(725)));
    outputs(1833) <= (layer6_outputs(399)) xor (layer6_outputs(1269));
    outputs(1834) <= not(layer6_outputs(2449));
    outputs(1835) <= (layer6_outputs(844)) and not (layer6_outputs(574));
    outputs(1836) <= not((layer6_outputs(1692)) or (layer6_outputs(2072)));
    outputs(1837) <= not(layer6_outputs(586));
    outputs(1838) <= (layer6_outputs(1897)) and (layer6_outputs(142));
    outputs(1839) <= (layer6_outputs(13)) or (layer6_outputs(1736));
    outputs(1840) <= layer6_outputs(366);
    outputs(1841) <= not((layer6_outputs(1469)) xor (layer6_outputs(771)));
    outputs(1842) <= not(layer6_outputs(842));
    outputs(1843) <= not((layer6_outputs(1486)) xor (layer6_outputs(2446)));
    outputs(1844) <= (layer6_outputs(2495)) and not (layer6_outputs(543));
    outputs(1845) <= not((layer6_outputs(1067)) or (layer6_outputs(2218)));
    outputs(1846) <= not(layer6_outputs(614)) or (layer6_outputs(2147));
    outputs(1847) <= layer6_outputs(1786);
    outputs(1848) <= not(layer6_outputs(804));
    outputs(1849) <= layer6_outputs(1035);
    outputs(1850) <= not((layer6_outputs(904)) or (layer6_outputs(2035)));
    outputs(1851) <= (layer6_outputs(1392)) and not (layer6_outputs(2072));
    outputs(1852) <= not(layer6_outputs(320));
    outputs(1853) <= not(layer6_outputs(1413));
    outputs(1854) <= not((layer6_outputs(2470)) or (layer6_outputs(1970)));
    outputs(1855) <= not((layer6_outputs(601)) xor (layer6_outputs(1274)));
    outputs(1856) <= (layer6_outputs(1906)) xor (layer6_outputs(2113));
    outputs(1857) <= (layer6_outputs(837)) or (layer6_outputs(2318));
    outputs(1858) <= not(layer6_outputs(2128));
    outputs(1859) <= layer6_outputs(2189);
    outputs(1860) <= not(layer6_outputs(258));
    outputs(1861) <= not(layer6_outputs(1936));
    outputs(1862) <= not(layer6_outputs(1058));
    outputs(1863) <= (layer6_outputs(1122)) and (layer6_outputs(1263));
    outputs(1864) <= layer6_outputs(1156);
    outputs(1865) <= layer6_outputs(97);
    outputs(1866) <= (layer6_outputs(2019)) or (layer6_outputs(673));
    outputs(1867) <= not((layer6_outputs(1271)) xor (layer6_outputs(675)));
    outputs(1868) <= not((layer6_outputs(993)) or (layer6_outputs(535)));
    outputs(1869) <= (layer6_outputs(1325)) xor (layer6_outputs(1237));
    outputs(1870) <= not((layer6_outputs(328)) or (layer6_outputs(2528)));
    outputs(1871) <= not(layer6_outputs(1993));
    outputs(1872) <= not(layer6_outputs(17));
    outputs(1873) <= (layer6_outputs(1825)) xor (layer6_outputs(432));
    outputs(1874) <= (layer6_outputs(1122)) and not (layer6_outputs(805));
    outputs(1875) <= (layer6_outputs(1611)) xor (layer6_outputs(2140));
    outputs(1876) <= (layer6_outputs(1130)) and (layer6_outputs(1712));
    outputs(1877) <= not(layer6_outputs(1179)) or (layer6_outputs(2499));
    outputs(1878) <= layer6_outputs(883);
    outputs(1879) <= layer6_outputs(1555);
    outputs(1880) <= not(layer6_outputs(2479));
    outputs(1881) <= (layer6_outputs(601)) and not (layer6_outputs(1314));
    outputs(1882) <= layer6_outputs(81);
    outputs(1883) <= not(layer6_outputs(355));
    outputs(1884) <= layer6_outputs(1819);
    outputs(1885) <= not((layer6_outputs(1983)) or (layer6_outputs(548)));
    outputs(1886) <= not(layer6_outputs(1784));
    outputs(1887) <= not(layer6_outputs(1326));
    outputs(1888) <= layer6_outputs(506);
    outputs(1889) <= not(layer6_outputs(2100));
    outputs(1890) <= (layer6_outputs(2556)) and not (layer6_outputs(440));
    outputs(1891) <= layer6_outputs(1028);
    outputs(1892) <= layer6_outputs(494);
    outputs(1893) <= not((layer6_outputs(513)) xor (layer6_outputs(1933)));
    outputs(1894) <= not((layer6_outputs(1233)) or (layer6_outputs(1678)));
    outputs(1895) <= not(layer6_outputs(2362));
    outputs(1896) <= layer6_outputs(427);
    outputs(1897) <= not((layer6_outputs(1909)) xor (layer6_outputs(2361)));
    outputs(1898) <= (layer6_outputs(1804)) xor (layer6_outputs(1097));
    outputs(1899) <= not((layer6_outputs(878)) or (layer6_outputs(260)));
    outputs(1900) <= layer6_outputs(1710);
    outputs(1901) <= layer6_outputs(1066);
    outputs(1902) <= (layer6_outputs(2306)) and not (layer6_outputs(2460));
    outputs(1903) <= layer6_outputs(1699);
    outputs(1904) <= (layer6_outputs(2258)) xor (layer6_outputs(2372));
    outputs(1905) <= not(layer6_outputs(25));
    outputs(1906) <= not(layer6_outputs(797));
    outputs(1907) <= not((layer6_outputs(442)) xor (layer6_outputs(1283)));
    outputs(1908) <= not(layer6_outputs(230));
    outputs(1909) <= not(layer6_outputs(323)) or (layer6_outputs(2437));
    outputs(1910) <= not(layer6_outputs(1520));
    outputs(1911) <= not((layer6_outputs(1940)) xor (layer6_outputs(2082)));
    outputs(1912) <= layer6_outputs(1629);
    outputs(1913) <= layer6_outputs(2131);
    outputs(1914) <= (layer6_outputs(2141)) and (layer6_outputs(1548));
    outputs(1915) <= layer6_outputs(1361);
    outputs(1916) <= (layer6_outputs(2252)) xor (layer6_outputs(308));
    outputs(1917) <= not(layer6_outputs(1181)) or (layer6_outputs(110));
    outputs(1918) <= not(layer6_outputs(2277));
    outputs(1919) <= layer6_outputs(40);
    outputs(1920) <= (layer6_outputs(1247)) and not (layer6_outputs(316));
    outputs(1921) <= not(layer6_outputs(344));
    outputs(1922) <= (layer6_outputs(562)) xor (layer6_outputs(1034));
    outputs(1923) <= not(layer6_outputs(1149));
    outputs(1924) <= layer6_outputs(2130);
    outputs(1925) <= layer6_outputs(2299);
    outputs(1926) <= not(layer6_outputs(1391));
    outputs(1927) <= layer6_outputs(2326);
    outputs(1928) <= not((layer6_outputs(2266)) or (layer6_outputs(2412)));
    outputs(1929) <= not((layer6_outputs(2289)) or (layer6_outputs(94)));
    outputs(1930) <= (layer6_outputs(299)) xor (layer6_outputs(1875));
    outputs(1931) <= layer6_outputs(676);
    outputs(1932) <= layer6_outputs(1758);
    outputs(1933) <= layer6_outputs(1919);
    outputs(1934) <= not(layer6_outputs(2394));
    outputs(1935) <= not(layer6_outputs(1815)) or (layer6_outputs(742));
    outputs(1936) <= not((layer6_outputs(1205)) or (layer6_outputs(237)));
    outputs(1937) <= (layer6_outputs(14)) and not (layer6_outputs(1321));
    outputs(1938) <= (layer6_outputs(269)) and not (layer6_outputs(1232));
    outputs(1939) <= layer6_outputs(57);
    outputs(1940) <= layer6_outputs(1505);
    outputs(1941) <= not((layer6_outputs(688)) or (layer6_outputs(392)));
    outputs(1942) <= not(layer6_outputs(34));
    outputs(1943) <= (layer6_outputs(2138)) and not (layer6_outputs(2128));
    outputs(1944) <= not(layer6_outputs(18));
    outputs(1945) <= not(layer6_outputs(2056));
    outputs(1946) <= (layer6_outputs(1156)) and (layer6_outputs(1468));
    outputs(1947) <= (layer6_outputs(669)) and (layer6_outputs(2369));
    outputs(1948) <= (layer6_outputs(1716)) and (layer6_outputs(1734));
    outputs(1949) <= (layer6_outputs(1448)) xor (layer6_outputs(1908));
    outputs(1950) <= not((layer6_outputs(2349)) xor (layer6_outputs(2145)));
    outputs(1951) <= layer6_outputs(2214);
    outputs(1952) <= not((layer6_outputs(2546)) xor (layer6_outputs(2336)));
    outputs(1953) <= not(layer6_outputs(254));
    outputs(1954) <= not(layer6_outputs(1442));
    outputs(1955) <= (layer6_outputs(1886)) and not (layer6_outputs(1463));
    outputs(1956) <= (layer6_outputs(2084)) and not (layer6_outputs(2034));
    outputs(1957) <= not((layer6_outputs(704)) xor (layer6_outputs(493)));
    outputs(1958) <= not((layer6_outputs(644)) or (layer6_outputs(296)));
    outputs(1959) <= (layer6_outputs(2367)) xor (layer6_outputs(1760));
    outputs(1960) <= not(layer6_outputs(874));
    outputs(1961) <= not((layer6_outputs(2557)) or (layer6_outputs(274)));
    outputs(1962) <= not((layer6_outputs(2438)) xor (layer6_outputs(2199)));
    outputs(1963) <= not((layer6_outputs(80)) xor (layer6_outputs(2281)));
    outputs(1964) <= (layer6_outputs(2315)) and not (layer6_outputs(89));
    outputs(1965) <= layer6_outputs(2068);
    outputs(1966) <= not(layer6_outputs(2045));
    outputs(1967) <= layer6_outputs(2265);
    outputs(1968) <= (layer6_outputs(96)) xor (layer6_outputs(1210));
    outputs(1969) <= layer6_outputs(1543);
    outputs(1970) <= not((layer6_outputs(2038)) or (layer6_outputs(1590)));
    outputs(1971) <= layer6_outputs(908);
    outputs(1972) <= not(layer6_outputs(409));
    outputs(1973) <= (layer6_outputs(2434)) and (layer6_outputs(2327));
    outputs(1974) <= (layer6_outputs(2112)) and (layer6_outputs(1513));
    outputs(1975) <= (layer6_outputs(1296)) and not (layer6_outputs(2428));
    outputs(1976) <= not(layer6_outputs(963)) or (layer6_outputs(2261));
    outputs(1977) <= layer6_outputs(2037);
    outputs(1978) <= (layer6_outputs(2178)) and (layer6_outputs(2551));
    outputs(1979) <= layer6_outputs(1493);
    outputs(1980) <= not(layer6_outputs(680));
    outputs(1981) <= not((layer6_outputs(1086)) xor (layer6_outputs(1857)));
    outputs(1982) <= layer6_outputs(1727);
    outputs(1983) <= layer6_outputs(1216);
    outputs(1984) <= layer6_outputs(524);
    outputs(1985) <= not((layer6_outputs(622)) xor (layer6_outputs(1763)));
    outputs(1986) <= not(layer6_outputs(1485));
    outputs(1987) <= not(layer6_outputs(1478)) or (layer6_outputs(825));
    outputs(1988) <= not((layer6_outputs(607)) xor (layer6_outputs(498)));
    outputs(1989) <= layer6_outputs(937);
    outputs(1990) <= layer6_outputs(836);
    outputs(1991) <= not((layer6_outputs(747)) and (layer6_outputs(278)));
    outputs(1992) <= not((layer6_outputs(338)) or (layer6_outputs(1025)));
    outputs(1993) <= (layer6_outputs(2352)) xor (layer6_outputs(1132));
    outputs(1994) <= layer6_outputs(2241);
    outputs(1995) <= (layer6_outputs(353)) and (layer6_outputs(1943));
    outputs(1996) <= not(layer6_outputs(714));
    outputs(1997) <= not(layer6_outputs(609));
    outputs(1998) <= not(layer6_outputs(2409));
    outputs(1999) <= (layer6_outputs(2535)) and (layer6_outputs(2297));
    outputs(2000) <= (layer6_outputs(865)) xor (layer6_outputs(2405));
    outputs(2001) <= layer6_outputs(1151);
    outputs(2002) <= layer6_outputs(2031);
    outputs(2003) <= layer6_outputs(1656);
    outputs(2004) <= layer6_outputs(1907);
    outputs(2005) <= layer6_outputs(1694);
    outputs(2006) <= layer6_outputs(76);
    outputs(2007) <= not(layer6_outputs(1201));
    outputs(2008) <= not((layer6_outputs(2388)) or (layer6_outputs(1973)));
    outputs(2009) <= (layer6_outputs(1368)) and not (layer6_outputs(2076));
    outputs(2010) <= (layer6_outputs(1659)) xor (layer6_outputs(709));
    outputs(2011) <= layer6_outputs(1416);
    outputs(2012) <= not(layer6_outputs(2007));
    outputs(2013) <= not((layer6_outputs(2498)) or (layer6_outputs(1256)));
    outputs(2014) <= not(layer6_outputs(665)) or (layer6_outputs(370));
    outputs(2015) <= layer6_outputs(2488);
    outputs(2016) <= (layer6_outputs(2413)) and not (layer6_outputs(1024));
    outputs(2017) <= layer6_outputs(434);
    outputs(2018) <= not((layer6_outputs(11)) xor (layer6_outputs(1743)));
    outputs(2019) <= layer6_outputs(2535);
    outputs(2020) <= not(layer6_outputs(726));
    outputs(2021) <= (layer6_outputs(1052)) and not (layer6_outputs(2291));
    outputs(2022) <= not((layer6_outputs(2108)) xor (layer6_outputs(138)));
    outputs(2023) <= layer6_outputs(1998);
    outputs(2024) <= (layer6_outputs(1036)) xor (layer6_outputs(2440));
    outputs(2025) <= (layer6_outputs(2471)) and (layer6_outputs(1732));
    outputs(2026) <= (layer6_outputs(1792)) and not (layer6_outputs(1070));
    outputs(2027) <= not(layer6_outputs(1997));
    outputs(2028) <= not(layer6_outputs(1288)) or (layer6_outputs(1717));
    outputs(2029) <= layer6_outputs(651);
    outputs(2030) <= (layer6_outputs(2117)) and not (layer6_outputs(459));
    outputs(2031) <= layer6_outputs(2242);
    outputs(2032) <= not(layer6_outputs(2555));
    outputs(2033) <= not((layer6_outputs(282)) or (layer6_outputs(1903)));
    outputs(2034) <= (layer6_outputs(26)) and not (layer6_outputs(1936));
    outputs(2035) <= (layer6_outputs(1817)) and (layer6_outputs(1821));
    outputs(2036) <= not(layer6_outputs(547));
    outputs(2037) <= not((layer6_outputs(1450)) or (layer6_outputs(454)));
    outputs(2038) <= (layer6_outputs(1872)) xor (layer6_outputs(2513));
    outputs(2039) <= not(layer6_outputs(1262));
    outputs(2040) <= not((layer6_outputs(1313)) xor (layer6_outputs(2102)));
    outputs(2041) <= layer6_outputs(352);
    outputs(2042) <= (layer6_outputs(1307)) and not (layer6_outputs(767));
    outputs(2043) <= not((layer6_outputs(535)) or (layer6_outputs(1521)));
    outputs(2044) <= layer6_outputs(231);
    outputs(2045) <= not(layer6_outputs(2050)) or (layer6_outputs(1887));
    outputs(2046) <= (layer6_outputs(2396)) and (layer6_outputs(1075));
    outputs(2047) <= (layer6_outputs(1661)) and (layer6_outputs(31));
    outputs(2048) <= layer6_outputs(41);
    outputs(2049) <= layer6_outputs(270);
    outputs(2050) <= not(layer6_outputs(1792));
    outputs(2051) <= not((layer6_outputs(917)) or (layer6_outputs(1586)));
    outputs(2052) <= (layer6_outputs(945)) xor (layer6_outputs(1245));
    outputs(2053) <= (layer6_outputs(1270)) xor (layer6_outputs(478));
    outputs(2054) <= not((layer6_outputs(410)) xor (layer6_outputs(920)));
    outputs(2055) <= layer6_outputs(1001);
    outputs(2056) <= not((layer6_outputs(1770)) xor (layer6_outputs(2109)));
    outputs(2057) <= not(layer6_outputs(988));
    outputs(2058) <= layer6_outputs(528);
    outputs(2059) <= not((layer6_outputs(778)) xor (layer6_outputs(2163)));
    outputs(2060) <= layer6_outputs(1527);
    outputs(2061) <= not((layer6_outputs(932)) or (layer6_outputs(1890)));
    outputs(2062) <= not(layer6_outputs(71));
    outputs(2063) <= not((layer6_outputs(49)) or (layer6_outputs(1860)));
    outputs(2064) <= (layer6_outputs(1169)) and not (layer6_outputs(427));
    outputs(2065) <= not((layer6_outputs(798)) xor (layer6_outputs(2443)));
    outputs(2066) <= not(layer6_outputs(604));
    outputs(2067) <= not(layer6_outputs(1313));
    outputs(2068) <= (layer6_outputs(2230)) xor (layer6_outputs(1444));
    outputs(2069) <= layer6_outputs(281);
    outputs(2070) <= layer6_outputs(2467);
    outputs(2071) <= layer6_outputs(1624);
    outputs(2072) <= (layer6_outputs(1206)) xor (layer6_outputs(226));
    outputs(2073) <= layer6_outputs(710);
    outputs(2074) <= not(layer6_outputs(2012));
    outputs(2075) <= layer6_outputs(231);
    outputs(2076) <= not(layer6_outputs(277));
    outputs(2077) <= layer6_outputs(733);
    outputs(2078) <= not((layer6_outputs(205)) xor (layer6_outputs(894)));
    outputs(2079) <= not(layer6_outputs(1581));
    outputs(2080) <= layer6_outputs(2287);
    outputs(2081) <= not(layer6_outputs(1613)) or (layer6_outputs(2518));
    outputs(2082) <= layer6_outputs(1597);
    outputs(2083) <= not(layer6_outputs(2366));
    outputs(2084) <= (layer6_outputs(84)) and not (layer6_outputs(2279));
    outputs(2085) <= not(layer6_outputs(1064));
    outputs(2086) <= layer6_outputs(2521);
    outputs(2087) <= not((layer6_outputs(1356)) xor (layer6_outputs(1751)));
    outputs(2088) <= not(layer6_outputs(855)) or (layer6_outputs(967));
    outputs(2089) <= not(layer6_outputs(405));
    outputs(2090) <= layer6_outputs(188);
    outputs(2091) <= (layer6_outputs(1217)) and not (layer6_outputs(1068));
    outputs(2092) <= not((layer6_outputs(1)) xor (layer6_outputs(287)));
    outputs(2093) <= (layer6_outputs(130)) and not (layer6_outputs(108));
    outputs(2094) <= layer6_outputs(2510);
    outputs(2095) <= layer6_outputs(1153);
    outputs(2096) <= not(layer6_outputs(233));
    outputs(2097) <= not((layer6_outputs(1573)) and (layer6_outputs(2195)));
    outputs(2098) <= not(layer6_outputs(2225));
    outputs(2099) <= layer6_outputs(213);
    outputs(2100) <= layer6_outputs(983);
    outputs(2101) <= layer6_outputs(432);
    outputs(2102) <= not(layer6_outputs(2364));
    outputs(2103) <= (layer6_outputs(1187)) xor (layer6_outputs(1959));
    outputs(2104) <= not(layer6_outputs(1946));
    outputs(2105) <= not((layer6_outputs(139)) or (layer6_outputs(2150)));
    outputs(2106) <= layer6_outputs(1038);
    outputs(2107) <= layer6_outputs(1471);
    outputs(2108) <= (layer6_outputs(595)) xor (layer6_outputs(305));
    outputs(2109) <= not(layer6_outputs(1144));
    outputs(2110) <= not(layer6_outputs(763));
    outputs(2111) <= layer6_outputs(1923);
    outputs(2112) <= not(layer6_outputs(347)) or (layer6_outputs(218));
    outputs(2113) <= layer6_outputs(1618);
    outputs(2114) <= layer6_outputs(1466);
    outputs(2115) <= not(layer6_outputs(2508));
    outputs(2116) <= not(layer6_outputs(244));
    outputs(2117) <= not((layer6_outputs(1207)) xor (layer6_outputs(1965)));
    outputs(2118) <= layer6_outputs(1770);
    outputs(2119) <= not(layer6_outputs(1192));
    outputs(2120) <= not((layer6_outputs(43)) xor (layer6_outputs(349)));
    outputs(2121) <= layer6_outputs(1813);
    outputs(2122) <= not(layer6_outputs(302));
    outputs(2123) <= (layer6_outputs(431)) or (layer6_outputs(767));
    outputs(2124) <= (layer6_outputs(715)) and not (layer6_outputs(1406));
    outputs(2125) <= not(layer6_outputs(243));
    outputs(2126) <= layer6_outputs(1985);
    outputs(2127) <= layer6_outputs(1562);
    outputs(2128) <= (layer6_outputs(1491)) xor (layer6_outputs(1816));
    outputs(2129) <= not(layer6_outputs(933));
    outputs(2130) <= layer6_outputs(84);
    outputs(2131) <= not((layer6_outputs(1700)) or (layer6_outputs(2150)));
    outputs(2132) <= layer6_outputs(529);
    outputs(2133) <= layer6_outputs(1317);
    outputs(2134) <= not((layer6_outputs(1606)) or (layer6_outputs(2194)));
    outputs(2135) <= not(layer6_outputs(1148));
    outputs(2136) <= not(layer6_outputs(1579));
    outputs(2137) <= (layer6_outputs(1037)) and not (layer6_outputs(92));
    outputs(2138) <= not((layer6_outputs(400)) or (layer6_outputs(1974)));
    outputs(2139) <= not(layer6_outputs(363));
    outputs(2140) <= not(layer6_outputs(2098));
    outputs(2141) <= not(layer6_outputs(1822));
    outputs(2142) <= layer6_outputs(256);
    outputs(2143) <= layer6_outputs(2533);
    outputs(2144) <= not((layer6_outputs(1453)) xor (layer6_outputs(4)));
    outputs(2145) <= not(layer6_outputs(1745));
    outputs(2146) <= (layer6_outputs(418)) and not (layer6_outputs(2080));
    outputs(2147) <= not(layer6_outputs(934));
    outputs(2148) <= layer6_outputs(1985);
    outputs(2149) <= not((layer6_outputs(327)) xor (layer6_outputs(551)));
    outputs(2150) <= (layer6_outputs(721)) or (layer6_outputs(178));
    outputs(2151) <= layer6_outputs(1475);
    outputs(2152) <= (layer6_outputs(1086)) xor (layer6_outputs(658));
    outputs(2153) <= not(layer6_outputs(1986));
    outputs(2154) <= not((layer6_outputs(379)) xor (layer6_outputs(761)));
    outputs(2155) <= (layer6_outputs(400)) xor (layer6_outputs(55));
    outputs(2156) <= layer6_outputs(944);
    outputs(2157) <= layer6_outputs(2143);
    outputs(2158) <= not((layer6_outputs(757)) xor (layer6_outputs(468)));
    outputs(2159) <= not(layer6_outputs(366));
    outputs(2160) <= not(layer6_outputs(1285));
    outputs(2161) <= (layer6_outputs(297)) and not (layer6_outputs(450));
    outputs(2162) <= not((layer6_outputs(361)) or (layer6_outputs(2516)));
    outputs(2163) <= not(layer6_outputs(2509));
    outputs(2164) <= not(layer6_outputs(469)) or (layer6_outputs(549));
    outputs(2165) <= not(layer6_outputs(2290));
    outputs(2166) <= not((layer6_outputs(1999)) xor (layer6_outputs(1463)));
    outputs(2167) <= layer6_outputs(1585);
    outputs(2168) <= (layer6_outputs(2296)) and not (layer6_outputs(2316));
    outputs(2169) <= layer6_outputs(572);
    outputs(2170) <= layer6_outputs(1988);
    outputs(2171) <= not(layer6_outputs(1150));
    outputs(2172) <= layer6_outputs(68);
    outputs(2173) <= layer6_outputs(284);
    outputs(2174) <= not(layer6_outputs(2216));
    outputs(2175) <= (layer6_outputs(2205)) and not (layer6_outputs(810));
    outputs(2176) <= (layer6_outputs(1013)) xor (layer6_outputs(1402));
    outputs(2177) <= not((layer6_outputs(2333)) xor (layer6_outputs(205)));
    outputs(2178) <= layer6_outputs(1774);
    outputs(2179) <= not((layer6_outputs(1932)) and (layer6_outputs(1333)));
    outputs(2180) <= (layer6_outputs(719)) and not (layer6_outputs(219));
    outputs(2181) <= not(layer6_outputs(1070));
    outputs(2182) <= not((layer6_outputs(739)) xor (layer6_outputs(957)));
    outputs(2183) <= not(layer6_outputs(2516));
    outputs(2184) <= layer6_outputs(1236);
    outputs(2185) <= layer6_outputs(1485);
    outputs(2186) <= layer6_outputs(1211);
    outputs(2187) <= not(layer6_outputs(475));
    outputs(2188) <= (layer6_outputs(87)) and not (layer6_outputs(951));
    outputs(2189) <= (layer6_outputs(2390)) xor (layer6_outputs(2358));
    outputs(2190) <= not(layer6_outputs(833));
    outputs(2191) <= layer6_outputs(943);
    outputs(2192) <= layer6_outputs(2384);
    outputs(2193) <= layer6_outputs(1128);
    outputs(2194) <= not(layer6_outputs(288)) or (layer6_outputs(996));
    outputs(2195) <= not(layer6_outputs(847));
    outputs(2196) <= layer6_outputs(332);
    outputs(2197) <= (layer6_outputs(1149)) and not (layer6_outputs(855));
    outputs(2198) <= not((layer6_outputs(841)) xor (layer6_outputs(549)));
    outputs(2199) <= not(layer6_outputs(1637));
    outputs(2200) <= (layer6_outputs(495)) and not (layer6_outputs(929));
    outputs(2201) <= not(layer6_outputs(1043));
    outputs(2202) <= not(layer6_outputs(2101));
    outputs(2203) <= (layer6_outputs(2193)) or (layer6_outputs(589));
    outputs(2204) <= not(layer6_outputs(2493)) or (layer6_outputs(2313));
    outputs(2205) <= (layer6_outputs(1883)) xor (layer6_outputs(1839));
    outputs(2206) <= layer6_outputs(2152);
    outputs(2207) <= layer6_outputs(2289);
    outputs(2208) <= layer6_outputs(1459);
    outputs(2209) <= (layer6_outputs(1720)) xor (layer6_outputs(1697));
    outputs(2210) <= layer6_outputs(2478);
    outputs(2211) <= layer6_outputs(1800);
    outputs(2212) <= not(layer6_outputs(834));
    outputs(2213) <= not(layer6_outputs(512));
    outputs(2214) <= (layer6_outputs(150)) and not (layer6_outputs(1008));
    outputs(2215) <= not(layer6_outputs(1975));
    outputs(2216) <= not(layer6_outputs(615));
    outputs(2217) <= not(layer6_outputs(112));
    outputs(2218) <= layer6_outputs(2380);
    outputs(2219) <= not(layer6_outputs(743));
    outputs(2220) <= not((layer6_outputs(1275)) xor (layer6_outputs(2033)));
    outputs(2221) <= layer6_outputs(2380);
    outputs(2222) <= (layer6_outputs(1976)) and not (layer6_outputs(2039));
    outputs(2223) <= layer6_outputs(1217);
    outputs(2224) <= layer6_outputs(429);
    outputs(2225) <= layer6_outputs(1821);
    outputs(2226) <= not(layer6_outputs(413));
    outputs(2227) <= (layer6_outputs(1421)) xor (layer6_outputs(430));
    outputs(2228) <= not((layer6_outputs(1401)) xor (layer6_outputs(747)));
    outputs(2229) <= not(layer6_outputs(1417));
    outputs(2230) <= not(layer6_outputs(2210));
    outputs(2231) <= not(layer6_outputs(2288));
    outputs(2232) <= not((layer6_outputs(271)) xor (layer6_outputs(2473)));
    outputs(2233) <= not(layer6_outputs(1978));
    outputs(2234) <= (layer6_outputs(722)) and not (layer6_outputs(744));
    outputs(2235) <= (layer6_outputs(1660)) xor (layer6_outputs(760));
    outputs(2236) <= not((layer6_outputs(217)) xor (layer6_outputs(1019)));
    outputs(2237) <= not(layer6_outputs(2415));
    outputs(2238) <= layer6_outputs(2521);
    outputs(2239) <= not(layer6_outputs(1645));
    outputs(2240) <= (layer6_outputs(1351)) xor (layer6_outputs(1845));
    outputs(2241) <= (layer6_outputs(685)) and not (layer6_outputs(991));
    outputs(2242) <= layer6_outputs(1919);
    outputs(2243) <= layer6_outputs(1805);
    outputs(2244) <= not((layer6_outputs(269)) and (layer6_outputs(2503)));
    outputs(2245) <= not(layer6_outputs(1811));
    outputs(2246) <= not((layer6_outputs(865)) xor (layer6_outputs(444)));
    outputs(2247) <= (layer6_outputs(1746)) and not (layer6_outputs(1161));
    outputs(2248) <= (layer6_outputs(284)) and not (layer6_outputs(1902));
    outputs(2249) <= not(layer6_outputs(1289));
    outputs(2250) <= layer6_outputs(944);
    outputs(2251) <= layer6_outputs(642);
    outputs(2252) <= not(layer6_outputs(2541));
    outputs(2253) <= layer6_outputs(1931);
    outputs(2254) <= not(layer6_outputs(1489));
    outputs(2255) <= (layer6_outputs(800)) and not (layer6_outputs(330));
    outputs(2256) <= not(layer6_outputs(2084));
    outputs(2257) <= layer6_outputs(1420);
    outputs(2258) <= layer6_outputs(1206);
    outputs(2259) <= (layer6_outputs(1612)) xor (layer6_outputs(325));
    outputs(2260) <= layer6_outputs(1335);
    outputs(2261) <= not(layer6_outputs(2198)) or (layer6_outputs(2360));
    outputs(2262) <= not((layer6_outputs(2263)) xor (layer6_outputs(1163)));
    outputs(2263) <= not((layer6_outputs(394)) xor (layer6_outputs(1350)));
    outputs(2264) <= layer6_outputs(1722);
    outputs(2265) <= not(layer6_outputs(71));
    outputs(2266) <= (layer6_outputs(2001)) and not (layer6_outputs(1014));
    outputs(2267) <= not(layer6_outputs(612));
    outputs(2268) <= layer6_outputs(852);
    outputs(2269) <= not(layer6_outputs(1116));
    outputs(2270) <= layer6_outputs(1229);
    outputs(2271) <= layer6_outputs(246);
    outputs(2272) <= layer6_outputs(1633);
    outputs(2273) <= (layer6_outputs(83)) and (layer6_outputs(1891));
    outputs(2274) <= not((layer6_outputs(2121)) xor (layer6_outputs(557)));
    outputs(2275) <= layer6_outputs(2113);
    outputs(2276) <= layer6_outputs(900);
    outputs(2277) <= (layer6_outputs(1785)) and not (layer6_outputs(314));
    outputs(2278) <= not(layer6_outputs(2362));
    outputs(2279) <= layer6_outputs(1190);
    outputs(2280) <= (layer6_outputs(2184)) and (layer6_outputs(716));
    outputs(2281) <= layer6_outputs(936);
    outputs(2282) <= (layer6_outputs(224)) xor (layer6_outputs(359));
    outputs(2283) <= (layer6_outputs(1872)) and (layer6_outputs(670));
    outputs(2284) <= not(layer6_outputs(1440));
    outputs(2285) <= not(layer6_outputs(2052));
    outputs(2286) <= not(layer6_outputs(1074));
    outputs(2287) <= not(layer6_outputs(1565));
    outputs(2288) <= not(layer6_outputs(2411));
    outputs(2289) <= layer6_outputs(1532);
    outputs(2290) <= (layer6_outputs(455)) xor (layer6_outputs(1335));
    outputs(2291) <= layer6_outputs(960);
    outputs(2292) <= layer6_outputs(1441);
    outputs(2293) <= not(layer6_outputs(558));
    outputs(2294) <= layer6_outputs(1807);
    outputs(2295) <= (layer6_outputs(238)) and not (layer6_outputs(2093));
    outputs(2296) <= not(layer6_outputs(243));
    outputs(2297) <= (layer6_outputs(1123)) xor (layer6_outputs(776));
    outputs(2298) <= not(layer6_outputs(2298));
    outputs(2299) <= (layer6_outputs(1276)) xor (layer6_outputs(2036));
    outputs(2300) <= not(layer6_outputs(1925));
    outputs(2301) <= layer6_outputs(681);
    outputs(2302) <= not(layer6_outputs(1197));
    outputs(2303) <= not(layer6_outputs(553));
    outputs(2304) <= (layer6_outputs(2328)) xor (layer6_outputs(1062));
    outputs(2305) <= not((layer6_outputs(2393)) and (layer6_outputs(1111)));
    outputs(2306) <= layer6_outputs(673);
    outputs(2307) <= (layer6_outputs(813)) and not (layer6_outputs(560));
    outputs(2308) <= layer6_outputs(1081);
    outputs(2309) <= not((layer6_outputs(131)) xor (layer6_outputs(2212)));
    outputs(2310) <= layer6_outputs(837);
    outputs(2311) <= not((layer6_outputs(1642)) xor (layer6_outputs(1448)));
    outputs(2312) <= not((layer6_outputs(882)) or (layer6_outputs(509)));
    outputs(2313) <= not((layer6_outputs(1762)) xor (layer6_outputs(498)));
    outputs(2314) <= not(layer6_outputs(711));
    outputs(2315) <= (layer6_outputs(2108)) xor (layer6_outputs(1517));
    outputs(2316) <= (layer6_outputs(1863)) xor (layer6_outputs(1421));
    outputs(2317) <= layer6_outputs(1118);
    outputs(2318) <= layer6_outputs(982);
    outputs(2319) <= not((layer6_outputs(64)) or (layer6_outputs(402)));
    outputs(2320) <= not((layer6_outputs(2342)) xor (layer6_outputs(1569)));
    outputs(2321) <= layer6_outputs(2198);
    outputs(2322) <= layer6_outputs(1724);
    outputs(2323) <= not(layer6_outputs(1839));
    outputs(2324) <= layer6_outputs(56);
    outputs(2325) <= (layer6_outputs(774)) and not (layer6_outputs(559));
    outputs(2326) <= layer6_outputs(1066);
    outputs(2327) <= layer6_outputs(999);
    outputs(2328) <= not(layer6_outputs(2296));
    outputs(2329) <= not(layer6_outputs(1020));
    outputs(2330) <= (layer6_outputs(2330)) xor (layer6_outputs(306));
    outputs(2331) <= layer6_outputs(8);
    outputs(2332) <= (layer6_outputs(1852)) and not (layer6_outputs(1418));
    outputs(2333) <= (layer6_outputs(2273)) xor (layer6_outputs(230));
    outputs(2334) <= (layer6_outputs(781)) or (layer6_outputs(98));
    outputs(2335) <= (layer6_outputs(726)) and (layer6_outputs(1361));
    outputs(2336) <= not(layer6_outputs(212));
    outputs(2337) <= not((layer6_outputs(1165)) xor (layer6_outputs(801)));
    outputs(2338) <= not(layer6_outputs(2181));
    outputs(2339) <= layer6_outputs(1009);
    outputs(2340) <= not(layer6_outputs(1587));
    outputs(2341) <= layer6_outputs(1843);
    outputs(2342) <= layer6_outputs(1826);
    outputs(2343) <= not(layer6_outputs(294));
    outputs(2344) <= (layer6_outputs(1427)) and not (layer6_outputs(2402));
    outputs(2345) <= not((layer6_outputs(661)) xor (layer6_outputs(2405)));
    outputs(2346) <= not(layer6_outputs(341));
    outputs(2347) <= layer6_outputs(214);
    outputs(2348) <= not(layer6_outputs(734));
    outputs(2349) <= layer6_outputs(29);
    outputs(2350) <= not(layer6_outputs(1337));
    outputs(2351) <= (layer6_outputs(1432)) and not (layer6_outputs(530));
    outputs(2352) <= not((layer6_outputs(1159)) xor (layer6_outputs(2321)));
    outputs(2353) <= not(layer6_outputs(822));
    outputs(2354) <= not(layer6_outputs(270));
    outputs(2355) <= not(layer6_outputs(2010));
    outputs(2356) <= not(layer6_outputs(1172));
    outputs(2357) <= layer6_outputs(1734);
    outputs(2358) <= (layer6_outputs(949)) and not (layer6_outputs(1585));
    outputs(2359) <= not(layer6_outputs(1371));
    outputs(2360) <= (layer6_outputs(351)) and not (layer6_outputs(116));
    outputs(2361) <= not(layer6_outputs(363));
    outputs(2362) <= (layer6_outputs(193)) and (layer6_outputs(1615));
    outputs(2363) <= not((layer6_outputs(802)) or (layer6_outputs(93)));
    outputs(2364) <= layer6_outputs(737);
    outputs(2365) <= layer6_outputs(1085);
    outputs(2366) <= not(layer6_outputs(985));
    outputs(2367) <= layer6_outputs(669);
    outputs(2368) <= not((layer6_outputs(1017)) xor (layer6_outputs(660)));
    outputs(2369) <= layer6_outputs(461);
    outputs(2370) <= not(layer6_outputs(128));
    outputs(2371) <= not((layer6_outputs(1008)) or (layer6_outputs(612)));
    outputs(2372) <= not(layer6_outputs(2416));
    outputs(2373) <= not(layer6_outputs(356));
    outputs(2374) <= layer6_outputs(1834);
    outputs(2375) <= (layer6_outputs(1160)) xor (layer6_outputs(361));
    outputs(2376) <= layer6_outputs(1800);
    outputs(2377) <= not(layer6_outputs(144));
    outputs(2378) <= not(layer6_outputs(1605));
    outputs(2379) <= layer6_outputs(1698);
    outputs(2380) <= not(layer6_outputs(1781));
    outputs(2381) <= layer6_outputs(161);
    outputs(2382) <= not(layer6_outputs(775));
    outputs(2383) <= not((layer6_outputs(1682)) or (layer6_outputs(974)));
    outputs(2384) <= not(layer6_outputs(1316));
    outputs(2385) <= not(layer6_outputs(2412));
    outputs(2386) <= layer6_outputs(1137);
    outputs(2387) <= (layer6_outputs(2379)) and not (layer6_outputs(1133));
    outputs(2388) <= (layer6_outputs(2253)) and not (layer6_outputs(1393));
    outputs(2389) <= (layer6_outputs(1174)) or (layer6_outputs(1830));
    outputs(2390) <= layer6_outputs(343);
    outputs(2391) <= not((layer6_outputs(318)) or (layer6_outputs(411)));
    outputs(2392) <= (layer6_outputs(542)) and (layer6_outputs(56));
    outputs(2393) <= layer6_outputs(1631);
    outputs(2394) <= not(layer6_outputs(714));
    outputs(2395) <= not(layer6_outputs(287));
    outputs(2396) <= not(layer6_outputs(356));
    outputs(2397) <= (layer6_outputs(1416)) and (layer6_outputs(2005));
    outputs(2398) <= (layer6_outputs(373)) and (layer6_outputs(1565));
    outputs(2399) <= not(layer6_outputs(1405));
    outputs(2400) <= layer6_outputs(1598);
    outputs(2401) <= not((layer6_outputs(1236)) or (layer6_outputs(974)));
    outputs(2402) <= not((layer6_outputs(1672)) xor (layer6_outputs(1477)));
    outputs(2403) <= not(layer6_outputs(2239));
    outputs(2404) <= (layer6_outputs(2211)) xor (layer6_outputs(2273));
    outputs(2405) <= not(layer6_outputs(1049)) or (layer6_outputs(2464));
    outputs(2406) <= layer6_outputs(1909);
    outputs(2407) <= layer6_outputs(2525);
    outputs(2408) <= layer6_outputs(960);
    outputs(2409) <= not(layer6_outputs(2493));
    outputs(2410) <= layer6_outputs(1707);
    outputs(2411) <= not(layer6_outputs(1041));
    outputs(2412) <= not(layer6_outputs(454));
    outputs(2413) <= (layer6_outputs(2223)) or (layer6_outputs(1241));
    outputs(2414) <= layer6_outputs(12);
    outputs(2415) <= layer6_outputs(2415);
    outputs(2416) <= not(layer6_outputs(2158));
    outputs(2417) <= (layer6_outputs(1508)) xor (layer6_outputs(2019));
    outputs(2418) <= (layer6_outputs(718)) xor (layer6_outputs(1951));
    outputs(2419) <= layer6_outputs(1007);
    outputs(2420) <= (layer6_outputs(1823)) and (layer6_outputs(351));
    outputs(2421) <= layer6_outputs(810);
    outputs(2422) <= not((layer6_outputs(2311)) or (layer6_outputs(1691)));
    outputs(2423) <= not(layer6_outputs(1732));
    outputs(2424) <= (layer6_outputs(1408)) and not (layer6_outputs(1833));
    outputs(2425) <= layer6_outputs(1078);
    outputs(2426) <= not((layer6_outputs(1295)) or (layer6_outputs(1238)));
    outputs(2427) <= layer6_outputs(1051);
    outputs(2428) <= not((layer6_outputs(1892)) or (layer6_outputs(1227)));
    outputs(2429) <= layer6_outputs(1530);
    outputs(2430) <= (layer6_outputs(830)) xor (layer6_outputs(2486));
    outputs(2431) <= layer6_outputs(2346);
    outputs(2432) <= not(layer6_outputs(1045));
    outputs(2433) <= not((layer6_outputs(2081)) or (layer6_outputs(1136)));
    outputs(2434) <= (layer6_outputs(1558)) xor (layer6_outputs(247));
    outputs(2435) <= layer6_outputs(970);
    outputs(2436) <= layer6_outputs(2448);
    outputs(2437) <= not(layer6_outputs(403));
    outputs(2438) <= not(layer6_outputs(598));
    outputs(2439) <= (layer6_outputs(779)) or (layer6_outputs(1877));
    outputs(2440) <= layer6_outputs(1928);
    outputs(2441) <= (layer6_outputs(2217)) xor (layer6_outputs(2340));
    outputs(2442) <= layer6_outputs(2205);
    outputs(2443) <= layer6_outputs(1575);
    outputs(2444) <= (layer6_outputs(2237)) and (layer6_outputs(1927));
    outputs(2445) <= not(layer6_outputs(1454));
    outputs(2446) <= not(layer6_outputs(73));
    outputs(2447) <= layer6_outputs(1596);
    outputs(2448) <= (layer6_outputs(769)) xor (layer6_outputs(681));
    outputs(2449) <= (layer6_outputs(755)) and not (layer6_outputs(1951));
    outputs(2450) <= (layer6_outputs(1228)) and not (layer6_outputs(247));
    outputs(2451) <= layer6_outputs(20);
    outputs(2452) <= layer6_outputs(170);
    outputs(2453) <= (layer6_outputs(719)) xor (layer6_outputs(1802));
    outputs(2454) <= not(layer6_outputs(483));
    outputs(2455) <= (layer6_outputs(2271)) and not (layer6_outputs(1996));
    outputs(2456) <= layer6_outputs(336);
    outputs(2457) <= not(layer6_outputs(2450));
    outputs(2458) <= not((layer6_outputs(1511)) or (layer6_outputs(2392)));
    outputs(2459) <= layer6_outputs(793);
    outputs(2460) <= (layer6_outputs(677)) and not (layer6_outputs(1177));
    outputs(2461) <= layer6_outputs(1067);
    outputs(2462) <= layer6_outputs(1336);
    outputs(2463) <= not((layer6_outputs(2049)) or (layer6_outputs(1095)));
    outputs(2464) <= (layer6_outputs(2069)) and not (layer6_outputs(114));
    outputs(2465) <= layer6_outputs(2298);
    outputs(2466) <= not(layer6_outputs(358));
    outputs(2467) <= layer6_outputs(1218);
    outputs(2468) <= not(layer6_outputs(124));
    outputs(2469) <= not(layer6_outputs(1590));
    outputs(2470) <= (layer6_outputs(1687)) xor (layer6_outputs(147));
    outputs(2471) <= not(layer6_outputs(2034));
    outputs(2472) <= not(layer6_outputs(1517));
    outputs(2473) <= not((layer6_outputs(2099)) or (layer6_outputs(1711)));
    outputs(2474) <= not(layer6_outputs(2010));
    outputs(2475) <= not(layer6_outputs(1443));
    outputs(2476) <= layer6_outputs(2173);
    outputs(2477) <= layer6_outputs(1281);
    outputs(2478) <= not(layer6_outputs(577));
    outputs(2479) <= layer6_outputs(983);
    outputs(2480) <= (layer6_outputs(317)) and not (layer6_outputs(1930));
    outputs(2481) <= (layer6_outputs(1608)) xor (layer6_outputs(1630));
    outputs(2482) <= (layer6_outputs(843)) or (layer6_outputs(1761));
    outputs(2483) <= layer6_outputs(1269);
    outputs(2484) <= not(layer6_outputs(1960));
    outputs(2485) <= not((layer6_outputs(2014)) or (layer6_outputs(1623)));
    outputs(2486) <= layer6_outputs(774);
    outputs(2487) <= (layer6_outputs(1998)) and not (layer6_outputs(2038));
    outputs(2488) <= (layer6_outputs(1322)) and not (layer6_outputs(437));
    outputs(2489) <= not(layer6_outputs(1524));
    outputs(2490) <= not((layer6_outputs(792)) xor (layer6_outputs(1808)));
    outputs(2491) <= not(layer6_outputs(1026));
    outputs(2492) <= not((layer6_outputs(559)) and (layer6_outputs(1704)));
    outputs(2493) <= (layer6_outputs(1537)) or (layer6_outputs(1741));
    outputs(2494) <= not(layer6_outputs(2461));
    outputs(2495) <= not((layer6_outputs(2075)) or (layer6_outputs(992)));
    outputs(2496) <= not((layer6_outputs(764)) xor (layer6_outputs(2042)));
    outputs(2497) <= not(layer6_outputs(667));
    outputs(2498) <= not(layer6_outputs(1848)) or (layer6_outputs(1916));
    outputs(2499) <= (layer6_outputs(1560)) xor (layer6_outputs(1458));
    outputs(2500) <= layer6_outputs(129);
    outputs(2501) <= layer6_outputs(554);
    outputs(2502) <= not(layer6_outputs(1782));
    outputs(2503) <= not((layer6_outputs(191)) or (layer6_outputs(867)));
    outputs(2504) <= not(layer6_outputs(692));
    outputs(2505) <= layer6_outputs(1245);
    outputs(2506) <= (layer6_outputs(1175)) or (layer6_outputs(981));
    outputs(2507) <= not(layer6_outputs(1167));
    outputs(2508) <= not(layer6_outputs(122));
    outputs(2509) <= (layer6_outputs(1852)) or (layer6_outputs(1249));
    outputs(2510) <= (layer6_outputs(998)) and not (layer6_outputs(483));
    outputs(2511) <= not(layer6_outputs(1299));
    outputs(2512) <= not(layer6_outputs(2148));
    outputs(2513) <= layer6_outputs(2185);
    outputs(2514) <= not(layer6_outputs(2171));
    outputs(2515) <= layer6_outputs(858);
    outputs(2516) <= not(layer6_outputs(947));
    outputs(2517) <= (layer6_outputs(1415)) and not (layer6_outputs(643));
    outputs(2518) <= (layer6_outputs(86)) xor (layer6_outputs(1506));
    outputs(2519) <= not(layer6_outputs(1479));
    outputs(2520) <= layer6_outputs(1584);
    outputs(2521) <= not(layer6_outputs(804));
    outputs(2522) <= layer6_outputs(1107);
    outputs(2523) <= (layer6_outputs(2023)) xor (layer6_outputs(1055));
    outputs(2524) <= not(layer6_outputs(801)) or (layer6_outputs(1518));
    outputs(2525) <= not(layer6_outputs(212));
    outputs(2526) <= not(layer6_outputs(594)) or (layer6_outputs(1377));
    outputs(2527) <= (layer6_outputs(1879)) and (layer6_outputs(1078));
    outputs(2528) <= layer6_outputs(2285);
    outputs(2529) <= not(layer6_outputs(114));
    outputs(2530) <= not(layer6_outputs(2378));
    outputs(2531) <= (layer6_outputs(2039)) and (layer6_outputs(2213));
    outputs(2532) <= not(layer6_outputs(1973));
    outputs(2533) <= not(layer6_outputs(1324));
    outputs(2534) <= (layer6_outputs(306)) and (layer6_outputs(1688));
    outputs(2535) <= not(layer6_outputs(1400));
    outputs(2536) <= layer6_outputs(1153);
    outputs(2537) <= not((layer6_outputs(615)) xor (layer6_outputs(2024)));
    outputs(2538) <= not(layer6_outputs(240));
    outputs(2539) <= layer6_outputs(1254);
    outputs(2540) <= not((layer6_outputs(2125)) or (layer6_outputs(875)));
    outputs(2541) <= not((layer6_outputs(2359)) xor (layer6_outputs(2462)));
    outputs(2542) <= not(layer6_outputs(2071));
    outputs(2543) <= layer6_outputs(848);
    outputs(2544) <= layer6_outputs(572);
    outputs(2545) <= not(layer6_outputs(2152));
    outputs(2546) <= not(layer6_outputs(1812));
    outputs(2547) <= not(layer6_outputs(197));
    outputs(2548) <= (layer6_outputs(1082)) and not (layer6_outputs(994));
    outputs(2549) <= not(layer6_outputs(2040));
    outputs(2550) <= layer6_outputs(502);
    outputs(2551) <= (layer6_outputs(281)) and (layer6_outputs(2119));
    outputs(2552) <= layer6_outputs(1356);
    outputs(2553) <= layer6_outputs(1377);
    outputs(2554) <= not(layer6_outputs(1266));
    outputs(2555) <= not(layer6_outputs(2536));
    outputs(2556) <= not(layer6_outputs(2244)) or (layer6_outputs(2293));
    outputs(2557) <= not(layer6_outputs(1291)) or (layer6_outputs(2159));
    outputs(2558) <= not((layer6_outputs(183)) xor (layer6_outputs(2346)));
    outputs(2559) <= (layer6_outputs(1553)) xor (layer6_outputs(1234));

end Behavioral;
