library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(12799 downto 0);

begin

    layer0_outputs(0) <= (inputs(233)) or (inputs(14));
    layer0_outputs(1) <= not((inputs(176)) or (inputs(218)));
    layer0_outputs(2) <= not((inputs(222)) and (inputs(24)));
    layer0_outputs(3) <= not((inputs(4)) xor (inputs(163)));
    layer0_outputs(4) <= not((inputs(24)) xor (inputs(19)));
    layer0_outputs(5) <= not((inputs(119)) or (inputs(9)));
    layer0_outputs(6) <= inputs(31);
    layer0_outputs(7) <= (inputs(191)) and not (inputs(31));
    layer0_outputs(8) <= inputs(193);
    layer0_outputs(9) <= inputs(119);
    layer0_outputs(10) <= (inputs(79)) or (inputs(124));
    layer0_outputs(11) <= not((inputs(5)) xor (inputs(238)));
    layer0_outputs(12) <= (inputs(163)) or (inputs(185));
    layer0_outputs(13) <= (inputs(142)) or (inputs(72));
    layer0_outputs(14) <= not(inputs(101));
    layer0_outputs(15) <= (inputs(66)) or (inputs(20));
    layer0_outputs(16) <= (inputs(64)) and (inputs(79));
    layer0_outputs(17) <= not((inputs(213)) xor (inputs(181)));
    layer0_outputs(18) <= (inputs(144)) xor (inputs(96));
    layer0_outputs(19) <= not((inputs(118)) xor (inputs(101)));
    layer0_outputs(20) <= not(inputs(40));
    layer0_outputs(21) <= (inputs(105)) and not (inputs(149));
    layer0_outputs(22) <= (inputs(0)) xor (inputs(148));
    layer0_outputs(23) <= not(inputs(30)) or (inputs(213));
    layer0_outputs(24) <= (inputs(48)) or (inputs(232));
    layer0_outputs(25) <= not((inputs(198)) or (inputs(189)));
    layer0_outputs(26) <= (inputs(92)) and (inputs(103));
    layer0_outputs(27) <= not((inputs(182)) or (inputs(88)));
    layer0_outputs(28) <= (inputs(233)) and not (inputs(48));
    layer0_outputs(29) <= '1';
    layer0_outputs(30) <= (inputs(71)) xor (inputs(55));
    layer0_outputs(31) <= not((inputs(26)) xor (inputs(241)));
    layer0_outputs(32) <= inputs(122);
    layer0_outputs(33) <= not((inputs(166)) xor (inputs(165)));
    layer0_outputs(34) <= (inputs(171)) xor (inputs(175));
    layer0_outputs(35) <= (inputs(161)) or (inputs(209));
    layer0_outputs(36) <= inputs(171);
    layer0_outputs(37) <= inputs(191);
    layer0_outputs(38) <= (inputs(219)) or (inputs(19));
    layer0_outputs(39) <= (inputs(172)) or (inputs(112));
    layer0_outputs(40) <= not(inputs(196)) or (inputs(14));
    layer0_outputs(41) <= (inputs(204)) or (inputs(41));
    layer0_outputs(42) <= not((inputs(189)) xor (inputs(194)));
    layer0_outputs(43) <= not((inputs(125)) xor (inputs(138)));
    layer0_outputs(44) <= (inputs(243)) or (inputs(195));
    layer0_outputs(45) <= not((inputs(193)) xor (inputs(8)));
    layer0_outputs(46) <= (inputs(233)) or (inputs(95));
    layer0_outputs(47) <= not((inputs(4)) and (inputs(35)));
    layer0_outputs(48) <= not(inputs(214)) or (inputs(162));
    layer0_outputs(49) <= inputs(119);
    layer0_outputs(50) <= (inputs(135)) and not (inputs(77));
    layer0_outputs(51) <= not((inputs(187)) xor (inputs(75)));
    layer0_outputs(52) <= inputs(117);
    layer0_outputs(53) <= inputs(97);
    layer0_outputs(54) <= not(inputs(40));
    layer0_outputs(55) <= (inputs(171)) xor (inputs(98));
    layer0_outputs(56) <= (inputs(145)) xor (inputs(191));
    layer0_outputs(57) <= (inputs(14)) xor (inputs(242));
    layer0_outputs(58) <= not(inputs(21)) or (inputs(81));
    layer0_outputs(59) <= (inputs(37)) and not (inputs(246));
    layer0_outputs(60) <= (inputs(240)) or (inputs(237));
    layer0_outputs(61) <= not(inputs(105));
    layer0_outputs(62) <= '0';
    layer0_outputs(63) <= not(inputs(250)) or (inputs(16));
    layer0_outputs(64) <= not(inputs(98)) or (inputs(235));
    layer0_outputs(65) <= not((inputs(169)) xor (inputs(209)));
    layer0_outputs(66) <= not(inputs(33));
    layer0_outputs(67) <= (inputs(254)) and (inputs(7));
    layer0_outputs(68) <= not(inputs(117)) or (inputs(95));
    layer0_outputs(69) <= (inputs(189)) xor (inputs(39));
    layer0_outputs(70) <= (inputs(56)) or (inputs(97));
    layer0_outputs(71) <= not((inputs(9)) xor (inputs(184)));
    layer0_outputs(72) <= (inputs(19)) and (inputs(232));
    layer0_outputs(73) <= '0';
    layer0_outputs(74) <= not(inputs(78));
    layer0_outputs(75) <= inputs(252);
    layer0_outputs(76) <= inputs(132);
    layer0_outputs(77) <= not((inputs(36)) or (inputs(186)));
    layer0_outputs(78) <= not((inputs(221)) xor (inputs(86)));
    layer0_outputs(79) <= not((inputs(15)) xor (inputs(144)));
    layer0_outputs(80) <= inputs(140);
    layer0_outputs(81) <= not(inputs(150)) or (inputs(159));
    layer0_outputs(82) <= (inputs(13)) and (inputs(78));
    layer0_outputs(83) <= not(inputs(214)) or (inputs(194));
    layer0_outputs(84) <= not((inputs(155)) xor (inputs(134)));
    layer0_outputs(85) <= not(inputs(133));
    layer0_outputs(86) <= (inputs(18)) and not (inputs(115));
    layer0_outputs(87) <= inputs(106);
    layer0_outputs(88) <= inputs(125);
    layer0_outputs(89) <= not((inputs(209)) or (inputs(190)));
    layer0_outputs(90) <= not(inputs(217));
    layer0_outputs(91) <= (inputs(136)) and not (inputs(6));
    layer0_outputs(92) <= not((inputs(197)) or (inputs(161)));
    layer0_outputs(93) <= (inputs(20)) and (inputs(155));
    layer0_outputs(94) <= (inputs(28)) and not (inputs(105));
    layer0_outputs(95) <= (inputs(37)) and not (inputs(24));
    layer0_outputs(96) <= inputs(100);
    layer0_outputs(97) <= not(inputs(99)) or (inputs(159));
    layer0_outputs(98) <= not(inputs(9));
    layer0_outputs(99) <= (inputs(195)) and (inputs(120));
    layer0_outputs(100) <= not(inputs(210));
    layer0_outputs(101) <= (inputs(222)) or (inputs(135));
    layer0_outputs(102) <= not(inputs(245)) or (inputs(61));
    layer0_outputs(103) <= not(inputs(207));
    layer0_outputs(104) <= inputs(153);
    layer0_outputs(105) <= inputs(252);
    layer0_outputs(106) <= not(inputs(150));
    layer0_outputs(107) <= not(inputs(155));
    layer0_outputs(108) <= not(inputs(131));
    layer0_outputs(109) <= (inputs(103)) and not (inputs(17));
    layer0_outputs(110) <= inputs(155);
    layer0_outputs(111) <= not(inputs(14));
    layer0_outputs(112) <= inputs(10);
    layer0_outputs(113) <= not((inputs(54)) and (inputs(54)));
    layer0_outputs(114) <= (inputs(132)) or (inputs(210));
    layer0_outputs(115) <= not((inputs(209)) and (inputs(162)));
    layer0_outputs(116) <= inputs(140);
    layer0_outputs(117) <= (inputs(200)) xor (inputs(215));
    layer0_outputs(118) <= not((inputs(235)) and (inputs(80)));
    layer0_outputs(119) <= inputs(92);
    layer0_outputs(120) <= (inputs(71)) or (inputs(71));
    layer0_outputs(121) <= not((inputs(66)) or (inputs(33)));
    layer0_outputs(122) <= not(inputs(55));
    layer0_outputs(123) <= (inputs(82)) or (inputs(86));
    layer0_outputs(124) <= inputs(111);
    layer0_outputs(125) <= (inputs(8)) and not (inputs(169));
    layer0_outputs(126) <= (inputs(204)) and not (inputs(129));
    layer0_outputs(127) <= (inputs(117)) and not (inputs(80));
    layer0_outputs(128) <= (inputs(34)) or (inputs(219));
    layer0_outputs(129) <= (inputs(225)) or (inputs(101));
    layer0_outputs(130) <= not((inputs(71)) or (inputs(177)));
    layer0_outputs(131) <= (inputs(21)) or (inputs(210));
    layer0_outputs(132) <= (inputs(120)) xor (inputs(101));
    layer0_outputs(133) <= (inputs(125)) xor (inputs(27));
    layer0_outputs(134) <= not((inputs(234)) xor (inputs(178)));
    layer0_outputs(135) <= (inputs(64)) xor (inputs(47));
    layer0_outputs(136) <= not(inputs(166));
    layer0_outputs(137) <= inputs(232);
    layer0_outputs(138) <= inputs(86);
    layer0_outputs(139) <= not((inputs(213)) xor (inputs(18)));
    layer0_outputs(140) <= (inputs(18)) and (inputs(16));
    layer0_outputs(141) <= (inputs(8)) or (inputs(98));
    layer0_outputs(142) <= not(inputs(77));
    layer0_outputs(143) <= not(inputs(184)) or (inputs(235));
    layer0_outputs(144) <= not((inputs(55)) or (inputs(2)));
    layer0_outputs(145) <= not((inputs(49)) xor (inputs(173)));
    layer0_outputs(146) <= inputs(149);
    layer0_outputs(147) <= not(inputs(139));
    layer0_outputs(148) <= not(inputs(118));
    layer0_outputs(149) <= not((inputs(1)) xor (inputs(218)));
    layer0_outputs(150) <= not(inputs(231));
    layer0_outputs(151) <= (inputs(60)) and not (inputs(177));
    layer0_outputs(152) <= not((inputs(244)) or (inputs(169)));
    layer0_outputs(153) <= inputs(142);
    layer0_outputs(154) <= not(inputs(122));
    layer0_outputs(155) <= not(inputs(182)) or (inputs(46));
    layer0_outputs(156) <= not(inputs(56));
    layer0_outputs(157) <= inputs(205);
    layer0_outputs(158) <= inputs(18);
    layer0_outputs(159) <= not(inputs(222));
    layer0_outputs(160) <= (inputs(53)) xor (inputs(186));
    layer0_outputs(161) <= (inputs(234)) and not (inputs(110));
    layer0_outputs(162) <= not((inputs(243)) xor (inputs(29)));
    layer0_outputs(163) <= '0';
    layer0_outputs(164) <= not((inputs(233)) xor (inputs(223)));
    layer0_outputs(165) <= (inputs(81)) xor (inputs(167));
    layer0_outputs(166) <= not(inputs(88));
    layer0_outputs(167) <= not((inputs(88)) or (inputs(52)));
    layer0_outputs(168) <= not((inputs(194)) and (inputs(242)));
    layer0_outputs(169) <= (inputs(217)) xor (inputs(1));
    layer0_outputs(170) <= not(inputs(158));
    layer0_outputs(171) <= not(inputs(173));
    layer0_outputs(172) <= (inputs(108)) or (inputs(157));
    layer0_outputs(173) <= (inputs(26)) or (inputs(173));
    layer0_outputs(174) <= not(inputs(237));
    layer0_outputs(175) <= (inputs(214)) or (inputs(52));
    layer0_outputs(176) <= inputs(21);
    layer0_outputs(177) <= not((inputs(189)) or (inputs(54)));
    layer0_outputs(178) <= inputs(61);
    layer0_outputs(179) <= inputs(44);
    layer0_outputs(180) <= (inputs(152)) or (inputs(162));
    layer0_outputs(181) <= (inputs(139)) xor (inputs(240));
    layer0_outputs(182) <= not((inputs(85)) and (inputs(250)));
    layer0_outputs(183) <= inputs(43);
    layer0_outputs(184) <= not((inputs(13)) or (inputs(140)));
    layer0_outputs(185) <= inputs(141);
    layer0_outputs(186) <= not(inputs(169));
    layer0_outputs(187) <= not((inputs(60)) xor (inputs(80)));
    layer0_outputs(188) <= inputs(139);
    layer0_outputs(189) <= inputs(171);
    layer0_outputs(190) <= not((inputs(145)) xor (inputs(145)));
    layer0_outputs(191) <= (inputs(99)) and not (inputs(132));
    layer0_outputs(192) <= not(inputs(180)) or (inputs(218));
    layer0_outputs(193) <= inputs(77);
    layer0_outputs(194) <= inputs(105);
    layer0_outputs(195) <= not(inputs(66));
    layer0_outputs(196) <= not(inputs(12)) or (inputs(132));
    layer0_outputs(197) <= inputs(151);
    layer0_outputs(198) <= (inputs(64)) and not (inputs(88));
    layer0_outputs(199) <= not((inputs(26)) or (inputs(177)));
    layer0_outputs(200) <= inputs(85);
    layer0_outputs(201) <= (inputs(235)) and not (inputs(144));
    layer0_outputs(202) <= (inputs(172)) or (inputs(194));
    layer0_outputs(203) <= not((inputs(39)) xor (inputs(21)));
    layer0_outputs(204) <= not((inputs(205)) or (inputs(147)));
    layer0_outputs(205) <= (inputs(93)) or (inputs(229));
    layer0_outputs(206) <= not(inputs(15)) or (inputs(177));
    layer0_outputs(207) <= inputs(160);
    layer0_outputs(208) <= not((inputs(55)) or (inputs(199)));
    layer0_outputs(209) <= (inputs(16)) xor (inputs(190));
    layer0_outputs(210) <= inputs(131);
    layer0_outputs(211) <= not(inputs(181)) or (inputs(146));
    layer0_outputs(212) <= not(inputs(59));
    layer0_outputs(213) <= (inputs(245)) and (inputs(237));
    layer0_outputs(214) <= (inputs(230)) or (inputs(204));
    layer0_outputs(215) <= not((inputs(75)) xor (inputs(61)));
    layer0_outputs(216) <= (inputs(29)) or (inputs(157));
    layer0_outputs(217) <= (inputs(180)) and not (inputs(223));
    layer0_outputs(218) <= not(inputs(231)) or (inputs(188));
    layer0_outputs(219) <= not(inputs(216));
    layer0_outputs(220) <= not(inputs(85));
    layer0_outputs(221) <= not(inputs(83)) or (inputs(136));
    layer0_outputs(222) <= (inputs(69)) and not (inputs(21));
    layer0_outputs(223) <= not((inputs(171)) xor (inputs(117)));
    layer0_outputs(224) <= inputs(171);
    layer0_outputs(225) <= not((inputs(23)) or (inputs(154)));
    layer0_outputs(226) <= (inputs(118)) xor (inputs(235));
    layer0_outputs(227) <= not((inputs(101)) or (inputs(145)));
    layer0_outputs(228) <= inputs(77);
    layer0_outputs(229) <= (inputs(129)) and not (inputs(42));
    layer0_outputs(230) <= '0';
    layer0_outputs(231) <= not(inputs(213));
    layer0_outputs(232) <= not((inputs(116)) and (inputs(238)));
    layer0_outputs(233) <= not(inputs(199)) or (inputs(255));
    layer0_outputs(234) <= not(inputs(102));
    layer0_outputs(235) <= inputs(13);
    layer0_outputs(236) <= '1';
    layer0_outputs(237) <= not((inputs(167)) xor (inputs(207)));
    layer0_outputs(238) <= not((inputs(227)) or (inputs(211)));
    layer0_outputs(239) <= not((inputs(244)) or (inputs(47)));
    layer0_outputs(240) <= (inputs(178)) and (inputs(243));
    layer0_outputs(241) <= '1';
    layer0_outputs(242) <= (inputs(147)) xor (inputs(53));
    layer0_outputs(243) <= inputs(66);
    layer0_outputs(244) <= (inputs(237)) and not (inputs(253));
    layer0_outputs(245) <= (inputs(143)) and not (inputs(188));
    layer0_outputs(246) <= (inputs(12)) or (inputs(249));
    layer0_outputs(247) <= inputs(249);
    layer0_outputs(248) <= not(inputs(199));
    layer0_outputs(249) <= (inputs(46)) xor (inputs(74));
    layer0_outputs(250) <= (inputs(44)) or (inputs(139));
    layer0_outputs(251) <= not((inputs(239)) xor (inputs(42)));
    layer0_outputs(252) <= '1';
    layer0_outputs(253) <= (inputs(200)) or (inputs(182));
    layer0_outputs(254) <= (inputs(209)) or (inputs(56));
    layer0_outputs(255) <= inputs(13);
    layer0_outputs(256) <= not(inputs(192));
    layer0_outputs(257) <= not(inputs(151)) or (inputs(232));
    layer0_outputs(258) <= not(inputs(97)) or (inputs(238));
    layer0_outputs(259) <= (inputs(203)) or (inputs(110));
    layer0_outputs(260) <= not((inputs(237)) xor (inputs(35)));
    layer0_outputs(261) <= (inputs(209)) and (inputs(95));
    layer0_outputs(262) <= (inputs(222)) xor (inputs(103));
    layer0_outputs(263) <= not((inputs(176)) or (inputs(100)));
    layer0_outputs(264) <= (inputs(156)) or (inputs(248));
    layer0_outputs(265) <= not(inputs(134)) or (inputs(236));
    layer0_outputs(266) <= not(inputs(56));
    layer0_outputs(267) <= (inputs(73)) and not (inputs(25));
    layer0_outputs(268) <= (inputs(18)) and not (inputs(220));
    layer0_outputs(269) <= not((inputs(194)) xor (inputs(28)));
    layer0_outputs(270) <= not(inputs(212));
    layer0_outputs(271) <= '1';
    layer0_outputs(272) <= not(inputs(131)) or (inputs(254));
    layer0_outputs(273) <= inputs(83);
    layer0_outputs(274) <= not((inputs(94)) xor (inputs(219)));
    layer0_outputs(275) <= (inputs(194)) xor (inputs(44));
    layer0_outputs(276) <= (inputs(221)) and not (inputs(225));
    layer0_outputs(277) <= not((inputs(232)) or (inputs(193)));
    layer0_outputs(278) <= '1';
    layer0_outputs(279) <= (inputs(219)) and not (inputs(237));
    layer0_outputs(280) <= not(inputs(198)) or (inputs(207));
    layer0_outputs(281) <= (inputs(180)) and not (inputs(100));
    layer0_outputs(282) <= not(inputs(163)) or (inputs(79));
    layer0_outputs(283) <= not(inputs(241));
    layer0_outputs(284) <= inputs(215);
    layer0_outputs(285) <= not((inputs(22)) xor (inputs(206)));
    layer0_outputs(286) <= '1';
    layer0_outputs(287) <= not(inputs(164));
    layer0_outputs(288) <= inputs(247);
    layer0_outputs(289) <= not(inputs(200)) or (inputs(62));
    layer0_outputs(290) <= '0';
    layer0_outputs(291) <= not((inputs(23)) or (inputs(221)));
    layer0_outputs(292) <= not((inputs(235)) or (inputs(181)));
    layer0_outputs(293) <= not(inputs(28)) or (inputs(243));
    layer0_outputs(294) <= not(inputs(157));
    layer0_outputs(295) <= not((inputs(183)) or (inputs(80)));
    layer0_outputs(296) <= not((inputs(214)) and (inputs(124)));
    layer0_outputs(297) <= inputs(153);
    layer0_outputs(298) <= not((inputs(177)) xor (inputs(194)));
    layer0_outputs(299) <= not((inputs(51)) or (inputs(121)));
    layer0_outputs(300) <= not(inputs(245)) or (inputs(178));
    layer0_outputs(301) <= (inputs(240)) and not (inputs(109));
    layer0_outputs(302) <= '0';
    layer0_outputs(303) <= not(inputs(196)) or (inputs(37));
    layer0_outputs(304) <= not(inputs(224));
    layer0_outputs(305) <= (inputs(74)) xor (inputs(217));
    layer0_outputs(306) <= inputs(89);
    layer0_outputs(307) <= (inputs(165)) and not (inputs(242));
    layer0_outputs(308) <= not((inputs(168)) xor (inputs(10)));
    layer0_outputs(309) <= not((inputs(66)) xor (inputs(84)));
    layer0_outputs(310) <= (inputs(27)) and not (inputs(18));
    layer0_outputs(311) <= (inputs(41)) xor (inputs(166));
    layer0_outputs(312) <= inputs(47);
    layer0_outputs(313) <= '0';
    layer0_outputs(314) <= not(inputs(10)) or (inputs(127));
    layer0_outputs(315) <= (inputs(61)) xor (inputs(243));
    layer0_outputs(316) <= inputs(170);
    layer0_outputs(317) <= not(inputs(30)) or (inputs(84));
    layer0_outputs(318) <= (inputs(243)) xor (inputs(154));
    layer0_outputs(319) <= (inputs(87)) and not (inputs(220));
    layer0_outputs(320) <= not(inputs(114)) or (inputs(224));
    layer0_outputs(321) <= not(inputs(152));
    layer0_outputs(322) <= not((inputs(163)) xor (inputs(155)));
    layer0_outputs(323) <= (inputs(254)) and not (inputs(0));
    layer0_outputs(324) <= inputs(152);
    layer0_outputs(325) <= inputs(211);
    layer0_outputs(326) <= not(inputs(152));
    layer0_outputs(327) <= inputs(120);
    layer0_outputs(328) <= inputs(119);
    layer0_outputs(329) <= not((inputs(153)) xor (inputs(82)));
    layer0_outputs(330) <= not(inputs(150));
    layer0_outputs(331) <= not((inputs(254)) and (inputs(244)));
    layer0_outputs(332) <= (inputs(249)) and not (inputs(84));
    layer0_outputs(333) <= (inputs(238)) or (inputs(183));
    layer0_outputs(334) <= not(inputs(166));
    layer0_outputs(335) <= not(inputs(88));
    layer0_outputs(336) <= not(inputs(216)) or (inputs(246));
    layer0_outputs(337) <= not(inputs(37)) or (inputs(184));
    layer0_outputs(338) <= (inputs(127)) xor (inputs(148));
    layer0_outputs(339) <= inputs(170);
    layer0_outputs(340) <= inputs(48);
    layer0_outputs(341) <= inputs(15);
    layer0_outputs(342) <= (inputs(30)) and not (inputs(63));
    layer0_outputs(343) <= '1';
    layer0_outputs(344) <= (inputs(102)) and not (inputs(235));
    layer0_outputs(345) <= not((inputs(91)) xor (inputs(7)));
    layer0_outputs(346) <= (inputs(33)) xor (inputs(235));
    layer0_outputs(347) <= not(inputs(211));
    layer0_outputs(348) <= (inputs(80)) xor (inputs(108));
    layer0_outputs(349) <= not((inputs(147)) or (inputs(216)));
    layer0_outputs(350) <= not(inputs(139));
    layer0_outputs(351) <= not((inputs(144)) xor (inputs(110)));
    layer0_outputs(352) <= (inputs(239)) and not (inputs(254));
    layer0_outputs(353) <= not((inputs(49)) xor (inputs(230)));
    layer0_outputs(354) <= (inputs(241)) xor (inputs(73));
    layer0_outputs(355) <= (inputs(24)) and not (inputs(245));
    layer0_outputs(356) <= not((inputs(112)) and (inputs(227)));
    layer0_outputs(357) <= not((inputs(159)) xor (inputs(202)));
    layer0_outputs(358) <= not((inputs(128)) or (inputs(60)));
    layer0_outputs(359) <= (inputs(6)) or (inputs(220));
    layer0_outputs(360) <= not((inputs(192)) or (inputs(137)));
    layer0_outputs(361) <= not((inputs(154)) xor (inputs(71)));
    layer0_outputs(362) <= (inputs(229)) and not (inputs(49));
    layer0_outputs(363) <= (inputs(42)) or (inputs(166));
    layer0_outputs(364) <= (inputs(197)) or (inputs(0));
    layer0_outputs(365) <= not((inputs(191)) and (inputs(98)));
    layer0_outputs(366) <= '0';
    layer0_outputs(367) <= not(inputs(84)) or (inputs(71));
    layer0_outputs(368) <= not(inputs(89)) or (inputs(96));
    layer0_outputs(369) <= '1';
    layer0_outputs(370) <= not(inputs(115));
    layer0_outputs(371) <= not(inputs(141));
    layer0_outputs(372) <= not((inputs(34)) xor (inputs(162)));
    layer0_outputs(373) <= (inputs(252)) or (inputs(7));
    layer0_outputs(374) <= '0';
    layer0_outputs(375) <= not(inputs(255)) or (inputs(209));
    layer0_outputs(376) <= not((inputs(139)) xor (inputs(13)));
    layer0_outputs(377) <= inputs(108);
    layer0_outputs(378) <= (inputs(168)) or (inputs(168));
    layer0_outputs(379) <= not(inputs(154)) or (inputs(231));
    layer0_outputs(380) <= inputs(100);
    layer0_outputs(381) <= not(inputs(231));
    layer0_outputs(382) <= '1';
    layer0_outputs(383) <= (inputs(245)) and (inputs(100));
    layer0_outputs(384) <= not(inputs(91));
    layer0_outputs(385) <= '1';
    layer0_outputs(386) <= (inputs(5)) and (inputs(254));
    layer0_outputs(387) <= (inputs(61)) and not (inputs(180));
    layer0_outputs(388) <= not(inputs(167));
    layer0_outputs(389) <= (inputs(161)) xor (inputs(58));
    layer0_outputs(390) <= not((inputs(92)) or (inputs(235)));
    layer0_outputs(391) <= (inputs(239)) and not (inputs(198));
    layer0_outputs(392) <= (inputs(153)) and not (inputs(217));
    layer0_outputs(393) <= inputs(64);
    layer0_outputs(394) <= not((inputs(79)) and (inputs(208)));
    layer0_outputs(395) <= inputs(254);
    layer0_outputs(396) <= inputs(186);
    layer0_outputs(397) <= (inputs(242)) and not (inputs(193));
    layer0_outputs(398) <= not((inputs(255)) xor (inputs(100)));
    layer0_outputs(399) <= inputs(182);
    layer0_outputs(400) <= not(inputs(153)) or (inputs(221));
    layer0_outputs(401) <= not((inputs(213)) or (inputs(231)));
    layer0_outputs(402) <= not((inputs(43)) xor (inputs(154)));
    layer0_outputs(403) <= not(inputs(163)) or (inputs(225));
    layer0_outputs(404) <= not(inputs(171)) or (inputs(249));
    layer0_outputs(405) <= (inputs(18)) xor (inputs(104));
    layer0_outputs(406) <= not((inputs(51)) xor (inputs(14)));
    layer0_outputs(407) <= (inputs(184)) and not (inputs(249));
    layer0_outputs(408) <= not(inputs(125));
    layer0_outputs(409) <= inputs(181);
    layer0_outputs(410) <= (inputs(246)) and not (inputs(174));
    layer0_outputs(411) <= (inputs(120)) and not (inputs(187));
    layer0_outputs(412) <= (inputs(232)) and (inputs(193));
    layer0_outputs(413) <= not((inputs(17)) or (inputs(53)));
    layer0_outputs(414) <= not((inputs(84)) or (inputs(1)));
    layer0_outputs(415) <= (inputs(102)) and not (inputs(25));
    layer0_outputs(416) <= (inputs(23)) and not (inputs(250));
    layer0_outputs(417) <= (inputs(128)) and (inputs(135));
    layer0_outputs(418) <= '1';
    layer0_outputs(419) <= inputs(244);
    layer0_outputs(420) <= not((inputs(77)) xor (inputs(46)));
    layer0_outputs(421) <= (inputs(131)) or (inputs(208));
    layer0_outputs(422) <= (inputs(119)) or (inputs(55));
    layer0_outputs(423) <= not(inputs(219));
    layer0_outputs(424) <= not((inputs(77)) xor (inputs(51)));
    layer0_outputs(425) <= (inputs(17)) or (inputs(139));
    layer0_outputs(426) <= inputs(165);
    layer0_outputs(427) <= not((inputs(120)) xor (inputs(100)));
    layer0_outputs(428) <= not((inputs(192)) and (inputs(193)));
    layer0_outputs(429) <= not((inputs(98)) or (inputs(227)));
    layer0_outputs(430) <= not(inputs(214));
    layer0_outputs(431) <= not(inputs(213)) or (inputs(141));
    layer0_outputs(432) <= not((inputs(6)) or (inputs(162)));
    layer0_outputs(433) <= not((inputs(95)) xor (inputs(213)));
    layer0_outputs(434) <= (inputs(210)) xor (inputs(100));
    layer0_outputs(435) <= (inputs(177)) and not (inputs(228));
    layer0_outputs(436) <= not(inputs(191));
    layer0_outputs(437) <= not((inputs(179)) xor (inputs(44)));
    layer0_outputs(438) <= inputs(67);
    layer0_outputs(439) <= not(inputs(197));
    layer0_outputs(440) <= inputs(51);
    layer0_outputs(441) <= not(inputs(163)) or (inputs(233));
    layer0_outputs(442) <= not(inputs(216)) or (inputs(6));
    layer0_outputs(443) <= not(inputs(175)) or (inputs(196));
    layer0_outputs(444) <= not(inputs(220));
    layer0_outputs(445) <= not((inputs(139)) xor (inputs(249)));
    layer0_outputs(446) <= inputs(135);
    layer0_outputs(447) <= not((inputs(196)) or (inputs(2)));
    layer0_outputs(448) <= (inputs(34)) and not (inputs(42));
    layer0_outputs(449) <= not((inputs(21)) or (inputs(165)));
    layer0_outputs(450) <= inputs(48);
    layer0_outputs(451) <= not(inputs(213));
    layer0_outputs(452) <= not((inputs(109)) or (inputs(17)));
    layer0_outputs(453) <= (inputs(63)) and (inputs(188));
    layer0_outputs(454) <= inputs(149);
    layer0_outputs(455) <= not(inputs(25)) or (inputs(94));
    layer0_outputs(456) <= not(inputs(178));
    layer0_outputs(457) <= not((inputs(191)) xor (inputs(141)));
    layer0_outputs(458) <= not((inputs(135)) xor (inputs(2)));
    layer0_outputs(459) <= (inputs(63)) xor (inputs(242));
    layer0_outputs(460) <= not(inputs(231)) or (inputs(80));
    layer0_outputs(461) <= not(inputs(198)) or (inputs(159));
    layer0_outputs(462) <= not(inputs(113));
    layer0_outputs(463) <= (inputs(123)) and (inputs(155));
    layer0_outputs(464) <= inputs(48);
    layer0_outputs(465) <= (inputs(168)) xor (inputs(148));
    layer0_outputs(466) <= not(inputs(43)) or (inputs(147));
    layer0_outputs(467) <= (inputs(136)) or (inputs(104));
    layer0_outputs(468) <= (inputs(206)) or (inputs(189));
    layer0_outputs(469) <= (inputs(116)) and not (inputs(22));
    layer0_outputs(470) <= not(inputs(163));
    layer0_outputs(471) <= not((inputs(252)) or (inputs(146)));
    layer0_outputs(472) <= (inputs(181)) and not (inputs(208));
    layer0_outputs(473) <= not((inputs(231)) or (inputs(236)));
    layer0_outputs(474) <= not((inputs(208)) or (inputs(241)));
    layer0_outputs(475) <= inputs(125);
    layer0_outputs(476) <= not((inputs(101)) or (inputs(68)));
    layer0_outputs(477) <= not(inputs(138)) or (inputs(124));
    layer0_outputs(478) <= (inputs(21)) or (inputs(94));
    layer0_outputs(479) <= inputs(123);
    layer0_outputs(480) <= not((inputs(153)) or (inputs(236)));
    layer0_outputs(481) <= not((inputs(138)) xor (inputs(149)));
    layer0_outputs(482) <= (inputs(92)) and (inputs(121));
    layer0_outputs(483) <= not(inputs(164)) or (inputs(160));
    layer0_outputs(484) <= not(inputs(158));
    layer0_outputs(485) <= (inputs(5)) and not (inputs(12));
    layer0_outputs(486) <= (inputs(190)) or (inputs(84));
    layer0_outputs(487) <= not((inputs(26)) xor (inputs(6)));
    layer0_outputs(488) <= not((inputs(56)) xor (inputs(222)));
    layer0_outputs(489) <= inputs(98);
    layer0_outputs(490) <= (inputs(174)) or (inputs(181));
    layer0_outputs(491) <= inputs(241);
    layer0_outputs(492) <= not(inputs(17)) or (inputs(212));
    layer0_outputs(493) <= inputs(74);
    layer0_outputs(494) <= not(inputs(225)) or (inputs(20));
    layer0_outputs(495) <= not((inputs(225)) xor (inputs(61)));
    layer0_outputs(496) <= not(inputs(56));
    layer0_outputs(497) <= (inputs(124)) or (inputs(227));
    layer0_outputs(498) <= not(inputs(228)) or (inputs(194));
    layer0_outputs(499) <= (inputs(92)) and not (inputs(138));
    layer0_outputs(500) <= not(inputs(69));
    layer0_outputs(501) <= not((inputs(126)) or (inputs(56)));
    layer0_outputs(502) <= not((inputs(112)) and (inputs(49)));
    layer0_outputs(503) <= not((inputs(200)) or (inputs(6)));
    layer0_outputs(504) <= inputs(133);
    layer0_outputs(505) <= (inputs(166)) and not (inputs(54));
    layer0_outputs(506) <= inputs(121);
    layer0_outputs(507) <= (inputs(169)) and not (inputs(83));
    layer0_outputs(508) <= (inputs(188)) and not (inputs(247));
    layer0_outputs(509) <= not((inputs(199)) or (inputs(41)));
    layer0_outputs(510) <= (inputs(181)) and not (inputs(57));
    layer0_outputs(511) <= not((inputs(84)) xor (inputs(204)));
    layer0_outputs(512) <= not((inputs(11)) or (inputs(106)));
    layer0_outputs(513) <= not((inputs(20)) or (inputs(16)));
    layer0_outputs(514) <= not((inputs(162)) xor (inputs(202)));
    layer0_outputs(515) <= inputs(116);
    layer0_outputs(516) <= not((inputs(29)) or (inputs(184)));
    layer0_outputs(517) <= inputs(43);
    layer0_outputs(518) <= (inputs(155)) xor (inputs(253));
    layer0_outputs(519) <= not(inputs(167));
    layer0_outputs(520) <= (inputs(17)) or (inputs(22));
    layer0_outputs(521) <= inputs(155);
    layer0_outputs(522) <= not((inputs(2)) xor (inputs(17)));
    layer0_outputs(523) <= (inputs(112)) and not (inputs(19));
    layer0_outputs(524) <= (inputs(10)) or (inputs(124));
    layer0_outputs(525) <= (inputs(196)) or (inputs(162));
    layer0_outputs(526) <= not((inputs(250)) or (inputs(140)));
    layer0_outputs(527) <= (inputs(41)) xor (inputs(212));
    layer0_outputs(528) <= (inputs(16)) and (inputs(253));
    layer0_outputs(529) <= inputs(119);
    layer0_outputs(530) <= not(inputs(10)) or (inputs(175));
    layer0_outputs(531) <= not(inputs(245));
    layer0_outputs(532) <= inputs(68);
    layer0_outputs(533) <= inputs(140);
    layer0_outputs(534) <= not((inputs(45)) or (inputs(136)));
    layer0_outputs(535) <= inputs(252);
    layer0_outputs(536) <= inputs(215);
    layer0_outputs(537) <= not(inputs(182)) or (inputs(114));
    layer0_outputs(538) <= not((inputs(31)) xor (inputs(82)));
    layer0_outputs(539) <= not((inputs(138)) xor (inputs(81)));
    layer0_outputs(540) <= not((inputs(33)) xor (inputs(39)));
    layer0_outputs(541) <= (inputs(218)) and not (inputs(255));
    layer0_outputs(542) <= not(inputs(241)) or (inputs(144));
    layer0_outputs(543) <= inputs(94);
    layer0_outputs(544) <= not((inputs(147)) or (inputs(116)));
    layer0_outputs(545) <= (inputs(123)) xor (inputs(175));
    layer0_outputs(546) <= (inputs(174)) or (inputs(157));
    layer0_outputs(547) <= inputs(16);
    layer0_outputs(548) <= inputs(57);
    layer0_outputs(549) <= not(inputs(223)) or (inputs(127));
    layer0_outputs(550) <= (inputs(18)) xor (inputs(92));
    layer0_outputs(551) <= not((inputs(231)) or (inputs(136)));
    layer0_outputs(552) <= (inputs(245)) or (inputs(185));
    layer0_outputs(553) <= not(inputs(141));
    layer0_outputs(554) <= (inputs(252)) and (inputs(65));
    layer0_outputs(555) <= not((inputs(44)) or (inputs(10)));
    layer0_outputs(556) <= not((inputs(182)) xor (inputs(51)));
    layer0_outputs(557) <= (inputs(232)) xor (inputs(160));
    layer0_outputs(558) <= (inputs(122)) or (inputs(38));
    layer0_outputs(559) <= (inputs(25)) and not (inputs(76));
    layer0_outputs(560) <= inputs(164);
    layer0_outputs(561) <= '0';
    layer0_outputs(562) <= (inputs(21)) and not (inputs(1));
    layer0_outputs(563) <= not(inputs(50));
    layer0_outputs(564) <= not(inputs(107)) or (inputs(51));
    layer0_outputs(565) <= not(inputs(208));
    layer0_outputs(566) <= inputs(182);
    layer0_outputs(567) <= (inputs(140)) or (inputs(163));
    layer0_outputs(568) <= not((inputs(180)) or (inputs(98)));
    layer0_outputs(569) <= not(inputs(179));
    layer0_outputs(570) <= not(inputs(227));
    layer0_outputs(571) <= not((inputs(30)) xor (inputs(253)));
    layer0_outputs(572) <= (inputs(209)) xor (inputs(86));
    layer0_outputs(573) <= inputs(147);
    layer0_outputs(574) <= not((inputs(181)) or (inputs(197)));
    layer0_outputs(575) <= (inputs(41)) and not (inputs(194));
    layer0_outputs(576) <= (inputs(106)) or (inputs(36));
    layer0_outputs(577) <= (inputs(211)) and not (inputs(27));
    layer0_outputs(578) <= (inputs(20)) or (inputs(51));
    layer0_outputs(579) <= '1';
    layer0_outputs(580) <= (inputs(8)) and not (inputs(32));
    layer0_outputs(581) <= (inputs(153)) and not (inputs(171));
    layer0_outputs(582) <= '1';
    layer0_outputs(583) <= not((inputs(241)) or (inputs(182)));
    layer0_outputs(584) <= inputs(173);
    layer0_outputs(585) <= not(inputs(68));
    layer0_outputs(586) <= (inputs(200)) or (inputs(61));
    layer0_outputs(587) <= not((inputs(245)) or (inputs(120)));
    layer0_outputs(588) <= not((inputs(134)) xor (inputs(231)));
    layer0_outputs(589) <= not((inputs(218)) or (inputs(30)));
    layer0_outputs(590) <= (inputs(129)) or (inputs(92));
    layer0_outputs(591) <= not((inputs(208)) xor (inputs(86)));
    layer0_outputs(592) <= (inputs(187)) xor (inputs(41));
    layer0_outputs(593) <= (inputs(1)) and (inputs(7));
    layer0_outputs(594) <= not(inputs(178));
    layer0_outputs(595) <= (inputs(220)) and not (inputs(192));
    layer0_outputs(596) <= not(inputs(213));
    layer0_outputs(597) <= inputs(149);
    layer0_outputs(598) <= (inputs(204)) and not (inputs(97));
    layer0_outputs(599) <= (inputs(119)) and not (inputs(53));
    layer0_outputs(600) <= not((inputs(99)) and (inputs(48)));
    layer0_outputs(601) <= (inputs(120)) and not (inputs(122));
    layer0_outputs(602) <= '1';
    layer0_outputs(603) <= not(inputs(49)) or (inputs(207));
    layer0_outputs(604) <= inputs(92);
    layer0_outputs(605) <= '1';
    layer0_outputs(606) <= (inputs(184)) and not (inputs(12));
    layer0_outputs(607) <= not((inputs(119)) or (inputs(139)));
    layer0_outputs(608) <= (inputs(168)) and not (inputs(157));
    layer0_outputs(609) <= not((inputs(189)) or (inputs(123)));
    layer0_outputs(610) <= (inputs(109)) xor (inputs(226));
    layer0_outputs(611) <= (inputs(103)) and not (inputs(206));
    layer0_outputs(612) <= not(inputs(231));
    layer0_outputs(613) <= (inputs(247)) xor (inputs(253));
    layer0_outputs(614) <= not(inputs(102)) or (inputs(46));
    layer0_outputs(615) <= not(inputs(124));
    layer0_outputs(616) <= inputs(67);
    layer0_outputs(617) <= not((inputs(23)) xor (inputs(87)));
    layer0_outputs(618) <= not(inputs(89));
    layer0_outputs(619) <= (inputs(89)) and not (inputs(247));
    layer0_outputs(620) <= not(inputs(232)) or (inputs(185));
    layer0_outputs(621) <= inputs(137);
    layer0_outputs(622) <= not(inputs(230));
    layer0_outputs(623) <= inputs(215);
    layer0_outputs(624) <= not(inputs(106));
    layer0_outputs(625) <= not(inputs(88));
    layer0_outputs(626) <= not(inputs(116));
    layer0_outputs(627) <= (inputs(79)) and not (inputs(112));
    layer0_outputs(628) <= (inputs(184)) and (inputs(68));
    layer0_outputs(629) <= (inputs(247)) xor (inputs(43));
    layer0_outputs(630) <= not(inputs(168));
    layer0_outputs(631) <= not(inputs(247)) or (inputs(126));
    layer0_outputs(632) <= (inputs(195)) or (inputs(44));
    layer0_outputs(633) <= inputs(252);
    layer0_outputs(634) <= not((inputs(196)) xor (inputs(140)));
    layer0_outputs(635) <= not(inputs(36)) or (inputs(41));
    layer0_outputs(636) <= (inputs(86)) or (inputs(139));
    layer0_outputs(637) <= (inputs(137)) and (inputs(118));
    layer0_outputs(638) <= (inputs(37)) and (inputs(96));
    layer0_outputs(639) <= (inputs(187)) and not (inputs(252));
    layer0_outputs(640) <= not(inputs(23)) or (inputs(245));
    layer0_outputs(641) <= (inputs(53)) or (inputs(214));
    layer0_outputs(642) <= inputs(127);
    layer0_outputs(643) <= '1';
    layer0_outputs(644) <= not((inputs(223)) or (inputs(91)));
    layer0_outputs(645) <= (inputs(28)) and not (inputs(19));
    layer0_outputs(646) <= not(inputs(80));
    layer0_outputs(647) <= (inputs(233)) xor (inputs(197));
    layer0_outputs(648) <= inputs(166);
    layer0_outputs(649) <= inputs(77);
    layer0_outputs(650) <= (inputs(150)) and not (inputs(195));
    layer0_outputs(651) <= inputs(67);
    layer0_outputs(652) <= '0';
    layer0_outputs(653) <= (inputs(195)) or (inputs(199));
    layer0_outputs(654) <= inputs(112);
    layer0_outputs(655) <= not((inputs(192)) and (inputs(79)));
    layer0_outputs(656) <= not((inputs(225)) or (inputs(81)));
    layer0_outputs(657) <= inputs(151);
    layer0_outputs(658) <= (inputs(83)) or (inputs(213));
    layer0_outputs(659) <= '1';
    layer0_outputs(660) <= (inputs(78)) and (inputs(32));
    layer0_outputs(661) <= (inputs(106)) and not (inputs(140));
    layer0_outputs(662) <= not(inputs(89)) or (inputs(99));
    layer0_outputs(663) <= not((inputs(171)) or (inputs(81)));
    layer0_outputs(664) <= (inputs(166)) xor (inputs(52));
    layer0_outputs(665) <= (inputs(213)) or (inputs(213));
    layer0_outputs(666) <= not((inputs(204)) or (inputs(203)));
    layer0_outputs(667) <= not(inputs(100));
    layer0_outputs(668) <= '1';
    layer0_outputs(669) <= (inputs(109)) or (inputs(172));
    layer0_outputs(670) <= (inputs(18)) xor (inputs(96));
    layer0_outputs(671) <= (inputs(93)) and not (inputs(111));
    layer0_outputs(672) <= (inputs(65)) xor (inputs(164));
    layer0_outputs(673) <= inputs(15);
    layer0_outputs(674) <= '1';
    layer0_outputs(675) <= inputs(205);
    layer0_outputs(676) <= not(inputs(231)) or (inputs(244));
    layer0_outputs(677) <= not((inputs(213)) xor (inputs(249)));
    layer0_outputs(678) <= not((inputs(151)) or (inputs(38)));
    layer0_outputs(679) <= (inputs(248)) xor (inputs(201));
    layer0_outputs(680) <= not((inputs(208)) and (inputs(188)));
    layer0_outputs(681) <= not(inputs(215));
    layer0_outputs(682) <= inputs(151);
    layer0_outputs(683) <= (inputs(72)) and not (inputs(167));
    layer0_outputs(684) <= (inputs(247)) or (inputs(169));
    layer0_outputs(685) <= (inputs(121)) and not (inputs(44));
    layer0_outputs(686) <= (inputs(1)) xor (inputs(152));
    layer0_outputs(687) <= (inputs(166)) xor (inputs(28));
    layer0_outputs(688) <= (inputs(25)) xor (inputs(254));
    layer0_outputs(689) <= not((inputs(18)) or (inputs(231)));
    layer0_outputs(690) <= (inputs(194)) xor (inputs(205));
    layer0_outputs(691) <= (inputs(241)) xor (inputs(200));
    layer0_outputs(692) <= not(inputs(130));
    layer0_outputs(693) <= not((inputs(37)) xor (inputs(70)));
    layer0_outputs(694) <= (inputs(254)) and not (inputs(7));
    layer0_outputs(695) <= inputs(54);
    layer0_outputs(696) <= not(inputs(131));
    layer0_outputs(697) <= '0';
    layer0_outputs(698) <= (inputs(216)) xor (inputs(16));
    layer0_outputs(699) <= not((inputs(57)) xor (inputs(93)));
    layer0_outputs(700) <= (inputs(44)) xor (inputs(188));
    layer0_outputs(701) <= not((inputs(9)) xor (inputs(216)));
    layer0_outputs(702) <= inputs(117);
    layer0_outputs(703) <= not(inputs(114));
    layer0_outputs(704) <= (inputs(35)) xor (inputs(51));
    layer0_outputs(705) <= not(inputs(153)) or (inputs(191));
    layer0_outputs(706) <= (inputs(64)) and not (inputs(199));
    layer0_outputs(707) <= not(inputs(168)) or (inputs(155));
    layer0_outputs(708) <= not(inputs(104));
    layer0_outputs(709) <= not((inputs(55)) or (inputs(41)));
    layer0_outputs(710) <= not((inputs(212)) xor (inputs(171)));
    layer0_outputs(711) <= not((inputs(114)) or (inputs(61)));
    layer0_outputs(712) <= (inputs(228)) and not (inputs(146));
    layer0_outputs(713) <= (inputs(4)) and not (inputs(1));
    layer0_outputs(714) <= inputs(76);
    layer0_outputs(715) <= '0';
    layer0_outputs(716) <= not((inputs(221)) and (inputs(147)));
    layer0_outputs(717) <= not(inputs(156)) or (inputs(221));
    layer0_outputs(718) <= not((inputs(55)) or (inputs(93)));
    layer0_outputs(719) <= (inputs(54)) or (inputs(110));
    layer0_outputs(720) <= (inputs(90)) xor (inputs(250));
    layer0_outputs(721) <= not((inputs(25)) xor (inputs(77)));
    layer0_outputs(722) <= (inputs(131)) xor (inputs(32));
    layer0_outputs(723) <= not((inputs(125)) or (inputs(10)));
    layer0_outputs(724) <= (inputs(29)) and not (inputs(51));
    layer0_outputs(725) <= not((inputs(163)) or (inputs(213)));
    layer0_outputs(726) <= not(inputs(7));
    layer0_outputs(727) <= not((inputs(229)) xor (inputs(142)));
    layer0_outputs(728) <= (inputs(168)) or (inputs(5));
    layer0_outputs(729) <= not((inputs(43)) xor (inputs(41)));
    layer0_outputs(730) <= inputs(80);
    layer0_outputs(731) <= '0';
    layer0_outputs(732) <= not((inputs(94)) or (inputs(185)));
    layer0_outputs(733) <= not((inputs(136)) or (inputs(125)));
    layer0_outputs(734) <= not(inputs(7)) or (inputs(127));
    layer0_outputs(735) <= not((inputs(197)) xor (inputs(100)));
    layer0_outputs(736) <= '0';
    layer0_outputs(737) <= not(inputs(40));
    layer0_outputs(738) <= inputs(43);
    layer0_outputs(739) <= (inputs(219)) xor (inputs(129));
    layer0_outputs(740) <= not(inputs(168)) or (inputs(158));
    layer0_outputs(741) <= not(inputs(27)) or (inputs(82));
    layer0_outputs(742) <= not(inputs(40));
    layer0_outputs(743) <= not((inputs(129)) xor (inputs(221)));
    layer0_outputs(744) <= (inputs(60)) or (inputs(106));
    layer0_outputs(745) <= not((inputs(161)) xor (inputs(157)));
    layer0_outputs(746) <= (inputs(215)) xor (inputs(96));
    layer0_outputs(747) <= '1';
    layer0_outputs(748) <= not(inputs(44)) or (inputs(37));
    layer0_outputs(749) <= (inputs(205)) and not (inputs(97));
    layer0_outputs(750) <= (inputs(172)) and not (inputs(23));
    layer0_outputs(751) <= '0';
    layer0_outputs(752) <= not(inputs(176));
    layer0_outputs(753) <= (inputs(235)) and (inputs(221));
    layer0_outputs(754) <= inputs(169);
    layer0_outputs(755) <= not((inputs(110)) or (inputs(81)));
    layer0_outputs(756) <= (inputs(86)) or (inputs(1));
    layer0_outputs(757) <= not(inputs(72));
    layer0_outputs(758) <= not(inputs(187)) or (inputs(10));
    layer0_outputs(759) <= (inputs(122)) or (inputs(47));
    layer0_outputs(760) <= (inputs(74)) or (inputs(91));
    layer0_outputs(761) <= inputs(169);
    layer0_outputs(762) <= (inputs(85)) and not (inputs(134));
    layer0_outputs(763) <= inputs(131);
    layer0_outputs(764) <= (inputs(198)) or (inputs(179));
    layer0_outputs(765) <= not((inputs(196)) xor (inputs(230)));
    layer0_outputs(766) <= not((inputs(52)) and (inputs(52)));
    layer0_outputs(767) <= (inputs(118)) or (inputs(80));
    layer0_outputs(768) <= (inputs(135)) xor (inputs(10));
    layer0_outputs(769) <= not((inputs(160)) or (inputs(103)));
    layer0_outputs(770) <= not((inputs(194)) xor (inputs(54)));
    layer0_outputs(771) <= not((inputs(101)) or (inputs(235)));
    layer0_outputs(772) <= (inputs(142)) or (inputs(49));
    layer0_outputs(773) <= (inputs(73)) xor (inputs(237));
    layer0_outputs(774) <= not(inputs(255)) or (inputs(123));
    layer0_outputs(775) <= inputs(113);
    layer0_outputs(776) <= '1';
    layer0_outputs(777) <= not(inputs(133)) or (inputs(97));
    layer0_outputs(778) <= not(inputs(41)) or (inputs(113));
    layer0_outputs(779) <= not(inputs(39));
    layer0_outputs(780) <= (inputs(21)) or (inputs(124));
    layer0_outputs(781) <= not(inputs(251)) or (inputs(130));
    layer0_outputs(782) <= (inputs(66)) xor (inputs(208));
    layer0_outputs(783) <= (inputs(179)) and not (inputs(202));
    layer0_outputs(784) <= inputs(34);
    layer0_outputs(785) <= inputs(89);
    layer0_outputs(786) <= not((inputs(108)) and (inputs(228)));
    layer0_outputs(787) <= not((inputs(191)) xor (inputs(156)));
    layer0_outputs(788) <= inputs(55);
    layer0_outputs(789) <= (inputs(160)) or (inputs(141));
    layer0_outputs(790) <= inputs(183);
    layer0_outputs(791) <= inputs(191);
    layer0_outputs(792) <= not(inputs(105));
    layer0_outputs(793) <= not(inputs(223));
    layer0_outputs(794) <= '0';
    layer0_outputs(795) <= (inputs(100)) and not (inputs(63));
    layer0_outputs(796) <= not((inputs(13)) and (inputs(66)));
    layer0_outputs(797) <= (inputs(211)) and not (inputs(95));
    layer0_outputs(798) <= inputs(69);
    layer0_outputs(799) <= (inputs(46)) xor (inputs(119));
    layer0_outputs(800) <= (inputs(60)) xor (inputs(44));
    layer0_outputs(801) <= not(inputs(112));
    layer0_outputs(802) <= not(inputs(66));
    layer0_outputs(803) <= not(inputs(70));
    layer0_outputs(804) <= '0';
    layer0_outputs(805) <= inputs(62);
    layer0_outputs(806) <= not(inputs(114)) or (inputs(11));
    layer0_outputs(807) <= inputs(97);
    layer0_outputs(808) <= (inputs(65)) or (inputs(70));
    layer0_outputs(809) <= not((inputs(211)) or (inputs(158)));
    layer0_outputs(810) <= not((inputs(80)) xor (inputs(39)));
    layer0_outputs(811) <= not(inputs(177));
    layer0_outputs(812) <= (inputs(37)) and (inputs(31));
    layer0_outputs(813) <= not(inputs(233));
    layer0_outputs(814) <= (inputs(50)) or (inputs(145));
    layer0_outputs(815) <= inputs(81);
    layer0_outputs(816) <= not((inputs(99)) xor (inputs(198)));
    layer0_outputs(817) <= not((inputs(41)) or (inputs(152)));
    layer0_outputs(818) <= not(inputs(102));
    layer0_outputs(819) <= not((inputs(217)) or (inputs(109)));
    layer0_outputs(820) <= (inputs(28)) xor (inputs(235));
    layer0_outputs(821) <= '1';
    layer0_outputs(822) <= inputs(150);
    layer0_outputs(823) <= not((inputs(114)) xor (inputs(97)));
    layer0_outputs(824) <= '1';
    layer0_outputs(825) <= (inputs(17)) and not (inputs(138));
    layer0_outputs(826) <= inputs(102);
    layer0_outputs(827) <= (inputs(56)) xor (inputs(127));
    layer0_outputs(828) <= not((inputs(105)) xor (inputs(219)));
    layer0_outputs(829) <= inputs(239);
    layer0_outputs(830) <= (inputs(18)) and not (inputs(211));
    layer0_outputs(831) <= not(inputs(127)) or (inputs(3));
    layer0_outputs(832) <= (inputs(67)) and not (inputs(96));
    layer0_outputs(833) <= (inputs(109)) or (inputs(38));
    layer0_outputs(834) <= (inputs(175)) and not (inputs(248));
    layer0_outputs(835) <= (inputs(92)) and not (inputs(219));
    layer0_outputs(836) <= not(inputs(240)) or (inputs(78));
    layer0_outputs(837) <= inputs(216);
    layer0_outputs(838) <= (inputs(199)) xor (inputs(207));
    layer0_outputs(839) <= (inputs(176)) and not (inputs(130));
    layer0_outputs(840) <= (inputs(204)) xor (inputs(172));
    layer0_outputs(841) <= not(inputs(61)) or (inputs(245));
    layer0_outputs(842) <= not((inputs(108)) or (inputs(56)));
    layer0_outputs(843) <= not((inputs(220)) xor (inputs(157)));
    layer0_outputs(844) <= (inputs(239)) or (inputs(82));
    layer0_outputs(845) <= (inputs(157)) and not (inputs(80));
    layer0_outputs(846) <= not((inputs(52)) and (inputs(141)));
    layer0_outputs(847) <= (inputs(108)) xor (inputs(225));
    layer0_outputs(848) <= (inputs(209)) or (inputs(77));
    layer0_outputs(849) <= not(inputs(55)) or (inputs(239));
    layer0_outputs(850) <= not((inputs(70)) or (inputs(174)));
    layer0_outputs(851) <= (inputs(137)) and not (inputs(213));
    layer0_outputs(852) <= not(inputs(164));
    layer0_outputs(853) <= inputs(34);
    layer0_outputs(854) <= (inputs(72)) or (inputs(211));
    layer0_outputs(855) <= (inputs(137)) and not (inputs(21));
    layer0_outputs(856) <= not(inputs(89));
    layer0_outputs(857) <= not(inputs(41)) or (inputs(171));
    layer0_outputs(858) <= not(inputs(154));
    layer0_outputs(859) <= (inputs(70)) xor (inputs(128));
    layer0_outputs(860) <= not(inputs(163));
    layer0_outputs(861) <= (inputs(232)) xor (inputs(193));
    layer0_outputs(862) <= (inputs(149)) and not (inputs(245));
    layer0_outputs(863) <= not((inputs(98)) xor (inputs(2)));
    layer0_outputs(864) <= '1';
    layer0_outputs(865) <= (inputs(177)) and not (inputs(183));
    layer0_outputs(866) <= (inputs(232)) and not (inputs(218));
    layer0_outputs(867) <= (inputs(216)) or (inputs(211));
    layer0_outputs(868) <= not((inputs(169)) xor (inputs(202)));
    layer0_outputs(869) <= inputs(47);
    layer0_outputs(870) <= not((inputs(118)) xor (inputs(186)));
    layer0_outputs(871) <= not(inputs(2));
    layer0_outputs(872) <= (inputs(228)) xor (inputs(215));
    layer0_outputs(873) <= not(inputs(245)) or (inputs(226));
    layer0_outputs(874) <= not((inputs(192)) and (inputs(244)));
    layer0_outputs(875) <= inputs(83);
    layer0_outputs(876) <= not(inputs(56));
    layer0_outputs(877) <= not(inputs(25)) or (inputs(42));
    layer0_outputs(878) <= not((inputs(129)) or (inputs(70)));
    layer0_outputs(879) <= not((inputs(75)) xor (inputs(209)));
    layer0_outputs(880) <= not(inputs(188)) or (inputs(142));
    layer0_outputs(881) <= (inputs(162)) or (inputs(173));
    layer0_outputs(882) <= not(inputs(91));
    layer0_outputs(883) <= (inputs(225)) and not (inputs(211));
    layer0_outputs(884) <= not((inputs(126)) or (inputs(153)));
    layer0_outputs(885) <= not((inputs(42)) or (inputs(186)));
    layer0_outputs(886) <= not((inputs(25)) xor (inputs(21)));
    layer0_outputs(887) <= not(inputs(4));
    layer0_outputs(888) <= not(inputs(140)) or (inputs(203));
    layer0_outputs(889) <= (inputs(5)) or (inputs(20));
    layer0_outputs(890) <= not((inputs(233)) xor (inputs(198)));
    layer0_outputs(891) <= (inputs(206)) xor (inputs(81));
    layer0_outputs(892) <= not((inputs(17)) xor (inputs(73)));
    layer0_outputs(893) <= not((inputs(193)) or (inputs(170)));
    layer0_outputs(894) <= (inputs(229)) or (inputs(53));
    layer0_outputs(895) <= not(inputs(101));
    layer0_outputs(896) <= inputs(136);
    layer0_outputs(897) <= (inputs(58)) and not (inputs(229));
    layer0_outputs(898) <= (inputs(176)) or (inputs(44));
    layer0_outputs(899) <= (inputs(10)) or (inputs(71));
    layer0_outputs(900) <= (inputs(53)) and not (inputs(210));
    layer0_outputs(901) <= not(inputs(19));
    layer0_outputs(902) <= not(inputs(103));
    layer0_outputs(903) <= not(inputs(120)) or (inputs(194));
    layer0_outputs(904) <= (inputs(101)) and not (inputs(230));
    layer0_outputs(905) <= not(inputs(174)) or (inputs(47));
    layer0_outputs(906) <= (inputs(0)) and (inputs(3));
    layer0_outputs(907) <= not(inputs(179)) or (inputs(128));
    layer0_outputs(908) <= not((inputs(43)) or (inputs(157)));
    layer0_outputs(909) <= '1';
    layer0_outputs(910) <= not((inputs(68)) xor (inputs(79)));
    layer0_outputs(911) <= '0';
    layer0_outputs(912) <= not(inputs(198)) or (inputs(131));
    layer0_outputs(913) <= not(inputs(209)) or (inputs(249));
    layer0_outputs(914) <= not(inputs(171)) or (inputs(177));
    layer0_outputs(915) <= (inputs(174)) and not (inputs(248));
    layer0_outputs(916) <= (inputs(72)) or (inputs(247));
    layer0_outputs(917) <= not(inputs(147));
    layer0_outputs(918) <= not((inputs(191)) or (inputs(106)));
    layer0_outputs(919) <= (inputs(181)) and not (inputs(148));
    layer0_outputs(920) <= not(inputs(140));
    layer0_outputs(921) <= (inputs(61)) or (inputs(139));
    layer0_outputs(922) <= (inputs(56)) or (inputs(57));
    layer0_outputs(923) <= '1';
    layer0_outputs(924) <= (inputs(226)) and not (inputs(155));
    layer0_outputs(925) <= (inputs(112)) or (inputs(110));
    layer0_outputs(926) <= '1';
    layer0_outputs(927) <= '1';
    layer0_outputs(928) <= not((inputs(221)) xor (inputs(88)));
    layer0_outputs(929) <= not((inputs(139)) or (inputs(239)));
    layer0_outputs(930) <= (inputs(222)) or (inputs(26));
    layer0_outputs(931) <= (inputs(60)) or (inputs(156));
    layer0_outputs(932) <= '0';
    layer0_outputs(933) <= not((inputs(79)) or (inputs(64)));
    layer0_outputs(934) <= not(inputs(149)) or (inputs(123));
    layer0_outputs(935) <= not(inputs(167));
    layer0_outputs(936) <= inputs(88);
    layer0_outputs(937) <= (inputs(166)) and not (inputs(246));
    layer0_outputs(938) <= not(inputs(166));
    layer0_outputs(939) <= not((inputs(105)) xor (inputs(107)));
    layer0_outputs(940) <= (inputs(27)) xor (inputs(228));
    layer0_outputs(941) <= inputs(105);
    layer0_outputs(942) <= not(inputs(234)) or (inputs(145));
    layer0_outputs(943) <= inputs(70);
    layer0_outputs(944) <= not((inputs(2)) and (inputs(61)));
    layer0_outputs(945) <= (inputs(23)) xor (inputs(99));
    layer0_outputs(946) <= inputs(81);
    layer0_outputs(947) <= (inputs(113)) and (inputs(62));
    layer0_outputs(948) <= '0';
    layer0_outputs(949) <= not(inputs(132)) or (inputs(73));
    layer0_outputs(950) <= not((inputs(77)) or (inputs(65)));
    layer0_outputs(951) <= not((inputs(14)) xor (inputs(70)));
    layer0_outputs(952) <= inputs(236);
    layer0_outputs(953) <= inputs(91);
    layer0_outputs(954) <= (inputs(64)) and not (inputs(197));
    layer0_outputs(955) <= inputs(119);
    layer0_outputs(956) <= (inputs(127)) xor (inputs(196));
    layer0_outputs(957) <= not(inputs(73));
    layer0_outputs(958) <= (inputs(76)) xor (inputs(192));
    layer0_outputs(959) <= inputs(55);
    layer0_outputs(960) <= inputs(152);
    layer0_outputs(961) <= not((inputs(159)) xor (inputs(254)));
    layer0_outputs(962) <= inputs(86);
    layer0_outputs(963) <= not((inputs(110)) xor (inputs(192)));
    layer0_outputs(964) <= not((inputs(87)) or (inputs(206)));
    layer0_outputs(965) <= not((inputs(44)) xor (inputs(53)));
    layer0_outputs(966) <= not((inputs(112)) xor (inputs(178)));
    layer0_outputs(967) <= not((inputs(98)) xor (inputs(38)));
    layer0_outputs(968) <= (inputs(43)) and not (inputs(70));
    layer0_outputs(969) <= (inputs(2)) and not (inputs(112));
    layer0_outputs(970) <= not((inputs(207)) or (inputs(4)));
    layer0_outputs(971) <= not(inputs(29));
    layer0_outputs(972) <= not(inputs(206)) or (inputs(32));
    layer0_outputs(973) <= not((inputs(129)) xor (inputs(84)));
    layer0_outputs(974) <= '0';
    layer0_outputs(975) <= not(inputs(172)) or (inputs(107));
    layer0_outputs(976) <= inputs(205);
    layer0_outputs(977) <= (inputs(65)) or (inputs(202));
    layer0_outputs(978) <= (inputs(30)) or (inputs(125));
    layer0_outputs(979) <= (inputs(233)) and not (inputs(226));
    layer0_outputs(980) <= not(inputs(71));
    layer0_outputs(981) <= (inputs(48)) and not (inputs(173));
    layer0_outputs(982) <= not(inputs(88)) or (inputs(242));
    layer0_outputs(983) <= not(inputs(108));
    layer0_outputs(984) <= not(inputs(103));
    layer0_outputs(985) <= not((inputs(192)) xor (inputs(236)));
    layer0_outputs(986) <= not(inputs(72));
    layer0_outputs(987) <= (inputs(214)) xor (inputs(27));
    layer0_outputs(988) <= inputs(88);
    layer0_outputs(989) <= inputs(74);
    layer0_outputs(990) <= not((inputs(162)) or (inputs(136)));
    layer0_outputs(991) <= not(inputs(15));
    layer0_outputs(992) <= (inputs(128)) and not (inputs(34));
    layer0_outputs(993) <= (inputs(11)) xor (inputs(218));
    layer0_outputs(994) <= (inputs(82)) or (inputs(195));
    layer0_outputs(995) <= inputs(167);
    layer0_outputs(996) <= not((inputs(244)) xor (inputs(102)));
    layer0_outputs(997) <= not((inputs(128)) or (inputs(136)));
    layer0_outputs(998) <= not(inputs(120)) or (inputs(176));
    layer0_outputs(999) <= not(inputs(184)) or (inputs(193));
    layer0_outputs(1000) <= not(inputs(108)) or (inputs(37));
    layer0_outputs(1001) <= not(inputs(41)) or (inputs(67));
    layer0_outputs(1002) <= not(inputs(102));
    layer0_outputs(1003) <= (inputs(10)) or (inputs(100));
    layer0_outputs(1004) <= (inputs(39)) or (inputs(231));
    layer0_outputs(1005) <= inputs(132);
    layer0_outputs(1006) <= not(inputs(59));
    layer0_outputs(1007) <= inputs(100);
    layer0_outputs(1008) <= not((inputs(217)) or (inputs(60)));
    layer0_outputs(1009) <= (inputs(183)) and not (inputs(1));
    layer0_outputs(1010) <= (inputs(11)) or (inputs(75));
    layer0_outputs(1011) <= '0';
    layer0_outputs(1012) <= (inputs(196)) and not (inputs(115));
    layer0_outputs(1013) <= (inputs(162)) xor (inputs(137));
    layer0_outputs(1014) <= inputs(150);
    layer0_outputs(1015) <= (inputs(121)) or (inputs(26));
    layer0_outputs(1016) <= inputs(84);
    layer0_outputs(1017) <= not(inputs(116)) or (inputs(250));
    layer0_outputs(1018) <= (inputs(196)) and not (inputs(174));
    layer0_outputs(1019) <= not((inputs(194)) or (inputs(230)));
    layer0_outputs(1020) <= (inputs(71)) xor (inputs(100));
    layer0_outputs(1021) <= inputs(86);
    layer0_outputs(1022) <= (inputs(28)) and not (inputs(255));
    layer0_outputs(1023) <= not(inputs(142)) or (inputs(122));
    layer0_outputs(1024) <= not(inputs(144)) or (inputs(213));
    layer0_outputs(1025) <= (inputs(205)) xor (inputs(75));
    layer0_outputs(1026) <= (inputs(83)) xor (inputs(170));
    layer0_outputs(1027) <= (inputs(184)) or (inputs(179));
    layer0_outputs(1028) <= (inputs(155)) or (inputs(44));
    layer0_outputs(1029) <= not((inputs(2)) xor (inputs(164)));
    layer0_outputs(1030) <= (inputs(104)) or (inputs(184));
    layer0_outputs(1031) <= not(inputs(186));
    layer0_outputs(1032) <= (inputs(76)) and not (inputs(251));
    layer0_outputs(1033) <= (inputs(227)) and (inputs(35));
    layer0_outputs(1034) <= (inputs(81)) xor (inputs(254));
    layer0_outputs(1035) <= not((inputs(168)) or (inputs(3)));
    layer0_outputs(1036) <= (inputs(104)) and not (inputs(229));
    layer0_outputs(1037) <= not(inputs(130));
    layer0_outputs(1038) <= not((inputs(142)) xor (inputs(33)));
    layer0_outputs(1039) <= (inputs(140)) and not (inputs(3));
    layer0_outputs(1040) <= not(inputs(40)) or (inputs(174));
    layer0_outputs(1041) <= not(inputs(223));
    layer0_outputs(1042) <= (inputs(25)) and (inputs(145));
    layer0_outputs(1043) <= (inputs(114)) or (inputs(19));
    layer0_outputs(1044) <= (inputs(233)) and not (inputs(46));
    layer0_outputs(1045) <= (inputs(135)) or (inputs(233));
    layer0_outputs(1046) <= (inputs(255)) xor (inputs(11));
    layer0_outputs(1047) <= not((inputs(239)) xor (inputs(150)));
    layer0_outputs(1048) <= not(inputs(10));
    layer0_outputs(1049) <= not(inputs(133)) or (inputs(207));
    layer0_outputs(1050) <= not(inputs(30));
    layer0_outputs(1051) <= not((inputs(41)) or (inputs(36)));
    layer0_outputs(1052) <= (inputs(159)) and not (inputs(126));
    layer0_outputs(1053) <= not((inputs(179)) or (inputs(197)));
    layer0_outputs(1054) <= (inputs(36)) or (inputs(162));
    layer0_outputs(1055) <= not(inputs(164));
    layer0_outputs(1056) <= (inputs(45)) xor (inputs(81));
    layer0_outputs(1057) <= (inputs(24)) and (inputs(174));
    layer0_outputs(1058) <= (inputs(181)) and not (inputs(44));
    layer0_outputs(1059) <= not((inputs(202)) or (inputs(62)));
    layer0_outputs(1060) <= not(inputs(124)) or (inputs(219));
    layer0_outputs(1061) <= not(inputs(27));
    layer0_outputs(1062) <= not(inputs(141));
    layer0_outputs(1063) <= not(inputs(55)) or (inputs(79));
    layer0_outputs(1064) <= inputs(43);
    layer0_outputs(1065) <= '0';
    layer0_outputs(1066) <= (inputs(174)) xor (inputs(100));
    layer0_outputs(1067) <= not(inputs(135)) or (inputs(89));
    layer0_outputs(1068) <= (inputs(180)) and not (inputs(222));
    layer0_outputs(1069) <= (inputs(67)) or (inputs(151));
    layer0_outputs(1070) <= (inputs(226)) and not (inputs(113));
    layer0_outputs(1071) <= not(inputs(62)) or (inputs(158));
    layer0_outputs(1072) <= not((inputs(238)) or (inputs(35)));
    layer0_outputs(1073) <= not(inputs(21));
    layer0_outputs(1074) <= '1';
    layer0_outputs(1075) <= not(inputs(148)) or (inputs(28));
    layer0_outputs(1076) <= (inputs(66)) or (inputs(215));
    layer0_outputs(1077) <= not(inputs(76));
    layer0_outputs(1078) <= (inputs(63)) or (inputs(68));
    layer0_outputs(1079) <= (inputs(154)) and not (inputs(78));
    layer0_outputs(1080) <= not(inputs(32));
    layer0_outputs(1081) <= (inputs(49)) or (inputs(78));
    layer0_outputs(1082) <= (inputs(89)) or (inputs(249));
    layer0_outputs(1083) <= (inputs(43)) xor (inputs(32));
    layer0_outputs(1084) <= not((inputs(251)) or (inputs(224)));
    layer0_outputs(1085) <= not(inputs(114)) or (inputs(62));
    layer0_outputs(1086) <= not(inputs(134)) or (inputs(166));
    layer0_outputs(1087) <= not((inputs(149)) or (inputs(93)));
    layer0_outputs(1088) <= '1';
    layer0_outputs(1089) <= (inputs(170)) or (inputs(85));
    layer0_outputs(1090) <= not((inputs(237)) xor (inputs(36)));
    layer0_outputs(1091) <= (inputs(125)) and not (inputs(83));
    layer0_outputs(1092) <= not(inputs(46));
    layer0_outputs(1093) <= not(inputs(91));
    layer0_outputs(1094) <= '0';
    layer0_outputs(1095) <= (inputs(62)) and not (inputs(193));
    layer0_outputs(1096) <= not((inputs(61)) xor (inputs(187)));
    layer0_outputs(1097) <= (inputs(135)) and (inputs(59));
    layer0_outputs(1098) <= (inputs(103)) or (inputs(69));
    layer0_outputs(1099) <= (inputs(89)) and not (inputs(23));
    layer0_outputs(1100) <= not(inputs(163)) or (inputs(165));
    layer0_outputs(1101) <= not(inputs(132)) or (inputs(63));
    layer0_outputs(1102) <= (inputs(78)) xor (inputs(128));
    layer0_outputs(1103) <= inputs(133);
    layer0_outputs(1104) <= (inputs(186)) or (inputs(190));
    layer0_outputs(1105) <= not((inputs(11)) xor (inputs(5)));
    layer0_outputs(1106) <= not((inputs(93)) and (inputs(12)));
    layer0_outputs(1107) <= not((inputs(66)) and (inputs(249)));
    layer0_outputs(1108) <= '1';
    layer0_outputs(1109) <= not((inputs(223)) and (inputs(178)));
    layer0_outputs(1110) <= not(inputs(120));
    layer0_outputs(1111) <= (inputs(205)) or (inputs(166));
    layer0_outputs(1112) <= inputs(173);
    layer0_outputs(1113) <= (inputs(191)) and not (inputs(236));
    layer0_outputs(1114) <= not(inputs(22)) or (inputs(147));
    layer0_outputs(1115) <= (inputs(101)) or (inputs(78));
    layer0_outputs(1116) <= (inputs(198)) xor (inputs(218));
    layer0_outputs(1117) <= not(inputs(103));
    layer0_outputs(1118) <= '1';
    layer0_outputs(1119) <= (inputs(221)) and (inputs(82));
    layer0_outputs(1120) <= (inputs(6)) or (inputs(64));
    layer0_outputs(1121) <= not((inputs(44)) or (inputs(118)));
    layer0_outputs(1122) <= '1';
    layer0_outputs(1123) <= (inputs(4)) and (inputs(184));
    layer0_outputs(1124) <= not((inputs(114)) xor (inputs(116)));
    layer0_outputs(1125) <= (inputs(47)) and (inputs(38));
    layer0_outputs(1126) <= not(inputs(61));
    layer0_outputs(1127) <= not((inputs(139)) or (inputs(241)));
    layer0_outputs(1128) <= (inputs(149)) or (inputs(247));
    layer0_outputs(1129) <= (inputs(18)) or (inputs(219));
    layer0_outputs(1130) <= (inputs(195)) or (inputs(232));
    layer0_outputs(1131) <= not(inputs(182)) or (inputs(243));
    layer0_outputs(1132) <= not(inputs(124));
    layer0_outputs(1133) <= not(inputs(217)) or (inputs(32));
    layer0_outputs(1134) <= not((inputs(157)) or (inputs(37)));
    layer0_outputs(1135) <= inputs(105);
    layer0_outputs(1136) <= not((inputs(150)) xor (inputs(226)));
    layer0_outputs(1137) <= '1';
    layer0_outputs(1138) <= inputs(197);
    layer0_outputs(1139) <= not((inputs(32)) xor (inputs(139)));
    layer0_outputs(1140) <= inputs(57);
    layer0_outputs(1141) <= inputs(47);
    layer0_outputs(1142) <= not(inputs(56)) or (inputs(220));
    layer0_outputs(1143) <= not(inputs(90));
    layer0_outputs(1144) <= (inputs(175)) and (inputs(193));
    layer0_outputs(1145) <= inputs(26);
    layer0_outputs(1146) <= not((inputs(77)) and (inputs(12)));
    layer0_outputs(1147) <= not(inputs(156));
    layer0_outputs(1148) <= not(inputs(113));
    layer0_outputs(1149) <= not(inputs(142)) or (inputs(52));
    layer0_outputs(1150) <= (inputs(154)) and not (inputs(4));
    layer0_outputs(1151) <= not(inputs(40));
    layer0_outputs(1152) <= not(inputs(231));
    layer0_outputs(1153) <= not((inputs(20)) and (inputs(59)));
    layer0_outputs(1154) <= (inputs(249)) or (inputs(234));
    layer0_outputs(1155) <= not(inputs(242)) or (inputs(66));
    layer0_outputs(1156) <= not(inputs(64));
    layer0_outputs(1157) <= (inputs(172)) or (inputs(182));
    layer0_outputs(1158) <= not(inputs(152)) or (inputs(223));
    layer0_outputs(1159) <= inputs(133);
    layer0_outputs(1160) <= not((inputs(75)) or (inputs(5)));
    layer0_outputs(1161) <= (inputs(118)) and not (inputs(209));
    layer0_outputs(1162) <= (inputs(219)) xor (inputs(186));
    layer0_outputs(1163) <= (inputs(86)) and not (inputs(241));
    layer0_outputs(1164) <= not(inputs(201));
    layer0_outputs(1165) <= not((inputs(111)) xor (inputs(153)));
    layer0_outputs(1166) <= (inputs(196)) or (inputs(38));
    layer0_outputs(1167) <= not((inputs(135)) or (inputs(111)));
    layer0_outputs(1168) <= (inputs(98)) xor (inputs(170));
    layer0_outputs(1169) <= not(inputs(122));
    layer0_outputs(1170) <= (inputs(0)) xor (inputs(173));
    layer0_outputs(1171) <= '1';
    layer0_outputs(1172) <= not((inputs(117)) or (inputs(107)));
    layer0_outputs(1173) <= (inputs(138)) and not (inputs(159));
    layer0_outputs(1174) <= (inputs(34)) and not (inputs(115));
    layer0_outputs(1175) <= (inputs(188)) and not (inputs(132));
    layer0_outputs(1176) <= not(inputs(71)) or (inputs(8));
    layer0_outputs(1177) <= inputs(247);
    layer0_outputs(1178) <= not((inputs(39)) or (inputs(1)));
    layer0_outputs(1179) <= not(inputs(212)) or (inputs(194));
    layer0_outputs(1180) <= (inputs(206)) xor (inputs(148));
    layer0_outputs(1181) <= not(inputs(227)) or (inputs(221));
    layer0_outputs(1182) <= (inputs(18)) and not (inputs(93));
    layer0_outputs(1183) <= (inputs(201)) xor (inputs(127));
    layer0_outputs(1184) <= (inputs(36)) xor (inputs(56));
    layer0_outputs(1185) <= not((inputs(5)) xor (inputs(9)));
    layer0_outputs(1186) <= (inputs(217)) and not (inputs(247));
    layer0_outputs(1187) <= (inputs(249)) or (inputs(190));
    layer0_outputs(1188) <= (inputs(20)) xor (inputs(69));
    layer0_outputs(1189) <= (inputs(117)) or (inputs(119));
    layer0_outputs(1190) <= inputs(38);
    layer0_outputs(1191) <= not((inputs(146)) or (inputs(122)));
    layer0_outputs(1192) <= (inputs(10)) xor (inputs(43));
    layer0_outputs(1193) <= not(inputs(99));
    layer0_outputs(1194) <= (inputs(222)) or (inputs(56));
    layer0_outputs(1195) <= not((inputs(58)) or (inputs(148)));
    layer0_outputs(1196) <= not((inputs(75)) and (inputs(193)));
    layer0_outputs(1197) <= not((inputs(18)) or (inputs(168)));
    layer0_outputs(1198) <= inputs(255);
    layer0_outputs(1199) <= not(inputs(212));
    layer0_outputs(1200) <= (inputs(87)) xor (inputs(244));
    layer0_outputs(1201) <= not((inputs(224)) xor (inputs(104)));
    layer0_outputs(1202) <= '1';
    layer0_outputs(1203) <= not(inputs(149));
    layer0_outputs(1204) <= inputs(236);
    layer0_outputs(1205) <= (inputs(126)) and not (inputs(81));
    layer0_outputs(1206) <= (inputs(32)) xor (inputs(237));
    layer0_outputs(1207) <= not((inputs(120)) xor (inputs(141)));
    layer0_outputs(1208) <= inputs(193);
    layer0_outputs(1209) <= (inputs(150)) and not (inputs(243));
    layer0_outputs(1210) <= not(inputs(41));
    layer0_outputs(1211) <= (inputs(188)) or (inputs(155));
    layer0_outputs(1212) <= (inputs(132)) or (inputs(142));
    layer0_outputs(1213) <= not((inputs(59)) xor (inputs(104)));
    layer0_outputs(1214) <= not(inputs(109));
    layer0_outputs(1215) <= not(inputs(92)) or (inputs(205));
    layer0_outputs(1216) <= not(inputs(207));
    layer0_outputs(1217) <= inputs(166);
    layer0_outputs(1218) <= not(inputs(50)) or (inputs(32));
    layer0_outputs(1219) <= not(inputs(46));
    layer0_outputs(1220) <= not(inputs(37));
    layer0_outputs(1221) <= (inputs(62)) and (inputs(20));
    layer0_outputs(1222) <= not((inputs(108)) or (inputs(224)));
    layer0_outputs(1223) <= inputs(139);
    layer0_outputs(1224) <= not((inputs(2)) xor (inputs(199)));
    layer0_outputs(1225) <= not((inputs(106)) xor (inputs(148)));
    layer0_outputs(1226) <= inputs(132);
    layer0_outputs(1227) <= (inputs(105)) and (inputs(89));
    layer0_outputs(1228) <= not(inputs(28));
    layer0_outputs(1229) <= not((inputs(148)) xor (inputs(84)));
    layer0_outputs(1230) <= (inputs(122)) and not (inputs(40));
    layer0_outputs(1231) <= not((inputs(211)) or (inputs(187)));
    layer0_outputs(1232) <= not((inputs(224)) or (inputs(42)));
    layer0_outputs(1233) <= not(inputs(217));
    layer0_outputs(1234) <= not((inputs(79)) xor (inputs(121)));
    layer0_outputs(1235) <= not(inputs(107)) or (inputs(191));
    layer0_outputs(1236) <= (inputs(129)) and not (inputs(162));
    layer0_outputs(1237) <= (inputs(117)) and not (inputs(234));
    layer0_outputs(1238) <= (inputs(202)) xor (inputs(181));
    layer0_outputs(1239) <= not(inputs(152)) or (inputs(136));
    layer0_outputs(1240) <= not(inputs(73));
    layer0_outputs(1241) <= not(inputs(210));
    layer0_outputs(1242) <= (inputs(38)) or (inputs(8));
    layer0_outputs(1243) <= not(inputs(66)) or (inputs(96));
    layer0_outputs(1244) <= inputs(237);
    layer0_outputs(1245) <= not((inputs(158)) or (inputs(48)));
    layer0_outputs(1246) <= not((inputs(208)) xor (inputs(171)));
    layer0_outputs(1247) <= not((inputs(56)) xor (inputs(99)));
    layer0_outputs(1248) <= not((inputs(186)) xor (inputs(72)));
    layer0_outputs(1249) <= (inputs(104)) and not (inputs(147));
    layer0_outputs(1250) <= (inputs(1)) or (inputs(218));
    layer0_outputs(1251) <= inputs(249);
    layer0_outputs(1252) <= '0';
    layer0_outputs(1253) <= (inputs(25)) and not (inputs(20));
    layer0_outputs(1254) <= (inputs(109)) xor (inputs(176));
    layer0_outputs(1255) <= (inputs(192)) xor (inputs(42));
    layer0_outputs(1256) <= not((inputs(72)) xor (inputs(171)));
    layer0_outputs(1257) <= not(inputs(138)) or (inputs(150));
    layer0_outputs(1258) <= not((inputs(146)) or (inputs(96)));
    layer0_outputs(1259) <= (inputs(158)) and not (inputs(217));
    layer0_outputs(1260) <= not((inputs(98)) and (inputs(250)));
    layer0_outputs(1261) <= inputs(35);
    layer0_outputs(1262) <= not(inputs(135)) or (inputs(222));
    layer0_outputs(1263) <= not(inputs(11));
    layer0_outputs(1264) <= inputs(231);
    layer0_outputs(1265) <= not((inputs(184)) xor (inputs(35)));
    layer0_outputs(1266) <= inputs(136);
    layer0_outputs(1267) <= not((inputs(73)) or (inputs(14)));
    layer0_outputs(1268) <= not((inputs(206)) or (inputs(146)));
    layer0_outputs(1269) <= (inputs(158)) and not (inputs(129));
    layer0_outputs(1270) <= inputs(27);
    layer0_outputs(1271) <= not((inputs(28)) and (inputs(159)));
    layer0_outputs(1272) <= not((inputs(238)) or (inputs(51)));
    layer0_outputs(1273) <= (inputs(138)) and not (inputs(85));
    layer0_outputs(1274) <= not((inputs(190)) or (inputs(214)));
    layer0_outputs(1275) <= not(inputs(121));
    layer0_outputs(1276) <= inputs(83);
    layer0_outputs(1277) <= inputs(236);
    layer0_outputs(1278) <= not(inputs(228));
    layer0_outputs(1279) <= (inputs(49)) and (inputs(218));
    layer0_outputs(1280) <= not((inputs(105)) xor (inputs(74)));
    layer0_outputs(1281) <= not((inputs(144)) or (inputs(57)));
    layer0_outputs(1282) <= (inputs(86)) or (inputs(233));
    layer0_outputs(1283) <= not(inputs(75));
    layer0_outputs(1284) <= (inputs(20)) and not (inputs(10));
    layer0_outputs(1285) <= not(inputs(162));
    layer0_outputs(1286) <= inputs(165);
    layer0_outputs(1287) <= not(inputs(85)) or (inputs(176));
    layer0_outputs(1288) <= not(inputs(183)) or (inputs(191));
    layer0_outputs(1289) <= (inputs(222)) or (inputs(37));
    layer0_outputs(1290) <= not((inputs(90)) xor (inputs(243)));
    layer0_outputs(1291) <= not((inputs(161)) xor (inputs(103)));
    layer0_outputs(1292) <= not((inputs(97)) or (inputs(60)));
    layer0_outputs(1293) <= (inputs(167)) and not (inputs(225));
    layer0_outputs(1294) <= (inputs(244)) xor (inputs(166));
    layer0_outputs(1295) <= (inputs(180)) or (inputs(170));
    layer0_outputs(1296) <= inputs(134);
    layer0_outputs(1297) <= inputs(101);
    layer0_outputs(1298) <= inputs(223);
    layer0_outputs(1299) <= not(inputs(26)) or (inputs(223));
    layer0_outputs(1300) <= not(inputs(40)) or (inputs(205));
    layer0_outputs(1301) <= inputs(117);
    layer0_outputs(1302) <= (inputs(147)) xor (inputs(44));
    layer0_outputs(1303) <= (inputs(247)) and not (inputs(186));
    layer0_outputs(1304) <= inputs(37);
    layer0_outputs(1305) <= not(inputs(41));
    layer0_outputs(1306) <= not(inputs(154));
    layer0_outputs(1307) <= (inputs(122)) and not (inputs(40));
    layer0_outputs(1308) <= (inputs(132)) and not (inputs(172));
    layer0_outputs(1309) <= not((inputs(33)) xor (inputs(98)));
    layer0_outputs(1310) <= not(inputs(245));
    layer0_outputs(1311) <= not((inputs(211)) or (inputs(187)));
    layer0_outputs(1312) <= not((inputs(59)) or (inputs(17)));
    layer0_outputs(1313) <= not((inputs(3)) and (inputs(250)));
    layer0_outputs(1314) <= inputs(19);
    layer0_outputs(1315) <= not(inputs(149)) or (inputs(35));
    layer0_outputs(1316) <= (inputs(162)) or (inputs(170));
    layer0_outputs(1317) <= (inputs(36)) or (inputs(240));
    layer0_outputs(1318) <= inputs(136);
    layer0_outputs(1319) <= inputs(5);
    layer0_outputs(1320) <= not(inputs(79));
    layer0_outputs(1321) <= (inputs(85)) or (inputs(229));
    layer0_outputs(1322) <= not(inputs(230));
    layer0_outputs(1323) <= (inputs(106)) xor (inputs(4));
    layer0_outputs(1324) <= inputs(52);
    layer0_outputs(1325) <= inputs(189);
    layer0_outputs(1326) <= not(inputs(244));
    layer0_outputs(1327) <= not(inputs(234));
    layer0_outputs(1328) <= (inputs(254)) and not (inputs(82));
    layer0_outputs(1329) <= not(inputs(166));
    layer0_outputs(1330) <= not(inputs(214)) or (inputs(51));
    layer0_outputs(1331) <= not((inputs(123)) xor (inputs(86)));
    layer0_outputs(1332) <= not((inputs(131)) xor (inputs(210)));
    layer0_outputs(1333) <= (inputs(124)) or (inputs(141));
    layer0_outputs(1334) <= (inputs(138)) or (inputs(87));
    layer0_outputs(1335) <= not(inputs(179));
    layer0_outputs(1336) <= inputs(177);
    layer0_outputs(1337) <= (inputs(182)) or (inputs(51));
    layer0_outputs(1338) <= not((inputs(83)) or (inputs(76)));
    layer0_outputs(1339) <= (inputs(73)) and not (inputs(5));
    layer0_outputs(1340) <= (inputs(14)) and (inputs(67));
    layer0_outputs(1341) <= not((inputs(83)) or (inputs(153)));
    layer0_outputs(1342) <= inputs(149);
    layer0_outputs(1343) <= not((inputs(224)) xor (inputs(118)));
    layer0_outputs(1344) <= not(inputs(61)) or (inputs(128));
    layer0_outputs(1345) <= not((inputs(198)) and (inputs(112)));
    layer0_outputs(1346) <= not(inputs(165));
    layer0_outputs(1347) <= not(inputs(167));
    layer0_outputs(1348) <= inputs(149);
    layer0_outputs(1349) <= inputs(181);
    layer0_outputs(1350) <= (inputs(101)) and not (inputs(187));
    layer0_outputs(1351) <= (inputs(202)) and not (inputs(124));
    layer0_outputs(1352) <= '0';
    layer0_outputs(1353) <= (inputs(147)) xor (inputs(62));
    layer0_outputs(1354) <= (inputs(109)) xor (inputs(102));
    layer0_outputs(1355) <= not((inputs(54)) or (inputs(68)));
    layer0_outputs(1356) <= (inputs(204)) and not (inputs(1));
    layer0_outputs(1357) <= not(inputs(2));
    layer0_outputs(1358) <= (inputs(23)) or (inputs(113));
    layer0_outputs(1359) <= not((inputs(63)) and (inputs(237)));
    layer0_outputs(1360) <= not(inputs(27)) or (inputs(30));
    layer0_outputs(1361) <= not(inputs(85));
    layer0_outputs(1362) <= (inputs(86)) and not (inputs(117));
    layer0_outputs(1363) <= not((inputs(13)) or (inputs(200)));
    layer0_outputs(1364) <= (inputs(22)) and (inputs(229));
    layer0_outputs(1365) <= not((inputs(61)) or (inputs(95)));
    layer0_outputs(1366) <= (inputs(111)) and not (inputs(31));
    layer0_outputs(1367) <= (inputs(9)) or (inputs(238));
    layer0_outputs(1368) <= '1';
    layer0_outputs(1369) <= not(inputs(168));
    layer0_outputs(1370) <= inputs(51);
    layer0_outputs(1371) <= not(inputs(165));
    layer0_outputs(1372) <= inputs(38);
    layer0_outputs(1373) <= not(inputs(56)) or (inputs(3));
    layer0_outputs(1374) <= (inputs(188)) or (inputs(194));
    layer0_outputs(1375) <= not((inputs(41)) or (inputs(52)));
    layer0_outputs(1376) <= inputs(184);
    layer0_outputs(1377) <= (inputs(65)) and not (inputs(113));
    layer0_outputs(1378) <= '0';
    layer0_outputs(1379) <= not(inputs(78));
    layer0_outputs(1380) <= not(inputs(62)) or (inputs(81));
    layer0_outputs(1381) <= (inputs(255)) and not (inputs(197));
    layer0_outputs(1382) <= (inputs(218)) and not (inputs(134));
    layer0_outputs(1383) <= not(inputs(149));
    layer0_outputs(1384) <= inputs(41);
    layer0_outputs(1385) <= not((inputs(113)) and (inputs(253)));
    layer0_outputs(1386) <= not(inputs(137)) or (inputs(205));
    layer0_outputs(1387) <= not(inputs(155));
    layer0_outputs(1388) <= not(inputs(157));
    layer0_outputs(1389) <= (inputs(247)) or (inputs(165));
    layer0_outputs(1390) <= '1';
    layer0_outputs(1391) <= not(inputs(107)) or (inputs(173));
    layer0_outputs(1392) <= (inputs(197)) and not (inputs(109));
    layer0_outputs(1393) <= (inputs(190)) and (inputs(190));
    layer0_outputs(1394) <= (inputs(73)) xor (inputs(119));
    layer0_outputs(1395) <= not(inputs(229)) or (inputs(119));
    layer0_outputs(1396) <= not(inputs(114));
    layer0_outputs(1397) <= (inputs(10)) xor (inputs(215));
    layer0_outputs(1398) <= not((inputs(192)) or (inputs(23)));
    layer0_outputs(1399) <= (inputs(209)) or (inputs(88));
    layer0_outputs(1400) <= (inputs(43)) and not (inputs(251));
    layer0_outputs(1401) <= not((inputs(85)) and (inputs(85)));
    layer0_outputs(1402) <= not(inputs(213)) or (inputs(189));
    layer0_outputs(1403) <= not((inputs(189)) xor (inputs(96)));
    layer0_outputs(1404) <= (inputs(135)) and not (inputs(162));
    layer0_outputs(1405) <= not(inputs(149));
    layer0_outputs(1406) <= (inputs(55)) and not (inputs(30));
    layer0_outputs(1407) <= (inputs(25)) and not (inputs(210));
    layer0_outputs(1408) <= not((inputs(95)) or (inputs(27)));
    layer0_outputs(1409) <= (inputs(126)) and not (inputs(207));
    layer0_outputs(1410) <= (inputs(167)) xor (inputs(164));
    layer0_outputs(1411) <= (inputs(46)) xor (inputs(215));
    layer0_outputs(1412) <= inputs(56);
    layer0_outputs(1413) <= not(inputs(59));
    layer0_outputs(1414) <= '1';
    layer0_outputs(1415) <= not(inputs(215)) or (inputs(204));
    layer0_outputs(1416) <= not(inputs(34)) or (inputs(241));
    layer0_outputs(1417) <= inputs(103);
    layer0_outputs(1418) <= not(inputs(185));
    layer0_outputs(1419) <= '1';
    layer0_outputs(1420) <= not(inputs(105)) or (inputs(156));
    layer0_outputs(1421) <= (inputs(0)) and not (inputs(246));
    layer0_outputs(1422) <= '1';
    layer0_outputs(1423) <= not((inputs(29)) xor (inputs(100)));
    layer0_outputs(1424) <= (inputs(140)) or (inputs(208));
    layer0_outputs(1425) <= not(inputs(92));
    layer0_outputs(1426) <= not((inputs(175)) xor (inputs(219)));
    layer0_outputs(1427) <= not((inputs(76)) or (inputs(74)));
    layer0_outputs(1428) <= not(inputs(107));
    layer0_outputs(1429) <= not(inputs(135));
    layer0_outputs(1430) <= not(inputs(7));
    layer0_outputs(1431) <= (inputs(154)) or (inputs(5));
    layer0_outputs(1432) <= (inputs(43)) and not (inputs(177));
    layer0_outputs(1433) <= inputs(203);
    layer0_outputs(1434) <= (inputs(224)) xor (inputs(227));
    layer0_outputs(1435) <= (inputs(32)) xor (inputs(124));
    layer0_outputs(1436) <= not((inputs(168)) or (inputs(27)));
    layer0_outputs(1437) <= not((inputs(60)) xor (inputs(137)));
    layer0_outputs(1438) <= not(inputs(3));
    layer0_outputs(1439) <= (inputs(84)) or (inputs(20));
    layer0_outputs(1440) <= inputs(120);
    layer0_outputs(1441) <= (inputs(56)) xor (inputs(38));
    layer0_outputs(1442) <= inputs(154);
    layer0_outputs(1443) <= not((inputs(186)) or (inputs(186)));
    layer0_outputs(1444) <= (inputs(117)) and not (inputs(164));
    layer0_outputs(1445) <= (inputs(59)) or (inputs(139));
    layer0_outputs(1446) <= inputs(254);
    layer0_outputs(1447) <= (inputs(184)) or (inputs(192));
    layer0_outputs(1448) <= (inputs(91)) and not (inputs(247));
    layer0_outputs(1449) <= (inputs(211)) or (inputs(76));
    layer0_outputs(1450) <= (inputs(87)) and not (inputs(47));
    layer0_outputs(1451) <= (inputs(22)) and not (inputs(192));
    layer0_outputs(1452) <= (inputs(28)) and not (inputs(192));
    layer0_outputs(1453) <= '0';
    layer0_outputs(1454) <= (inputs(36)) and (inputs(224));
    layer0_outputs(1455) <= not(inputs(56)) or (inputs(80));
    layer0_outputs(1456) <= not(inputs(39)) or (inputs(82));
    layer0_outputs(1457) <= not((inputs(51)) and (inputs(65)));
    layer0_outputs(1458) <= not((inputs(243)) xor (inputs(191)));
    layer0_outputs(1459) <= inputs(190);
    layer0_outputs(1460) <= '1';
    layer0_outputs(1461) <= not((inputs(22)) or (inputs(229)));
    layer0_outputs(1462) <= (inputs(239)) xor (inputs(48));
    layer0_outputs(1463) <= not((inputs(173)) or (inputs(60)));
    layer0_outputs(1464) <= not((inputs(194)) or (inputs(132)));
    layer0_outputs(1465) <= not(inputs(167)) or (inputs(111));
    layer0_outputs(1466) <= '0';
    layer0_outputs(1467) <= (inputs(156)) xor (inputs(21));
    layer0_outputs(1468) <= '1';
    layer0_outputs(1469) <= inputs(120);
    layer0_outputs(1470) <= '1';
    layer0_outputs(1471) <= inputs(184);
    layer0_outputs(1472) <= (inputs(139)) xor (inputs(229));
    layer0_outputs(1473) <= (inputs(112)) xor (inputs(227));
    layer0_outputs(1474) <= inputs(115);
    layer0_outputs(1475) <= (inputs(80)) and (inputs(212));
    layer0_outputs(1476) <= not((inputs(252)) and (inputs(246)));
    layer0_outputs(1477) <= (inputs(85)) and not (inputs(17));
    layer0_outputs(1478) <= (inputs(68)) or (inputs(162));
    layer0_outputs(1479) <= not(inputs(181));
    layer0_outputs(1480) <= not(inputs(172));
    layer0_outputs(1481) <= inputs(210);
    layer0_outputs(1482) <= (inputs(69)) and not (inputs(66));
    layer0_outputs(1483) <= (inputs(220)) and not (inputs(92));
    layer0_outputs(1484) <= (inputs(210)) and not (inputs(24));
    layer0_outputs(1485) <= not((inputs(131)) or (inputs(227)));
    layer0_outputs(1486) <= not((inputs(192)) or (inputs(201)));
    layer0_outputs(1487) <= not(inputs(37));
    layer0_outputs(1488) <= not((inputs(172)) or (inputs(20)));
    layer0_outputs(1489) <= inputs(99);
    layer0_outputs(1490) <= (inputs(24)) or (inputs(156));
    layer0_outputs(1491) <= '0';
    layer0_outputs(1492) <= not((inputs(167)) or (inputs(42)));
    layer0_outputs(1493) <= (inputs(236)) and (inputs(11));
    layer0_outputs(1494) <= not(inputs(200));
    layer0_outputs(1495) <= (inputs(194)) and not (inputs(110));
    layer0_outputs(1496) <= not(inputs(179));
    layer0_outputs(1497) <= inputs(41);
    layer0_outputs(1498) <= not((inputs(232)) xor (inputs(239)));
    layer0_outputs(1499) <= not((inputs(143)) xor (inputs(217)));
    layer0_outputs(1500) <= not(inputs(35)) or (inputs(22));
    layer0_outputs(1501) <= not((inputs(113)) or (inputs(172)));
    layer0_outputs(1502) <= not((inputs(54)) or (inputs(143)));
    layer0_outputs(1503) <= '0';
    layer0_outputs(1504) <= not((inputs(179)) or (inputs(241)));
    layer0_outputs(1505) <= (inputs(59)) xor (inputs(163));
    layer0_outputs(1506) <= (inputs(183)) and not (inputs(9));
    layer0_outputs(1507) <= not((inputs(50)) xor (inputs(194)));
    layer0_outputs(1508) <= not(inputs(11)) or (inputs(155));
    layer0_outputs(1509) <= not(inputs(234));
    layer0_outputs(1510) <= not((inputs(11)) and (inputs(174)));
    layer0_outputs(1511) <= not(inputs(175));
    layer0_outputs(1512) <= (inputs(209)) and (inputs(191));
    layer0_outputs(1513) <= not(inputs(146)) or (inputs(94));
    layer0_outputs(1514) <= not((inputs(131)) xor (inputs(155)));
    layer0_outputs(1515) <= not(inputs(210)) or (inputs(115));
    layer0_outputs(1516) <= not(inputs(151)) or (inputs(132));
    layer0_outputs(1517) <= (inputs(190)) xor (inputs(128));
    layer0_outputs(1518) <= not(inputs(241));
    layer0_outputs(1519) <= (inputs(208)) or (inputs(127));
    layer0_outputs(1520) <= not(inputs(163)) or (inputs(102));
    layer0_outputs(1521) <= not(inputs(152)) or (inputs(32));
    layer0_outputs(1522) <= not((inputs(47)) xor (inputs(115)));
    layer0_outputs(1523) <= not(inputs(207));
    layer0_outputs(1524) <= inputs(151);
    layer0_outputs(1525) <= not((inputs(104)) xor (inputs(239)));
    layer0_outputs(1526) <= (inputs(155)) xor (inputs(62));
    layer0_outputs(1527) <= (inputs(55)) or (inputs(190));
    layer0_outputs(1528) <= '1';
    layer0_outputs(1529) <= (inputs(104)) xor (inputs(253));
    layer0_outputs(1530) <= (inputs(244)) xor (inputs(58));
    layer0_outputs(1531) <= (inputs(103)) and not (inputs(234));
    layer0_outputs(1532) <= (inputs(172)) and (inputs(252));
    layer0_outputs(1533) <= not((inputs(24)) xor (inputs(161)));
    layer0_outputs(1534) <= inputs(189);
    layer0_outputs(1535) <= not(inputs(134));
    layer0_outputs(1536) <= inputs(222);
    layer0_outputs(1537) <= not((inputs(102)) xor (inputs(70)));
    layer0_outputs(1538) <= not(inputs(26));
    layer0_outputs(1539) <= not((inputs(222)) xor (inputs(86)));
    layer0_outputs(1540) <= not((inputs(0)) xor (inputs(26)));
    layer0_outputs(1541) <= (inputs(213)) and not (inputs(3));
    layer0_outputs(1542) <= not(inputs(58));
    layer0_outputs(1543) <= not((inputs(227)) or (inputs(158)));
    layer0_outputs(1544) <= not(inputs(81)) or (inputs(17));
    layer0_outputs(1545) <= not((inputs(7)) or (inputs(202)));
    layer0_outputs(1546) <= (inputs(145)) or (inputs(212));
    layer0_outputs(1547) <= not((inputs(5)) or (inputs(252)));
    layer0_outputs(1548) <= (inputs(125)) or (inputs(123));
    layer0_outputs(1549) <= (inputs(219)) xor (inputs(159));
    layer0_outputs(1550) <= inputs(108);
    layer0_outputs(1551) <= not((inputs(153)) or (inputs(51)));
    layer0_outputs(1552) <= not((inputs(126)) xor (inputs(116)));
    layer0_outputs(1553) <= (inputs(75)) or (inputs(100));
    layer0_outputs(1554) <= not(inputs(108)) or (inputs(27));
    layer0_outputs(1555) <= not(inputs(89));
    layer0_outputs(1556) <= (inputs(102)) or (inputs(78));
    layer0_outputs(1557) <= inputs(138);
    layer0_outputs(1558) <= (inputs(165)) or (inputs(141));
    layer0_outputs(1559) <= not(inputs(151)) or (inputs(77));
    layer0_outputs(1560) <= (inputs(219)) or (inputs(107));
    layer0_outputs(1561) <= not((inputs(49)) and (inputs(241)));
    layer0_outputs(1562) <= (inputs(106)) xor (inputs(94));
    layer0_outputs(1563) <= not((inputs(164)) or (inputs(86)));
    layer0_outputs(1564) <= '0';
    layer0_outputs(1565) <= not(inputs(107));
    layer0_outputs(1566) <= (inputs(66)) xor (inputs(135));
    layer0_outputs(1567) <= not((inputs(184)) or (inputs(1)));
    layer0_outputs(1568) <= (inputs(80)) xor (inputs(3));
    layer0_outputs(1569) <= not(inputs(211)) or (inputs(145));
    layer0_outputs(1570) <= (inputs(149)) and not (inputs(159));
    layer0_outputs(1571) <= (inputs(98)) and not (inputs(129));
    layer0_outputs(1572) <= (inputs(89)) xor (inputs(168));
    layer0_outputs(1573) <= '0';
    layer0_outputs(1574) <= (inputs(13)) or (inputs(126));
    layer0_outputs(1575) <= inputs(229);
    layer0_outputs(1576) <= (inputs(56)) and not (inputs(254));
    layer0_outputs(1577) <= (inputs(154)) xor (inputs(155));
    layer0_outputs(1578) <= not(inputs(152));
    layer0_outputs(1579) <= not((inputs(221)) xor (inputs(41)));
    layer0_outputs(1580) <= not(inputs(4));
    layer0_outputs(1581) <= (inputs(111)) or (inputs(140));
    layer0_outputs(1582) <= (inputs(54)) and not (inputs(141));
    layer0_outputs(1583) <= not((inputs(190)) xor (inputs(118)));
    layer0_outputs(1584) <= not(inputs(66)) or (inputs(224));
    layer0_outputs(1585) <= not((inputs(101)) or (inputs(228)));
    layer0_outputs(1586) <= not((inputs(87)) and (inputs(18)));
    layer0_outputs(1587) <= not(inputs(9));
    layer0_outputs(1588) <= (inputs(86)) and not (inputs(51));
    layer0_outputs(1589) <= (inputs(206)) and not (inputs(208));
    layer0_outputs(1590) <= (inputs(119)) and (inputs(185));
    layer0_outputs(1591) <= not((inputs(53)) xor (inputs(45)));
    layer0_outputs(1592) <= (inputs(182)) or (inputs(18));
    layer0_outputs(1593) <= (inputs(138)) and not (inputs(63));
    layer0_outputs(1594) <= not(inputs(111));
    layer0_outputs(1595) <= (inputs(104)) xor (inputs(89));
    layer0_outputs(1596) <= not(inputs(139));
    layer0_outputs(1597) <= not((inputs(234)) xor (inputs(125)));
    layer0_outputs(1598) <= (inputs(246)) or (inputs(195));
    layer0_outputs(1599) <= '0';
    layer0_outputs(1600) <= (inputs(64)) and not (inputs(159));
    layer0_outputs(1601) <= (inputs(194)) or (inputs(70));
    layer0_outputs(1602) <= not(inputs(93));
    layer0_outputs(1603) <= (inputs(215)) and (inputs(135));
    layer0_outputs(1604) <= inputs(110);
    layer0_outputs(1605) <= (inputs(136)) xor (inputs(243));
    layer0_outputs(1606) <= not((inputs(32)) and (inputs(206)));
    layer0_outputs(1607) <= not(inputs(197)) or (inputs(249));
    layer0_outputs(1608) <= (inputs(117)) and not (inputs(133));
    layer0_outputs(1609) <= not((inputs(104)) or (inputs(251)));
    layer0_outputs(1610) <= (inputs(1)) and not (inputs(53));
    layer0_outputs(1611) <= not(inputs(220));
    layer0_outputs(1612) <= not(inputs(243)) or (inputs(63));
    layer0_outputs(1613) <= (inputs(245)) xor (inputs(228));
    layer0_outputs(1614) <= not((inputs(151)) xor (inputs(177)));
    layer0_outputs(1615) <= not(inputs(208));
    layer0_outputs(1616) <= (inputs(141)) or (inputs(2));
    layer0_outputs(1617) <= (inputs(9)) and not (inputs(44));
    layer0_outputs(1618) <= (inputs(37)) and not (inputs(244));
    layer0_outputs(1619) <= not(inputs(140)) or (inputs(25));
    layer0_outputs(1620) <= not(inputs(164));
    layer0_outputs(1621) <= not(inputs(114));
    layer0_outputs(1622) <= not(inputs(167));
    layer0_outputs(1623) <= (inputs(223)) and not (inputs(244));
    layer0_outputs(1624) <= '1';
    layer0_outputs(1625) <= not(inputs(232)) or (inputs(193));
    layer0_outputs(1626) <= inputs(14);
    layer0_outputs(1627) <= (inputs(120)) xor (inputs(24));
    layer0_outputs(1628) <= (inputs(232)) and (inputs(253));
    layer0_outputs(1629) <= not((inputs(51)) or (inputs(72)));
    layer0_outputs(1630) <= inputs(185);
    layer0_outputs(1631) <= not(inputs(167));
    layer0_outputs(1632) <= not((inputs(23)) xor (inputs(255)));
    layer0_outputs(1633) <= not((inputs(179)) or (inputs(60)));
    layer0_outputs(1634) <= not(inputs(11));
    layer0_outputs(1635) <= (inputs(40)) xor (inputs(215));
    layer0_outputs(1636) <= (inputs(86)) or (inputs(31));
    layer0_outputs(1637) <= not(inputs(246)) or (inputs(226));
    layer0_outputs(1638) <= (inputs(173)) or (inputs(86));
    layer0_outputs(1639) <= '1';
    layer0_outputs(1640) <= inputs(26);
    layer0_outputs(1641) <= not(inputs(237));
    layer0_outputs(1642) <= not(inputs(44)) or (inputs(91));
    layer0_outputs(1643) <= not((inputs(69)) xor (inputs(51)));
    layer0_outputs(1644) <= (inputs(90)) xor (inputs(130));
    layer0_outputs(1645) <= (inputs(97)) and (inputs(24));
    layer0_outputs(1646) <= not((inputs(155)) or (inputs(125)));
    layer0_outputs(1647) <= not(inputs(93));
    layer0_outputs(1648) <= not((inputs(53)) xor (inputs(79)));
    layer0_outputs(1649) <= (inputs(138)) xor (inputs(17));
    layer0_outputs(1650) <= (inputs(171)) xor (inputs(137));
    layer0_outputs(1651) <= not((inputs(143)) or (inputs(0)));
    layer0_outputs(1652) <= not((inputs(53)) xor (inputs(246)));
    layer0_outputs(1653) <= (inputs(228)) and (inputs(147));
    layer0_outputs(1654) <= not((inputs(87)) or (inputs(114)));
    layer0_outputs(1655) <= not((inputs(58)) or (inputs(249)));
    layer0_outputs(1656) <= (inputs(216)) xor (inputs(132));
    layer0_outputs(1657) <= (inputs(12)) and not (inputs(145));
    layer0_outputs(1658) <= not(inputs(80));
    layer0_outputs(1659) <= not((inputs(103)) xor (inputs(158)));
    layer0_outputs(1660) <= not((inputs(71)) xor (inputs(207)));
    layer0_outputs(1661) <= '1';
    layer0_outputs(1662) <= '1';
    layer0_outputs(1663) <= (inputs(153)) and not (inputs(221));
    layer0_outputs(1664) <= not((inputs(240)) or (inputs(198)));
    layer0_outputs(1665) <= not(inputs(69)) or (inputs(131));
    layer0_outputs(1666) <= not((inputs(166)) xor (inputs(236)));
    layer0_outputs(1667) <= not(inputs(213));
    layer0_outputs(1668) <= not((inputs(16)) or (inputs(233)));
    layer0_outputs(1669) <= '0';
    layer0_outputs(1670) <= inputs(189);
    layer0_outputs(1671) <= (inputs(57)) xor (inputs(124));
    layer0_outputs(1672) <= (inputs(217)) or (inputs(177));
    layer0_outputs(1673) <= (inputs(218)) or (inputs(215));
    layer0_outputs(1674) <= not((inputs(205)) or (inputs(38)));
    layer0_outputs(1675) <= '1';
    layer0_outputs(1676) <= not((inputs(77)) or (inputs(58)));
    layer0_outputs(1677) <= not((inputs(167)) or (inputs(234)));
    layer0_outputs(1678) <= (inputs(75)) and not (inputs(196));
    layer0_outputs(1679) <= (inputs(189)) or (inputs(190));
    layer0_outputs(1680) <= '1';
    layer0_outputs(1681) <= not((inputs(84)) xor (inputs(43)));
    layer0_outputs(1682) <= not((inputs(59)) xor (inputs(214)));
    layer0_outputs(1683) <= not((inputs(13)) xor (inputs(196)));
    layer0_outputs(1684) <= not(inputs(166));
    layer0_outputs(1685) <= (inputs(194)) xor (inputs(168));
    layer0_outputs(1686) <= not(inputs(230));
    layer0_outputs(1687) <= not((inputs(68)) xor (inputs(47)));
    layer0_outputs(1688) <= inputs(247);
    layer0_outputs(1689) <= not(inputs(131)) or (inputs(144));
    layer0_outputs(1690) <= not((inputs(13)) xor (inputs(159)));
    layer0_outputs(1691) <= not(inputs(81)) or (inputs(159));
    layer0_outputs(1692) <= not(inputs(183)) or (inputs(77));
    layer0_outputs(1693) <= not((inputs(141)) and (inputs(101)));
    layer0_outputs(1694) <= not(inputs(165)) or (inputs(82));
    layer0_outputs(1695) <= not(inputs(101));
    layer0_outputs(1696) <= not((inputs(6)) xor (inputs(103)));
    layer0_outputs(1697) <= not((inputs(8)) or (inputs(244)));
    layer0_outputs(1698) <= not(inputs(41)) or (inputs(93));
    layer0_outputs(1699) <= inputs(220);
    layer0_outputs(1700) <= (inputs(235)) xor (inputs(224));
    layer0_outputs(1701) <= not((inputs(24)) xor (inputs(248)));
    layer0_outputs(1702) <= not(inputs(53));
    layer0_outputs(1703) <= (inputs(254)) and (inputs(184));
    layer0_outputs(1704) <= inputs(11);
    layer0_outputs(1705) <= (inputs(60)) and not (inputs(254));
    layer0_outputs(1706) <= not((inputs(82)) or (inputs(164)));
    layer0_outputs(1707) <= (inputs(107)) or (inputs(201));
    layer0_outputs(1708) <= inputs(26);
    layer0_outputs(1709) <= not((inputs(122)) or (inputs(228)));
    layer0_outputs(1710) <= not(inputs(105)) or (inputs(79));
    layer0_outputs(1711) <= inputs(166);
    layer0_outputs(1712) <= inputs(126);
    layer0_outputs(1713) <= (inputs(64)) or (inputs(69));
    layer0_outputs(1714) <= not((inputs(131)) or (inputs(239)));
    layer0_outputs(1715) <= inputs(66);
    layer0_outputs(1716) <= (inputs(75)) or (inputs(203));
    layer0_outputs(1717) <= not(inputs(46));
    layer0_outputs(1718) <= not(inputs(234));
    layer0_outputs(1719) <= (inputs(118)) xor (inputs(240));
    layer0_outputs(1720) <= (inputs(95)) and not (inputs(0));
    layer0_outputs(1721) <= not((inputs(22)) or (inputs(83)));
    layer0_outputs(1722) <= (inputs(101)) and not (inputs(178));
    layer0_outputs(1723) <= inputs(92);
    layer0_outputs(1724) <= (inputs(156)) or (inputs(130));
    layer0_outputs(1725) <= not((inputs(94)) or (inputs(212)));
    layer0_outputs(1726) <= (inputs(119)) and not (inputs(185));
    layer0_outputs(1727) <= not((inputs(114)) or (inputs(249)));
    layer0_outputs(1728) <= (inputs(76)) xor (inputs(241));
    layer0_outputs(1729) <= not(inputs(72)) or (inputs(77));
    layer0_outputs(1730) <= inputs(203);
    layer0_outputs(1731) <= inputs(32);
    layer0_outputs(1732) <= inputs(10);
    layer0_outputs(1733) <= not(inputs(240));
    layer0_outputs(1734) <= not((inputs(114)) xor (inputs(150)));
    layer0_outputs(1735) <= not(inputs(233)) or (inputs(82));
    layer0_outputs(1736) <= not(inputs(88));
    layer0_outputs(1737) <= not(inputs(132)) or (inputs(195));
    layer0_outputs(1738) <= not((inputs(39)) or (inputs(37)));
    layer0_outputs(1739) <= not(inputs(158)) or (inputs(8));
    layer0_outputs(1740) <= not(inputs(202)) or (inputs(22));
    layer0_outputs(1741) <= inputs(230);
    layer0_outputs(1742) <= not(inputs(234));
    layer0_outputs(1743) <= not(inputs(202)) or (inputs(44));
    layer0_outputs(1744) <= not(inputs(8));
    layer0_outputs(1745) <= not(inputs(99));
    layer0_outputs(1746) <= (inputs(49)) and not (inputs(142));
    layer0_outputs(1747) <= not((inputs(30)) xor (inputs(52)));
    layer0_outputs(1748) <= (inputs(233)) xor (inputs(201));
    layer0_outputs(1749) <= not((inputs(77)) or (inputs(217)));
    layer0_outputs(1750) <= inputs(39);
    layer0_outputs(1751) <= not(inputs(234));
    layer0_outputs(1752) <= not((inputs(154)) xor (inputs(21)));
    layer0_outputs(1753) <= not(inputs(186));
    layer0_outputs(1754) <= not(inputs(119)) or (inputs(111));
    layer0_outputs(1755) <= (inputs(38)) and not (inputs(99));
    layer0_outputs(1756) <= (inputs(104)) or (inputs(212));
    layer0_outputs(1757) <= inputs(132);
    layer0_outputs(1758) <= not(inputs(75));
    layer0_outputs(1759) <= inputs(126);
    layer0_outputs(1760) <= (inputs(213)) or (inputs(44));
    layer0_outputs(1761) <= inputs(224);
    layer0_outputs(1762) <= (inputs(13)) and not (inputs(51));
    layer0_outputs(1763) <= (inputs(254)) and not (inputs(96));
    layer0_outputs(1764) <= not(inputs(169));
    layer0_outputs(1765) <= not(inputs(167)) or (inputs(112));
    layer0_outputs(1766) <= (inputs(16)) or (inputs(188));
    layer0_outputs(1767) <= not(inputs(132));
    layer0_outputs(1768) <= not(inputs(85));
    layer0_outputs(1769) <= inputs(167);
    layer0_outputs(1770) <= not((inputs(187)) or (inputs(163)));
    layer0_outputs(1771) <= (inputs(62)) and (inputs(251));
    layer0_outputs(1772) <= (inputs(74)) xor (inputs(143));
    layer0_outputs(1773) <= '0';
    layer0_outputs(1774) <= not((inputs(10)) xor (inputs(195)));
    layer0_outputs(1775) <= inputs(187);
    layer0_outputs(1776) <= inputs(214);
    layer0_outputs(1777) <= (inputs(79)) xor (inputs(3));
    layer0_outputs(1778) <= '1';
    layer0_outputs(1779) <= not((inputs(237)) xor (inputs(253)));
    layer0_outputs(1780) <= not(inputs(233));
    layer0_outputs(1781) <= not(inputs(180)) or (inputs(154));
    layer0_outputs(1782) <= not(inputs(229));
    layer0_outputs(1783) <= not((inputs(42)) xor (inputs(241)));
    layer0_outputs(1784) <= not(inputs(220)) or (inputs(7));
    layer0_outputs(1785) <= inputs(152);
    layer0_outputs(1786) <= not(inputs(105));
    layer0_outputs(1787) <= not((inputs(252)) or (inputs(125)));
    layer0_outputs(1788) <= (inputs(3)) and not (inputs(238));
    layer0_outputs(1789) <= not(inputs(122));
    layer0_outputs(1790) <= not((inputs(60)) or (inputs(151)));
    layer0_outputs(1791) <= inputs(57);
    layer0_outputs(1792) <= not((inputs(90)) xor (inputs(190)));
    layer0_outputs(1793) <= (inputs(83)) and not (inputs(62));
    layer0_outputs(1794) <= not(inputs(187));
    layer0_outputs(1795) <= '0';
    layer0_outputs(1796) <= (inputs(138)) and not (inputs(177));
    layer0_outputs(1797) <= not(inputs(133));
    layer0_outputs(1798) <= not(inputs(173));
    layer0_outputs(1799) <= not(inputs(133));
    layer0_outputs(1800) <= not(inputs(105)) or (inputs(235));
    layer0_outputs(1801) <= not(inputs(206)) or (inputs(20));
    layer0_outputs(1802) <= not(inputs(234)) or (inputs(87));
    layer0_outputs(1803) <= (inputs(244)) xor (inputs(104));
    layer0_outputs(1804) <= not(inputs(245));
    layer0_outputs(1805) <= (inputs(73)) and not (inputs(247));
    layer0_outputs(1806) <= (inputs(37)) or (inputs(186));
    layer0_outputs(1807) <= (inputs(166)) and not (inputs(90));
    layer0_outputs(1808) <= not(inputs(74));
    layer0_outputs(1809) <= not((inputs(248)) and (inputs(230)));
    layer0_outputs(1810) <= (inputs(96)) xor (inputs(168));
    layer0_outputs(1811) <= (inputs(36)) or (inputs(177));
    layer0_outputs(1812) <= not((inputs(172)) or (inputs(230)));
    layer0_outputs(1813) <= not((inputs(253)) xor (inputs(96)));
    layer0_outputs(1814) <= (inputs(245)) xor (inputs(70));
    layer0_outputs(1815) <= (inputs(45)) and (inputs(233));
    layer0_outputs(1816) <= not(inputs(100));
    layer0_outputs(1817) <= (inputs(189)) xor (inputs(101));
    layer0_outputs(1818) <= not((inputs(56)) and (inputs(11)));
    layer0_outputs(1819) <= not((inputs(255)) and (inputs(253)));
    layer0_outputs(1820) <= inputs(70);
    layer0_outputs(1821) <= (inputs(243)) xor (inputs(136));
    layer0_outputs(1822) <= inputs(123);
    layer0_outputs(1823) <= not(inputs(106));
    layer0_outputs(1824) <= not((inputs(254)) xor (inputs(119)));
    layer0_outputs(1825) <= not(inputs(93));
    layer0_outputs(1826) <= (inputs(105)) or (inputs(82));
    layer0_outputs(1827) <= (inputs(205)) and not (inputs(18));
    layer0_outputs(1828) <= (inputs(230)) and not (inputs(63));
    layer0_outputs(1829) <= not((inputs(76)) xor (inputs(197)));
    layer0_outputs(1830) <= (inputs(213)) or (inputs(131));
    layer0_outputs(1831) <= (inputs(154)) xor (inputs(172));
    layer0_outputs(1832) <= (inputs(240)) and not (inputs(210));
    layer0_outputs(1833) <= (inputs(156)) xor (inputs(89));
    layer0_outputs(1834) <= not(inputs(96));
    layer0_outputs(1835) <= not(inputs(219));
    layer0_outputs(1836) <= not((inputs(11)) xor (inputs(150)));
    layer0_outputs(1837) <= not((inputs(73)) xor (inputs(5)));
    layer0_outputs(1838) <= (inputs(142)) or (inputs(180));
    layer0_outputs(1839) <= (inputs(19)) or (inputs(104));
    layer0_outputs(1840) <= not((inputs(120)) or (inputs(235)));
    layer0_outputs(1841) <= not(inputs(227));
    layer0_outputs(1842) <= (inputs(75)) or (inputs(146));
    layer0_outputs(1843) <= inputs(230);
    layer0_outputs(1844) <= not(inputs(105));
    layer0_outputs(1845) <= '0';
    layer0_outputs(1846) <= inputs(20);
    layer0_outputs(1847) <= '0';
    layer0_outputs(1848) <= not(inputs(134)) or (inputs(53));
    layer0_outputs(1849) <= not(inputs(225));
    layer0_outputs(1850) <= not(inputs(76));
    layer0_outputs(1851) <= not(inputs(193));
    layer0_outputs(1852) <= not((inputs(79)) or (inputs(154)));
    layer0_outputs(1853) <= not(inputs(19));
    layer0_outputs(1854) <= (inputs(121)) and not (inputs(57));
    layer0_outputs(1855) <= (inputs(121)) or (inputs(179));
    layer0_outputs(1856) <= not((inputs(31)) xor (inputs(91)));
    layer0_outputs(1857) <= (inputs(88)) and not (inputs(14));
    layer0_outputs(1858) <= (inputs(162)) or (inputs(166));
    layer0_outputs(1859) <= inputs(236);
    layer0_outputs(1860) <= not(inputs(97)) or (inputs(126));
    layer0_outputs(1861) <= not(inputs(117)) or (inputs(180));
    layer0_outputs(1862) <= (inputs(157)) xor (inputs(231));
    layer0_outputs(1863) <= not(inputs(165));
    layer0_outputs(1864) <= (inputs(216)) and not (inputs(246));
    layer0_outputs(1865) <= not((inputs(12)) or (inputs(121)));
    layer0_outputs(1866) <= not(inputs(150)) or (inputs(8));
    layer0_outputs(1867) <= (inputs(145)) and not (inputs(236));
    layer0_outputs(1868) <= not((inputs(153)) xor (inputs(186)));
    layer0_outputs(1869) <= (inputs(51)) xor (inputs(230));
    layer0_outputs(1870) <= (inputs(208)) and not (inputs(65));
    layer0_outputs(1871) <= not((inputs(4)) and (inputs(177)));
    layer0_outputs(1872) <= (inputs(197)) and not (inputs(193));
    layer0_outputs(1873) <= (inputs(118)) and not (inputs(18));
    layer0_outputs(1874) <= not(inputs(175));
    layer0_outputs(1875) <= (inputs(136)) and not (inputs(162));
    layer0_outputs(1876) <= not((inputs(98)) xor (inputs(232)));
    layer0_outputs(1877) <= '0';
    layer0_outputs(1878) <= (inputs(193)) or (inputs(202));
    layer0_outputs(1879) <= not(inputs(189)) or (inputs(79));
    layer0_outputs(1880) <= not((inputs(148)) xor (inputs(47)));
    layer0_outputs(1881) <= not(inputs(43)) or (inputs(218));
    layer0_outputs(1882) <= (inputs(88)) and not (inputs(243));
    layer0_outputs(1883) <= (inputs(176)) and (inputs(36));
    layer0_outputs(1884) <= not((inputs(150)) or (inputs(143)));
    layer0_outputs(1885) <= (inputs(205)) or (inputs(210));
    layer0_outputs(1886) <= not(inputs(65)) or (inputs(57));
    layer0_outputs(1887) <= (inputs(36)) xor (inputs(62));
    layer0_outputs(1888) <= (inputs(225)) xor (inputs(138));
    layer0_outputs(1889) <= (inputs(57)) and not (inputs(45));
    layer0_outputs(1890) <= not((inputs(246)) or (inputs(70)));
    layer0_outputs(1891) <= not(inputs(220)) or (inputs(33));
    layer0_outputs(1892) <= (inputs(234)) and not (inputs(189));
    layer0_outputs(1893) <= (inputs(37)) and not (inputs(25));
    layer0_outputs(1894) <= not((inputs(51)) xor (inputs(176)));
    layer0_outputs(1895) <= not((inputs(69)) xor (inputs(3)));
    layer0_outputs(1896) <= (inputs(180)) or (inputs(110));
    layer0_outputs(1897) <= (inputs(223)) or (inputs(185));
    layer0_outputs(1898) <= (inputs(199)) and not (inputs(159));
    layer0_outputs(1899) <= (inputs(191)) or (inputs(109));
    layer0_outputs(1900) <= inputs(182);
    layer0_outputs(1901) <= (inputs(153)) and not (inputs(43));
    layer0_outputs(1902) <= not(inputs(137)) or (inputs(13));
    layer0_outputs(1903) <= (inputs(6)) and not (inputs(254));
    layer0_outputs(1904) <= inputs(169);
    layer0_outputs(1905) <= not(inputs(131)) or (inputs(159));
    layer0_outputs(1906) <= not((inputs(124)) xor (inputs(183)));
    layer0_outputs(1907) <= (inputs(141)) and not (inputs(142));
    layer0_outputs(1908) <= inputs(208);
    layer0_outputs(1909) <= (inputs(189)) xor (inputs(146));
    layer0_outputs(1910) <= not(inputs(10)) or (inputs(158));
    layer0_outputs(1911) <= (inputs(72)) or (inputs(82));
    layer0_outputs(1912) <= (inputs(56)) and not (inputs(131));
    layer0_outputs(1913) <= (inputs(115)) or (inputs(73));
    layer0_outputs(1914) <= (inputs(70)) and (inputs(12));
    layer0_outputs(1915) <= (inputs(71)) and not (inputs(212));
    layer0_outputs(1916) <= not(inputs(32));
    layer0_outputs(1917) <= not((inputs(24)) xor (inputs(9)));
    layer0_outputs(1918) <= inputs(196);
    layer0_outputs(1919) <= (inputs(14)) or (inputs(99));
    layer0_outputs(1920) <= (inputs(223)) xor (inputs(253));
    layer0_outputs(1921) <= (inputs(226)) xor (inputs(46));
    layer0_outputs(1922) <= inputs(131);
    layer0_outputs(1923) <= inputs(1);
    layer0_outputs(1924) <= (inputs(132)) and not (inputs(22));
    layer0_outputs(1925) <= not(inputs(150)) or (inputs(225));
    layer0_outputs(1926) <= not((inputs(166)) or (inputs(2)));
    layer0_outputs(1927) <= not(inputs(163));
    layer0_outputs(1928) <= not(inputs(94)) or (inputs(45));
    layer0_outputs(1929) <= inputs(137);
    layer0_outputs(1930) <= (inputs(145)) and (inputs(192));
    layer0_outputs(1931) <= not(inputs(75)) or (inputs(7));
    layer0_outputs(1932) <= not(inputs(22));
    layer0_outputs(1933) <= (inputs(175)) and not (inputs(114));
    layer0_outputs(1934) <= not((inputs(53)) xor (inputs(176)));
    layer0_outputs(1935) <= not(inputs(46));
    layer0_outputs(1936) <= not((inputs(101)) or (inputs(115)));
    layer0_outputs(1937) <= not((inputs(18)) xor (inputs(140)));
    layer0_outputs(1938) <= (inputs(1)) or (inputs(107));
    layer0_outputs(1939) <= '1';
    layer0_outputs(1940) <= not((inputs(235)) xor (inputs(44)));
    layer0_outputs(1941) <= (inputs(219)) or (inputs(175));
    layer0_outputs(1942) <= not(inputs(24));
    layer0_outputs(1943) <= not(inputs(122)) or (inputs(249));
    layer0_outputs(1944) <= inputs(126);
    layer0_outputs(1945) <= (inputs(74)) or (inputs(211));
    layer0_outputs(1946) <= not((inputs(235)) or (inputs(20)));
    layer0_outputs(1947) <= inputs(99);
    layer0_outputs(1948) <= not(inputs(169)) or (inputs(232));
    layer0_outputs(1949) <= not((inputs(142)) xor (inputs(8)));
    layer0_outputs(1950) <= inputs(135);
    layer0_outputs(1951) <= not((inputs(108)) or (inputs(54)));
    layer0_outputs(1952) <= not((inputs(89)) xor (inputs(106)));
    layer0_outputs(1953) <= not(inputs(184));
    layer0_outputs(1954) <= (inputs(162)) and not (inputs(160));
    layer0_outputs(1955) <= (inputs(146)) xor (inputs(211));
    layer0_outputs(1956) <= not(inputs(167));
    layer0_outputs(1957) <= not(inputs(218)) or (inputs(220));
    layer0_outputs(1958) <= not(inputs(144));
    layer0_outputs(1959) <= not((inputs(11)) or (inputs(253)));
    layer0_outputs(1960) <= (inputs(132)) or (inputs(183));
    layer0_outputs(1961) <= not((inputs(120)) or (inputs(189)));
    layer0_outputs(1962) <= (inputs(93)) and not (inputs(242));
    layer0_outputs(1963) <= (inputs(144)) or (inputs(77));
    layer0_outputs(1964) <= (inputs(164)) and not (inputs(60));
    layer0_outputs(1965) <= inputs(147);
    layer0_outputs(1966) <= not((inputs(137)) and (inputs(122)));
    layer0_outputs(1967) <= inputs(171);
    layer0_outputs(1968) <= not(inputs(105));
    layer0_outputs(1969) <= not((inputs(150)) or (inputs(183)));
    layer0_outputs(1970) <= not((inputs(230)) xor (inputs(14)));
    layer0_outputs(1971) <= (inputs(242)) or (inputs(250));
    layer0_outputs(1972) <= (inputs(114)) and not (inputs(112));
    layer0_outputs(1973) <= not((inputs(168)) or (inputs(36)));
    layer0_outputs(1974) <= (inputs(189)) and not (inputs(251));
    layer0_outputs(1975) <= inputs(167);
    layer0_outputs(1976) <= not((inputs(164)) or (inputs(243)));
    layer0_outputs(1977) <= not((inputs(60)) xor (inputs(215)));
    layer0_outputs(1978) <= not((inputs(122)) or (inputs(231)));
    layer0_outputs(1979) <= not(inputs(189));
    layer0_outputs(1980) <= (inputs(104)) and not (inputs(32));
    layer0_outputs(1981) <= (inputs(150)) and not (inputs(78));
    layer0_outputs(1982) <= not((inputs(240)) xor (inputs(100)));
    layer0_outputs(1983) <= not(inputs(75)) or (inputs(4));
    layer0_outputs(1984) <= inputs(38);
    layer0_outputs(1985) <= (inputs(182)) or (inputs(222));
    layer0_outputs(1986) <= (inputs(246)) or (inputs(39));
    layer0_outputs(1987) <= (inputs(136)) and not (inputs(52));
    layer0_outputs(1988) <= not((inputs(131)) xor (inputs(96)));
    layer0_outputs(1989) <= (inputs(92)) or (inputs(248));
    layer0_outputs(1990) <= not((inputs(186)) or (inputs(17)));
    layer0_outputs(1991) <= not(inputs(81)) or (inputs(2));
    layer0_outputs(1992) <= not((inputs(195)) or (inputs(95)));
    layer0_outputs(1993) <= not((inputs(172)) or (inputs(215)));
    layer0_outputs(1994) <= (inputs(170)) and not (inputs(251));
    layer0_outputs(1995) <= inputs(165);
    layer0_outputs(1996) <= (inputs(114)) or (inputs(180));
    layer0_outputs(1997) <= not((inputs(136)) or (inputs(130)));
    layer0_outputs(1998) <= (inputs(240)) or (inputs(165));
    layer0_outputs(1999) <= not((inputs(240)) or (inputs(174)));
    layer0_outputs(2000) <= not(inputs(6)) or (inputs(59));
    layer0_outputs(2001) <= (inputs(9)) xor (inputs(30));
    layer0_outputs(2002) <= (inputs(226)) and (inputs(104));
    layer0_outputs(2003) <= (inputs(117)) and not (inputs(225));
    layer0_outputs(2004) <= inputs(52);
    layer0_outputs(2005) <= not(inputs(31));
    layer0_outputs(2006) <= not((inputs(53)) or (inputs(158)));
    layer0_outputs(2007) <= not(inputs(68)) or (inputs(19));
    layer0_outputs(2008) <= not(inputs(108));
    layer0_outputs(2009) <= inputs(227);
    layer0_outputs(2010) <= not((inputs(74)) or (inputs(153)));
    layer0_outputs(2011) <= not((inputs(255)) xor (inputs(236)));
    layer0_outputs(2012) <= (inputs(1)) xor (inputs(103));
    layer0_outputs(2013) <= (inputs(37)) and (inputs(128));
    layer0_outputs(2014) <= (inputs(55)) xor (inputs(57));
    layer0_outputs(2015) <= inputs(25);
    layer0_outputs(2016) <= not(inputs(185));
    layer0_outputs(2017) <= (inputs(101)) and not (inputs(19));
    layer0_outputs(2018) <= not((inputs(27)) or (inputs(251)));
    layer0_outputs(2019) <= not(inputs(214));
    layer0_outputs(2020) <= not((inputs(194)) xor (inputs(75)));
    layer0_outputs(2021) <= inputs(134);
    layer0_outputs(2022) <= not(inputs(132));
    layer0_outputs(2023) <= (inputs(121)) and not (inputs(98));
    layer0_outputs(2024) <= not((inputs(81)) xor (inputs(148)));
    layer0_outputs(2025) <= (inputs(65)) and not (inputs(78));
    layer0_outputs(2026) <= not((inputs(36)) or (inputs(185)));
    layer0_outputs(2027) <= (inputs(96)) or (inputs(77));
    layer0_outputs(2028) <= (inputs(21)) or (inputs(197));
    layer0_outputs(2029) <= (inputs(68)) or (inputs(46));
    layer0_outputs(2030) <= inputs(126);
    layer0_outputs(2031) <= not((inputs(55)) xor (inputs(179)));
    layer0_outputs(2032) <= not((inputs(58)) xor (inputs(206)));
    layer0_outputs(2033) <= not(inputs(106)) or (inputs(186));
    layer0_outputs(2034) <= (inputs(103)) and not (inputs(46));
    layer0_outputs(2035) <= (inputs(212)) xor (inputs(250));
    layer0_outputs(2036) <= not(inputs(168)) or (inputs(94));
    layer0_outputs(2037) <= '0';
    layer0_outputs(2038) <= inputs(136);
    layer0_outputs(2039) <= (inputs(69)) or (inputs(124));
    layer0_outputs(2040) <= not(inputs(223)) or (inputs(61));
    layer0_outputs(2041) <= '0';
    layer0_outputs(2042) <= not(inputs(190));
    layer0_outputs(2043) <= not(inputs(73));
    layer0_outputs(2044) <= not((inputs(183)) and (inputs(230)));
    layer0_outputs(2045) <= not((inputs(187)) or (inputs(225)));
    layer0_outputs(2046) <= '1';
    layer0_outputs(2047) <= (inputs(159)) xor (inputs(82));
    layer0_outputs(2048) <= not(inputs(94)) or (inputs(48));
    layer0_outputs(2049) <= not(inputs(214)) or (inputs(245));
    layer0_outputs(2050) <= not(inputs(134));
    layer0_outputs(2051) <= not(inputs(242)) or (inputs(127));
    layer0_outputs(2052) <= (inputs(244)) xor (inputs(75));
    layer0_outputs(2053) <= '1';
    layer0_outputs(2054) <= not((inputs(115)) or (inputs(112)));
    layer0_outputs(2055) <= not((inputs(84)) xor (inputs(53)));
    layer0_outputs(2056) <= not((inputs(216)) xor (inputs(32)));
    layer0_outputs(2057) <= not((inputs(84)) or (inputs(252)));
    layer0_outputs(2058) <= (inputs(215)) and not (inputs(208));
    layer0_outputs(2059) <= (inputs(170)) or (inputs(226));
    layer0_outputs(2060) <= (inputs(110)) or (inputs(27));
    layer0_outputs(2061) <= not((inputs(43)) xor (inputs(77)));
    layer0_outputs(2062) <= not(inputs(43)) or (inputs(7));
    layer0_outputs(2063) <= (inputs(106)) and not (inputs(185));
    layer0_outputs(2064) <= not(inputs(6));
    layer0_outputs(2065) <= inputs(191);
    layer0_outputs(2066) <= inputs(179);
    layer0_outputs(2067) <= (inputs(170)) and not (inputs(221));
    layer0_outputs(2068) <= inputs(116);
    layer0_outputs(2069) <= not((inputs(53)) xor (inputs(208)));
    layer0_outputs(2070) <= (inputs(86)) or (inputs(108));
    layer0_outputs(2071) <= inputs(228);
    layer0_outputs(2072) <= (inputs(27)) xor (inputs(140));
    layer0_outputs(2073) <= not((inputs(240)) or (inputs(24)));
    layer0_outputs(2074) <= not((inputs(90)) xor (inputs(243)));
    layer0_outputs(2075) <= (inputs(8)) xor (inputs(44));
    layer0_outputs(2076) <= inputs(123);
    layer0_outputs(2077) <= not((inputs(85)) xor (inputs(106)));
    layer0_outputs(2078) <= not((inputs(250)) xor (inputs(184)));
    layer0_outputs(2079) <= not(inputs(60)) or (inputs(253));
    layer0_outputs(2080) <= (inputs(71)) and not (inputs(29));
    layer0_outputs(2081) <= inputs(53);
    layer0_outputs(2082) <= not((inputs(45)) xor (inputs(152)));
    layer0_outputs(2083) <= not(inputs(78));
    layer0_outputs(2084) <= not(inputs(28)) or (inputs(245));
    layer0_outputs(2085) <= not((inputs(70)) xor (inputs(200)));
    layer0_outputs(2086) <= (inputs(240)) xor (inputs(243));
    layer0_outputs(2087) <= (inputs(229)) and not (inputs(160));
    layer0_outputs(2088) <= not(inputs(89));
    layer0_outputs(2089) <= (inputs(81)) and not (inputs(218));
    layer0_outputs(2090) <= not((inputs(184)) or (inputs(30)));
    layer0_outputs(2091) <= (inputs(164)) and not (inputs(41));
    layer0_outputs(2092) <= '0';
    layer0_outputs(2093) <= not(inputs(168));
    layer0_outputs(2094) <= not((inputs(161)) and (inputs(66)));
    layer0_outputs(2095) <= inputs(42);
    layer0_outputs(2096) <= (inputs(10)) or (inputs(91));
    layer0_outputs(2097) <= not((inputs(49)) xor (inputs(61)));
    layer0_outputs(2098) <= (inputs(2)) or (inputs(190));
    layer0_outputs(2099) <= not(inputs(202)) or (inputs(22));
    layer0_outputs(2100) <= inputs(179);
    layer0_outputs(2101) <= not(inputs(255));
    layer0_outputs(2102) <= not((inputs(149)) or (inputs(39)));
    layer0_outputs(2103) <= (inputs(46)) and (inputs(41));
    layer0_outputs(2104) <= not((inputs(252)) or (inputs(15)));
    layer0_outputs(2105) <= inputs(227);
    layer0_outputs(2106) <= '1';
    layer0_outputs(2107) <= (inputs(167)) and not (inputs(155));
    layer0_outputs(2108) <= (inputs(98)) or (inputs(154));
    layer0_outputs(2109) <= not((inputs(73)) xor (inputs(208)));
    layer0_outputs(2110) <= (inputs(198)) xor (inputs(182));
    layer0_outputs(2111) <= (inputs(102)) and not (inputs(197));
    layer0_outputs(2112) <= (inputs(167)) and not (inputs(33));
    layer0_outputs(2113) <= not((inputs(104)) or (inputs(36)));
    layer0_outputs(2114) <= (inputs(174)) xor (inputs(159));
    layer0_outputs(2115) <= inputs(191);
    layer0_outputs(2116) <= (inputs(81)) or (inputs(237));
    layer0_outputs(2117) <= (inputs(217)) and not (inputs(15));
    layer0_outputs(2118) <= (inputs(223)) or (inputs(234));
    layer0_outputs(2119) <= inputs(131);
    layer0_outputs(2120) <= not(inputs(248));
    layer0_outputs(2121) <= not(inputs(57));
    layer0_outputs(2122) <= not(inputs(56));
    layer0_outputs(2123) <= (inputs(197)) or (inputs(180));
    layer0_outputs(2124) <= not((inputs(190)) xor (inputs(19)));
    layer0_outputs(2125) <= (inputs(185)) or (inputs(110));
    layer0_outputs(2126) <= not(inputs(220));
    layer0_outputs(2127) <= inputs(136);
    layer0_outputs(2128) <= not(inputs(235));
    layer0_outputs(2129) <= not(inputs(52)) or (inputs(246));
    layer0_outputs(2130) <= not(inputs(102)) or (inputs(110));
    layer0_outputs(2131) <= (inputs(39)) xor (inputs(95));
    layer0_outputs(2132) <= not(inputs(103));
    layer0_outputs(2133) <= (inputs(200)) xor (inputs(41));
    layer0_outputs(2134) <= not(inputs(201));
    layer0_outputs(2135) <= inputs(106);
    layer0_outputs(2136) <= not(inputs(170));
    layer0_outputs(2137) <= (inputs(117)) or (inputs(60));
    layer0_outputs(2138) <= not((inputs(111)) or (inputs(62)));
    layer0_outputs(2139) <= not((inputs(139)) xor (inputs(92)));
    layer0_outputs(2140) <= (inputs(130)) xor (inputs(49));
    layer0_outputs(2141) <= not((inputs(65)) xor (inputs(60)));
    layer0_outputs(2142) <= not((inputs(211)) and (inputs(37)));
    layer0_outputs(2143) <= not((inputs(19)) xor (inputs(119)));
    layer0_outputs(2144) <= not(inputs(110));
    layer0_outputs(2145) <= not(inputs(63));
    layer0_outputs(2146) <= not(inputs(117));
    layer0_outputs(2147) <= (inputs(40)) or (inputs(116));
    layer0_outputs(2148) <= not((inputs(204)) xor (inputs(88)));
    layer0_outputs(2149) <= not(inputs(40)) or (inputs(46));
    layer0_outputs(2150) <= not((inputs(88)) xor (inputs(118)));
    layer0_outputs(2151) <= '0';
    layer0_outputs(2152) <= (inputs(209)) or (inputs(0));
    layer0_outputs(2153) <= not(inputs(174)) or (inputs(82));
    layer0_outputs(2154) <= (inputs(87)) or (inputs(59));
    layer0_outputs(2155) <= not(inputs(233));
    layer0_outputs(2156) <= not((inputs(155)) or (inputs(129)));
    layer0_outputs(2157) <= inputs(161);
    layer0_outputs(2158) <= inputs(167);
    layer0_outputs(2159) <= not(inputs(141));
    layer0_outputs(2160) <= inputs(85);
    layer0_outputs(2161) <= inputs(227);
    layer0_outputs(2162) <= not((inputs(98)) or (inputs(12)));
    layer0_outputs(2163) <= not(inputs(228));
    layer0_outputs(2164) <= not(inputs(106)) or (inputs(173));
    layer0_outputs(2165) <= (inputs(210)) xor (inputs(5));
    layer0_outputs(2166) <= inputs(229);
    layer0_outputs(2167) <= not(inputs(217));
    layer0_outputs(2168) <= (inputs(2)) or (inputs(57));
    layer0_outputs(2169) <= not((inputs(207)) xor (inputs(62)));
    layer0_outputs(2170) <= (inputs(79)) xor (inputs(19));
    layer0_outputs(2171) <= (inputs(51)) and (inputs(173));
    layer0_outputs(2172) <= (inputs(171)) xor (inputs(154));
    layer0_outputs(2173) <= not(inputs(118));
    layer0_outputs(2174) <= not(inputs(226)) or (inputs(20));
    layer0_outputs(2175) <= (inputs(198)) and not (inputs(123));
    layer0_outputs(2176) <= not((inputs(105)) xor (inputs(76)));
    layer0_outputs(2177) <= (inputs(121)) or (inputs(22));
    layer0_outputs(2178) <= (inputs(139)) and not (inputs(88));
    layer0_outputs(2179) <= (inputs(118)) or (inputs(149));
    layer0_outputs(2180) <= not(inputs(24)) or (inputs(253));
    layer0_outputs(2181) <= (inputs(86)) xor (inputs(192));
    layer0_outputs(2182) <= not(inputs(70)) or (inputs(6));
    layer0_outputs(2183) <= not((inputs(93)) xor (inputs(41)));
    layer0_outputs(2184) <= not((inputs(59)) xor (inputs(92)));
    layer0_outputs(2185) <= not((inputs(76)) and (inputs(15)));
    layer0_outputs(2186) <= not(inputs(123)) or (inputs(173));
    layer0_outputs(2187) <= not((inputs(193)) xor (inputs(100)));
    layer0_outputs(2188) <= inputs(241);
    layer0_outputs(2189) <= (inputs(145)) or (inputs(24));
    layer0_outputs(2190) <= not(inputs(167));
    layer0_outputs(2191) <= inputs(138);
    layer0_outputs(2192) <= not(inputs(91));
    layer0_outputs(2193) <= (inputs(6)) or (inputs(23));
    layer0_outputs(2194) <= (inputs(25)) and (inputs(30));
    layer0_outputs(2195) <= (inputs(82)) and not (inputs(248));
    layer0_outputs(2196) <= '0';
    layer0_outputs(2197) <= not(inputs(189)) or (inputs(237));
    layer0_outputs(2198) <= (inputs(11)) xor (inputs(68));
    layer0_outputs(2199) <= not(inputs(124));
    layer0_outputs(2200) <= not((inputs(68)) or (inputs(54)));
    layer0_outputs(2201) <= '0';
    layer0_outputs(2202) <= (inputs(154)) and not (inputs(12));
    layer0_outputs(2203) <= not((inputs(38)) or (inputs(14)));
    layer0_outputs(2204) <= '1';
    layer0_outputs(2205) <= not(inputs(135)) or (inputs(172));
    layer0_outputs(2206) <= not((inputs(174)) xor (inputs(197)));
    layer0_outputs(2207) <= not((inputs(103)) xor (inputs(160)));
    layer0_outputs(2208) <= (inputs(107)) or (inputs(215));
    layer0_outputs(2209) <= not(inputs(92)) or (inputs(193));
    layer0_outputs(2210) <= '1';
    layer0_outputs(2211) <= not(inputs(48)) or (inputs(68));
    layer0_outputs(2212) <= (inputs(41)) and not (inputs(68));
    layer0_outputs(2213) <= not((inputs(23)) or (inputs(174)));
    layer0_outputs(2214) <= not((inputs(159)) xor (inputs(188)));
    layer0_outputs(2215) <= inputs(116);
    layer0_outputs(2216) <= not((inputs(59)) or (inputs(169)));
    layer0_outputs(2217) <= not(inputs(165)) or (inputs(115));
    layer0_outputs(2218) <= (inputs(37)) and not (inputs(125));
    layer0_outputs(2219) <= (inputs(22)) and (inputs(94));
    layer0_outputs(2220) <= (inputs(221)) and (inputs(191));
    layer0_outputs(2221) <= inputs(132);
    layer0_outputs(2222) <= '0';
    layer0_outputs(2223) <= not(inputs(104));
    layer0_outputs(2224) <= not((inputs(142)) or (inputs(185)));
    layer0_outputs(2225) <= (inputs(15)) xor (inputs(175));
    layer0_outputs(2226) <= inputs(102);
    layer0_outputs(2227) <= (inputs(122)) and not (inputs(122));
    layer0_outputs(2228) <= not((inputs(23)) xor (inputs(192)));
    layer0_outputs(2229) <= not(inputs(147)) or (inputs(109));
    layer0_outputs(2230) <= not(inputs(44));
    layer0_outputs(2231) <= not((inputs(60)) xor (inputs(196)));
    layer0_outputs(2232) <= (inputs(13)) or (inputs(212));
    layer0_outputs(2233) <= inputs(88);
    layer0_outputs(2234) <= not((inputs(137)) or (inputs(43)));
    layer0_outputs(2235) <= (inputs(126)) and not (inputs(240));
    layer0_outputs(2236) <= (inputs(75)) and not (inputs(48));
    layer0_outputs(2237) <= not(inputs(77)) or (inputs(145));
    layer0_outputs(2238) <= not(inputs(93)) or (inputs(249));
    layer0_outputs(2239) <= inputs(116);
    layer0_outputs(2240) <= (inputs(78)) xor (inputs(49));
    layer0_outputs(2241) <= not((inputs(142)) or (inputs(166)));
    layer0_outputs(2242) <= not((inputs(214)) xor (inputs(43)));
    layer0_outputs(2243) <= not((inputs(234)) and (inputs(126)));
    layer0_outputs(2244) <= not((inputs(158)) or (inputs(187)));
    layer0_outputs(2245) <= inputs(198);
    layer0_outputs(2246) <= (inputs(47)) and not (inputs(21));
    layer0_outputs(2247) <= (inputs(55)) or (inputs(24));
    layer0_outputs(2248) <= not(inputs(203)) or (inputs(193));
    layer0_outputs(2249) <= not((inputs(253)) or (inputs(200)));
    layer0_outputs(2250) <= not(inputs(247));
    layer0_outputs(2251) <= not(inputs(108));
    layer0_outputs(2252) <= (inputs(70)) and not (inputs(152));
    layer0_outputs(2253) <= inputs(166);
    layer0_outputs(2254) <= not(inputs(19));
    layer0_outputs(2255) <= (inputs(55)) and not (inputs(248));
    layer0_outputs(2256) <= '1';
    layer0_outputs(2257) <= not((inputs(91)) xor (inputs(28)));
    layer0_outputs(2258) <= '0';
    layer0_outputs(2259) <= inputs(133);
    layer0_outputs(2260) <= (inputs(16)) or (inputs(210));
    layer0_outputs(2261) <= not((inputs(101)) or (inputs(175)));
    layer0_outputs(2262) <= not(inputs(50));
    layer0_outputs(2263) <= (inputs(7)) xor (inputs(123));
    layer0_outputs(2264) <= not((inputs(61)) xor (inputs(175)));
    layer0_outputs(2265) <= inputs(100);
    layer0_outputs(2266) <= not(inputs(182));
    layer0_outputs(2267) <= not(inputs(102));
    layer0_outputs(2268) <= inputs(145);
    layer0_outputs(2269) <= not(inputs(131)) or (inputs(31));
    layer0_outputs(2270) <= not((inputs(105)) xor (inputs(66)));
    layer0_outputs(2271) <= not((inputs(138)) and (inputs(0)));
    layer0_outputs(2272) <= not(inputs(90));
    layer0_outputs(2273) <= (inputs(142)) or (inputs(248));
    layer0_outputs(2274) <= not(inputs(217));
    layer0_outputs(2275) <= (inputs(197)) xor (inputs(38));
    layer0_outputs(2276) <= not(inputs(87)) or (inputs(192));
    layer0_outputs(2277) <= not((inputs(49)) xor (inputs(110)));
    layer0_outputs(2278) <= inputs(230);
    layer0_outputs(2279) <= not(inputs(61)) or (inputs(174));
    layer0_outputs(2280) <= not(inputs(57)) or (inputs(192));
    layer0_outputs(2281) <= not(inputs(198)) or (inputs(164));
    layer0_outputs(2282) <= (inputs(192)) and not (inputs(83));
    layer0_outputs(2283) <= (inputs(189)) xor (inputs(197));
    layer0_outputs(2284) <= '0';
    layer0_outputs(2285) <= (inputs(55)) or (inputs(165));
    layer0_outputs(2286) <= not(inputs(228));
    layer0_outputs(2287) <= inputs(133);
    layer0_outputs(2288) <= not(inputs(105)) or (inputs(19));
    layer0_outputs(2289) <= not(inputs(236));
    layer0_outputs(2290) <= '0';
    layer0_outputs(2291) <= not(inputs(185)) or (inputs(239));
    layer0_outputs(2292) <= not((inputs(13)) xor (inputs(191)));
    layer0_outputs(2293) <= '0';
    layer0_outputs(2294) <= inputs(71);
    layer0_outputs(2295) <= not(inputs(110));
    layer0_outputs(2296) <= '0';
    layer0_outputs(2297) <= (inputs(164)) xor (inputs(153));
    layer0_outputs(2298) <= (inputs(199)) or (inputs(31));
    layer0_outputs(2299) <= (inputs(222)) xor (inputs(130));
    layer0_outputs(2300) <= not(inputs(25)) or (inputs(219));
    layer0_outputs(2301) <= (inputs(115)) and not (inputs(209));
    layer0_outputs(2302) <= not(inputs(13));
    layer0_outputs(2303) <= not(inputs(73));
    layer0_outputs(2304) <= (inputs(58)) xor (inputs(158));
    layer0_outputs(2305) <= (inputs(235)) and not (inputs(51));
    layer0_outputs(2306) <= (inputs(15)) or (inputs(25));
    layer0_outputs(2307) <= not(inputs(56));
    layer0_outputs(2308) <= (inputs(243)) or (inputs(138));
    layer0_outputs(2309) <= not(inputs(52)) or (inputs(75));
    layer0_outputs(2310) <= inputs(133);
    layer0_outputs(2311) <= not(inputs(185)) or (inputs(195));
    layer0_outputs(2312) <= not(inputs(246)) or (inputs(235));
    layer0_outputs(2313) <= (inputs(152)) and not (inputs(206));
    layer0_outputs(2314) <= inputs(128);
    layer0_outputs(2315) <= not((inputs(230)) xor (inputs(50)));
    layer0_outputs(2316) <= not((inputs(251)) or (inputs(109)));
    layer0_outputs(2317) <= not(inputs(238));
    layer0_outputs(2318) <= not(inputs(102)) or (inputs(194));
    layer0_outputs(2319) <= inputs(232);
    layer0_outputs(2320) <= '1';
    layer0_outputs(2321) <= not(inputs(161));
    layer0_outputs(2322) <= inputs(223);
    layer0_outputs(2323) <= not(inputs(89));
    layer0_outputs(2324) <= (inputs(249)) and not (inputs(220));
    layer0_outputs(2325) <= not((inputs(233)) or (inputs(24)));
    layer0_outputs(2326) <= not((inputs(236)) xor (inputs(58)));
    layer0_outputs(2327) <= (inputs(234)) or (inputs(236));
    layer0_outputs(2328) <= not(inputs(68)) or (inputs(34));
    layer0_outputs(2329) <= inputs(198);
    layer0_outputs(2330) <= (inputs(242)) and not (inputs(252));
    layer0_outputs(2331) <= (inputs(173)) and not (inputs(5));
    layer0_outputs(2332) <= (inputs(151)) and not (inputs(31));
    layer0_outputs(2333) <= (inputs(39)) and not (inputs(240));
    layer0_outputs(2334) <= (inputs(109)) and not (inputs(31));
    layer0_outputs(2335) <= (inputs(20)) or (inputs(103));
    layer0_outputs(2336) <= not(inputs(210)) or (inputs(154));
    layer0_outputs(2337) <= not(inputs(52));
    layer0_outputs(2338) <= not((inputs(243)) or (inputs(124)));
    layer0_outputs(2339) <= not((inputs(215)) or (inputs(172)));
    layer0_outputs(2340) <= inputs(146);
    layer0_outputs(2341) <= not(inputs(202));
    layer0_outputs(2342) <= (inputs(26)) and (inputs(19));
    layer0_outputs(2343) <= (inputs(201)) xor (inputs(129));
    layer0_outputs(2344) <= (inputs(32)) xor (inputs(44));
    layer0_outputs(2345) <= (inputs(196)) xor (inputs(223));
    layer0_outputs(2346) <= (inputs(69)) or (inputs(127));
    layer0_outputs(2347) <= inputs(118);
    layer0_outputs(2348) <= (inputs(40)) or (inputs(226));
    layer0_outputs(2349) <= not(inputs(41));
    layer0_outputs(2350) <= inputs(81);
    layer0_outputs(2351) <= not(inputs(137));
    layer0_outputs(2352) <= not((inputs(64)) or (inputs(179)));
    layer0_outputs(2353) <= not((inputs(109)) xor (inputs(212)));
    layer0_outputs(2354) <= not((inputs(86)) and (inputs(226)));
    layer0_outputs(2355) <= not((inputs(110)) and (inputs(244)));
    layer0_outputs(2356) <= not(inputs(203)) or (inputs(96));
    layer0_outputs(2357) <= (inputs(99)) and not (inputs(10));
    layer0_outputs(2358) <= inputs(251);
    layer0_outputs(2359) <= (inputs(47)) xor (inputs(110));
    layer0_outputs(2360) <= '0';
    layer0_outputs(2361) <= not((inputs(88)) xor (inputs(242)));
    layer0_outputs(2362) <= (inputs(214)) or (inputs(123));
    layer0_outputs(2363) <= (inputs(162)) and not (inputs(34));
    layer0_outputs(2364) <= not(inputs(204));
    layer0_outputs(2365) <= not(inputs(138));
    layer0_outputs(2366) <= inputs(21);
    layer0_outputs(2367) <= not((inputs(60)) xor (inputs(25)));
    layer0_outputs(2368) <= inputs(153);
    layer0_outputs(2369) <= not(inputs(79));
    layer0_outputs(2370) <= (inputs(124)) xor (inputs(210));
    layer0_outputs(2371) <= not((inputs(13)) or (inputs(107)));
    layer0_outputs(2372) <= not(inputs(162)) or (inputs(13));
    layer0_outputs(2373) <= not((inputs(247)) or (inputs(212)));
    layer0_outputs(2374) <= not(inputs(32)) or (inputs(97));
    layer0_outputs(2375) <= not((inputs(52)) or (inputs(184)));
    layer0_outputs(2376) <= not(inputs(238)) or (inputs(211));
    layer0_outputs(2377) <= inputs(117);
    layer0_outputs(2378) <= '1';
    layer0_outputs(2379) <= (inputs(222)) or (inputs(227));
    layer0_outputs(2380) <= (inputs(163)) and not (inputs(247));
    layer0_outputs(2381) <= not((inputs(171)) or (inputs(189)));
    layer0_outputs(2382) <= not(inputs(134));
    layer0_outputs(2383) <= (inputs(198)) xor (inputs(87));
    layer0_outputs(2384) <= inputs(168);
    layer0_outputs(2385) <= not((inputs(52)) and (inputs(43)));
    layer0_outputs(2386) <= inputs(50);
    layer0_outputs(2387) <= inputs(94);
    layer0_outputs(2388) <= not(inputs(135)) or (inputs(67));
    layer0_outputs(2389) <= not(inputs(113));
    layer0_outputs(2390) <= (inputs(49)) xor (inputs(142));
    layer0_outputs(2391) <= not(inputs(124)) or (inputs(253));
    layer0_outputs(2392) <= (inputs(172)) and not (inputs(114));
    layer0_outputs(2393) <= (inputs(91)) and (inputs(66));
    layer0_outputs(2394) <= not((inputs(243)) xor (inputs(97)));
    layer0_outputs(2395) <= inputs(181);
    layer0_outputs(2396) <= (inputs(14)) and (inputs(254));
    layer0_outputs(2397) <= not(inputs(98));
    layer0_outputs(2398) <= (inputs(230)) xor (inputs(178));
    layer0_outputs(2399) <= not(inputs(15));
    layer0_outputs(2400) <= not(inputs(157));
    layer0_outputs(2401) <= not((inputs(31)) xor (inputs(70)));
    layer0_outputs(2402) <= not(inputs(202));
    layer0_outputs(2403) <= not((inputs(179)) or (inputs(201)));
    layer0_outputs(2404) <= inputs(120);
    layer0_outputs(2405) <= (inputs(88)) and not (inputs(124));
    layer0_outputs(2406) <= not(inputs(233));
    layer0_outputs(2407) <= (inputs(80)) and not (inputs(12));
    layer0_outputs(2408) <= (inputs(107)) or (inputs(213));
    layer0_outputs(2409) <= (inputs(75)) or (inputs(177));
    layer0_outputs(2410) <= not(inputs(42)) or (inputs(111));
    layer0_outputs(2411) <= not((inputs(9)) xor (inputs(15)));
    layer0_outputs(2412) <= (inputs(172)) xor (inputs(7));
    layer0_outputs(2413) <= not(inputs(51));
    layer0_outputs(2414) <= '0';
    layer0_outputs(2415) <= not((inputs(139)) or (inputs(192)));
    layer0_outputs(2416) <= (inputs(78)) xor (inputs(39));
    layer0_outputs(2417) <= not((inputs(239)) or (inputs(117)));
    layer0_outputs(2418) <= (inputs(117)) and not (inputs(7));
    layer0_outputs(2419) <= inputs(121);
    layer0_outputs(2420) <= not(inputs(219));
    layer0_outputs(2421) <= (inputs(66)) or (inputs(229));
    layer0_outputs(2422) <= not(inputs(100)) or (inputs(248));
    layer0_outputs(2423) <= not(inputs(172));
    layer0_outputs(2424) <= not(inputs(170));
    layer0_outputs(2425) <= not(inputs(232));
    layer0_outputs(2426) <= not((inputs(49)) and (inputs(127)));
    layer0_outputs(2427) <= not((inputs(61)) xor (inputs(49)));
    layer0_outputs(2428) <= not((inputs(167)) or (inputs(50)));
    layer0_outputs(2429) <= '1';
    layer0_outputs(2430) <= inputs(25);
    layer0_outputs(2431) <= (inputs(237)) and (inputs(72));
    layer0_outputs(2432) <= (inputs(120)) xor (inputs(111));
    layer0_outputs(2433) <= inputs(214);
    layer0_outputs(2434) <= not((inputs(93)) xor (inputs(7)));
    layer0_outputs(2435) <= not(inputs(119)) or (inputs(26));
    layer0_outputs(2436) <= not((inputs(236)) xor (inputs(144)));
    layer0_outputs(2437) <= '1';
    layer0_outputs(2438) <= inputs(68);
    layer0_outputs(2439) <= (inputs(141)) and not (inputs(5));
    layer0_outputs(2440) <= not((inputs(214)) xor (inputs(217)));
    layer0_outputs(2441) <= '1';
    layer0_outputs(2442) <= not((inputs(70)) or (inputs(81)));
    layer0_outputs(2443) <= not((inputs(32)) or (inputs(129)));
    layer0_outputs(2444) <= inputs(152);
    layer0_outputs(2445) <= inputs(23);
    layer0_outputs(2446) <= not(inputs(17));
    layer0_outputs(2447) <= (inputs(139)) and not (inputs(202));
    layer0_outputs(2448) <= (inputs(207)) xor (inputs(174));
    layer0_outputs(2449) <= not((inputs(90)) or (inputs(12)));
    layer0_outputs(2450) <= (inputs(170)) and not (inputs(194));
    layer0_outputs(2451) <= (inputs(29)) and not (inputs(209));
    layer0_outputs(2452) <= not((inputs(108)) or (inputs(97)));
    layer0_outputs(2453) <= not(inputs(203));
    layer0_outputs(2454) <= not(inputs(111)) or (inputs(7));
    layer0_outputs(2455) <= not(inputs(133));
    layer0_outputs(2456) <= not(inputs(116));
    layer0_outputs(2457) <= inputs(206);
    layer0_outputs(2458) <= (inputs(90)) xor (inputs(31));
    layer0_outputs(2459) <= not(inputs(107));
    layer0_outputs(2460) <= '1';
    layer0_outputs(2461) <= not((inputs(253)) xor (inputs(204)));
    layer0_outputs(2462) <= not((inputs(54)) and (inputs(198)));
    layer0_outputs(2463) <= '1';
    layer0_outputs(2464) <= (inputs(165)) and not (inputs(179));
    layer0_outputs(2465) <= (inputs(13)) or (inputs(45));
    layer0_outputs(2466) <= (inputs(110)) xor (inputs(236));
    layer0_outputs(2467) <= not(inputs(137));
    layer0_outputs(2468) <= (inputs(110)) and not (inputs(20));
    layer0_outputs(2469) <= not((inputs(183)) xor (inputs(125)));
    layer0_outputs(2470) <= not(inputs(89));
    layer0_outputs(2471) <= (inputs(225)) and (inputs(221));
    layer0_outputs(2472) <= (inputs(203)) and not (inputs(241));
    layer0_outputs(2473) <= not((inputs(178)) xor (inputs(53)));
    layer0_outputs(2474) <= inputs(32);
    layer0_outputs(2475) <= '1';
    layer0_outputs(2476) <= inputs(69);
    layer0_outputs(2477) <= (inputs(148)) or (inputs(130));
    layer0_outputs(2478) <= not(inputs(171)) or (inputs(142));
    layer0_outputs(2479) <= (inputs(81)) or (inputs(195));
    layer0_outputs(2480) <= (inputs(20)) or (inputs(176));
    layer0_outputs(2481) <= not((inputs(175)) or (inputs(147)));
    layer0_outputs(2482) <= not(inputs(184));
    layer0_outputs(2483) <= inputs(100);
    layer0_outputs(2484) <= not(inputs(54)) or (inputs(20));
    layer0_outputs(2485) <= not((inputs(108)) and (inputs(111)));
    layer0_outputs(2486) <= (inputs(34)) or (inputs(92));
    layer0_outputs(2487) <= not(inputs(96));
    layer0_outputs(2488) <= not(inputs(89));
    layer0_outputs(2489) <= not((inputs(115)) or (inputs(134)));
    layer0_outputs(2490) <= not(inputs(91)) or (inputs(159));
    layer0_outputs(2491) <= (inputs(93)) xor (inputs(234));
    layer0_outputs(2492) <= (inputs(77)) xor (inputs(107));
    layer0_outputs(2493) <= (inputs(17)) or (inputs(148));
    layer0_outputs(2494) <= not((inputs(10)) or (inputs(185)));
    layer0_outputs(2495) <= not((inputs(65)) or (inputs(212)));
    layer0_outputs(2496) <= (inputs(170)) xor (inputs(135));
    layer0_outputs(2497) <= inputs(64);
    layer0_outputs(2498) <= (inputs(40)) and not (inputs(64));
    layer0_outputs(2499) <= not(inputs(105));
    layer0_outputs(2500) <= not(inputs(55)) or (inputs(144));
    layer0_outputs(2501) <= (inputs(8)) or (inputs(136));
    layer0_outputs(2502) <= (inputs(148)) or (inputs(12));
    layer0_outputs(2503) <= inputs(159);
    layer0_outputs(2504) <= inputs(66);
    layer0_outputs(2505) <= (inputs(184)) and not (inputs(68));
    layer0_outputs(2506) <= not(inputs(70)) or (inputs(187));
    layer0_outputs(2507) <= '1';
    layer0_outputs(2508) <= not((inputs(74)) xor (inputs(90)));
    layer0_outputs(2509) <= inputs(229);
    layer0_outputs(2510) <= (inputs(52)) and not (inputs(128));
    layer0_outputs(2511) <= not(inputs(95)) or (inputs(72));
    layer0_outputs(2512) <= inputs(33);
    layer0_outputs(2513) <= not((inputs(131)) and (inputs(169)));
    layer0_outputs(2514) <= (inputs(199)) and not (inputs(112));
    layer0_outputs(2515) <= (inputs(161)) xor (inputs(121));
    layer0_outputs(2516) <= not(inputs(19));
    layer0_outputs(2517) <= (inputs(151)) xor (inputs(85));
    layer0_outputs(2518) <= (inputs(141)) and not (inputs(159));
    layer0_outputs(2519) <= not((inputs(238)) xor (inputs(150)));
    layer0_outputs(2520) <= '1';
    layer0_outputs(2521) <= not((inputs(123)) or (inputs(37)));
    layer0_outputs(2522) <= not((inputs(36)) or (inputs(36)));
    layer0_outputs(2523) <= not(inputs(132));
    layer0_outputs(2524) <= not((inputs(27)) xor (inputs(63)));
    layer0_outputs(2525) <= not(inputs(185)) or (inputs(69));
    layer0_outputs(2526) <= (inputs(160)) xor (inputs(24));
    layer0_outputs(2527) <= not(inputs(53));
    layer0_outputs(2528) <= (inputs(41)) and not (inputs(25));
    layer0_outputs(2529) <= (inputs(193)) or (inputs(83));
    layer0_outputs(2530) <= not(inputs(54)) or (inputs(10));
    layer0_outputs(2531) <= inputs(103);
    layer0_outputs(2532) <= inputs(220);
    layer0_outputs(2533) <= not((inputs(201)) or (inputs(194)));
    layer0_outputs(2534) <= not((inputs(12)) xor (inputs(169)));
    layer0_outputs(2535) <= (inputs(165)) xor (inputs(111));
    layer0_outputs(2536) <= (inputs(212)) xor (inputs(156));
    layer0_outputs(2537) <= (inputs(49)) or (inputs(94));
    layer0_outputs(2538) <= (inputs(100)) and not (inputs(159));
    layer0_outputs(2539) <= not(inputs(56)) or (inputs(108));
    layer0_outputs(2540) <= (inputs(94)) and (inputs(33));
    layer0_outputs(2541) <= not((inputs(47)) xor (inputs(153)));
    layer0_outputs(2542) <= not((inputs(112)) xor (inputs(170)));
    layer0_outputs(2543) <= not((inputs(111)) or (inputs(199)));
    layer0_outputs(2544) <= (inputs(98)) or (inputs(209));
    layer0_outputs(2545) <= not((inputs(79)) or (inputs(87)));
    layer0_outputs(2546) <= not((inputs(156)) or (inputs(155)));
    layer0_outputs(2547) <= not(inputs(28)) or (inputs(48));
    layer0_outputs(2548) <= (inputs(48)) or (inputs(107));
    layer0_outputs(2549) <= not(inputs(167)) or (inputs(145));
    layer0_outputs(2550) <= not(inputs(230)) or (inputs(242));
    layer0_outputs(2551) <= not(inputs(85));
    layer0_outputs(2552) <= not((inputs(26)) xor (inputs(23)));
    layer0_outputs(2553) <= not(inputs(205)) or (inputs(93));
    layer0_outputs(2554) <= not((inputs(108)) or (inputs(51)));
    layer0_outputs(2555) <= not(inputs(185)) or (inputs(204));
    layer0_outputs(2556) <= (inputs(52)) and not (inputs(205));
    layer0_outputs(2557) <= not((inputs(242)) xor (inputs(59)));
    layer0_outputs(2558) <= not((inputs(155)) or (inputs(78)));
    layer0_outputs(2559) <= (inputs(116)) and not (inputs(130));
    layer0_outputs(2560) <= (inputs(146)) xor (inputs(200));
    layer0_outputs(2561) <= (inputs(91)) and not (inputs(51));
    layer0_outputs(2562) <= not(inputs(211));
    layer0_outputs(2563) <= not(inputs(49)) or (inputs(20));
    layer0_outputs(2564) <= (inputs(148)) or (inputs(253));
    layer0_outputs(2565) <= (inputs(38)) and not (inputs(129));
    layer0_outputs(2566) <= (inputs(45)) or (inputs(93));
    layer0_outputs(2567) <= not((inputs(201)) xor (inputs(17)));
    layer0_outputs(2568) <= not(inputs(83));
    layer0_outputs(2569) <= not(inputs(168)) or (inputs(116));
    layer0_outputs(2570) <= not(inputs(133)) or (inputs(159));
    layer0_outputs(2571) <= inputs(112);
    layer0_outputs(2572) <= not(inputs(133));
    layer0_outputs(2573) <= not((inputs(247)) xor (inputs(75)));
    layer0_outputs(2574) <= (inputs(223)) xor (inputs(215));
    layer0_outputs(2575) <= (inputs(225)) xor (inputs(239));
    layer0_outputs(2576) <= not(inputs(149)) or (inputs(230));
    layer0_outputs(2577) <= not(inputs(152));
    layer0_outputs(2578) <= not(inputs(42)) or (inputs(46));
    layer0_outputs(2579) <= not((inputs(25)) or (inputs(206)));
    layer0_outputs(2580) <= (inputs(152)) or (inputs(107));
    layer0_outputs(2581) <= not(inputs(222)) or (inputs(193));
    layer0_outputs(2582) <= (inputs(133)) and (inputs(107));
    layer0_outputs(2583) <= inputs(124);
    layer0_outputs(2584) <= not((inputs(49)) or (inputs(128)));
    layer0_outputs(2585) <= (inputs(199)) xor (inputs(178));
    layer0_outputs(2586) <= not(inputs(164)) or (inputs(29));
    layer0_outputs(2587) <= (inputs(171)) or (inputs(170));
    layer0_outputs(2588) <= (inputs(211)) or (inputs(90));
    layer0_outputs(2589) <= not((inputs(175)) xor (inputs(107)));
    layer0_outputs(2590) <= not((inputs(90)) or (inputs(194)));
    layer0_outputs(2591) <= (inputs(167)) and not (inputs(78));
    layer0_outputs(2592) <= not((inputs(129)) or (inputs(128)));
    layer0_outputs(2593) <= not(inputs(30));
    layer0_outputs(2594) <= not(inputs(133)) or (inputs(178));
    layer0_outputs(2595) <= not(inputs(230));
    layer0_outputs(2596) <= (inputs(91)) and not (inputs(242));
    layer0_outputs(2597) <= (inputs(124)) and (inputs(122));
    layer0_outputs(2598) <= not(inputs(195)) or (inputs(107));
    layer0_outputs(2599) <= (inputs(68)) and not (inputs(176));
    layer0_outputs(2600) <= not(inputs(151)) or (inputs(145));
    layer0_outputs(2601) <= not(inputs(106)) or (inputs(214));
    layer0_outputs(2602) <= not((inputs(141)) or (inputs(124)));
    layer0_outputs(2603) <= inputs(64);
    layer0_outputs(2604) <= not((inputs(158)) xor (inputs(161)));
    layer0_outputs(2605) <= inputs(95);
    layer0_outputs(2606) <= not(inputs(229));
    layer0_outputs(2607) <= '0';
    layer0_outputs(2608) <= not((inputs(91)) or (inputs(60)));
    layer0_outputs(2609) <= (inputs(216)) and not (inputs(248));
    layer0_outputs(2610) <= inputs(61);
    layer0_outputs(2611) <= not(inputs(152)) or (inputs(238));
    layer0_outputs(2612) <= not(inputs(45));
    layer0_outputs(2613) <= (inputs(105)) and not (inputs(52));
    layer0_outputs(2614) <= not(inputs(149)) or (inputs(234));
    layer0_outputs(2615) <= not((inputs(59)) or (inputs(185)));
    layer0_outputs(2616) <= not(inputs(235)) or (inputs(11));
    layer0_outputs(2617) <= not(inputs(120)) or (inputs(16));
    layer0_outputs(2618) <= (inputs(168)) or (inputs(7));
    layer0_outputs(2619) <= not((inputs(55)) or (inputs(107)));
    layer0_outputs(2620) <= not((inputs(69)) xor (inputs(8)));
    layer0_outputs(2621) <= (inputs(214)) and not (inputs(237));
    layer0_outputs(2622) <= not(inputs(57));
    layer0_outputs(2623) <= (inputs(119)) xor (inputs(100));
    layer0_outputs(2624) <= not((inputs(54)) xor (inputs(199)));
    layer0_outputs(2625) <= not(inputs(149));
    layer0_outputs(2626) <= (inputs(169)) and not (inputs(194));
    layer0_outputs(2627) <= not(inputs(28));
    layer0_outputs(2628) <= not(inputs(232));
    layer0_outputs(2629) <= not((inputs(128)) or (inputs(151)));
    layer0_outputs(2630) <= '0';
    layer0_outputs(2631) <= (inputs(196)) xor (inputs(159));
    layer0_outputs(2632) <= (inputs(237)) or (inputs(94));
    layer0_outputs(2633) <= not(inputs(248));
    layer0_outputs(2634) <= not(inputs(163)) or (inputs(235));
    layer0_outputs(2635) <= (inputs(37)) and not (inputs(213));
    layer0_outputs(2636) <= not((inputs(101)) xor (inputs(98)));
    layer0_outputs(2637) <= not((inputs(84)) xor (inputs(255)));
    layer0_outputs(2638) <= '1';
    layer0_outputs(2639) <= (inputs(245)) and not (inputs(42));
    layer0_outputs(2640) <= (inputs(67)) or (inputs(114));
    layer0_outputs(2641) <= (inputs(171)) xor (inputs(181));
    layer0_outputs(2642) <= (inputs(229)) and not (inputs(192));
    layer0_outputs(2643) <= (inputs(124)) or (inputs(35));
    layer0_outputs(2644) <= (inputs(216)) or (inputs(90));
    layer0_outputs(2645) <= (inputs(152)) xor (inputs(212));
    layer0_outputs(2646) <= inputs(101);
    layer0_outputs(2647) <= not((inputs(99)) xor (inputs(128)));
    layer0_outputs(2648) <= inputs(161);
    layer0_outputs(2649) <= not(inputs(172)) or (inputs(210));
    layer0_outputs(2650) <= (inputs(146)) or (inputs(192));
    layer0_outputs(2651) <= not(inputs(57)) or (inputs(130));
    layer0_outputs(2652) <= not(inputs(88)) or (inputs(241));
    layer0_outputs(2653) <= not(inputs(39)) or (inputs(46));
    layer0_outputs(2654) <= not(inputs(12));
    layer0_outputs(2655) <= (inputs(66)) or (inputs(63));
    layer0_outputs(2656) <= (inputs(154)) and not (inputs(115));
    layer0_outputs(2657) <= (inputs(47)) and not (inputs(112));
    layer0_outputs(2658) <= not((inputs(255)) or (inputs(99)));
    layer0_outputs(2659) <= inputs(72);
    layer0_outputs(2660) <= not(inputs(125));
    layer0_outputs(2661) <= not(inputs(4));
    layer0_outputs(2662) <= (inputs(252)) and not (inputs(115));
    layer0_outputs(2663) <= not((inputs(26)) or (inputs(124)));
    layer0_outputs(2664) <= (inputs(54)) and not (inputs(205));
    layer0_outputs(2665) <= not(inputs(204));
    layer0_outputs(2666) <= (inputs(222)) and (inputs(49));
    layer0_outputs(2667) <= not(inputs(230));
    layer0_outputs(2668) <= not((inputs(35)) or (inputs(229)));
    layer0_outputs(2669) <= not((inputs(117)) or (inputs(21)));
    layer0_outputs(2670) <= not((inputs(36)) or (inputs(71)));
    layer0_outputs(2671) <= not((inputs(250)) xor (inputs(204)));
    layer0_outputs(2672) <= (inputs(168)) xor (inputs(244));
    layer0_outputs(2673) <= (inputs(138)) and not (inputs(60));
    layer0_outputs(2674) <= (inputs(100)) or (inputs(207));
    layer0_outputs(2675) <= '0';
    layer0_outputs(2676) <= not((inputs(52)) or (inputs(68)));
    layer0_outputs(2677) <= inputs(235);
    layer0_outputs(2678) <= not((inputs(34)) xor (inputs(237)));
    layer0_outputs(2679) <= not((inputs(105)) xor (inputs(76)));
    layer0_outputs(2680) <= (inputs(169)) and not (inputs(254));
    layer0_outputs(2681) <= not((inputs(95)) xor (inputs(191)));
    layer0_outputs(2682) <= not((inputs(68)) xor (inputs(108)));
    layer0_outputs(2683) <= not((inputs(188)) or (inputs(10)));
    layer0_outputs(2684) <= not((inputs(194)) or (inputs(238)));
    layer0_outputs(2685) <= (inputs(115)) or (inputs(54));
    layer0_outputs(2686) <= inputs(106);
    layer0_outputs(2687) <= (inputs(209)) or (inputs(24));
    layer0_outputs(2688) <= not(inputs(165)) or (inputs(96));
    layer0_outputs(2689) <= inputs(102);
    layer0_outputs(2690) <= not((inputs(242)) and (inputs(145)));
    layer0_outputs(2691) <= inputs(55);
    layer0_outputs(2692) <= not((inputs(134)) xor (inputs(217)));
    layer0_outputs(2693) <= not((inputs(198)) or (inputs(182)));
    layer0_outputs(2694) <= not((inputs(209)) xor (inputs(112)));
    layer0_outputs(2695) <= not(inputs(42)) or (inputs(11));
    layer0_outputs(2696) <= (inputs(216)) and not (inputs(45));
    layer0_outputs(2697) <= (inputs(42)) xor (inputs(107));
    layer0_outputs(2698) <= not((inputs(82)) or (inputs(91)));
    layer0_outputs(2699) <= not((inputs(233)) xor (inputs(195)));
    layer0_outputs(2700) <= not(inputs(148));
    layer0_outputs(2701) <= (inputs(216)) and not (inputs(58));
    layer0_outputs(2702) <= (inputs(59)) and not (inputs(31));
    layer0_outputs(2703) <= not(inputs(135)) or (inputs(231));
    layer0_outputs(2704) <= not((inputs(253)) xor (inputs(134)));
    layer0_outputs(2705) <= (inputs(164)) or (inputs(123));
    layer0_outputs(2706) <= inputs(10);
    layer0_outputs(2707) <= not(inputs(235));
    layer0_outputs(2708) <= not((inputs(128)) or (inputs(156)));
    layer0_outputs(2709) <= not(inputs(65));
    layer0_outputs(2710) <= (inputs(22)) xor (inputs(238));
    layer0_outputs(2711) <= not((inputs(35)) or (inputs(91)));
    layer0_outputs(2712) <= (inputs(123)) xor (inputs(160));
    layer0_outputs(2713) <= not(inputs(10));
    layer0_outputs(2714) <= inputs(8);
    layer0_outputs(2715) <= (inputs(109)) or (inputs(112));
    layer0_outputs(2716) <= not(inputs(23)) or (inputs(7));
    layer0_outputs(2717) <= not((inputs(62)) or (inputs(234)));
    layer0_outputs(2718) <= not(inputs(176));
    layer0_outputs(2719) <= inputs(241);
    layer0_outputs(2720) <= not((inputs(137)) xor (inputs(206)));
    layer0_outputs(2721) <= (inputs(19)) xor (inputs(242));
    layer0_outputs(2722) <= inputs(125);
    layer0_outputs(2723) <= (inputs(37)) and not (inputs(41));
    layer0_outputs(2724) <= inputs(49);
    layer0_outputs(2725) <= inputs(164);
    layer0_outputs(2726) <= not(inputs(204));
    layer0_outputs(2727) <= not((inputs(206)) or (inputs(183)));
    layer0_outputs(2728) <= not(inputs(15));
    layer0_outputs(2729) <= inputs(141);
    layer0_outputs(2730) <= not((inputs(13)) or (inputs(88)));
    layer0_outputs(2731) <= (inputs(57)) xor (inputs(183));
    layer0_outputs(2732) <= inputs(55);
    layer0_outputs(2733) <= (inputs(89)) and not (inputs(14));
    layer0_outputs(2734) <= not((inputs(2)) or (inputs(14)));
    layer0_outputs(2735) <= not((inputs(192)) xor (inputs(178)));
    layer0_outputs(2736) <= (inputs(178)) or (inputs(128));
    layer0_outputs(2737) <= not((inputs(240)) or (inputs(196)));
    layer0_outputs(2738) <= not(inputs(166));
    layer0_outputs(2739) <= (inputs(5)) xor (inputs(111));
    layer0_outputs(2740) <= (inputs(237)) and not (inputs(62));
    layer0_outputs(2741) <= (inputs(191)) or (inputs(15));
    layer0_outputs(2742) <= (inputs(111)) or (inputs(25));
    layer0_outputs(2743) <= (inputs(123)) and not (inputs(174));
    layer0_outputs(2744) <= not(inputs(60)) or (inputs(51));
    layer0_outputs(2745) <= (inputs(25)) or (inputs(167));
    layer0_outputs(2746) <= not((inputs(71)) xor (inputs(96)));
    layer0_outputs(2747) <= (inputs(100)) xor (inputs(179));
    layer0_outputs(2748) <= inputs(196);
    layer0_outputs(2749) <= not((inputs(172)) or (inputs(29)));
    layer0_outputs(2750) <= (inputs(45)) or (inputs(219));
    layer0_outputs(2751) <= not((inputs(54)) or (inputs(37)));
    layer0_outputs(2752) <= not(inputs(107)) or (inputs(158));
    layer0_outputs(2753) <= not(inputs(40)) or (inputs(8));
    layer0_outputs(2754) <= inputs(119);
    layer0_outputs(2755) <= (inputs(218)) or (inputs(203));
    layer0_outputs(2756) <= not((inputs(54)) xor (inputs(87)));
    layer0_outputs(2757) <= (inputs(154)) or (inputs(142));
    layer0_outputs(2758) <= inputs(247);
    layer0_outputs(2759) <= not(inputs(198));
    layer0_outputs(2760) <= not(inputs(199)) or (inputs(226));
    layer0_outputs(2761) <= '1';
    layer0_outputs(2762) <= not((inputs(104)) or (inputs(104)));
    layer0_outputs(2763) <= (inputs(212)) and not (inputs(249));
    layer0_outputs(2764) <= (inputs(72)) xor (inputs(250));
    layer0_outputs(2765) <= not((inputs(204)) or (inputs(65)));
    layer0_outputs(2766) <= not(inputs(164));
    layer0_outputs(2767) <= '1';
    layer0_outputs(2768) <= inputs(151);
    layer0_outputs(2769) <= (inputs(29)) or (inputs(113));
    layer0_outputs(2770) <= '1';
    layer0_outputs(2771) <= not((inputs(62)) and (inputs(16)));
    layer0_outputs(2772) <= (inputs(219)) or (inputs(18));
    layer0_outputs(2773) <= inputs(212);
    layer0_outputs(2774) <= (inputs(184)) and not (inputs(73));
    layer0_outputs(2775) <= (inputs(63)) xor (inputs(130));
    layer0_outputs(2776) <= (inputs(88)) or (inputs(108));
    layer0_outputs(2777) <= not(inputs(248)) or (inputs(236));
    layer0_outputs(2778) <= not((inputs(240)) xor (inputs(181)));
    layer0_outputs(2779) <= (inputs(46)) or (inputs(167));
    layer0_outputs(2780) <= inputs(148);
    layer0_outputs(2781) <= inputs(74);
    layer0_outputs(2782) <= (inputs(76)) or (inputs(19));
    layer0_outputs(2783) <= not(inputs(198));
    layer0_outputs(2784) <= (inputs(222)) xor (inputs(59));
    layer0_outputs(2785) <= (inputs(130)) or (inputs(218));
    layer0_outputs(2786) <= not(inputs(246)) or (inputs(34));
    layer0_outputs(2787) <= not((inputs(27)) xor (inputs(131)));
    layer0_outputs(2788) <= not(inputs(112));
    layer0_outputs(2789) <= (inputs(153)) or (inputs(187));
    layer0_outputs(2790) <= (inputs(104)) or (inputs(233));
    layer0_outputs(2791) <= (inputs(45)) and not (inputs(146));
    layer0_outputs(2792) <= not(inputs(10));
    layer0_outputs(2793) <= (inputs(44)) and not (inputs(226));
    layer0_outputs(2794) <= not(inputs(205)) or (inputs(211));
    layer0_outputs(2795) <= not(inputs(249)) or (inputs(141));
    layer0_outputs(2796) <= (inputs(78)) and (inputs(155));
    layer0_outputs(2797) <= not((inputs(254)) and (inputs(146)));
    layer0_outputs(2798) <= not(inputs(251));
    layer0_outputs(2799) <= not((inputs(25)) or (inputs(34)));
    layer0_outputs(2800) <= not(inputs(115));
    layer0_outputs(2801) <= (inputs(4)) and (inputs(94));
    layer0_outputs(2802) <= (inputs(61)) xor (inputs(90));
    layer0_outputs(2803) <= not((inputs(7)) or (inputs(197)));
    layer0_outputs(2804) <= '0';
    layer0_outputs(2805) <= not(inputs(215));
    layer0_outputs(2806) <= not(inputs(106));
    layer0_outputs(2807) <= (inputs(87)) and not (inputs(50));
    layer0_outputs(2808) <= not(inputs(105));
    layer0_outputs(2809) <= (inputs(67)) or (inputs(134));
    layer0_outputs(2810) <= not((inputs(170)) and (inputs(46)));
    layer0_outputs(2811) <= inputs(54);
    layer0_outputs(2812) <= not((inputs(250)) xor (inputs(111)));
    layer0_outputs(2813) <= not((inputs(249)) xor (inputs(209)));
    layer0_outputs(2814) <= not((inputs(250)) or (inputs(164)));
    layer0_outputs(2815) <= not(inputs(51));
    layer0_outputs(2816) <= not(inputs(230));
    layer0_outputs(2817) <= not((inputs(69)) or (inputs(108)));
    layer0_outputs(2818) <= (inputs(179)) xor (inputs(181));
    layer0_outputs(2819) <= not(inputs(183)) or (inputs(240));
    layer0_outputs(2820) <= not((inputs(180)) or (inputs(144)));
    layer0_outputs(2821) <= not((inputs(146)) xor (inputs(184)));
    layer0_outputs(2822) <= not((inputs(173)) or (inputs(151)));
    layer0_outputs(2823) <= not((inputs(249)) or (inputs(184)));
    layer0_outputs(2824) <= inputs(41);
    layer0_outputs(2825) <= not((inputs(140)) xor (inputs(19)));
    layer0_outputs(2826) <= not((inputs(69)) xor (inputs(244)));
    layer0_outputs(2827) <= (inputs(69)) or (inputs(77));
    layer0_outputs(2828) <= not(inputs(152));
    layer0_outputs(2829) <= not(inputs(209));
    layer0_outputs(2830) <= (inputs(43)) xor (inputs(203));
    layer0_outputs(2831) <= not((inputs(122)) or (inputs(36)));
    layer0_outputs(2832) <= (inputs(36)) and not (inputs(122));
    layer0_outputs(2833) <= not(inputs(100));
    layer0_outputs(2834) <= (inputs(64)) xor (inputs(212));
    layer0_outputs(2835) <= not(inputs(212));
    layer0_outputs(2836) <= inputs(141);
    layer0_outputs(2837) <= not((inputs(11)) or (inputs(33)));
    layer0_outputs(2838) <= (inputs(156)) and not (inputs(157));
    layer0_outputs(2839) <= inputs(135);
    layer0_outputs(2840) <= not(inputs(139));
    layer0_outputs(2841) <= not(inputs(156)) or (inputs(219));
    layer0_outputs(2842) <= not(inputs(176)) or (inputs(81));
    layer0_outputs(2843) <= not(inputs(167)) or (inputs(33));
    layer0_outputs(2844) <= (inputs(212)) and not (inputs(64));
    layer0_outputs(2845) <= not((inputs(36)) or (inputs(52)));
    layer0_outputs(2846) <= not((inputs(196)) xor (inputs(42)));
    layer0_outputs(2847) <= not((inputs(15)) xor (inputs(153)));
    layer0_outputs(2848) <= not((inputs(58)) or (inputs(232)));
    layer0_outputs(2849) <= not((inputs(121)) xor (inputs(48)));
    layer0_outputs(2850) <= not((inputs(116)) or (inputs(255)));
    layer0_outputs(2851) <= not(inputs(146));
    layer0_outputs(2852) <= (inputs(205)) or (inputs(237));
    layer0_outputs(2853) <= inputs(245);
    layer0_outputs(2854) <= '0';
    layer0_outputs(2855) <= (inputs(193)) and not (inputs(162));
    layer0_outputs(2856) <= (inputs(40)) or (inputs(42));
    layer0_outputs(2857) <= not(inputs(125));
    layer0_outputs(2858) <= (inputs(205)) xor (inputs(237));
    layer0_outputs(2859) <= (inputs(97)) or (inputs(90));
    layer0_outputs(2860) <= inputs(47);
    layer0_outputs(2861) <= not((inputs(76)) xor (inputs(188)));
    layer0_outputs(2862) <= not(inputs(122));
    layer0_outputs(2863) <= not((inputs(43)) xor (inputs(133)));
    layer0_outputs(2864) <= (inputs(136)) and not (inputs(181));
    layer0_outputs(2865) <= not(inputs(120)) or (inputs(109));
    layer0_outputs(2866) <= not((inputs(175)) or (inputs(105)));
    layer0_outputs(2867) <= inputs(24);
    layer0_outputs(2868) <= inputs(157);
    layer0_outputs(2869) <= (inputs(86)) xor (inputs(238));
    layer0_outputs(2870) <= not(inputs(10)) or (inputs(99));
    layer0_outputs(2871) <= not(inputs(129)) or (inputs(11));
    layer0_outputs(2872) <= not((inputs(222)) xor (inputs(48)));
    layer0_outputs(2873) <= (inputs(235)) and not (inputs(224));
    layer0_outputs(2874) <= not(inputs(75));
    layer0_outputs(2875) <= inputs(6);
    layer0_outputs(2876) <= not((inputs(248)) and (inputs(213)));
    layer0_outputs(2877) <= not(inputs(149)) or (inputs(178));
    layer0_outputs(2878) <= not(inputs(101)) or (inputs(240));
    layer0_outputs(2879) <= inputs(35);
    layer0_outputs(2880) <= inputs(190);
    layer0_outputs(2881) <= not(inputs(106)) or (inputs(189));
    layer0_outputs(2882) <= not((inputs(252)) or (inputs(152)));
    layer0_outputs(2883) <= not((inputs(1)) or (inputs(59)));
    layer0_outputs(2884) <= '0';
    layer0_outputs(2885) <= (inputs(105)) or (inputs(154));
    layer0_outputs(2886) <= (inputs(192)) xor (inputs(16));
    layer0_outputs(2887) <= not((inputs(208)) or (inputs(40)));
    layer0_outputs(2888) <= inputs(40);
    layer0_outputs(2889) <= (inputs(199)) xor (inputs(207));
    layer0_outputs(2890) <= not((inputs(146)) and (inputs(224)));
    layer0_outputs(2891) <= not(inputs(170));
    layer0_outputs(2892) <= not(inputs(151));
    layer0_outputs(2893) <= (inputs(181)) and not (inputs(66));
    layer0_outputs(2894) <= not((inputs(221)) xor (inputs(168)));
    layer0_outputs(2895) <= not(inputs(191)) or (inputs(238));
    layer0_outputs(2896) <= not(inputs(78)) or (inputs(203));
    layer0_outputs(2897) <= (inputs(144)) xor (inputs(13));
    layer0_outputs(2898) <= not((inputs(176)) and (inputs(5)));
    layer0_outputs(2899) <= not(inputs(41)) or (inputs(27));
    layer0_outputs(2900) <= (inputs(216)) and not (inputs(45));
    layer0_outputs(2901) <= (inputs(28)) or (inputs(169));
    layer0_outputs(2902) <= (inputs(164)) or (inputs(67));
    layer0_outputs(2903) <= inputs(203);
    layer0_outputs(2904) <= not(inputs(27)) or (inputs(211));
    layer0_outputs(2905) <= (inputs(180)) xor (inputs(161));
    layer0_outputs(2906) <= not(inputs(102)) or (inputs(18));
    layer0_outputs(2907) <= (inputs(196)) and not (inputs(64));
    layer0_outputs(2908) <= not(inputs(44));
    layer0_outputs(2909) <= inputs(37);
    layer0_outputs(2910) <= not(inputs(202));
    layer0_outputs(2911) <= inputs(13);
    layer0_outputs(2912) <= not((inputs(202)) or (inputs(221)));
    layer0_outputs(2913) <= not(inputs(84)) or (inputs(67));
    layer0_outputs(2914) <= not((inputs(110)) or (inputs(164)));
    layer0_outputs(2915) <= not(inputs(70)) or (inputs(206));
    layer0_outputs(2916) <= not(inputs(67));
    layer0_outputs(2917) <= not((inputs(1)) and (inputs(14)));
    layer0_outputs(2918) <= not((inputs(165)) or (inputs(141)));
    layer0_outputs(2919) <= inputs(222);
    layer0_outputs(2920) <= inputs(162);
    layer0_outputs(2921) <= (inputs(97)) and not (inputs(115));
    layer0_outputs(2922) <= not((inputs(154)) or (inputs(66)));
    layer0_outputs(2923) <= (inputs(28)) xor (inputs(100));
    layer0_outputs(2924) <= not(inputs(254));
    layer0_outputs(2925) <= not(inputs(165)) or (inputs(71));
    layer0_outputs(2926) <= (inputs(228)) and not (inputs(189));
    layer0_outputs(2927) <= (inputs(149)) and not (inputs(35));
    layer0_outputs(2928) <= (inputs(145)) xor (inputs(239));
    layer0_outputs(2929) <= not(inputs(88)) or (inputs(57));
    layer0_outputs(2930) <= not(inputs(56)) or (inputs(9));
    layer0_outputs(2931) <= not(inputs(39));
    layer0_outputs(2932) <= (inputs(142)) xor (inputs(199));
    layer0_outputs(2933) <= not(inputs(91));
    layer0_outputs(2934) <= (inputs(254)) and (inputs(197));
    layer0_outputs(2935) <= inputs(164);
    layer0_outputs(2936) <= not((inputs(156)) xor (inputs(175)));
    layer0_outputs(2937) <= not(inputs(91)) or (inputs(125));
    layer0_outputs(2938) <= (inputs(200)) or (inputs(26));
    layer0_outputs(2939) <= (inputs(106)) and not (inputs(118));
    layer0_outputs(2940) <= not((inputs(108)) or (inputs(118)));
    layer0_outputs(2941) <= (inputs(56)) xor (inputs(120));
    layer0_outputs(2942) <= (inputs(182)) and not (inputs(153));
    layer0_outputs(2943) <= not((inputs(70)) or (inputs(39)));
    layer0_outputs(2944) <= not(inputs(115));
    layer0_outputs(2945) <= inputs(86);
    layer0_outputs(2946) <= inputs(150);
    layer0_outputs(2947) <= inputs(162);
    layer0_outputs(2948) <= inputs(99);
    layer0_outputs(2949) <= not((inputs(82)) xor (inputs(15)));
    layer0_outputs(2950) <= (inputs(136)) and not (inputs(171));
    layer0_outputs(2951) <= not((inputs(86)) and (inputs(81)));
    layer0_outputs(2952) <= '0';
    layer0_outputs(2953) <= not(inputs(73)) or (inputs(237));
    layer0_outputs(2954) <= (inputs(81)) or (inputs(89));
    layer0_outputs(2955) <= not((inputs(207)) or (inputs(222)));
    layer0_outputs(2956) <= not(inputs(104));
    layer0_outputs(2957) <= not((inputs(35)) or (inputs(196)));
    layer0_outputs(2958) <= not((inputs(215)) or (inputs(180)));
    layer0_outputs(2959) <= (inputs(216)) xor (inputs(96));
    layer0_outputs(2960) <= inputs(137);
    layer0_outputs(2961) <= not((inputs(29)) xor (inputs(205)));
    layer0_outputs(2962) <= not(inputs(26)) or (inputs(1));
    layer0_outputs(2963) <= (inputs(61)) or (inputs(240));
    layer0_outputs(2964) <= (inputs(57)) and not (inputs(64));
    layer0_outputs(2965) <= inputs(142);
    layer0_outputs(2966) <= inputs(66);
    layer0_outputs(2967) <= inputs(167);
    layer0_outputs(2968) <= (inputs(250)) and not (inputs(59));
    layer0_outputs(2969) <= not(inputs(118));
    layer0_outputs(2970) <= not((inputs(16)) xor (inputs(70)));
    layer0_outputs(2971) <= not(inputs(133));
    layer0_outputs(2972) <= not(inputs(206));
    layer0_outputs(2973) <= '1';
    layer0_outputs(2974) <= not(inputs(200)) or (inputs(89));
    layer0_outputs(2975) <= not(inputs(197));
    layer0_outputs(2976) <= not((inputs(55)) or (inputs(155)));
    layer0_outputs(2977) <= not(inputs(201));
    layer0_outputs(2978) <= (inputs(27)) and (inputs(58));
    layer0_outputs(2979) <= not((inputs(95)) xor (inputs(146)));
    layer0_outputs(2980) <= (inputs(159)) or (inputs(154));
    layer0_outputs(2981) <= not((inputs(106)) or (inputs(156)));
    layer0_outputs(2982) <= not(inputs(152));
    layer0_outputs(2983) <= (inputs(147)) xor (inputs(118));
    layer0_outputs(2984) <= not((inputs(41)) xor (inputs(207)));
    layer0_outputs(2985) <= (inputs(222)) xor (inputs(157));
    layer0_outputs(2986) <= not(inputs(9));
    layer0_outputs(2987) <= (inputs(88)) and not (inputs(123));
    layer0_outputs(2988) <= not(inputs(39)) or (inputs(111));
    layer0_outputs(2989) <= '1';
    layer0_outputs(2990) <= '0';
    layer0_outputs(2991) <= inputs(220);
    layer0_outputs(2992) <= (inputs(206)) xor (inputs(105));
    layer0_outputs(2993) <= (inputs(221)) or (inputs(44));
    layer0_outputs(2994) <= not((inputs(10)) or (inputs(214)));
    layer0_outputs(2995) <= (inputs(57)) and not (inputs(84));
    layer0_outputs(2996) <= not(inputs(78));
    layer0_outputs(2997) <= (inputs(80)) and not (inputs(65));
    layer0_outputs(2998) <= not(inputs(31)) or (inputs(143));
    layer0_outputs(2999) <= not(inputs(101)) or (inputs(157));
    layer0_outputs(3000) <= (inputs(232)) and not (inputs(164));
    layer0_outputs(3001) <= inputs(101);
    layer0_outputs(3002) <= (inputs(23)) xor (inputs(39));
    layer0_outputs(3003) <= not(inputs(50)) or (inputs(174));
    layer0_outputs(3004) <= not(inputs(68));
    layer0_outputs(3005) <= (inputs(143)) and not (inputs(248));
    layer0_outputs(3006) <= not(inputs(197)) or (inputs(169));
    layer0_outputs(3007) <= not((inputs(179)) or (inputs(148)));
    layer0_outputs(3008) <= inputs(77);
    layer0_outputs(3009) <= inputs(140);
    layer0_outputs(3010) <= inputs(42);
    layer0_outputs(3011) <= not(inputs(115)) or (inputs(11));
    layer0_outputs(3012) <= not(inputs(114)) or (inputs(80));
    layer0_outputs(3013) <= not(inputs(45)) or (inputs(113));
    layer0_outputs(3014) <= inputs(176);
    layer0_outputs(3015) <= (inputs(108)) xor (inputs(186));
    layer0_outputs(3016) <= not((inputs(135)) and (inputs(213)));
    layer0_outputs(3017) <= (inputs(214)) and not (inputs(204));
    layer0_outputs(3018) <= inputs(178);
    layer0_outputs(3019) <= (inputs(182)) xor (inputs(127));
    layer0_outputs(3020) <= not(inputs(96));
    layer0_outputs(3021) <= not(inputs(53));
    layer0_outputs(3022) <= not((inputs(184)) or (inputs(160)));
    layer0_outputs(3023) <= inputs(151);
    layer0_outputs(3024) <= (inputs(160)) or (inputs(197));
    layer0_outputs(3025) <= not((inputs(68)) or (inputs(173)));
    layer0_outputs(3026) <= inputs(108);
    layer0_outputs(3027) <= not((inputs(26)) xor (inputs(241)));
    layer0_outputs(3028) <= not((inputs(154)) xor (inputs(185)));
    layer0_outputs(3029) <= (inputs(233)) or (inputs(122));
    layer0_outputs(3030) <= (inputs(248)) and (inputs(78));
    layer0_outputs(3031) <= (inputs(183)) or (inputs(175));
    layer0_outputs(3032) <= not(inputs(124)) or (inputs(98));
    layer0_outputs(3033) <= (inputs(176)) and not (inputs(196));
    layer0_outputs(3034) <= not((inputs(103)) xor (inputs(218)));
    layer0_outputs(3035) <= not(inputs(108));
    layer0_outputs(3036) <= (inputs(63)) and not (inputs(29));
    layer0_outputs(3037) <= not((inputs(80)) and (inputs(113)));
    layer0_outputs(3038) <= (inputs(16)) and not (inputs(67));
    layer0_outputs(3039) <= (inputs(63)) and (inputs(208));
    layer0_outputs(3040) <= (inputs(216)) or (inputs(165));
    layer0_outputs(3041) <= not((inputs(166)) or (inputs(82)));
    layer0_outputs(3042) <= inputs(123);
    layer0_outputs(3043) <= not(inputs(238));
    layer0_outputs(3044) <= (inputs(20)) xor (inputs(60));
    layer0_outputs(3045) <= not((inputs(255)) xor (inputs(169)));
    layer0_outputs(3046) <= not((inputs(50)) xor (inputs(246)));
    layer0_outputs(3047) <= not(inputs(173));
    layer0_outputs(3048) <= not((inputs(211)) or (inputs(90)));
    layer0_outputs(3049) <= (inputs(217)) or (inputs(236));
    layer0_outputs(3050) <= inputs(182);
    layer0_outputs(3051) <= (inputs(75)) and not (inputs(47));
    layer0_outputs(3052) <= (inputs(130)) and not (inputs(86));
    layer0_outputs(3053) <= '1';
    layer0_outputs(3054) <= not(inputs(217)) or (inputs(51));
    layer0_outputs(3055) <= (inputs(135)) or (inputs(235));
    layer0_outputs(3056) <= not(inputs(98));
    layer0_outputs(3057) <= (inputs(229)) and not (inputs(128));
    layer0_outputs(3058) <= not(inputs(24)) or (inputs(146));
    layer0_outputs(3059) <= inputs(184);
    layer0_outputs(3060) <= inputs(103);
    layer0_outputs(3061) <= not(inputs(12)) or (inputs(126));
    layer0_outputs(3062) <= '1';
    layer0_outputs(3063) <= not(inputs(94));
    layer0_outputs(3064) <= (inputs(33)) xor (inputs(86));
    layer0_outputs(3065) <= not((inputs(254)) xor (inputs(123)));
    layer0_outputs(3066) <= inputs(241);
    layer0_outputs(3067) <= inputs(164);
    layer0_outputs(3068) <= (inputs(237)) or (inputs(119));
    layer0_outputs(3069) <= not((inputs(51)) or (inputs(153)));
    layer0_outputs(3070) <= (inputs(49)) or (inputs(151));
    layer0_outputs(3071) <= inputs(209);
    layer0_outputs(3072) <= (inputs(247)) or (inputs(237));
    layer0_outputs(3073) <= not(inputs(68)) or (inputs(207));
    layer0_outputs(3074) <= (inputs(137)) xor (inputs(1));
    layer0_outputs(3075) <= not(inputs(58)) or (inputs(98));
    layer0_outputs(3076) <= (inputs(147)) and not (inputs(36));
    layer0_outputs(3077) <= not(inputs(193));
    layer0_outputs(3078) <= (inputs(186)) and not (inputs(54));
    layer0_outputs(3079) <= (inputs(227)) or (inputs(228));
    layer0_outputs(3080) <= (inputs(15)) xor (inputs(1));
    layer0_outputs(3081) <= not(inputs(78)) or (inputs(36));
    layer0_outputs(3082) <= not((inputs(92)) or (inputs(211)));
    layer0_outputs(3083) <= not(inputs(93)) or (inputs(111));
    layer0_outputs(3084) <= inputs(70);
    layer0_outputs(3085) <= (inputs(74)) xor (inputs(246));
    layer0_outputs(3086) <= not(inputs(90)) or (inputs(239));
    layer0_outputs(3087) <= not(inputs(197)) or (inputs(227));
    layer0_outputs(3088) <= not((inputs(62)) and (inputs(145)));
    layer0_outputs(3089) <= '0';
    layer0_outputs(3090) <= not(inputs(137));
    layer0_outputs(3091) <= (inputs(110)) or (inputs(158));
    layer0_outputs(3092) <= (inputs(185)) and (inputs(146));
    layer0_outputs(3093) <= not(inputs(156));
    layer0_outputs(3094) <= (inputs(227)) or (inputs(137));
    layer0_outputs(3095) <= not(inputs(173)) or (inputs(225));
    layer0_outputs(3096) <= not(inputs(151));
    layer0_outputs(3097) <= not((inputs(94)) or (inputs(199)));
    layer0_outputs(3098) <= (inputs(142)) and not (inputs(85));
    layer0_outputs(3099) <= (inputs(73)) or (inputs(37));
    layer0_outputs(3100) <= (inputs(244)) or (inputs(162));
    layer0_outputs(3101) <= not((inputs(117)) or (inputs(46)));
    layer0_outputs(3102) <= not(inputs(72));
    layer0_outputs(3103) <= inputs(211);
    layer0_outputs(3104) <= not(inputs(228)) or (inputs(159));
    layer0_outputs(3105) <= not(inputs(121)) or (inputs(141));
    layer0_outputs(3106) <= (inputs(84)) xor (inputs(199));
    layer0_outputs(3107) <= '0';
    layer0_outputs(3108) <= inputs(121);
    layer0_outputs(3109) <= not(inputs(176)) or (inputs(45));
    layer0_outputs(3110) <= not(inputs(168)) or (inputs(195));
    layer0_outputs(3111) <= (inputs(148)) xor (inputs(5));
    layer0_outputs(3112) <= not((inputs(16)) xor (inputs(131)));
    layer0_outputs(3113) <= not(inputs(36));
    layer0_outputs(3114) <= not(inputs(200)) or (inputs(130));
    layer0_outputs(3115) <= (inputs(27)) xor (inputs(126));
    layer0_outputs(3116) <= not(inputs(115)) or (inputs(2));
    layer0_outputs(3117) <= not((inputs(211)) xor (inputs(50)));
    layer0_outputs(3118) <= not((inputs(130)) or (inputs(133)));
    layer0_outputs(3119) <= not(inputs(215)) or (inputs(254));
    layer0_outputs(3120) <= not(inputs(133));
    layer0_outputs(3121) <= (inputs(223)) or (inputs(47));
    layer0_outputs(3122) <= not(inputs(190)) or (inputs(252));
    layer0_outputs(3123) <= not(inputs(12));
    layer0_outputs(3124) <= (inputs(77)) and not (inputs(244));
    layer0_outputs(3125) <= not(inputs(183));
    layer0_outputs(3126) <= not((inputs(200)) xor (inputs(34)));
    layer0_outputs(3127) <= not((inputs(106)) or (inputs(147)));
    layer0_outputs(3128) <= not((inputs(236)) xor (inputs(232)));
    layer0_outputs(3129) <= (inputs(197)) xor (inputs(34));
    layer0_outputs(3130) <= not((inputs(178)) or (inputs(36)));
    layer0_outputs(3131) <= (inputs(109)) xor (inputs(116));
    layer0_outputs(3132) <= not((inputs(86)) xor (inputs(212)));
    layer0_outputs(3133) <= (inputs(33)) and not (inputs(126));
    layer0_outputs(3134) <= (inputs(204)) or (inputs(149));
    layer0_outputs(3135) <= not(inputs(138)) or (inputs(3));
    layer0_outputs(3136) <= not((inputs(146)) xor (inputs(74)));
    layer0_outputs(3137) <= not(inputs(121));
    layer0_outputs(3138) <= not(inputs(103));
    layer0_outputs(3139) <= not(inputs(148)) or (inputs(6));
    layer0_outputs(3140) <= not(inputs(214));
    layer0_outputs(3141) <= not((inputs(198)) and (inputs(91)));
    layer0_outputs(3142) <= (inputs(111)) or (inputs(110));
    layer0_outputs(3143) <= not(inputs(210)) or (inputs(189));
    layer0_outputs(3144) <= not(inputs(150));
    layer0_outputs(3145) <= inputs(133);
    layer0_outputs(3146) <= (inputs(38)) xor (inputs(26));
    layer0_outputs(3147) <= not((inputs(211)) or (inputs(68)));
    layer0_outputs(3148) <= not(inputs(87)) or (inputs(42));
    layer0_outputs(3149) <= not((inputs(83)) or (inputs(95)));
    layer0_outputs(3150) <= not(inputs(0));
    layer0_outputs(3151) <= not(inputs(232));
    layer0_outputs(3152) <= not(inputs(224));
    layer0_outputs(3153) <= (inputs(157)) and not (inputs(2));
    layer0_outputs(3154) <= not(inputs(14)) or (inputs(254));
    layer0_outputs(3155) <= not((inputs(42)) xor (inputs(127)));
    layer0_outputs(3156) <= (inputs(46)) and (inputs(64));
    layer0_outputs(3157) <= not((inputs(175)) or (inputs(91)));
    layer0_outputs(3158) <= not((inputs(147)) xor (inputs(50)));
    layer0_outputs(3159) <= (inputs(65)) and not (inputs(44));
    layer0_outputs(3160) <= not((inputs(52)) or (inputs(128)));
    layer0_outputs(3161) <= not(inputs(224));
    layer0_outputs(3162) <= inputs(137);
    layer0_outputs(3163) <= not(inputs(166));
    layer0_outputs(3164) <= (inputs(203)) and not (inputs(141));
    layer0_outputs(3165) <= not((inputs(59)) xor (inputs(16)));
    layer0_outputs(3166) <= not(inputs(11));
    layer0_outputs(3167) <= (inputs(242)) or (inputs(200));
    layer0_outputs(3168) <= (inputs(43)) and not (inputs(76));
    layer0_outputs(3169) <= not((inputs(34)) and (inputs(222)));
    layer0_outputs(3170) <= not((inputs(119)) or (inputs(44)));
    layer0_outputs(3171) <= not(inputs(86)) or (inputs(207));
    layer0_outputs(3172) <= (inputs(233)) and not (inputs(66));
    layer0_outputs(3173) <= not(inputs(192)) or (inputs(65));
    layer0_outputs(3174) <= not(inputs(118)) or (inputs(81));
    layer0_outputs(3175) <= (inputs(222)) and not (inputs(14));
    layer0_outputs(3176) <= not((inputs(57)) xor (inputs(66)));
    layer0_outputs(3177) <= not((inputs(104)) xor (inputs(144)));
    layer0_outputs(3178) <= (inputs(171)) and not (inputs(128));
    layer0_outputs(3179) <= (inputs(113)) xor (inputs(103));
    layer0_outputs(3180) <= not(inputs(31));
    layer0_outputs(3181) <= not(inputs(243));
    layer0_outputs(3182) <= not((inputs(51)) xor (inputs(234)));
    layer0_outputs(3183) <= not(inputs(242)) or (inputs(250));
    layer0_outputs(3184) <= not((inputs(228)) xor (inputs(143)));
    layer0_outputs(3185) <= not(inputs(13));
    layer0_outputs(3186) <= (inputs(77)) or (inputs(87));
    layer0_outputs(3187) <= (inputs(44)) or (inputs(140));
    layer0_outputs(3188) <= not(inputs(109)) or (inputs(13));
    layer0_outputs(3189) <= (inputs(63)) xor (inputs(250));
    layer0_outputs(3190) <= not(inputs(215));
    layer0_outputs(3191) <= not(inputs(121));
    layer0_outputs(3192) <= not((inputs(42)) or (inputs(22)));
    layer0_outputs(3193) <= (inputs(26)) xor (inputs(131));
    layer0_outputs(3194) <= inputs(31);
    layer0_outputs(3195) <= not((inputs(219)) or (inputs(109)));
    layer0_outputs(3196) <= not((inputs(91)) xor (inputs(53)));
    layer0_outputs(3197) <= not(inputs(232));
    layer0_outputs(3198) <= not(inputs(178)) or (inputs(121));
    layer0_outputs(3199) <= inputs(58);
    layer0_outputs(3200) <= '0';
    layer0_outputs(3201) <= not((inputs(48)) xor (inputs(230)));
    layer0_outputs(3202) <= inputs(8);
    layer0_outputs(3203) <= (inputs(187)) and not (inputs(6));
    layer0_outputs(3204) <= not(inputs(205));
    layer0_outputs(3205) <= inputs(13);
    layer0_outputs(3206) <= (inputs(43)) or (inputs(131));
    layer0_outputs(3207) <= not((inputs(65)) or (inputs(21)));
    layer0_outputs(3208) <= (inputs(138)) and not (inputs(194));
    layer0_outputs(3209) <= not((inputs(65)) and (inputs(35)));
    layer0_outputs(3210) <= not((inputs(152)) xor (inputs(235)));
    layer0_outputs(3211) <= (inputs(141)) and not (inputs(143));
    layer0_outputs(3212) <= not(inputs(137));
    layer0_outputs(3213) <= not(inputs(56));
    layer0_outputs(3214) <= not((inputs(57)) or (inputs(197)));
    layer0_outputs(3215) <= not(inputs(131)) or (inputs(208));
    layer0_outputs(3216) <= not(inputs(82));
    layer0_outputs(3217) <= (inputs(66)) xor (inputs(215));
    layer0_outputs(3218) <= not((inputs(154)) and (inputs(70)));
    layer0_outputs(3219) <= (inputs(43)) and not (inputs(145));
    layer0_outputs(3220) <= (inputs(198)) xor (inputs(197));
    layer0_outputs(3221) <= not(inputs(225));
    layer0_outputs(3222) <= (inputs(83)) or (inputs(105));
    layer0_outputs(3223) <= not((inputs(132)) or (inputs(38)));
    layer0_outputs(3224) <= (inputs(221)) or (inputs(39));
    layer0_outputs(3225) <= (inputs(130)) and not (inputs(237));
    layer0_outputs(3226) <= not(inputs(132)) or (inputs(37));
    layer0_outputs(3227) <= (inputs(186)) and not (inputs(241));
    layer0_outputs(3228) <= not(inputs(72)) or (inputs(225));
    layer0_outputs(3229) <= inputs(31);
    layer0_outputs(3230) <= inputs(132);
    layer0_outputs(3231) <= '1';
    layer0_outputs(3232) <= (inputs(91)) and not (inputs(151));
    layer0_outputs(3233) <= not(inputs(139));
    layer0_outputs(3234) <= (inputs(102)) or (inputs(158));
    layer0_outputs(3235) <= (inputs(174)) xor (inputs(145));
    layer0_outputs(3236) <= (inputs(141)) or (inputs(171));
    layer0_outputs(3237) <= inputs(196);
    layer0_outputs(3238) <= (inputs(174)) and not (inputs(220));
    layer0_outputs(3239) <= (inputs(162)) or (inputs(99));
    layer0_outputs(3240) <= inputs(20);
    layer0_outputs(3241) <= not((inputs(123)) xor (inputs(114)));
    layer0_outputs(3242) <= not(inputs(136));
    layer0_outputs(3243) <= not((inputs(221)) or (inputs(50)));
    layer0_outputs(3244) <= (inputs(252)) xor (inputs(166));
    layer0_outputs(3245) <= not(inputs(224)) or (inputs(7));
    layer0_outputs(3246) <= inputs(224);
    layer0_outputs(3247) <= (inputs(165)) or (inputs(100));
    layer0_outputs(3248) <= not((inputs(198)) or (inputs(157)));
    layer0_outputs(3249) <= not((inputs(169)) or (inputs(219)));
    layer0_outputs(3250) <= not(inputs(24));
    layer0_outputs(3251) <= (inputs(255)) and not (inputs(80));
    layer0_outputs(3252) <= inputs(39);
    layer0_outputs(3253) <= (inputs(183)) or (inputs(182));
    layer0_outputs(3254) <= (inputs(240)) xor (inputs(158));
    layer0_outputs(3255) <= not(inputs(142)) or (inputs(192));
    layer0_outputs(3256) <= inputs(40);
    layer0_outputs(3257) <= not(inputs(198));
    layer0_outputs(3258) <= (inputs(204)) and not (inputs(146));
    layer0_outputs(3259) <= (inputs(94)) or (inputs(154));
    layer0_outputs(3260) <= not((inputs(1)) xor (inputs(163)));
    layer0_outputs(3261) <= not(inputs(255)) or (inputs(9));
    layer0_outputs(3262) <= not((inputs(216)) or (inputs(217)));
    layer0_outputs(3263) <= not((inputs(123)) xor (inputs(168)));
    layer0_outputs(3264) <= not((inputs(138)) xor (inputs(122)));
    layer0_outputs(3265) <= not(inputs(118));
    layer0_outputs(3266) <= not(inputs(104)) or (inputs(84));
    layer0_outputs(3267) <= (inputs(3)) xor (inputs(125));
    layer0_outputs(3268) <= not((inputs(125)) xor (inputs(29)));
    layer0_outputs(3269) <= (inputs(12)) or (inputs(79));
    layer0_outputs(3270) <= (inputs(23)) or (inputs(141));
    layer0_outputs(3271) <= inputs(136);
    layer0_outputs(3272) <= '0';
    layer0_outputs(3273) <= not(inputs(174));
    layer0_outputs(3274) <= inputs(118);
    layer0_outputs(3275) <= (inputs(48)) or (inputs(48));
    layer0_outputs(3276) <= not(inputs(179));
    layer0_outputs(3277) <= not(inputs(45));
    layer0_outputs(3278) <= inputs(118);
    layer0_outputs(3279) <= (inputs(224)) or (inputs(0));
    layer0_outputs(3280) <= inputs(200);
    layer0_outputs(3281) <= not((inputs(249)) or (inputs(234)));
    layer0_outputs(3282) <= not((inputs(109)) or (inputs(52)));
    layer0_outputs(3283) <= not((inputs(91)) or (inputs(19)));
    layer0_outputs(3284) <= '1';
    layer0_outputs(3285) <= (inputs(245)) or (inputs(170));
    layer0_outputs(3286) <= '0';
    layer0_outputs(3287) <= not((inputs(195)) or (inputs(36)));
    layer0_outputs(3288) <= (inputs(232)) xor (inputs(17));
    layer0_outputs(3289) <= not((inputs(153)) xor (inputs(171)));
    layer0_outputs(3290) <= not(inputs(116)) or (inputs(192));
    layer0_outputs(3291) <= (inputs(83)) or (inputs(126));
    layer0_outputs(3292) <= not(inputs(84)) or (inputs(193));
    layer0_outputs(3293) <= '0';
    layer0_outputs(3294) <= not((inputs(152)) xor (inputs(65)));
    layer0_outputs(3295) <= not((inputs(27)) xor (inputs(241)));
    layer0_outputs(3296) <= inputs(148);
    layer0_outputs(3297) <= not((inputs(103)) or (inputs(113)));
    layer0_outputs(3298) <= not((inputs(145)) xor (inputs(35)));
    layer0_outputs(3299) <= (inputs(16)) or (inputs(25));
    layer0_outputs(3300) <= not(inputs(165));
    layer0_outputs(3301) <= (inputs(102)) and not (inputs(49));
    layer0_outputs(3302) <= not(inputs(154)) or (inputs(245));
    layer0_outputs(3303) <= not((inputs(182)) or (inputs(188)));
    layer0_outputs(3304) <= (inputs(96)) and not (inputs(208));
    layer0_outputs(3305) <= not(inputs(127));
    layer0_outputs(3306) <= (inputs(79)) and (inputs(201));
    layer0_outputs(3307) <= (inputs(56)) or (inputs(111));
    layer0_outputs(3308) <= (inputs(225)) and not (inputs(249));
    layer0_outputs(3309) <= (inputs(93)) or (inputs(159));
    layer0_outputs(3310) <= (inputs(30)) and not (inputs(29));
    layer0_outputs(3311) <= (inputs(92)) and (inputs(11));
    layer0_outputs(3312) <= not((inputs(158)) or (inputs(162)));
    layer0_outputs(3313) <= (inputs(104)) and not (inputs(223));
    layer0_outputs(3314) <= '0';
    layer0_outputs(3315) <= (inputs(226)) xor (inputs(110));
    layer0_outputs(3316) <= (inputs(84)) and not (inputs(136));
    layer0_outputs(3317) <= (inputs(171)) or (inputs(193));
    layer0_outputs(3318) <= (inputs(28)) or (inputs(250));
    layer0_outputs(3319) <= not((inputs(178)) xor (inputs(97)));
    layer0_outputs(3320) <= (inputs(201)) or (inputs(6));
    layer0_outputs(3321) <= (inputs(27)) xor (inputs(209));
    layer0_outputs(3322) <= not(inputs(40)) or (inputs(34));
    layer0_outputs(3323) <= not((inputs(119)) xor (inputs(44)));
    layer0_outputs(3324) <= not(inputs(107)) or (inputs(17));
    layer0_outputs(3325) <= not((inputs(138)) xor (inputs(32)));
    layer0_outputs(3326) <= not(inputs(187)) or (inputs(174));
    layer0_outputs(3327) <= (inputs(197)) and not (inputs(103));
    layer0_outputs(3328) <= not(inputs(146));
    layer0_outputs(3329) <= not(inputs(111)) or (inputs(29));
    layer0_outputs(3330) <= '1';
    layer0_outputs(3331) <= not((inputs(14)) xor (inputs(9)));
    layer0_outputs(3332) <= (inputs(124)) and (inputs(150));
    layer0_outputs(3333) <= not((inputs(23)) or (inputs(68)));
    layer0_outputs(3334) <= not(inputs(25)) or (inputs(97));
    layer0_outputs(3335) <= (inputs(126)) or (inputs(102));
    layer0_outputs(3336) <= not((inputs(177)) or (inputs(167)));
    layer0_outputs(3337) <= not(inputs(224)) or (inputs(68));
    layer0_outputs(3338) <= not((inputs(55)) and (inputs(56)));
    layer0_outputs(3339) <= (inputs(137)) xor (inputs(225));
    layer0_outputs(3340) <= inputs(117);
    layer0_outputs(3341) <= not(inputs(183));
    layer0_outputs(3342) <= not((inputs(145)) xor (inputs(142)));
    layer0_outputs(3343) <= (inputs(155)) xor (inputs(191));
    layer0_outputs(3344) <= not(inputs(153));
    layer0_outputs(3345) <= not((inputs(88)) xor (inputs(24)));
    layer0_outputs(3346) <= inputs(31);
    layer0_outputs(3347) <= (inputs(7)) or (inputs(107));
    layer0_outputs(3348) <= not((inputs(17)) or (inputs(72)));
    layer0_outputs(3349) <= inputs(229);
    layer0_outputs(3350) <= (inputs(187)) or (inputs(77));
    layer0_outputs(3351) <= '1';
    layer0_outputs(3352) <= not(inputs(149)) or (inputs(222));
    layer0_outputs(3353) <= not(inputs(84));
    layer0_outputs(3354) <= not((inputs(41)) or (inputs(110)));
    layer0_outputs(3355) <= (inputs(128)) or (inputs(242));
    layer0_outputs(3356) <= (inputs(217)) or (inputs(220));
    layer0_outputs(3357) <= not((inputs(223)) xor (inputs(119)));
    layer0_outputs(3358) <= not((inputs(26)) xor (inputs(162)));
    layer0_outputs(3359) <= (inputs(167)) xor (inputs(177));
    layer0_outputs(3360) <= not((inputs(22)) or (inputs(52)));
    layer0_outputs(3361) <= not((inputs(241)) or (inputs(106)));
    layer0_outputs(3362) <= (inputs(169)) xor (inputs(19));
    layer0_outputs(3363) <= inputs(52);
    layer0_outputs(3364) <= (inputs(198)) and not (inputs(129));
    layer0_outputs(3365) <= (inputs(213)) or (inputs(250));
    layer0_outputs(3366) <= (inputs(134)) or (inputs(221));
    layer0_outputs(3367) <= (inputs(205)) or (inputs(181));
    layer0_outputs(3368) <= not(inputs(212));
    layer0_outputs(3369) <= (inputs(73)) xor (inputs(180));
    layer0_outputs(3370) <= not((inputs(174)) or (inputs(133)));
    layer0_outputs(3371) <= (inputs(45)) or (inputs(234));
    layer0_outputs(3372) <= not((inputs(216)) xor (inputs(35)));
    layer0_outputs(3373) <= (inputs(28)) and not (inputs(178));
    layer0_outputs(3374) <= (inputs(215)) or (inputs(126));
    layer0_outputs(3375) <= not(inputs(215)) or (inputs(221));
    layer0_outputs(3376) <= not((inputs(151)) xor (inputs(31)));
    layer0_outputs(3377) <= inputs(114);
    layer0_outputs(3378) <= not(inputs(49)) or (inputs(51));
    layer0_outputs(3379) <= (inputs(206)) xor (inputs(101));
    layer0_outputs(3380) <= not(inputs(118)) or (inputs(209));
    layer0_outputs(3381) <= (inputs(229)) or (inputs(116));
    layer0_outputs(3382) <= (inputs(162)) or (inputs(94));
    layer0_outputs(3383) <= inputs(102);
    layer0_outputs(3384) <= (inputs(196)) xor (inputs(39));
    layer0_outputs(3385) <= not((inputs(65)) or (inputs(114)));
    layer0_outputs(3386) <= (inputs(177)) or (inputs(99));
    layer0_outputs(3387) <= not((inputs(213)) or (inputs(55)));
    layer0_outputs(3388) <= (inputs(249)) and not (inputs(128));
    layer0_outputs(3389) <= not((inputs(224)) or (inputs(243)));
    layer0_outputs(3390) <= '0';
    layer0_outputs(3391) <= (inputs(55)) and not (inputs(160));
    layer0_outputs(3392) <= not((inputs(33)) xor (inputs(212)));
    layer0_outputs(3393) <= (inputs(232)) xor (inputs(74));
    layer0_outputs(3394) <= not(inputs(120)) or (inputs(61));
    layer0_outputs(3395) <= not((inputs(135)) xor (inputs(9)));
    layer0_outputs(3396) <= not((inputs(46)) xor (inputs(112)));
    layer0_outputs(3397) <= inputs(180);
    layer0_outputs(3398) <= inputs(240);
    layer0_outputs(3399) <= not((inputs(51)) or (inputs(182)));
    layer0_outputs(3400) <= not(inputs(182)) or (inputs(155));
    layer0_outputs(3401) <= inputs(221);
    layer0_outputs(3402) <= (inputs(56)) xor (inputs(245));
    layer0_outputs(3403) <= not(inputs(230)) or (inputs(249));
    layer0_outputs(3404) <= inputs(40);
    layer0_outputs(3405) <= not((inputs(91)) and (inputs(26)));
    layer0_outputs(3406) <= not(inputs(180));
    layer0_outputs(3407) <= (inputs(73)) and (inputs(122));
    layer0_outputs(3408) <= not(inputs(47)) or (inputs(71));
    layer0_outputs(3409) <= not(inputs(129)) or (inputs(81));
    layer0_outputs(3410) <= (inputs(154)) or (inputs(14));
    layer0_outputs(3411) <= not((inputs(4)) xor (inputs(118)));
    layer0_outputs(3412) <= (inputs(89)) and not (inputs(148));
    layer0_outputs(3413) <= (inputs(111)) and not (inputs(174));
    layer0_outputs(3414) <= inputs(22);
    layer0_outputs(3415) <= not(inputs(68));
    layer0_outputs(3416) <= (inputs(23)) or (inputs(74));
    layer0_outputs(3417) <= (inputs(162)) and not (inputs(98));
    layer0_outputs(3418) <= '0';
    layer0_outputs(3419) <= (inputs(44)) and not (inputs(255));
    layer0_outputs(3420) <= (inputs(236)) xor (inputs(214));
    layer0_outputs(3421) <= not(inputs(134));
    layer0_outputs(3422) <= not((inputs(103)) or (inputs(143)));
    layer0_outputs(3423) <= (inputs(106)) xor (inputs(124));
    layer0_outputs(3424) <= inputs(255);
    layer0_outputs(3425) <= '1';
    layer0_outputs(3426) <= '1';
    layer0_outputs(3427) <= not((inputs(24)) or (inputs(53)));
    layer0_outputs(3428) <= not((inputs(39)) or (inputs(16)));
    layer0_outputs(3429) <= not(inputs(253)) or (inputs(145));
    layer0_outputs(3430) <= (inputs(254)) and not (inputs(4));
    layer0_outputs(3431) <= (inputs(123)) and (inputs(14));
    layer0_outputs(3432) <= (inputs(157)) and not (inputs(59));
    layer0_outputs(3433) <= inputs(102);
    layer0_outputs(3434) <= (inputs(60)) xor (inputs(85));
    layer0_outputs(3435) <= '1';
    layer0_outputs(3436) <= not((inputs(204)) xor (inputs(144)));
    layer0_outputs(3437) <= not((inputs(198)) or (inputs(179)));
    layer0_outputs(3438) <= inputs(189);
    layer0_outputs(3439) <= not(inputs(36)) or (inputs(159));
    layer0_outputs(3440) <= (inputs(101)) and not (inputs(173));
    layer0_outputs(3441) <= not((inputs(227)) xor (inputs(236)));
    layer0_outputs(3442) <= not((inputs(6)) xor (inputs(109)));
    layer0_outputs(3443) <= inputs(1);
    layer0_outputs(3444) <= not(inputs(78));
    layer0_outputs(3445) <= (inputs(224)) or (inputs(58));
    layer0_outputs(3446) <= (inputs(88)) or (inputs(108));
    layer0_outputs(3447) <= (inputs(150)) and not (inputs(78));
    layer0_outputs(3448) <= (inputs(138)) or (inputs(200));
    layer0_outputs(3449) <= (inputs(182)) or (inputs(92));
    layer0_outputs(3450) <= (inputs(17)) xor (inputs(230));
    layer0_outputs(3451) <= not((inputs(1)) or (inputs(41)));
    layer0_outputs(3452) <= not((inputs(8)) or (inputs(211)));
    layer0_outputs(3453) <= (inputs(227)) xor (inputs(201));
    layer0_outputs(3454) <= not(inputs(108));
    layer0_outputs(3455) <= (inputs(91)) or (inputs(25));
    layer0_outputs(3456) <= inputs(68);
    layer0_outputs(3457) <= (inputs(105)) or (inputs(211));
    layer0_outputs(3458) <= (inputs(161)) or (inputs(47));
    layer0_outputs(3459) <= not((inputs(198)) xor (inputs(126)));
    layer0_outputs(3460) <= not(inputs(174)) or (inputs(21));
    layer0_outputs(3461) <= inputs(148);
    layer0_outputs(3462) <= (inputs(90)) and not (inputs(164));
    layer0_outputs(3463) <= (inputs(75)) or (inputs(140));
    layer0_outputs(3464) <= not((inputs(104)) or (inputs(125)));
    layer0_outputs(3465) <= (inputs(217)) or (inputs(73));
    layer0_outputs(3466) <= not((inputs(122)) or (inputs(174)));
    layer0_outputs(3467) <= not((inputs(91)) or (inputs(82)));
    layer0_outputs(3468) <= not((inputs(18)) xor (inputs(124)));
    layer0_outputs(3469) <= not(inputs(170));
    layer0_outputs(3470) <= not((inputs(166)) or (inputs(210)));
    layer0_outputs(3471) <= not((inputs(120)) and (inputs(115)));
    layer0_outputs(3472) <= not(inputs(104)) or (inputs(176));
    layer0_outputs(3473) <= not(inputs(148));
    layer0_outputs(3474) <= not((inputs(245)) and (inputs(82)));
    layer0_outputs(3475) <= (inputs(242)) and not (inputs(186));
    layer0_outputs(3476) <= inputs(102);
    layer0_outputs(3477) <= (inputs(40)) or (inputs(20));
    layer0_outputs(3478) <= not((inputs(137)) or (inputs(119)));
    layer0_outputs(3479) <= not(inputs(70));
    layer0_outputs(3480) <= not(inputs(150)) or (inputs(163));
    layer0_outputs(3481) <= '0';
    layer0_outputs(3482) <= (inputs(120)) and not (inputs(19));
    layer0_outputs(3483) <= not(inputs(141));
    layer0_outputs(3484) <= inputs(121);
    layer0_outputs(3485) <= (inputs(95)) and not (inputs(241));
    layer0_outputs(3486) <= not(inputs(254));
    layer0_outputs(3487) <= '1';
    layer0_outputs(3488) <= not((inputs(143)) or (inputs(24)));
    layer0_outputs(3489) <= not(inputs(141));
    layer0_outputs(3490) <= not((inputs(136)) and (inputs(215)));
    layer0_outputs(3491) <= not(inputs(73)) or (inputs(174));
    layer0_outputs(3492) <= not((inputs(47)) or (inputs(181)));
    layer0_outputs(3493) <= (inputs(110)) xor (inputs(213));
    layer0_outputs(3494) <= (inputs(66)) and not (inputs(26));
    layer0_outputs(3495) <= inputs(236);
    layer0_outputs(3496) <= (inputs(74)) xor (inputs(220));
    layer0_outputs(3497) <= (inputs(240)) xor (inputs(20));
    layer0_outputs(3498) <= not((inputs(164)) or (inputs(230)));
    layer0_outputs(3499) <= not(inputs(159));
    layer0_outputs(3500) <= (inputs(196)) xor (inputs(6));
    layer0_outputs(3501) <= not((inputs(213)) or (inputs(37)));
    layer0_outputs(3502) <= (inputs(226)) xor (inputs(200));
    layer0_outputs(3503) <= not(inputs(253));
    layer0_outputs(3504) <= (inputs(50)) or (inputs(147));
    layer0_outputs(3505) <= not(inputs(225)) or (inputs(38));
    layer0_outputs(3506) <= not(inputs(25)) or (inputs(82));
    layer0_outputs(3507) <= not((inputs(67)) or (inputs(106)));
    layer0_outputs(3508) <= (inputs(15)) and not (inputs(209));
    layer0_outputs(3509) <= not((inputs(234)) or (inputs(234)));
    layer0_outputs(3510) <= (inputs(70)) and not (inputs(77));
    layer0_outputs(3511) <= (inputs(50)) xor (inputs(231));
    layer0_outputs(3512) <= '0';
    layer0_outputs(3513) <= not((inputs(152)) xor (inputs(208)));
    layer0_outputs(3514) <= not((inputs(158)) or (inputs(67)));
    layer0_outputs(3515) <= not((inputs(80)) xor (inputs(107)));
    layer0_outputs(3516) <= (inputs(0)) and not (inputs(143));
    layer0_outputs(3517) <= not((inputs(154)) or (inputs(75)));
    layer0_outputs(3518) <= (inputs(73)) and not (inputs(143));
    layer0_outputs(3519) <= '0';
    layer0_outputs(3520) <= not(inputs(86)) or (inputs(65));
    layer0_outputs(3521) <= not((inputs(9)) or (inputs(125)));
    layer0_outputs(3522) <= not((inputs(84)) or (inputs(63)));
    layer0_outputs(3523) <= not((inputs(176)) or (inputs(95)));
    layer0_outputs(3524) <= (inputs(133)) or (inputs(125));
    layer0_outputs(3525) <= (inputs(28)) or (inputs(123));
    layer0_outputs(3526) <= (inputs(121)) or (inputs(240));
    layer0_outputs(3527) <= not(inputs(218)) or (inputs(13));
    layer0_outputs(3528) <= not(inputs(52)) or (inputs(172));
    layer0_outputs(3529) <= not(inputs(156));
    layer0_outputs(3530) <= inputs(210);
    layer0_outputs(3531) <= not(inputs(216));
    layer0_outputs(3532) <= inputs(17);
    layer0_outputs(3533) <= not((inputs(139)) or (inputs(153)));
    layer0_outputs(3534) <= inputs(121);
    layer0_outputs(3535) <= not(inputs(116)) or (inputs(98));
    layer0_outputs(3536) <= not((inputs(198)) xor (inputs(50)));
    layer0_outputs(3537) <= inputs(42);
    layer0_outputs(3538) <= (inputs(129)) and not (inputs(176));
    layer0_outputs(3539) <= inputs(92);
    layer0_outputs(3540) <= (inputs(120)) xor (inputs(245));
    layer0_outputs(3541) <= not(inputs(247));
    layer0_outputs(3542) <= (inputs(86)) or (inputs(68));
    layer0_outputs(3543) <= '1';
    layer0_outputs(3544) <= inputs(176);
    layer0_outputs(3545) <= not((inputs(233)) or (inputs(184)));
    layer0_outputs(3546) <= not(inputs(205)) or (inputs(54));
    layer0_outputs(3547) <= not((inputs(40)) xor (inputs(143)));
    layer0_outputs(3548) <= (inputs(67)) and not (inputs(29));
    layer0_outputs(3549) <= (inputs(184)) xor (inputs(112));
    layer0_outputs(3550) <= inputs(62);
    layer0_outputs(3551) <= not((inputs(90)) and (inputs(74)));
    layer0_outputs(3552) <= (inputs(85)) xor (inputs(102));
    layer0_outputs(3553) <= not(inputs(148));
    layer0_outputs(3554) <= not((inputs(177)) and (inputs(24)));
    layer0_outputs(3555) <= inputs(136);
    layer0_outputs(3556) <= inputs(138);
    layer0_outputs(3557) <= not(inputs(204));
    layer0_outputs(3558) <= not(inputs(214));
    layer0_outputs(3559) <= (inputs(126)) or (inputs(78));
    layer0_outputs(3560) <= (inputs(230)) and not (inputs(20));
    layer0_outputs(3561) <= not((inputs(102)) xor (inputs(115)));
    layer0_outputs(3562) <= '0';
    layer0_outputs(3563) <= inputs(165);
    layer0_outputs(3564) <= not((inputs(221)) and (inputs(9)));
    layer0_outputs(3565) <= '0';
    layer0_outputs(3566) <= not(inputs(80));
    layer0_outputs(3567) <= (inputs(166)) or (inputs(98));
    layer0_outputs(3568) <= not(inputs(255)) or (inputs(64));
    layer0_outputs(3569) <= not(inputs(45));
    layer0_outputs(3570) <= not((inputs(85)) xor (inputs(98)));
    layer0_outputs(3571) <= (inputs(238)) and not (inputs(161));
    layer0_outputs(3572) <= not((inputs(208)) or (inputs(68)));
    layer0_outputs(3573) <= (inputs(39)) xor (inputs(86));
    layer0_outputs(3574) <= not(inputs(74));
    layer0_outputs(3575) <= (inputs(44)) and not (inputs(205));
    layer0_outputs(3576) <= not(inputs(53));
    layer0_outputs(3577) <= (inputs(193)) or (inputs(135));
    layer0_outputs(3578) <= not(inputs(186));
    layer0_outputs(3579) <= not(inputs(3)) or (inputs(255));
    layer0_outputs(3580) <= (inputs(101)) or (inputs(147));
    layer0_outputs(3581) <= inputs(107);
    layer0_outputs(3582) <= not((inputs(149)) or (inputs(82)));
    layer0_outputs(3583) <= not(inputs(106));
    layer0_outputs(3584) <= not((inputs(214)) xor (inputs(110)));
    layer0_outputs(3585) <= not(inputs(76));
    layer0_outputs(3586) <= not((inputs(161)) xor (inputs(86)));
    layer0_outputs(3587) <= not((inputs(91)) xor (inputs(50)));
    layer0_outputs(3588) <= not((inputs(74)) or (inputs(240)));
    layer0_outputs(3589) <= (inputs(41)) and not (inputs(163));
    layer0_outputs(3590) <= not((inputs(32)) or (inputs(226)));
    layer0_outputs(3591) <= inputs(136);
    layer0_outputs(3592) <= not((inputs(50)) xor (inputs(193)));
    layer0_outputs(3593) <= not((inputs(144)) or (inputs(138)));
    layer0_outputs(3594) <= inputs(249);
    layer0_outputs(3595) <= not(inputs(98));
    layer0_outputs(3596) <= not(inputs(149)) or (inputs(199));
    layer0_outputs(3597) <= (inputs(172)) and not (inputs(34));
    layer0_outputs(3598) <= not(inputs(41)) or (inputs(18));
    layer0_outputs(3599) <= (inputs(150)) or (inputs(97));
    layer0_outputs(3600) <= not((inputs(88)) or (inputs(231)));
    layer0_outputs(3601) <= not((inputs(102)) xor (inputs(53)));
    layer0_outputs(3602) <= not(inputs(105));
    layer0_outputs(3603) <= '0';
    layer0_outputs(3604) <= inputs(169);
    layer0_outputs(3605) <= (inputs(236)) or (inputs(134));
    layer0_outputs(3606) <= not(inputs(255));
    layer0_outputs(3607) <= not((inputs(7)) xor (inputs(219)));
    layer0_outputs(3608) <= not((inputs(87)) or (inputs(1)));
    layer0_outputs(3609) <= inputs(134);
    layer0_outputs(3610) <= inputs(104);
    layer0_outputs(3611) <= not(inputs(3)) or (inputs(250));
    layer0_outputs(3612) <= not(inputs(49)) or (inputs(29));
    layer0_outputs(3613) <= (inputs(236)) or (inputs(139));
    layer0_outputs(3614) <= inputs(191);
    layer0_outputs(3615) <= not((inputs(116)) or (inputs(47)));
    layer0_outputs(3616) <= (inputs(44)) and not (inputs(248));
    layer0_outputs(3617) <= not(inputs(48));
    layer0_outputs(3618) <= not((inputs(180)) or (inputs(53)));
    layer0_outputs(3619) <= not((inputs(48)) xor (inputs(184)));
    layer0_outputs(3620) <= not((inputs(21)) or (inputs(239)));
    layer0_outputs(3621) <= (inputs(107)) xor (inputs(112));
    layer0_outputs(3622) <= (inputs(169)) or (inputs(80));
    layer0_outputs(3623) <= not(inputs(160)) or (inputs(79));
    layer0_outputs(3624) <= (inputs(32)) xor (inputs(184));
    layer0_outputs(3625) <= not(inputs(97));
    layer0_outputs(3626) <= not(inputs(67));
    layer0_outputs(3627) <= (inputs(29)) or (inputs(138));
    layer0_outputs(3628) <= not((inputs(50)) or (inputs(210)));
    layer0_outputs(3629) <= (inputs(245)) and not (inputs(195));
    layer0_outputs(3630) <= inputs(166);
    layer0_outputs(3631) <= not((inputs(144)) xor (inputs(96)));
    layer0_outputs(3632) <= not(inputs(84));
    layer0_outputs(3633) <= not(inputs(91)) or (inputs(194));
    layer0_outputs(3634) <= not((inputs(216)) or (inputs(34)));
    layer0_outputs(3635) <= inputs(56);
    layer0_outputs(3636) <= not(inputs(87)) or (inputs(223));
    layer0_outputs(3637) <= not(inputs(111)) or (inputs(112));
    layer0_outputs(3638) <= not(inputs(69));
    layer0_outputs(3639) <= (inputs(166)) or (inputs(189));
    layer0_outputs(3640) <= not((inputs(164)) or (inputs(92)));
    layer0_outputs(3641) <= (inputs(105)) and not (inputs(21));
    layer0_outputs(3642) <= inputs(120);
    layer0_outputs(3643) <= not(inputs(131)) or (inputs(188));
    layer0_outputs(3644) <= not(inputs(166)) or (inputs(21));
    layer0_outputs(3645) <= (inputs(221)) and (inputs(9));
    layer0_outputs(3646) <= (inputs(85)) and (inputs(119));
    layer0_outputs(3647) <= inputs(231);
    layer0_outputs(3648) <= (inputs(104)) or (inputs(194));
    layer0_outputs(3649) <= not(inputs(116)) or (inputs(6));
    layer0_outputs(3650) <= not(inputs(64));
    layer0_outputs(3651) <= (inputs(110)) and not (inputs(34));
    layer0_outputs(3652) <= inputs(60);
    layer0_outputs(3653) <= not((inputs(45)) or (inputs(135)));
    layer0_outputs(3654) <= (inputs(216)) and not (inputs(228));
    layer0_outputs(3655) <= inputs(114);
    layer0_outputs(3656) <= not(inputs(132));
    layer0_outputs(3657) <= (inputs(19)) and not (inputs(255));
    layer0_outputs(3658) <= '1';
    layer0_outputs(3659) <= not(inputs(8));
    layer0_outputs(3660) <= '0';
    layer0_outputs(3661) <= (inputs(177)) or (inputs(143));
    layer0_outputs(3662) <= inputs(129);
    layer0_outputs(3663) <= not((inputs(130)) or (inputs(219)));
    layer0_outputs(3664) <= not(inputs(168));
    layer0_outputs(3665) <= not((inputs(192)) xor (inputs(67)));
    layer0_outputs(3666) <= inputs(58);
    layer0_outputs(3667) <= '1';
    layer0_outputs(3668) <= not((inputs(147)) or (inputs(115)));
    layer0_outputs(3669) <= not((inputs(12)) xor (inputs(126)));
    layer0_outputs(3670) <= (inputs(4)) or (inputs(151));
    layer0_outputs(3671) <= not(inputs(166));
    layer0_outputs(3672) <= not(inputs(29)) or (inputs(250));
    layer0_outputs(3673) <= not(inputs(183)) or (inputs(84));
    layer0_outputs(3674) <= (inputs(76)) or (inputs(56));
    layer0_outputs(3675) <= inputs(94);
    layer0_outputs(3676) <= (inputs(252)) xor (inputs(84));
    layer0_outputs(3677) <= not((inputs(114)) or (inputs(160)));
    layer0_outputs(3678) <= (inputs(178)) or (inputs(220));
    layer0_outputs(3679) <= '0';
    layer0_outputs(3680) <= not((inputs(219)) xor (inputs(3)));
    layer0_outputs(3681) <= '0';
    layer0_outputs(3682) <= (inputs(172)) or (inputs(233));
    layer0_outputs(3683) <= '0';
    layer0_outputs(3684) <= inputs(57);
    layer0_outputs(3685) <= not((inputs(140)) xor (inputs(189)));
    layer0_outputs(3686) <= (inputs(203)) or (inputs(167));
    layer0_outputs(3687) <= (inputs(126)) or (inputs(177));
    layer0_outputs(3688) <= not(inputs(123)) or (inputs(109));
    layer0_outputs(3689) <= not((inputs(235)) and (inputs(241)));
    layer0_outputs(3690) <= not(inputs(117));
    layer0_outputs(3691) <= not(inputs(168)) or (inputs(174));
    layer0_outputs(3692) <= not(inputs(142)) or (inputs(26));
    layer0_outputs(3693) <= not(inputs(196)) or (inputs(173));
    layer0_outputs(3694) <= inputs(18);
    layer0_outputs(3695) <= (inputs(72)) xor (inputs(136));
    layer0_outputs(3696) <= not(inputs(146)) or (inputs(211));
    layer0_outputs(3697) <= not(inputs(135)) or (inputs(241));
    layer0_outputs(3698) <= not((inputs(17)) or (inputs(152)));
    layer0_outputs(3699) <= not((inputs(1)) xor (inputs(66)));
    layer0_outputs(3700) <= inputs(134);
    layer0_outputs(3701) <= inputs(194);
    layer0_outputs(3702) <= (inputs(189)) xor (inputs(151));
    layer0_outputs(3703) <= not(inputs(5));
    layer0_outputs(3704) <= (inputs(153)) and not (inputs(187));
    layer0_outputs(3705) <= not((inputs(38)) or (inputs(202)));
    layer0_outputs(3706) <= '0';
    layer0_outputs(3707) <= not(inputs(51));
    layer0_outputs(3708) <= (inputs(223)) and (inputs(239));
    layer0_outputs(3709) <= not((inputs(154)) xor (inputs(227)));
    layer0_outputs(3710) <= not((inputs(9)) xor (inputs(51)));
    layer0_outputs(3711) <= not(inputs(247)) or (inputs(219));
    layer0_outputs(3712) <= not((inputs(72)) or (inputs(155)));
    layer0_outputs(3713) <= (inputs(219)) and not (inputs(239));
    layer0_outputs(3714) <= not((inputs(53)) xor (inputs(16)));
    layer0_outputs(3715) <= (inputs(6)) and not (inputs(96));
    layer0_outputs(3716) <= (inputs(205)) and not (inputs(0));
    layer0_outputs(3717) <= not(inputs(84)) or (inputs(157));
    layer0_outputs(3718) <= inputs(99);
    layer0_outputs(3719) <= not(inputs(121)) or (inputs(145));
    layer0_outputs(3720) <= '0';
    layer0_outputs(3721) <= not((inputs(246)) and (inputs(239)));
    layer0_outputs(3722) <= (inputs(80)) xor (inputs(28));
    layer0_outputs(3723) <= (inputs(45)) or (inputs(105));
    layer0_outputs(3724) <= inputs(26);
    layer0_outputs(3725) <= not(inputs(17));
    layer0_outputs(3726) <= (inputs(139)) and not (inputs(246));
    layer0_outputs(3727) <= inputs(188);
    layer0_outputs(3728) <= '0';
    layer0_outputs(3729) <= not((inputs(117)) xor (inputs(144)));
    layer0_outputs(3730) <= (inputs(27)) or (inputs(241));
    layer0_outputs(3731) <= not((inputs(75)) or (inputs(199)));
    layer0_outputs(3732) <= not((inputs(35)) xor (inputs(68)));
    layer0_outputs(3733) <= not((inputs(247)) or (inputs(252)));
    layer0_outputs(3734) <= (inputs(139)) and not (inputs(224));
    layer0_outputs(3735) <= not(inputs(199)) or (inputs(80));
    layer0_outputs(3736) <= inputs(16);
    layer0_outputs(3737) <= not((inputs(13)) or (inputs(50)));
    layer0_outputs(3738) <= inputs(149);
    layer0_outputs(3739) <= '0';
    layer0_outputs(3740) <= '0';
    layer0_outputs(3741) <= '1';
    layer0_outputs(3742) <= (inputs(174)) and not (inputs(34));
    layer0_outputs(3743) <= not(inputs(184)) or (inputs(29));
    layer0_outputs(3744) <= (inputs(169)) and not (inputs(58));
    layer0_outputs(3745) <= not((inputs(141)) or (inputs(140)));
    layer0_outputs(3746) <= (inputs(85)) and not (inputs(190));
    layer0_outputs(3747) <= inputs(156);
    layer0_outputs(3748) <= not((inputs(158)) or (inputs(40)));
    layer0_outputs(3749) <= not(inputs(217)) or (inputs(43));
    layer0_outputs(3750) <= not((inputs(89)) xor (inputs(131)));
    layer0_outputs(3751) <= not((inputs(119)) or (inputs(204)));
    layer0_outputs(3752) <= not((inputs(212)) or (inputs(176)));
    layer0_outputs(3753) <= (inputs(196)) xor (inputs(28));
    layer0_outputs(3754) <= (inputs(116)) xor (inputs(154));
    layer0_outputs(3755) <= (inputs(117)) and not (inputs(229));
    layer0_outputs(3756) <= not(inputs(130)) or (inputs(19));
    layer0_outputs(3757) <= not((inputs(68)) xor (inputs(18)));
    layer0_outputs(3758) <= inputs(157);
    layer0_outputs(3759) <= not(inputs(40)) or (inputs(44));
    layer0_outputs(3760) <= (inputs(71)) and not (inputs(171));
    layer0_outputs(3761) <= not((inputs(188)) xor (inputs(252)));
    layer0_outputs(3762) <= not((inputs(175)) xor (inputs(115)));
    layer0_outputs(3763) <= not(inputs(60));
    layer0_outputs(3764) <= (inputs(114)) xor (inputs(73));
    layer0_outputs(3765) <= not(inputs(173)) or (inputs(160));
    layer0_outputs(3766) <= not(inputs(23));
    layer0_outputs(3767) <= (inputs(14)) and (inputs(96));
    layer0_outputs(3768) <= (inputs(165)) xor (inputs(62));
    layer0_outputs(3769) <= not(inputs(135));
    layer0_outputs(3770) <= (inputs(96)) xor (inputs(46));
    layer0_outputs(3771) <= not(inputs(89)) or (inputs(151));
    layer0_outputs(3772) <= (inputs(110)) and not (inputs(17));
    layer0_outputs(3773) <= not((inputs(190)) or (inputs(196)));
    layer0_outputs(3774) <= (inputs(37)) or (inputs(13));
    layer0_outputs(3775) <= (inputs(166)) and not (inputs(140));
    layer0_outputs(3776) <= not((inputs(183)) xor (inputs(175)));
    layer0_outputs(3777) <= (inputs(204)) or (inputs(187));
    layer0_outputs(3778) <= (inputs(179)) and not (inputs(44));
    layer0_outputs(3779) <= inputs(1);
    layer0_outputs(3780) <= '0';
    layer0_outputs(3781) <= not(inputs(137));
    layer0_outputs(3782) <= not(inputs(69));
    layer0_outputs(3783) <= not((inputs(175)) xor (inputs(57)));
    layer0_outputs(3784) <= not(inputs(155));
    layer0_outputs(3785) <= inputs(137);
    layer0_outputs(3786) <= not((inputs(180)) xor (inputs(44)));
    layer0_outputs(3787) <= not(inputs(134)) or (inputs(211));
    layer0_outputs(3788) <= inputs(231);
    layer0_outputs(3789) <= not(inputs(122));
    layer0_outputs(3790) <= not((inputs(22)) or (inputs(246)));
    layer0_outputs(3791) <= not(inputs(50));
    layer0_outputs(3792) <= not(inputs(90)) or (inputs(193));
    layer0_outputs(3793) <= not(inputs(243));
    layer0_outputs(3794) <= not(inputs(122)) or (inputs(182));
    layer0_outputs(3795) <= (inputs(119)) xor (inputs(28));
    layer0_outputs(3796) <= not((inputs(142)) xor (inputs(22)));
    layer0_outputs(3797) <= not((inputs(15)) xor (inputs(124)));
    layer0_outputs(3798) <= inputs(168);
    layer0_outputs(3799) <= not((inputs(200)) xor (inputs(35)));
    layer0_outputs(3800) <= not(inputs(110));
    layer0_outputs(3801) <= inputs(29);
    layer0_outputs(3802) <= not(inputs(182));
    layer0_outputs(3803) <= not(inputs(85)) or (inputs(111));
    layer0_outputs(3804) <= (inputs(218)) or (inputs(197));
    layer0_outputs(3805) <= '1';
    layer0_outputs(3806) <= (inputs(106)) or (inputs(71));
    layer0_outputs(3807) <= inputs(61);
    layer0_outputs(3808) <= inputs(61);
    layer0_outputs(3809) <= (inputs(54)) or (inputs(251));
    layer0_outputs(3810) <= (inputs(135)) and not (inputs(232));
    layer0_outputs(3811) <= not(inputs(94)) or (inputs(146));
    layer0_outputs(3812) <= not((inputs(198)) xor (inputs(31)));
    layer0_outputs(3813) <= inputs(34);
    layer0_outputs(3814) <= not(inputs(99));
    layer0_outputs(3815) <= (inputs(97)) or (inputs(29));
    layer0_outputs(3816) <= (inputs(184)) xor (inputs(222));
    layer0_outputs(3817) <= not(inputs(239)) or (inputs(208));
    layer0_outputs(3818) <= (inputs(129)) or (inputs(107));
    layer0_outputs(3819) <= (inputs(39)) or (inputs(54));
    layer0_outputs(3820) <= not(inputs(167));
    layer0_outputs(3821) <= (inputs(147)) and not (inputs(12));
    layer0_outputs(3822) <= inputs(106);
    layer0_outputs(3823) <= not(inputs(97)) or (inputs(186));
    layer0_outputs(3824) <= (inputs(92)) and not (inputs(71));
    layer0_outputs(3825) <= (inputs(197)) or (inputs(161));
    layer0_outputs(3826) <= (inputs(4)) xor (inputs(134));
    layer0_outputs(3827) <= (inputs(136)) xor (inputs(222));
    layer0_outputs(3828) <= inputs(182);
    layer0_outputs(3829) <= inputs(69);
    layer0_outputs(3830) <= not((inputs(207)) or (inputs(90)));
    layer0_outputs(3831) <= not(inputs(215)) or (inputs(188));
    layer0_outputs(3832) <= inputs(104);
    layer0_outputs(3833) <= not((inputs(178)) or (inputs(239)));
    layer0_outputs(3834) <= not(inputs(138));
    layer0_outputs(3835) <= '1';
    layer0_outputs(3836) <= (inputs(98)) xor (inputs(55));
    layer0_outputs(3837) <= not(inputs(247)) or (inputs(190));
    layer0_outputs(3838) <= (inputs(66)) or (inputs(97));
    layer0_outputs(3839) <= not(inputs(242)) or (inputs(128));
    layer0_outputs(3840) <= not(inputs(188));
    layer0_outputs(3841) <= '0';
    layer0_outputs(3842) <= '1';
    layer0_outputs(3843) <= '1';
    layer0_outputs(3844) <= (inputs(203)) or (inputs(38));
    layer0_outputs(3845) <= (inputs(84)) and not (inputs(175));
    layer0_outputs(3846) <= not((inputs(59)) xor (inputs(161)));
    layer0_outputs(3847) <= (inputs(127)) and not (inputs(233));
    layer0_outputs(3848) <= (inputs(96)) and not (inputs(254));
    layer0_outputs(3849) <= not((inputs(117)) or (inputs(149)));
    layer0_outputs(3850) <= inputs(163);
    layer0_outputs(3851) <= not(inputs(62)) or (inputs(227));
    layer0_outputs(3852) <= (inputs(189)) or (inputs(248));
    layer0_outputs(3853) <= (inputs(123)) and not (inputs(205));
    layer0_outputs(3854) <= (inputs(91)) and not (inputs(212));
    layer0_outputs(3855) <= not((inputs(123)) or (inputs(96)));
    layer0_outputs(3856) <= inputs(90);
    layer0_outputs(3857) <= not((inputs(143)) or (inputs(215)));
    layer0_outputs(3858) <= not(inputs(6)) or (inputs(26));
    layer0_outputs(3859) <= not((inputs(43)) or (inputs(12)));
    layer0_outputs(3860) <= not((inputs(154)) or (inputs(22)));
    layer0_outputs(3861) <= (inputs(248)) and not (inputs(176));
    layer0_outputs(3862) <= not(inputs(203)) or (inputs(246));
    layer0_outputs(3863) <= not(inputs(64)) or (inputs(20));
    layer0_outputs(3864) <= not(inputs(24)) or (inputs(143));
    layer0_outputs(3865) <= inputs(241);
    layer0_outputs(3866) <= inputs(139);
    layer0_outputs(3867) <= not(inputs(211));
    layer0_outputs(3868) <= (inputs(138)) and not (inputs(13));
    layer0_outputs(3869) <= not(inputs(25));
    layer0_outputs(3870) <= not(inputs(105)) or (inputs(100));
    layer0_outputs(3871) <= not((inputs(27)) and (inputs(32)));
    layer0_outputs(3872) <= (inputs(119)) xor (inputs(149));
    layer0_outputs(3873) <= not(inputs(187)) or (inputs(206));
    layer0_outputs(3874) <= (inputs(91)) xor (inputs(0));
    layer0_outputs(3875) <= not((inputs(219)) xor (inputs(231)));
    layer0_outputs(3876) <= not(inputs(31)) or (inputs(48));
    layer0_outputs(3877) <= not(inputs(162)) or (inputs(206));
    layer0_outputs(3878) <= not((inputs(195)) or (inputs(212)));
    layer0_outputs(3879) <= (inputs(236)) xor (inputs(239));
    layer0_outputs(3880) <= (inputs(141)) or (inputs(66));
    layer0_outputs(3881) <= not(inputs(58)) or (inputs(228));
    layer0_outputs(3882) <= not(inputs(212));
    layer0_outputs(3883) <= inputs(200);
    layer0_outputs(3884) <= not(inputs(142)) or (inputs(47));
    layer0_outputs(3885) <= not(inputs(89));
    layer0_outputs(3886) <= not((inputs(122)) xor (inputs(227)));
    layer0_outputs(3887) <= not((inputs(198)) xor (inputs(32)));
    layer0_outputs(3888) <= (inputs(75)) and not (inputs(66));
    layer0_outputs(3889) <= not(inputs(98));
    layer0_outputs(3890) <= not((inputs(81)) xor (inputs(36)));
    layer0_outputs(3891) <= not(inputs(207)) or (inputs(224));
    layer0_outputs(3892) <= not(inputs(74)) or (inputs(44));
    layer0_outputs(3893) <= (inputs(223)) and not (inputs(18));
    layer0_outputs(3894) <= inputs(137);
    layer0_outputs(3895) <= not(inputs(122));
    layer0_outputs(3896) <= not((inputs(119)) or (inputs(13)));
    layer0_outputs(3897) <= (inputs(65)) xor (inputs(135));
    layer0_outputs(3898) <= not(inputs(138));
    layer0_outputs(3899) <= not(inputs(40));
    layer0_outputs(3900) <= not(inputs(188));
    layer0_outputs(3901) <= not((inputs(234)) xor (inputs(152)));
    layer0_outputs(3902) <= (inputs(254)) or (inputs(150));
    layer0_outputs(3903) <= inputs(185);
    layer0_outputs(3904) <= (inputs(134)) and not (inputs(66));
    layer0_outputs(3905) <= (inputs(108)) or (inputs(196));
    layer0_outputs(3906) <= (inputs(162)) or (inputs(213));
    layer0_outputs(3907) <= (inputs(85)) or (inputs(249));
    layer0_outputs(3908) <= not((inputs(44)) xor (inputs(9)));
    layer0_outputs(3909) <= (inputs(252)) and (inputs(176));
    layer0_outputs(3910) <= (inputs(151)) or (inputs(190));
    layer0_outputs(3911) <= (inputs(59)) and not (inputs(249));
    layer0_outputs(3912) <= (inputs(30)) xor (inputs(188));
    layer0_outputs(3913) <= not(inputs(74));
    layer0_outputs(3914) <= not(inputs(159));
    layer0_outputs(3915) <= (inputs(123)) or (inputs(71));
    layer0_outputs(3916) <= not(inputs(62));
    layer0_outputs(3917) <= '0';
    layer0_outputs(3918) <= not((inputs(1)) or (inputs(15)));
    layer0_outputs(3919) <= inputs(117);
    layer0_outputs(3920) <= (inputs(107)) and not (inputs(145));
    layer0_outputs(3921) <= not((inputs(150)) or (inputs(207)));
    layer0_outputs(3922) <= not(inputs(191)) or (inputs(129));
    layer0_outputs(3923) <= (inputs(24)) or (inputs(173));
    layer0_outputs(3924) <= '0';
    layer0_outputs(3925) <= (inputs(93)) or (inputs(58));
    layer0_outputs(3926) <= (inputs(139)) or (inputs(198));
    layer0_outputs(3927) <= not(inputs(109));
    layer0_outputs(3928) <= (inputs(174)) or (inputs(198));
    layer0_outputs(3929) <= (inputs(210)) and not (inputs(97));
    layer0_outputs(3930) <= not((inputs(143)) xor (inputs(100)));
    layer0_outputs(3931) <= inputs(88);
    layer0_outputs(3932) <= (inputs(145)) and (inputs(247));
    layer0_outputs(3933) <= not(inputs(231)) or (inputs(209));
    layer0_outputs(3934) <= not(inputs(42)) or (inputs(222));
    layer0_outputs(3935) <= (inputs(234)) and not (inputs(223));
    layer0_outputs(3936) <= not((inputs(225)) and (inputs(132)));
    layer0_outputs(3937) <= (inputs(198)) xor (inputs(118));
    layer0_outputs(3938) <= not((inputs(80)) or (inputs(11)));
    layer0_outputs(3939) <= (inputs(124)) or (inputs(108));
    layer0_outputs(3940) <= (inputs(93)) or (inputs(67));
    layer0_outputs(3941) <= '1';
    layer0_outputs(3942) <= not(inputs(67));
    layer0_outputs(3943) <= (inputs(100)) and not (inputs(103));
    layer0_outputs(3944) <= not(inputs(120));
    layer0_outputs(3945) <= (inputs(158)) and not (inputs(48));
    layer0_outputs(3946) <= '1';
    layer0_outputs(3947) <= (inputs(105)) and (inputs(120));
    layer0_outputs(3948) <= not(inputs(53)) or (inputs(204));
    layer0_outputs(3949) <= (inputs(202)) and not (inputs(140));
    layer0_outputs(3950) <= (inputs(38)) and not (inputs(2));
    layer0_outputs(3951) <= not(inputs(35)) or (inputs(140));
    layer0_outputs(3952) <= (inputs(102)) and not (inputs(67));
    layer0_outputs(3953) <= (inputs(135)) xor (inputs(39));
    layer0_outputs(3954) <= (inputs(29)) and (inputs(110));
    layer0_outputs(3955) <= (inputs(225)) and not (inputs(65));
    layer0_outputs(3956) <= not((inputs(93)) xor (inputs(248)));
    layer0_outputs(3957) <= (inputs(81)) or (inputs(77));
    layer0_outputs(3958) <= inputs(182);
    layer0_outputs(3959) <= (inputs(21)) and not (inputs(254));
    layer0_outputs(3960) <= not((inputs(225)) xor (inputs(14)));
    layer0_outputs(3961) <= inputs(119);
    layer0_outputs(3962) <= (inputs(71)) xor (inputs(72));
    layer0_outputs(3963) <= not(inputs(75));
    layer0_outputs(3964) <= '1';
    layer0_outputs(3965) <= (inputs(32)) xor (inputs(166));
    layer0_outputs(3966) <= (inputs(203)) and not (inputs(95));
    layer0_outputs(3967) <= (inputs(169)) and not (inputs(71));
    layer0_outputs(3968) <= (inputs(239)) xor (inputs(182));
    layer0_outputs(3969) <= (inputs(200)) or (inputs(211));
    layer0_outputs(3970) <= not(inputs(195));
    layer0_outputs(3971) <= not(inputs(227));
    layer0_outputs(3972) <= inputs(76);
    layer0_outputs(3973) <= not((inputs(112)) xor (inputs(188)));
    layer0_outputs(3974) <= not((inputs(112)) or (inputs(104)));
    layer0_outputs(3975) <= (inputs(76)) or (inputs(119));
    layer0_outputs(3976) <= (inputs(94)) and not (inputs(224));
    layer0_outputs(3977) <= not(inputs(170)) or (inputs(234));
    layer0_outputs(3978) <= (inputs(197)) xor (inputs(236));
    layer0_outputs(3979) <= inputs(67);
    layer0_outputs(3980) <= not((inputs(232)) or (inputs(66)));
    layer0_outputs(3981) <= not(inputs(219)) or (inputs(175));
    layer0_outputs(3982) <= (inputs(161)) and (inputs(236));
    layer0_outputs(3983) <= '1';
    layer0_outputs(3984) <= not(inputs(72));
    layer0_outputs(3985) <= (inputs(62)) or (inputs(112));
    layer0_outputs(3986) <= (inputs(216)) xor (inputs(25));
    layer0_outputs(3987) <= not((inputs(67)) and (inputs(174)));
    layer0_outputs(3988) <= not(inputs(185));
    layer0_outputs(3989) <= (inputs(217)) and not (inputs(250));
    layer0_outputs(3990) <= not(inputs(75)) or (inputs(235));
    layer0_outputs(3991) <= not((inputs(117)) xor (inputs(34)));
    layer0_outputs(3992) <= (inputs(182)) and not (inputs(145));
    layer0_outputs(3993) <= inputs(71);
    layer0_outputs(3994) <= (inputs(144)) or (inputs(170));
    layer0_outputs(3995) <= (inputs(242)) xor (inputs(70));
    layer0_outputs(3996) <= not((inputs(16)) xor (inputs(57)));
    layer0_outputs(3997) <= (inputs(227)) and (inputs(70));
    layer0_outputs(3998) <= not((inputs(30)) or (inputs(38)));
    layer0_outputs(3999) <= not((inputs(73)) and (inputs(235)));
    layer0_outputs(4000) <= inputs(183);
    layer0_outputs(4001) <= not((inputs(207)) xor (inputs(133)));
    layer0_outputs(4002) <= not((inputs(111)) xor (inputs(126)));
    layer0_outputs(4003) <= (inputs(225)) xor (inputs(123));
    layer0_outputs(4004) <= not(inputs(136)) or (inputs(31));
    layer0_outputs(4005) <= (inputs(195)) or (inputs(199));
    layer0_outputs(4006) <= not(inputs(86));
    layer0_outputs(4007) <= (inputs(208)) xor (inputs(107));
    layer0_outputs(4008) <= not(inputs(238));
    layer0_outputs(4009) <= not((inputs(200)) and (inputs(91)));
    layer0_outputs(4010) <= inputs(29);
    layer0_outputs(4011) <= (inputs(121)) and not (inputs(24));
    layer0_outputs(4012) <= not(inputs(145));
    layer0_outputs(4013) <= not(inputs(118)) or (inputs(158));
    layer0_outputs(4014) <= not(inputs(84));
    layer0_outputs(4015) <= not(inputs(25)) or (inputs(218));
    layer0_outputs(4016) <= (inputs(17)) xor (inputs(219));
    layer0_outputs(4017) <= (inputs(17)) or (inputs(42));
    layer0_outputs(4018) <= not(inputs(160));
    layer0_outputs(4019) <= not((inputs(201)) xor (inputs(80)));
    layer0_outputs(4020) <= not((inputs(128)) or (inputs(165)));
    layer0_outputs(4021) <= (inputs(39)) or (inputs(118));
    layer0_outputs(4022) <= (inputs(1)) xor (inputs(229));
    layer0_outputs(4023) <= inputs(198);
    layer0_outputs(4024) <= not((inputs(67)) xor (inputs(252)));
    layer0_outputs(4025) <= '0';
    layer0_outputs(4026) <= inputs(121);
    layer0_outputs(4027) <= not(inputs(185)) or (inputs(4));
    layer0_outputs(4028) <= not(inputs(62)) or (inputs(207));
    layer0_outputs(4029) <= not((inputs(234)) or (inputs(204)));
    layer0_outputs(4030) <= not(inputs(234)) or (inputs(158));
    layer0_outputs(4031) <= not((inputs(79)) and (inputs(237)));
    layer0_outputs(4032) <= not((inputs(224)) xor (inputs(169)));
    layer0_outputs(4033) <= not((inputs(63)) or (inputs(177)));
    layer0_outputs(4034) <= (inputs(93)) or (inputs(202));
    layer0_outputs(4035) <= not((inputs(220)) or (inputs(207)));
    layer0_outputs(4036) <= inputs(174);
    layer0_outputs(4037) <= (inputs(10)) or (inputs(39));
    layer0_outputs(4038) <= inputs(38);
    layer0_outputs(4039) <= not(inputs(72)) or (inputs(217));
    layer0_outputs(4040) <= not(inputs(197)) or (inputs(34));
    layer0_outputs(4041) <= (inputs(7)) xor (inputs(180));
    layer0_outputs(4042) <= not(inputs(167));
    layer0_outputs(4043) <= '0';
    layer0_outputs(4044) <= not(inputs(175)) or (inputs(50));
    layer0_outputs(4045) <= (inputs(149)) or (inputs(189));
    layer0_outputs(4046) <= not((inputs(118)) or (inputs(11)));
    layer0_outputs(4047) <= (inputs(55)) or (inputs(245));
    layer0_outputs(4048) <= (inputs(74)) or (inputs(179));
    layer0_outputs(4049) <= inputs(54);
    layer0_outputs(4050) <= (inputs(81)) xor (inputs(28));
    layer0_outputs(4051) <= (inputs(131)) and not (inputs(17));
    layer0_outputs(4052) <= (inputs(161)) xor (inputs(109));
    layer0_outputs(4053) <= inputs(44);
    layer0_outputs(4054) <= (inputs(233)) xor (inputs(217));
    layer0_outputs(4055) <= not(inputs(126)) or (inputs(128));
    layer0_outputs(4056) <= not(inputs(195));
    layer0_outputs(4057) <= not((inputs(33)) xor (inputs(59)));
    layer0_outputs(4058) <= inputs(221);
    layer0_outputs(4059) <= not(inputs(122));
    layer0_outputs(4060) <= not(inputs(198)) or (inputs(131));
    layer0_outputs(4061) <= (inputs(30)) and not (inputs(114));
    layer0_outputs(4062) <= not((inputs(180)) xor (inputs(183)));
    layer0_outputs(4063) <= not(inputs(253));
    layer0_outputs(4064) <= not(inputs(4)) or (inputs(158));
    layer0_outputs(4065) <= not((inputs(86)) xor (inputs(76)));
    layer0_outputs(4066) <= not((inputs(31)) and (inputs(112)));
    layer0_outputs(4067) <= (inputs(179)) or (inputs(21));
    layer0_outputs(4068) <= not((inputs(200)) xor (inputs(98)));
    layer0_outputs(4069) <= not(inputs(74)) or (inputs(180));
    layer0_outputs(4070) <= not(inputs(229));
    layer0_outputs(4071) <= inputs(134);
    layer0_outputs(4072) <= not((inputs(172)) or (inputs(63)));
    layer0_outputs(4073) <= '1';
    layer0_outputs(4074) <= not(inputs(27));
    layer0_outputs(4075) <= inputs(12);
    layer0_outputs(4076) <= (inputs(171)) and not (inputs(84));
    layer0_outputs(4077) <= not((inputs(40)) or (inputs(56)));
    layer0_outputs(4078) <= (inputs(246)) and (inputs(16));
    layer0_outputs(4079) <= not(inputs(105));
    layer0_outputs(4080) <= (inputs(186)) and not (inputs(48));
    layer0_outputs(4081) <= not((inputs(192)) or (inputs(196)));
    layer0_outputs(4082) <= (inputs(169)) or (inputs(95));
    layer0_outputs(4083) <= '0';
    layer0_outputs(4084) <= (inputs(117)) or (inputs(138));
    layer0_outputs(4085) <= (inputs(161)) or (inputs(92));
    layer0_outputs(4086) <= (inputs(78)) and not (inputs(252));
    layer0_outputs(4087) <= not(inputs(201));
    layer0_outputs(4088) <= (inputs(103)) xor (inputs(221));
    layer0_outputs(4089) <= not((inputs(150)) xor (inputs(157)));
    layer0_outputs(4090) <= (inputs(93)) xor (inputs(81));
    layer0_outputs(4091) <= inputs(180);
    layer0_outputs(4092) <= (inputs(90)) xor (inputs(251));
    layer0_outputs(4093) <= not(inputs(158));
    layer0_outputs(4094) <= not(inputs(66));
    layer0_outputs(4095) <= (inputs(173)) and (inputs(202));
    layer0_outputs(4096) <= (inputs(112)) and not (inputs(127));
    layer0_outputs(4097) <= inputs(19);
    layer0_outputs(4098) <= not((inputs(115)) or (inputs(134)));
    layer0_outputs(4099) <= (inputs(12)) or (inputs(94));
    layer0_outputs(4100) <= not(inputs(67)) or (inputs(133));
    layer0_outputs(4101) <= not((inputs(231)) and (inputs(59)));
    layer0_outputs(4102) <= (inputs(43)) or (inputs(104));
    layer0_outputs(4103) <= inputs(139);
    layer0_outputs(4104) <= (inputs(12)) xor (inputs(0));
    layer0_outputs(4105) <= not(inputs(102));
    layer0_outputs(4106) <= not((inputs(191)) or (inputs(137)));
    layer0_outputs(4107) <= (inputs(210)) xor (inputs(125));
    layer0_outputs(4108) <= not(inputs(214));
    layer0_outputs(4109) <= inputs(91);
    layer0_outputs(4110) <= not((inputs(191)) xor (inputs(118)));
    layer0_outputs(4111) <= (inputs(220)) and not (inputs(156));
    layer0_outputs(4112) <= inputs(25);
    layer0_outputs(4113) <= not(inputs(13)) or (inputs(222));
    layer0_outputs(4114) <= not((inputs(139)) xor (inputs(230)));
    layer0_outputs(4115) <= not((inputs(127)) or (inputs(227)));
    layer0_outputs(4116) <= not((inputs(73)) or (inputs(179)));
    layer0_outputs(4117) <= not((inputs(196)) xor (inputs(49)));
    layer0_outputs(4118) <= not(inputs(139));
    layer0_outputs(4119) <= not((inputs(255)) or (inputs(32)));
    layer0_outputs(4120) <= (inputs(216)) xor (inputs(125));
    layer0_outputs(4121) <= (inputs(13)) and not (inputs(221));
    layer0_outputs(4122) <= '1';
    layer0_outputs(4123) <= (inputs(239)) and not (inputs(64));
    layer0_outputs(4124) <= (inputs(159)) xor (inputs(156));
    layer0_outputs(4125) <= (inputs(128)) or (inputs(237));
    layer0_outputs(4126) <= not(inputs(61));
    layer0_outputs(4127) <= not(inputs(186));
    layer0_outputs(4128) <= (inputs(46)) and not (inputs(192));
    layer0_outputs(4129) <= inputs(75);
    layer0_outputs(4130) <= (inputs(200)) and not (inputs(36));
    layer0_outputs(4131) <= (inputs(118)) and not (inputs(209));
    layer0_outputs(4132) <= not(inputs(151));
    layer0_outputs(4133) <= (inputs(182)) or (inputs(179));
    layer0_outputs(4134) <= not((inputs(82)) or (inputs(161)));
    layer0_outputs(4135) <= inputs(140);
    layer0_outputs(4136) <= inputs(166);
    layer0_outputs(4137) <= not((inputs(253)) xor (inputs(0)));
    layer0_outputs(4138) <= not(inputs(183));
    layer0_outputs(4139) <= not((inputs(78)) xor (inputs(28)));
    layer0_outputs(4140) <= (inputs(89)) and not (inputs(14));
    layer0_outputs(4141) <= not(inputs(68)) or (inputs(240));
    layer0_outputs(4142) <= inputs(110);
    layer0_outputs(4143) <= not(inputs(201));
    layer0_outputs(4144) <= not(inputs(44));
    layer0_outputs(4145) <= (inputs(18)) xor (inputs(29));
    layer0_outputs(4146) <= (inputs(246)) or (inputs(156));
    layer0_outputs(4147) <= (inputs(27)) xor (inputs(122));
    layer0_outputs(4148) <= not((inputs(157)) or (inputs(0)));
    layer0_outputs(4149) <= (inputs(55)) or (inputs(53));
    layer0_outputs(4150) <= (inputs(92)) and (inputs(74));
    layer0_outputs(4151) <= not((inputs(60)) or (inputs(231)));
    layer0_outputs(4152) <= inputs(123);
    layer0_outputs(4153) <= not((inputs(199)) or (inputs(0)));
    layer0_outputs(4154) <= not(inputs(212));
    layer0_outputs(4155) <= (inputs(103)) or (inputs(118));
    layer0_outputs(4156) <= (inputs(75)) and not (inputs(158));
    layer0_outputs(4157) <= inputs(4);
    layer0_outputs(4158) <= (inputs(154)) and not (inputs(195));
    layer0_outputs(4159) <= (inputs(245)) xor (inputs(153));
    layer0_outputs(4160) <= inputs(198);
    layer0_outputs(4161) <= not(inputs(122));
    layer0_outputs(4162) <= (inputs(18)) and not (inputs(225));
    layer0_outputs(4163) <= not(inputs(56));
    layer0_outputs(4164) <= not(inputs(105));
    layer0_outputs(4165) <= not((inputs(135)) xor (inputs(87)));
    layer0_outputs(4166) <= not((inputs(82)) or (inputs(187)));
    layer0_outputs(4167) <= not(inputs(122));
    layer0_outputs(4168) <= inputs(122);
    layer0_outputs(4169) <= (inputs(250)) and (inputs(238));
    layer0_outputs(4170) <= '1';
    layer0_outputs(4171) <= (inputs(169)) and not (inputs(220));
    layer0_outputs(4172) <= inputs(38);
    layer0_outputs(4173) <= (inputs(132)) or (inputs(6));
    layer0_outputs(4174) <= not(inputs(105)) or (inputs(133));
    layer0_outputs(4175) <= not((inputs(8)) xor (inputs(48)));
    layer0_outputs(4176) <= not(inputs(68));
    layer0_outputs(4177) <= not((inputs(95)) xor (inputs(180)));
    layer0_outputs(4178) <= not(inputs(152)) or (inputs(24));
    layer0_outputs(4179) <= not(inputs(125));
    layer0_outputs(4180) <= inputs(156);
    layer0_outputs(4181) <= not((inputs(1)) xor (inputs(151)));
    layer0_outputs(4182) <= (inputs(89)) xor (inputs(177));
    layer0_outputs(4183) <= not((inputs(26)) xor (inputs(112)));
    layer0_outputs(4184) <= (inputs(62)) or (inputs(250));
    layer0_outputs(4185) <= (inputs(35)) xor (inputs(42));
    layer0_outputs(4186) <= not(inputs(40));
    layer0_outputs(4187) <= not((inputs(206)) or (inputs(240)));
    layer0_outputs(4188) <= not(inputs(137)) or (inputs(46));
    layer0_outputs(4189) <= not((inputs(206)) or (inputs(195)));
    layer0_outputs(4190) <= not(inputs(100)) or (inputs(187));
    layer0_outputs(4191) <= inputs(3);
    layer0_outputs(4192) <= inputs(227);
    layer0_outputs(4193) <= inputs(28);
    layer0_outputs(4194) <= (inputs(133)) or (inputs(115));
    layer0_outputs(4195) <= not(inputs(74)) or (inputs(239));
    layer0_outputs(4196) <= (inputs(174)) and not (inputs(7));
    layer0_outputs(4197) <= (inputs(51)) and not (inputs(255));
    layer0_outputs(4198) <= not(inputs(171)) or (inputs(90));
    layer0_outputs(4199) <= not(inputs(5)) or (inputs(144));
    layer0_outputs(4200) <= (inputs(235)) and not (inputs(173));
    layer0_outputs(4201) <= not(inputs(121)) or (inputs(157));
    layer0_outputs(4202) <= (inputs(129)) or (inputs(85));
    layer0_outputs(4203) <= not(inputs(46));
    layer0_outputs(4204) <= (inputs(42)) xor (inputs(220));
    layer0_outputs(4205) <= not((inputs(42)) or (inputs(181)));
    layer0_outputs(4206) <= not((inputs(223)) and (inputs(192)));
    layer0_outputs(4207) <= (inputs(59)) or (inputs(190));
    layer0_outputs(4208) <= (inputs(78)) or (inputs(122));
    layer0_outputs(4209) <= not(inputs(137));
    layer0_outputs(4210) <= not((inputs(20)) xor (inputs(26)));
    layer0_outputs(4211) <= (inputs(46)) xor (inputs(232));
    layer0_outputs(4212) <= (inputs(103)) and not (inputs(32));
    layer0_outputs(4213) <= (inputs(101)) and not (inputs(83));
    layer0_outputs(4214) <= (inputs(218)) and not (inputs(229));
    layer0_outputs(4215) <= (inputs(163)) or (inputs(79));
    layer0_outputs(4216) <= (inputs(21)) xor (inputs(184));
    layer0_outputs(4217) <= not(inputs(213)) or (inputs(22));
    layer0_outputs(4218) <= inputs(130);
    layer0_outputs(4219) <= not(inputs(151));
    layer0_outputs(4220) <= (inputs(48)) xor (inputs(115));
    layer0_outputs(4221) <= not((inputs(187)) or (inputs(171)));
    layer0_outputs(4222) <= (inputs(105)) or (inputs(246));
    layer0_outputs(4223) <= (inputs(166)) and not (inputs(91));
    layer0_outputs(4224) <= inputs(56);
    layer0_outputs(4225) <= not((inputs(202)) xor (inputs(82)));
    layer0_outputs(4226) <= (inputs(174)) xor (inputs(169));
    layer0_outputs(4227) <= not((inputs(35)) or (inputs(187)));
    layer0_outputs(4228) <= not(inputs(71)) or (inputs(220));
    layer0_outputs(4229) <= (inputs(165)) or (inputs(216));
    layer0_outputs(4230) <= (inputs(183)) and not (inputs(106));
    layer0_outputs(4231) <= inputs(219);
    layer0_outputs(4232) <= not(inputs(196)) or (inputs(162));
    layer0_outputs(4233) <= inputs(153);
    layer0_outputs(4234) <= (inputs(17)) xor (inputs(152));
    layer0_outputs(4235) <= not(inputs(44));
    layer0_outputs(4236) <= (inputs(26)) xor (inputs(104));
    layer0_outputs(4237) <= '0';
    layer0_outputs(4238) <= (inputs(135)) or (inputs(223));
    layer0_outputs(4239) <= not(inputs(134));
    layer0_outputs(4240) <= inputs(166);
    layer0_outputs(4241) <= not(inputs(60));
    layer0_outputs(4242) <= not((inputs(210)) or (inputs(106)));
    layer0_outputs(4243) <= inputs(119);
    layer0_outputs(4244) <= not(inputs(44)) or (inputs(176));
    layer0_outputs(4245) <= not((inputs(209)) xor (inputs(98)));
    layer0_outputs(4246) <= (inputs(82)) xor (inputs(162));
    layer0_outputs(4247) <= not(inputs(2)) or (inputs(81));
    layer0_outputs(4248) <= not((inputs(100)) xor (inputs(61)));
    layer0_outputs(4249) <= not((inputs(199)) xor (inputs(34)));
    layer0_outputs(4250) <= '0';
    layer0_outputs(4251) <= not((inputs(188)) xor (inputs(87)));
    layer0_outputs(4252) <= not(inputs(146)) or (inputs(236));
    layer0_outputs(4253) <= (inputs(38)) or (inputs(35));
    layer0_outputs(4254) <= (inputs(149)) and not (inputs(84));
    layer0_outputs(4255) <= not(inputs(12)) or (inputs(221));
    layer0_outputs(4256) <= not(inputs(156)) or (inputs(36));
    layer0_outputs(4257) <= inputs(151);
    layer0_outputs(4258) <= not((inputs(83)) xor (inputs(14)));
    layer0_outputs(4259) <= not(inputs(58));
    layer0_outputs(4260) <= inputs(143);
    layer0_outputs(4261) <= inputs(137);
    layer0_outputs(4262) <= '1';
    layer0_outputs(4263) <= not((inputs(176)) xor (inputs(123)));
    layer0_outputs(4264) <= not(inputs(127));
    layer0_outputs(4265) <= '0';
    layer0_outputs(4266) <= not(inputs(100)) or (inputs(31));
    layer0_outputs(4267) <= (inputs(15)) xor (inputs(43));
    layer0_outputs(4268) <= (inputs(79)) or (inputs(193));
    layer0_outputs(4269) <= inputs(195);
    layer0_outputs(4270) <= '1';
    layer0_outputs(4271) <= not(inputs(219)) or (inputs(236));
    layer0_outputs(4272) <= not((inputs(107)) or (inputs(37)));
    layer0_outputs(4273) <= (inputs(177)) or (inputs(142));
    layer0_outputs(4274) <= not(inputs(68));
    layer0_outputs(4275) <= (inputs(169)) xor (inputs(246));
    layer0_outputs(4276) <= not(inputs(150));
    layer0_outputs(4277) <= not((inputs(114)) or (inputs(206)));
    layer0_outputs(4278) <= not(inputs(56));
    layer0_outputs(4279) <= not((inputs(150)) xor (inputs(95)));
    layer0_outputs(4280) <= (inputs(170)) and not (inputs(155));
    layer0_outputs(4281) <= not((inputs(223)) or (inputs(69)));
    layer0_outputs(4282) <= (inputs(201)) xor (inputs(88));
    layer0_outputs(4283) <= (inputs(86)) xor (inputs(40));
    layer0_outputs(4284) <= not(inputs(139)) or (inputs(220));
    layer0_outputs(4285) <= inputs(122);
    layer0_outputs(4286) <= (inputs(146)) xor (inputs(158));
    layer0_outputs(4287) <= '1';
    layer0_outputs(4288) <= not((inputs(162)) xor (inputs(112)));
    layer0_outputs(4289) <= inputs(136);
    layer0_outputs(4290) <= not(inputs(164)) or (inputs(130));
    layer0_outputs(4291) <= not((inputs(16)) or (inputs(188)));
    layer0_outputs(4292) <= not(inputs(72)) or (inputs(143));
    layer0_outputs(4293) <= (inputs(152)) and not (inputs(67));
    layer0_outputs(4294) <= not(inputs(186)) or (inputs(15));
    layer0_outputs(4295) <= not((inputs(37)) xor (inputs(231)));
    layer0_outputs(4296) <= not((inputs(189)) or (inputs(73)));
    layer0_outputs(4297) <= (inputs(122)) or (inputs(210));
    layer0_outputs(4298) <= not(inputs(90));
    layer0_outputs(4299) <= not(inputs(233)) or (inputs(67));
    layer0_outputs(4300) <= not(inputs(125));
    layer0_outputs(4301) <= not((inputs(146)) or (inputs(202)));
    layer0_outputs(4302) <= not(inputs(154)) or (inputs(146));
    layer0_outputs(4303) <= (inputs(46)) xor (inputs(26));
    layer0_outputs(4304) <= inputs(12);
    layer0_outputs(4305) <= (inputs(160)) or (inputs(85));
    layer0_outputs(4306) <= inputs(211);
    layer0_outputs(4307) <= (inputs(87)) xor (inputs(163));
    layer0_outputs(4308) <= not(inputs(190));
    layer0_outputs(4309) <= (inputs(158)) xor (inputs(99));
    layer0_outputs(4310) <= not(inputs(167));
    layer0_outputs(4311) <= not(inputs(60));
    layer0_outputs(4312) <= (inputs(202)) and not (inputs(35));
    layer0_outputs(4313) <= inputs(105);
    layer0_outputs(4314) <= inputs(229);
    layer0_outputs(4315) <= (inputs(254)) or (inputs(161));
    layer0_outputs(4316) <= (inputs(55)) and not (inputs(125));
    layer0_outputs(4317) <= not(inputs(128)) or (inputs(115));
    layer0_outputs(4318) <= (inputs(134)) or (inputs(252));
    layer0_outputs(4319) <= inputs(77);
    layer0_outputs(4320) <= (inputs(106)) and not (inputs(171));
    layer0_outputs(4321) <= not((inputs(74)) xor (inputs(8)));
    layer0_outputs(4322) <= not((inputs(88)) or (inputs(211)));
    layer0_outputs(4323) <= (inputs(213)) and not (inputs(27));
    layer0_outputs(4324) <= (inputs(180)) xor (inputs(175));
    layer0_outputs(4325) <= not(inputs(91)) or (inputs(235));
    layer0_outputs(4326) <= not(inputs(57));
    layer0_outputs(4327) <= inputs(14);
    layer0_outputs(4328) <= inputs(125);
    layer0_outputs(4329) <= (inputs(51)) or (inputs(68));
    layer0_outputs(4330) <= '0';
    layer0_outputs(4331) <= inputs(139);
    layer0_outputs(4332) <= (inputs(55)) and (inputs(242));
    layer0_outputs(4333) <= not(inputs(133)) or (inputs(82));
    layer0_outputs(4334) <= not(inputs(198));
    layer0_outputs(4335) <= not((inputs(24)) xor (inputs(77)));
    layer0_outputs(4336) <= '1';
    layer0_outputs(4337) <= not(inputs(127)) or (inputs(45));
    layer0_outputs(4338) <= not(inputs(131)) or (inputs(176));
    layer0_outputs(4339) <= not((inputs(2)) or (inputs(121)));
    layer0_outputs(4340) <= (inputs(78)) and not (inputs(175));
    layer0_outputs(4341) <= not(inputs(73)) or (inputs(18));
    layer0_outputs(4342) <= not((inputs(129)) xor (inputs(68)));
    layer0_outputs(4343) <= inputs(154);
    layer0_outputs(4344) <= not(inputs(164)) or (inputs(200));
    layer0_outputs(4345) <= not((inputs(139)) xor (inputs(165)));
    layer0_outputs(4346) <= '1';
    layer0_outputs(4347) <= not((inputs(136)) or (inputs(66)));
    layer0_outputs(4348) <= not(inputs(118));
    layer0_outputs(4349) <= inputs(167);
    layer0_outputs(4350) <= (inputs(213)) and not (inputs(183));
    layer0_outputs(4351) <= (inputs(182)) or (inputs(62));
    layer0_outputs(4352) <= (inputs(28)) and not (inputs(35));
    layer0_outputs(4353) <= (inputs(124)) and (inputs(206));
    layer0_outputs(4354) <= not(inputs(245));
    layer0_outputs(4355) <= not(inputs(61));
    layer0_outputs(4356) <= (inputs(55)) and not (inputs(99));
    layer0_outputs(4357) <= (inputs(8)) and not (inputs(238));
    layer0_outputs(4358) <= (inputs(139)) or (inputs(85));
    layer0_outputs(4359) <= (inputs(205)) and not (inputs(98));
    layer0_outputs(4360) <= not((inputs(223)) xor (inputs(204)));
    layer0_outputs(4361) <= not(inputs(52));
    layer0_outputs(4362) <= not((inputs(110)) or (inputs(116)));
    layer0_outputs(4363) <= (inputs(52)) and (inputs(67));
    layer0_outputs(4364) <= not((inputs(233)) or (inputs(68)));
    layer0_outputs(4365) <= inputs(183);
    layer0_outputs(4366) <= (inputs(238)) and not (inputs(29));
    layer0_outputs(4367) <= (inputs(240)) and not (inputs(62));
    layer0_outputs(4368) <= not(inputs(217)) or (inputs(222));
    layer0_outputs(4369) <= not(inputs(89));
    layer0_outputs(4370) <= not((inputs(157)) xor (inputs(254)));
    layer0_outputs(4371) <= (inputs(148)) or (inputs(251));
    layer0_outputs(4372) <= (inputs(58)) and not (inputs(110));
    layer0_outputs(4373) <= not((inputs(121)) or (inputs(232)));
    layer0_outputs(4374) <= '0';
    layer0_outputs(4375) <= not((inputs(174)) xor (inputs(15)));
    layer0_outputs(4376) <= not((inputs(170)) xor (inputs(213)));
    layer0_outputs(4377) <= (inputs(193)) xor (inputs(71));
    layer0_outputs(4378) <= not((inputs(94)) xor (inputs(130)));
    layer0_outputs(4379) <= (inputs(67)) and not (inputs(80));
    layer0_outputs(4380) <= not(inputs(28)) or (inputs(242));
    layer0_outputs(4381) <= (inputs(173)) and (inputs(32));
    layer0_outputs(4382) <= (inputs(173)) and not (inputs(0));
    layer0_outputs(4383) <= (inputs(29)) and not (inputs(127));
    layer0_outputs(4384) <= inputs(29);
    layer0_outputs(4385) <= not(inputs(180));
    layer0_outputs(4386) <= not(inputs(100));
    layer0_outputs(4387) <= (inputs(51)) and not (inputs(5));
    layer0_outputs(4388) <= (inputs(91)) or (inputs(239));
    layer0_outputs(4389) <= not((inputs(68)) or (inputs(113)));
    layer0_outputs(4390) <= (inputs(215)) xor (inputs(217));
    layer0_outputs(4391) <= '1';
    layer0_outputs(4392) <= not((inputs(55)) and (inputs(56)));
    layer0_outputs(4393) <= not((inputs(219)) xor (inputs(21)));
    layer0_outputs(4394) <= not(inputs(107));
    layer0_outputs(4395) <= inputs(87);
    layer0_outputs(4396) <= (inputs(14)) and (inputs(234));
    layer0_outputs(4397) <= (inputs(176)) and not (inputs(183));
    layer0_outputs(4398) <= (inputs(60)) or (inputs(197));
    layer0_outputs(4399) <= (inputs(34)) and not (inputs(217));
    layer0_outputs(4400) <= not(inputs(201)) or (inputs(146));
    layer0_outputs(4401) <= not(inputs(214)) or (inputs(190));
    layer0_outputs(4402) <= (inputs(56)) and not (inputs(175));
    layer0_outputs(4403) <= not(inputs(167));
    layer0_outputs(4404) <= (inputs(190)) and not (inputs(248));
    layer0_outputs(4405) <= not((inputs(137)) and (inputs(222)));
    layer0_outputs(4406) <= not(inputs(150)) or (inputs(48));
    layer0_outputs(4407) <= not((inputs(49)) or (inputs(45)));
    layer0_outputs(4408) <= not((inputs(243)) or (inputs(185)));
    layer0_outputs(4409) <= inputs(139);
    layer0_outputs(4410) <= not((inputs(154)) or (inputs(20)));
    layer0_outputs(4411) <= not((inputs(156)) or (inputs(95)));
    layer0_outputs(4412) <= (inputs(8)) or (inputs(217));
    layer0_outputs(4413) <= (inputs(100)) xor (inputs(9));
    layer0_outputs(4414) <= not(inputs(69));
    layer0_outputs(4415) <= (inputs(145)) and not (inputs(57));
    layer0_outputs(4416) <= (inputs(214)) and not (inputs(220));
    layer0_outputs(4417) <= not(inputs(101));
    layer0_outputs(4418) <= (inputs(177)) or (inputs(155));
    layer0_outputs(4419) <= (inputs(137)) and not (inputs(21));
    layer0_outputs(4420) <= not((inputs(249)) xor (inputs(167)));
    layer0_outputs(4421) <= (inputs(83)) and not (inputs(18));
    layer0_outputs(4422) <= not(inputs(148)) or (inputs(111));
    layer0_outputs(4423) <= not(inputs(200)) or (inputs(0));
    layer0_outputs(4424) <= (inputs(33)) or (inputs(226));
    layer0_outputs(4425) <= (inputs(57)) or (inputs(187));
    layer0_outputs(4426) <= not(inputs(54));
    layer0_outputs(4427) <= not((inputs(93)) xor (inputs(218)));
    layer0_outputs(4428) <= (inputs(9)) or (inputs(168));
    layer0_outputs(4429) <= inputs(174);
    layer0_outputs(4430) <= (inputs(221)) and (inputs(146));
    layer0_outputs(4431) <= not((inputs(127)) xor (inputs(239)));
    layer0_outputs(4432) <= inputs(104);
    layer0_outputs(4433) <= (inputs(139)) and (inputs(16));
    layer0_outputs(4434) <= not(inputs(151));
    layer0_outputs(4435) <= (inputs(34)) xor (inputs(20));
    layer0_outputs(4436) <= inputs(106);
    layer0_outputs(4437) <= (inputs(5)) or (inputs(40));
    layer0_outputs(4438) <= inputs(56);
    layer0_outputs(4439) <= not(inputs(104));
    layer0_outputs(4440) <= not((inputs(8)) or (inputs(171)));
    layer0_outputs(4441) <= not((inputs(70)) xor (inputs(26)));
    layer0_outputs(4442) <= (inputs(208)) xor (inputs(168));
    layer0_outputs(4443) <= '1';
    layer0_outputs(4444) <= (inputs(22)) and not (inputs(79));
    layer0_outputs(4445) <= inputs(190);
    layer0_outputs(4446) <= not(inputs(199)) or (inputs(39));
    layer0_outputs(4447) <= not(inputs(25)) or (inputs(73));
    layer0_outputs(4448) <= not((inputs(74)) or (inputs(176)));
    layer0_outputs(4449) <= inputs(243);
    layer0_outputs(4450) <= (inputs(25)) or (inputs(13));
    layer0_outputs(4451) <= not((inputs(188)) or (inputs(71)));
    layer0_outputs(4452) <= not((inputs(81)) xor (inputs(178)));
    layer0_outputs(4453) <= not(inputs(203)) or (inputs(82));
    layer0_outputs(4454) <= not((inputs(198)) xor (inputs(4)));
    layer0_outputs(4455) <= not(inputs(108));
    layer0_outputs(4456) <= (inputs(136)) and not (inputs(232));
    layer0_outputs(4457) <= (inputs(118)) xor (inputs(141));
    layer0_outputs(4458) <= (inputs(133)) xor (inputs(161));
    layer0_outputs(4459) <= not((inputs(69)) or (inputs(186)));
    layer0_outputs(4460) <= not((inputs(226)) or (inputs(215)));
    layer0_outputs(4461) <= not((inputs(28)) or (inputs(201)));
    layer0_outputs(4462) <= not(inputs(15));
    layer0_outputs(4463) <= not((inputs(211)) xor (inputs(112)));
    layer0_outputs(4464) <= (inputs(219)) and not (inputs(127));
    layer0_outputs(4465) <= not((inputs(22)) or (inputs(143)));
    layer0_outputs(4466) <= (inputs(166)) xor (inputs(96));
    layer0_outputs(4467) <= (inputs(111)) and not (inputs(161));
    layer0_outputs(4468) <= (inputs(248)) and not (inputs(112));
    layer0_outputs(4469) <= (inputs(215)) and not (inputs(0));
    layer0_outputs(4470) <= inputs(76);
    layer0_outputs(4471) <= (inputs(137)) and not (inputs(82));
    layer0_outputs(4472) <= inputs(139);
    layer0_outputs(4473) <= not((inputs(173)) xor (inputs(66)));
    layer0_outputs(4474) <= (inputs(231)) xor (inputs(218));
    layer0_outputs(4475) <= (inputs(121)) xor (inputs(227));
    layer0_outputs(4476) <= (inputs(196)) or (inputs(57));
    layer0_outputs(4477) <= inputs(134);
    layer0_outputs(4478) <= (inputs(77)) and not (inputs(142));
    layer0_outputs(4479) <= not(inputs(138));
    layer0_outputs(4480) <= not((inputs(85)) or (inputs(73)));
    layer0_outputs(4481) <= inputs(171);
    layer0_outputs(4482) <= not((inputs(168)) and (inputs(184)));
    layer0_outputs(4483) <= not(inputs(227)) or (inputs(240));
    layer0_outputs(4484) <= not(inputs(56)) or (inputs(231));
    layer0_outputs(4485) <= (inputs(94)) or (inputs(84));
    layer0_outputs(4486) <= (inputs(110)) xor (inputs(33));
    layer0_outputs(4487) <= not(inputs(76)) or (inputs(32));
    layer0_outputs(4488) <= not((inputs(122)) xor (inputs(160)));
    layer0_outputs(4489) <= not(inputs(113)) or (inputs(66));
    layer0_outputs(4490) <= (inputs(123)) and not (inputs(162));
    layer0_outputs(4491) <= (inputs(229)) and not (inputs(99));
    layer0_outputs(4492) <= (inputs(21)) xor (inputs(42));
    layer0_outputs(4493) <= not((inputs(94)) xor (inputs(6)));
    layer0_outputs(4494) <= (inputs(235)) xor (inputs(233));
    layer0_outputs(4495) <= inputs(159);
    layer0_outputs(4496) <= not(inputs(85));
    layer0_outputs(4497) <= (inputs(142)) and (inputs(7));
    layer0_outputs(4498) <= not((inputs(181)) xor (inputs(63)));
    layer0_outputs(4499) <= inputs(34);
    layer0_outputs(4500) <= (inputs(240)) xor (inputs(91));
    layer0_outputs(4501) <= not((inputs(60)) or (inputs(167)));
    layer0_outputs(4502) <= (inputs(26)) or (inputs(180));
    layer0_outputs(4503) <= (inputs(169)) and not (inputs(62));
    layer0_outputs(4504) <= (inputs(212)) or (inputs(140));
    layer0_outputs(4505) <= not((inputs(203)) or (inputs(205)));
    layer0_outputs(4506) <= not(inputs(114)) or (inputs(46));
    layer0_outputs(4507) <= not(inputs(96));
    layer0_outputs(4508) <= not(inputs(147));
    layer0_outputs(4509) <= inputs(47);
    layer0_outputs(4510) <= not((inputs(159)) and (inputs(193)));
    layer0_outputs(4511) <= inputs(34);
    layer0_outputs(4512) <= (inputs(82)) xor (inputs(60));
    layer0_outputs(4513) <= (inputs(239)) and not (inputs(141));
    layer0_outputs(4514) <= not(inputs(85)) or (inputs(34));
    layer0_outputs(4515) <= not((inputs(110)) or (inputs(221)));
    layer0_outputs(4516) <= not((inputs(75)) or (inputs(237)));
    layer0_outputs(4517) <= (inputs(212)) xor (inputs(132));
    layer0_outputs(4518) <= (inputs(45)) and (inputs(160));
    layer0_outputs(4519) <= not(inputs(237));
    layer0_outputs(4520) <= not((inputs(166)) xor (inputs(253)));
    layer0_outputs(4521) <= (inputs(108)) or (inputs(46));
    layer0_outputs(4522) <= not((inputs(7)) xor (inputs(114)));
    layer0_outputs(4523) <= not((inputs(58)) or (inputs(239)));
    layer0_outputs(4524) <= not((inputs(125)) and (inputs(10)));
    layer0_outputs(4525) <= (inputs(144)) or (inputs(164));
    layer0_outputs(4526) <= (inputs(185)) xor (inputs(169));
    layer0_outputs(4527) <= not(inputs(33)) or (inputs(30));
    layer0_outputs(4528) <= (inputs(250)) and (inputs(226));
    layer0_outputs(4529) <= not(inputs(57));
    layer0_outputs(4530) <= inputs(108);
    layer0_outputs(4531) <= not(inputs(6)) or (inputs(49));
    layer0_outputs(4532) <= not(inputs(228)) or (inputs(209));
    layer0_outputs(4533) <= not((inputs(148)) xor (inputs(151)));
    layer0_outputs(4534) <= not(inputs(200)) or (inputs(95));
    layer0_outputs(4535) <= inputs(230);
    layer0_outputs(4536) <= (inputs(136)) and not (inputs(205));
    layer0_outputs(4537) <= inputs(61);
    layer0_outputs(4538) <= not((inputs(195)) xor (inputs(83)));
    layer0_outputs(4539) <= not(inputs(138));
    layer0_outputs(4540) <= not(inputs(53)) or (inputs(240));
    layer0_outputs(4541) <= not((inputs(149)) or (inputs(106)));
    layer0_outputs(4542) <= not((inputs(94)) or (inputs(44)));
    layer0_outputs(4543) <= inputs(237);
    layer0_outputs(4544) <= '1';
    layer0_outputs(4545) <= not((inputs(54)) xor (inputs(64)));
    layer0_outputs(4546) <= not((inputs(116)) or (inputs(93)));
    layer0_outputs(4547) <= not((inputs(221)) or (inputs(182)));
    layer0_outputs(4548) <= (inputs(0)) xor (inputs(44));
    layer0_outputs(4549) <= not((inputs(178)) xor (inputs(72)));
    layer0_outputs(4550) <= not(inputs(139));
    layer0_outputs(4551) <= (inputs(54)) and not (inputs(145));
    layer0_outputs(4552) <= not(inputs(109)) or (inputs(227));
    layer0_outputs(4553) <= not(inputs(198));
    layer0_outputs(4554) <= (inputs(211)) and not (inputs(123));
    layer0_outputs(4555) <= (inputs(9)) and (inputs(245));
    layer0_outputs(4556) <= not(inputs(137));
    layer0_outputs(4557) <= inputs(126);
    layer0_outputs(4558) <= (inputs(58)) xor (inputs(56));
    layer0_outputs(4559) <= '0';
    layer0_outputs(4560) <= not(inputs(88)) or (inputs(26));
    layer0_outputs(4561) <= not((inputs(232)) or (inputs(196)));
    layer0_outputs(4562) <= not(inputs(22)) or (inputs(92));
    layer0_outputs(4563) <= not(inputs(102)) or (inputs(20));
    layer0_outputs(4564) <= not(inputs(150));
    layer0_outputs(4565) <= not((inputs(17)) xor (inputs(166)));
    layer0_outputs(4566) <= not((inputs(19)) and (inputs(19)));
    layer0_outputs(4567) <= (inputs(211)) xor (inputs(112));
    layer0_outputs(4568) <= (inputs(161)) xor (inputs(83));
    layer0_outputs(4569) <= not(inputs(97));
    layer0_outputs(4570) <= inputs(36);
    layer0_outputs(4571) <= not((inputs(127)) or (inputs(185)));
    layer0_outputs(4572) <= (inputs(4)) and (inputs(28));
    layer0_outputs(4573) <= (inputs(233)) xor (inputs(219));
    layer0_outputs(4574) <= (inputs(197)) and not (inputs(64));
    layer0_outputs(4575) <= inputs(168);
    layer0_outputs(4576) <= not(inputs(163));
    layer0_outputs(4577) <= inputs(157);
    layer0_outputs(4578) <= not(inputs(73)) or (inputs(196));
    layer0_outputs(4579) <= not(inputs(71));
    layer0_outputs(4580) <= (inputs(209)) and (inputs(2));
    layer0_outputs(4581) <= (inputs(126)) and not (inputs(33));
    layer0_outputs(4582) <= not((inputs(222)) or (inputs(131)));
    layer0_outputs(4583) <= not((inputs(36)) xor (inputs(250)));
    layer0_outputs(4584) <= '1';
    layer0_outputs(4585) <= not(inputs(165));
    layer0_outputs(4586) <= (inputs(18)) and not (inputs(64));
    layer0_outputs(4587) <= '0';
    layer0_outputs(4588) <= not(inputs(103)) or (inputs(255));
    layer0_outputs(4589) <= (inputs(247)) and not (inputs(80));
    layer0_outputs(4590) <= not((inputs(243)) and (inputs(243)));
    layer0_outputs(4591) <= not((inputs(89)) and (inputs(252)));
    layer0_outputs(4592) <= not(inputs(73)) or (inputs(77));
    layer0_outputs(4593) <= inputs(176);
    layer0_outputs(4594) <= (inputs(44)) xor (inputs(1));
    layer0_outputs(4595) <= (inputs(195)) xor (inputs(69));
    layer0_outputs(4596) <= (inputs(191)) and not (inputs(158));
    layer0_outputs(4597) <= inputs(88);
    layer0_outputs(4598) <= not((inputs(12)) and (inputs(6)));
    layer0_outputs(4599) <= not((inputs(145)) xor (inputs(137)));
    layer0_outputs(4600) <= not(inputs(138));
    layer0_outputs(4601) <= (inputs(53)) xor (inputs(252));
    layer0_outputs(4602) <= not(inputs(47));
    layer0_outputs(4603) <= not((inputs(158)) or (inputs(172)));
    layer0_outputs(4604) <= not(inputs(67));
    layer0_outputs(4605) <= (inputs(80)) and not (inputs(0));
    layer0_outputs(4606) <= (inputs(100)) and not (inputs(172));
    layer0_outputs(4607) <= (inputs(107)) and not (inputs(241));
    layer0_outputs(4608) <= not(inputs(203)) or (inputs(21));
    layer0_outputs(4609) <= not(inputs(100));
    layer0_outputs(4610) <= not((inputs(145)) xor (inputs(53)));
    layer0_outputs(4611) <= (inputs(54)) or (inputs(241));
    layer0_outputs(4612) <= (inputs(156)) or (inputs(155));
    layer0_outputs(4613) <= not((inputs(140)) or (inputs(61)));
    layer0_outputs(4614) <= not((inputs(157)) or (inputs(237)));
    layer0_outputs(4615) <= (inputs(239)) xor (inputs(172));
    layer0_outputs(4616) <= not(inputs(188)) or (inputs(237));
    layer0_outputs(4617) <= not((inputs(179)) or (inputs(194)));
    layer0_outputs(4618) <= not(inputs(197));
    layer0_outputs(4619) <= not((inputs(162)) xor (inputs(221)));
    layer0_outputs(4620) <= '0';
    layer0_outputs(4621) <= (inputs(87)) and not (inputs(54));
    layer0_outputs(4622) <= inputs(134);
    layer0_outputs(4623) <= (inputs(101)) or (inputs(233));
    layer0_outputs(4624) <= (inputs(214)) or (inputs(11));
    layer0_outputs(4625) <= not((inputs(121)) xor (inputs(1)));
    layer0_outputs(4626) <= not(inputs(179)) or (inputs(191));
    layer0_outputs(4627) <= not((inputs(90)) xor (inputs(11)));
    layer0_outputs(4628) <= not(inputs(136)) or (inputs(86));
    layer0_outputs(4629) <= not((inputs(138)) or (inputs(161)));
    layer0_outputs(4630) <= (inputs(55)) and (inputs(39));
    layer0_outputs(4631) <= not((inputs(254)) or (inputs(244)));
    layer0_outputs(4632) <= (inputs(145)) xor (inputs(185));
    layer0_outputs(4633) <= (inputs(186)) xor (inputs(95));
    layer0_outputs(4634) <= not(inputs(105));
    layer0_outputs(4635) <= not(inputs(154));
    layer0_outputs(4636) <= (inputs(180)) xor (inputs(111));
    layer0_outputs(4637) <= not(inputs(58));
    layer0_outputs(4638) <= (inputs(105)) and not (inputs(30));
    layer0_outputs(4639) <= not((inputs(154)) xor (inputs(80)));
    layer0_outputs(4640) <= not(inputs(232));
    layer0_outputs(4641) <= not((inputs(37)) xor (inputs(63)));
    layer0_outputs(4642) <= (inputs(138)) xor (inputs(46));
    layer0_outputs(4643) <= (inputs(87)) and not (inputs(130));
    layer0_outputs(4644) <= not(inputs(232)) or (inputs(162));
    layer0_outputs(4645) <= not(inputs(198)) or (inputs(218));
    layer0_outputs(4646) <= '0';
    layer0_outputs(4647) <= not(inputs(61)) or (inputs(47));
    layer0_outputs(4648) <= (inputs(134)) and (inputs(241));
    layer0_outputs(4649) <= (inputs(142)) or (inputs(97));
    layer0_outputs(4650) <= not((inputs(206)) or (inputs(190)));
    layer0_outputs(4651) <= (inputs(35)) and not (inputs(125));
    layer0_outputs(4652) <= not((inputs(116)) and (inputs(187)));
    layer0_outputs(4653) <= inputs(196);
    layer0_outputs(4654) <= inputs(117);
    layer0_outputs(4655) <= not(inputs(124));
    layer0_outputs(4656) <= not(inputs(110)) or (inputs(34));
    layer0_outputs(4657) <= (inputs(34)) or (inputs(66));
    layer0_outputs(4658) <= (inputs(204)) or (inputs(137));
    layer0_outputs(4659) <= not(inputs(204)) or (inputs(10));
    layer0_outputs(4660) <= not(inputs(78));
    layer0_outputs(4661) <= not((inputs(118)) xor (inputs(28)));
    layer0_outputs(4662) <= inputs(86);
    layer0_outputs(4663) <= not(inputs(237)) or (inputs(113));
    layer0_outputs(4664) <= (inputs(140)) and not (inputs(207));
    layer0_outputs(4665) <= not((inputs(88)) or (inputs(240)));
    layer0_outputs(4666) <= not(inputs(159)) or (inputs(209));
    layer0_outputs(4667) <= not(inputs(31));
    layer0_outputs(4668) <= not(inputs(254)) or (inputs(29));
    layer0_outputs(4669) <= not((inputs(176)) xor (inputs(12)));
    layer0_outputs(4670) <= (inputs(37)) or (inputs(230));
    layer0_outputs(4671) <= not(inputs(197)) or (inputs(239));
    layer0_outputs(4672) <= not(inputs(113)) or (inputs(48));
    layer0_outputs(4673) <= not(inputs(100));
    layer0_outputs(4674) <= not(inputs(214));
    layer0_outputs(4675) <= not(inputs(195));
    layer0_outputs(4676) <= (inputs(254)) or (inputs(52));
    layer0_outputs(4677) <= inputs(122);
    layer0_outputs(4678) <= not((inputs(10)) xor (inputs(131)));
    layer0_outputs(4679) <= inputs(169);
    layer0_outputs(4680) <= (inputs(53)) xor (inputs(92));
    layer0_outputs(4681) <= not((inputs(152)) or (inputs(121)));
    layer0_outputs(4682) <= not((inputs(101)) xor (inputs(221)));
    layer0_outputs(4683) <= (inputs(167)) and not (inputs(230));
    layer0_outputs(4684) <= not((inputs(222)) xor (inputs(153)));
    layer0_outputs(4685) <= not((inputs(45)) xor (inputs(81)));
    layer0_outputs(4686) <= (inputs(0)) xor (inputs(132));
    layer0_outputs(4687) <= not(inputs(22)) or (inputs(22));
    layer0_outputs(4688) <= (inputs(216)) and not (inputs(89));
    layer0_outputs(4689) <= not((inputs(28)) xor (inputs(50)));
    layer0_outputs(4690) <= not(inputs(129)) or (inputs(173));
    layer0_outputs(4691) <= not((inputs(192)) or (inputs(155)));
    layer0_outputs(4692) <= '1';
    layer0_outputs(4693) <= not(inputs(247));
    layer0_outputs(4694) <= (inputs(113)) and not (inputs(130));
    layer0_outputs(4695) <= (inputs(126)) and (inputs(65));
    layer0_outputs(4696) <= inputs(240);
    layer0_outputs(4697) <= inputs(185);
    layer0_outputs(4698) <= inputs(231);
    layer0_outputs(4699) <= not((inputs(97)) or (inputs(160)));
    layer0_outputs(4700) <= (inputs(138)) or (inputs(207));
    layer0_outputs(4701) <= not(inputs(146));
    layer0_outputs(4702) <= (inputs(159)) and not (inputs(62));
    layer0_outputs(4703) <= (inputs(85)) xor (inputs(20));
    layer0_outputs(4704) <= not(inputs(167)) or (inputs(230));
    layer0_outputs(4705) <= (inputs(190)) and not (inputs(169));
    layer0_outputs(4706) <= (inputs(250)) xor (inputs(126));
    layer0_outputs(4707) <= (inputs(117)) and not (inputs(195));
    layer0_outputs(4708) <= (inputs(215)) or (inputs(39));
    layer0_outputs(4709) <= not(inputs(185)) or (inputs(152));
    layer0_outputs(4710) <= (inputs(230)) and not (inputs(197));
    layer0_outputs(4711) <= '0';
    layer0_outputs(4712) <= (inputs(134)) and not (inputs(231));
    layer0_outputs(4713) <= inputs(79);
    layer0_outputs(4714) <= not((inputs(154)) xor (inputs(116)));
    layer0_outputs(4715) <= not((inputs(27)) or (inputs(239)));
    layer0_outputs(4716) <= (inputs(71)) and (inputs(41));
    layer0_outputs(4717) <= (inputs(235)) or (inputs(118));
    layer0_outputs(4718) <= (inputs(99)) or (inputs(251));
    layer0_outputs(4719) <= (inputs(248)) or (inputs(117));
    layer0_outputs(4720) <= inputs(236);
    layer0_outputs(4721) <= (inputs(126)) and not (inputs(47));
    layer0_outputs(4722) <= (inputs(131)) or (inputs(181));
    layer0_outputs(4723) <= not((inputs(38)) or (inputs(121)));
    layer0_outputs(4724) <= not(inputs(234)) or (inputs(158));
    layer0_outputs(4725) <= (inputs(72)) xor (inputs(198));
    layer0_outputs(4726) <= not((inputs(108)) and (inputs(3)));
    layer0_outputs(4727) <= inputs(93);
    layer0_outputs(4728) <= not(inputs(238));
    layer0_outputs(4729) <= not(inputs(230));
    layer0_outputs(4730) <= '1';
    layer0_outputs(4731) <= not((inputs(59)) or (inputs(123)));
    layer0_outputs(4732) <= inputs(203);
    layer0_outputs(4733) <= not(inputs(234));
    layer0_outputs(4734) <= (inputs(197)) or (inputs(170));
    layer0_outputs(4735) <= (inputs(73)) and not (inputs(84));
    layer0_outputs(4736) <= inputs(179);
    layer0_outputs(4737) <= not(inputs(234));
    layer0_outputs(4738) <= (inputs(11)) and not (inputs(66));
    layer0_outputs(4739) <= not((inputs(200)) xor (inputs(23)));
    layer0_outputs(4740) <= not(inputs(41));
    layer0_outputs(4741) <= not((inputs(119)) xor (inputs(254)));
    layer0_outputs(4742) <= not((inputs(222)) and (inputs(237)));
    layer0_outputs(4743) <= (inputs(85)) xor (inputs(103));
    layer0_outputs(4744) <= not(inputs(181));
    layer0_outputs(4745) <= not(inputs(138)) or (inputs(40));
    layer0_outputs(4746) <= not((inputs(2)) xor (inputs(177)));
    layer0_outputs(4747) <= '0';
    layer0_outputs(4748) <= (inputs(132)) and not (inputs(194));
    layer0_outputs(4749) <= not((inputs(248)) xor (inputs(51)));
    layer0_outputs(4750) <= not(inputs(92));
    layer0_outputs(4751) <= not(inputs(171));
    layer0_outputs(4752) <= not(inputs(195)) or (inputs(147));
    layer0_outputs(4753) <= not(inputs(82)) or (inputs(24));
    layer0_outputs(4754) <= (inputs(94)) xor (inputs(188));
    layer0_outputs(4755) <= not(inputs(137));
    layer0_outputs(4756) <= not(inputs(225));
    layer0_outputs(4757) <= not(inputs(92)) or (inputs(173));
    layer0_outputs(4758) <= not(inputs(179)) or (inputs(229));
    layer0_outputs(4759) <= not((inputs(79)) and (inputs(112)));
    layer0_outputs(4760) <= not(inputs(156));
    layer0_outputs(4761) <= inputs(185);
    layer0_outputs(4762) <= not(inputs(156));
    layer0_outputs(4763) <= (inputs(111)) and (inputs(30));
    layer0_outputs(4764) <= not((inputs(176)) xor (inputs(212)));
    layer0_outputs(4765) <= not(inputs(42));
    layer0_outputs(4766) <= (inputs(102)) or (inputs(180));
    layer0_outputs(4767) <= (inputs(184)) and not (inputs(83));
    layer0_outputs(4768) <= not((inputs(254)) and (inputs(34)));
    layer0_outputs(4769) <= '1';
    layer0_outputs(4770) <= not(inputs(200));
    layer0_outputs(4771) <= not(inputs(55));
    layer0_outputs(4772) <= inputs(133);
    layer0_outputs(4773) <= (inputs(185)) or (inputs(147));
    layer0_outputs(4774) <= not((inputs(132)) or (inputs(160)));
    layer0_outputs(4775) <= not((inputs(106)) and (inputs(16)));
    layer0_outputs(4776) <= not(inputs(50));
    layer0_outputs(4777) <= (inputs(186)) or (inputs(26));
    layer0_outputs(4778) <= not(inputs(251)) or (inputs(128));
    layer0_outputs(4779) <= (inputs(204)) xor (inputs(142));
    layer0_outputs(4780) <= (inputs(43)) or (inputs(61));
    layer0_outputs(4781) <= not((inputs(139)) xor (inputs(53)));
    layer0_outputs(4782) <= inputs(167);
    layer0_outputs(4783) <= not((inputs(128)) xor (inputs(234)));
    layer0_outputs(4784) <= not((inputs(165)) xor (inputs(50)));
    layer0_outputs(4785) <= not((inputs(10)) xor (inputs(58)));
    layer0_outputs(4786) <= not((inputs(18)) or (inputs(185)));
    layer0_outputs(4787) <= not(inputs(110));
    layer0_outputs(4788) <= (inputs(179)) or (inputs(38));
    layer0_outputs(4789) <= not(inputs(42));
    layer0_outputs(4790) <= not(inputs(59)) or (inputs(27));
    layer0_outputs(4791) <= inputs(119);
    layer0_outputs(4792) <= (inputs(162)) or (inputs(75));
    layer0_outputs(4793) <= (inputs(229)) or (inputs(248));
    layer0_outputs(4794) <= '0';
    layer0_outputs(4795) <= not((inputs(61)) or (inputs(27)));
    layer0_outputs(4796) <= (inputs(133)) and not (inputs(249));
    layer0_outputs(4797) <= not((inputs(56)) or (inputs(199)));
    layer0_outputs(4798) <= (inputs(65)) and not (inputs(161));
    layer0_outputs(4799) <= not((inputs(151)) or (inputs(46)));
    layer0_outputs(4800) <= (inputs(191)) or (inputs(220));
    layer0_outputs(4801) <= (inputs(87)) and not (inputs(227));
    layer0_outputs(4802) <= not((inputs(254)) xor (inputs(33)));
    layer0_outputs(4803) <= inputs(213);
    layer0_outputs(4804) <= (inputs(116)) xor (inputs(62));
    layer0_outputs(4805) <= not(inputs(141));
    layer0_outputs(4806) <= not(inputs(15));
    layer0_outputs(4807) <= not(inputs(122));
    layer0_outputs(4808) <= inputs(213);
    layer0_outputs(4809) <= not((inputs(166)) and (inputs(225)));
    layer0_outputs(4810) <= not(inputs(128));
    layer0_outputs(4811) <= not(inputs(74)) or (inputs(159));
    layer0_outputs(4812) <= not(inputs(123)) or (inputs(66));
    layer0_outputs(4813) <= inputs(40);
    layer0_outputs(4814) <= (inputs(106)) and not (inputs(78));
    layer0_outputs(4815) <= not(inputs(167));
    layer0_outputs(4816) <= inputs(108);
    layer0_outputs(4817) <= inputs(147);
    layer0_outputs(4818) <= not(inputs(134));
    layer0_outputs(4819) <= (inputs(237)) and not (inputs(190));
    layer0_outputs(4820) <= (inputs(50)) and not (inputs(1));
    layer0_outputs(4821) <= not(inputs(40));
    layer0_outputs(4822) <= (inputs(41)) and not (inputs(208));
    layer0_outputs(4823) <= (inputs(82)) xor (inputs(23));
    layer0_outputs(4824) <= inputs(123);
    layer0_outputs(4825) <= not((inputs(205)) xor (inputs(214)));
    layer0_outputs(4826) <= (inputs(69)) xor (inputs(212));
    layer0_outputs(4827) <= (inputs(23)) xor (inputs(227));
    layer0_outputs(4828) <= (inputs(76)) xor (inputs(183));
    layer0_outputs(4829) <= (inputs(152)) xor (inputs(225));
    layer0_outputs(4830) <= (inputs(237)) or (inputs(110));
    layer0_outputs(4831) <= (inputs(165)) and not (inputs(42));
    layer0_outputs(4832) <= (inputs(56)) or (inputs(75));
    layer0_outputs(4833) <= (inputs(114)) and not (inputs(28));
    layer0_outputs(4834) <= inputs(176);
    layer0_outputs(4835) <= not((inputs(170)) xor (inputs(225)));
    layer0_outputs(4836) <= '1';
    layer0_outputs(4837) <= (inputs(49)) and (inputs(145));
    layer0_outputs(4838) <= not((inputs(128)) xor (inputs(74)));
    layer0_outputs(4839) <= (inputs(58)) xor (inputs(60));
    layer0_outputs(4840) <= not((inputs(220)) xor (inputs(243)));
    layer0_outputs(4841) <= not(inputs(4));
    layer0_outputs(4842) <= '1';
    layer0_outputs(4843) <= not(inputs(101));
    layer0_outputs(4844) <= not(inputs(55)) or (inputs(127));
    layer0_outputs(4845) <= (inputs(86)) and not (inputs(47));
    layer0_outputs(4846) <= (inputs(221)) and not (inputs(29));
    layer0_outputs(4847) <= not(inputs(186));
    layer0_outputs(4848) <= (inputs(149)) or (inputs(46));
    layer0_outputs(4849) <= not(inputs(92)) or (inputs(224));
    layer0_outputs(4850) <= (inputs(95)) or (inputs(100));
    layer0_outputs(4851) <= (inputs(12)) and not (inputs(206));
    layer0_outputs(4852) <= (inputs(142)) xor (inputs(44));
    layer0_outputs(4853) <= not(inputs(136)) or (inputs(43));
    layer0_outputs(4854) <= not(inputs(176));
    layer0_outputs(4855) <= inputs(57);
    layer0_outputs(4856) <= (inputs(188)) or (inputs(163));
    layer0_outputs(4857) <= (inputs(55)) xor (inputs(7));
    layer0_outputs(4858) <= (inputs(139)) and not (inputs(126));
    layer0_outputs(4859) <= not((inputs(35)) and (inputs(157)));
    layer0_outputs(4860) <= (inputs(42)) and (inputs(247));
    layer0_outputs(4861) <= not(inputs(199));
    layer0_outputs(4862) <= not(inputs(87));
    layer0_outputs(4863) <= (inputs(241)) and not (inputs(4));
    layer0_outputs(4864) <= not(inputs(228)) or (inputs(24));
    layer0_outputs(4865) <= (inputs(20)) or (inputs(184));
    layer0_outputs(4866) <= not((inputs(160)) or (inputs(201)));
    layer0_outputs(4867) <= not(inputs(106));
    layer0_outputs(4868) <= not(inputs(59));
    layer0_outputs(4869) <= not(inputs(47));
    layer0_outputs(4870) <= '0';
    layer0_outputs(4871) <= (inputs(150)) and not (inputs(215));
    layer0_outputs(4872) <= not((inputs(3)) and (inputs(113)));
    layer0_outputs(4873) <= not((inputs(86)) or (inputs(169)));
    layer0_outputs(4874) <= (inputs(65)) xor (inputs(152));
    layer0_outputs(4875) <= not(inputs(184)) or (inputs(70));
    layer0_outputs(4876) <= not(inputs(251));
    layer0_outputs(4877) <= inputs(186);
    layer0_outputs(4878) <= (inputs(178)) or (inputs(163));
    layer0_outputs(4879) <= not(inputs(249)) or (inputs(21));
    layer0_outputs(4880) <= not(inputs(133)) or (inputs(22));
    layer0_outputs(4881) <= not(inputs(133));
    layer0_outputs(4882) <= not(inputs(72));
    layer0_outputs(4883) <= inputs(231);
    layer0_outputs(4884) <= '0';
    layer0_outputs(4885) <= not((inputs(150)) and (inputs(172)));
    layer0_outputs(4886) <= inputs(74);
    layer0_outputs(4887) <= not((inputs(77)) or (inputs(241)));
    layer0_outputs(4888) <= (inputs(2)) or (inputs(10));
    layer0_outputs(4889) <= not(inputs(160)) or (inputs(3));
    layer0_outputs(4890) <= (inputs(64)) xor (inputs(229));
    layer0_outputs(4891) <= not((inputs(182)) or (inputs(26)));
    layer0_outputs(4892) <= not(inputs(69));
    layer0_outputs(4893) <= not(inputs(134)) or (inputs(237));
    layer0_outputs(4894) <= not(inputs(251)) or (inputs(219));
    layer0_outputs(4895) <= not(inputs(105)) or (inputs(88));
    layer0_outputs(4896) <= inputs(6);
    layer0_outputs(4897) <= not((inputs(242)) or (inputs(243)));
    layer0_outputs(4898) <= not((inputs(251)) or (inputs(187)));
    layer0_outputs(4899) <= '1';
    layer0_outputs(4900) <= inputs(239);
    layer0_outputs(4901) <= (inputs(150)) and not (inputs(78));
    layer0_outputs(4902) <= inputs(219);
    layer0_outputs(4903) <= (inputs(138)) and not (inputs(162));
    layer0_outputs(4904) <= not(inputs(181));
    layer0_outputs(4905) <= not((inputs(42)) xor (inputs(40)));
    layer0_outputs(4906) <= (inputs(186)) and not (inputs(17));
    layer0_outputs(4907) <= (inputs(200)) or (inputs(26));
    layer0_outputs(4908) <= not((inputs(86)) xor (inputs(252)));
    layer0_outputs(4909) <= not(inputs(34));
    layer0_outputs(4910) <= inputs(138);
    layer0_outputs(4911) <= not((inputs(192)) or (inputs(126)));
    layer0_outputs(4912) <= (inputs(111)) and not (inputs(236));
    layer0_outputs(4913) <= not((inputs(171)) xor (inputs(93)));
    layer0_outputs(4914) <= (inputs(3)) and not (inputs(199));
    layer0_outputs(4915) <= not((inputs(67)) or (inputs(223)));
    layer0_outputs(4916) <= not(inputs(64)) or (inputs(6));
    layer0_outputs(4917) <= (inputs(110)) or (inputs(136));
    layer0_outputs(4918) <= not(inputs(180)) or (inputs(4));
    layer0_outputs(4919) <= (inputs(51)) xor (inputs(122));
    layer0_outputs(4920) <= (inputs(106)) or (inputs(50));
    layer0_outputs(4921) <= not(inputs(255));
    layer0_outputs(4922) <= (inputs(73)) and not (inputs(98));
    layer0_outputs(4923) <= (inputs(242)) and not (inputs(20));
    layer0_outputs(4924) <= (inputs(94)) and not (inputs(141));
    layer0_outputs(4925) <= not((inputs(211)) xor (inputs(188)));
    layer0_outputs(4926) <= not((inputs(179)) or (inputs(178)));
    layer0_outputs(4927) <= (inputs(132)) and not (inputs(81));
    layer0_outputs(4928) <= not((inputs(202)) or (inputs(229)));
    layer0_outputs(4929) <= (inputs(100)) and not (inputs(11));
    layer0_outputs(4930) <= inputs(119);
    layer0_outputs(4931) <= (inputs(58)) and not (inputs(30));
    layer0_outputs(4932) <= not(inputs(219)) or (inputs(8));
    layer0_outputs(4933) <= not(inputs(54)) or (inputs(220));
    layer0_outputs(4934) <= not((inputs(129)) or (inputs(83)));
    layer0_outputs(4935) <= not(inputs(133)) or (inputs(64));
    layer0_outputs(4936) <= not(inputs(254));
    layer0_outputs(4937) <= (inputs(193)) or (inputs(119));
    layer0_outputs(4938) <= inputs(125);
    layer0_outputs(4939) <= (inputs(80)) and (inputs(81));
    layer0_outputs(4940) <= not((inputs(248)) xor (inputs(163)));
    layer0_outputs(4941) <= (inputs(12)) and not (inputs(248));
    layer0_outputs(4942) <= (inputs(177)) and not (inputs(249));
    layer0_outputs(4943) <= (inputs(196)) and not (inputs(168));
    layer0_outputs(4944) <= not(inputs(55));
    layer0_outputs(4945) <= not(inputs(15));
    layer0_outputs(4946) <= not(inputs(40));
    layer0_outputs(4947) <= not(inputs(37)) or (inputs(34));
    layer0_outputs(4948) <= not((inputs(215)) or (inputs(47)));
    layer0_outputs(4949) <= inputs(117);
    layer0_outputs(4950) <= not((inputs(147)) xor (inputs(118)));
    layer0_outputs(4951) <= (inputs(20)) and not (inputs(142));
    layer0_outputs(4952) <= not(inputs(32)) or (inputs(96));
    layer0_outputs(4953) <= inputs(152);
    layer0_outputs(4954) <= not(inputs(154));
    layer0_outputs(4955) <= not((inputs(132)) and (inputs(138)));
    layer0_outputs(4956) <= not((inputs(55)) xor (inputs(190)));
    layer0_outputs(4957) <= not((inputs(167)) or (inputs(67)));
    layer0_outputs(4958) <= (inputs(127)) or (inputs(38));
    layer0_outputs(4959) <= inputs(36);
    layer0_outputs(4960) <= not((inputs(121)) and (inputs(105)));
    layer0_outputs(4961) <= (inputs(103)) and (inputs(136));
    layer0_outputs(4962) <= (inputs(203)) or (inputs(165));
    layer0_outputs(4963) <= not((inputs(87)) xor (inputs(253)));
    layer0_outputs(4964) <= (inputs(47)) and not (inputs(212));
    layer0_outputs(4965) <= not(inputs(121)) or (inputs(22));
    layer0_outputs(4966) <= not((inputs(90)) or (inputs(216)));
    layer0_outputs(4967) <= not((inputs(251)) xor (inputs(24)));
    layer0_outputs(4968) <= not(inputs(199));
    layer0_outputs(4969) <= (inputs(84)) xor (inputs(253));
    layer0_outputs(4970) <= not(inputs(75)) or (inputs(243));
    layer0_outputs(4971) <= not(inputs(136)) or (inputs(62));
    layer0_outputs(4972) <= inputs(92);
    layer0_outputs(4973) <= (inputs(157)) or (inputs(39));
    layer0_outputs(4974) <= not((inputs(242)) or (inputs(57)));
    layer0_outputs(4975) <= not((inputs(249)) or (inputs(77)));
    layer0_outputs(4976) <= inputs(89);
    layer0_outputs(4977) <= not(inputs(79));
    layer0_outputs(4978) <= inputs(213);
    layer0_outputs(4979) <= '0';
    layer0_outputs(4980) <= inputs(204);
    layer0_outputs(4981) <= not((inputs(112)) or (inputs(210)));
    layer0_outputs(4982) <= (inputs(40)) and not (inputs(190));
    layer0_outputs(4983) <= inputs(183);
    layer0_outputs(4984) <= not(inputs(8)) or (inputs(78));
    layer0_outputs(4985) <= not((inputs(153)) or (inputs(189)));
    layer0_outputs(4986) <= inputs(214);
    layer0_outputs(4987) <= (inputs(218)) and not (inputs(2));
    layer0_outputs(4988) <= inputs(163);
    layer0_outputs(4989) <= not((inputs(243)) and (inputs(194)));
    layer0_outputs(4990) <= (inputs(183)) xor (inputs(120));
    layer0_outputs(4991) <= not(inputs(101)) or (inputs(255));
    layer0_outputs(4992) <= not(inputs(149)) or (inputs(173));
    layer0_outputs(4993) <= inputs(132);
    layer0_outputs(4994) <= not(inputs(147));
    layer0_outputs(4995) <= not(inputs(97));
    layer0_outputs(4996) <= not(inputs(41));
    layer0_outputs(4997) <= (inputs(213)) or (inputs(63));
    layer0_outputs(4998) <= (inputs(151)) xor (inputs(211));
    layer0_outputs(4999) <= '0';
    layer0_outputs(5000) <= (inputs(168)) and not (inputs(95));
    layer0_outputs(5001) <= (inputs(55)) or (inputs(201));
    layer0_outputs(5002) <= (inputs(104)) and not (inputs(179));
    layer0_outputs(5003) <= (inputs(211)) or (inputs(228));
    layer0_outputs(5004) <= not(inputs(99));
    layer0_outputs(5005) <= not((inputs(148)) or (inputs(77)));
    layer0_outputs(5006) <= (inputs(168)) or (inputs(82));
    layer0_outputs(5007) <= not((inputs(98)) or (inputs(42)));
    layer0_outputs(5008) <= (inputs(82)) and not (inputs(28));
    layer0_outputs(5009) <= not(inputs(201));
    layer0_outputs(5010) <= inputs(62);
    layer0_outputs(5011) <= (inputs(34)) xor (inputs(9));
    layer0_outputs(5012) <= not(inputs(120));
    layer0_outputs(5013) <= inputs(41);
    layer0_outputs(5014) <= (inputs(36)) or (inputs(9));
    layer0_outputs(5015) <= not((inputs(149)) xor (inputs(222)));
    layer0_outputs(5016) <= (inputs(249)) or (inputs(117));
    layer0_outputs(5017) <= not((inputs(223)) or (inputs(112)));
    layer0_outputs(5018) <= not((inputs(84)) xor (inputs(166)));
    layer0_outputs(5019) <= '1';
    layer0_outputs(5020) <= (inputs(179)) and (inputs(239));
    layer0_outputs(5021) <= not((inputs(39)) xor (inputs(122)));
    layer0_outputs(5022) <= inputs(150);
    layer0_outputs(5023) <= not((inputs(204)) xor (inputs(73)));
    layer0_outputs(5024) <= inputs(232);
    layer0_outputs(5025) <= (inputs(254)) and (inputs(20));
    layer0_outputs(5026) <= not(inputs(125)) or (inputs(207));
    layer0_outputs(5027) <= not((inputs(68)) xor (inputs(172)));
    layer0_outputs(5028) <= (inputs(101)) and not (inputs(195));
    layer0_outputs(5029) <= (inputs(18)) xor (inputs(117));
    layer0_outputs(5030) <= (inputs(18)) xor (inputs(102));
    layer0_outputs(5031) <= not(inputs(174)) or (inputs(17));
    layer0_outputs(5032) <= inputs(124);
    layer0_outputs(5033) <= not(inputs(114)) or (inputs(207));
    layer0_outputs(5034) <= '1';
    layer0_outputs(5035) <= (inputs(104)) or (inputs(189));
    layer0_outputs(5036) <= (inputs(139)) xor (inputs(220));
    layer0_outputs(5037) <= inputs(77);
    layer0_outputs(5038) <= not(inputs(83)) or (inputs(69));
    layer0_outputs(5039) <= (inputs(188)) xor (inputs(151));
    layer0_outputs(5040) <= not(inputs(76));
    layer0_outputs(5041) <= (inputs(102)) and not (inputs(26));
    layer0_outputs(5042) <= (inputs(159)) xor (inputs(179));
    layer0_outputs(5043) <= (inputs(138)) and not (inputs(202));
    layer0_outputs(5044) <= inputs(229);
    layer0_outputs(5045) <= not(inputs(86)) or (inputs(182));
    layer0_outputs(5046) <= not((inputs(67)) or (inputs(249)));
    layer0_outputs(5047) <= not(inputs(27));
    layer0_outputs(5048) <= inputs(138);
    layer0_outputs(5049) <= (inputs(208)) or (inputs(215));
    layer0_outputs(5050) <= inputs(119);
    layer0_outputs(5051) <= (inputs(28)) and not (inputs(185));
    layer0_outputs(5052) <= inputs(134);
    layer0_outputs(5053) <= not((inputs(20)) or (inputs(183)));
    layer0_outputs(5054) <= not(inputs(166));
    layer0_outputs(5055) <= not(inputs(109));
    layer0_outputs(5056) <= inputs(42);
    layer0_outputs(5057) <= not((inputs(110)) or (inputs(161)));
    layer0_outputs(5058) <= (inputs(175)) xor (inputs(42));
    layer0_outputs(5059) <= not((inputs(254)) or (inputs(187)));
    layer0_outputs(5060) <= '0';
    layer0_outputs(5061) <= (inputs(5)) xor (inputs(61));
    layer0_outputs(5062) <= not(inputs(139));
    layer0_outputs(5063) <= not(inputs(153));
    layer0_outputs(5064) <= (inputs(136)) xor (inputs(49));
    layer0_outputs(5065) <= not((inputs(8)) or (inputs(103)));
    layer0_outputs(5066) <= (inputs(14)) or (inputs(108));
    layer0_outputs(5067) <= not(inputs(70));
    layer0_outputs(5068) <= not(inputs(192));
    layer0_outputs(5069) <= (inputs(41)) or (inputs(5));
    layer0_outputs(5070) <= not(inputs(164)) or (inputs(110));
    layer0_outputs(5071) <= not((inputs(128)) xor (inputs(54)));
    layer0_outputs(5072) <= not((inputs(218)) or (inputs(113)));
    layer0_outputs(5073) <= not(inputs(179)) or (inputs(219));
    layer0_outputs(5074) <= not((inputs(223)) or (inputs(50)));
    layer0_outputs(5075) <= not(inputs(22)) or (inputs(236));
    layer0_outputs(5076) <= not((inputs(119)) xor (inputs(64)));
    layer0_outputs(5077) <= (inputs(213)) and (inputs(239));
    layer0_outputs(5078) <= not(inputs(6)) or (inputs(16));
    layer0_outputs(5079) <= inputs(28);
    layer0_outputs(5080) <= not(inputs(220));
    layer0_outputs(5081) <= not((inputs(60)) or (inputs(32)));
    layer0_outputs(5082) <= inputs(77);
    layer0_outputs(5083) <= not((inputs(12)) xor (inputs(201)));
    layer0_outputs(5084) <= (inputs(238)) xor (inputs(152));
    layer0_outputs(5085) <= not(inputs(232)) or (inputs(75));
    layer0_outputs(5086) <= inputs(9);
    layer0_outputs(5087) <= not(inputs(148));
    layer0_outputs(5088) <= (inputs(249)) or (inputs(231));
    layer0_outputs(5089) <= (inputs(189)) or (inputs(131));
    layer0_outputs(5090) <= (inputs(212)) or (inputs(211));
    layer0_outputs(5091) <= not(inputs(179)) or (inputs(206));
    layer0_outputs(5092) <= not(inputs(57));
    layer0_outputs(5093) <= not((inputs(118)) or (inputs(20)));
    layer0_outputs(5094) <= not((inputs(79)) or (inputs(211)));
    layer0_outputs(5095) <= inputs(204);
    layer0_outputs(5096) <= (inputs(218)) xor (inputs(148));
    layer0_outputs(5097) <= not(inputs(42)) or (inputs(209));
    layer0_outputs(5098) <= not(inputs(162)) or (inputs(252));
    layer0_outputs(5099) <= not((inputs(249)) and (inputs(221)));
    layer0_outputs(5100) <= inputs(192);
    layer0_outputs(5101) <= not((inputs(223)) or (inputs(182)));
    layer0_outputs(5102) <= inputs(90);
    layer0_outputs(5103) <= (inputs(6)) or (inputs(25));
    layer0_outputs(5104) <= (inputs(212)) and not (inputs(190));
    layer0_outputs(5105) <= not((inputs(123)) or (inputs(16)));
    layer0_outputs(5106) <= (inputs(137)) or (inputs(99));
    layer0_outputs(5107) <= (inputs(129)) xor (inputs(66));
    layer0_outputs(5108) <= not((inputs(105)) or (inputs(176)));
    layer0_outputs(5109) <= not((inputs(244)) or (inputs(186)));
    layer0_outputs(5110) <= (inputs(105)) and not (inputs(1));
    layer0_outputs(5111) <= inputs(10);
    layer0_outputs(5112) <= not((inputs(35)) and (inputs(248)));
    layer0_outputs(5113) <= not(inputs(95));
    layer0_outputs(5114) <= (inputs(136)) and not (inputs(128));
    layer0_outputs(5115) <= not(inputs(109)) or (inputs(14));
    layer0_outputs(5116) <= not((inputs(237)) or (inputs(201)));
    layer0_outputs(5117) <= (inputs(242)) and not (inputs(250));
    layer0_outputs(5118) <= (inputs(119)) or (inputs(159));
    layer0_outputs(5119) <= (inputs(72)) and not (inputs(46));
    layer0_outputs(5120) <= (inputs(138)) and not (inputs(96));
    layer0_outputs(5121) <= (inputs(117)) or (inputs(240));
    layer0_outputs(5122) <= (inputs(92)) and not (inputs(19));
    layer0_outputs(5123) <= (inputs(208)) xor (inputs(236));
    layer0_outputs(5124) <= (inputs(45)) xor (inputs(250));
    layer0_outputs(5125) <= (inputs(4)) and not (inputs(25));
    layer0_outputs(5126) <= (inputs(219)) and not (inputs(131));
    layer0_outputs(5127) <= not((inputs(155)) xor (inputs(100)));
    layer0_outputs(5128) <= (inputs(15)) or (inputs(68));
    layer0_outputs(5129) <= not(inputs(104));
    layer0_outputs(5130) <= not(inputs(228)) or (inputs(90));
    layer0_outputs(5131) <= '0';
    layer0_outputs(5132) <= inputs(104);
    layer0_outputs(5133) <= (inputs(50)) or (inputs(89));
    layer0_outputs(5134) <= (inputs(214)) or (inputs(250));
    layer0_outputs(5135) <= not(inputs(151));
    layer0_outputs(5136) <= not((inputs(77)) or (inputs(54)));
    layer0_outputs(5137) <= not((inputs(251)) xor (inputs(107)));
    layer0_outputs(5138) <= (inputs(108)) or (inputs(164));
    layer0_outputs(5139) <= inputs(202);
    layer0_outputs(5140) <= not((inputs(146)) or (inputs(235)));
    layer0_outputs(5141) <= not(inputs(155)) or (inputs(237));
    layer0_outputs(5142) <= not((inputs(136)) or (inputs(136)));
    layer0_outputs(5143) <= (inputs(230)) and not (inputs(95));
    layer0_outputs(5144) <= not(inputs(165));
    layer0_outputs(5145) <= (inputs(232)) or (inputs(136));
    layer0_outputs(5146) <= not((inputs(191)) or (inputs(102)));
    layer0_outputs(5147) <= '1';
    layer0_outputs(5148) <= not((inputs(77)) or (inputs(148)));
    layer0_outputs(5149) <= inputs(148);
    layer0_outputs(5150) <= not((inputs(182)) and (inputs(170)));
    layer0_outputs(5151) <= (inputs(176)) and (inputs(33));
    layer0_outputs(5152) <= not((inputs(42)) or (inputs(55)));
    layer0_outputs(5153) <= not((inputs(161)) xor (inputs(157)));
    layer0_outputs(5154) <= not((inputs(201)) xor (inputs(160)));
    layer0_outputs(5155) <= (inputs(180)) and not (inputs(29));
    layer0_outputs(5156) <= (inputs(189)) or (inputs(40));
    layer0_outputs(5157) <= (inputs(22)) and (inputs(254));
    layer0_outputs(5158) <= (inputs(72)) and not (inputs(163));
    layer0_outputs(5159) <= inputs(216);
    layer0_outputs(5160) <= not(inputs(251)) or (inputs(36));
    layer0_outputs(5161) <= not((inputs(229)) or (inputs(98)));
    layer0_outputs(5162) <= inputs(199);
    layer0_outputs(5163) <= inputs(161);
    layer0_outputs(5164) <= not(inputs(248));
    layer0_outputs(5165) <= not(inputs(167)) or (inputs(76));
    layer0_outputs(5166) <= not(inputs(35));
    layer0_outputs(5167) <= not((inputs(72)) xor (inputs(33)));
    layer0_outputs(5168) <= (inputs(1)) or (inputs(236));
    layer0_outputs(5169) <= inputs(146);
    layer0_outputs(5170) <= (inputs(146)) xor (inputs(15));
    layer0_outputs(5171) <= (inputs(200)) and not (inputs(66));
    layer0_outputs(5172) <= not((inputs(123)) xor (inputs(254)));
    layer0_outputs(5173) <= not(inputs(73)) or (inputs(65));
    layer0_outputs(5174) <= '0';
    layer0_outputs(5175) <= (inputs(195)) or (inputs(189));
    layer0_outputs(5176) <= inputs(36);
    layer0_outputs(5177) <= (inputs(17)) xor (inputs(121));
    layer0_outputs(5178) <= (inputs(111)) xor (inputs(24));
    layer0_outputs(5179) <= not(inputs(83)) or (inputs(215));
    layer0_outputs(5180) <= not((inputs(144)) and (inputs(130)));
    layer0_outputs(5181) <= not((inputs(118)) xor (inputs(65)));
    layer0_outputs(5182) <= not((inputs(173)) xor (inputs(87)));
    layer0_outputs(5183) <= (inputs(197)) or (inputs(170));
    layer0_outputs(5184) <= not((inputs(6)) xor (inputs(92)));
    layer0_outputs(5185) <= (inputs(133)) and not (inputs(133));
    layer0_outputs(5186) <= (inputs(145)) or (inputs(176));
    layer0_outputs(5187) <= '0';
    layer0_outputs(5188) <= (inputs(42)) and (inputs(25));
    layer0_outputs(5189) <= not((inputs(114)) xor (inputs(251)));
    layer0_outputs(5190) <= (inputs(72)) or (inputs(255));
    layer0_outputs(5191) <= (inputs(134)) xor (inputs(148));
    layer0_outputs(5192) <= not(inputs(173));
    layer0_outputs(5193) <= not(inputs(253)) or (inputs(242));
    layer0_outputs(5194) <= inputs(139);
    layer0_outputs(5195) <= not(inputs(151));
    layer0_outputs(5196) <= not((inputs(37)) or (inputs(132)));
    layer0_outputs(5197) <= not((inputs(45)) or (inputs(149)));
    layer0_outputs(5198) <= not(inputs(12));
    layer0_outputs(5199) <= inputs(163);
    layer0_outputs(5200) <= not(inputs(139)) or (inputs(185));
    layer0_outputs(5201) <= not(inputs(119));
    layer0_outputs(5202) <= inputs(119);
    layer0_outputs(5203) <= (inputs(35)) and (inputs(94));
    layer0_outputs(5204) <= (inputs(133)) and not (inputs(146));
    layer0_outputs(5205) <= not(inputs(153));
    layer0_outputs(5206) <= '1';
    layer0_outputs(5207) <= not(inputs(72)) or (inputs(248));
    layer0_outputs(5208) <= not((inputs(76)) xor (inputs(182)));
    layer0_outputs(5209) <= not(inputs(28));
    layer0_outputs(5210) <= inputs(168);
    layer0_outputs(5211) <= not((inputs(149)) or (inputs(248)));
    layer0_outputs(5212) <= not((inputs(28)) xor (inputs(24)));
    layer0_outputs(5213) <= not((inputs(158)) or (inputs(99)));
    layer0_outputs(5214) <= not((inputs(58)) xor (inputs(133)));
    layer0_outputs(5215) <= not((inputs(174)) and (inputs(211)));
    layer0_outputs(5216) <= not(inputs(75));
    layer0_outputs(5217) <= not(inputs(58)) or (inputs(22));
    layer0_outputs(5218) <= not((inputs(190)) or (inputs(160)));
    layer0_outputs(5219) <= (inputs(168)) or (inputs(132));
    layer0_outputs(5220) <= not(inputs(15));
    layer0_outputs(5221) <= not(inputs(118)) or (inputs(14));
    layer0_outputs(5222) <= inputs(202);
    layer0_outputs(5223) <= not((inputs(94)) xor (inputs(144)));
    layer0_outputs(5224) <= not(inputs(163));
    layer0_outputs(5225) <= inputs(151);
    layer0_outputs(5226) <= not(inputs(172));
    layer0_outputs(5227) <= not((inputs(249)) or (inputs(169)));
    layer0_outputs(5228) <= (inputs(144)) or (inputs(11));
    layer0_outputs(5229) <= not((inputs(11)) or (inputs(132)));
    layer0_outputs(5230) <= not((inputs(165)) or (inputs(67)));
    layer0_outputs(5231) <= not(inputs(147)) or (inputs(244));
    layer0_outputs(5232) <= (inputs(150)) or (inputs(41));
    layer0_outputs(5233) <= not((inputs(126)) xor (inputs(76)));
    layer0_outputs(5234) <= not(inputs(20));
    layer0_outputs(5235) <= (inputs(101)) or (inputs(27));
    layer0_outputs(5236) <= (inputs(214)) xor (inputs(58));
    layer0_outputs(5237) <= not((inputs(25)) or (inputs(149)));
    layer0_outputs(5238) <= (inputs(253)) xor (inputs(49));
    layer0_outputs(5239) <= (inputs(23)) and not (inputs(212));
    layer0_outputs(5240) <= (inputs(204)) or (inputs(46));
    layer0_outputs(5241) <= (inputs(199)) or (inputs(241));
    layer0_outputs(5242) <= (inputs(215)) or (inputs(34));
    layer0_outputs(5243) <= (inputs(63)) xor (inputs(136));
    layer0_outputs(5244) <= not((inputs(116)) xor (inputs(44)));
    layer0_outputs(5245) <= not(inputs(149)) or (inputs(39));
    layer0_outputs(5246) <= not(inputs(50)) or (inputs(93));
    layer0_outputs(5247) <= (inputs(204)) and (inputs(13));
    layer0_outputs(5248) <= (inputs(199)) and not (inputs(217));
    layer0_outputs(5249) <= not((inputs(2)) xor (inputs(217)));
    layer0_outputs(5250) <= inputs(217);
    layer0_outputs(5251) <= inputs(165);
    layer0_outputs(5252) <= (inputs(150)) and not (inputs(46));
    layer0_outputs(5253) <= (inputs(214)) xor (inputs(64));
    layer0_outputs(5254) <= inputs(195);
    layer0_outputs(5255) <= not((inputs(191)) or (inputs(170)));
    layer0_outputs(5256) <= not((inputs(65)) xor (inputs(19)));
    layer0_outputs(5257) <= (inputs(31)) xor (inputs(233));
    layer0_outputs(5258) <= (inputs(85)) and not (inputs(77));
    layer0_outputs(5259) <= not((inputs(33)) or (inputs(228)));
    layer0_outputs(5260) <= (inputs(76)) or (inputs(25));
    layer0_outputs(5261) <= not(inputs(107)) or (inputs(160));
    layer0_outputs(5262) <= not(inputs(150));
    layer0_outputs(5263) <= not((inputs(120)) or (inputs(228)));
    layer0_outputs(5264) <= not(inputs(18));
    layer0_outputs(5265) <= (inputs(50)) and (inputs(47));
    layer0_outputs(5266) <= not((inputs(176)) or (inputs(136)));
    layer0_outputs(5267) <= (inputs(74)) and not (inputs(255));
    layer0_outputs(5268) <= (inputs(132)) or (inputs(92));
    layer0_outputs(5269) <= (inputs(182)) and not (inputs(184));
    layer0_outputs(5270) <= not((inputs(73)) or (inputs(1)));
    layer0_outputs(5271) <= not((inputs(186)) or (inputs(40)));
    layer0_outputs(5272) <= not((inputs(213)) or (inputs(84)));
    layer0_outputs(5273) <= '1';
    layer0_outputs(5274) <= inputs(107);
    layer0_outputs(5275) <= not(inputs(148)) or (inputs(107));
    layer0_outputs(5276) <= (inputs(193)) or (inputs(40));
    layer0_outputs(5277) <= inputs(40);
    layer0_outputs(5278) <= inputs(195);
    layer0_outputs(5279) <= not(inputs(255));
    layer0_outputs(5280) <= inputs(73);
    layer0_outputs(5281) <= (inputs(218)) or (inputs(31));
    layer0_outputs(5282) <= (inputs(143)) xor (inputs(38));
    layer0_outputs(5283) <= (inputs(73)) xor (inputs(235));
    layer0_outputs(5284) <= not(inputs(45));
    layer0_outputs(5285) <= inputs(170);
    layer0_outputs(5286) <= not((inputs(200)) and (inputs(213)));
    layer0_outputs(5287) <= inputs(140);
    layer0_outputs(5288) <= (inputs(157)) or (inputs(108));
    layer0_outputs(5289) <= (inputs(104)) xor (inputs(134));
    layer0_outputs(5290) <= not((inputs(243)) xor (inputs(105)));
    layer0_outputs(5291) <= not(inputs(22));
    layer0_outputs(5292) <= inputs(150);
    layer0_outputs(5293) <= not(inputs(168)) or (inputs(180));
    layer0_outputs(5294) <= not(inputs(238)) or (inputs(43));
    layer0_outputs(5295) <= inputs(196);
    layer0_outputs(5296) <= inputs(24);
    layer0_outputs(5297) <= '0';
    layer0_outputs(5298) <= not((inputs(215)) xor (inputs(24)));
    layer0_outputs(5299) <= not(inputs(121)) or (inputs(176));
    layer0_outputs(5300) <= not(inputs(109));
    layer0_outputs(5301) <= not((inputs(165)) or (inputs(124)));
    layer0_outputs(5302) <= '0';
    layer0_outputs(5303) <= not(inputs(98));
    layer0_outputs(5304) <= not((inputs(83)) or (inputs(71)));
    layer0_outputs(5305) <= inputs(86);
    layer0_outputs(5306) <= not(inputs(102)) or (inputs(125));
    layer0_outputs(5307) <= not((inputs(9)) and (inputs(2)));
    layer0_outputs(5308) <= not(inputs(152));
    layer0_outputs(5309) <= '0';
    layer0_outputs(5310) <= not((inputs(6)) xor (inputs(231)));
    layer0_outputs(5311) <= '0';
    layer0_outputs(5312) <= (inputs(225)) or (inputs(54));
    layer0_outputs(5313) <= inputs(34);
    layer0_outputs(5314) <= not(inputs(115));
    layer0_outputs(5315) <= inputs(50);
    layer0_outputs(5316) <= not((inputs(162)) or (inputs(69)));
    layer0_outputs(5317) <= not((inputs(238)) xor (inputs(166)));
    layer0_outputs(5318) <= (inputs(113)) xor (inputs(162));
    layer0_outputs(5319) <= not((inputs(188)) xor (inputs(194)));
    layer0_outputs(5320) <= not((inputs(64)) and (inputs(33)));
    layer0_outputs(5321) <= not(inputs(185)) or (inputs(89));
    layer0_outputs(5322) <= inputs(125);
    layer0_outputs(5323) <= not(inputs(98)) or (inputs(226));
    layer0_outputs(5324) <= (inputs(122)) or (inputs(143));
    layer0_outputs(5325) <= not(inputs(89)) or (inputs(116));
    layer0_outputs(5326) <= (inputs(100)) or (inputs(221));
    layer0_outputs(5327) <= (inputs(133)) and not (inputs(230));
    layer0_outputs(5328) <= not(inputs(87)) or (inputs(254));
    layer0_outputs(5329) <= inputs(119);
    layer0_outputs(5330) <= (inputs(115)) xor (inputs(5));
    layer0_outputs(5331) <= (inputs(235)) and not (inputs(66));
    layer0_outputs(5332) <= not(inputs(41)) or (inputs(25));
    layer0_outputs(5333) <= (inputs(244)) and not (inputs(64));
    layer0_outputs(5334) <= (inputs(55)) and not (inputs(162));
    layer0_outputs(5335) <= (inputs(154)) xor (inputs(117));
    layer0_outputs(5336) <= (inputs(158)) or (inputs(185));
    layer0_outputs(5337) <= not(inputs(249));
    layer0_outputs(5338) <= (inputs(170)) and not (inputs(245));
    layer0_outputs(5339) <= not((inputs(161)) and (inputs(61)));
    layer0_outputs(5340) <= not(inputs(33)) or (inputs(126));
    layer0_outputs(5341) <= (inputs(255)) and (inputs(42));
    layer0_outputs(5342) <= not(inputs(171)) or (inputs(221));
    layer0_outputs(5343) <= not((inputs(54)) or (inputs(76)));
    layer0_outputs(5344) <= '1';
    layer0_outputs(5345) <= not(inputs(132)) or (inputs(247));
    layer0_outputs(5346) <= (inputs(195)) and not (inputs(175));
    layer0_outputs(5347) <= (inputs(181)) xor (inputs(72));
    layer0_outputs(5348) <= inputs(158);
    layer0_outputs(5349) <= (inputs(125)) and (inputs(76));
    layer0_outputs(5350) <= inputs(92);
    layer0_outputs(5351) <= not(inputs(180));
    layer0_outputs(5352) <= '1';
    layer0_outputs(5353) <= inputs(107);
    layer0_outputs(5354) <= (inputs(140)) and not (inputs(237));
    layer0_outputs(5355) <= not(inputs(126)) or (inputs(48));
    layer0_outputs(5356) <= (inputs(161)) xor (inputs(70));
    layer0_outputs(5357) <= not((inputs(28)) xor (inputs(37)));
    layer0_outputs(5358) <= not((inputs(72)) or (inputs(172)));
    layer0_outputs(5359) <= not((inputs(46)) xor (inputs(149)));
    layer0_outputs(5360) <= not((inputs(231)) xor (inputs(51)));
    layer0_outputs(5361) <= (inputs(123)) or (inputs(115));
    layer0_outputs(5362) <= inputs(105);
    layer0_outputs(5363) <= (inputs(104)) and not (inputs(70));
    layer0_outputs(5364) <= inputs(33);
    layer0_outputs(5365) <= (inputs(117)) and not (inputs(156));
    layer0_outputs(5366) <= inputs(85);
    layer0_outputs(5367) <= (inputs(14)) and not (inputs(27));
    layer0_outputs(5368) <= not(inputs(71)) or (inputs(157));
    layer0_outputs(5369) <= (inputs(153)) and not (inputs(204));
    layer0_outputs(5370) <= (inputs(44)) or (inputs(255));
    layer0_outputs(5371) <= (inputs(68)) xor (inputs(39));
    layer0_outputs(5372) <= (inputs(188)) or (inputs(10));
    layer0_outputs(5373) <= (inputs(30)) or (inputs(162));
    layer0_outputs(5374) <= (inputs(57)) and not (inputs(70));
    layer0_outputs(5375) <= not(inputs(80));
    layer0_outputs(5376) <= (inputs(193)) xor (inputs(185));
    layer0_outputs(5377) <= not(inputs(89));
    layer0_outputs(5378) <= not(inputs(189));
    layer0_outputs(5379) <= not(inputs(71));
    layer0_outputs(5380) <= (inputs(152)) and not (inputs(158));
    layer0_outputs(5381) <= (inputs(62)) or (inputs(52));
    layer0_outputs(5382) <= (inputs(93)) and not (inputs(251));
    layer0_outputs(5383) <= '0';
    layer0_outputs(5384) <= inputs(59);
    layer0_outputs(5385) <= (inputs(254)) xor (inputs(202));
    layer0_outputs(5386) <= not((inputs(120)) or (inputs(189)));
    layer0_outputs(5387) <= not((inputs(147)) xor (inputs(91)));
    layer0_outputs(5388) <= inputs(131);
    layer0_outputs(5389) <= not(inputs(102)) or (inputs(108));
    layer0_outputs(5390) <= (inputs(220)) xor (inputs(118));
    layer0_outputs(5391) <= (inputs(103)) or (inputs(31));
    layer0_outputs(5392) <= not(inputs(148));
    layer0_outputs(5393) <= (inputs(225)) and (inputs(190));
    layer0_outputs(5394) <= not((inputs(63)) xor (inputs(84)));
    layer0_outputs(5395) <= not((inputs(54)) or (inputs(107)));
    layer0_outputs(5396) <= inputs(143);
    layer0_outputs(5397) <= (inputs(197)) xor (inputs(182));
    layer0_outputs(5398) <= inputs(196);
    layer0_outputs(5399) <= '1';
    layer0_outputs(5400) <= not(inputs(53)) or (inputs(177));
    layer0_outputs(5401) <= inputs(178);
    layer0_outputs(5402) <= inputs(152);
    layer0_outputs(5403) <= not((inputs(252)) or (inputs(156)));
    layer0_outputs(5404) <= (inputs(214)) or (inputs(155));
    layer0_outputs(5405) <= not((inputs(70)) xor (inputs(31)));
    layer0_outputs(5406) <= not(inputs(180));
    layer0_outputs(5407) <= not(inputs(151)) or (inputs(72));
    layer0_outputs(5408) <= not((inputs(183)) xor (inputs(216)));
    layer0_outputs(5409) <= (inputs(123)) and not (inputs(119));
    layer0_outputs(5410) <= not(inputs(29)) or (inputs(9));
    layer0_outputs(5411) <= (inputs(182)) or (inputs(112));
    layer0_outputs(5412) <= not((inputs(154)) or (inputs(255)));
    layer0_outputs(5413) <= (inputs(213)) or (inputs(53));
    layer0_outputs(5414) <= not((inputs(129)) xor (inputs(133)));
    layer0_outputs(5415) <= not(inputs(171)) or (inputs(18));
    layer0_outputs(5416) <= not(inputs(69)) or (inputs(140));
    layer0_outputs(5417) <= not((inputs(223)) xor (inputs(124)));
    layer0_outputs(5418) <= not((inputs(10)) or (inputs(5)));
    layer0_outputs(5419) <= (inputs(161)) or (inputs(199));
    layer0_outputs(5420) <= not(inputs(173)) or (inputs(112));
    layer0_outputs(5421) <= (inputs(166)) and not (inputs(208));
    layer0_outputs(5422) <= '0';
    layer0_outputs(5423) <= not(inputs(155));
    layer0_outputs(5424) <= not(inputs(170));
    layer0_outputs(5425) <= not(inputs(39));
    layer0_outputs(5426) <= not(inputs(96));
    layer0_outputs(5427) <= (inputs(65)) or (inputs(220));
    layer0_outputs(5428) <= (inputs(180)) or (inputs(134));
    layer0_outputs(5429) <= (inputs(36)) and not (inputs(255));
    layer0_outputs(5430) <= (inputs(172)) and not (inputs(146));
    layer0_outputs(5431) <= not(inputs(217)) or (inputs(89));
    layer0_outputs(5432) <= not(inputs(52));
    layer0_outputs(5433) <= inputs(172);
    layer0_outputs(5434) <= inputs(181);
    layer0_outputs(5435) <= inputs(61);
    layer0_outputs(5436) <= not(inputs(100)) or (inputs(210));
    layer0_outputs(5437) <= inputs(143);
    layer0_outputs(5438) <= not(inputs(153));
    layer0_outputs(5439) <= not((inputs(189)) or (inputs(166)));
    layer0_outputs(5440) <= (inputs(114)) and not (inputs(238));
    layer0_outputs(5441) <= (inputs(73)) and not (inputs(110));
    layer0_outputs(5442) <= inputs(218);
    layer0_outputs(5443) <= not((inputs(102)) or (inputs(96)));
    layer0_outputs(5444) <= (inputs(172)) xor (inputs(42));
    layer0_outputs(5445) <= (inputs(16)) xor (inputs(212));
    layer0_outputs(5446) <= (inputs(225)) and not (inputs(159));
    layer0_outputs(5447) <= (inputs(151)) or (inputs(39));
    layer0_outputs(5448) <= (inputs(68)) and not (inputs(28));
    layer0_outputs(5449) <= not((inputs(178)) and (inputs(15)));
    layer0_outputs(5450) <= '1';
    layer0_outputs(5451) <= (inputs(71)) and not (inputs(203));
    layer0_outputs(5452) <= (inputs(3)) or (inputs(58));
    layer0_outputs(5453) <= (inputs(88)) xor (inputs(195));
    layer0_outputs(5454) <= (inputs(132)) and not (inputs(81));
    layer0_outputs(5455) <= not(inputs(23));
    layer0_outputs(5456) <= not(inputs(170)) or (inputs(75));
    layer0_outputs(5457) <= not((inputs(231)) or (inputs(253)));
    layer0_outputs(5458) <= not(inputs(127));
    layer0_outputs(5459) <= (inputs(157)) or (inputs(126));
    layer0_outputs(5460) <= '0';
    layer0_outputs(5461) <= inputs(121);
    layer0_outputs(5462) <= (inputs(252)) and not (inputs(152));
    layer0_outputs(5463) <= (inputs(160)) or (inputs(52));
    layer0_outputs(5464) <= not(inputs(187)) or (inputs(4));
    layer0_outputs(5465) <= not(inputs(63)) or (inputs(174));
    layer0_outputs(5466) <= not(inputs(146)) or (inputs(124));
    layer0_outputs(5467) <= (inputs(74)) xor (inputs(105));
    layer0_outputs(5468) <= not((inputs(123)) or (inputs(244)));
    layer0_outputs(5469) <= (inputs(182)) and not (inputs(87));
    layer0_outputs(5470) <= (inputs(123)) or (inputs(102));
    layer0_outputs(5471) <= (inputs(3)) and not (inputs(34));
    layer0_outputs(5472) <= not((inputs(109)) or (inputs(225)));
    layer0_outputs(5473) <= inputs(134);
    layer0_outputs(5474) <= not(inputs(116));
    layer0_outputs(5475) <= inputs(125);
    layer0_outputs(5476) <= not((inputs(222)) xor (inputs(147)));
    layer0_outputs(5477) <= '0';
    layer0_outputs(5478) <= (inputs(112)) or (inputs(40));
    layer0_outputs(5479) <= not(inputs(217)) or (inputs(199));
    layer0_outputs(5480) <= inputs(40);
    layer0_outputs(5481) <= inputs(202);
    layer0_outputs(5482) <= inputs(7);
    layer0_outputs(5483) <= not(inputs(253)) or (inputs(206));
    layer0_outputs(5484) <= (inputs(206)) or (inputs(127));
    layer0_outputs(5485) <= (inputs(184)) and not (inputs(253));
    layer0_outputs(5486) <= not(inputs(93)) or (inputs(29));
    layer0_outputs(5487) <= inputs(143);
    layer0_outputs(5488) <= not((inputs(14)) xor (inputs(154)));
    layer0_outputs(5489) <= not((inputs(121)) or (inputs(255)));
    layer0_outputs(5490) <= (inputs(102)) and not (inputs(4));
    layer0_outputs(5491) <= (inputs(63)) and not (inputs(160));
    layer0_outputs(5492) <= (inputs(195)) and not (inputs(78));
    layer0_outputs(5493) <= not((inputs(4)) xor (inputs(80)));
    layer0_outputs(5494) <= inputs(232);
    layer0_outputs(5495) <= not((inputs(133)) xor (inputs(238)));
    layer0_outputs(5496) <= (inputs(112)) or (inputs(215));
    layer0_outputs(5497) <= (inputs(185)) or (inputs(6));
    layer0_outputs(5498) <= not(inputs(104));
    layer0_outputs(5499) <= not((inputs(151)) or (inputs(30)));
    layer0_outputs(5500) <= inputs(151);
    layer0_outputs(5501) <= not(inputs(175));
    layer0_outputs(5502) <= not(inputs(12));
    layer0_outputs(5503) <= inputs(88);
    layer0_outputs(5504) <= not((inputs(155)) xor (inputs(52)));
    layer0_outputs(5505) <= not((inputs(47)) and (inputs(159)));
    layer0_outputs(5506) <= not(inputs(166)) or (inputs(94));
    layer0_outputs(5507) <= not(inputs(195)) or (inputs(158));
    layer0_outputs(5508) <= not(inputs(123)) or (inputs(161));
    layer0_outputs(5509) <= (inputs(56)) and not (inputs(51));
    layer0_outputs(5510) <= not(inputs(254));
    layer0_outputs(5511) <= not((inputs(140)) xor (inputs(207)));
    layer0_outputs(5512) <= (inputs(114)) and not (inputs(243));
    layer0_outputs(5513) <= not(inputs(214)) or (inputs(60));
    layer0_outputs(5514) <= not(inputs(89));
    layer0_outputs(5515) <= (inputs(157)) and (inputs(162));
    layer0_outputs(5516) <= not((inputs(32)) xor (inputs(132)));
    layer0_outputs(5517) <= (inputs(214)) or (inputs(195));
    layer0_outputs(5518) <= not(inputs(158));
    layer0_outputs(5519) <= (inputs(128)) or (inputs(32));
    layer0_outputs(5520) <= inputs(131);
    layer0_outputs(5521) <= (inputs(23)) and not (inputs(52));
    layer0_outputs(5522) <= not(inputs(13));
    layer0_outputs(5523) <= not(inputs(215)) or (inputs(45));
    layer0_outputs(5524) <= not((inputs(98)) and (inputs(11)));
    layer0_outputs(5525) <= (inputs(237)) xor (inputs(134));
    layer0_outputs(5526) <= not(inputs(231)) or (inputs(21));
    layer0_outputs(5527) <= (inputs(159)) xor (inputs(233));
    layer0_outputs(5528) <= '1';
    layer0_outputs(5529) <= not((inputs(244)) or (inputs(38)));
    layer0_outputs(5530) <= (inputs(38)) or (inputs(37));
    layer0_outputs(5531) <= inputs(90);
    layer0_outputs(5532) <= '1';
    layer0_outputs(5533) <= '1';
    layer0_outputs(5534) <= (inputs(186)) or (inputs(97));
    layer0_outputs(5535) <= not(inputs(134)) or (inputs(190));
    layer0_outputs(5536) <= (inputs(72)) xor (inputs(157));
    layer0_outputs(5537) <= not(inputs(104));
    layer0_outputs(5538) <= not((inputs(80)) or (inputs(40)));
    layer0_outputs(5539) <= (inputs(86)) xor (inputs(171));
    layer0_outputs(5540) <= (inputs(121)) or (inputs(31));
    layer0_outputs(5541) <= inputs(247);
    layer0_outputs(5542) <= not(inputs(132));
    layer0_outputs(5543) <= '1';
    layer0_outputs(5544) <= (inputs(187)) and not (inputs(48));
    layer0_outputs(5545) <= (inputs(167)) and (inputs(232));
    layer0_outputs(5546) <= '1';
    layer0_outputs(5547) <= (inputs(103)) and not (inputs(67));
    layer0_outputs(5548) <= '0';
    layer0_outputs(5549) <= not((inputs(108)) xor (inputs(12)));
    layer0_outputs(5550) <= not((inputs(250)) xor (inputs(237)));
    layer0_outputs(5551) <= not(inputs(212)) or (inputs(21));
    layer0_outputs(5552) <= (inputs(52)) or (inputs(35));
    layer0_outputs(5553) <= not((inputs(252)) or (inputs(153)));
    layer0_outputs(5554) <= (inputs(156)) or (inputs(11));
    layer0_outputs(5555) <= inputs(167);
    layer0_outputs(5556) <= not((inputs(223)) xor (inputs(43)));
    layer0_outputs(5557) <= (inputs(136)) or (inputs(226));
    layer0_outputs(5558) <= not(inputs(76));
    layer0_outputs(5559) <= not(inputs(152)) or (inputs(231));
    layer0_outputs(5560) <= (inputs(160)) and not (inputs(250));
    layer0_outputs(5561) <= not(inputs(120));
    layer0_outputs(5562) <= (inputs(66)) xor (inputs(23));
    layer0_outputs(5563) <= inputs(171);
    layer0_outputs(5564) <= (inputs(34)) and (inputs(106));
    layer0_outputs(5565) <= not((inputs(35)) or (inputs(39)));
    layer0_outputs(5566) <= not((inputs(109)) and (inputs(59)));
    layer0_outputs(5567) <= not((inputs(222)) or (inputs(163)));
    layer0_outputs(5568) <= not((inputs(160)) xor (inputs(39)));
    layer0_outputs(5569) <= not(inputs(96));
    layer0_outputs(5570) <= not((inputs(120)) or (inputs(183)));
    layer0_outputs(5571) <= not(inputs(84)) or (inputs(238));
    layer0_outputs(5572) <= inputs(190);
    layer0_outputs(5573) <= not((inputs(202)) or (inputs(93)));
    layer0_outputs(5574) <= not((inputs(156)) xor (inputs(108)));
    layer0_outputs(5575) <= (inputs(222)) xor (inputs(218));
    layer0_outputs(5576) <= inputs(167);
    layer0_outputs(5577) <= not(inputs(151));
    layer0_outputs(5578) <= (inputs(39)) or (inputs(129));
    layer0_outputs(5579) <= (inputs(45)) xor (inputs(249));
    layer0_outputs(5580) <= inputs(131);
    layer0_outputs(5581) <= not((inputs(43)) or (inputs(212)));
    layer0_outputs(5582) <= (inputs(149)) and not (inputs(212));
    layer0_outputs(5583) <= not(inputs(206)) or (inputs(243));
    layer0_outputs(5584) <= (inputs(120)) xor (inputs(79));
    layer0_outputs(5585) <= (inputs(20)) xor (inputs(196));
    layer0_outputs(5586) <= not(inputs(224)) or (inputs(80));
    layer0_outputs(5587) <= (inputs(67)) or (inputs(158));
    layer0_outputs(5588) <= (inputs(38)) xor (inputs(197));
    layer0_outputs(5589) <= (inputs(144)) or (inputs(169));
    layer0_outputs(5590) <= (inputs(71)) and not (inputs(192));
    layer0_outputs(5591) <= inputs(153);
    layer0_outputs(5592) <= (inputs(155)) xor (inputs(138));
    layer0_outputs(5593) <= not((inputs(100)) xor (inputs(190)));
    layer0_outputs(5594) <= not(inputs(89)) or (inputs(237));
    layer0_outputs(5595) <= (inputs(106)) and not (inputs(131));
    layer0_outputs(5596) <= inputs(96);
    layer0_outputs(5597) <= not(inputs(74));
    layer0_outputs(5598) <= (inputs(163)) and not (inputs(33));
    layer0_outputs(5599) <= not(inputs(41));
    layer0_outputs(5600) <= (inputs(169)) or (inputs(189));
    layer0_outputs(5601) <= inputs(137);
    layer0_outputs(5602) <= not((inputs(75)) and (inputs(217)));
    layer0_outputs(5603) <= not(inputs(61)) or (inputs(236));
    layer0_outputs(5604) <= (inputs(81)) or (inputs(90));
    layer0_outputs(5605) <= (inputs(63)) xor (inputs(120));
    layer0_outputs(5606) <= (inputs(71)) xor (inputs(255));
    layer0_outputs(5607) <= not(inputs(212)) or (inputs(4));
    layer0_outputs(5608) <= not(inputs(122));
    layer0_outputs(5609) <= not((inputs(30)) xor (inputs(175)));
    layer0_outputs(5610) <= not((inputs(164)) or (inputs(36)));
    layer0_outputs(5611) <= (inputs(71)) and not (inputs(167));
    layer0_outputs(5612) <= not(inputs(152));
    layer0_outputs(5613) <= not(inputs(59)) or (inputs(35));
    layer0_outputs(5614) <= not(inputs(187));
    layer0_outputs(5615) <= not((inputs(57)) xor (inputs(70)));
    layer0_outputs(5616) <= not(inputs(118));
    layer0_outputs(5617) <= not((inputs(7)) or (inputs(143)));
    layer0_outputs(5618) <= '1';
    layer0_outputs(5619) <= not(inputs(69));
    layer0_outputs(5620) <= not((inputs(162)) xor (inputs(230)));
    layer0_outputs(5621) <= not(inputs(117)) or (inputs(15));
    layer0_outputs(5622) <= (inputs(149)) xor (inputs(141));
    layer0_outputs(5623) <= not((inputs(209)) xor (inputs(226)));
    layer0_outputs(5624) <= (inputs(43)) xor (inputs(130));
    layer0_outputs(5625) <= not(inputs(170));
    layer0_outputs(5626) <= (inputs(184)) xor (inputs(216));
    layer0_outputs(5627) <= (inputs(11)) and not (inputs(144));
    layer0_outputs(5628) <= not((inputs(138)) xor (inputs(242)));
    layer0_outputs(5629) <= not(inputs(119));
    layer0_outputs(5630) <= (inputs(145)) or (inputs(200));
    layer0_outputs(5631) <= not((inputs(8)) xor (inputs(235)));
    layer0_outputs(5632) <= not((inputs(20)) xor (inputs(203)));
    layer0_outputs(5633) <= not(inputs(231));
    layer0_outputs(5634) <= not((inputs(7)) or (inputs(113)));
    layer0_outputs(5635) <= (inputs(40)) and not (inputs(186));
    layer0_outputs(5636) <= inputs(133);
    layer0_outputs(5637) <= (inputs(85)) xor (inputs(92));
    layer0_outputs(5638) <= (inputs(164)) xor (inputs(51));
    layer0_outputs(5639) <= (inputs(140)) or (inputs(25));
    layer0_outputs(5640) <= (inputs(188)) or (inputs(178));
    layer0_outputs(5641) <= inputs(219);
    layer0_outputs(5642) <= (inputs(80)) and not (inputs(193));
    layer0_outputs(5643) <= not(inputs(107)) or (inputs(218));
    layer0_outputs(5644) <= not(inputs(202));
    layer0_outputs(5645) <= not((inputs(55)) xor (inputs(170)));
    layer0_outputs(5646) <= not(inputs(46));
    layer0_outputs(5647) <= not((inputs(125)) or (inputs(76)));
    layer0_outputs(5648) <= not((inputs(13)) xor (inputs(52)));
    layer0_outputs(5649) <= '0';
    layer0_outputs(5650) <= inputs(56);
    layer0_outputs(5651) <= (inputs(114)) and not (inputs(37));
    layer0_outputs(5652) <= (inputs(28)) and not (inputs(143));
    layer0_outputs(5653) <= not(inputs(253));
    layer0_outputs(5654) <= (inputs(93)) or (inputs(85));
    layer0_outputs(5655) <= not(inputs(221));
    layer0_outputs(5656) <= not((inputs(211)) xor (inputs(127)));
    layer0_outputs(5657) <= (inputs(52)) or (inputs(153));
    layer0_outputs(5658) <= (inputs(40)) and not (inputs(88));
    layer0_outputs(5659) <= (inputs(249)) and not (inputs(129));
    layer0_outputs(5660) <= inputs(117);
    layer0_outputs(5661) <= '1';
    layer0_outputs(5662) <= inputs(150);
    layer0_outputs(5663) <= not((inputs(152)) or (inputs(206)));
    layer0_outputs(5664) <= (inputs(85)) xor (inputs(191));
    layer0_outputs(5665) <= (inputs(76)) and not (inputs(87));
    layer0_outputs(5666) <= not((inputs(97)) xor (inputs(205)));
    layer0_outputs(5667) <= (inputs(115)) or (inputs(230));
    layer0_outputs(5668) <= not(inputs(159));
    layer0_outputs(5669) <= not((inputs(178)) or (inputs(2)));
    layer0_outputs(5670) <= inputs(105);
    layer0_outputs(5671) <= (inputs(90)) and not (inputs(43));
    layer0_outputs(5672) <= (inputs(84)) xor (inputs(132));
    layer0_outputs(5673) <= not((inputs(60)) and (inputs(127)));
    layer0_outputs(5674) <= (inputs(43)) and not (inputs(239));
    layer0_outputs(5675) <= (inputs(251)) and (inputs(95));
    layer0_outputs(5676) <= not(inputs(37));
    layer0_outputs(5677) <= not((inputs(134)) or (inputs(205)));
    layer0_outputs(5678) <= (inputs(226)) or (inputs(143));
    layer0_outputs(5679) <= not((inputs(138)) xor (inputs(228)));
    layer0_outputs(5680) <= not(inputs(55));
    layer0_outputs(5681) <= not(inputs(60)) or (inputs(37));
    layer0_outputs(5682) <= not(inputs(210)) or (inputs(245));
    layer0_outputs(5683) <= not((inputs(205)) xor (inputs(10)));
    layer0_outputs(5684) <= not(inputs(78)) or (inputs(62));
    layer0_outputs(5685) <= (inputs(169)) and not (inputs(46));
    layer0_outputs(5686) <= not(inputs(35));
    layer0_outputs(5687) <= (inputs(233)) and not (inputs(250));
    layer0_outputs(5688) <= not((inputs(209)) or (inputs(238)));
    layer0_outputs(5689) <= (inputs(96)) and not (inputs(1));
    layer0_outputs(5690) <= not(inputs(202)) or (inputs(225));
    layer0_outputs(5691) <= (inputs(180)) or (inputs(19));
    layer0_outputs(5692) <= inputs(53);
    layer0_outputs(5693) <= not((inputs(233)) or (inputs(150)));
    layer0_outputs(5694) <= not(inputs(169));
    layer0_outputs(5695) <= (inputs(205)) or (inputs(65));
    layer0_outputs(5696) <= not(inputs(9)) or (inputs(81));
    layer0_outputs(5697) <= not((inputs(128)) or (inputs(229)));
    layer0_outputs(5698) <= inputs(109);
    layer0_outputs(5699) <= not(inputs(178)) or (inputs(206));
    layer0_outputs(5700) <= (inputs(229)) and not (inputs(232));
    layer0_outputs(5701) <= (inputs(194)) or (inputs(23));
    layer0_outputs(5702) <= (inputs(63)) xor (inputs(93));
    layer0_outputs(5703) <= not(inputs(94)) or (inputs(80));
    layer0_outputs(5704) <= not((inputs(142)) xor (inputs(193)));
    layer0_outputs(5705) <= not(inputs(86));
    layer0_outputs(5706) <= inputs(198);
    layer0_outputs(5707) <= inputs(58);
    layer0_outputs(5708) <= (inputs(57)) xor (inputs(38));
    layer0_outputs(5709) <= not(inputs(180)) or (inputs(88));
    layer0_outputs(5710) <= inputs(101);
    layer0_outputs(5711) <= (inputs(119)) or (inputs(38));
    layer0_outputs(5712) <= (inputs(5)) xor (inputs(220));
    layer0_outputs(5713) <= (inputs(217)) and not (inputs(200));
    layer0_outputs(5714) <= inputs(123);
    layer0_outputs(5715) <= (inputs(21)) xor (inputs(147));
    layer0_outputs(5716) <= not((inputs(153)) or (inputs(74)));
    layer0_outputs(5717) <= inputs(113);
    layer0_outputs(5718) <= '1';
    layer0_outputs(5719) <= not((inputs(225)) xor (inputs(171)));
    layer0_outputs(5720) <= not(inputs(217)) or (inputs(11));
    layer0_outputs(5721) <= not((inputs(243)) or (inputs(87)));
    layer0_outputs(5722) <= not(inputs(218));
    layer0_outputs(5723) <= not(inputs(58));
    layer0_outputs(5724) <= (inputs(65)) and not (inputs(5));
    layer0_outputs(5725) <= not(inputs(10));
    layer0_outputs(5726) <= (inputs(194)) and (inputs(239));
    layer0_outputs(5727) <= (inputs(116)) and not (inputs(193));
    layer0_outputs(5728) <= not((inputs(253)) or (inputs(181)));
    layer0_outputs(5729) <= (inputs(16)) and not (inputs(141));
    layer0_outputs(5730) <= not((inputs(191)) and (inputs(110)));
    layer0_outputs(5731) <= inputs(61);
    layer0_outputs(5732) <= (inputs(175)) xor (inputs(82));
    layer0_outputs(5733) <= inputs(13);
    layer0_outputs(5734) <= (inputs(140)) and not (inputs(238));
    layer0_outputs(5735) <= not(inputs(83));
    layer0_outputs(5736) <= not(inputs(164));
    layer0_outputs(5737) <= not((inputs(24)) xor (inputs(181)));
    layer0_outputs(5738) <= (inputs(74)) or (inputs(194));
    layer0_outputs(5739) <= not((inputs(99)) or (inputs(232)));
    layer0_outputs(5740) <= not((inputs(78)) or (inputs(77)));
    layer0_outputs(5741) <= not(inputs(6));
    layer0_outputs(5742) <= (inputs(149)) or (inputs(7));
    layer0_outputs(5743) <= not(inputs(188));
    layer0_outputs(5744) <= not((inputs(177)) or (inputs(24)));
    layer0_outputs(5745) <= inputs(87);
    layer0_outputs(5746) <= '0';
    layer0_outputs(5747) <= (inputs(179)) xor (inputs(1));
    layer0_outputs(5748) <= not(inputs(74)) or (inputs(42));
    layer0_outputs(5749) <= inputs(101);
    layer0_outputs(5750) <= (inputs(116)) and not (inputs(172));
    layer0_outputs(5751) <= (inputs(232)) and not (inputs(219));
    layer0_outputs(5752) <= not((inputs(173)) xor (inputs(59)));
    layer0_outputs(5753) <= (inputs(199)) xor (inputs(134));
    layer0_outputs(5754) <= not(inputs(53)) or (inputs(15));
    layer0_outputs(5755) <= not(inputs(60));
    layer0_outputs(5756) <= not(inputs(51));
    layer0_outputs(5757) <= '1';
    layer0_outputs(5758) <= inputs(246);
    layer0_outputs(5759) <= not(inputs(188)) or (inputs(146));
    layer0_outputs(5760) <= (inputs(0)) or (inputs(127));
    layer0_outputs(5761) <= not((inputs(102)) or (inputs(155)));
    layer0_outputs(5762) <= not(inputs(101));
    layer0_outputs(5763) <= not(inputs(138)) or (inputs(21));
    layer0_outputs(5764) <= not((inputs(251)) xor (inputs(167)));
    layer0_outputs(5765) <= inputs(23);
    layer0_outputs(5766) <= not((inputs(144)) xor (inputs(39)));
    layer0_outputs(5767) <= inputs(113);
    layer0_outputs(5768) <= not((inputs(70)) or (inputs(213)));
    layer0_outputs(5769) <= (inputs(125)) or (inputs(90));
    layer0_outputs(5770) <= not((inputs(64)) xor (inputs(19)));
    layer0_outputs(5771) <= '1';
    layer0_outputs(5772) <= (inputs(114)) or (inputs(221));
    layer0_outputs(5773) <= not((inputs(125)) or (inputs(90)));
    layer0_outputs(5774) <= not(inputs(77)) or (inputs(1));
    layer0_outputs(5775) <= inputs(103);
    layer0_outputs(5776) <= not(inputs(149));
    layer0_outputs(5777) <= (inputs(122)) or (inputs(109));
    layer0_outputs(5778) <= (inputs(133)) xor (inputs(12));
    layer0_outputs(5779) <= not(inputs(85));
    layer0_outputs(5780) <= (inputs(27)) xor (inputs(156));
    layer0_outputs(5781) <= (inputs(203)) and not (inputs(22));
    layer0_outputs(5782) <= not(inputs(213));
    layer0_outputs(5783) <= (inputs(174)) xor (inputs(202));
    layer0_outputs(5784) <= '1';
    layer0_outputs(5785) <= (inputs(55)) xor (inputs(93));
    layer0_outputs(5786) <= not((inputs(234)) xor (inputs(43)));
    layer0_outputs(5787) <= (inputs(233)) xor (inputs(42));
    layer0_outputs(5788) <= not(inputs(24)) or (inputs(255));
    layer0_outputs(5789) <= (inputs(92)) and not (inputs(15));
    layer0_outputs(5790) <= not((inputs(175)) or (inputs(179)));
    layer0_outputs(5791) <= (inputs(137)) xor (inputs(242));
    layer0_outputs(5792) <= not(inputs(136)) or (inputs(131));
    layer0_outputs(5793) <= (inputs(101)) or (inputs(129));
    layer0_outputs(5794) <= (inputs(189)) or (inputs(202));
    layer0_outputs(5795) <= not((inputs(147)) or (inputs(125)));
    layer0_outputs(5796) <= not((inputs(251)) and (inputs(4)));
    layer0_outputs(5797) <= (inputs(250)) or (inputs(76));
    layer0_outputs(5798) <= not(inputs(14));
    layer0_outputs(5799) <= (inputs(245)) or (inputs(129));
    layer0_outputs(5800) <= (inputs(224)) xor (inputs(135));
    layer0_outputs(5801) <= not((inputs(151)) or (inputs(28)));
    layer0_outputs(5802) <= not((inputs(193)) and (inputs(198)));
    layer0_outputs(5803) <= not(inputs(143)) or (inputs(4));
    layer0_outputs(5804) <= not(inputs(94)) or (inputs(64));
    layer0_outputs(5805) <= not((inputs(30)) or (inputs(234)));
    layer0_outputs(5806) <= (inputs(217)) xor (inputs(88));
    layer0_outputs(5807) <= not(inputs(230)) or (inputs(49));
    layer0_outputs(5808) <= not((inputs(145)) xor (inputs(183)));
    layer0_outputs(5809) <= '1';
    layer0_outputs(5810) <= '1';
    layer0_outputs(5811) <= (inputs(252)) and not (inputs(3));
    layer0_outputs(5812) <= (inputs(65)) xor (inputs(217));
    layer0_outputs(5813) <= not((inputs(107)) or (inputs(211)));
    layer0_outputs(5814) <= inputs(19);
    layer0_outputs(5815) <= (inputs(208)) and not (inputs(187));
    layer0_outputs(5816) <= (inputs(242)) and not (inputs(207));
    layer0_outputs(5817) <= not((inputs(197)) xor (inputs(161)));
    layer0_outputs(5818) <= (inputs(116)) xor (inputs(1));
    layer0_outputs(5819) <= '1';
    layer0_outputs(5820) <= not(inputs(121));
    layer0_outputs(5821) <= inputs(153);
    layer0_outputs(5822) <= not(inputs(79));
    layer0_outputs(5823) <= inputs(99);
    layer0_outputs(5824) <= not((inputs(76)) xor (inputs(229)));
    layer0_outputs(5825) <= (inputs(159)) xor (inputs(134));
    layer0_outputs(5826) <= not((inputs(99)) or (inputs(209)));
    layer0_outputs(5827) <= (inputs(16)) or (inputs(213));
    layer0_outputs(5828) <= (inputs(156)) and not (inputs(184));
    layer0_outputs(5829) <= (inputs(191)) and not (inputs(207));
    layer0_outputs(5830) <= (inputs(254)) and not (inputs(83));
    layer0_outputs(5831) <= (inputs(233)) xor (inputs(164));
    layer0_outputs(5832) <= not(inputs(84));
    layer0_outputs(5833) <= not(inputs(52));
    layer0_outputs(5834) <= (inputs(193)) or (inputs(219));
    layer0_outputs(5835) <= not((inputs(146)) xor (inputs(158)));
    layer0_outputs(5836) <= inputs(147);
    layer0_outputs(5837) <= not((inputs(69)) xor (inputs(24)));
    layer0_outputs(5838) <= not(inputs(201)) or (inputs(8));
    layer0_outputs(5839) <= (inputs(162)) xor (inputs(189));
    layer0_outputs(5840) <= (inputs(134)) and not (inputs(190));
    layer0_outputs(5841) <= (inputs(79)) xor (inputs(6));
    layer0_outputs(5842) <= (inputs(21)) and not (inputs(223));
    layer0_outputs(5843) <= (inputs(23)) or (inputs(137));
    layer0_outputs(5844) <= inputs(189);
    layer0_outputs(5845) <= '0';
    layer0_outputs(5846) <= not((inputs(64)) or (inputs(209)));
    layer0_outputs(5847) <= not(inputs(11));
    layer0_outputs(5848) <= (inputs(215)) or (inputs(161));
    layer0_outputs(5849) <= not(inputs(167));
    layer0_outputs(5850) <= not(inputs(89));
    layer0_outputs(5851) <= not(inputs(201)) or (inputs(90));
    layer0_outputs(5852) <= (inputs(10)) and not (inputs(20));
    layer0_outputs(5853) <= (inputs(178)) or (inputs(71));
    layer0_outputs(5854) <= not((inputs(205)) and (inputs(224)));
    layer0_outputs(5855) <= (inputs(183)) xor (inputs(13));
    layer0_outputs(5856) <= not((inputs(27)) xor (inputs(87)));
    layer0_outputs(5857) <= (inputs(135)) xor (inputs(152));
    layer0_outputs(5858) <= not(inputs(147));
    layer0_outputs(5859) <= inputs(23);
    layer0_outputs(5860) <= (inputs(165)) and not (inputs(205));
    layer0_outputs(5861) <= inputs(189);
    layer0_outputs(5862) <= (inputs(172)) and not (inputs(210));
    layer0_outputs(5863) <= '1';
    layer0_outputs(5864) <= not(inputs(133));
    layer0_outputs(5865) <= not((inputs(239)) or (inputs(46)));
    layer0_outputs(5866) <= not((inputs(119)) or (inputs(143)));
    layer0_outputs(5867) <= not(inputs(218));
    layer0_outputs(5868) <= '1';
    layer0_outputs(5869) <= not(inputs(8));
    layer0_outputs(5870) <= not((inputs(222)) and (inputs(174)));
    layer0_outputs(5871) <= not(inputs(36)) or (inputs(143));
    layer0_outputs(5872) <= inputs(133);
    layer0_outputs(5873) <= not((inputs(210)) xor (inputs(38)));
    layer0_outputs(5874) <= not(inputs(118)) or (inputs(226));
    layer0_outputs(5875) <= not(inputs(57));
    layer0_outputs(5876) <= not((inputs(218)) or (inputs(111)));
    layer0_outputs(5877) <= (inputs(86)) xor (inputs(83));
    layer0_outputs(5878) <= not(inputs(154));
    layer0_outputs(5879) <= inputs(33);
    layer0_outputs(5880) <= inputs(196);
    layer0_outputs(5881) <= not((inputs(54)) or (inputs(106)));
    layer0_outputs(5882) <= not(inputs(121));
    layer0_outputs(5883) <= (inputs(171)) and not (inputs(161));
    layer0_outputs(5884) <= not((inputs(247)) xor (inputs(11)));
    layer0_outputs(5885) <= (inputs(216)) or (inputs(90));
    layer0_outputs(5886) <= not((inputs(204)) xor (inputs(0)));
    layer0_outputs(5887) <= not((inputs(21)) or (inputs(71)));
    layer0_outputs(5888) <= not(inputs(174));
    layer0_outputs(5889) <= '1';
    layer0_outputs(5890) <= not(inputs(132));
    layer0_outputs(5891) <= not((inputs(52)) and (inputs(32)));
    layer0_outputs(5892) <= (inputs(148)) xor (inputs(101));
    layer0_outputs(5893) <= (inputs(73)) xor (inputs(129));
    layer0_outputs(5894) <= (inputs(108)) and not (inputs(82));
    layer0_outputs(5895) <= (inputs(14)) or (inputs(234));
    layer0_outputs(5896) <= not((inputs(193)) xor (inputs(157)));
    layer0_outputs(5897) <= not((inputs(134)) or (inputs(69)));
    layer0_outputs(5898) <= not(inputs(41));
    layer0_outputs(5899) <= (inputs(126)) and (inputs(8));
    layer0_outputs(5900) <= (inputs(91)) or (inputs(15));
    layer0_outputs(5901) <= not(inputs(199)) or (inputs(52));
    layer0_outputs(5902) <= (inputs(136)) or (inputs(255));
    layer0_outputs(5903) <= not((inputs(207)) xor (inputs(35)));
    layer0_outputs(5904) <= (inputs(198)) or (inputs(194));
    layer0_outputs(5905) <= (inputs(134)) or (inputs(251));
    layer0_outputs(5906) <= not(inputs(155)) or (inputs(51));
    layer0_outputs(5907) <= (inputs(162)) or (inputs(132));
    layer0_outputs(5908) <= (inputs(124)) or (inputs(199));
    layer0_outputs(5909) <= (inputs(201)) xor (inputs(3));
    layer0_outputs(5910) <= not((inputs(86)) and (inputs(121)));
    layer0_outputs(5911) <= (inputs(98)) xor (inputs(87));
    layer0_outputs(5912) <= inputs(122);
    layer0_outputs(5913) <= (inputs(6)) or (inputs(109));
    layer0_outputs(5914) <= not(inputs(218)) or (inputs(240));
    layer0_outputs(5915) <= not((inputs(19)) xor (inputs(132)));
    layer0_outputs(5916) <= (inputs(233)) and not (inputs(3));
    layer0_outputs(5917) <= not(inputs(219));
    layer0_outputs(5918) <= not((inputs(55)) xor (inputs(85)));
    layer0_outputs(5919) <= not(inputs(95));
    layer0_outputs(5920) <= (inputs(107)) and not (inputs(210));
    layer0_outputs(5921) <= not(inputs(101)) or (inputs(133));
    layer0_outputs(5922) <= inputs(72);
    layer0_outputs(5923) <= not((inputs(133)) xor (inputs(0)));
    layer0_outputs(5924) <= not(inputs(182)) or (inputs(54));
    layer0_outputs(5925) <= not((inputs(109)) xor (inputs(71)));
    layer0_outputs(5926) <= inputs(82);
    layer0_outputs(5927) <= not(inputs(214));
    layer0_outputs(5928) <= not((inputs(148)) or (inputs(6)));
    layer0_outputs(5929) <= '0';
    layer0_outputs(5930) <= inputs(150);
    layer0_outputs(5931) <= inputs(137);
    layer0_outputs(5932) <= not((inputs(219)) xor (inputs(217)));
    layer0_outputs(5933) <= inputs(28);
    layer0_outputs(5934) <= inputs(75);
    layer0_outputs(5935) <= (inputs(229)) or (inputs(220));
    layer0_outputs(5936) <= '0';
    layer0_outputs(5937) <= not(inputs(116));
    layer0_outputs(5938) <= not(inputs(76));
    layer0_outputs(5939) <= (inputs(39)) xor (inputs(26));
    layer0_outputs(5940) <= not((inputs(123)) and (inputs(75)));
    layer0_outputs(5941) <= not((inputs(238)) or (inputs(77)));
    layer0_outputs(5942) <= not(inputs(88));
    layer0_outputs(5943) <= not(inputs(48));
    layer0_outputs(5944) <= '0';
    layer0_outputs(5945) <= not((inputs(224)) or (inputs(173)));
    layer0_outputs(5946) <= inputs(192);
    layer0_outputs(5947) <= (inputs(233)) or (inputs(148));
    layer0_outputs(5948) <= not((inputs(48)) or (inputs(124)));
    layer0_outputs(5949) <= inputs(218);
    layer0_outputs(5950) <= not(inputs(123));
    layer0_outputs(5951) <= (inputs(110)) and not (inputs(203));
    layer0_outputs(5952) <= (inputs(78)) and not (inputs(244));
    layer0_outputs(5953) <= inputs(34);
    layer0_outputs(5954) <= not((inputs(169)) or (inputs(172)));
    layer0_outputs(5955) <= inputs(215);
    layer0_outputs(5956) <= not(inputs(102));
    layer0_outputs(5957) <= not((inputs(252)) or (inputs(94)));
    layer0_outputs(5958) <= (inputs(56)) or (inputs(218));
    layer0_outputs(5959) <= '0';
    layer0_outputs(5960) <= not((inputs(212)) or (inputs(175)));
    layer0_outputs(5961) <= not(inputs(48)) or (inputs(203));
    layer0_outputs(5962) <= not((inputs(91)) or (inputs(47)));
    layer0_outputs(5963) <= (inputs(29)) and not (inputs(65));
    layer0_outputs(5964) <= not(inputs(20));
    layer0_outputs(5965) <= not((inputs(21)) or (inputs(54)));
    layer0_outputs(5966) <= not((inputs(17)) and (inputs(31)));
    layer0_outputs(5967) <= not((inputs(105)) xor (inputs(112)));
    layer0_outputs(5968) <= (inputs(133)) and not (inputs(179));
    layer0_outputs(5969) <= not((inputs(182)) or (inputs(94)));
    layer0_outputs(5970) <= (inputs(27)) or (inputs(119));
    layer0_outputs(5971) <= (inputs(203)) and (inputs(251));
    layer0_outputs(5972) <= '1';
    layer0_outputs(5973) <= '1';
    layer0_outputs(5974) <= not(inputs(144)) or (inputs(80));
    layer0_outputs(5975) <= (inputs(132)) and not (inputs(227));
    layer0_outputs(5976) <= (inputs(126)) or (inputs(87));
    layer0_outputs(5977) <= (inputs(151)) xor (inputs(238));
    layer0_outputs(5978) <= inputs(55);
    layer0_outputs(5979) <= not((inputs(228)) or (inputs(78)));
    layer0_outputs(5980) <= not((inputs(196)) or (inputs(223)));
    layer0_outputs(5981) <= not(inputs(210));
    layer0_outputs(5982) <= not(inputs(190)) or (inputs(5));
    layer0_outputs(5983) <= '0';
    layer0_outputs(5984) <= not((inputs(178)) or (inputs(242)));
    layer0_outputs(5985) <= (inputs(171)) and not (inputs(128));
    layer0_outputs(5986) <= (inputs(78)) xor (inputs(57));
    layer0_outputs(5987) <= not((inputs(254)) xor (inputs(232)));
    layer0_outputs(5988) <= not(inputs(114)) or (inputs(254));
    layer0_outputs(5989) <= not(inputs(168)) or (inputs(26));
    layer0_outputs(5990) <= not(inputs(229));
    layer0_outputs(5991) <= (inputs(8)) or (inputs(110));
    layer0_outputs(5992) <= (inputs(185)) and (inputs(86));
    layer0_outputs(5993) <= (inputs(150)) or (inputs(25));
    layer0_outputs(5994) <= not((inputs(207)) xor (inputs(108)));
    layer0_outputs(5995) <= not((inputs(10)) or (inputs(141)));
    layer0_outputs(5996) <= not(inputs(118)) or (inputs(93));
    layer0_outputs(5997) <= not((inputs(166)) xor (inputs(104)));
    layer0_outputs(5998) <= '0';
    layer0_outputs(5999) <= not(inputs(145)) or (inputs(55));
    layer0_outputs(6000) <= inputs(17);
    layer0_outputs(6001) <= (inputs(241)) xor (inputs(62));
    layer0_outputs(6002) <= (inputs(109)) and not (inputs(12));
    layer0_outputs(6003) <= inputs(107);
    layer0_outputs(6004) <= (inputs(124)) or (inputs(125));
    layer0_outputs(6005) <= (inputs(166)) or (inputs(29));
    layer0_outputs(6006) <= inputs(107);
    layer0_outputs(6007) <= (inputs(60)) or (inputs(175));
    layer0_outputs(6008) <= not((inputs(109)) xor (inputs(171)));
    layer0_outputs(6009) <= not((inputs(80)) xor (inputs(130)));
    layer0_outputs(6010) <= not((inputs(246)) or (inputs(132)));
    layer0_outputs(6011) <= (inputs(74)) and not (inputs(45));
    layer0_outputs(6012) <= not((inputs(233)) or (inputs(20)));
    layer0_outputs(6013) <= not(inputs(229));
    layer0_outputs(6014) <= (inputs(184)) or (inputs(98));
    layer0_outputs(6015) <= (inputs(57)) and not (inputs(255));
    layer0_outputs(6016) <= not((inputs(73)) or (inputs(188)));
    layer0_outputs(6017) <= (inputs(162)) or (inputs(250));
    layer0_outputs(6018) <= '0';
    layer0_outputs(6019) <= inputs(118);
    layer0_outputs(6020) <= (inputs(56)) or (inputs(78));
    layer0_outputs(6021) <= not((inputs(243)) xor (inputs(75)));
    layer0_outputs(6022) <= not((inputs(163)) xor (inputs(195)));
    layer0_outputs(6023) <= '1';
    layer0_outputs(6024) <= not((inputs(62)) and (inputs(158)));
    layer0_outputs(6025) <= not((inputs(173)) or (inputs(250)));
    layer0_outputs(6026) <= not((inputs(178)) xor (inputs(239)));
    layer0_outputs(6027) <= not(inputs(172)) or (inputs(251));
    layer0_outputs(6028) <= (inputs(33)) and (inputs(142));
    layer0_outputs(6029) <= (inputs(29)) xor (inputs(5));
    layer0_outputs(6030) <= not((inputs(114)) or (inputs(106)));
    layer0_outputs(6031) <= (inputs(233)) xor (inputs(75));
    layer0_outputs(6032) <= (inputs(221)) xor (inputs(189));
    layer0_outputs(6033) <= (inputs(60)) and not (inputs(9));
    layer0_outputs(6034) <= not(inputs(138));
    layer0_outputs(6035) <= (inputs(39)) or (inputs(39));
    layer0_outputs(6036) <= not(inputs(201));
    layer0_outputs(6037) <= '1';
    layer0_outputs(6038) <= (inputs(255)) and not (inputs(238));
    layer0_outputs(6039) <= not(inputs(180));
    layer0_outputs(6040) <= (inputs(73)) xor (inputs(114));
    layer0_outputs(6041) <= '1';
    layer0_outputs(6042) <= (inputs(180)) xor (inputs(134));
    layer0_outputs(6043) <= not(inputs(156)) or (inputs(254));
    layer0_outputs(6044) <= not((inputs(26)) xor (inputs(23)));
    layer0_outputs(6045) <= (inputs(247)) xor (inputs(170));
    layer0_outputs(6046) <= not((inputs(203)) xor (inputs(195)));
    layer0_outputs(6047) <= not((inputs(174)) xor (inputs(52)));
    layer0_outputs(6048) <= not(inputs(128)) or (inputs(15));
    layer0_outputs(6049) <= (inputs(47)) xor (inputs(146));
    layer0_outputs(6050) <= not(inputs(85)) or (inputs(163));
    layer0_outputs(6051) <= not(inputs(201));
    layer0_outputs(6052) <= (inputs(168)) and not (inputs(80));
    layer0_outputs(6053) <= not(inputs(183)) or (inputs(163));
    layer0_outputs(6054) <= (inputs(117)) and not (inputs(143));
    layer0_outputs(6055) <= '1';
    layer0_outputs(6056) <= not(inputs(61)) or (inputs(50));
    layer0_outputs(6057) <= not(inputs(186)) or (inputs(82));
    layer0_outputs(6058) <= inputs(216);
    layer0_outputs(6059) <= inputs(179);
    layer0_outputs(6060) <= not((inputs(100)) xor (inputs(37)));
    layer0_outputs(6061) <= '1';
    layer0_outputs(6062) <= not(inputs(158)) or (inputs(42));
    layer0_outputs(6063) <= (inputs(88)) and not (inputs(29));
    layer0_outputs(6064) <= not((inputs(119)) xor (inputs(35)));
    layer0_outputs(6065) <= (inputs(70)) xor (inputs(144));
    layer0_outputs(6066) <= not((inputs(116)) xor (inputs(4)));
    layer0_outputs(6067) <= (inputs(241)) or (inputs(90));
    layer0_outputs(6068) <= (inputs(43)) and not (inputs(19));
    layer0_outputs(6069) <= inputs(16);
    layer0_outputs(6070) <= inputs(241);
    layer0_outputs(6071) <= (inputs(170)) xor (inputs(233));
    layer0_outputs(6072) <= (inputs(110)) or (inputs(216));
    layer0_outputs(6073) <= '0';
    layer0_outputs(6074) <= (inputs(210)) xor (inputs(170));
    layer0_outputs(6075) <= inputs(24);
    layer0_outputs(6076) <= not(inputs(51));
    layer0_outputs(6077) <= not((inputs(87)) or (inputs(113)));
    layer0_outputs(6078) <= (inputs(200)) and not (inputs(196));
    layer0_outputs(6079) <= (inputs(85)) or (inputs(6));
    layer0_outputs(6080) <= not((inputs(6)) xor (inputs(160)));
    layer0_outputs(6081) <= not(inputs(245)) or (inputs(27));
    layer0_outputs(6082) <= not((inputs(172)) or (inputs(211)));
    layer0_outputs(6083) <= not(inputs(173));
    layer0_outputs(6084) <= (inputs(58)) and not (inputs(45));
    layer0_outputs(6085) <= not((inputs(68)) or (inputs(171)));
    layer0_outputs(6086) <= not((inputs(124)) and (inputs(61)));
    layer0_outputs(6087) <= inputs(196);
    layer0_outputs(6088) <= not((inputs(176)) xor (inputs(68)));
    layer0_outputs(6089) <= not((inputs(45)) xor (inputs(85)));
    layer0_outputs(6090) <= (inputs(170)) and not (inputs(77));
    layer0_outputs(6091) <= not((inputs(55)) or (inputs(53)));
    layer0_outputs(6092) <= (inputs(210)) or (inputs(142));
    layer0_outputs(6093) <= not((inputs(232)) or (inputs(75)));
    layer0_outputs(6094) <= not((inputs(62)) and (inputs(79)));
    layer0_outputs(6095) <= (inputs(115)) and not (inputs(127));
    layer0_outputs(6096) <= not(inputs(72));
    layer0_outputs(6097) <= not((inputs(115)) xor (inputs(192)));
    layer0_outputs(6098) <= not(inputs(55));
    layer0_outputs(6099) <= (inputs(238)) xor (inputs(104));
    layer0_outputs(6100) <= (inputs(132)) or (inputs(176));
    layer0_outputs(6101) <= inputs(187);
    layer0_outputs(6102) <= not((inputs(235)) or (inputs(188)));
    layer0_outputs(6103) <= (inputs(38)) and not (inputs(13));
    layer0_outputs(6104) <= '0';
    layer0_outputs(6105) <= (inputs(130)) and not (inputs(177));
    layer0_outputs(6106) <= (inputs(6)) xor (inputs(62));
    layer0_outputs(6107) <= '1';
    layer0_outputs(6108) <= (inputs(61)) or (inputs(49));
    layer0_outputs(6109) <= inputs(169);
    layer0_outputs(6110) <= inputs(104);
    layer0_outputs(6111) <= not(inputs(66));
    layer0_outputs(6112) <= (inputs(78)) and (inputs(227));
    layer0_outputs(6113) <= not((inputs(239)) xor (inputs(4)));
    layer0_outputs(6114) <= inputs(202);
    layer0_outputs(6115) <= not((inputs(38)) and (inputs(82)));
    layer0_outputs(6116) <= not((inputs(188)) or (inputs(50)));
    layer0_outputs(6117) <= not((inputs(233)) or (inputs(245)));
    layer0_outputs(6118) <= not((inputs(228)) and (inputs(238)));
    layer0_outputs(6119) <= not((inputs(98)) or (inputs(29)));
    layer0_outputs(6120) <= (inputs(95)) xor (inputs(90));
    layer0_outputs(6121) <= not(inputs(181)) or (inputs(28));
    layer0_outputs(6122) <= inputs(46);
    layer0_outputs(6123) <= (inputs(154)) and not (inputs(44));
    layer0_outputs(6124) <= inputs(30);
    layer0_outputs(6125) <= (inputs(93)) and not (inputs(9));
    layer0_outputs(6126) <= inputs(22);
    layer0_outputs(6127) <= not(inputs(31));
    layer0_outputs(6128) <= (inputs(28)) and (inputs(26));
    layer0_outputs(6129) <= (inputs(186)) xor (inputs(30));
    layer0_outputs(6130) <= not(inputs(122));
    layer0_outputs(6131) <= inputs(57);
    layer0_outputs(6132) <= (inputs(123)) and not (inputs(36));
    layer0_outputs(6133) <= inputs(55);
    layer0_outputs(6134) <= not((inputs(2)) xor (inputs(59)));
    layer0_outputs(6135) <= not(inputs(149)) or (inputs(130));
    layer0_outputs(6136) <= (inputs(145)) or (inputs(150));
    layer0_outputs(6137) <= (inputs(232)) or (inputs(212));
    layer0_outputs(6138) <= (inputs(149)) xor (inputs(242));
    layer0_outputs(6139) <= (inputs(49)) or (inputs(180));
    layer0_outputs(6140) <= not(inputs(198)) or (inputs(94));
    layer0_outputs(6141) <= (inputs(118)) or (inputs(119));
    layer0_outputs(6142) <= (inputs(21)) and not (inputs(98));
    layer0_outputs(6143) <= '0';
    layer0_outputs(6144) <= (inputs(207)) and (inputs(93));
    layer0_outputs(6145) <= not(inputs(143)) or (inputs(17));
    layer0_outputs(6146) <= not(inputs(105)) or (inputs(94));
    layer0_outputs(6147) <= (inputs(62)) xor (inputs(195));
    layer0_outputs(6148) <= not((inputs(99)) and (inputs(241)));
    layer0_outputs(6149) <= (inputs(121)) and not (inputs(177));
    layer0_outputs(6150) <= not((inputs(219)) or (inputs(152)));
    layer0_outputs(6151) <= (inputs(215)) and not (inputs(16));
    layer0_outputs(6152) <= inputs(93);
    layer0_outputs(6153) <= (inputs(23)) and (inputs(190));
    layer0_outputs(6154) <= not(inputs(69));
    layer0_outputs(6155) <= inputs(224);
    layer0_outputs(6156) <= '0';
    layer0_outputs(6157) <= inputs(124);
    layer0_outputs(6158) <= inputs(115);
    layer0_outputs(6159) <= inputs(91);
    layer0_outputs(6160) <= not((inputs(82)) xor (inputs(158)));
    layer0_outputs(6161) <= (inputs(85)) xor (inputs(147));
    layer0_outputs(6162) <= not(inputs(20)) or (inputs(49));
    layer0_outputs(6163) <= not((inputs(41)) xor (inputs(165)));
    layer0_outputs(6164) <= (inputs(195)) and not (inputs(30));
    layer0_outputs(6165) <= '1';
    layer0_outputs(6166) <= not(inputs(183)) or (inputs(172));
    layer0_outputs(6167) <= not(inputs(60)) or (inputs(1));
    layer0_outputs(6168) <= (inputs(100)) or (inputs(106));
    layer0_outputs(6169) <= (inputs(103)) and not (inputs(6));
    layer0_outputs(6170) <= (inputs(32)) xor (inputs(185));
    layer0_outputs(6171) <= (inputs(204)) and not (inputs(131));
    layer0_outputs(6172) <= (inputs(66)) and not (inputs(224));
    layer0_outputs(6173) <= inputs(218);
    layer0_outputs(6174) <= inputs(18);
    layer0_outputs(6175) <= not((inputs(170)) xor (inputs(181)));
    layer0_outputs(6176) <= (inputs(126)) and not (inputs(27));
    layer0_outputs(6177) <= (inputs(116)) or (inputs(52));
    layer0_outputs(6178) <= (inputs(182)) xor (inputs(212));
    layer0_outputs(6179) <= '0';
    layer0_outputs(6180) <= (inputs(120)) and not (inputs(39));
    layer0_outputs(6181) <= '0';
    layer0_outputs(6182) <= not(inputs(151)) or (inputs(208));
    layer0_outputs(6183) <= (inputs(55)) or (inputs(242));
    layer0_outputs(6184) <= inputs(232);
    layer0_outputs(6185) <= inputs(148);
    layer0_outputs(6186) <= (inputs(67)) xor (inputs(2));
    layer0_outputs(6187) <= (inputs(113)) xor (inputs(216));
    layer0_outputs(6188) <= inputs(213);
    layer0_outputs(6189) <= inputs(3);
    layer0_outputs(6190) <= not(inputs(106)) or (inputs(95));
    layer0_outputs(6191) <= (inputs(183)) and not (inputs(216));
    layer0_outputs(6192) <= (inputs(154)) xor (inputs(203));
    layer0_outputs(6193) <= not(inputs(0));
    layer0_outputs(6194) <= not((inputs(96)) or (inputs(110)));
    layer0_outputs(6195) <= (inputs(81)) and (inputs(12));
    layer0_outputs(6196) <= inputs(124);
    layer0_outputs(6197) <= not(inputs(69));
    layer0_outputs(6198) <= inputs(181);
    layer0_outputs(6199) <= (inputs(254)) or (inputs(143));
    layer0_outputs(6200) <= not(inputs(121));
    layer0_outputs(6201) <= (inputs(164)) and (inputs(3));
    layer0_outputs(6202) <= not(inputs(181)) or (inputs(203));
    layer0_outputs(6203) <= (inputs(227)) and not (inputs(83));
    layer0_outputs(6204) <= (inputs(133)) or (inputs(148));
    layer0_outputs(6205) <= not(inputs(111));
    layer0_outputs(6206) <= not((inputs(181)) xor (inputs(183)));
    layer0_outputs(6207) <= (inputs(72)) and not (inputs(52));
    layer0_outputs(6208) <= (inputs(95)) or (inputs(187));
    layer0_outputs(6209) <= inputs(155);
    layer0_outputs(6210) <= (inputs(165)) and not (inputs(235));
    layer0_outputs(6211) <= not((inputs(86)) or (inputs(29)));
    layer0_outputs(6212) <= inputs(159);
    layer0_outputs(6213) <= not((inputs(255)) or (inputs(161)));
    layer0_outputs(6214) <= not((inputs(148)) or (inputs(145)));
    layer0_outputs(6215) <= (inputs(86)) and not (inputs(12));
    layer0_outputs(6216) <= not(inputs(123));
    layer0_outputs(6217) <= (inputs(36)) xor (inputs(62));
    layer0_outputs(6218) <= (inputs(54)) or (inputs(88));
    layer0_outputs(6219) <= (inputs(19)) xor (inputs(109));
    layer0_outputs(6220) <= (inputs(63)) xor (inputs(140));
    layer0_outputs(6221) <= (inputs(181)) and not (inputs(194));
    layer0_outputs(6222) <= not((inputs(6)) or (inputs(35)));
    layer0_outputs(6223) <= (inputs(218)) or (inputs(187));
    layer0_outputs(6224) <= (inputs(0)) or (inputs(1));
    layer0_outputs(6225) <= '1';
    layer0_outputs(6226) <= not((inputs(156)) or (inputs(105)));
    layer0_outputs(6227) <= not((inputs(199)) xor (inputs(95)));
    layer0_outputs(6228) <= not(inputs(89)) or (inputs(255));
    layer0_outputs(6229) <= not((inputs(185)) or (inputs(211)));
    layer0_outputs(6230) <= not(inputs(220));
    layer0_outputs(6231) <= (inputs(26)) or (inputs(27));
    layer0_outputs(6232) <= not((inputs(114)) xor (inputs(242)));
    layer0_outputs(6233) <= not((inputs(71)) xor (inputs(87)));
    layer0_outputs(6234) <= '0';
    layer0_outputs(6235) <= (inputs(169)) or (inputs(241));
    layer0_outputs(6236) <= '0';
    layer0_outputs(6237) <= not((inputs(227)) or (inputs(156)));
    layer0_outputs(6238) <= (inputs(169)) and not (inputs(247));
    layer0_outputs(6239) <= not((inputs(203)) or (inputs(37)));
    layer0_outputs(6240) <= not(inputs(141)) or (inputs(14));
    layer0_outputs(6241) <= not(inputs(35));
    layer0_outputs(6242) <= not(inputs(120)) or (inputs(117));
    layer0_outputs(6243) <= (inputs(202)) xor (inputs(124));
    layer0_outputs(6244) <= (inputs(139)) xor (inputs(187));
    layer0_outputs(6245) <= not((inputs(47)) xor (inputs(166)));
    layer0_outputs(6246) <= (inputs(168)) xor (inputs(137));
    layer0_outputs(6247) <= (inputs(247)) and not (inputs(128));
    layer0_outputs(6248) <= not((inputs(71)) or (inputs(33)));
    layer0_outputs(6249) <= not(inputs(109)) or (inputs(201));
    layer0_outputs(6250) <= inputs(221);
    layer0_outputs(6251) <= (inputs(128)) xor (inputs(212));
    layer0_outputs(6252) <= not((inputs(30)) or (inputs(39)));
    layer0_outputs(6253) <= inputs(67);
    layer0_outputs(6254) <= (inputs(197)) and not (inputs(114));
    layer0_outputs(6255) <= (inputs(141)) xor (inputs(26));
    layer0_outputs(6256) <= not((inputs(170)) or (inputs(227)));
    layer0_outputs(6257) <= not(inputs(84));
    layer0_outputs(6258) <= not(inputs(173)) or (inputs(10));
    layer0_outputs(6259) <= not(inputs(6)) or (inputs(255));
    layer0_outputs(6260) <= not(inputs(42)) or (inputs(130));
    layer0_outputs(6261) <= not((inputs(103)) xor (inputs(231)));
    layer0_outputs(6262) <= not(inputs(137));
    layer0_outputs(6263) <= (inputs(254)) xor (inputs(60));
    layer0_outputs(6264) <= not((inputs(203)) xor (inputs(118)));
    layer0_outputs(6265) <= inputs(14);
    layer0_outputs(6266) <= not((inputs(197)) or (inputs(203)));
    layer0_outputs(6267) <= (inputs(21)) or (inputs(242));
    layer0_outputs(6268) <= not(inputs(76)) or (inputs(223));
    layer0_outputs(6269) <= inputs(120);
    layer0_outputs(6270) <= '0';
    layer0_outputs(6271) <= not(inputs(48)) or (inputs(26));
    layer0_outputs(6272) <= not(inputs(113));
    layer0_outputs(6273) <= inputs(111);
    layer0_outputs(6274) <= not(inputs(228));
    layer0_outputs(6275) <= '1';
    layer0_outputs(6276) <= not((inputs(61)) and (inputs(73)));
    layer0_outputs(6277) <= (inputs(121)) and not (inputs(6));
    layer0_outputs(6278) <= (inputs(199)) and not (inputs(168));
    layer0_outputs(6279) <= (inputs(229)) xor (inputs(176));
    layer0_outputs(6280) <= not((inputs(118)) or (inputs(104)));
    layer0_outputs(6281) <= not((inputs(150)) or (inputs(121)));
    layer0_outputs(6282) <= not(inputs(31)) or (inputs(164));
    layer0_outputs(6283) <= (inputs(214)) and not (inputs(124));
    layer0_outputs(6284) <= (inputs(48)) or (inputs(193));
    layer0_outputs(6285) <= not(inputs(126)) or (inputs(112));
    layer0_outputs(6286) <= (inputs(218)) xor (inputs(69));
    layer0_outputs(6287) <= inputs(97);
    layer0_outputs(6288) <= (inputs(223)) xor (inputs(109));
    layer0_outputs(6289) <= '1';
    layer0_outputs(6290) <= inputs(87);
    layer0_outputs(6291) <= not((inputs(194)) xor (inputs(228)));
    layer0_outputs(6292) <= inputs(33);
    layer0_outputs(6293) <= inputs(16);
    layer0_outputs(6294) <= inputs(12);
    layer0_outputs(6295) <= (inputs(218)) xor (inputs(122));
    layer0_outputs(6296) <= inputs(180);
    layer0_outputs(6297) <= not(inputs(203)) or (inputs(100));
    layer0_outputs(6298) <= (inputs(159)) xor (inputs(198));
    layer0_outputs(6299) <= (inputs(72)) and not (inputs(50));
    layer0_outputs(6300) <= (inputs(103)) xor (inputs(189));
    layer0_outputs(6301) <= (inputs(184)) xor (inputs(136));
    layer0_outputs(6302) <= (inputs(60)) and not (inputs(29));
    layer0_outputs(6303) <= not(inputs(22));
    layer0_outputs(6304) <= (inputs(36)) or (inputs(168));
    layer0_outputs(6305) <= (inputs(1)) or (inputs(56));
    layer0_outputs(6306) <= not((inputs(82)) or (inputs(211)));
    layer0_outputs(6307) <= inputs(129);
    layer0_outputs(6308) <= not(inputs(56)) or (inputs(149));
    layer0_outputs(6309) <= not(inputs(134)) or (inputs(65));
    layer0_outputs(6310) <= (inputs(242)) and not (inputs(7));
    layer0_outputs(6311) <= (inputs(18)) and not (inputs(35));
    layer0_outputs(6312) <= inputs(57);
    layer0_outputs(6313) <= (inputs(100)) xor (inputs(102));
    layer0_outputs(6314) <= (inputs(14)) or (inputs(247));
    layer0_outputs(6315) <= (inputs(147)) xor (inputs(231));
    layer0_outputs(6316) <= not(inputs(17));
    layer0_outputs(6317) <= (inputs(94)) and not (inputs(22));
    layer0_outputs(6318) <= inputs(131);
    layer0_outputs(6319) <= not((inputs(239)) xor (inputs(84)));
    layer0_outputs(6320) <= not((inputs(60)) xor (inputs(41)));
    layer0_outputs(6321) <= (inputs(40)) xor (inputs(122));
    layer0_outputs(6322) <= not(inputs(25));
    layer0_outputs(6323) <= (inputs(151)) and not (inputs(148));
    layer0_outputs(6324) <= (inputs(133)) and not (inputs(197));
    layer0_outputs(6325) <= (inputs(86)) or (inputs(102));
    layer0_outputs(6326) <= not((inputs(100)) or (inputs(115)));
    layer0_outputs(6327) <= (inputs(219)) and not (inputs(96));
    layer0_outputs(6328) <= (inputs(105)) xor (inputs(76));
    layer0_outputs(6329) <= (inputs(203)) xor (inputs(69));
    layer0_outputs(6330) <= not((inputs(59)) or (inputs(3)));
    layer0_outputs(6331) <= not((inputs(64)) and (inputs(7)));
    layer0_outputs(6332) <= inputs(66);
    layer0_outputs(6333) <= not((inputs(14)) xor (inputs(169)));
    layer0_outputs(6334) <= (inputs(52)) and not (inputs(93));
    layer0_outputs(6335) <= inputs(101);
    layer0_outputs(6336) <= not((inputs(173)) or (inputs(58)));
    layer0_outputs(6337) <= inputs(231);
    layer0_outputs(6338) <= (inputs(34)) and (inputs(1));
    layer0_outputs(6339) <= (inputs(219)) xor (inputs(189));
    layer0_outputs(6340) <= '0';
    layer0_outputs(6341) <= inputs(217);
    layer0_outputs(6342) <= not(inputs(36));
    layer0_outputs(6343) <= (inputs(187)) or (inputs(78));
    layer0_outputs(6344) <= inputs(93);
    layer0_outputs(6345) <= (inputs(51)) and not (inputs(109));
    layer0_outputs(6346) <= not(inputs(171));
    layer0_outputs(6347) <= not(inputs(153)) or (inputs(167));
    layer0_outputs(6348) <= not(inputs(243));
    layer0_outputs(6349) <= (inputs(249)) and (inputs(2));
    layer0_outputs(6350) <= (inputs(171)) and not (inputs(236));
    layer0_outputs(6351) <= inputs(254);
    layer0_outputs(6352) <= inputs(131);
    layer0_outputs(6353) <= not(inputs(115)) or (inputs(81));
    layer0_outputs(6354) <= not((inputs(107)) or (inputs(165)));
    layer0_outputs(6355) <= inputs(157);
    layer0_outputs(6356) <= '1';
    layer0_outputs(6357) <= not((inputs(178)) or (inputs(236)));
    layer0_outputs(6358) <= not((inputs(175)) or (inputs(82)));
    layer0_outputs(6359) <= not(inputs(188));
    layer0_outputs(6360) <= inputs(239);
    layer0_outputs(6361) <= (inputs(91)) and (inputs(224));
    layer0_outputs(6362) <= (inputs(61)) or (inputs(99));
    layer0_outputs(6363) <= not(inputs(186)) or (inputs(26));
    layer0_outputs(6364) <= (inputs(231)) and (inputs(17));
    layer0_outputs(6365) <= inputs(225);
    layer0_outputs(6366) <= (inputs(202)) and not (inputs(148));
    layer0_outputs(6367) <= not((inputs(168)) and (inputs(91)));
    layer0_outputs(6368) <= not((inputs(129)) or (inputs(239)));
    layer0_outputs(6369) <= (inputs(248)) or (inputs(85));
    layer0_outputs(6370) <= not(inputs(137));
    layer0_outputs(6371) <= not((inputs(72)) xor (inputs(146)));
    layer0_outputs(6372) <= (inputs(210)) or (inputs(181));
    layer0_outputs(6373) <= (inputs(153)) xor (inputs(243));
    layer0_outputs(6374) <= inputs(63);
    layer0_outputs(6375) <= (inputs(133)) or (inputs(31));
    layer0_outputs(6376) <= inputs(107);
    layer0_outputs(6377) <= not(inputs(181));
    layer0_outputs(6378) <= (inputs(111)) and not (inputs(37));
    layer0_outputs(6379) <= not((inputs(0)) xor (inputs(224)));
    layer0_outputs(6380) <= (inputs(36)) and not (inputs(197));
    layer0_outputs(6381) <= (inputs(178)) or (inputs(63));
    layer0_outputs(6382) <= (inputs(196)) or (inputs(179));
    layer0_outputs(6383) <= not((inputs(107)) and (inputs(232)));
    layer0_outputs(6384) <= not(inputs(102));
    layer0_outputs(6385) <= (inputs(101)) and not (inputs(65));
    layer0_outputs(6386) <= (inputs(195)) or (inputs(180));
    layer0_outputs(6387) <= (inputs(174)) or (inputs(12));
    layer0_outputs(6388) <= (inputs(117)) and not (inputs(107));
    layer0_outputs(6389) <= inputs(181);
    layer0_outputs(6390) <= inputs(153);
    layer0_outputs(6391) <= (inputs(169)) and not (inputs(81));
    layer0_outputs(6392) <= (inputs(174)) and not (inputs(208));
    layer0_outputs(6393) <= not(inputs(161));
    layer0_outputs(6394) <= (inputs(133)) or (inputs(78));
    layer0_outputs(6395) <= inputs(64);
    layer0_outputs(6396) <= '0';
    layer0_outputs(6397) <= not(inputs(233)) or (inputs(180));
    layer0_outputs(6398) <= (inputs(144)) or (inputs(217));
    layer0_outputs(6399) <= (inputs(39)) or (inputs(26));
    layer0_outputs(6400) <= (inputs(250)) and (inputs(189));
    layer0_outputs(6401) <= not(inputs(109)) or (inputs(94));
    layer0_outputs(6402) <= not(inputs(72));
    layer0_outputs(6403) <= not((inputs(59)) and (inputs(76)));
    layer0_outputs(6404) <= inputs(252);
    layer0_outputs(6405) <= '0';
    layer0_outputs(6406) <= not(inputs(236));
    layer0_outputs(6407) <= (inputs(79)) xor (inputs(160));
    layer0_outputs(6408) <= (inputs(133)) xor (inputs(98));
    layer0_outputs(6409) <= '1';
    layer0_outputs(6410) <= '0';
    layer0_outputs(6411) <= not((inputs(224)) or (inputs(218)));
    layer0_outputs(6412) <= (inputs(231)) xor (inputs(29));
    layer0_outputs(6413) <= (inputs(12)) and not (inputs(145));
    layer0_outputs(6414) <= not(inputs(153));
    layer0_outputs(6415) <= not((inputs(29)) xor (inputs(125)));
    layer0_outputs(6416) <= (inputs(83)) and not (inputs(190));
    layer0_outputs(6417) <= not((inputs(231)) or (inputs(186)));
    layer0_outputs(6418) <= not(inputs(134));
    layer0_outputs(6419) <= '1';
    layer0_outputs(6420) <= (inputs(222)) and not (inputs(89));
    layer0_outputs(6421) <= not((inputs(11)) or (inputs(117)));
    layer0_outputs(6422) <= (inputs(162)) xor (inputs(199));
    layer0_outputs(6423) <= not(inputs(238));
    layer0_outputs(6424) <= (inputs(138)) xor (inputs(172));
    layer0_outputs(6425) <= not(inputs(6));
    layer0_outputs(6426) <= inputs(238);
    layer0_outputs(6427) <= (inputs(4)) and not (inputs(0));
    layer0_outputs(6428) <= inputs(150);
    layer0_outputs(6429) <= '1';
    layer0_outputs(6430) <= inputs(61);
    layer0_outputs(6431) <= '0';
    layer0_outputs(6432) <= not(inputs(18));
    layer0_outputs(6433) <= not((inputs(179)) or (inputs(74)));
    layer0_outputs(6434) <= (inputs(217)) or (inputs(190));
    layer0_outputs(6435) <= not((inputs(169)) xor (inputs(171)));
    layer0_outputs(6436) <= '1';
    layer0_outputs(6437) <= not((inputs(44)) xor (inputs(116)));
    layer0_outputs(6438) <= (inputs(7)) xor (inputs(40));
    layer0_outputs(6439) <= not(inputs(132));
    layer0_outputs(6440) <= not((inputs(61)) or (inputs(83)));
    layer0_outputs(6441) <= not((inputs(223)) xor (inputs(15)));
    layer0_outputs(6442) <= (inputs(52)) xor (inputs(56));
    layer0_outputs(6443) <= not(inputs(216));
    layer0_outputs(6444) <= inputs(232);
    layer0_outputs(6445) <= not(inputs(134));
    layer0_outputs(6446) <= inputs(103);
    layer0_outputs(6447) <= inputs(200);
    layer0_outputs(6448) <= '1';
    layer0_outputs(6449) <= (inputs(96)) or (inputs(30));
    layer0_outputs(6450) <= (inputs(189)) xor (inputs(95));
    layer0_outputs(6451) <= (inputs(120)) xor (inputs(142));
    layer0_outputs(6452) <= not(inputs(122)) or (inputs(50));
    layer0_outputs(6453) <= not(inputs(199));
    layer0_outputs(6454) <= not(inputs(86));
    layer0_outputs(6455) <= (inputs(95)) and not (inputs(241));
    layer0_outputs(6456) <= (inputs(239)) and not (inputs(12));
    layer0_outputs(6457) <= not((inputs(170)) or (inputs(236)));
    layer0_outputs(6458) <= not((inputs(168)) xor (inputs(147)));
    layer0_outputs(6459) <= (inputs(66)) xor (inputs(4));
    layer0_outputs(6460) <= not((inputs(47)) xor (inputs(142)));
    layer0_outputs(6461) <= not(inputs(217)) or (inputs(147));
    layer0_outputs(6462) <= inputs(173);
    layer0_outputs(6463) <= not((inputs(235)) or (inputs(190)));
    layer0_outputs(6464) <= (inputs(171)) xor (inputs(95));
    layer0_outputs(6465) <= not(inputs(115));
    layer0_outputs(6466) <= not(inputs(194)) or (inputs(91));
    layer0_outputs(6467) <= inputs(243);
    layer0_outputs(6468) <= not((inputs(22)) and (inputs(174)));
    layer0_outputs(6469) <= inputs(214);
    layer0_outputs(6470) <= (inputs(235)) or (inputs(98));
    layer0_outputs(6471) <= inputs(152);
    layer0_outputs(6472) <= (inputs(40)) or (inputs(185));
    layer0_outputs(6473) <= (inputs(218)) and (inputs(198));
    layer0_outputs(6474) <= not(inputs(19));
    layer0_outputs(6475) <= (inputs(137)) or (inputs(163));
    layer0_outputs(6476) <= not((inputs(31)) xor (inputs(85)));
    layer0_outputs(6477) <= (inputs(181)) xor (inputs(43));
    layer0_outputs(6478) <= (inputs(12)) and (inputs(254));
    layer0_outputs(6479) <= not(inputs(250));
    layer0_outputs(6480) <= inputs(28);
    layer0_outputs(6481) <= not(inputs(25));
    layer0_outputs(6482) <= not(inputs(218)) or (inputs(244));
    layer0_outputs(6483) <= not(inputs(197));
    layer0_outputs(6484) <= not(inputs(210));
    layer0_outputs(6485) <= (inputs(235)) and not (inputs(129));
    layer0_outputs(6486) <= (inputs(74)) or (inputs(79));
    layer0_outputs(6487) <= not(inputs(122)) or (inputs(68));
    layer0_outputs(6488) <= not((inputs(144)) xor (inputs(228)));
    layer0_outputs(6489) <= (inputs(108)) and not (inputs(15));
    layer0_outputs(6490) <= not(inputs(95));
    layer0_outputs(6491) <= not(inputs(119));
    layer0_outputs(6492) <= not((inputs(253)) and (inputs(226)));
    layer0_outputs(6493) <= (inputs(132)) and not (inputs(43));
    layer0_outputs(6494) <= not(inputs(48));
    layer0_outputs(6495) <= (inputs(109)) or (inputs(8));
    layer0_outputs(6496) <= not(inputs(24));
    layer0_outputs(6497) <= (inputs(156)) and not (inputs(94));
    layer0_outputs(6498) <= (inputs(71)) xor (inputs(127));
    layer0_outputs(6499) <= not((inputs(96)) xor (inputs(195)));
    layer0_outputs(6500) <= (inputs(88)) xor (inputs(253));
    layer0_outputs(6501) <= (inputs(145)) or (inputs(60));
    layer0_outputs(6502) <= not(inputs(250));
    layer0_outputs(6503) <= (inputs(205)) xor (inputs(47));
    layer0_outputs(6504) <= not((inputs(125)) or (inputs(116)));
    layer0_outputs(6505) <= '0';
    layer0_outputs(6506) <= not(inputs(152)) or (inputs(102));
    layer0_outputs(6507) <= not(inputs(130));
    layer0_outputs(6508) <= (inputs(171)) and not (inputs(17));
    layer0_outputs(6509) <= not(inputs(34)) or (inputs(253));
    layer0_outputs(6510) <= not(inputs(59));
    layer0_outputs(6511) <= not((inputs(17)) xor (inputs(119)));
    layer0_outputs(6512) <= '0';
    layer0_outputs(6513) <= not((inputs(73)) xor (inputs(139)));
    layer0_outputs(6514) <= (inputs(34)) or (inputs(14));
    layer0_outputs(6515) <= (inputs(255)) or (inputs(129));
    layer0_outputs(6516) <= (inputs(74)) or (inputs(69));
    layer0_outputs(6517) <= not(inputs(117));
    layer0_outputs(6518) <= (inputs(208)) xor (inputs(35));
    layer0_outputs(6519) <= (inputs(62)) xor (inputs(121));
    layer0_outputs(6520) <= not(inputs(101)) or (inputs(140));
    layer0_outputs(6521) <= (inputs(81)) and not (inputs(147));
    layer0_outputs(6522) <= '0';
    layer0_outputs(6523) <= (inputs(154)) and not (inputs(65));
    layer0_outputs(6524) <= (inputs(83)) and not (inputs(19));
    layer0_outputs(6525) <= (inputs(105)) or (inputs(151));
    layer0_outputs(6526) <= (inputs(198)) xor (inputs(188));
    layer0_outputs(6527) <= (inputs(38)) and not (inputs(65));
    layer0_outputs(6528) <= '1';
    layer0_outputs(6529) <= (inputs(125)) xor (inputs(247));
    layer0_outputs(6530) <= (inputs(39)) or (inputs(89));
    layer0_outputs(6531) <= (inputs(208)) and not (inputs(116));
    layer0_outputs(6532) <= inputs(179);
    layer0_outputs(6533) <= not(inputs(90)) or (inputs(42));
    layer0_outputs(6534) <= '1';
    layer0_outputs(6535) <= (inputs(43)) and not (inputs(144));
    layer0_outputs(6536) <= not(inputs(240)) or (inputs(238));
    layer0_outputs(6537) <= not(inputs(50));
    layer0_outputs(6538) <= inputs(217);
    layer0_outputs(6539) <= (inputs(110)) or (inputs(15));
    layer0_outputs(6540) <= not(inputs(157));
    layer0_outputs(6541) <= (inputs(177)) xor (inputs(138));
    layer0_outputs(6542) <= not(inputs(202));
    layer0_outputs(6543) <= not(inputs(121)) or (inputs(92));
    layer0_outputs(6544) <= not((inputs(160)) or (inputs(228)));
    layer0_outputs(6545) <= not(inputs(248));
    layer0_outputs(6546) <= not(inputs(119));
    layer0_outputs(6547) <= inputs(126);
    layer0_outputs(6548) <= '1';
    layer0_outputs(6549) <= not(inputs(137));
    layer0_outputs(6550) <= not((inputs(236)) or (inputs(169)));
    layer0_outputs(6551) <= not((inputs(64)) xor (inputs(21)));
    layer0_outputs(6552) <= not(inputs(66));
    layer0_outputs(6553) <= not(inputs(129));
    layer0_outputs(6554) <= not(inputs(172));
    layer0_outputs(6555) <= not(inputs(135));
    layer0_outputs(6556) <= not(inputs(118));
    layer0_outputs(6557) <= (inputs(75)) xor (inputs(185));
    layer0_outputs(6558) <= not((inputs(157)) or (inputs(219)));
    layer0_outputs(6559) <= not(inputs(148));
    layer0_outputs(6560) <= inputs(180);
    layer0_outputs(6561) <= inputs(204);
    layer0_outputs(6562) <= '1';
    layer0_outputs(6563) <= not(inputs(200));
    layer0_outputs(6564) <= inputs(24);
    layer0_outputs(6565) <= not((inputs(111)) or (inputs(55)));
    layer0_outputs(6566) <= not(inputs(134)) or (inputs(83));
    layer0_outputs(6567) <= (inputs(83)) xor (inputs(160));
    layer0_outputs(6568) <= '1';
    layer0_outputs(6569) <= (inputs(158)) or (inputs(132));
    layer0_outputs(6570) <= not((inputs(206)) xor (inputs(196)));
    layer0_outputs(6571) <= inputs(106);
    layer0_outputs(6572) <= (inputs(255)) and (inputs(206));
    layer0_outputs(6573) <= (inputs(195)) xor (inputs(87));
    layer0_outputs(6574) <= (inputs(178)) or (inputs(17));
    layer0_outputs(6575) <= (inputs(71)) xor (inputs(180));
    layer0_outputs(6576) <= not((inputs(121)) or (inputs(63)));
    layer0_outputs(6577) <= (inputs(175)) xor (inputs(76));
    layer0_outputs(6578) <= (inputs(208)) xor (inputs(30));
    layer0_outputs(6579) <= (inputs(236)) or (inputs(215));
    layer0_outputs(6580) <= not((inputs(145)) or (inputs(32)));
    layer0_outputs(6581) <= not(inputs(228)) or (inputs(80));
    layer0_outputs(6582) <= '0';
    layer0_outputs(6583) <= not(inputs(205));
    layer0_outputs(6584) <= not(inputs(86)) or (inputs(190));
    layer0_outputs(6585) <= inputs(176);
    layer0_outputs(6586) <= not((inputs(120)) or (inputs(101)));
    layer0_outputs(6587) <= inputs(137);
    layer0_outputs(6588) <= (inputs(123)) or (inputs(117));
    layer0_outputs(6589) <= (inputs(148)) and not (inputs(246));
    layer0_outputs(6590) <= (inputs(100)) and not (inputs(112));
    layer0_outputs(6591) <= (inputs(187)) or (inputs(18));
    layer0_outputs(6592) <= not((inputs(107)) or (inputs(244)));
    layer0_outputs(6593) <= (inputs(88)) and (inputs(74));
    layer0_outputs(6594) <= inputs(110);
    layer0_outputs(6595) <= '1';
    layer0_outputs(6596) <= not(inputs(212));
    layer0_outputs(6597) <= not(inputs(118)) or (inputs(42));
    layer0_outputs(6598) <= not(inputs(1)) or (inputs(183));
    layer0_outputs(6599) <= (inputs(187)) or (inputs(40));
    layer0_outputs(6600) <= not(inputs(133));
    layer0_outputs(6601) <= (inputs(104)) and not (inputs(64));
    layer0_outputs(6602) <= not(inputs(164)) or (inputs(234));
    layer0_outputs(6603) <= not(inputs(253));
    layer0_outputs(6604) <= (inputs(206)) and not (inputs(125));
    layer0_outputs(6605) <= not((inputs(198)) or (inputs(197)));
    layer0_outputs(6606) <= not((inputs(212)) or (inputs(100)));
    layer0_outputs(6607) <= not(inputs(236)) or (inputs(60));
    layer0_outputs(6608) <= not(inputs(167)) or (inputs(161));
    layer0_outputs(6609) <= not(inputs(197));
    layer0_outputs(6610) <= not(inputs(137));
    layer0_outputs(6611) <= not(inputs(215));
    layer0_outputs(6612) <= (inputs(178)) and not (inputs(65));
    layer0_outputs(6613) <= (inputs(210)) and not (inputs(238));
    layer0_outputs(6614) <= not(inputs(213)) or (inputs(220));
    layer0_outputs(6615) <= inputs(117);
    layer0_outputs(6616) <= not((inputs(203)) xor (inputs(164)));
    layer0_outputs(6617) <= (inputs(155)) xor (inputs(156));
    layer0_outputs(6618) <= not((inputs(149)) or (inputs(126)));
    layer0_outputs(6619) <= inputs(115);
    layer0_outputs(6620) <= not(inputs(235)) or (inputs(52));
    layer0_outputs(6621) <= not(inputs(243));
    layer0_outputs(6622) <= not(inputs(134)) or (inputs(14));
    layer0_outputs(6623) <= '1';
    layer0_outputs(6624) <= not(inputs(53));
    layer0_outputs(6625) <= not(inputs(70));
    layer0_outputs(6626) <= not((inputs(108)) or (inputs(155)));
    layer0_outputs(6627) <= not(inputs(112));
    layer0_outputs(6628) <= inputs(19);
    layer0_outputs(6629) <= not(inputs(187)) or (inputs(98));
    layer0_outputs(6630) <= not(inputs(186)) or (inputs(89));
    layer0_outputs(6631) <= not((inputs(197)) or (inputs(48)));
    layer0_outputs(6632) <= (inputs(21)) or (inputs(47));
    layer0_outputs(6633) <= (inputs(101)) xor (inputs(152));
    layer0_outputs(6634) <= inputs(156);
    layer0_outputs(6635) <= not(inputs(198)) or (inputs(28));
    layer0_outputs(6636) <= (inputs(140)) and (inputs(124));
    layer0_outputs(6637) <= not((inputs(169)) xor (inputs(188)));
    layer0_outputs(6638) <= (inputs(206)) xor (inputs(191));
    layer0_outputs(6639) <= (inputs(7)) xor (inputs(206));
    layer0_outputs(6640) <= not((inputs(174)) or (inputs(181)));
    layer0_outputs(6641) <= not((inputs(211)) or (inputs(29)));
    layer0_outputs(6642) <= (inputs(60)) or (inputs(49));
    layer0_outputs(6643) <= not(inputs(104));
    layer0_outputs(6644) <= not((inputs(231)) or (inputs(134)));
    layer0_outputs(6645) <= not(inputs(78));
    layer0_outputs(6646) <= inputs(59);
    layer0_outputs(6647) <= (inputs(211)) and not (inputs(124));
    layer0_outputs(6648) <= not(inputs(251));
    layer0_outputs(6649) <= inputs(43);
    layer0_outputs(6650) <= inputs(227);
    layer0_outputs(6651) <= not(inputs(151));
    layer0_outputs(6652) <= not((inputs(135)) or (inputs(255)));
    layer0_outputs(6653) <= not(inputs(126)) or (inputs(241));
    layer0_outputs(6654) <= inputs(150);
    layer0_outputs(6655) <= '1';
    layer0_outputs(6656) <= inputs(144);
    layer0_outputs(6657) <= (inputs(121)) and not (inputs(7));
    layer0_outputs(6658) <= (inputs(184)) and not (inputs(124));
    layer0_outputs(6659) <= (inputs(241)) xor (inputs(7));
    layer0_outputs(6660) <= '0';
    layer0_outputs(6661) <= (inputs(44)) xor (inputs(114));
    layer0_outputs(6662) <= not(inputs(175));
    layer0_outputs(6663) <= not(inputs(181));
    layer0_outputs(6664) <= not((inputs(22)) or (inputs(80)));
    layer0_outputs(6665) <= not((inputs(238)) or (inputs(10)));
    layer0_outputs(6666) <= not(inputs(118));
    layer0_outputs(6667) <= (inputs(176)) and not (inputs(17));
    layer0_outputs(6668) <= (inputs(204)) and not (inputs(205));
    layer0_outputs(6669) <= not(inputs(105)) or (inputs(28));
    layer0_outputs(6670) <= (inputs(68)) or (inputs(231));
    layer0_outputs(6671) <= (inputs(66)) and not (inputs(176));
    layer0_outputs(6672) <= not((inputs(59)) xor (inputs(188)));
    layer0_outputs(6673) <= inputs(107);
    layer0_outputs(6674) <= not((inputs(134)) xor (inputs(26)));
    layer0_outputs(6675) <= (inputs(150)) and not (inputs(207));
    layer0_outputs(6676) <= (inputs(75)) xor (inputs(47));
    layer0_outputs(6677) <= not(inputs(229)) or (inputs(210));
    layer0_outputs(6678) <= (inputs(157)) or (inputs(195));
    layer0_outputs(6679) <= not((inputs(61)) or (inputs(29)));
    layer0_outputs(6680) <= inputs(78);
    layer0_outputs(6681) <= (inputs(185)) and not (inputs(81));
    layer0_outputs(6682) <= not((inputs(153)) xor (inputs(96)));
    layer0_outputs(6683) <= not(inputs(131)) or (inputs(20));
    layer0_outputs(6684) <= not(inputs(114));
    layer0_outputs(6685) <= (inputs(224)) xor (inputs(250));
    layer0_outputs(6686) <= not(inputs(115));
    layer0_outputs(6687) <= not(inputs(108));
    layer0_outputs(6688) <= (inputs(197)) or (inputs(183));
    layer0_outputs(6689) <= (inputs(230)) and not (inputs(11));
    layer0_outputs(6690) <= (inputs(178)) and not (inputs(143));
    layer0_outputs(6691) <= not(inputs(97)) or (inputs(241));
    layer0_outputs(6692) <= (inputs(236)) or (inputs(236));
    layer0_outputs(6693) <= (inputs(193)) and not (inputs(84));
    layer0_outputs(6694) <= not(inputs(55));
    layer0_outputs(6695) <= (inputs(85)) and not (inputs(36));
    layer0_outputs(6696) <= not((inputs(223)) or (inputs(101)));
    layer0_outputs(6697) <= not(inputs(211));
    layer0_outputs(6698) <= '0';
    layer0_outputs(6699) <= (inputs(240)) xor (inputs(85));
    layer0_outputs(6700) <= not((inputs(103)) xor (inputs(196)));
    layer0_outputs(6701) <= (inputs(224)) and (inputs(86));
    layer0_outputs(6702) <= not(inputs(196)) or (inputs(127));
    layer0_outputs(6703) <= (inputs(145)) xor (inputs(236));
    layer0_outputs(6704) <= (inputs(205)) xor (inputs(59));
    layer0_outputs(6705) <= not(inputs(136)) or (inputs(80));
    layer0_outputs(6706) <= (inputs(3)) or (inputs(229));
    layer0_outputs(6707) <= not(inputs(90)) or (inputs(119));
    layer0_outputs(6708) <= (inputs(104)) or (inputs(63));
    layer0_outputs(6709) <= not((inputs(92)) xor (inputs(6)));
    layer0_outputs(6710) <= not(inputs(183));
    layer0_outputs(6711) <= inputs(24);
    layer0_outputs(6712) <= (inputs(140)) or (inputs(124));
    layer0_outputs(6713) <= inputs(107);
    layer0_outputs(6714) <= '0';
    layer0_outputs(6715) <= not((inputs(181)) or (inputs(132)));
    layer0_outputs(6716) <= not(inputs(78)) or (inputs(31));
    layer0_outputs(6717) <= inputs(134);
    layer0_outputs(6718) <= inputs(180);
    layer0_outputs(6719) <= inputs(185);
    layer0_outputs(6720) <= '0';
    layer0_outputs(6721) <= (inputs(158)) or (inputs(39));
    layer0_outputs(6722) <= (inputs(157)) and (inputs(174));
    layer0_outputs(6723) <= inputs(121);
    layer0_outputs(6724) <= not(inputs(85));
    layer0_outputs(6725) <= (inputs(25)) xor (inputs(128));
    layer0_outputs(6726) <= (inputs(18)) and not (inputs(43));
    layer0_outputs(6727) <= (inputs(216)) or (inputs(180));
    layer0_outputs(6728) <= (inputs(174)) or (inputs(189));
    layer0_outputs(6729) <= (inputs(7)) and not (inputs(35));
    layer0_outputs(6730) <= not(inputs(168));
    layer0_outputs(6731) <= not((inputs(216)) or (inputs(251)));
    layer0_outputs(6732) <= not((inputs(22)) and (inputs(192)));
    layer0_outputs(6733) <= (inputs(207)) and (inputs(116));
    layer0_outputs(6734) <= (inputs(99)) or (inputs(28));
    layer0_outputs(6735) <= (inputs(128)) and not (inputs(14));
    layer0_outputs(6736) <= (inputs(171)) and not (inputs(131));
    layer0_outputs(6737) <= not((inputs(237)) and (inputs(190)));
    layer0_outputs(6738) <= (inputs(17)) xor (inputs(129));
    layer0_outputs(6739) <= (inputs(170)) xor (inputs(91));
    layer0_outputs(6740) <= (inputs(51)) or (inputs(218));
    layer0_outputs(6741) <= not(inputs(157));
    layer0_outputs(6742) <= (inputs(103)) and not (inputs(30));
    layer0_outputs(6743) <= (inputs(253)) or (inputs(124));
    layer0_outputs(6744) <= inputs(213);
    layer0_outputs(6745) <= not(inputs(213));
    layer0_outputs(6746) <= inputs(117);
    layer0_outputs(6747) <= (inputs(60)) or (inputs(97));
    layer0_outputs(6748) <= (inputs(89)) and not (inputs(13));
    layer0_outputs(6749) <= not((inputs(2)) and (inputs(95)));
    layer0_outputs(6750) <= (inputs(240)) or (inputs(5));
    layer0_outputs(6751) <= inputs(41);
    layer0_outputs(6752) <= (inputs(136)) and not (inputs(117));
    layer0_outputs(6753) <= (inputs(165)) or (inputs(99));
    layer0_outputs(6754) <= not((inputs(32)) and (inputs(6)));
    layer0_outputs(6755) <= inputs(114);
    layer0_outputs(6756) <= not(inputs(39));
    layer0_outputs(6757) <= (inputs(25)) or (inputs(233));
    layer0_outputs(6758) <= (inputs(19)) and not (inputs(18));
    layer0_outputs(6759) <= not(inputs(56)) or (inputs(133));
    layer0_outputs(6760) <= not((inputs(98)) xor (inputs(79)));
    layer0_outputs(6761) <= (inputs(127)) and not (inputs(113));
    layer0_outputs(6762) <= not(inputs(135));
    layer0_outputs(6763) <= '1';
    layer0_outputs(6764) <= (inputs(16)) and not (inputs(173));
    layer0_outputs(6765) <= inputs(251);
    layer0_outputs(6766) <= (inputs(158)) xor (inputs(93));
    layer0_outputs(6767) <= (inputs(154)) or (inputs(94));
    layer0_outputs(6768) <= not(inputs(6)) or (inputs(238));
    layer0_outputs(6769) <= (inputs(170)) or (inputs(23));
    layer0_outputs(6770) <= (inputs(120)) xor (inputs(34));
    layer0_outputs(6771) <= (inputs(97)) xor (inputs(209));
    layer0_outputs(6772) <= inputs(76);
    layer0_outputs(6773) <= (inputs(165)) xor (inputs(186));
    layer0_outputs(6774) <= inputs(90);
    layer0_outputs(6775) <= (inputs(18)) and (inputs(64));
    layer0_outputs(6776) <= not(inputs(190)) or (inputs(0));
    layer0_outputs(6777) <= inputs(176);
    layer0_outputs(6778) <= (inputs(159)) or (inputs(89));
    layer0_outputs(6779) <= (inputs(188)) and not (inputs(28));
    layer0_outputs(6780) <= inputs(247);
    layer0_outputs(6781) <= (inputs(152)) or (inputs(5));
    layer0_outputs(6782) <= inputs(89);
    layer0_outputs(6783) <= (inputs(122)) xor (inputs(77));
    layer0_outputs(6784) <= not(inputs(38));
    layer0_outputs(6785) <= not((inputs(219)) or (inputs(37)));
    layer0_outputs(6786) <= not((inputs(200)) or (inputs(229)));
    layer0_outputs(6787) <= (inputs(157)) and not (inputs(227));
    layer0_outputs(6788) <= not(inputs(119)) or (inputs(17));
    layer0_outputs(6789) <= (inputs(178)) or (inputs(163));
    layer0_outputs(6790) <= (inputs(114)) and (inputs(249));
    layer0_outputs(6791) <= not(inputs(59)) or (inputs(18));
    layer0_outputs(6792) <= (inputs(239)) or (inputs(106));
    layer0_outputs(6793) <= not((inputs(174)) or (inputs(213)));
    layer0_outputs(6794) <= not(inputs(209)) or (inputs(9));
    layer0_outputs(6795) <= not(inputs(133)) or (inputs(143));
    layer0_outputs(6796) <= (inputs(117)) and not (inputs(5));
    layer0_outputs(6797) <= (inputs(21)) or (inputs(59));
    layer0_outputs(6798) <= (inputs(131)) xor (inputs(223));
    layer0_outputs(6799) <= (inputs(202)) and not (inputs(133));
    layer0_outputs(6800) <= not(inputs(122)) or (inputs(65));
    layer0_outputs(6801) <= not(inputs(119));
    layer0_outputs(6802) <= not((inputs(153)) and (inputs(160)));
    layer0_outputs(6803) <= (inputs(2)) and not (inputs(5));
    layer0_outputs(6804) <= not((inputs(213)) xor (inputs(57)));
    layer0_outputs(6805) <= '0';
    layer0_outputs(6806) <= (inputs(100)) and not (inputs(98));
    layer0_outputs(6807) <= not((inputs(206)) xor (inputs(148)));
    layer0_outputs(6808) <= (inputs(199)) or (inputs(26));
    layer0_outputs(6809) <= inputs(72);
    layer0_outputs(6810) <= inputs(141);
    layer0_outputs(6811) <= inputs(144);
    layer0_outputs(6812) <= not(inputs(153));
    layer0_outputs(6813) <= not(inputs(240)) or (inputs(143));
    layer0_outputs(6814) <= not((inputs(74)) xor (inputs(244)));
    layer0_outputs(6815) <= (inputs(66)) xor (inputs(243));
    layer0_outputs(6816) <= (inputs(128)) xor (inputs(107));
    layer0_outputs(6817) <= (inputs(11)) and (inputs(241));
    layer0_outputs(6818) <= not(inputs(205)) or (inputs(9));
    layer0_outputs(6819) <= inputs(216);
    layer0_outputs(6820) <= inputs(117);
    layer0_outputs(6821) <= inputs(61);
    layer0_outputs(6822) <= (inputs(182)) and not (inputs(215));
    layer0_outputs(6823) <= (inputs(139)) and not (inputs(95));
    layer0_outputs(6824) <= not(inputs(123));
    layer0_outputs(6825) <= not(inputs(105));
    layer0_outputs(6826) <= not(inputs(212));
    layer0_outputs(6827) <= (inputs(146)) and not (inputs(18));
    layer0_outputs(6828) <= (inputs(139)) and not (inputs(164));
    layer0_outputs(6829) <= not(inputs(255)) or (inputs(103));
    layer0_outputs(6830) <= (inputs(225)) or (inputs(142));
    layer0_outputs(6831) <= not((inputs(194)) xor (inputs(31)));
    layer0_outputs(6832) <= not(inputs(178));
    layer0_outputs(6833) <= (inputs(225)) or (inputs(89));
    layer0_outputs(6834) <= '1';
    layer0_outputs(6835) <= (inputs(37)) and not (inputs(96));
    layer0_outputs(6836) <= not((inputs(58)) xor (inputs(55)));
    layer0_outputs(6837) <= not((inputs(52)) xor (inputs(248)));
    layer0_outputs(6838) <= not(inputs(148)) or (inputs(30));
    layer0_outputs(6839) <= '0';
    layer0_outputs(6840) <= not((inputs(131)) or (inputs(158)));
    layer0_outputs(6841) <= not(inputs(88)) or (inputs(8));
    layer0_outputs(6842) <= (inputs(214)) and not (inputs(240));
    layer0_outputs(6843) <= (inputs(160)) xor (inputs(193));
    layer0_outputs(6844) <= (inputs(4)) and not (inputs(255));
    layer0_outputs(6845) <= (inputs(182)) and not (inputs(227));
    layer0_outputs(6846) <= not((inputs(200)) xor (inputs(236)));
    layer0_outputs(6847) <= (inputs(73)) xor (inputs(57));
    layer0_outputs(6848) <= not(inputs(143)) or (inputs(124));
    layer0_outputs(6849) <= (inputs(210)) xor (inputs(224));
    layer0_outputs(6850) <= (inputs(238)) or (inputs(193));
    layer0_outputs(6851) <= '1';
    layer0_outputs(6852) <= (inputs(252)) and not (inputs(22));
    layer0_outputs(6853) <= not((inputs(243)) xor (inputs(51)));
    layer0_outputs(6854) <= not((inputs(158)) and (inputs(255)));
    layer0_outputs(6855) <= inputs(55);
    layer0_outputs(6856) <= not(inputs(195));
    layer0_outputs(6857) <= (inputs(6)) and (inputs(64));
    layer0_outputs(6858) <= inputs(151);
    layer0_outputs(6859) <= not((inputs(147)) or (inputs(142)));
    layer0_outputs(6860) <= inputs(61);
    layer0_outputs(6861) <= (inputs(28)) or (inputs(4));
    layer0_outputs(6862) <= not(inputs(38)) or (inputs(245));
    layer0_outputs(6863) <= not((inputs(47)) or (inputs(34)));
    layer0_outputs(6864) <= inputs(207);
    layer0_outputs(6865) <= not(inputs(56)) or (inputs(96));
    layer0_outputs(6866) <= (inputs(251)) or (inputs(235));
    layer0_outputs(6867) <= (inputs(231)) and not (inputs(33));
    layer0_outputs(6868) <= (inputs(94)) and not (inputs(239));
    layer0_outputs(6869) <= not(inputs(182)) or (inputs(242));
    layer0_outputs(6870) <= not(inputs(118)) or (inputs(205));
    layer0_outputs(6871) <= not(inputs(118)) or (inputs(81));
    layer0_outputs(6872) <= not(inputs(252)) or (inputs(195));
    layer0_outputs(6873) <= inputs(62);
    layer0_outputs(6874) <= inputs(131);
    layer0_outputs(6875) <= not((inputs(0)) or (inputs(225)));
    layer0_outputs(6876) <= not(inputs(100));
    layer0_outputs(6877) <= '1';
    layer0_outputs(6878) <= not(inputs(87));
    layer0_outputs(6879) <= (inputs(180)) or (inputs(205));
    layer0_outputs(6880) <= '0';
    layer0_outputs(6881) <= not((inputs(65)) or (inputs(88)));
    layer0_outputs(6882) <= (inputs(65)) or (inputs(176));
    layer0_outputs(6883) <= not((inputs(250)) or (inputs(151)));
    layer0_outputs(6884) <= not((inputs(38)) xor (inputs(153)));
    layer0_outputs(6885) <= not((inputs(67)) xor (inputs(98)));
    layer0_outputs(6886) <= (inputs(232)) xor (inputs(65));
    layer0_outputs(6887) <= (inputs(224)) and not (inputs(131));
    layer0_outputs(6888) <= not((inputs(68)) or (inputs(29)));
    layer0_outputs(6889) <= (inputs(53)) and not (inputs(80));
    layer0_outputs(6890) <= not(inputs(193)) or (inputs(65));
    layer0_outputs(6891) <= not(inputs(186));
    layer0_outputs(6892) <= not(inputs(129)) or (inputs(250));
    layer0_outputs(6893) <= (inputs(80)) and (inputs(246));
    layer0_outputs(6894) <= (inputs(116)) xor (inputs(68));
    layer0_outputs(6895) <= (inputs(187)) and not (inputs(179));
    layer0_outputs(6896) <= not((inputs(133)) and (inputs(165)));
    layer0_outputs(6897) <= not((inputs(86)) or (inputs(175)));
    layer0_outputs(6898) <= not(inputs(196)) or (inputs(16));
    layer0_outputs(6899) <= not(inputs(106)) or (inputs(28));
    layer0_outputs(6900) <= not(inputs(165));
    layer0_outputs(6901) <= (inputs(167)) and not (inputs(180));
    layer0_outputs(6902) <= (inputs(160)) and not (inputs(10));
    layer0_outputs(6903) <= (inputs(244)) or (inputs(105));
    layer0_outputs(6904) <= not(inputs(101));
    layer0_outputs(6905) <= not((inputs(21)) or (inputs(240)));
    layer0_outputs(6906) <= (inputs(0)) and not (inputs(252));
    layer0_outputs(6907) <= not(inputs(49));
    layer0_outputs(6908) <= (inputs(171)) or (inputs(244));
    layer0_outputs(6909) <= inputs(181);
    layer0_outputs(6910) <= not(inputs(102)) or (inputs(82));
    layer0_outputs(6911) <= inputs(28);
    layer0_outputs(6912) <= (inputs(87)) xor (inputs(240));
    layer0_outputs(6913) <= not(inputs(137)) or (inputs(147));
    layer0_outputs(6914) <= not((inputs(205)) or (inputs(19)));
    layer0_outputs(6915) <= (inputs(166)) or (inputs(177));
    layer0_outputs(6916) <= (inputs(200)) or (inputs(156));
    layer0_outputs(6917) <= (inputs(203)) and (inputs(183));
    layer0_outputs(6918) <= (inputs(175)) or (inputs(2));
    layer0_outputs(6919) <= inputs(120);
    layer0_outputs(6920) <= not(inputs(102));
    layer0_outputs(6921) <= (inputs(110)) and (inputs(0));
    layer0_outputs(6922) <= (inputs(92)) and (inputs(147));
    layer0_outputs(6923) <= (inputs(144)) and not (inputs(248));
    layer0_outputs(6924) <= not(inputs(23));
    layer0_outputs(6925) <= inputs(128);
    layer0_outputs(6926) <= not((inputs(181)) or (inputs(203)));
    layer0_outputs(6927) <= not(inputs(247)) or (inputs(16));
    layer0_outputs(6928) <= not((inputs(11)) and (inputs(215)));
    layer0_outputs(6929) <= not(inputs(185));
    layer0_outputs(6930) <= not((inputs(197)) xor (inputs(198)));
    layer0_outputs(6931) <= not(inputs(66));
    layer0_outputs(6932) <= (inputs(235)) or (inputs(214));
    layer0_outputs(6933) <= not(inputs(105));
    layer0_outputs(6934) <= inputs(31);
    layer0_outputs(6935) <= inputs(127);
    layer0_outputs(6936) <= not(inputs(245));
    layer0_outputs(6937) <= not(inputs(184)) or (inputs(14));
    layer0_outputs(6938) <= (inputs(74)) and not (inputs(247));
    layer0_outputs(6939) <= inputs(90);
    layer0_outputs(6940) <= (inputs(80)) and not (inputs(207));
    layer0_outputs(6941) <= not(inputs(81));
    layer0_outputs(6942) <= not((inputs(112)) or (inputs(108)));
    layer0_outputs(6943) <= (inputs(211)) and not (inputs(49));
    layer0_outputs(6944) <= (inputs(9)) xor (inputs(217));
    layer0_outputs(6945) <= not(inputs(122));
    layer0_outputs(6946) <= (inputs(53)) xor (inputs(57));
    layer0_outputs(6947) <= (inputs(179)) xor (inputs(41));
    layer0_outputs(6948) <= inputs(226);
    layer0_outputs(6949) <= inputs(230);
    layer0_outputs(6950) <= not((inputs(243)) or (inputs(166)));
    layer0_outputs(6951) <= (inputs(55)) xor (inputs(43));
    layer0_outputs(6952) <= (inputs(102)) and not (inputs(174));
    layer0_outputs(6953) <= not(inputs(18)) or (inputs(174));
    layer0_outputs(6954) <= not(inputs(27)) or (inputs(139));
    layer0_outputs(6955) <= inputs(153);
    layer0_outputs(6956) <= not(inputs(84)) or (inputs(252));
    layer0_outputs(6957) <= not((inputs(140)) xor (inputs(125)));
    layer0_outputs(6958) <= (inputs(84)) and (inputs(32));
    layer0_outputs(6959) <= (inputs(197)) or (inputs(72));
    layer0_outputs(6960) <= not(inputs(108)) or (inputs(227));
    layer0_outputs(6961) <= inputs(229);
    layer0_outputs(6962) <= not(inputs(57)) or (inputs(172));
    layer0_outputs(6963) <= (inputs(101)) and not (inputs(228));
    layer0_outputs(6964) <= (inputs(46)) xor (inputs(92));
    layer0_outputs(6965) <= inputs(73);
    layer0_outputs(6966) <= inputs(153);
    layer0_outputs(6967) <= not(inputs(98)) or (inputs(23));
    layer0_outputs(6968) <= (inputs(3)) and (inputs(2));
    layer0_outputs(6969) <= not(inputs(9)) or (inputs(208));
    layer0_outputs(6970) <= (inputs(243)) and not (inputs(15));
    layer0_outputs(6971) <= not((inputs(31)) xor (inputs(121)));
    layer0_outputs(6972) <= not((inputs(120)) or (inputs(190)));
    layer0_outputs(6973) <= inputs(49);
    layer0_outputs(6974) <= (inputs(197)) and not (inputs(96));
    layer0_outputs(6975) <= (inputs(199)) xor (inputs(206));
    layer0_outputs(6976) <= (inputs(71)) and not (inputs(156));
    layer0_outputs(6977) <= not(inputs(141));
    layer0_outputs(6978) <= not(inputs(49)) or (inputs(239));
    layer0_outputs(6979) <= not((inputs(196)) or (inputs(12)));
    layer0_outputs(6980) <= (inputs(169)) or (inputs(95));
    layer0_outputs(6981) <= not(inputs(116));
    layer0_outputs(6982) <= '0';
    layer0_outputs(6983) <= (inputs(233)) and not (inputs(176));
    layer0_outputs(6984) <= not((inputs(58)) xor (inputs(251)));
    layer0_outputs(6985) <= inputs(224);
    layer0_outputs(6986) <= not(inputs(158)) or (inputs(60));
    layer0_outputs(6987) <= inputs(107);
    layer0_outputs(6988) <= not(inputs(52));
    layer0_outputs(6989) <= not(inputs(62)) or (inputs(17));
    layer0_outputs(6990) <= (inputs(37)) xor (inputs(76));
    layer0_outputs(6991) <= not(inputs(253)) or (inputs(230));
    layer0_outputs(6992) <= (inputs(45)) or (inputs(12));
    layer0_outputs(6993) <= not(inputs(82));
    layer0_outputs(6994) <= (inputs(97)) and (inputs(207));
    layer0_outputs(6995) <= inputs(155);
    layer0_outputs(6996) <= not(inputs(104)) or (inputs(131));
    layer0_outputs(6997) <= inputs(117);
    layer0_outputs(6998) <= not(inputs(153)) or (inputs(75));
    layer0_outputs(6999) <= not(inputs(149));
    layer0_outputs(7000) <= (inputs(223)) xor (inputs(233));
    layer0_outputs(7001) <= not((inputs(88)) or (inputs(23)));
    layer0_outputs(7002) <= not((inputs(205)) or (inputs(98)));
    layer0_outputs(7003) <= not(inputs(177)) or (inputs(13));
    layer0_outputs(7004) <= not((inputs(66)) xor (inputs(19)));
    layer0_outputs(7005) <= '1';
    layer0_outputs(7006) <= (inputs(214)) xor (inputs(193));
    layer0_outputs(7007) <= (inputs(106)) and not (inputs(34));
    layer0_outputs(7008) <= not(inputs(109)) or (inputs(26));
    layer0_outputs(7009) <= (inputs(175)) or (inputs(1));
    layer0_outputs(7010) <= not(inputs(233));
    layer0_outputs(7011) <= inputs(116);
    layer0_outputs(7012) <= (inputs(248)) xor (inputs(59));
    layer0_outputs(7013) <= (inputs(54)) xor (inputs(187));
    layer0_outputs(7014) <= not(inputs(135));
    layer0_outputs(7015) <= inputs(125);
    layer0_outputs(7016) <= '1';
    layer0_outputs(7017) <= not(inputs(133)) or (inputs(211));
    layer0_outputs(7018) <= not(inputs(54));
    layer0_outputs(7019) <= '1';
    layer0_outputs(7020) <= not((inputs(184)) or (inputs(16)));
    layer0_outputs(7021) <= not(inputs(43));
    layer0_outputs(7022) <= '0';
    layer0_outputs(7023) <= not((inputs(22)) xor (inputs(27)));
    layer0_outputs(7024) <= not((inputs(234)) xor (inputs(216)));
    layer0_outputs(7025) <= not(inputs(242)) or (inputs(31));
    layer0_outputs(7026) <= not((inputs(248)) or (inputs(74)));
    layer0_outputs(7027) <= not(inputs(215));
    layer0_outputs(7028) <= not((inputs(64)) xor (inputs(16)));
    layer0_outputs(7029) <= '0';
    layer0_outputs(7030) <= inputs(198);
    layer0_outputs(7031) <= (inputs(72)) xor (inputs(183));
    layer0_outputs(7032) <= not((inputs(230)) xor (inputs(202)));
    layer0_outputs(7033) <= (inputs(216)) and not (inputs(158));
    layer0_outputs(7034) <= not((inputs(198)) or (inputs(94)));
    layer0_outputs(7035) <= (inputs(226)) and not (inputs(21));
    layer0_outputs(7036) <= (inputs(78)) and not (inputs(34));
    layer0_outputs(7037) <= inputs(60);
    layer0_outputs(7038) <= not((inputs(88)) xor (inputs(244)));
    layer0_outputs(7039) <= (inputs(217)) and not (inputs(141));
    layer0_outputs(7040) <= not((inputs(110)) xor (inputs(111)));
    layer0_outputs(7041) <= (inputs(159)) and not (inputs(139));
    layer0_outputs(7042) <= (inputs(149)) and not (inputs(242));
    layer0_outputs(7043) <= not((inputs(241)) xor (inputs(102)));
    layer0_outputs(7044) <= not(inputs(123)) or (inputs(217));
    layer0_outputs(7045) <= (inputs(60)) or (inputs(245));
    layer0_outputs(7046) <= not((inputs(118)) or (inputs(164)));
    layer0_outputs(7047) <= not(inputs(76));
    layer0_outputs(7048) <= inputs(160);
    layer0_outputs(7049) <= not((inputs(214)) or (inputs(229)));
    layer0_outputs(7050) <= (inputs(243)) and (inputs(42));
    layer0_outputs(7051) <= not(inputs(135)) or (inputs(43));
    layer0_outputs(7052) <= not((inputs(147)) xor (inputs(112)));
    layer0_outputs(7053) <= inputs(79);
    layer0_outputs(7054) <= not(inputs(235));
    layer0_outputs(7055) <= (inputs(234)) or (inputs(94));
    layer0_outputs(7056) <= not((inputs(185)) or (inputs(7)));
    layer0_outputs(7057) <= (inputs(165)) xor (inputs(35));
    layer0_outputs(7058) <= (inputs(144)) and not (inputs(127));
    layer0_outputs(7059) <= not(inputs(58)) or (inputs(65));
    layer0_outputs(7060) <= not((inputs(100)) or (inputs(250)));
    layer0_outputs(7061) <= '0';
    layer0_outputs(7062) <= (inputs(183)) and not (inputs(63));
    layer0_outputs(7063) <= not(inputs(129)) or (inputs(198));
    layer0_outputs(7064) <= not(inputs(154));
    layer0_outputs(7065) <= not(inputs(52));
    layer0_outputs(7066) <= (inputs(196)) or (inputs(207));
    layer0_outputs(7067) <= (inputs(205)) xor (inputs(108));
    layer0_outputs(7068) <= '1';
    layer0_outputs(7069) <= (inputs(202)) and not (inputs(142));
    layer0_outputs(7070) <= (inputs(88)) and not (inputs(158));
    layer0_outputs(7071) <= not(inputs(228)) or (inputs(2));
    layer0_outputs(7072) <= not(inputs(228)) or (inputs(111));
    layer0_outputs(7073) <= not((inputs(219)) or (inputs(155)));
    layer0_outputs(7074) <= not((inputs(169)) or (inputs(4)));
    layer0_outputs(7075) <= inputs(229);
    layer0_outputs(7076) <= not(inputs(87));
    layer0_outputs(7077) <= (inputs(246)) and (inputs(63));
    layer0_outputs(7078) <= not(inputs(128)) or (inputs(31));
    layer0_outputs(7079) <= (inputs(156)) or (inputs(41));
    layer0_outputs(7080) <= not((inputs(192)) xor (inputs(117)));
    layer0_outputs(7081) <= not(inputs(213));
    layer0_outputs(7082) <= (inputs(165)) and not (inputs(39));
    layer0_outputs(7083) <= not(inputs(122)) or (inputs(127));
    layer0_outputs(7084) <= (inputs(39)) and not (inputs(249));
    layer0_outputs(7085) <= inputs(245);
    layer0_outputs(7086) <= not(inputs(166)) or (inputs(102));
    layer0_outputs(7087) <= inputs(72);
    layer0_outputs(7088) <= inputs(99);
    layer0_outputs(7089) <= not(inputs(89));
    layer0_outputs(7090) <= '1';
    layer0_outputs(7091) <= inputs(152);
    layer0_outputs(7092) <= not(inputs(189)) or (inputs(76));
    layer0_outputs(7093) <= (inputs(215)) and not (inputs(28));
    layer0_outputs(7094) <= inputs(93);
    layer0_outputs(7095) <= inputs(192);
    layer0_outputs(7096) <= (inputs(251)) or (inputs(96));
    layer0_outputs(7097) <= (inputs(4)) or (inputs(129));
    layer0_outputs(7098) <= inputs(58);
    layer0_outputs(7099) <= not((inputs(33)) xor (inputs(43)));
    layer0_outputs(7100) <= not((inputs(64)) or (inputs(95)));
    layer0_outputs(7101) <= inputs(204);
    layer0_outputs(7102) <= (inputs(200)) xor (inputs(38));
    layer0_outputs(7103) <= '1';
    layer0_outputs(7104) <= not((inputs(222)) or (inputs(211)));
    layer0_outputs(7105) <= not((inputs(2)) or (inputs(51)));
    layer0_outputs(7106) <= not(inputs(146)) or (inputs(255));
    layer0_outputs(7107) <= not(inputs(99)) or (inputs(81));
    layer0_outputs(7108) <= (inputs(90)) xor (inputs(11));
    layer0_outputs(7109) <= inputs(75);
    layer0_outputs(7110) <= not((inputs(108)) xor (inputs(79)));
    layer0_outputs(7111) <= '0';
    layer0_outputs(7112) <= (inputs(202)) xor (inputs(63));
    layer0_outputs(7113) <= '0';
    layer0_outputs(7114) <= inputs(96);
    layer0_outputs(7115) <= (inputs(136)) or (inputs(234));
    layer0_outputs(7116) <= (inputs(137)) and not (inputs(170));
    layer0_outputs(7117) <= (inputs(83)) or (inputs(79));
    layer0_outputs(7118) <= (inputs(14)) or (inputs(175));
    layer0_outputs(7119) <= (inputs(204)) and not (inputs(204));
    layer0_outputs(7120) <= (inputs(45)) xor (inputs(243));
    layer0_outputs(7121) <= inputs(90);
    layer0_outputs(7122) <= not((inputs(62)) or (inputs(185)));
    layer0_outputs(7123) <= not((inputs(74)) xor (inputs(237)));
    layer0_outputs(7124) <= not(inputs(141));
    layer0_outputs(7125) <= not((inputs(167)) or (inputs(125)));
    layer0_outputs(7126) <= not(inputs(200)) or (inputs(235));
    layer0_outputs(7127) <= not(inputs(91)) or (inputs(16));
    layer0_outputs(7128) <= not(inputs(91));
    layer0_outputs(7129) <= not(inputs(123)) or (inputs(32));
    layer0_outputs(7130) <= inputs(101);
    layer0_outputs(7131) <= (inputs(174)) or (inputs(124));
    layer0_outputs(7132) <= inputs(152);
    layer0_outputs(7133) <= not((inputs(104)) xor (inputs(44)));
    layer0_outputs(7134) <= (inputs(42)) or (inputs(7));
    layer0_outputs(7135) <= (inputs(158)) xor (inputs(156));
    layer0_outputs(7136) <= not(inputs(230));
    layer0_outputs(7137) <= not((inputs(129)) or (inputs(193)));
    layer0_outputs(7138) <= not((inputs(16)) xor (inputs(123)));
    layer0_outputs(7139) <= (inputs(29)) or (inputs(244));
    layer0_outputs(7140) <= (inputs(219)) and (inputs(95));
    layer0_outputs(7141) <= not((inputs(136)) and (inputs(5)));
    layer0_outputs(7142) <= (inputs(99)) and not (inputs(195));
    layer0_outputs(7143) <= (inputs(88)) and not (inputs(69));
    layer0_outputs(7144) <= not(inputs(201)) or (inputs(57));
    layer0_outputs(7145) <= '0';
    layer0_outputs(7146) <= (inputs(72)) or (inputs(93));
    layer0_outputs(7147) <= not(inputs(117));
    layer0_outputs(7148) <= (inputs(27)) and not (inputs(17));
    layer0_outputs(7149) <= (inputs(247)) xor (inputs(74));
    layer0_outputs(7150) <= not(inputs(90));
    layer0_outputs(7151) <= not(inputs(71)) or (inputs(177));
    layer0_outputs(7152) <= not(inputs(104)) or (inputs(187));
    layer0_outputs(7153) <= not(inputs(74)) or (inputs(6));
    layer0_outputs(7154) <= not(inputs(93));
    layer0_outputs(7155) <= inputs(138);
    layer0_outputs(7156) <= (inputs(38)) or (inputs(149));
    layer0_outputs(7157) <= not((inputs(182)) or (inputs(37)));
    layer0_outputs(7158) <= (inputs(179)) and not (inputs(131));
    layer0_outputs(7159) <= inputs(71);
    layer0_outputs(7160) <= inputs(116);
    layer0_outputs(7161) <= not(inputs(189));
    layer0_outputs(7162) <= not((inputs(86)) xor (inputs(225)));
    layer0_outputs(7163) <= not(inputs(21)) or (inputs(192));
    layer0_outputs(7164) <= not(inputs(251)) or (inputs(22));
    layer0_outputs(7165) <= not(inputs(103));
    layer0_outputs(7166) <= not((inputs(60)) or (inputs(151)));
    layer0_outputs(7167) <= (inputs(109)) or (inputs(11));
    layer0_outputs(7168) <= not((inputs(30)) or (inputs(30)));
    layer0_outputs(7169) <= '1';
    layer0_outputs(7170) <= (inputs(76)) or (inputs(83));
    layer0_outputs(7171) <= not((inputs(101)) xor (inputs(251)));
    layer0_outputs(7172) <= not((inputs(246)) xor (inputs(8)));
    layer0_outputs(7173) <= (inputs(164)) xor (inputs(55));
    layer0_outputs(7174) <= not((inputs(133)) or (inputs(192)));
    layer0_outputs(7175) <= (inputs(145)) xor (inputs(75));
    layer0_outputs(7176) <= not((inputs(23)) xor (inputs(250)));
    layer0_outputs(7177) <= (inputs(225)) and (inputs(199));
    layer0_outputs(7178) <= '0';
    layer0_outputs(7179) <= (inputs(135)) or (inputs(78));
    layer0_outputs(7180) <= inputs(151);
    layer0_outputs(7181) <= (inputs(214)) or (inputs(92));
    layer0_outputs(7182) <= inputs(164);
    layer0_outputs(7183) <= not(inputs(185));
    layer0_outputs(7184) <= not(inputs(148));
    layer0_outputs(7185) <= not(inputs(138)) or (inputs(190));
    layer0_outputs(7186) <= not(inputs(112)) or (inputs(22));
    layer0_outputs(7187) <= not(inputs(85));
    layer0_outputs(7188) <= not(inputs(125));
    layer0_outputs(7189) <= (inputs(70)) or (inputs(109));
    layer0_outputs(7190) <= inputs(230);
    layer0_outputs(7191) <= (inputs(103)) xor (inputs(97));
    layer0_outputs(7192) <= not((inputs(250)) xor (inputs(106)));
    layer0_outputs(7193) <= not(inputs(143)) or (inputs(28));
    layer0_outputs(7194) <= (inputs(165)) and not (inputs(251));
    layer0_outputs(7195) <= not((inputs(126)) or (inputs(135)));
    layer0_outputs(7196) <= (inputs(199)) or (inputs(25));
    layer0_outputs(7197) <= inputs(154);
    layer0_outputs(7198) <= not((inputs(146)) xor (inputs(58)));
    layer0_outputs(7199) <= not(inputs(199)) or (inputs(18));
    layer0_outputs(7200) <= '1';
    layer0_outputs(7201) <= not(inputs(125)) or (inputs(9));
    layer0_outputs(7202) <= not(inputs(233)) or (inputs(193));
    layer0_outputs(7203) <= not((inputs(165)) or (inputs(53)));
    layer0_outputs(7204) <= inputs(131);
    layer0_outputs(7205) <= (inputs(209)) xor (inputs(121));
    layer0_outputs(7206) <= (inputs(203)) or (inputs(5));
    layer0_outputs(7207) <= not(inputs(213));
    layer0_outputs(7208) <= '0';
    layer0_outputs(7209) <= (inputs(158)) xor (inputs(224));
    layer0_outputs(7210) <= not(inputs(215));
    layer0_outputs(7211) <= (inputs(92)) or (inputs(62));
    layer0_outputs(7212) <= not(inputs(16));
    layer0_outputs(7213) <= not((inputs(225)) xor (inputs(185)));
    layer0_outputs(7214) <= (inputs(226)) or (inputs(220));
    layer0_outputs(7215) <= not((inputs(187)) xor (inputs(196)));
    layer0_outputs(7216) <= (inputs(233)) or (inputs(69));
    layer0_outputs(7217) <= inputs(173);
    layer0_outputs(7218) <= not(inputs(103));
    layer0_outputs(7219) <= not((inputs(22)) xor (inputs(130)));
    layer0_outputs(7220) <= (inputs(106)) and not (inputs(203));
    layer0_outputs(7221) <= not((inputs(177)) or (inputs(137)));
    layer0_outputs(7222) <= (inputs(214)) and not (inputs(156));
    layer0_outputs(7223) <= (inputs(10)) or (inputs(52));
    layer0_outputs(7224) <= not(inputs(84));
    layer0_outputs(7225) <= not((inputs(190)) xor (inputs(254)));
    layer0_outputs(7226) <= not(inputs(35)) or (inputs(109));
    layer0_outputs(7227) <= not(inputs(239));
    layer0_outputs(7228) <= (inputs(170)) xor (inputs(12));
    layer0_outputs(7229) <= (inputs(132)) and not (inputs(24));
    layer0_outputs(7230) <= not((inputs(17)) or (inputs(218)));
    layer0_outputs(7231) <= not((inputs(36)) xor (inputs(181)));
    layer0_outputs(7232) <= inputs(149);
    layer0_outputs(7233) <= not((inputs(37)) or (inputs(111)));
    layer0_outputs(7234) <= not((inputs(79)) xor (inputs(61)));
    layer0_outputs(7235) <= (inputs(190)) or (inputs(213));
    layer0_outputs(7236) <= (inputs(183)) or (inputs(147));
    layer0_outputs(7237) <= inputs(5);
    layer0_outputs(7238) <= not((inputs(129)) xor (inputs(201)));
    layer0_outputs(7239) <= not(inputs(194));
    layer0_outputs(7240) <= inputs(82);
    layer0_outputs(7241) <= '1';
    layer0_outputs(7242) <= (inputs(10)) and not (inputs(208));
    layer0_outputs(7243) <= inputs(97);
    layer0_outputs(7244) <= '1';
    layer0_outputs(7245) <= not(inputs(207)) or (inputs(78));
    layer0_outputs(7246) <= not(inputs(2)) or (inputs(45));
    layer0_outputs(7247) <= '1';
    layer0_outputs(7248) <= (inputs(69)) and not (inputs(108));
    layer0_outputs(7249) <= not(inputs(244));
    layer0_outputs(7250) <= not((inputs(81)) xor (inputs(249)));
    layer0_outputs(7251) <= (inputs(153)) and not (inputs(240));
    layer0_outputs(7252) <= not((inputs(131)) or (inputs(226)));
    layer0_outputs(7253) <= not(inputs(200));
    layer0_outputs(7254) <= (inputs(19)) or (inputs(152));
    layer0_outputs(7255) <= inputs(197);
    layer0_outputs(7256) <= not(inputs(182)) or (inputs(91));
    layer0_outputs(7257) <= not(inputs(27)) or (inputs(31));
    layer0_outputs(7258) <= (inputs(175)) xor (inputs(179));
    layer0_outputs(7259) <= not(inputs(117)) or (inputs(38));
    layer0_outputs(7260) <= (inputs(46)) and not (inputs(145));
    layer0_outputs(7261) <= not(inputs(227)) or (inputs(251));
    layer0_outputs(7262) <= not((inputs(229)) xor (inputs(240)));
    layer0_outputs(7263) <= inputs(247);
    layer0_outputs(7264) <= not((inputs(54)) or (inputs(83)));
    layer0_outputs(7265) <= (inputs(178)) or (inputs(199));
    layer0_outputs(7266) <= (inputs(35)) and not (inputs(219));
    layer0_outputs(7267) <= not(inputs(200));
    layer0_outputs(7268) <= not((inputs(215)) or (inputs(17)));
    layer0_outputs(7269) <= (inputs(55)) or (inputs(227));
    layer0_outputs(7270) <= inputs(108);
    layer0_outputs(7271) <= inputs(209);
    layer0_outputs(7272) <= inputs(208);
    layer0_outputs(7273) <= not(inputs(90));
    layer0_outputs(7274) <= (inputs(121)) or (inputs(230));
    layer0_outputs(7275) <= (inputs(69)) or (inputs(191));
    layer0_outputs(7276) <= '0';
    layer0_outputs(7277) <= (inputs(228)) or (inputs(173));
    layer0_outputs(7278) <= (inputs(167)) or (inputs(43));
    layer0_outputs(7279) <= not(inputs(132)) or (inputs(235));
    layer0_outputs(7280) <= not(inputs(69));
    layer0_outputs(7281) <= (inputs(27)) and (inputs(142));
    layer0_outputs(7282) <= not(inputs(24));
    layer0_outputs(7283) <= not((inputs(19)) xor (inputs(28)));
    layer0_outputs(7284) <= not((inputs(220)) xor (inputs(219)));
    layer0_outputs(7285) <= not((inputs(192)) xor (inputs(179)));
    layer0_outputs(7286) <= (inputs(27)) and not (inputs(25));
    layer0_outputs(7287) <= not((inputs(67)) xor (inputs(194)));
    layer0_outputs(7288) <= not(inputs(122));
    layer0_outputs(7289) <= not(inputs(195)) or (inputs(226));
    layer0_outputs(7290) <= not((inputs(197)) xor (inputs(18)));
    layer0_outputs(7291) <= (inputs(46)) or (inputs(131));
    layer0_outputs(7292) <= not((inputs(202)) xor (inputs(190)));
    layer0_outputs(7293) <= inputs(75);
    layer0_outputs(7294) <= not(inputs(180)) or (inputs(17));
    layer0_outputs(7295) <= not((inputs(172)) or (inputs(200)));
    layer0_outputs(7296) <= inputs(121);
    layer0_outputs(7297) <= not((inputs(186)) and (inputs(211)));
    layer0_outputs(7298) <= (inputs(166)) or (inputs(124));
    layer0_outputs(7299) <= not((inputs(150)) or (inputs(168)));
    layer0_outputs(7300) <= not(inputs(119)) or (inputs(177));
    layer0_outputs(7301) <= (inputs(172)) or (inputs(29));
    layer0_outputs(7302) <= not((inputs(5)) or (inputs(98)));
    layer0_outputs(7303) <= not(inputs(80));
    layer0_outputs(7304) <= (inputs(130)) or (inputs(243));
    layer0_outputs(7305) <= (inputs(42)) and not (inputs(223));
    layer0_outputs(7306) <= (inputs(245)) or (inputs(68));
    layer0_outputs(7307) <= not(inputs(102));
    layer0_outputs(7308) <= not(inputs(196)) or (inputs(119));
    layer0_outputs(7309) <= (inputs(231)) or (inputs(57));
    layer0_outputs(7310) <= not((inputs(68)) or (inputs(42)));
    layer0_outputs(7311) <= not((inputs(155)) xor (inputs(103)));
    layer0_outputs(7312) <= not((inputs(144)) or (inputs(85)));
    layer0_outputs(7313) <= not(inputs(93));
    layer0_outputs(7314) <= not(inputs(133));
    layer0_outputs(7315) <= (inputs(94)) xor (inputs(106));
    layer0_outputs(7316) <= (inputs(122)) and not (inputs(208));
    layer0_outputs(7317) <= not(inputs(137));
    layer0_outputs(7318) <= not(inputs(153)) or (inputs(25));
    layer0_outputs(7319) <= not((inputs(73)) xor (inputs(217)));
    layer0_outputs(7320) <= (inputs(204)) xor (inputs(89));
    layer0_outputs(7321) <= not(inputs(232));
    layer0_outputs(7322) <= not(inputs(59)) or (inputs(112));
    layer0_outputs(7323) <= inputs(201);
    layer0_outputs(7324) <= inputs(36);
    layer0_outputs(7325) <= not((inputs(181)) xor (inputs(126)));
    layer0_outputs(7326) <= inputs(147);
    layer0_outputs(7327) <= (inputs(250)) and not (inputs(253));
    layer0_outputs(7328) <= inputs(61);
    layer0_outputs(7329) <= (inputs(161)) or (inputs(230));
    layer0_outputs(7330) <= '1';
    layer0_outputs(7331) <= not((inputs(22)) xor (inputs(108)));
    layer0_outputs(7332) <= (inputs(163)) xor (inputs(143));
    layer0_outputs(7333) <= (inputs(41)) and (inputs(149));
    layer0_outputs(7334) <= inputs(108);
    layer0_outputs(7335) <= not(inputs(91)) or (inputs(242));
    layer0_outputs(7336) <= not((inputs(48)) xor (inputs(249)));
    layer0_outputs(7337) <= not(inputs(120));
    layer0_outputs(7338) <= not((inputs(61)) or (inputs(187)));
    layer0_outputs(7339) <= (inputs(190)) and not (inputs(101));
    layer0_outputs(7340) <= not((inputs(82)) or (inputs(106)));
    layer0_outputs(7341) <= not(inputs(98)) or (inputs(20));
    layer0_outputs(7342) <= (inputs(179)) xor (inputs(244));
    layer0_outputs(7343) <= (inputs(201)) xor (inputs(106));
    layer0_outputs(7344) <= not((inputs(172)) and (inputs(85)));
    layer0_outputs(7345) <= (inputs(90)) or (inputs(195));
    layer0_outputs(7346) <= not((inputs(93)) xor (inputs(26)));
    layer0_outputs(7347) <= not(inputs(173));
    layer0_outputs(7348) <= inputs(137);
    layer0_outputs(7349) <= not((inputs(80)) xor (inputs(155)));
    layer0_outputs(7350) <= (inputs(132)) xor (inputs(89));
    layer0_outputs(7351) <= '1';
    layer0_outputs(7352) <= not(inputs(189)) or (inputs(179));
    layer0_outputs(7353) <= not(inputs(35));
    layer0_outputs(7354) <= not(inputs(224)) or (inputs(114));
    layer0_outputs(7355) <= not((inputs(124)) and (inputs(201)));
    layer0_outputs(7356) <= not(inputs(157)) or (inputs(76));
    layer0_outputs(7357) <= not((inputs(237)) or (inputs(228)));
    layer0_outputs(7358) <= not(inputs(74)) or (inputs(131));
    layer0_outputs(7359) <= not((inputs(253)) xor (inputs(8)));
    layer0_outputs(7360) <= not(inputs(227)) or (inputs(43));
    layer0_outputs(7361) <= inputs(133);
    layer0_outputs(7362) <= '1';
    layer0_outputs(7363) <= (inputs(62)) or (inputs(100));
    layer0_outputs(7364) <= not(inputs(8));
    layer0_outputs(7365) <= inputs(95);
    layer0_outputs(7366) <= (inputs(103)) and not (inputs(142));
    layer0_outputs(7367) <= (inputs(130)) or (inputs(154));
    layer0_outputs(7368) <= (inputs(173)) and not (inputs(15));
    layer0_outputs(7369) <= (inputs(17)) xor (inputs(213));
    layer0_outputs(7370) <= (inputs(5)) or (inputs(39));
    layer0_outputs(7371) <= not(inputs(253)) or (inputs(209));
    layer0_outputs(7372) <= not(inputs(121));
    layer0_outputs(7373) <= not(inputs(175));
    layer0_outputs(7374) <= not(inputs(71)) or (inputs(125));
    layer0_outputs(7375) <= not(inputs(141)) or (inputs(144));
    layer0_outputs(7376) <= not((inputs(153)) xor (inputs(135)));
    layer0_outputs(7377) <= not(inputs(167));
    layer0_outputs(7378) <= not((inputs(201)) or (inputs(53)));
    layer0_outputs(7379) <= inputs(12);
    layer0_outputs(7380) <= not(inputs(206)) or (inputs(81));
    layer0_outputs(7381) <= (inputs(59)) or (inputs(103));
    layer0_outputs(7382) <= inputs(157);
    layer0_outputs(7383) <= (inputs(199)) or (inputs(85));
    layer0_outputs(7384) <= inputs(4);
    layer0_outputs(7385) <= not(inputs(102));
    layer0_outputs(7386) <= not((inputs(184)) and (inputs(139)));
    layer0_outputs(7387) <= (inputs(161)) and not (inputs(14));
    layer0_outputs(7388) <= inputs(120);
    layer0_outputs(7389) <= not(inputs(230));
    layer0_outputs(7390) <= not(inputs(218));
    layer0_outputs(7391) <= (inputs(236)) or (inputs(99));
    layer0_outputs(7392) <= '1';
    layer0_outputs(7393) <= not(inputs(155));
    layer0_outputs(7394) <= not((inputs(222)) xor (inputs(68)));
    layer0_outputs(7395) <= not(inputs(173));
    layer0_outputs(7396) <= (inputs(240)) or (inputs(125));
    layer0_outputs(7397) <= not(inputs(168)) or (inputs(216));
    layer0_outputs(7398) <= (inputs(149)) and not (inputs(160));
    layer0_outputs(7399) <= not(inputs(27));
    layer0_outputs(7400) <= not(inputs(99)) or (inputs(0));
    layer0_outputs(7401) <= not((inputs(3)) or (inputs(252)));
    layer0_outputs(7402) <= inputs(70);
    layer0_outputs(7403) <= not((inputs(57)) and (inputs(91)));
    layer0_outputs(7404) <= not((inputs(226)) xor (inputs(178)));
    layer0_outputs(7405) <= (inputs(74)) and not (inputs(209));
    layer0_outputs(7406) <= (inputs(46)) xor (inputs(43));
    layer0_outputs(7407) <= not(inputs(102));
    layer0_outputs(7408) <= (inputs(12)) or (inputs(111));
    layer0_outputs(7409) <= (inputs(81)) xor (inputs(136));
    layer0_outputs(7410) <= not((inputs(62)) xor (inputs(198)));
    layer0_outputs(7411) <= (inputs(112)) xor (inputs(40));
    layer0_outputs(7412) <= inputs(25);
    layer0_outputs(7413) <= (inputs(101)) and not (inputs(26));
    layer0_outputs(7414) <= (inputs(83)) xor (inputs(6));
    layer0_outputs(7415) <= (inputs(192)) and not (inputs(30));
    layer0_outputs(7416) <= not((inputs(18)) xor (inputs(76)));
    layer0_outputs(7417) <= (inputs(203)) and not (inputs(172));
    layer0_outputs(7418) <= not((inputs(30)) or (inputs(8)));
    layer0_outputs(7419) <= not(inputs(3));
    layer0_outputs(7420) <= not((inputs(81)) xor (inputs(166)));
    layer0_outputs(7421) <= not(inputs(244));
    layer0_outputs(7422) <= (inputs(38)) xor (inputs(13));
    layer0_outputs(7423) <= not((inputs(81)) xor (inputs(216)));
    layer0_outputs(7424) <= (inputs(176)) xor (inputs(243));
    layer0_outputs(7425) <= not(inputs(202));
    layer0_outputs(7426) <= not((inputs(51)) or (inputs(0)));
    layer0_outputs(7427) <= not((inputs(81)) and (inputs(85)));
    layer0_outputs(7428) <= (inputs(57)) and not (inputs(182));
    layer0_outputs(7429) <= not((inputs(183)) or (inputs(161)));
    layer0_outputs(7430) <= (inputs(149)) and not (inputs(159));
    layer0_outputs(7431) <= (inputs(169)) and (inputs(171));
    layer0_outputs(7432) <= inputs(128);
    layer0_outputs(7433) <= not((inputs(19)) xor (inputs(60)));
    layer0_outputs(7434) <= (inputs(201)) xor (inputs(238));
    layer0_outputs(7435) <= not((inputs(82)) or (inputs(139)));
    layer0_outputs(7436) <= '1';
    layer0_outputs(7437) <= (inputs(199)) and (inputs(106));
    layer0_outputs(7438) <= '1';
    layer0_outputs(7439) <= not((inputs(2)) xor (inputs(177)));
    layer0_outputs(7440) <= not(inputs(139));
    layer0_outputs(7441) <= not(inputs(16)) or (inputs(90));
    layer0_outputs(7442) <= inputs(23);
    layer0_outputs(7443) <= not(inputs(116)) or (inputs(50));
    layer0_outputs(7444) <= inputs(86);
    layer0_outputs(7445) <= not(inputs(189)) or (inputs(87));
    layer0_outputs(7446) <= not((inputs(195)) or (inputs(159)));
    layer0_outputs(7447) <= not((inputs(153)) or (inputs(64)));
    layer0_outputs(7448) <= not((inputs(126)) or (inputs(18)));
    layer0_outputs(7449) <= (inputs(121)) and not (inputs(103));
    layer0_outputs(7450) <= (inputs(237)) xor (inputs(151));
    layer0_outputs(7451) <= (inputs(4)) or (inputs(176));
    layer0_outputs(7452) <= not(inputs(38)) or (inputs(244));
    layer0_outputs(7453) <= not(inputs(176)) or (inputs(98));
    layer0_outputs(7454) <= not((inputs(69)) and (inputs(218)));
    layer0_outputs(7455) <= not(inputs(28)) or (inputs(185));
    layer0_outputs(7456) <= not((inputs(200)) or (inputs(235)));
    layer0_outputs(7457) <= '0';
    layer0_outputs(7458) <= (inputs(3)) and (inputs(15));
    layer0_outputs(7459) <= not(inputs(55));
    layer0_outputs(7460) <= not((inputs(7)) or (inputs(64)));
    layer0_outputs(7461) <= (inputs(144)) and not (inputs(142));
    layer0_outputs(7462) <= not(inputs(163));
    layer0_outputs(7463) <= (inputs(160)) or (inputs(15));
    layer0_outputs(7464) <= (inputs(57)) and not (inputs(45));
    layer0_outputs(7465) <= (inputs(45)) or (inputs(43));
    layer0_outputs(7466) <= inputs(40);
    layer0_outputs(7467) <= (inputs(231)) or (inputs(100));
    layer0_outputs(7468) <= not((inputs(236)) or (inputs(72)));
    layer0_outputs(7469) <= (inputs(70)) and not (inputs(41));
    layer0_outputs(7470) <= (inputs(60)) or (inputs(113));
    layer0_outputs(7471) <= not((inputs(152)) xor (inputs(176)));
    layer0_outputs(7472) <= (inputs(55)) xor (inputs(196));
    layer0_outputs(7473) <= not(inputs(246)) or (inputs(35));
    layer0_outputs(7474) <= (inputs(161)) and not (inputs(94));
    layer0_outputs(7475) <= not(inputs(228)) or (inputs(203));
    layer0_outputs(7476) <= not((inputs(87)) xor (inputs(16)));
    layer0_outputs(7477) <= (inputs(252)) and not (inputs(66));
    layer0_outputs(7478) <= not(inputs(241)) or (inputs(33));
    layer0_outputs(7479) <= (inputs(101)) xor (inputs(56));
    layer0_outputs(7480) <= not(inputs(90));
    layer0_outputs(7481) <= not((inputs(193)) or (inputs(189)));
    layer0_outputs(7482) <= (inputs(52)) or (inputs(48));
    layer0_outputs(7483) <= not((inputs(116)) or (inputs(37)));
    layer0_outputs(7484) <= (inputs(108)) or (inputs(27));
    layer0_outputs(7485) <= inputs(170);
    layer0_outputs(7486) <= not((inputs(25)) or (inputs(204)));
    layer0_outputs(7487) <= (inputs(128)) xor (inputs(138));
    layer0_outputs(7488) <= inputs(199);
    layer0_outputs(7489) <= '1';
    layer0_outputs(7490) <= '1';
    layer0_outputs(7491) <= (inputs(42)) or (inputs(220));
    layer0_outputs(7492) <= inputs(167);
    layer0_outputs(7493) <= not(inputs(179)) or (inputs(97));
    layer0_outputs(7494) <= not((inputs(66)) and (inputs(208)));
    layer0_outputs(7495) <= not(inputs(58));
    layer0_outputs(7496) <= not(inputs(252));
    layer0_outputs(7497) <= inputs(197);
    layer0_outputs(7498) <= (inputs(4)) and not (inputs(62));
    layer0_outputs(7499) <= not((inputs(40)) or (inputs(23)));
    layer0_outputs(7500) <= (inputs(215)) or (inputs(65));
    layer0_outputs(7501) <= not(inputs(218));
    layer0_outputs(7502) <= not(inputs(184)) or (inputs(214));
    layer0_outputs(7503) <= not(inputs(162)) or (inputs(228));
    layer0_outputs(7504) <= (inputs(209)) xor (inputs(136));
    layer0_outputs(7505) <= not((inputs(141)) xor (inputs(38)));
    layer0_outputs(7506) <= not((inputs(170)) xor (inputs(137)));
    layer0_outputs(7507) <= (inputs(231)) and not (inputs(11));
    layer0_outputs(7508) <= inputs(198);
    layer0_outputs(7509) <= (inputs(205)) or (inputs(226));
    layer0_outputs(7510) <= not(inputs(196));
    layer0_outputs(7511) <= not((inputs(241)) xor (inputs(207)));
    layer0_outputs(7512) <= (inputs(153)) xor (inputs(112));
    layer0_outputs(7513) <= not(inputs(152)) or (inputs(67));
    layer0_outputs(7514) <= (inputs(73)) xor (inputs(192));
    layer0_outputs(7515) <= (inputs(216)) or (inputs(194));
    layer0_outputs(7516) <= inputs(253);
    layer0_outputs(7517) <= not(inputs(63)) or (inputs(65));
    layer0_outputs(7518) <= not((inputs(78)) or (inputs(216)));
    layer0_outputs(7519) <= not(inputs(100));
    layer0_outputs(7520) <= (inputs(149)) xor (inputs(193));
    layer0_outputs(7521) <= (inputs(24)) or (inputs(153));
    layer0_outputs(7522) <= not((inputs(188)) and (inputs(176)));
    layer0_outputs(7523) <= '0';
    layer0_outputs(7524) <= not((inputs(229)) or (inputs(248)));
    layer0_outputs(7525) <= (inputs(114)) or (inputs(116));
    layer0_outputs(7526) <= not((inputs(69)) and (inputs(106)));
    layer0_outputs(7527) <= not(inputs(55)) or (inputs(123));
    layer0_outputs(7528) <= not((inputs(78)) xor (inputs(216)));
    layer0_outputs(7529) <= inputs(79);
    layer0_outputs(7530) <= not(inputs(15));
    layer0_outputs(7531) <= (inputs(7)) or (inputs(193));
    layer0_outputs(7532) <= not(inputs(48)) or (inputs(112));
    layer0_outputs(7533) <= not(inputs(195));
    layer0_outputs(7534) <= not(inputs(120));
    layer0_outputs(7535) <= inputs(34);
    layer0_outputs(7536) <= (inputs(221)) and not (inputs(3));
    layer0_outputs(7537) <= not(inputs(140));
    layer0_outputs(7538) <= '1';
    layer0_outputs(7539) <= (inputs(183)) or (inputs(211));
    layer0_outputs(7540) <= not((inputs(71)) or (inputs(74)));
    layer0_outputs(7541) <= (inputs(249)) or (inputs(84));
    layer0_outputs(7542) <= not((inputs(81)) xor (inputs(45)));
    layer0_outputs(7543) <= (inputs(149)) and not (inputs(62));
    layer0_outputs(7544) <= (inputs(162)) and (inputs(245));
    layer0_outputs(7545) <= not((inputs(0)) xor (inputs(50)));
    layer0_outputs(7546) <= (inputs(43)) and (inputs(70));
    layer0_outputs(7547) <= inputs(170);
    layer0_outputs(7548) <= not(inputs(180)) or (inputs(144));
    layer0_outputs(7549) <= inputs(250);
    layer0_outputs(7550) <= (inputs(168)) and not (inputs(252));
    layer0_outputs(7551) <= (inputs(38)) or (inputs(194));
    layer0_outputs(7552) <= (inputs(187)) or (inputs(160));
    layer0_outputs(7553) <= not((inputs(118)) xor (inputs(43)));
    layer0_outputs(7554) <= not(inputs(77));
    layer0_outputs(7555) <= inputs(125);
    layer0_outputs(7556) <= (inputs(36)) and not (inputs(210));
    layer0_outputs(7557) <= not(inputs(52));
    layer0_outputs(7558) <= (inputs(71)) and not (inputs(6));
    layer0_outputs(7559) <= not(inputs(16));
    layer0_outputs(7560) <= not(inputs(52));
    layer0_outputs(7561) <= (inputs(181)) xor (inputs(242));
    layer0_outputs(7562) <= inputs(121);
    layer0_outputs(7563) <= inputs(148);
    layer0_outputs(7564) <= not(inputs(85));
    layer0_outputs(7565) <= (inputs(81)) or (inputs(228));
    layer0_outputs(7566) <= (inputs(21)) or (inputs(202));
    layer0_outputs(7567) <= not((inputs(184)) xor (inputs(192)));
    layer0_outputs(7568) <= not(inputs(23)) or (inputs(238));
    layer0_outputs(7569) <= (inputs(176)) and not (inputs(144));
    layer0_outputs(7570) <= inputs(255);
    layer0_outputs(7571) <= not(inputs(133));
    layer0_outputs(7572) <= '0';
    layer0_outputs(7573) <= '1';
    layer0_outputs(7574) <= (inputs(209)) and not (inputs(144));
    layer0_outputs(7575) <= not((inputs(144)) xor (inputs(31)));
    layer0_outputs(7576) <= (inputs(30)) xor (inputs(71));
    layer0_outputs(7577) <= inputs(85);
    layer0_outputs(7578) <= inputs(118);
    layer0_outputs(7579) <= (inputs(38)) xor (inputs(135));
    layer0_outputs(7580) <= (inputs(207)) xor (inputs(107));
    layer0_outputs(7581) <= inputs(108);
    layer0_outputs(7582) <= not((inputs(64)) or (inputs(166)));
    layer0_outputs(7583) <= not((inputs(190)) or (inputs(52)));
    layer0_outputs(7584) <= not((inputs(56)) or (inputs(188)));
    layer0_outputs(7585) <= (inputs(112)) xor (inputs(153));
    layer0_outputs(7586) <= '0';
    layer0_outputs(7587) <= not(inputs(146));
    layer0_outputs(7588) <= (inputs(236)) and not (inputs(228));
    layer0_outputs(7589) <= inputs(91);
    layer0_outputs(7590) <= (inputs(1)) xor (inputs(150));
    layer0_outputs(7591) <= (inputs(180)) or (inputs(202));
    layer0_outputs(7592) <= not((inputs(206)) and (inputs(63)));
    layer0_outputs(7593) <= not(inputs(175)) or (inputs(65));
    layer0_outputs(7594) <= not((inputs(45)) or (inputs(217)));
    layer0_outputs(7595) <= (inputs(33)) and not (inputs(20));
    layer0_outputs(7596) <= inputs(61);
    layer0_outputs(7597) <= inputs(25);
    layer0_outputs(7598) <= not(inputs(32)) or (inputs(49));
    layer0_outputs(7599) <= (inputs(46)) xor (inputs(212));
    layer0_outputs(7600) <= inputs(106);
    layer0_outputs(7601) <= not((inputs(35)) xor (inputs(169)));
    layer0_outputs(7602) <= not((inputs(35)) and (inputs(32)));
    layer0_outputs(7603) <= inputs(116);
    layer0_outputs(7604) <= (inputs(187)) and not (inputs(213));
    layer0_outputs(7605) <= (inputs(63)) xor (inputs(105));
    layer0_outputs(7606) <= not((inputs(123)) xor (inputs(105)));
    layer0_outputs(7607) <= not(inputs(165));
    layer0_outputs(7608) <= not((inputs(230)) or (inputs(234)));
    layer0_outputs(7609) <= inputs(181);
    layer0_outputs(7610) <= not(inputs(170)) or (inputs(28));
    layer0_outputs(7611) <= (inputs(225)) and not (inputs(9));
    layer0_outputs(7612) <= not(inputs(196));
    layer0_outputs(7613) <= not((inputs(128)) xor (inputs(158)));
    layer0_outputs(7614) <= not(inputs(85));
    layer0_outputs(7615) <= not((inputs(213)) or (inputs(80)));
    layer0_outputs(7616) <= (inputs(93)) or (inputs(126));
    layer0_outputs(7617) <= not(inputs(132)) or (inputs(194));
    layer0_outputs(7618) <= (inputs(198)) xor (inputs(214));
    layer0_outputs(7619) <= not((inputs(217)) xor (inputs(182)));
    layer0_outputs(7620) <= inputs(212);
    layer0_outputs(7621) <= inputs(165);
    layer0_outputs(7622) <= '1';
    layer0_outputs(7623) <= (inputs(27)) or (inputs(15));
    layer0_outputs(7624) <= inputs(241);
    layer0_outputs(7625) <= (inputs(248)) or (inputs(64));
    layer0_outputs(7626) <= not(inputs(116)) or (inputs(38));
    layer0_outputs(7627) <= inputs(166);
    layer0_outputs(7628) <= (inputs(101)) or (inputs(140));
    layer0_outputs(7629) <= not((inputs(36)) xor (inputs(83)));
    layer0_outputs(7630) <= not((inputs(15)) and (inputs(191)));
    layer0_outputs(7631) <= inputs(16);
    layer0_outputs(7632) <= inputs(120);
    layer0_outputs(7633) <= not((inputs(152)) xor (inputs(169)));
    layer0_outputs(7634) <= not(inputs(66));
    layer0_outputs(7635) <= not(inputs(25));
    layer0_outputs(7636) <= not(inputs(117)) or (inputs(154));
    layer0_outputs(7637) <= not((inputs(37)) or (inputs(94)));
    layer0_outputs(7638) <= not((inputs(42)) or (inputs(187)));
    layer0_outputs(7639) <= inputs(115);
    layer0_outputs(7640) <= '1';
    layer0_outputs(7641) <= (inputs(159)) xor (inputs(137));
    layer0_outputs(7642) <= '0';
    layer0_outputs(7643) <= not(inputs(179)) or (inputs(63));
    layer0_outputs(7644) <= not((inputs(234)) or (inputs(13)));
    layer0_outputs(7645) <= not(inputs(120));
    layer0_outputs(7646) <= '1';
    layer0_outputs(7647) <= (inputs(117)) xor (inputs(244));
    layer0_outputs(7648) <= (inputs(145)) xor (inputs(232));
    layer0_outputs(7649) <= (inputs(215)) and not (inputs(21));
    layer0_outputs(7650) <= not(inputs(219)) or (inputs(95));
    layer0_outputs(7651) <= not((inputs(131)) or (inputs(17)));
    layer0_outputs(7652) <= not((inputs(208)) xor (inputs(2)));
    layer0_outputs(7653) <= inputs(228);
    layer0_outputs(7654) <= (inputs(42)) xor (inputs(2));
    layer0_outputs(7655) <= not(inputs(111));
    layer0_outputs(7656) <= not(inputs(196));
    layer0_outputs(7657) <= not((inputs(138)) xor (inputs(37)));
    layer0_outputs(7658) <= (inputs(158)) xor (inputs(60));
    layer0_outputs(7659) <= not((inputs(226)) xor (inputs(45)));
    layer0_outputs(7660) <= inputs(24);
    layer0_outputs(7661) <= not(inputs(204)) or (inputs(35));
    layer0_outputs(7662) <= (inputs(186)) xor (inputs(9));
    layer0_outputs(7663) <= not(inputs(135));
    layer0_outputs(7664) <= not(inputs(230));
    layer0_outputs(7665) <= inputs(56);
    layer0_outputs(7666) <= '1';
    layer0_outputs(7667) <= not(inputs(90));
    layer0_outputs(7668) <= inputs(132);
    layer0_outputs(7669) <= not(inputs(120)) or (inputs(174));
    layer0_outputs(7670) <= (inputs(200)) or (inputs(30));
    layer0_outputs(7671) <= not(inputs(229)) or (inputs(3));
    layer0_outputs(7672) <= (inputs(158)) xor (inputs(155));
    layer0_outputs(7673) <= not((inputs(84)) xor (inputs(108)));
    layer0_outputs(7674) <= not((inputs(59)) xor (inputs(186)));
    layer0_outputs(7675) <= not(inputs(100));
    layer0_outputs(7676) <= not((inputs(3)) xor (inputs(60)));
    layer0_outputs(7677) <= (inputs(171)) and not (inputs(77));
    layer0_outputs(7678) <= not(inputs(208)) or (inputs(65));
    layer0_outputs(7679) <= not(inputs(105)) or (inputs(157));
    layer0_outputs(7680) <= not(inputs(12)) or (inputs(128));
    layer0_outputs(7681) <= (inputs(182)) and not (inputs(228));
    layer0_outputs(7682) <= not(inputs(87)) or (inputs(165));
    layer0_outputs(7683) <= not(inputs(203)) or (inputs(1));
    layer0_outputs(7684) <= not(inputs(197));
    layer0_outputs(7685) <= (inputs(160)) and not (inputs(155));
    layer0_outputs(7686) <= not((inputs(219)) and (inputs(51)));
    layer0_outputs(7687) <= not((inputs(109)) or (inputs(170)));
    layer0_outputs(7688) <= inputs(228);
    layer0_outputs(7689) <= not((inputs(71)) or (inputs(120)));
    layer0_outputs(7690) <= '1';
    layer0_outputs(7691) <= not((inputs(28)) or (inputs(242)));
    layer0_outputs(7692) <= (inputs(84)) xor (inputs(114));
    layer0_outputs(7693) <= inputs(168);
    layer0_outputs(7694) <= not((inputs(62)) xor (inputs(26)));
    layer0_outputs(7695) <= not(inputs(160)) or (inputs(18));
    layer0_outputs(7696) <= (inputs(48)) or (inputs(23));
    layer0_outputs(7697) <= '0';
    layer0_outputs(7698) <= (inputs(119)) and not (inputs(143));
    layer0_outputs(7699) <= not(inputs(165));
    layer0_outputs(7700) <= not(inputs(17));
    layer0_outputs(7701) <= not(inputs(174));
    layer0_outputs(7702) <= not(inputs(181));
    layer0_outputs(7703) <= not((inputs(170)) xor (inputs(203)));
    layer0_outputs(7704) <= (inputs(5)) or (inputs(156));
    layer0_outputs(7705) <= not((inputs(83)) or (inputs(9)));
    layer0_outputs(7706) <= not((inputs(254)) xor (inputs(24)));
    layer0_outputs(7707) <= (inputs(11)) and not (inputs(246));
    layer0_outputs(7708) <= (inputs(33)) or (inputs(78));
    layer0_outputs(7709) <= not((inputs(36)) or (inputs(182)));
    layer0_outputs(7710) <= (inputs(135)) xor (inputs(34));
    layer0_outputs(7711) <= (inputs(172)) or (inputs(82));
    layer0_outputs(7712) <= inputs(64);
    layer0_outputs(7713) <= not((inputs(7)) xor (inputs(102)));
    layer0_outputs(7714) <= (inputs(211)) or (inputs(228));
    layer0_outputs(7715) <= inputs(122);
    layer0_outputs(7716) <= inputs(77);
    layer0_outputs(7717) <= (inputs(14)) and not (inputs(47));
    layer0_outputs(7718) <= not(inputs(208));
    layer0_outputs(7719) <= inputs(10);
    layer0_outputs(7720) <= not((inputs(2)) and (inputs(170)));
    layer0_outputs(7721) <= not(inputs(214));
    layer0_outputs(7722) <= '1';
    layer0_outputs(7723) <= not(inputs(165)) or (inputs(236));
    layer0_outputs(7724) <= inputs(120);
    layer0_outputs(7725) <= not((inputs(158)) or (inputs(157)));
    layer0_outputs(7726) <= (inputs(8)) and not (inputs(144));
    layer0_outputs(7727) <= not((inputs(90)) or (inputs(164)));
    layer0_outputs(7728) <= (inputs(197)) or (inputs(222));
    layer0_outputs(7729) <= not((inputs(142)) xor (inputs(105)));
    layer0_outputs(7730) <= not(inputs(198)) or (inputs(144));
    layer0_outputs(7731) <= '1';
    layer0_outputs(7732) <= not((inputs(159)) or (inputs(231)));
    layer0_outputs(7733) <= (inputs(87)) and not (inputs(176));
    layer0_outputs(7734) <= '1';
    layer0_outputs(7735) <= (inputs(114)) xor (inputs(197));
    layer0_outputs(7736) <= not((inputs(208)) xor (inputs(187)));
    layer0_outputs(7737) <= (inputs(140)) and not (inputs(143));
    layer0_outputs(7738) <= (inputs(180)) and not (inputs(150));
    layer0_outputs(7739) <= not(inputs(173));
    layer0_outputs(7740) <= (inputs(194)) or (inputs(204));
    layer0_outputs(7741) <= not(inputs(102));
    layer0_outputs(7742) <= not(inputs(139)) or (inputs(241));
    layer0_outputs(7743) <= not(inputs(70)) or (inputs(163));
    layer0_outputs(7744) <= inputs(175);
    layer0_outputs(7745) <= not((inputs(174)) or (inputs(201)));
    layer0_outputs(7746) <= (inputs(92)) and not (inputs(240));
    layer0_outputs(7747) <= (inputs(226)) xor (inputs(13));
    layer0_outputs(7748) <= (inputs(208)) or (inputs(122));
    layer0_outputs(7749) <= not(inputs(120));
    layer0_outputs(7750) <= (inputs(100)) or (inputs(145));
    layer0_outputs(7751) <= (inputs(168)) or (inputs(150));
    layer0_outputs(7752) <= not((inputs(247)) xor (inputs(70)));
    layer0_outputs(7753) <= inputs(180);
    layer0_outputs(7754) <= not((inputs(19)) xor (inputs(103)));
    layer0_outputs(7755) <= not(inputs(237)) or (inputs(11));
    layer0_outputs(7756) <= inputs(177);
    layer0_outputs(7757) <= inputs(28);
    layer0_outputs(7758) <= '0';
    layer0_outputs(7759) <= (inputs(106)) and not (inputs(186));
    layer0_outputs(7760) <= (inputs(186)) xor (inputs(33));
    layer0_outputs(7761) <= inputs(145);
    layer0_outputs(7762) <= (inputs(193)) or (inputs(237));
    layer0_outputs(7763) <= not((inputs(182)) or (inputs(36)));
    layer0_outputs(7764) <= not(inputs(94)) or (inputs(219));
    layer0_outputs(7765) <= not((inputs(232)) or (inputs(251)));
    layer0_outputs(7766) <= not((inputs(206)) or (inputs(87)));
    layer0_outputs(7767) <= (inputs(186)) xor (inputs(5));
    layer0_outputs(7768) <= (inputs(104)) xor (inputs(145));
    layer0_outputs(7769) <= inputs(94);
    layer0_outputs(7770) <= (inputs(25)) xor (inputs(67));
    layer0_outputs(7771) <= not(inputs(16));
    layer0_outputs(7772) <= (inputs(138)) or (inputs(177));
    layer0_outputs(7773) <= not((inputs(68)) and (inputs(175)));
    layer0_outputs(7774) <= (inputs(208)) and not (inputs(237));
    layer0_outputs(7775) <= (inputs(20)) and (inputs(35));
    layer0_outputs(7776) <= (inputs(36)) or (inputs(185));
    layer0_outputs(7777) <= not(inputs(83)) or (inputs(216));
    layer0_outputs(7778) <= inputs(61);
    layer0_outputs(7779) <= not(inputs(76));
    layer0_outputs(7780) <= not(inputs(93));
    layer0_outputs(7781) <= not(inputs(126));
    layer0_outputs(7782) <= (inputs(247)) and not (inputs(250));
    layer0_outputs(7783) <= not((inputs(124)) or (inputs(98)));
    layer0_outputs(7784) <= (inputs(77)) and not (inputs(228));
    layer0_outputs(7785) <= inputs(71);
    layer0_outputs(7786) <= (inputs(62)) or (inputs(149));
    layer0_outputs(7787) <= (inputs(225)) or (inputs(151));
    layer0_outputs(7788) <= not(inputs(182)) or (inputs(130));
    layer0_outputs(7789) <= not(inputs(75)) or (inputs(46));
    layer0_outputs(7790) <= (inputs(59)) xor (inputs(32));
    layer0_outputs(7791) <= (inputs(136)) and not (inputs(163));
    layer0_outputs(7792) <= (inputs(94)) and not (inputs(141));
    layer0_outputs(7793) <= inputs(139);
    layer0_outputs(7794) <= inputs(215);
    layer0_outputs(7795) <= (inputs(68)) xor (inputs(232));
    layer0_outputs(7796) <= inputs(221);
    layer0_outputs(7797) <= (inputs(160)) xor (inputs(88));
    layer0_outputs(7798) <= inputs(207);
    layer0_outputs(7799) <= not((inputs(251)) xor (inputs(168)));
    layer0_outputs(7800) <= (inputs(144)) xor (inputs(233));
    layer0_outputs(7801) <= not((inputs(183)) xor (inputs(184)));
    layer0_outputs(7802) <= (inputs(67)) and not (inputs(206));
    layer0_outputs(7803) <= (inputs(162)) and not (inputs(225));
    layer0_outputs(7804) <= inputs(36);
    layer0_outputs(7805) <= (inputs(157)) and not (inputs(157));
    layer0_outputs(7806) <= (inputs(137)) xor (inputs(28));
    layer0_outputs(7807) <= not(inputs(241));
    layer0_outputs(7808) <= (inputs(167)) and not (inputs(234));
    layer0_outputs(7809) <= not(inputs(128)) or (inputs(178));
    layer0_outputs(7810) <= not(inputs(195)) or (inputs(82));
    layer0_outputs(7811) <= (inputs(99)) or (inputs(100));
    layer0_outputs(7812) <= not(inputs(214));
    layer0_outputs(7813) <= not(inputs(21)) or (inputs(244));
    layer0_outputs(7814) <= inputs(60);
    layer0_outputs(7815) <= (inputs(204)) and not (inputs(63));
    layer0_outputs(7816) <= not((inputs(53)) xor (inputs(65)));
    layer0_outputs(7817) <= not(inputs(7));
    layer0_outputs(7818) <= not((inputs(140)) or (inputs(201)));
    layer0_outputs(7819) <= not((inputs(38)) xor (inputs(113)));
    layer0_outputs(7820) <= not((inputs(153)) xor (inputs(26)));
    layer0_outputs(7821) <= not((inputs(34)) or (inputs(181)));
    layer0_outputs(7822) <= (inputs(86)) and not (inputs(68));
    layer0_outputs(7823) <= not((inputs(30)) or (inputs(181)));
    layer0_outputs(7824) <= not(inputs(176));
    layer0_outputs(7825) <= not((inputs(92)) or (inputs(170)));
    layer0_outputs(7826) <= (inputs(114)) or (inputs(15));
    layer0_outputs(7827) <= not(inputs(229)) or (inputs(80));
    layer0_outputs(7828) <= (inputs(11)) xor (inputs(77));
    layer0_outputs(7829) <= (inputs(126)) and not (inputs(160));
    layer0_outputs(7830) <= not(inputs(149));
    layer0_outputs(7831) <= not(inputs(218));
    layer0_outputs(7832) <= not(inputs(250));
    layer0_outputs(7833) <= (inputs(79)) and not (inputs(127));
    layer0_outputs(7834) <= not((inputs(232)) and (inputs(228)));
    layer0_outputs(7835) <= not((inputs(216)) or (inputs(76)));
    layer0_outputs(7836) <= not((inputs(187)) xor (inputs(99)));
    layer0_outputs(7837) <= (inputs(28)) xor (inputs(244));
    layer0_outputs(7838) <= not(inputs(173)) or (inputs(130));
    layer0_outputs(7839) <= inputs(196);
    layer0_outputs(7840) <= inputs(149);
    layer0_outputs(7841) <= not(inputs(149));
    layer0_outputs(7842) <= not(inputs(50));
    layer0_outputs(7843) <= not((inputs(112)) or (inputs(90)));
    layer0_outputs(7844) <= not(inputs(158)) or (inputs(74));
    layer0_outputs(7845) <= not((inputs(188)) or (inputs(194)));
    layer0_outputs(7846) <= (inputs(117)) or (inputs(116));
    layer0_outputs(7847) <= not(inputs(231));
    layer0_outputs(7848) <= not((inputs(174)) or (inputs(152)));
    layer0_outputs(7849) <= not((inputs(253)) and (inputs(92)));
    layer0_outputs(7850) <= '0';
    layer0_outputs(7851) <= inputs(69);
    layer0_outputs(7852) <= not((inputs(219)) or (inputs(252)));
    layer0_outputs(7853) <= (inputs(207)) and not (inputs(4));
    layer0_outputs(7854) <= (inputs(60)) and (inputs(201));
    layer0_outputs(7855) <= (inputs(85)) and not (inputs(117));
    layer0_outputs(7856) <= (inputs(64)) and (inputs(255));
    layer0_outputs(7857) <= inputs(97);
    layer0_outputs(7858) <= (inputs(119)) or (inputs(165));
    layer0_outputs(7859) <= (inputs(239)) and not (inputs(204));
    layer0_outputs(7860) <= not(inputs(104));
    layer0_outputs(7861) <= not(inputs(210));
    layer0_outputs(7862) <= (inputs(182)) and not (inputs(195));
    layer0_outputs(7863) <= not((inputs(160)) xor (inputs(250)));
    layer0_outputs(7864) <= not(inputs(203)) or (inputs(226));
    layer0_outputs(7865) <= not(inputs(197)) or (inputs(204));
    layer0_outputs(7866) <= not((inputs(130)) or (inputs(205)));
    layer0_outputs(7867) <= not((inputs(40)) or (inputs(124)));
    layer0_outputs(7868) <= not((inputs(153)) or (inputs(137)));
    layer0_outputs(7869) <= (inputs(84)) and not (inputs(242));
    layer0_outputs(7870) <= not(inputs(136)) or (inputs(211));
    layer0_outputs(7871) <= not(inputs(203)) or (inputs(13));
    layer0_outputs(7872) <= '1';
    layer0_outputs(7873) <= not(inputs(187));
    layer0_outputs(7874) <= not((inputs(6)) and (inputs(145)));
    layer0_outputs(7875) <= (inputs(234)) xor (inputs(249));
    layer0_outputs(7876) <= (inputs(2)) xor (inputs(232));
    layer0_outputs(7877) <= inputs(55);
    layer0_outputs(7878) <= inputs(167);
    layer0_outputs(7879) <= (inputs(40)) or (inputs(207));
    layer0_outputs(7880) <= not(inputs(178));
    layer0_outputs(7881) <= (inputs(204)) and not (inputs(208));
    layer0_outputs(7882) <= not((inputs(41)) or (inputs(55)));
    layer0_outputs(7883) <= (inputs(15)) and (inputs(192));
    layer0_outputs(7884) <= (inputs(28)) and not (inputs(240));
    layer0_outputs(7885) <= not((inputs(149)) or (inputs(69)));
    layer0_outputs(7886) <= not(inputs(38));
    layer0_outputs(7887) <= not((inputs(185)) and (inputs(83)));
    layer0_outputs(7888) <= (inputs(89)) or (inputs(173));
    layer0_outputs(7889) <= (inputs(163)) or (inputs(137));
    layer0_outputs(7890) <= (inputs(49)) or (inputs(169));
    layer0_outputs(7891) <= inputs(57);
    layer0_outputs(7892) <= not((inputs(213)) or (inputs(134)));
    layer0_outputs(7893) <= (inputs(130)) or (inputs(207));
    layer0_outputs(7894) <= not((inputs(203)) or (inputs(70)));
    layer0_outputs(7895) <= (inputs(27)) or (inputs(125));
    layer0_outputs(7896) <= not(inputs(144));
    layer0_outputs(7897) <= not((inputs(185)) xor (inputs(113)));
    layer0_outputs(7898) <= '0';
    layer0_outputs(7899) <= not((inputs(27)) or (inputs(12)));
    layer0_outputs(7900) <= (inputs(19)) and (inputs(245));
    layer0_outputs(7901) <= not(inputs(122));
    layer0_outputs(7902) <= not(inputs(165));
    layer0_outputs(7903) <= '0';
    layer0_outputs(7904) <= not((inputs(44)) and (inputs(106)));
    layer0_outputs(7905) <= not(inputs(204)) or (inputs(211));
    layer0_outputs(7906) <= (inputs(31)) or (inputs(249));
    layer0_outputs(7907) <= not(inputs(6));
    layer0_outputs(7908) <= (inputs(157)) and not (inputs(33));
    layer0_outputs(7909) <= (inputs(80)) or (inputs(199));
    layer0_outputs(7910) <= not((inputs(82)) or (inputs(111)));
    layer0_outputs(7911) <= (inputs(30)) and (inputs(15));
    layer0_outputs(7912) <= (inputs(230)) xor (inputs(41));
    layer0_outputs(7913) <= inputs(136);
    layer0_outputs(7914) <= not(inputs(110));
    layer0_outputs(7915) <= not(inputs(148)) or (inputs(246));
    layer0_outputs(7916) <= (inputs(35)) xor (inputs(206));
    layer0_outputs(7917) <= not(inputs(58)) or (inputs(45));
    layer0_outputs(7918) <= (inputs(73)) or (inputs(244));
    layer0_outputs(7919) <= inputs(85);
    layer0_outputs(7920) <= (inputs(195)) and not (inputs(82));
    layer0_outputs(7921) <= '1';
    layer0_outputs(7922) <= not(inputs(162));
    layer0_outputs(7923) <= not(inputs(225));
    layer0_outputs(7924) <= (inputs(131)) or (inputs(132));
    layer0_outputs(7925) <= (inputs(172)) or (inputs(176));
    layer0_outputs(7926) <= not((inputs(177)) and (inputs(158)));
    layer0_outputs(7927) <= not(inputs(239)) or (inputs(224));
    layer0_outputs(7928) <= (inputs(185)) and not (inputs(98));
    layer0_outputs(7929) <= (inputs(207)) or (inputs(77));
    layer0_outputs(7930) <= not(inputs(28));
    layer0_outputs(7931) <= inputs(197);
    layer0_outputs(7932) <= inputs(96);
    layer0_outputs(7933) <= not(inputs(121)) or (inputs(125));
    layer0_outputs(7934) <= not((inputs(0)) or (inputs(71)));
    layer0_outputs(7935) <= (inputs(23)) xor (inputs(246));
    layer0_outputs(7936) <= not((inputs(57)) xor (inputs(142)));
    layer0_outputs(7937) <= not((inputs(225)) xor (inputs(99)));
    layer0_outputs(7938) <= not(inputs(81));
    layer0_outputs(7939) <= (inputs(154)) xor (inputs(187));
    layer0_outputs(7940) <= not(inputs(228));
    layer0_outputs(7941) <= (inputs(163)) or (inputs(239));
    layer0_outputs(7942) <= inputs(11);
    layer0_outputs(7943) <= not((inputs(163)) or (inputs(186)));
    layer0_outputs(7944) <= not(inputs(149)) or (inputs(159));
    layer0_outputs(7945) <= not((inputs(134)) xor (inputs(96)));
    layer0_outputs(7946) <= (inputs(141)) or (inputs(128));
    layer0_outputs(7947) <= (inputs(216)) or (inputs(170));
    layer0_outputs(7948) <= not((inputs(100)) or (inputs(90)));
    layer0_outputs(7949) <= not(inputs(70)) or (inputs(175));
    layer0_outputs(7950) <= not(inputs(3)) or (inputs(140));
    layer0_outputs(7951) <= not(inputs(81));
    layer0_outputs(7952) <= inputs(231);
    layer0_outputs(7953) <= (inputs(39)) and not (inputs(247));
    layer0_outputs(7954) <= (inputs(92)) and not (inputs(211));
    layer0_outputs(7955) <= not((inputs(13)) and (inputs(11)));
    layer0_outputs(7956) <= (inputs(115)) and not (inputs(112));
    layer0_outputs(7957) <= (inputs(213)) xor (inputs(140));
    layer0_outputs(7958) <= not((inputs(73)) xor (inputs(248)));
    layer0_outputs(7959) <= inputs(102);
    layer0_outputs(7960) <= (inputs(243)) and not (inputs(234));
    layer0_outputs(7961) <= (inputs(94)) and not (inputs(42));
    layer0_outputs(7962) <= (inputs(63)) and not (inputs(228));
    layer0_outputs(7963) <= '0';
    layer0_outputs(7964) <= '1';
    layer0_outputs(7965) <= not(inputs(106)) or (inputs(141));
    layer0_outputs(7966) <= not((inputs(125)) or (inputs(156)));
    layer0_outputs(7967) <= (inputs(212)) xor (inputs(203));
    layer0_outputs(7968) <= (inputs(154)) and not (inputs(5));
    layer0_outputs(7969) <= inputs(62);
    layer0_outputs(7970) <= not((inputs(111)) or (inputs(118)));
    layer0_outputs(7971) <= not(inputs(147));
    layer0_outputs(7972) <= not((inputs(161)) xor (inputs(123)));
    layer0_outputs(7973) <= not((inputs(64)) xor (inputs(194)));
    layer0_outputs(7974) <= not(inputs(56));
    layer0_outputs(7975) <= not((inputs(9)) or (inputs(255)));
    layer0_outputs(7976) <= (inputs(130)) or (inputs(116));
    layer0_outputs(7977) <= not(inputs(58)) or (inputs(244));
    layer0_outputs(7978) <= (inputs(145)) xor (inputs(91));
    layer0_outputs(7979) <= inputs(109);
    layer0_outputs(7980) <= (inputs(149)) or (inputs(210));
    layer0_outputs(7981) <= not(inputs(196));
    layer0_outputs(7982) <= not(inputs(205));
    layer0_outputs(7983) <= (inputs(173)) or (inputs(87));
    layer0_outputs(7984) <= (inputs(193)) or (inputs(8));
    layer0_outputs(7985) <= (inputs(76)) or (inputs(186));
    layer0_outputs(7986) <= inputs(121);
    layer0_outputs(7987) <= not(inputs(191));
    layer0_outputs(7988) <= not((inputs(224)) and (inputs(123)));
    layer0_outputs(7989) <= (inputs(31)) and not (inputs(17));
    layer0_outputs(7990) <= inputs(179);
    layer0_outputs(7991) <= not(inputs(165));
    layer0_outputs(7992) <= not((inputs(83)) or (inputs(112)));
    layer0_outputs(7993) <= (inputs(117)) or (inputs(161));
    layer0_outputs(7994) <= (inputs(197)) or (inputs(82));
    layer0_outputs(7995) <= not((inputs(228)) or (inputs(21)));
    layer0_outputs(7996) <= not((inputs(82)) or (inputs(123)));
    layer0_outputs(7997) <= (inputs(45)) or (inputs(255));
    layer0_outputs(7998) <= (inputs(85)) and not (inputs(211));
    layer0_outputs(7999) <= inputs(242);
    layer0_outputs(8000) <= (inputs(30)) or (inputs(53));
    layer0_outputs(8001) <= (inputs(2)) and not (inputs(63));
    layer0_outputs(8002) <= inputs(136);
    layer0_outputs(8003) <= (inputs(144)) and not (inputs(176));
    layer0_outputs(8004) <= not(inputs(119));
    layer0_outputs(8005) <= (inputs(238)) and (inputs(212));
    layer0_outputs(8006) <= (inputs(88)) and not (inputs(255));
    layer0_outputs(8007) <= (inputs(106)) or (inputs(229));
    layer0_outputs(8008) <= not((inputs(18)) xor (inputs(164)));
    layer0_outputs(8009) <= not(inputs(214)) or (inputs(105));
    layer0_outputs(8010) <= not(inputs(94));
    layer0_outputs(8011) <= not((inputs(250)) and (inputs(143)));
    layer0_outputs(8012) <= (inputs(53)) xor (inputs(70));
    layer0_outputs(8013) <= not((inputs(134)) or (inputs(220)));
    layer0_outputs(8014) <= (inputs(76)) and not (inputs(46));
    layer0_outputs(8015) <= not(inputs(36));
    layer0_outputs(8016) <= (inputs(152)) and not (inputs(160));
    layer0_outputs(8017) <= not(inputs(13)) or (inputs(0));
    layer0_outputs(8018) <= not((inputs(104)) or (inputs(0)));
    layer0_outputs(8019) <= '1';
    layer0_outputs(8020) <= inputs(18);
    layer0_outputs(8021) <= (inputs(32)) or (inputs(232));
    layer0_outputs(8022) <= (inputs(45)) and (inputs(235));
    layer0_outputs(8023) <= not((inputs(111)) or (inputs(43)));
    layer0_outputs(8024) <= not((inputs(155)) xor (inputs(254)));
    layer0_outputs(8025) <= not(inputs(179));
    layer0_outputs(8026) <= '0';
    layer0_outputs(8027) <= '0';
    layer0_outputs(8028) <= (inputs(155)) and not (inputs(246));
    layer0_outputs(8029) <= not((inputs(244)) xor (inputs(71)));
    layer0_outputs(8030) <= not(inputs(64));
    layer0_outputs(8031) <= inputs(155);
    layer0_outputs(8032) <= not((inputs(96)) and (inputs(201)));
    layer0_outputs(8033) <= (inputs(81)) xor (inputs(153));
    layer0_outputs(8034) <= (inputs(135)) and not (inputs(42));
    layer0_outputs(8035) <= (inputs(165)) or (inputs(217));
    layer0_outputs(8036) <= not(inputs(157));
    layer0_outputs(8037) <= (inputs(100)) xor (inputs(99));
    layer0_outputs(8038) <= not(inputs(38));
    layer0_outputs(8039) <= (inputs(69)) and not (inputs(52));
    layer0_outputs(8040) <= (inputs(178)) and not (inputs(97));
    layer0_outputs(8041) <= (inputs(60)) and not (inputs(36));
    layer0_outputs(8042) <= not(inputs(186));
    layer0_outputs(8043) <= (inputs(67)) and not (inputs(115));
    layer0_outputs(8044) <= (inputs(140)) or (inputs(109));
    layer0_outputs(8045) <= not((inputs(52)) xor (inputs(145)));
    layer0_outputs(8046) <= not(inputs(49));
    layer0_outputs(8047) <= (inputs(168)) or (inputs(67));
    layer0_outputs(8048) <= inputs(48);
    layer0_outputs(8049) <= not((inputs(250)) xor (inputs(255)));
    layer0_outputs(8050) <= (inputs(101)) and not (inputs(12));
    layer0_outputs(8051) <= (inputs(41)) and not (inputs(210));
    layer0_outputs(8052) <= not(inputs(172));
    layer0_outputs(8053) <= not(inputs(74)) or (inputs(193));
    layer0_outputs(8054) <= (inputs(15)) or (inputs(135));
    layer0_outputs(8055) <= '1';
    layer0_outputs(8056) <= not((inputs(246)) or (inputs(17)));
    layer0_outputs(8057) <= not((inputs(65)) and (inputs(115)));
    layer0_outputs(8058) <= (inputs(153)) xor (inputs(246));
    layer0_outputs(8059) <= not((inputs(194)) or (inputs(172)));
    layer0_outputs(8060) <= not(inputs(141));
    layer0_outputs(8061) <= (inputs(72)) or (inputs(196));
    layer0_outputs(8062) <= not((inputs(1)) or (inputs(77)));
    layer0_outputs(8063) <= not((inputs(17)) xor (inputs(160)));
    layer0_outputs(8064) <= (inputs(181)) and not (inputs(67));
    layer0_outputs(8065) <= inputs(88);
    layer0_outputs(8066) <= not(inputs(186)) or (inputs(42));
    layer0_outputs(8067) <= not(inputs(73)) or (inputs(240));
    layer0_outputs(8068) <= (inputs(160)) xor (inputs(186));
    layer0_outputs(8069) <= not((inputs(76)) xor (inputs(45)));
    layer0_outputs(8070) <= (inputs(15)) xor (inputs(148));
    layer0_outputs(8071) <= not((inputs(93)) or (inputs(36)));
    layer0_outputs(8072) <= not(inputs(57));
    layer0_outputs(8073) <= (inputs(124)) xor (inputs(142));
    layer0_outputs(8074) <= '1';
    layer0_outputs(8075) <= not((inputs(25)) or (inputs(153)));
    layer0_outputs(8076) <= not(inputs(69)) or (inputs(191));
    layer0_outputs(8077) <= (inputs(207)) or (inputs(207));
    layer0_outputs(8078) <= not(inputs(79));
    layer0_outputs(8079) <= (inputs(179)) xor (inputs(140));
    layer0_outputs(8080) <= not(inputs(183));
    layer0_outputs(8081) <= not((inputs(113)) or (inputs(158)));
    layer0_outputs(8082) <= (inputs(12)) or (inputs(138));
    layer0_outputs(8083) <= inputs(127);
    layer0_outputs(8084) <= not((inputs(139)) xor (inputs(37)));
    layer0_outputs(8085) <= inputs(135);
    layer0_outputs(8086) <= '0';
    layer0_outputs(8087) <= (inputs(128)) xor (inputs(89));
    layer0_outputs(8088) <= not((inputs(199)) or (inputs(68)));
    layer0_outputs(8089) <= not((inputs(151)) xor (inputs(125)));
    layer0_outputs(8090) <= (inputs(138)) and not (inputs(11));
    layer0_outputs(8091) <= (inputs(69)) xor (inputs(173));
    layer0_outputs(8092) <= not((inputs(248)) or (inputs(47)));
    layer0_outputs(8093) <= not(inputs(162));
    layer0_outputs(8094) <= not(inputs(71)) or (inputs(127));
    layer0_outputs(8095) <= inputs(232);
    layer0_outputs(8096) <= inputs(61);
    layer0_outputs(8097) <= not(inputs(178)) or (inputs(17));
    layer0_outputs(8098) <= inputs(222);
    layer0_outputs(8099) <= not((inputs(238)) xor (inputs(39)));
    layer0_outputs(8100) <= not((inputs(153)) or (inputs(36)));
    layer0_outputs(8101) <= not((inputs(70)) xor (inputs(98)));
    layer0_outputs(8102) <= (inputs(63)) or (inputs(229));
    layer0_outputs(8103) <= not(inputs(134));
    layer0_outputs(8104) <= (inputs(54)) and not (inputs(34));
    layer0_outputs(8105) <= not(inputs(99));
    layer0_outputs(8106) <= (inputs(247)) and (inputs(41));
    layer0_outputs(8107) <= (inputs(11)) and (inputs(15));
    layer0_outputs(8108) <= (inputs(72)) and (inputs(108));
    layer0_outputs(8109) <= (inputs(126)) and not (inputs(63));
    layer0_outputs(8110) <= not((inputs(63)) or (inputs(181)));
    layer0_outputs(8111) <= (inputs(176)) or (inputs(195));
    layer0_outputs(8112) <= inputs(177);
    layer0_outputs(8113) <= (inputs(10)) xor (inputs(140));
    layer0_outputs(8114) <= inputs(230);
    layer0_outputs(8115) <= inputs(219);
    layer0_outputs(8116) <= '1';
    layer0_outputs(8117) <= (inputs(63)) or (inputs(65));
    layer0_outputs(8118) <= not(inputs(164)) or (inputs(230));
    layer0_outputs(8119) <= not(inputs(169));
    layer0_outputs(8120) <= (inputs(122)) xor (inputs(32));
    layer0_outputs(8121) <= inputs(101);
    layer0_outputs(8122) <= not((inputs(87)) or (inputs(229)));
    layer0_outputs(8123) <= not((inputs(127)) or (inputs(201)));
    layer0_outputs(8124) <= not((inputs(241)) and (inputs(223)));
    layer0_outputs(8125) <= (inputs(18)) and (inputs(230));
    layer0_outputs(8126) <= not((inputs(189)) or (inputs(163)));
    layer0_outputs(8127) <= (inputs(109)) xor (inputs(205));
    layer0_outputs(8128) <= not((inputs(45)) xor (inputs(237)));
    layer0_outputs(8129) <= not(inputs(72));
    layer0_outputs(8130) <= not(inputs(137)) or (inputs(253));
    layer0_outputs(8131) <= '1';
    layer0_outputs(8132) <= not((inputs(241)) xor (inputs(214)));
    layer0_outputs(8133) <= (inputs(25)) and not (inputs(212));
    layer0_outputs(8134) <= not((inputs(31)) or (inputs(135)));
    layer0_outputs(8135) <= (inputs(118)) and not (inputs(89));
    layer0_outputs(8136) <= not(inputs(148)) or (inputs(22));
    layer0_outputs(8137) <= (inputs(52)) or (inputs(222));
    layer0_outputs(8138) <= inputs(211);
    layer0_outputs(8139) <= not(inputs(3)) or (inputs(5));
    layer0_outputs(8140) <= not((inputs(144)) and (inputs(232)));
    layer0_outputs(8141) <= (inputs(142)) or (inputs(150));
    layer0_outputs(8142) <= (inputs(108)) xor (inputs(97));
    layer0_outputs(8143) <= (inputs(217)) xor (inputs(48));
    layer0_outputs(8144) <= not(inputs(249)) or (inputs(27));
    layer0_outputs(8145) <= (inputs(33)) xor (inputs(69));
    layer0_outputs(8146) <= not(inputs(149)) or (inputs(189));
    layer0_outputs(8147) <= (inputs(231)) and not (inputs(236));
    layer0_outputs(8148) <= (inputs(124)) or (inputs(245));
    layer0_outputs(8149) <= not(inputs(183)) or (inputs(228));
    layer0_outputs(8150) <= (inputs(235)) or (inputs(148));
    layer0_outputs(8151) <= not((inputs(10)) or (inputs(31)));
    layer0_outputs(8152) <= (inputs(179)) or (inputs(203));
    layer0_outputs(8153) <= not(inputs(214)) or (inputs(93));
    layer0_outputs(8154) <= not(inputs(228)) or (inputs(126));
    layer0_outputs(8155) <= not((inputs(113)) and (inputs(1)));
    layer0_outputs(8156) <= not(inputs(106));
    layer0_outputs(8157) <= not((inputs(203)) or (inputs(123)));
    layer0_outputs(8158) <= not(inputs(135));
    layer0_outputs(8159) <= inputs(118);
    layer0_outputs(8160) <= not(inputs(75)) or (inputs(45));
    layer0_outputs(8161) <= '1';
    layer0_outputs(8162) <= not(inputs(137)) or (inputs(231));
    layer0_outputs(8163) <= (inputs(151)) or (inputs(27));
    layer0_outputs(8164) <= inputs(156);
    layer0_outputs(8165) <= not((inputs(223)) or (inputs(88)));
    layer0_outputs(8166) <= '0';
    layer0_outputs(8167) <= (inputs(71)) and not (inputs(23));
    layer0_outputs(8168) <= '0';
    layer0_outputs(8169) <= (inputs(143)) or (inputs(182));
    layer0_outputs(8170) <= '0';
    layer0_outputs(8171) <= (inputs(165)) xor (inputs(110));
    layer0_outputs(8172) <= not(inputs(126)) or (inputs(222));
    layer0_outputs(8173) <= not(inputs(120));
    layer0_outputs(8174) <= '0';
    layer0_outputs(8175) <= inputs(228);
    layer0_outputs(8176) <= '1';
    layer0_outputs(8177) <= (inputs(240)) and not (inputs(175));
    layer0_outputs(8178) <= inputs(67);
    layer0_outputs(8179) <= not(inputs(138));
    layer0_outputs(8180) <= not(inputs(149));
    layer0_outputs(8181) <= not(inputs(251)) or (inputs(224));
    layer0_outputs(8182) <= (inputs(149)) or (inputs(107));
    layer0_outputs(8183) <= (inputs(129)) or (inputs(63));
    layer0_outputs(8184) <= not((inputs(93)) or (inputs(213)));
    layer0_outputs(8185) <= not((inputs(181)) xor (inputs(27)));
    layer0_outputs(8186) <= not((inputs(19)) and (inputs(38)));
    layer0_outputs(8187) <= not(inputs(249));
    layer0_outputs(8188) <= inputs(82);
    layer0_outputs(8189) <= (inputs(84)) or (inputs(175));
    layer0_outputs(8190) <= not(inputs(53)) or (inputs(247));
    layer0_outputs(8191) <= (inputs(228)) or (inputs(132));
    layer0_outputs(8192) <= not((inputs(230)) xor (inputs(16)));
    layer0_outputs(8193) <= inputs(255);
    layer0_outputs(8194) <= not(inputs(81));
    layer0_outputs(8195) <= not(inputs(33)) or (inputs(33));
    layer0_outputs(8196) <= inputs(180);
    layer0_outputs(8197) <= not((inputs(136)) or (inputs(32)));
    layer0_outputs(8198) <= not((inputs(72)) xor (inputs(161)));
    layer0_outputs(8199) <= (inputs(227)) and (inputs(110));
    layer0_outputs(8200) <= not((inputs(90)) xor (inputs(248)));
    layer0_outputs(8201) <= (inputs(195)) and (inputs(162));
    layer0_outputs(8202) <= (inputs(32)) and (inputs(254));
    layer0_outputs(8203) <= inputs(86);
    layer0_outputs(8204) <= (inputs(179)) xor (inputs(150));
    layer0_outputs(8205) <= (inputs(251)) or (inputs(70));
    layer0_outputs(8206) <= not(inputs(209));
    layer0_outputs(8207) <= (inputs(217)) and not (inputs(97));
    layer0_outputs(8208) <= not(inputs(77));
    layer0_outputs(8209) <= '1';
    layer0_outputs(8210) <= not((inputs(92)) xor (inputs(71)));
    layer0_outputs(8211) <= not((inputs(215)) xor (inputs(170)));
    layer0_outputs(8212) <= inputs(79);
    layer0_outputs(8213) <= (inputs(133)) and not (inputs(50));
    layer0_outputs(8214) <= not(inputs(100));
    layer0_outputs(8215) <= not((inputs(49)) xor (inputs(69)));
    layer0_outputs(8216) <= '0';
    layer0_outputs(8217) <= not(inputs(88));
    layer0_outputs(8218) <= (inputs(141)) or (inputs(250));
    layer0_outputs(8219) <= not((inputs(2)) xor (inputs(255)));
    layer0_outputs(8220) <= (inputs(227)) and not (inputs(95));
    layer0_outputs(8221) <= (inputs(2)) and (inputs(217));
    layer0_outputs(8222) <= inputs(144);
    layer0_outputs(8223) <= not(inputs(169)) or (inputs(49));
    layer0_outputs(8224) <= not((inputs(185)) or (inputs(201)));
    layer0_outputs(8225) <= (inputs(5)) xor (inputs(101));
    layer0_outputs(8226) <= '0';
    layer0_outputs(8227) <= not((inputs(111)) and (inputs(4)));
    layer0_outputs(8228) <= not(inputs(254));
    layer0_outputs(8229) <= (inputs(240)) and not (inputs(63));
    layer0_outputs(8230) <= inputs(88);
    layer0_outputs(8231) <= not(inputs(133)) or (inputs(141));
    layer0_outputs(8232) <= (inputs(48)) and not (inputs(65));
    layer0_outputs(8233) <= (inputs(138)) and not (inputs(251));
    layer0_outputs(8234) <= not(inputs(234));
    layer0_outputs(8235) <= not(inputs(105));
    layer0_outputs(8236) <= '1';
    layer0_outputs(8237) <= not((inputs(99)) xor (inputs(228)));
    layer0_outputs(8238) <= not((inputs(225)) or (inputs(253)));
    layer0_outputs(8239) <= not(inputs(24));
    layer0_outputs(8240) <= (inputs(222)) or (inputs(116));
    layer0_outputs(8241) <= (inputs(119)) and not (inputs(19));
    layer0_outputs(8242) <= (inputs(38)) xor (inputs(79));
    layer0_outputs(8243) <= '0';
    layer0_outputs(8244) <= not((inputs(135)) and (inputs(106)));
    layer0_outputs(8245) <= '1';
    layer0_outputs(8246) <= (inputs(202)) xor (inputs(135));
    layer0_outputs(8247) <= inputs(234);
    layer0_outputs(8248) <= not(inputs(217));
    layer0_outputs(8249) <= (inputs(242)) and (inputs(146));
    layer0_outputs(8250) <= not((inputs(155)) xor (inputs(165)));
    layer0_outputs(8251) <= inputs(18);
    layer0_outputs(8252) <= not(inputs(165));
    layer0_outputs(8253) <= '0';
    layer0_outputs(8254) <= (inputs(71)) and not (inputs(160));
    layer0_outputs(8255) <= (inputs(36)) xor (inputs(105));
    layer0_outputs(8256) <= inputs(9);
    layer0_outputs(8257) <= (inputs(47)) and not (inputs(95));
    layer0_outputs(8258) <= not((inputs(214)) or (inputs(176)));
    layer0_outputs(8259) <= not(inputs(99));
    layer0_outputs(8260) <= (inputs(135)) and not (inputs(198));
    layer0_outputs(8261) <= (inputs(155)) and not (inputs(236));
    layer0_outputs(8262) <= not(inputs(4));
    layer0_outputs(8263) <= not(inputs(11)) or (inputs(16));
    layer0_outputs(8264) <= not(inputs(141));
    layer0_outputs(8265) <= not((inputs(80)) xor (inputs(141)));
    layer0_outputs(8266) <= (inputs(10)) or (inputs(207));
    layer0_outputs(8267) <= not(inputs(213)) or (inputs(64));
    layer0_outputs(8268) <= (inputs(226)) xor (inputs(178));
    layer0_outputs(8269) <= not((inputs(224)) or (inputs(27)));
    layer0_outputs(8270) <= not((inputs(212)) or (inputs(160)));
    layer0_outputs(8271) <= not((inputs(228)) xor (inputs(66)));
    layer0_outputs(8272) <= not((inputs(65)) xor (inputs(78)));
    layer0_outputs(8273) <= not((inputs(166)) xor (inputs(246)));
    layer0_outputs(8274) <= (inputs(183)) and not (inputs(86));
    layer0_outputs(8275) <= (inputs(9)) or (inputs(163));
    layer0_outputs(8276) <= (inputs(230)) and not (inputs(238));
    layer0_outputs(8277) <= (inputs(185)) xor (inputs(11));
    layer0_outputs(8278) <= not(inputs(165)) or (inputs(155));
    layer0_outputs(8279) <= (inputs(189)) xor (inputs(48));
    layer0_outputs(8280) <= (inputs(160)) or (inputs(119));
    layer0_outputs(8281) <= not((inputs(39)) or (inputs(221)));
    layer0_outputs(8282) <= (inputs(67)) and not (inputs(234));
    layer0_outputs(8283) <= not(inputs(235)) or (inputs(65));
    layer0_outputs(8284) <= (inputs(170)) xor (inputs(101));
    layer0_outputs(8285) <= (inputs(237)) and not (inputs(142));
    layer0_outputs(8286) <= not(inputs(156)) or (inputs(164));
    layer0_outputs(8287) <= not((inputs(88)) xor (inputs(90)));
    layer0_outputs(8288) <= not(inputs(254)) or (inputs(22));
    layer0_outputs(8289) <= '1';
    layer0_outputs(8290) <= not((inputs(13)) and (inputs(231)));
    layer0_outputs(8291) <= not(inputs(114));
    layer0_outputs(8292) <= (inputs(208)) and not (inputs(209));
    layer0_outputs(8293) <= inputs(246);
    layer0_outputs(8294) <= not(inputs(90)) or (inputs(68));
    layer0_outputs(8295) <= inputs(117);
    layer0_outputs(8296) <= (inputs(83)) and not (inputs(78));
    layer0_outputs(8297) <= not(inputs(155)) or (inputs(111));
    layer0_outputs(8298) <= not((inputs(165)) or (inputs(18)));
    layer0_outputs(8299) <= '0';
    layer0_outputs(8300) <= not(inputs(212)) or (inputs(63));
    layer0_outputs(8301) <= inputs(20);
    layer0_outputs(8302) <= (inputs(167)) xor (inputs(245));
    layer0_outputs(8303) <= not((inputs(52)) or (inputs(34)));
    layer0_outputs(8304) <= (inputs(181)) or (inputs(196));
    layer0_outputs(8305) <= not(inputs(149));
    layer0_outputs(8306) <= (inputs(18)) xor (inputs(175));
    layer0_outputs(8307) <= not(inputs(222)) or (inputs(161));
    layer0_outputs(8308) <= (inputs(22)) and not (inputs(128));
    layer0_outputs(8309) <= not(inputs(103));
    layer0_outputs(8310) <= not(inputs(184)) or (inputs(140));
    layer0_outputs(8311) <= inputs(26);
    layer0_outputs(8312) <= '0';
    layer0_outputs(8313) <= inputs(190);
    layer0_outputs(8314) <= not((inputs(253)) xor (inputs(133)));
    layer0_outputs(8315) <= not((inputs(49)) or (inputs(232)));
    layer0_outputs(8316) <= (inputs(231)) and not (inputs(254));
    layer0_outputs(8317) <= (inputs(144)) or (inputs(130));
    layer0_outputs(8318) <= not((inputs(204)) or (inputs(244)));
    layer0_outputs(8319) <= not((inputs(103)) xor (inputs(48)));
    layer0_outputs(8320) <= (inputs(117)) and not (inputs(251));
    layer0_outputs(8321) <= (inputs(6)) xor (inputs(106));
    layer0_outputs(8322) <= not((inputs(22)) and (inputs(67)));
    layer0_outputs(8323) <= inputs(215);
    layer0_outputs(8324) <= not(inputs(218)) or (inputs(3));
    layer0_outputs(8325) <= not(inputs(104)) or (inputs(52));
    layer0_outputs(8326) <= inputs(184);
    layer0_outputs(8327) <= not((inputs(134)) xor (inputs(127)));
    layer0_outputs(8328) <= (inputs(164)) or (inputs(77));
    layer0_outputs(8329) <= (inputs(253)) or (inputs(168));
    layer0_outputs(8330) <= (inputs(6)) xor (inputs(164));
    layer0_outputs(8331) <= (inputs(3)) xor (inputs(179));
    layer0_outputs(8332) <= not((inputs(23)) and (inputs(88)));
    layer0_outputs(8333) <= not(inputs(3));
    layer0_outputs(8334) <= not((inputs(193)) and (inputs(185)));
    layer0_outputs(8335) <= not((inputs(69)) or (inputs(221)));
    layer0_outputs(8336) <= not((inputs(249)) or (inputs(237)));
    layer0_outputs(8337) <= not((inputs(186)) and (inputs(195)));
    layer0_outputs(8338) <= not(inputs(135));
    layer0_outputs(8339) <= inputs(40);
    layer0_outputs(8340) <= inputs(113);
    layer0_outputs(8341) <= not(inputs(44));
    layer0_outputs(8342) <= inputs(143);
    layer0_outputs(8343) <= not((inputs(134)) or (inputs(97)));
    layer0_outputs(8344) <= not((inputs(235)) xor (inputs(223)));
    layer0_outputs(8345) <= '0';
    layer0_outputs(8346) <= (inputs(156)) and not (inputs(207));
    layer0_outputs(8347) <= not((inputs(83)) xor (inputs(60)));
    layer0_outputs(8348) <= not((inputs(215)) and (inputs(170)));
    layer0_outputs(8349) <= (inputs(129)) or (inputs(133));
    layer0_outputs(8350) <= (inputs(233)) xor (inputs(79));
    layer0_outputs(8351) <= '0';
    layer0_outputs(8352) <= inputs(129);
    layer0_outputs(8353) <= '1';
    layer0_outputs(8354) <= (inputs(15)) and (inputs(152));
    layer0_outputs(8355) <= inputs(77);
    layer0_outputs(8356) <= (inputs(49)) or (inputs(3));
    layer0_outputs(8357) <= not((inputs(241)) or (inputs(134)));
    layer0_outputs(8358) <= not(inputs(60)) or (inputs(16));
    layer0_outputs(8359) <= inputs(181);
    layer0_outputs(8360) <= not(inputs(135));
    layer0_outputs(8361) <= not(inputs(75));
    layer0_outputs(8362) <= not((inputs(29)) or (inputs(183)));
    layer0_outputs(8363) <= (inputs(240)) and not (inputs(10));
    layer0_outputs(8364) <= inputs(183);
    layer0_outputs(8365) <= (inputs(194)) or (inputs(9));
    layer0_outputs(8366) <= inputs(118);
    layer0_outputs(8367) <= (inputs(93)) or (inputs(121));
    layer0_outputs(8368) <= not(inputs(57)) or (inputs(20));
    layer0_outputs(8369) <= not(inputs(59)) or (inputs(44));
    layer0_outputs(8370) <= (inputs(101)) and not (inputs(23));
    layer0_outputs(8371) <= not(inputs(226));
    layer0_outputs(8372) <= not(inputs(0)) or (inputs(14));
    layer0_outputs(8373) <= (inputs(57)) and not (inputs(64));
    layer0_outputs(8374) <= inputs(206);
    layer0_outputs(8375) <= (inputs(192)) xor (inputs(188));
    layer0_outputs(8376) <= not((inputs(89)) or (inputs(180)));
    layer0_outputs(8377) <= not((inputs(200)) xor (inputs(221)));
    layer0_outputs(8378) <= inputs(156);
    layer0_outputs(8379) <= (inputs(52)) and not (inputs(7));
    layer0_outputs(8380) <= (inputs(216)) and not (inputs(186));
    layer0_outputs(8381) <= not(inputs(248)) or (inputs(246));
    layer0_outputs(8382) <= not(inputs(60)) or (inputs(82));
    layer0_outputs(8383) <= (inputs(100)) and not (inputs(254));
    layer0_outputs(8384) <= not(inputs(85));
    layer0_outputs(8385) <= '1';
    layer0_outputs(8386) <= not(inputs(80)) or (inputs(7));
    layer0_outputs(8387) <= not((inputs(164)) xor (inputs(151)));
    layer0_outputs(8388) <= not((inputs(115)) xor (inputs(50)));
    layer0_outputs(8389) <= not((inputs(165)) or (inputs(116)));
    layer0_outputs(8390) <= not((inputs(83)) or (inputs(197)));
    layer0_outputs(8391) <= (inputs(7)) and (inputs(210));
    layer0_outputs(8392) <= (inputs(193)) and (inputs(28));
    layer0_outputs(8393) <= inputs(55);
    layer0_outputs(8394) <= not((inputs(88)) xor (inputs(76)));
    layer0_outputs(8395) <= (inputs(163)) and not (inputs(228));
    layer0_outputs(8396) <= not(inputs(192));
    layer0_outputs(8397) <= not(inputs(106));
    layer0_outputs(8398) <= not(inputs(58)) or (inputs(218));
    layer0_outputs(8399) <= not((inputs(2)) or (inputs(137)));
    layer0_outputs(8400) <= (inputs(233)) and not (inputs(51));
    layer0_outputs(8401) <= (inputs(63)) and not (inputs(206));
    layer0_outputs(8402) <= not((inputs(92)) xor (inputs(202)));
    layer0_outputs(8403) <= (inputs(106)) and not (inputs(211));
    layer0_outputs(8404) <= not((inputs(142)) or (inputs(40)));
    layer0_outputs(8405) <= (inputs(140)) and not (inputs(99));
    layer0_outputs(8406) <= inputs(229);
    layer0_outputs(8407) <= (inputs(111)) xor (inputs(184));
    layer0_outputs(8408) <= not(inputs(179));
    layer0_outputs(8409) <= not((inputs(76)) xor (inputs(208)));
    layer0_outputs(8410) <= not(inputs(196));
    layer0_outputs(8411) <= not(inputs(151));
    layer0_outputs(8412) <= (inputs(218)) and not (inputs(206));
    layer0_outputs(8413) <= inputs(88);
    layer0_outputs(8414) <= inputs(162);
    layer0_outputs(8415) <= not((inputs(194)) and (inputs(70)));
    layer0_outputs(8416) <= (inputs(236)) xor (inputs(209));
    layer0_outputs(8417) <= inputs(110);
    layer0_outputs(8418) <= (inputs(233)) xor (inputs(160));
    layer0_outputs(8419) <= inputs(72);
    layer0_outputs(8420) <= inputs(166);
    layer0_outputs(8421) <= not((inputs(84)) xor (inputs(164)));
    layer0_outputs(8422) <= not((inputs(71)) or (inputs(21)));
    layer0_outputs(8423) <= not(inputs(109));
    layer0_outputs(8424) <= (inputs(84)) xor (inputs(41));
    layer0_outputs(8425) <= not((inputs(232)) or (inputs(87)));
    layer0_outputs(8426) <= (inputs(22)) and not (inputs(227));
    layer0_outputs(8427) <= not((inputs(111)) xor (inputs(65)));
    layer0_outputs(8428) <= not(inputs(87));
    layer0_outputs(8429) <= not(inputs(253)) or (inputs(43));
    layer0_outputs(8430) <= (inputs(70)) xor (inputs(85));
    layer0_outputs(8431) <= not(inputs(127)) or (inputs(223));
    layer0_outputs(8432) <= '1';
    layer0_outputs(8433) <= (inputs(167)) xor (inputs(234));
    layer0_outputs(8434) <= (inputs(212)) and not (inputs(205));
    layer0_outputs(8435) <= (inputs(78)) and (inputs(30));
    layer0_outputs(8436) <= not(inputs(105));
    layer0_outputs(8437) <= (inputs(189)) xor (inputs(68));
    layer0_outputs(8438) <= '1';
    layer0_outputs(8439) <= (inputs(19)) and not (inputs(222));
    layer0_outputs(8440) <= not(inputs(42));
    layer0_outputs(8441) <= not(inputs(190));
    layer0_outputs(8442) <= (inputs(125)) or (inputs(151));
    layer0_outputs(8443) <= not(inputs(188)) or (inputs(253));
    layer0_outputs(8444) <= not((inputs(58)) xor (inputs(50)));
    layer0_outputs(8445) <= not(inputs(117)) or (inputs(3));
    layer0_outputs(8446) <= (inputs(117)) and not (inputs(145));
    layer0_outputs(8447) <= (inputs(77)) xor (inputs(104));
    layer0_outputs(8448) <= not(inputs(60));
    layer0_outputs(8449) <= inputs(57);
    layer0_outputs(8450) <= not((inputs(34)) xor (inputs(93)));
    layer0_outputs(8451) <= (inputs(251)) xor (inputs(162));
    layer0_outputs(8452) <= '0';
    layer0_outputs(8453) <= (inputs(226)) and not (inputs(157));
    layer0_outputs(8454) <= not(inputs(14));
    layer0_outputs(8455) <= not((inputs(64)) or (inputs(215)));
    layer0_outputs(8456) <= (inputs(223)) or (inputs(155));
    layer0_outputs(8457) <= (inputs(137)) xor (inputs(126));
    layer0_outputs(8458) <= (inputs(165)) and not (inputs(211));
    layer0_outputs(8459) <= not(inputs(181)) or (inputs(210));
    layer0_outputs(8460) <= not((inputs(237)) or (inputs(122)));
    layer0_outputs(8461) <= not(inputs(203));
    layer0_outputs(8462) <= '1';
    layer0_outputs(8463) <= not((inputs(128)) xor (inputs(180)));
    layer0_outputs(8464) <= not((inputs(119)) or (inputs(4)));
    layer0_outputs(8465) <= inputs(67);
    layer0_outputs(8466) <= not((inputs(128)) xor (inputs(105)));
    layer0_outputs(8467) <= (inputs(48)) and not (inputs(204));
    layer0_outputs(8468) <= not(inputs(105));
    layer0_outputs(8469) <= '1';
    layer0_outputs(8470) <= not((inputs(80)) or (inputs(77)));
    layer0_outputs(8471) <= not(inputs(143));
    layer0_outputs(8472) <= (inputs(180)) or (inputs(92));
    layer0_outputs(8473) <= not(inputs(173));
    layer0_outputs(8474) <= (inputs(22)) and not (inputs(208));
    layer0_outputs(8475) <= inputs(120);
    layer0_outputs(8476) <= (inputs(24)) or (inputs(37));
    layer0_outputs(8477) <= inputs(38);
    layer0_outputs(8478) <= not((inputs(189)) xor (inputs(235)));
    layer0_outputs(8479) <= (inputs(250)) and (inputs(143));
    layer0_outputs(8480) <= inputs(135);
    layer0_outputs(8481) <= not(inputs(70));
    layer0_outputs(8482) <= inputs(172);
    layer0_outputs(8483) <= not(inputs(136));
    layer0_outputs(8484) <= (inputs(176)) xor (inputs(180));
    layer0_outputs(8485) <= inputs(177);
    layer0_outputs(8486) <= not(inputs(20));
    layer0_outputs(8487) <= not((inputs(196)) or (inputs(232)));
    layer0_outputs(8488) <= (inputs(29)) or (inputs(122));
    layer0_outputs(8489) <= inputs(121);
    layer0_outputs(8490) <= not(inputs(120));
    layer0_outputs(8491) <= (inputs(2)) or (inputs(78));
    layer0_outputs(8492) <= (inputs(86)) and not (inputs(180));
    layer0_outputs(8493) <= inputs(148);
    layer0_outputs(8494) <= not(inputs(140));
    layer0_outputs(8495) <= inputs(11);
    layer0_outputs(8496) <= not(inputs(72)) or (inputs(61));
    layer0_outputs(8497) <= not(inputs(160)) or (inputs(228));
    layer0_outputs(8498) <= not((inputs(82)) or (inputs(239)));
    layer0_outputs(8499) <= (inputs(227)) or (inputs(6));
    layer0_outputs(8500) <= inputs(107);
    layer0_outputs(8501) <= not(inputs(167)) or (inputs(205));
    layer0_outputs(8502) <= not((inputs(77)) or (inputs(111)));
    layer0_outputs(8503) <= (inputs(62)) and not (inputs(174));
    layer0_outputs(8504) <= inputs(43);
    layer0_outputs(8505) <= (inputs(213)) xor (inputs(184));
    layer0_outputs(8506) <= (inputs(202)) and not (inputs(99));
    layer0_outputs(8507) <= not(inputs(246));
    layer0_outputs(8508) <= (inputs(184)) and not (inputs(180));
    layer0_outputs(8509) <= not((inputs(28)) xor (inputs(155)));
    layer0_outputs(8510) <= (inputs(173)) and not (inputs(201));
    layer0_outputs(8511) <= not(inputs(136)) or (inputs(127));
    layer0_outputs(8512) <= (inputs(202)) or (inputs(41));
    layer0_outputs(8513) <= (inputs(130)) or (inputs(209));
    layer0_outputs(8514) <= (inputs(233)) xor (inputs(0));
    layer0_outputs(8515) <= not((inputs(87)) or (inputs(207)));
    layer0_outputs(8516) <= (inputs(45)) and not (inputs(31));
    layer0_outputs(8517) <= (inputs(36)) or (inputs(234));
    layer0_outputs(8518) <= not(inputs(242));
    layer0_outputs(8519) <= (inputs(6)) or (inputs(218));
    layer0_outputs(8520) <= not(inputs(98));
    layer0_outputs(8521) <= inputs(10);
    layer0_outputs(8522) <= not(inputs(110)) or (inputs(227));
    layer0_outputs(8523) <= not((inputs(145)) xor (inputs(39)));
    layer0_outputs(8524) <= (inputs(41)) xor (inputs(103));
    layer0_outputs(8525) <= not(inputs(42));
    layer0_outputs(8526) <= inputs(48);
    layer0_outputs(8527) <= (inputs(70)) or (inputs(188));
    layer0_outputs(8528) <= (inputs(56)) or (inputs(171));
    layer0_outputs(8529) <= not((inputs(201)) xor (inputs(86)));
    layer0_outputs(8530) <= (inputs(185)) or (inputs(80));
    layer0_outputs(8531) <= '0';
    layer0_outputs(8532) <= (inputs(70)) xor (inputs(100));
    layer0_outputs(8533) <= inputs(101);
    layer0_outputs(8534) <= not((inputs(148)) xor (inputs(163)));
    layer0_outputs(8535) <= (inputs(183)) and not (inputs(145));
    layer0_outputs(8536) <= not((inputs(40)) or (inputs(211)));
    layer0_outputs(8537) <= inputs(71);
    layer0_outputs(8538) <= not((inputs(143)) or (inputs(176)));
    layer0_outputs(8539) <= not(inputs(23));
    layer0_outputs(8540) <= (inputs(61)) xor (inputs(198));
    layer0_outputs(8541) <= not(inputs(84));
    layer0_outputs(8542) <= not(inputs(120)) or (inputs(204));
    layer0_outputs(8543) <= not((inputs(175)) or (inputs(138)));
    layer0_outputs(8544) <= inputs(109);
    layer0_outputs(8545) <= inputs(152);
    layer0_outputs(8546) <= inputs(229);
    layer0_outputs(8547) <= (inputs(227)) and not (inputs(6));
    layer0_outputs(8548) <= not((inputs(233)) or (inputs(187)));
    layer0_outputs(8549) <= inputs(74);
    layer0_outputs(8550) <= not((inputs(118)) xor (inputs(29)));
    layer0_outputs(8551) <= inputs(53);
    layer0_outputs(8552) <= not(inputs(166));
    layer0_outputs(8553) <= not((inputs(100)) or (inputs(131)));
    layer0_outputs(8554) <= not((inputs(41)) or (inputs(200)));
    layer0_outputs(8555) <= (inputs(254)) and (inputs(208));
    layer0_outputs(8556) <= not(inputs(8));
    layer0_outputs(8557) <= (inputs(123)) or (inputs(234));
    layer0_outputs(8558) <= (inputs(142)) xor (inputs(154));
    layer0_outputs(8559) <= not((inputs(174)) or (inputs(158)));
    layer0_outputs(8560) <= inputs(32);
    layer0_outputs(8561) <= not((inputs(141)) and (inputs(242)));
    layer0_outputs(8562) <= not((inputs(128)) and (inputs(10)));
    layer0_outputs(8563) <= (inputs(54)) and not (inputs(47));
    layer0_outputs(8564) <= (inputs(239)) and not (inputs(13));
    layer0_outputs(8565) <= (inputs(171)) or (inputs(121));
    layer0_outputs(8566) <= (inputs(62)) and not (inputs(245));
    layer0_outputs(8567) <= (inputs(65)) xor (inputs(223));
    layer0_outputs(8568) <= not((inputs(163)) xor (inputs(57)));
    layer0_outputs(8569) <= (inputs(242)) and (inputs(81));
    layer0_outputs(8570) <= not(inputs(151));
    layer0_outputs(8571) <= inputs(76);
    layer0_outputs(8572) <= not((inputs(99)) xor (inputs(38)));
    layer0_outputs(8573) <= inputs(58);
    layer0_outputs(8574) <= '0';
    layer0_outputs(8575) <= not((inputs(72)) xor (inputs(196)));
    layer0_outputs(8576) <= inputs(122);
    layer0_outputs(8577) <= not((inputs(210)) or (inputs(59)));
    layer0_outputs(8578) <= not(inputs(182));
    layer0_outputs(8579) <= '0';
    layer0_outputs(8580) <= (inputs(8)) and not (inputs(164));
    layer0_outputs(8581) <= not(inputs(192));
    layer0_outputs(8582) <= not((inputs(165)) xor (inputs(27)));
    layer0_outputs(8583) <= (inputs(226)) or (inputs(20));
    layer0_outputs(8584) <= inputs(89);
    layer0_outputs(8585) <= inputs(43);
    layer0_outputs(8586) <= not(inputs(163)) or (inputs(30));
    layer0_outputs(8587) <= '0';
    layer0_outputs(8588) <= (inputs(93)) xor (inputs(97));
    layer0_outputs(8589) <= inputs(156);
    layer0_outputs(8590) <= (inputs(200)) or (inputs(10));
    layer0_outputs(8591) <= not(inputs(171)) or (inputs(93));
    layer0_outputs(8592) <= not((inputs(84)) or (inputs(250)));
    layer0_outputs(8593) <= not(inputs(0));
    layer0_outputs(8594) <= not((inputs(57)) or (inputs(77)));
    layer0_outputs(8595) <= not((inputs(255)) xor (inputs(59)));
    layer0_outputs(8596) <= inputs(151);
    layer0_outputs(8597) <= inputs(86);
    layer0_outputs(8598) <= not(inputs(29)) or (inputs(48));
    layer0_outputs(8599) <= not((inputs(74)) or (inputs(64)));
    layer0_outputs(8600) <= (inputs(43)) or (inputs(141));
    layer0_outputs(8601) <= not(inputs(68));
    layer0_outputs(8602) <= (inputs(131)) and not (inputs(127));
    layer0_outputs(8603) <= not((inputs(86)) or (inputs(45)));
    layer0_outputs(8604) <= not(inputs(92));
    layer0_outputs(8605) <= (inputs(207)) and not (inputs(124));
    layer0_outputs(8606) <= not(inputs(213));
    layer0_outputs(8607) <= (inputs(121)) or (inputs(177));
    layer0_outputs(8608) <= not(inputs(197)) or (inputs(230));
    layer0_outputs(8609) <= (inputs(124)) or (inputs(15));
    layer0_outputs(8610) <= (inputs(10)) xor (inputs(168));
    layer0_outputs(8611) <= not((inputs(231)) or (inputs(105)));
    layer0_outputs(8612) <= not(inputs(134));
    layer0_outputs(8613) <= (inputs(69)) xor (inputs(46));
    layer0_outputs(8614) <= not((inputs(149)) and (inputs(197)));
    layer0_outputs(8615) <= (inputs(24)) xor (inputs(229));
    layer0_outputs(8616) <= not((inputs(209)) or (inputs(25)));
    layer0_outputs(8617) <= (inputs(231)) xor (inputs(158));
    layer0_outputs(8618) <= not((inputs(107)) or (inputs(97)));
    layer0_outputs(8619) <= not((inputs(92)) xor (inputs(150)));
    layer0_outputs(8620) <= (inputs(220)) and not (inputs(70));
    layer0_outputs(8621) <= not(inputs(102)) or (inputs(239));
    layer0_outputs(8622) <= (inputs(68)) and not (inputs(218));
    layer0_outputs(8623) <= (inputs(91)) or (inputs(163));
    layer0_outputs(8624) <= not(inputs(151)) or (inputs(2));
    layer0_outputs(8625) <= (inputs(118)) and not (inputs(83));
    layer0_outputs(8626) <= not(inputs(164)) or (inputs(205));
    layer0_outputs(8627) <= (inputs(92)) and not (inputs(113));
    layer0_outputs(8628) <= (inputs(3)) or (inputs(164));
    layer0_outputs(8629) <= (inputs(142)) and not (inputs(234));
    layer0_outputs(8630) <= not((inputs(154)) or (inputs(2)));
    layer0_outputs(8631) <= not((inputs(49)) xor (inputs(152)));
    layer0_outputs(8632) <= not((inputs(242)) xor (inputs(220)));
    layer0_outputs(8633) <= (inputs(101)) and not (inputs(239));
    layer0_outputs(8634) <= inputs(64);
    layer0_outputs(8635) <= (inputs(247)) or (inputs(85));
    layer0_outputs(8636) <= not((inputs(2)) and (inputs(1)));
    layer0_outputs(8637) <= not(inputs(196));
    layer0_outputs(8638) <= (inputs(211)) and not (inputs(236));
    layer0_outputs(8639) <= '1';
    layer0_outputs(8640) <= not((inputs(128)) and (inputs(247)));
    layer0_outputs(8641) <= not(inputs(121)) or (inputs(92));
    layer0_outputs(8642) <= (inputs(216)) or (inputs(245));
    layer0_outputs(8643) <= not((inputs(174)) xor (inputs(118)));
    layer0_outputs(8644) <= not(inputs(47)) or (inputs(29));
    layer0_outputs(8645) <= not((inputs(195)) xor (inputs(155)));
    layer0_outputs(8646) <= (inputs(87)) and not (inputs(161));
    layer0_outputs(8647) <= (inputs(152)) and not (inputs(145));
    layer0_outputs(8648) <= '1';
    layer0_outputs(8649) <= '1';
    layer0_outputs(8650) <= not((inputs(249)) xor (inputs(120)));
    layer0_outputs(8651) <= inputs(232);
    layer0_outputs(8652) <= (inputs(83)) and not (inputs(146));
    layer0_outputs(8653) <= not((inputs(247)) xor (inputs(197)));
    layer0_outputs(8654) <= not(inputs(93));
    layer0_outputs(8655) <= (inputs(77)) and (inputs(177));
    layer0_outputs(8656) <= not(inputs(205));
    layer0_outputs(8657) <= not(inputs(157));
    layer0_outputs(8658) <= (inputs(39)) and not (inputs(79));
    layer0_outputs(8659) <= not(inputs(14));
    layer0_outputs(8660) <= not((inputs(69)) or (inputs(90)));
    layer0_outputs(8661) <= not(inputs(182));
    layer0_outputs(8662) <= not(inputs(124));
    layer0_outputs(8663) <= (inputs(212)) and not (inputs(50));
    layer0_outputs(8664) <= not(inputs(16));
    layer0_outputs(8665) <= not(inputs(56));
    layer0_outputs(8666) <= not(inputs(192)) or (inputs(175));
    layer0_outputs(8667) <= '1';
    layer0_outputs(8668) <= (inputs(167)) and not (inputs(92));
    layer0_outputs(8669) <= not((inputs(15)) xor (inputs(191)));
    layer0_outputs(8670) <= inputs(2);
    layer0_outputs(8671) <= not((inputs(38)) or (inputs(57)));
    layer0_outputs(8672) <= (inputs(17)) xor (inputs(11));
    layer0_outputs(8673) <= (inputs(121)) and not (inputs(208));
    layer0_outputs(8674) <= not(inputs(236));
    layer0_outputs(8675) <= (inputs(162)) xor (inputs(208));
    layer0_outputs(8676) <= inputs(255);
    layer0_outputs(8677) <= '1';
    layer0_outputs(8678) <= (inputs(122)) or (inputs(133));
    layer0_outputs(8679) <= (inputs(196)) or (inputs(202));
    layer0_outputs(8680) <= not(inputs(219)) or (inputs(202));
    layer0_outputs(8681) <= not((inputs(13)) and (inputs(2)));
    layer0_outputs(8682) <= not((inputs(131)) or (inputs(217)));
    layer0_outputs(8683) <= not((inputs(116)) and (inputs(163)));
    layer0_outputs(8684) <= not((inputs(55)) or (inputs(108)));
    layer0_outputs(8685) <= not(inputs(122)) or (inputs(88));
    layer0_outputs(8686) <= (inputs(188)) xor (inputs(37));
    layer0_outputs(8687) <= (inputs(220)) or (inputs(63));
    layer0_outputs(8688) <= (inputs(107)) and not (inputs(47));
    layer0_outputs(8689) <= (inputs(83)) and (inputs(81));
    layer0_outputs(8690) <= '0';
    layer0_outputs(8691) <= not(inputs(72));
    layer0_outputs(8692) <= not((inputs(241)) xor (inputs(39)));
    layer0_outputs(8693) <= (inputs(234)) or (inputs(91));
    layer0_outputs(8694) <= (inputs(20)) or (inputs(49));
    layer0_outputs(8695) <= inputs(133);
    layer0_outputs(8696) <= not((inputs(77)) and (inputs(244)));
    layer0_outputs(8697) <= (inputs(87)) and not (inputs(25));
    layer0_outputs(8698) <= not(inputs(21)) or (inputs(160));
    layer0_outputs(8699) <= not((inputs(216)) xor (inputs(3)));
    layer0_outputs(8700) <= not((inputs(57)) xor (inputs(234)));
    layer0_outputs(8701) <= not(inputs(162)) or (inputs(48));
    layer0_outputs(8702) <= not(inputs(73));
    layer0_outputs(8703) <= inputs(186);
    layer0_outputs(8704) <= not(inputs(150));
    layer0_outputs(8705) <= (inputs(50)) xor (inputs(170));
    layer0_outputs(8706) <= (inputs(56)) or (inputs(217));
    layer0_outputs(8707) <= not((inputs(200)) xor (inputs(35)));
    layer0_outputs(8708) <= not((inputs(145)) xor (inputs(30)));
    layer0_outputs(8709) <= (inputs(98)) xor (inputs(197));
    layer0_outputs(8710) <= (inputs(143)) or (inputs(164));
    layer0_outputs(8711) <= (inputs(154)) and not (inputs(38));
    layer0_outputs(8712) <= '1';
    layer0_outputs(8713) <= (inputs(31)) xor (inputs(18));
    layer0_outputs(8714) <= not((inputs(228)) xor (inputs(97)));
    layer0_outputs(8715) <= inputs(52);
    layer0_outputs(8716) <= not((inputs(20)) xor (inputs(107)));
    layer0_outputs(8717) <= not(inputs(77));
    layer0_outputs(8718) <= (inputs(196)) xor (inputs(227));
    layer0_outputs(8719) <= (inputs(9)) and not (inputs(3));
    layer0_outputs(8720) <= not(inputs(134)) or (inputs(211));
    layer0_outputs(8721) <= (inputs(210)) xor (inputs(145));
    layer0_outputs(8722) <= not(inputs(4));
    layer0_outputs(8723) <= not((inputs(141)) or (inputs(213)));
    layer0_outputs(8724) <= not((inputs(213)) or (inputs(81)));
    layer0_outputs(8725) <= (inputs(175)) or (inputs(37));
    layer0_outputs(8726) <= inputs(197);
    layer0_outputs(8727) <= not(inputs(87));
    layer0_outputs(8728) <= (inputs(62)) and (inputs(235));
    layer0_outputs(8729) <= '1';
    layer0_outputs(8730) <= (inputs(164)) and not (inputs(115));
    layer0_outputs(8731) <= (inputs(209)) xor (inputs(75));
    layer0_outputs(8732) <= (inputs(173)) and not (inputs(75));
    layer0_outputs(8733) <= (inputs(27)) and not (inputs(219));
    layer0_outputs(8734) <= not(inputs(182));
    layer0_outputs(8735) <= inputs(156);
    layer0_outputs(8736) <= '0';
    layer0_outputs(8737) <= (inputs(155)) and not (inputs(63));
    layer0_outputs(8738) <= '0';
    layer0_outputs(8739) <= not((inputs(134)) or (inputs(111)));
    layer0_outputs(8740) <= not(inputs(202));
    layer0_outputs(8741) <= (inputs(218)) or (inputs(227));
    layer0_outputs(8742) <= (inputs(181)) xor (inputs(193));
    layer0_outputs(8743) <= (inputs(134)) and not (inputs(67));
    layer0_outputs(8744) <= '0';
    layer0_outputs(8745) <= not(inputs(23));
    layer0_outputs(8746) <= not(inputs(165)) or (inputs(76));
    layer0_outputs(8747) <= (inputs(170)) or (inputs(54));
    layer0_outputs(8748) <= (inputs(231)) xor (inputs(89));
    layer0_outputs(8749) <= not((inputs(215)) or (inputs(4)));
    layer0_outputs(8750) <= not((inputs(77)) or (inputs(119)));
    layer0_outputs(8751) <= inputs(154);
    layer0_outputs(8752) <= inputs(98);
    layer0_outputs(8753) <= (inputs(164)) and not (inputs(194));
    layer0_outputs(8754) <= (inputs(53)) xor (inputs(172));
    layer0_outputs(8755) <= not((inputs(19)) and (inputs(57)));
    layer0_outputs(8756) <= inputs(162);
    layer0_outputs(8757) <= not(inputs(206)) or (inputs(178));
    layer0_outputs(8758) <= not(inputs(150));
    layer0_outputs(8759) <= (inputs(198)) or (inputs(140));
    layer0_outputs(8760) <= not(inputs(138));
    layer0_outputs(8761) <= inputs(200);
    layer0_outputs(8762) <= (inputs(216)) and not (inputs(210));
    layer0_outputs(8763) <= inputs(0);
    layer0_outputs(8764) <= not(inputs(76));
    layer0_outputs(8765) <= '1';
    layer0_outputs(8766) <= not((inputs(115)) or (inputs(120)));
    layer0_outputs(8767) <= inputs(74);
    layer0_outputs(8768) <= not(inputs(216));
    layer0_outputs(8769) <= not((inputs(9)) and (inputs(234)));
    layer0_outputs(8770) <= not(inputs(56));
    layer0_outputs(8771) <= '0';
    layer0_outputs(8772) <= (inputs(242)) and not (inputs(243));
    layer0_outputs(8773) <= inputs(148);
    layer0_outputs(8774) <= not((inputs(132)) xor (inputs(154)));
    layer0_outputs(8775) <= inputs(164);
    layer0_outputs(8776) <= not(inputs(165)) or (inputs(25));
    layer0_outputs(8777) <= (inputs(186)) or (inputs(231));
    layer0_outputs(8778) <= inputs(204);
    layer0_outputs(8779) <= not((inputs(203)) xor (inputs(93)));
    layer0_outputs(8780) <= (inputs(109)) or (inputs(108));
    layer0_outputs(8781) <= (inputs(123)) xor (inputs(90));
    layer0_outputs(8782) <= inputs(252);
    layer0_outputs(8783) <= (inputs(58)) and (inputs(9));
    layer0_outputs(8784) <= (inputs(165)) xor (inputs(108));
    layer0_outputs(8785) <= (inputs(56)) or (inputs(110));
    layer0_outputs(8786) <= not(inputs(218)) or (inputs(231));
    layer0_outputs(8787) <= not((inputs(68)) xor (inputs(132)));
    layer0_outputs(8788) <= (inputs(197)) xor (inputs(130));
    layer0_outputs(8789) <= not(inputs(110)) or (inputs(54));
    layer0_outputs(8790) <= not((inputs(38)) or (inputs(201)));
    layer0_outputs(8791) <= (inputs(103)) or (inputs(145));
    layer0_outputs(8792) <= not(inputs(6)) or (inputs(5));
    layer0_outputs(8793) <= not((inputs(104)) xor (inputs(63)));
    layer0_outputs(8794) <= (inputs(117)) xor (inputs(5));
    layer0_outputs(8795) <= not((inputs(191)) or (inputs(153)));
    layer0_outputs(8796) <= not(inputs(135)) or (inputs(184));
    layer0_outputs(8797) <= not((inputs(225)) or (inputs(207)));
    layer0_outputs(8798) <= (inputs(135)) and not (inputs(66));
    layer0_outputs(8799) <= (inputs(243)) and not (inputs(13));
    layer0_outputs(8800) <= (inputs(145)) xor (inputs(156));
    layer0_outputs(8801) <= not((inputs(185)) xor (inputs(96)));
    layer0_outputs(8802) <= (inputs(177)) and not (inputs(157));
    layer0_outputs(8803) <= not((inputs(201)) or (inputs(223)));
    layer0_outputs(8804) <= not(inputs(108)) or (inputs(134));
    layer0_outputs(8805) <= (inputs(94)) or (inputs(119));
    layer0_outputs(8806) <= '1';
    layer0_outputs(8807) <= (inputs(197)) and not (inputs(241));
    layer0_outputs(8808) <= (inputs(157)) and not (inputs(91));
    layer0_outputs(8809) <= '1';
    layer0_outputs(8810) <= (inputs(174)) and (inputs(48));
    layer0_outputs(8811) <= not(inputs(129)) or (inputs(22));
    layer0_outputs(8812) <= (inputs(230)) xor (inputs(217));
    layer0_outputs(8813) <= inputs(162);
    layer0_outputs(8814) <= (inputs(147)) or (inputs(69));
    layer0_outputs(8815) <= inputs(115);
    layer0_outputs(8816) <= not((inputs(54)) or (inputs(92)));
    layer0_outputs(8817) <= '0';
    layer0_outputs(8818) <= (inputs(45)) and not (inputs(60));
    layer0_outputs(8819) <= not(inputs(75)) or (inputs(214));
    layer0_outputs(8820) <= not((inputs(223)) and (inputs(126)));
    layer0_outputs(8821) <= (inputs(88)) and not (inputs(21));
    layer0_outputs(8822) <= (inputs(168)) and not (inputs(16));
    layer0_outputs(8823) <= not((inputs(94)) or (inputs(15)));
    layer0_outputs(8824) <= not(inputs(220));
    layer0_outputs(8825) <= not(inputs(181));
    layer0_outputs(8826) <= not((inputs(0)) xor (inputs(184)));
    layer0_outputs(8827) <= not((inputs(225)) and (inputs(46)));
    layer0_outputs(8828) <= (inputs(69)) and not (inputs(127));
    layer0_outputs(8829) <= (inputs(203)) xor (inputs(54));
    layer0_outputs(8830) <= (inputs(178)) and not (inputs(222));
    layer0_outputs(8831) <= not(inputs(137)) or (inputs(213));
    layer0_outputs(8832) <= not(inputs(11));
    layer0_outputs(8833) <= not((inputs(0)) xor (inputs(34)));
    layer0_outputs(8834) <= not((inputs(47)) xor (inputs(177)));
    layer0_outputs(8835) <= inputs(8);
    layer0_outputs(8836) <= (inputs(214)) or (inputs(210));
    layer0_outputs(8837) <= (inputs(213)) or (inputs(89));
    layer0_outputs(8838) <= not(inputs(217)) or (inputs(238));
    layer0_outputs(8839) <= not((inputs(250)) or (inputs(187)));
    layer0_outputs(8840) <= not(inputs(200)) or (inputs(95));
    layer0_outputs(8841) <= not((inputs(29)) or (inputs(196)));
    layer0_outputs(8842) <= not(inputs(147)) or (inputs(63));
    layer0_outputs(8843) <= not((inputs(155)) and (inputs(170)));
    layer0_outputs(8844) <= (inputs(166)) xor (inputs(33));
    layer0_outputs(8845) <= (inputs(108)) and not (inputs(177));
    layer0_outputs(8846) <= (inputs(104)) xor (inputs(81));
    layer0_outputs(8847) <= (inputs(151)) and not (inputs(226));
    layer0_outputs(8848) <= not(inputs(1)) or (inputs(145));
    layer0_outputs(8849) <= not((inputs(168)) or (inputs(250)));
    layer0_outputs(8850) <= (inputs(150)) and not (inputs(123));
    layer0_outputs(8851) <= (inputs(4)) or (inputs(57));
    layer0_outputs(8852) <= (inputs(197)) and not (inputs(178));
    layer0_outputs(8853) <= not(inputs(23));
    layer0_outputs(8854) <= not(inputs(181));
    layer0_outputs(8855) <= not(inputs(154));
    layer0_outputs(8856) <= not(inputs(113));
    layer0_outputs(8857) <= (inputs(146)) and not (inputs(161));
    layer0_outputs(8858) <= (inputs(230)) and not (inputs(0));
    layer0_outputs(8859) <= not(inputs(69)) or (inputs(7));
    layer0_outputs(8860) <= inputs(53);
    layer0_outputs(8861) <= (inputs(48)) xor (inputs(51));
    layer0_outputs(8862) <= inputs(169);
    layer0_outputs(8863) <= (inputs(216)) or (inputs(82));
    layer0_outputs(8864) <= not((inputs(103)) or (inputs(163)));
    layer0_outputs(8865) <= inputs(153);
    layer0_outputs(8866) <= inputs(13);
    layer0_outputs(8867) <= (inputs(67)) and not (inputs(70));
    layer0_outputs(8868) <= not(inputs(184));
    layer0_outputs(8869) <= (inputs(42)) xor (inputs(180));
    layer0_outputs(8870) <= '0';
    layer0_outputs(8871) <= not((inputs(254)) and (inputs(46)));
    layer0_outputs(8872) <= not(inputs(214)) or (inputs(120));
    layer0_outputs(8873) <= (inputs(99)) or (inputs(78));
    layer0_outputs(8874) <= not((inputs(157)) or (inputs(163)));
    layer0_outputs(8875) <= not(inputs(41)) or (inputs(3));
    layer0_outputs(8876) <= (inputs(74)) and not (inputs(245));
    layer0_outputs(8877) <= not((inputs(80)) xor (inputs(87)));
    layer0_outputs(8878) <= (inputs(35)) or (inputs(187));
    layer0_outputs(8879) <= (inputs(174)) and not (inputs(32));
    layer0_outputs(8880) <= inputs(44);
    layer0_outputs(8881) <= (inputs(123)) and not (inputs(160));
    layer0_outputs(8882) <= inputs(138);
    layer0_outputs(8883) <= inputs(181);
    layer0_outputs(8884) <= not(inputs(45));
    layer0_outputs(8885) <= (inputs(147)) xor (inputs(210));
    layer0_outputs(8886) <= not(inputs(1)) or (inputs(237));
    layer0_outputs(8887) <= (inputs(76)) xor (inputs(89));
    layer0_outputs(8888) <= (inputs(104)) xor (inputs(18));
    layer0_outputs(8889) <= not((inputs(12)) or (inputs(21)));
    layer0_outputs(8890) <= not((inputs(121)) xor (inputs(33)));
    layer0_outputs(8891) <= (inputs(98)) or (inputs(43));
    layer0_outputs(8892) <= (inputs(182)) and not (inputs(34));
    layer0_outputs(8893) <= not(inputs(117));
    layer0_outputs(8894) <= (inputs(133)) and not (inputs(105));
    layer0_outputs(8895) <= (inputs(200)) and not (inputs(223));
    layer0_outputs(8896) <= inputs(161);
    layer0_outputs(8897) <= (inputs(153)) and not (inputs(117));
    layer0_outputs(8898) <= (inputs(30)) and not (inputs(192));
    layer0_outputs(8899) <= not((inputs(254)) xor (inputs(86)));
    layer0_outputs(8900) <= (inputs(24)) xor (inputs(248));
    layer0_outputs(8901) <= not(inputs(101));
    layer0_outputs(8902) <= '0';
    layer0_outputs(8903) <= not((inputs(76)) xor (inputs(182)));
    layer0_outputs(8904) <= (inputs(189)) xor (inputs(237));
    layer0_outputs(8905) <= not(inputs(193));
    layer0_outputs(8906) <= not((inputs(82)) xor (inputs(81)));
    layer0_outputs(8907) <= not((inputs(0)) xor (inputs(9)));
    layer0_outputs(8908) <= inputs(183);
    layer0_outputs(8909) <= not(inputs(130));
    layer0_outputs(8910) <= (inputs(180)) or (inputs(163));
    layer0_outputs(8911) <= inputs(3);
    layer0_outputs(8912) <= '0';
    layer0_outputs(8913) <= not((inputs(63)) xor (inputs(50)));
    layer0_outputs(8914) <= not((inputs(82)) or (inputs(221)));
    layer0_outputs(8915) <= not((inputs(99)) and (inputs(64)));
    layer0_outputs(8916) <= (inputs(255)) xor (inputs(66));
    layer0_outputs(8917) <= inputs(85);
    layer0_outputs(8918) <= (inputs(42)) and (inputs(65));
    layer0_outputs(8919) <= (inputs(201)) and not (inputs(8));
    layer0_outputs(8920) <= not((inputs(183)) or (inputs(244)));
    layer0_outputs(8921) <= (inputs(227)) or (inputs(84));
    layer0_outputs(8922) <= (inputs(76)) or (inputs(211));
    layer0_outputs(8923) <= (inputs(255)) and (inputs(97));
    layer0_outputs(8924) <= (inputs(104)) xor (inputs(100));
    layer0_outputs(8925) <= inputs(253);
    layer0_outputs(8926) <= not((inputs(55)) and (inputs(168)));
    layer0_outputs(8927) <= (inputs(204)) and not (inputs(129));
    layer0_outputs(8928) <= inputs(139);
    layer0_outputs(8929) <= not(inputs(138)) or (inputs(181));
    layer0_outputs(8930) <= not((inputs(162)) xor (inputs(60)));
    layer0_outputs(8931) <= (inputs(172)) and not (inputs(81));
    layer0_outputs(8932) <= (inputs(242)) or (inputs(53));
    layer0_outputs(8933) <= not((inputs(62)) xor (inputs(238)));
    layer0_outputs(8934) <= not(inputs(66));
    layer0_outputs(8935) <= (inputs(44)) and not (inputs(144));
    layer0_outputs(8936) <= not(inputs(121));
    layer0_outputs(8937) <= not(inputs(115));
    layer0_outputs(8938) <= not(inputs(71));
    layer0_outputs(8939) <= not(inputs(122)) or (inputs(226));
    layer0_outputs(8940) <= inputs(19);
    layer0_outputs(8941) <= (inputs(187)) xor (inputs(158));
    layer0_outputs(8942) <= inputs(135);
    layer0_outputs(8943) <= not(inputs(131)) or (inputs(192));
    layer0_outputs(8944) <= (inputs(7)) xor (inputs(179));
    layer0_outputs(8945) <= not((inputs(141)) or (inputs(12)));
    layer0_outputs(8946) <= not((inputs(198)) or (inputs(13)));
    layer0_outputs(8947) <= (inputs(153)) or (inputs(130));
    layer0_outputs(8948) <= inputs(206);
    layer0_outputs(8949) <= inputs(157);
    layer0_outputs(8950) <= inputs(173);
    layer0_outputs(8951) <= (inputs(156)) and not (inputs(244));
    layer0_outputs(8952) <= '0';
    layer0_outputs(8953) <= (inputs(226)) xor (inputs(61));
    layer0_outputs(8954) <= not(inputs(149));
    layer0_outputs(8955) <= not((inputs(225)) xor (inputs(83)));
    layer0_outputs(8956) <= inputs(146);
    layer0_outputs(8957) <= not(inputs(209));
    layer0_outputs(8958) <= not((inputs(91)) xor (inputs(157)));
    layer0_outputs(8959) <= not((inputs(108)) or (inputs(23)));
    layer0_outputs(8960) <= (inputs(158)) and (inputs(219));
    layer0_outputs(8961) <= not(inputs(153));
    layer0_outputs(8962) <= (inputs(254)) and not (inputs(64));
    layer0_outputs(8963) <= not(inputs(147)) or (inputs(5));
    layer0_outputs(8964) <= not((inputs(193)) xor (inputs(168)));
    layer0_outputs(8965) <= '1';
    layer0_outputs(8966) <= (inputs(128)) or (inputs(3));
    layer0_outputs(8967) <= '0';
    layer0_outputs(8968) <= not(inputs(5)) or (inputs(84));
    layer0_outputs(8969) <= (inputs(221)) and not (inputs(20));
    layer0_outputs(8970) <= not(inputs(225)) or (inputs(171));
    layer0_outputs(8971) <= (inputs(70)) xor (inputs(107));
    layer0_outputs(8972) <= '1';
    layer0_outputs(8973) <= not(inputs(109)) or (inputs(251));
    layer0_outputs(8974) <= inputs(233);
    layer0_outputs(8975) <= (inputs(10)) or (inputs(28));
    layer0_outputs(8976) <= not((inputs(212)) or (inputs(170)));
    layer0_outputs(8977) <= not(inputs(136));
    layer0_outputs(8978) <= not((inputs(224)) or (inputs(205)));
    layer0_outputs(8979) <= not((inputs(157)) and (inputs(4)));
    layer0_outputs(8980) <= inputs(203);
    layer0_outputs(8981) <= (inputs(43)) and not (inputs(53));
    layer0_outputs(8982) <= not(inputs(37));
    layer0_outputs(8983) <= not(inputs(100)) or (inputs(191));
    layer0_outputs(8984) <= not(inputs(64)) or (inputs(2));
    layer0_outputs(8985) <= (inputs(73)) and not (inputs(231));
    layer0_outputs(8986) <= (inputs(19)) xor (inputs(185));
    layer0_outputs(8987) <= (inputs(23)) and (inputs(23));
    layer0_outputs(8988) <= (inputs(253)) and not (inputs(5));
    layer0_outputs(8989) <= not((inputs(229)) xor (inputs(97)));
    layer0_outputs(8990) <= (inputs(39)) and not (inputs(220));
    layer0_outputs(8991) <= not(inputs(120)) or (inputs(95));
    layer0_outputs(8992) <= (inputs(21)) or (inputs(251));
    layer0_outputs(8993) <= (inputs(85)) and not (inputs(23));
    layer0_outputs(8994) <= (inputs(175)) or (inputs(21));
    layer0_outputs(8995) <= (inputs(140)) or (inputs(157));
    layer0_outputs(8996) <= (inputs(53)) and not (inputs(47));
    layer0_outputs(8997) <= not(inputs(117)) or (inputs(51));
    layer0_outputs(8998) <= inputs(171);
    layer0_outputs(8999) <= (inputs(164)) and not (inputs(19));
    layer0_outputs(9000) <= (inputs(198)) or (inputs(163));
    layer0_outputs(9001) <= (inputs(133)) xor (inputs(191));
    layer0_outputs(9002) <= not((inputs(89)) xor (inputs(142)));
    layer0_outputs(9003) <= (inputs(99)) or (inputs(249));
    layer0_outputs(9004) <= inputs(11);
    layer0_outputs(9005) <= not((inputs(240)) xor (inputs(144)));
    layer0_outputs(9006) <= inputs(84);
    layer0_outputs(9007) <= not((inputs(253)) and (inputs(14)));
    layer0_outputs(9008) <= not(inputs(103)) or (inputs(231));
    layer0_outputs(9009) <= (inputs(51)) and not (inputs(237));
    layer0_outputs(9010) <= not(inputs(22));
    layer0_outputs(9011) <= '1';
    layer0_outputs(9012) <= (inputs(189)) xor (inputs(31));
    layer0_outputs(9013) <= (inputs(87)) and not (inputs(76));
    layer0_outputs(9014) <= not((inputs(53)) and (inputs(201)));
    layer0_outputs(9015) <= not(inputs(147));
    layer0_outputs(9016) <= not((inputs(234)) or (inputs(85)));
    layer0_outputs(9017) <= inputs(181);
    layer0_outputs(9018) <= not((inputs(133)) xor (inputs(196)));
    layer0_outputs(9019) <= not(inputs(152));
    layer0_outputs(9020) <= inputs(167);
    layer0_outputs(9021) <= (inputs(25)) or (inputs(117));
    layer0_outputs(9022) <= not((inputs(38)) or (inputs(146)));
    layer0_outputs(9023) <= not(inputs(48)) or (inputs(8));
    layer0_outputs(9024) <= (inputs(132)) and not (inputs(142));
    layer0_outputs(9025) <= (inputs(145)) and not (inputs(13));
    layer0_outputs(9026) <= not(inputs(202)) or (inputs(101));
    layer0_outputs(9027) <= (inputs(78)) and (inputs(14));
    layer0_outputs(9028) <= not((inputs(141)) or (inputs(141)));
    layer0_outputs(9029) <= (inputs(208)) and not (inputs(142));
    layer0_outputs(9030) <= (inputs(206)) xor (inputs(121));
    layer0_outputs(9031) <= (inputs(0)) xor (inputs(73));
    layer0_outputs(9032) <= not(inputs(40));
    layer0_outputs(9033) <= inputs(212);
    layer0_outputs(9034) <= inputs(187);
    layer0_outputs(9035) <= (inputs(148)) xor (inputs(78));
    layer0_outputs(9036) <= (inputs(40)) or (inputs(164));
    layer0_outputs(9037) <= not((inputs(135)) or (inputs(26)));
    layer0_outputs(9038) <= not(inputs(122));
    layer0_outputs(9039) <= not((inputs(109)) or (inputs(229)));
    layer0_outputs(9040) <= (inputs(41)) or (inputs(156));
    layer0_outputs(9041) <= inputs(44);
    layer0_outputs(9042) <= (inputs(50)) xor (inputs(220));
    layer0_outputs(9043) <= not((inputs(116)) or (inputs(252)));
    layer0_outputs(9044) <= not((inputs(148)) or (inputs(157)));
    layer0_outputs(9045) <= (inputs(25)) or (inputs(188));
    layer0_outputs(9046) <= '1';
    layer0_outputs(9047) <= not(inputs(37));
    layer0_outputs(9048) <= (inputs(219)) and not (inputs(247));
    layer0_outputs(9049) <= (inputs(204)) and not (inputs(22));
    layer0_outputs(9050) <= '0';
    layer0_outputs(9051) <= (inputs(6)) xor (inputs(132));
    layer0_outputs(9052) <= not(inputs(34)) or (inputs(205));
    layer0_outputs(9053) <= (inputs(209)) xor (inputs(230));
    layer0_outputs(9054) <= not((inputs(167)) xor (inputs(17)));
    layer0_outputs(9055) <= (inputs(83)) and (inputs(81));
    layer0_outputs(9056) <= (inputs(57)) xor (inputs(60));
    layer0_outputs(9057) <= (inputs(165)) and not (inputs(24));
    layer0_outputs(9058) <= (inputs(122)) and not (inputs(243));
    layer0_outputs(9059) <= not(inputs(90)) or (inputs(176));
    layer0_outputs(9060) <= (inputs(128)) xor (inputs(216));
    layer0_outputs(9061) <= inputs(86);
    layer0_outputs(9062) <= '1';
    layer0_outputs(9063) <= (inputs(196)) and not (inputs(4));
    layer0_outputs(9064) <= not((inputs(60)) xor (inputs(77)));
    layer0_outputs(9065) <= (inputs(184)) and (inputs(113));
    layer0_outputs(9066) <= '1';
    layer0_outputs(9067) <= not(inputs(194));
    layer0_outputs(9068) <= (inputs(231)) xor (inputs(14));
    layer0_outputs(9069) <= not((inputs(242)) or (inputs(71)));
    layer0_outputs(9070) <= inputs(171);
    layer0_outputs(9071) <= (inputs(137)) xor (inputs(51));
    layer0_outputs(9072) <= inputs(119);
    layer0_outputs(9073) <= not(inputs(220)) or (inputs(36));
    layer0_outputs(9074) <= not(inputs(231));
    layer0_outputs(9075) <= (inputs(3)) and not (inputs(155));
    layer0_outputs(9076) <= inputs(215);
    layer0_outputs(9077) <= not(inputs(195)) or (inputs(160));
    layer0_outputs(9078) <= (inputs(130)) or (inputs(239));
    layer0_outputs(9079) <= not(inputs(85));
    layer0_outputs(9080) <= not((inputs(121)) or (inputs(114)));
    layer0_outputs(9081) <= not(inputs(47));
    layer0_outputs(9082) <= inputs(163);
    layer0_outputs(9083) <= (inputs(125)) or (inputs(236));
    layer0_outputs(9084) <= (inputs(202)) xor (inputs(201));
    layer0_outputs(9085) <= (inputs(52)) and not (inputs(113));
    layer0_outputs(9086) <= (inputs(50)) or (inputs(232));
    layer0_outputs(9087) <= inputs(179);
    layer0_outputs(9088) <= not((inputs(110)) xor (inputs(76)));
    layer0_outputs(9089) <= (inputs(223)) or (inputs(251));
    layer0_outputs(9090) <= inputs(182);
    layer0_outputs(9091) <= inputs(67);
    layer0_outputs(9092) <= not(inputs(117));
    layer0_outputs(9093) <= not((inputs(166)) or (inputs(251)));
    layer0_outputs(9094) <= (inputs(108)) or (inputs(164));
    layer0_outputs(9095) <= not(inputs(93));
    layer0_outputs(9096) <= (inputs(37)) or (inputs(89));
    layer0_outputs(9097) <= (inputs(172)) and not (inputs(244));
    layer0_outputs(9098) <= not(inputs(72)) or (inputs(87));
    layer0_outputs(9099) <= not((inputs(54)) or (inputs(234)));
    layer0_outputs(9100) <= inputs(57);
    layer0_outputs(9101) <= inputs(118);
    layer0_outputs(9102) <= not((inputs(127)) or (inputs(70)));
    layer0_outputs(9103) <= not((inputs(239)) xor (inputs(167)));
    layer0_outputs(9104) <= (inputs(187)) xor (inputs(197));
    layer0_outputs(9105) <= not(inputs(213)) or (inputs(23));
    layer0_outputs(9106) <= (inputs(72)) or (inputs(130));
    layer0_outputs(9107) <= not((inputs(166)) xor (inputs(135)));
    layer0_outputs(9108) <= (inputs(9)) or (inputs(1));
    layer0_outputs(9109) <= (inputs(172)) and not (inputs(45));
    layer0_outputs(9110) <= (inputs(160)) or (inputs(0));
    layer0_outputs(9111) <= (inputs(215)) or (inputs(182));
    layer0_outputs(9112) <= (inputs(127)) and not (inputs(14));
    layer0_outputs(9113) <= (inputs(69)) or (inputs(81));
    layer0_outputs(9114) <= inputs(91);
    layer0_outputs(9115) <= '1';
    layer0_outputs(9116) <= not((inputs(51)) xor (inputs(137)));
    layer0_outputs(9117) <= not(inputs(133)) or (inputs(230));
    layer0_outputs(9118) <= (inputs(250)) or (inputs(188));
    layer0_outputs(9119) <= not((inputs(135)) xor (inputs(147)));
    layer0_outputs(9120) <= not((inputs(236)) or (inputs(23)));
    layer0_outputs(9121) <= (inputs(202)) and not (inputs(111));
    layer0_outputs(9122) <= not(inputs(216));
    layer0_outputs(9123) <= not((inputs(163)) xor (inputs(21)));
    layer0_outputs(9124) <= inputs(94);
    layer0_outputs(9125) <= (inputs(237)) and not (inputs(136));
    layer0_outputs(9126) <= (inputs(39)) and not (inputs(63));
    layer0_outputs(9127) <= not((inputs(131)) xor (inputs(50)));
    layer0_outputs(9128) <= (inputs(238)) or (inputs(37));
    layer0_outputs(9129) <= (inputs(73)) and not (inputs(125));
    layer0_outputs(9130) <= not((inputs(31)) or (inputs(42)));
    layer0_outputs(9131) <= not(inputs(216)) or (inputs(45));
    layer0_outputs(9132) <= not(inputs(152));
    layer0_outputs(9133) <= not(inputs(170)) or (inputs(165));
    layer0_outputs(9134) <= (inputs(188)) and not (inputs(26));
    layer0_outputs(9135) <= (inputs(173)) xor (inputs(21));
    layer0_outputs(9136) <= not((inputs(104)) or (inputs(160)));
    layer0_outputs(9137) <= not((inputs(183)) xor (inputs(147)));
    layer0_outputs(9138) <= not(inputs(89));
    layer0_outputs(9139) <= inputs(238);
    layer0_outputs(9140) <= not(inputs(6));
    layer0_outputs(9141) <= not(inputs(139)) or (inputs(111));
    layer0_outputs(9142) <= not(inputs(171));
    layer0_outputs(9143) <= not(inputs(102)) or (inputs(140));
    layer0_outputs(9144) <= (inputs(143)) or (inputs(89));
    layer0_outputs(9145) <= (inputs(84)) and not (inputs(230));
    layer0_outputs(9146) <= not(inputs(176));
    layer0_outputs(9147) <= (inputs(212)) xor (inputs(33));
    layer0_outputs(9148) <= (inputs(129)) or (inputs(46));
    layer0_outputs(9149) <= not((inputs(104)) xor (inputs(176)));
    layer0_outputs(9150) <= (inputs(156)) xor (inputs(213));
    layer0_outputs(9151) <= (inputs(184)) xor (inputs(5));
    layer0_outputs(9152) <= inputs(13);
    layer0_outputs(9153) <= (inputs(68)) or (inputs(146));
    layer0_outputs(9154) <= not(inputs(3)) or (inputs(25));
    layer0_outputs(9155) <= (inputs(126)) or (inputs(38));
    layer0_outputs(9156) <= (inputs(84)) xor (inputs(243));
    layer0_outputs(9157) <= not(inputs(32));
    layer0_outputs(9158) <= (inputs(157)) xor (inputs(52));
    layer0_outputs(9159) <= not((inputs(48)) xor (inputs(109)));
    layer0_outputs(9160) <= (inputs(74)) and not (inputs(52));
    layer0_outputs(9161) <= (inputs(5)) or (inputs(226));
    layer0_outputs(9162) <= not(inputs(167)) or (inputs(226));
    layer0_outputs(9163) <= not((inputs(200)) xor (inputs(92)));
    layer0_outputs(9164) <= not((inputs(171)) or (inputs(145)));
    layer0_outputs(9165) <= inputs(15);
    layer0_outputs(9166) <= (inputs(91)) xor (inputs(64));
    layer0_outputs(9167) <= '1';
    layer0_outputs(9168) <= inputs(101);
    layer0_outputs(9169) <= not(inputs(210)) or (inputs(74));
    layer0_outputs(9170) <= (inputs(31)) and not (inputs(1));
    layer0_outputs(9171) <= not((inputs(91)) xor (inputs(149)));
    layer0_outputs(9172) <= (inputs(26)) and (inputs(245));
    layer0_outputs(9173) <= inputs(80);
    layer0_outputs(9174) <= not(inputs(105)) or (inputs(83));
    layer0_outputs(9175) <= not(inputs(187));
    layer0_outputs(9176) <= '0';
    layer0_outputs(9177) <= not(inputs(132));
    layer0_outputs(9178) <= not(inputs(243));
    layer0_outputs(9179) <= inputs(121);
    layer0_outputs(9180) <= not(inputs(208)) or (inputs(131));
    layer0_outputs(9181) <= not(inputs(136));
    layer0_outputs(9182) <= not(inputs(102));
    layer0_outputs(9183) <= (inputs(153)) xor (inputs(16));
    layer0_outputs(9184) <= not((inputs(134)) and (inputs(78)));
    layer0_outputs(9185) <= (inputs(25)) and (inputs(53));
    layer0_outputs(9186) <= not((inputs(131)) xor (inputs(136)));
    layer0_outputs(9187) <= not(inputs(165));
    layer0_outputs(9188) <= (inputs(54)) or (inputs(14));
    layer0_outputs(9189) <= (inputs(127)) and not (inputs(46));
    layer0_outputs(9190) <= (inputs(202)) and not (inputs(101));
    layer0_outputs(9191) <= inputs(144);
    layer0_outputs(9192) <= not((inputs(169)) or (inputs(179)));
    layer0_outputs(9193) <= (inputs(204)) or (inputs(163));
    layer0_outputs(9194) <= not((inputs(132)) xor (inputs(108)));
    layer0_outputs(9195) <= (inputs(201)) and not (inputs(220));
    layer0_outputs(9196) <= not(inputs(103));
    layer0_outputs(9197) <= not((inputs(52)) and (inputs(46)));
    layer0_outputs(9198) <= '0';
    layer0_outputs(9199) <= inputs(64);
    layer0_outputs(9200) <= not(inputs(182));
    layer0_outputs(9201) <= '1';
    layer0_outputs(9202) <= inputs(101);
    layer0_outputs(9203) <= (inputs(43)) and not (inputs(30));
    layer0_outputs(9204) <= not(inputs(26)) or (inputs(47));
    layer0_outputs(9205) <= (inputs(187)) and not (inputs(61));
    layer0_outputs(9206) <= not((inputs(141)) xor (inputs(8)));
    layer0_outputs(9207) <= inputs(38);
    layer0_outputs(9208) <= not((inputs(130)) or (inputs(149)));
    layer0_outputs(9209) <= inputs(120);
    layer0_outputs(9210) <= not(inputs(239)) or (inputs(218));
    layer0_outputs(9211) <= inputs(78);
    layer0_outputs(9212) <= inputs(212);
    layer0_outputs(9213) <= not(inputs(32)) or (inputs(222));
    layer0_outputs(9214) <= not((inputs(203)) or (inputs(104)));
    layer0_outputs(9215) <= not(inputs(177));
    layer0_outputs(9216) <= not(inputs(153)) or (inputs(235));
    layer0_outputs(9217) <= not(inputs(72)) or (inputs(195));
    layer0_outputs(9218) <= (inputs(29)) and not (inputs(75));
    layer0_outputs(9219) <= (inputs(44)) and not (inputs(147));
    layer0_outputs(9220) <= inputs(230);
    layer0_outputs(9221) <= (inputs(112)) or (inputs(43));
    layer0_outputs(9222) <= not((inputs(191)) or (inputs(115)));
    layer0_outputs(9223) <= (inputs(134)) xor (inputs(150));
    layer0_outputs(9224) <= not(inputs(65)) or (inputs(212));
    layer0_outputs(9225) <= not((inputs(115)) or (inputs(165)));
    layer0_outputs(9226) <= not((inputs(101)) or (inputs(130)));
    layer0_outputs(9227) <= not(inputs(120)) or (inputs(225));
    layer0_outputs(9228) <= (inputs(197)) xor (inputs(78));
    layer0_outputs(9229) <= (inputs(42)) and not (inputs(96));
    layer0_outputs(9230) <= inputs(122);
    layer0_outputs(9231) <= not((inputs(26)) and (inputs(154)));
    layer0_outputs(9232) <= not((inputs(158)) xor (inputs(51)));
    layer0_outputs(9233) <= inputs(184);
    layer0_outputs(9234) <= inputs(62);
    layer0_outputs(9235) <= not(inputs(70)) or (inputs(159));
    layer0_outputs(9236) <= not(inputs(10));
    layer0_outputs(9237) <= (inputs(147)) and not (inputs(217));
    layer0_outputs(9238) <= inputs(151);
    layer0_outputs(9239) <= not((inputs(162)) or (inputs(48)));
    layer0_outputs(9240) <= not(inputs(41));
    layer0_outputs(9241) <= inputs(189);
    layer0_outputs(9242) <= not((inputs(68)) or (inputs(215)));
    layer0_outputs(9243) <= (inputs(137)) and not (inputs(49));
    layer0_outputs(9244) <= not(inputs(30));
    layer0_outputs(9245) <= not(inputs(72));
    layer0_outputs(9246) <= not((inputs(234)) xor (inputs(132)));
    layer0_outputs(9247) <= inputs(215);
    layer0_outputs(9248) <= not((inputs(212)) or (inputs(153)));
    layer0_outputs(9249) <= not(inputs(120));
    layer0_outputs(9250) <= not((inputs(88)) or (inputs(26)));
    layer0_outputs(9251) <= inputs(152);
    layer0_outputs(9252) <= (inputs(43)) and not (inputs(64));
    layer0_outputs(9253) <= (inputs(208)) xor (inputs(167));
    layer0_outputs(9254) <= (inputs(171)) and not (inputs(30));
    layer0_outputs(9255) <= inputs(234);
    layer0_outputs(9256) <= (inputs(130)) or (inputs(62));
    layer0_outputs(9257) <= not((inputs(248)) or (inputs(188)));
    layer0_outputs(9258) <= (inputs(160)) or (inputs(54));
    layer0_outputs(9259) <= not(inputs(8));
    layer0_outputs(9260) <= (inputs(112)) and not (inputs(21));
    layer0_outputs(9261) <= (inputs(1)) or (inputs(83));
    layer0_outputs(9262) <= not(inputs(211)) or (inputs(251));
    layer0_outputs(9263) <= not((inputs(219)) or (inputs(12)));
    layer0_outputs(9264) <= inputs(85);
    layer0_outputs(9265) <= not((inputs(20)) xor (inputs(40)));
    layer0_outputs(9266) <= (inputs(4)) or (inputs(22));
    layer0_outputs(9267) <= not(inputs(93));
    layer0_outputs(9268) <= (inputs(195)) and (inputs(209));
    layer0_outputs(9269) <= not((inputs(35)) xor (inputs(202)));
    layer0_outputs(9270) <= not((inputs(89)) or (inputs(235)));
    layer0_outputs(9271) <= (inputs(39)) and not (inputs(180));
    layer0_outputs(9272) <= not(inputs(21)) or (inputs(229));
    layer0_outputs(9273) <= not(inputs(121));
    layer0_outputs(9274) <= '0';
    layer0_outputs(9275) <= (inputs(255)) or (inputs(199));
    layer0_outputs(9276) <= not((inputs(115)) or (inputs(86)));
    layer0_outputs(9277) <= (inputs(189)) and (inputs(111));
    layer0_outputs(9278) <= not((inputs(88)) xor (inputs(156)));
    layer0_outputs(9279) <= not((inputs(150)) or (inputs(37)));
    layer0_outputs(9280) <= '0';
    layer0_outputs(9281) <= not(inputs(122)) or (inputs(183));
    layer0_outputs(9282) <= (inputs(78)) and not (inputs(103));
    layer0_outputs(9283) <= not((inputs(187)) or (inputs(197)));
    layer0_outputs(9284) <= (inputs(184)) xor (inputs(156));
    layer0_outputs(9285) <= inputs(137);
    layer0_outputs(9286) <= (inputs(207)) and not (inputs(249));
    layer0_outputs(9287) <= not((inputs(237)) or (inputs(69)));
    layer0_outputs(9288) <= not((inputs(57)) or (inputs(206)));
    layer0_outputs(9289) <= (inputs(3)) and not (inputs(207));
    layer0_outputs(9290) <= '0';
    layer0_outputs(9291) <= not(inputs(115));
    layer0_outputs(9292) <= not(inputs(37));
    layer0_outputs(9293) <= not(inputs(147));
    layer0_outputs(9294) <= inputs(25);
    layer0_outputs(9295) <= not(inputs(125));
    layer0_outputs(9296) <= inputs(138);
    layer0_outputs(9297) <= (inputs(74)) and not (inputs(58));
    layer0_outputs(9298) <= not((inputs(157)) xor (inputs(100)));
    layer0_outputs(9299) <= not(inputs(182));
    layer0_outputs(9300) <= inputs(249);
    layer0_outputs(9301) <= (inputs(217)) and not (inputs(44));
    layer0_outputs(9302) <= (inputs(118)) or (inputs(134));
    layer0_outputs(9303) <= (inputs(164)) xor (inputs(51));
    layer0_outputs(9304) <= not(inputs(223)) or (inputs(4));
    layer0_outputs(9305) <= inputs(173);
    layer0_outputs(9306) <= inputs(102);
    layer0_outputs(9307) <= inputs(130);
    layer0_outputs(9308) <= not(inputs(69)) or (inputs(116));
    layer0_outputs(9309) <= '0';
    layer0_outputs(9310) <= not((inputs(7)) xor (inputs(230)));
    layer0_outputs(9311) <= (inputs(218)) or (inputs(119));
    layer0_outputs(9312) <= (inputs(172)) or (inputs(125));
    layer0_outputs(9313) <= (inputs(90)) and not (inputs(109));
    layer0_outputs(9314) <= not(inputs(169));
    layer0_outputs(9315) <= (inputs(10)) or (inputs(211));
    layer0_outputs(9316) <= not(inputs(194)) or (inputs(143));
    layer0_outputs(9317) <= (inputs(118)) or (inputs(243));
    layer0_outputs(9318) <= (inputs(216)) and not (inputs(77));
    layer0_outputs(9319) <= (inputs(250)) and (inputs(86));
    layer0_outputs(9320) <= (inputs(167)) xor (inputs(27));
    layer0_outputs(9321) <= (inputs(7)) and not (inputs(159));
    layer0_outputs(9322) <= inputs(96);
    layer0_outputs(9323) <= (inputs(188)) or (inputs(37));
    layer0_outputs(9324) <= '0';
    layer0_outputs(9325) <= not(inputs(177)) or (inputs(122));
    layer0_outputs(9326) <= '1';
    layer0_outputs(9327) <= not(inputs(233));
    layer0_outputs(9328) <= not((inputs(231)) or (inputs(20)));
    layer0_outputs(9329) <= (inputs(41)) or (inputs(13));
    layer0_outputs(9330) <= not(inputs(109)) or (inputs(30));
    layer0_outputs(9331) <= (inputs(111)) and not (inputs(85));
    layer0_outputs(9332) <= (inputs(183)) and not (inputs(127));
    layer0_outputs(9333) <= not((inputs(101)) xor (inputs(110)));
    layer0_outputs(9334) <= not((inputs(81)) xor (inputs(216)));
    layer0_outputs(9335) <= (inputs(89)) xor (inputs(73));
    layer0_outputs(9336) <= (inputs(118)) and not (inputs(152));
    layer0_outputs(9337) <= not((inputs(54)) xor (inputs(172)));
    layer0_outputs(9338) <= (inputs(17)) xor (inputs(57));
    layer0_outputs(9339) <= (inputs(37)) xor (inputs(54));
    layer0_outputs(9340) <= inputs(6);
    layer0_outputs(9341) <= (inputs(235)) and not (inputs(52));
    layer0_outputs(9342) <= not(inputs(197)) or (inputs(21));
    layer0_outputs(9343) <= not(inputs(36));
    layer0_outputs(9344) <= (inputs(218)) and (inputs(198));
    layer0_outputs(9345) <= not((inputs(212)) or (inputs(251)));
    layer0_outputs(9346) <= (inputs(104)) and not (inputs(19));
    layer0_outputs(9347) <= (inputs(151)) and not (inputs(93));
    layer0_outputs(9348) <= (inputs(202)) or (inputs(12));
    layer0_outputs(9349) <= not((inputs(19)) or (inputs(93)));
    layer0_outputs(9350) <= '1';
    layer0_outputs(9351) <= not(inputs(249));
    layer0_outputs(9352) <= not((inputs(103)) xor (inputs(71)));
    layer0_outputs(9353) <= (inputs(150)) and not (inputs(185));
    layer0_outputs(9354) <= not((inputs(100)) or (inputs(59)));
    layer0_outputs(9355) <= not(inputs(86)) or (inputs(7));
    layer0_outputs(9356) <= not(inputs(29));
    layer0_outputs(9357) <= inputs(141);
    layer0_outputs(9358) <= not(inputs(1)) or (inputs(9));
    layer0_outputs(9359) <= not(inputs(123)) or (inputs(95));
    layer0_outputs(9360) <= not(inputs(164));
    layer0_outputs(9361) <= inputs(171);
    layer0_outputs(9362) <= inputs(151);
    layer0_outputs(9363) <= '0';
    layer0_outputs(9364) <= not(inputs(196));
    layer0_outputs(9365) <= not((inputs(233)) and (inputs(53)));
    layer0_outputs(9366) <= not(inputs(11));
    layer0_outputs(9367) <= inputs(72);
    layer0_outputs(9368) <= not((inputs(245)) xor (inputs(8)));
    layer0_outputs(9369) <= not((inputs(239)) or (inputs(74)));
    layer0_outputs(9370) <= (inputs(148)) xor (inputs(143));
    layer0_outputs(9371) <= not((inputs(123)) xor (inputs(12)));
    layer0_outputs(9372) <= not(inputs(171)) or (inputs(167));
    layer0_outputs(9373) <= not((inputs(21)) xor (inputs(247)));
    layer0_outputs(9374) <= not(inputs(142)) or (inputs(151));
    layer0_outputs(9375) <= not((inputs(233)) or (inputs(37)));
    layer0_outputs(9376) <= '0';
    layer0_outputs(9377) <= not(inputs(110));
    layer0_outputs(9378) <= not((inputs(83)) or (inputs(186)));
    layer0_outputs(9379) <= inputs(117);
    layer0_outputs(9380) <= not((inputs(181)) or (inputs(40)));
    layer0_outputs(9381) <= not((inputs(75)) and (inputs(13)));
    layer0_outputs(9382) <= (inputs(182)) or (inputs(97));
    layer0_outputs(9383) <= (inputs(74)) or (inputs(227));
    layer0_outputs(9384) <= not(inputs(187)) or (inputs(40));
    layer0_outputs(9385) <= (inputs(30)) and not (inputs(16));
    layer0_outputs(9386) <= (inputs(34)) xor (inputs(134));
    layer0_outputs(9387) <= (inputs(106)) and not (inputs(165));
    layer0_outputs(9388) <= not(inputs(0));
    layer0_outputs(9389) <= '0';
    layer0_outputs(9390) <= '1';
    layer0_outputs(9391) <= (inputs(9)) and (inputs(22));
    layer0_outputs(9392) <= not((inputs(165)) or (inputs(80)));
    layer0_outputs(9393) <= not(inputs(120));
    layer0_outputs(9394) <= not(inputs(121)) or (inputs(212));
    layer0_outputs(9395) <= (inputs(202)) xor (inputs(74));
    layer0_outputs(9396) <= not(inputs(131)) or (inputs(178));
    layer0_outputs(9397) <= inputs(135);
    layer0_outputs(9398) <= (inputs(211)) xor (inputs(215));
    layer0_outputs(9399) <= not((inputs(142)) xor (inputs(190)));
    layer0_outputs(9400) <= (inputs(238)) and (inputs(26));
    layer0_outputs(9401) <= not((inputs(211)) or (inputs(24)));
    layer0_outputs(9402) <= inputs(224);
    layer0_outputs(9403) <= not((inputs(21)) or (inputs(204)));
    layer0_outputs(9404) <= not(inputs(215)) or (inputs(14));
    layer0_outputs(9405) <= inputs(86);
    layer0_outputs(9406) <= not((inputs(249)) and (inputs(113)));
    layer0_outputs(9407) <= not(inputs(235)) or (inputs(143));
    layer0_outputs(9408) <= not((inputs(230)) xor (inputs(218)));
    layer0_outputs(9409) <= (inputs(231)) or (inputs(66));
    layer0_outputs(9410) <= '0';
    layer0_outputs(9411) <= not(inputs(66));
    layer0_outputs(9412) <= inputs(105);
    layer0_outputs(9413) <= (inputs(217)) or (inputs(125));
    layer0_outputs(9414) <= (inputs(168)) and not (inputs(73));
    layer0_outputs(9415) <= not(inputs(124)) or (inputs(9));
    layer0_outputs(9416) <= inputs(104);
    layer0_outputs(9417) <= not(inputs(182));
    layer0_outputs(9418) <= (inputs(218)) xor (inputs(184));
    layer0_outputs(9419) <= (inputs(46)) xor (inputs(211));
    layer0_outputs(9420) <= not((inputs(57)) xor (inputs(221)));
    layer0_outputs(9421) <= (inputs(222)) or (inputs(157));
    layer0_outputs(9422) <= not(inputs(184)) or (inputs(128));
    layer0_outputs(9423) <= inputs(135);
    layer0_outputs(9424) <= inputs(41);
    layer0_outputs(9425) <= not(inputs(166));
    layer0_outputs(9426) <= not(inputs(150));
    layer0_outputs(9427) <= (inputs(77)) xor (inputs(200));
    layer0_outputs(9428) <= not((inputs(82)) or (inputs(182)));
    layer0_outputs(9429) <= not((inputs(37)) or (inputs(90)));
    layer0_outputs(9430) <= (inputs(26)) and not (inputs(188));
    layer0_outputs(9431) <= not((inputs(5)) or (inputs(226)));
    layer0_outputs(9432) <= (inputs(162)) xor (inputs(140));
    layer0_outputs(9433) <= '0';
    layer0_outputs(9434) <= (inputs(174)) and not (inputs(24));
    layer0_outputs(9435) <= not((inputs(174)) or (inputs(147)));
    layer0_outputs(9436) <= not((inputs(202)) xor (inputs(17)));
    layer0_outputs(9437) <= (inputs(86)) and not (inputs(230));
    layer0_outputs(9438) <= (inputs(230)) xor (inputs(241));
    layer0_outputs(9439) <= not(inputs(119));
    layer0_outputs(9440) <= not(inputs(168));
    layer0_outputs(9441) <= not((inputs(145)) and (inputs(135)));
    layer0_outputs(9442) <= inputs(245);
    layer0_outputs(9443) <= not(inputs(73));
    layer0_outputs(9444) <= not((inputs(194)) or (inputs(196)));
    layer0_outputs(9445) <= not((inputs(240)) xor (inputs(86)));
    layer0_outputs(9446) <= not(inputs(169));
    layer0_outputs(9447) <= (inputs(171)) xor (inputs(86));
    layer0_outputs(9448) <= (inputs(138)) and not (inputs(243));
    layer0_outputs(9449) <= not(inputs(249)) or (inputs(158));
    layer0_outputs(9450) <= inputs(143);
    layer0_outputs(9451) <= (inputs(185)) and not (inputs(8));
    layer0_outputs(9452) <= not((inputs(109)) or (inputs(124)));
    layer0_outputs(9453) <= not((inputs(170)) or (inputs(155)));
    layer0_outputs(9454) <= not((inputs(93)) xor (inputs(252)));
    layer0_outputs(9455) <= (inputs(213)) and not (inputs(17));
    layer0_outputs(9456) <= not(inputs(214)) or (inputs(95));
    layer0_outputs(9457) <= not(inputs(179)) or (inputs(126));
    layer0_outputs(9458) <= '0';
    layer0_outputs(9459) <= not(inputs(136));
    layer0_outputs(9460) <= not(inputs(74)) or (inputs(229));
    layer0_outputs(9461) <= (inputs(199)) and not (inputs(159));
    layer0_outputs(9462) <= not(inputs(148)) or (inputs(95));
    layer0_outputs(9463) <= not(inputs(213)) or (inputs(206));
    layer0_outputs(9464) <= '0';
    layer0_outputs(9465) <= not(inputs(151)) or (inputs(227));
    layer0_outputs(9466) <= not(inputs(218)) or (inputs(249));
    layer0_outputs(9467) <= not(inputs(206));
    layer0_outputs(9468) <= not(inputs(60)) or (inputs(130));
    layer0_outputs(9469) <= not(inputs(189));
    layer0_outputs(9470) <= (inputs(10)) xor (inputs(168));
    layer0_outputs(9471) <= not(inputs(110)) or (inputs(203));
    layer0_outputs(9472) <= inputs(76);
    layer0_outputs(9473) <= not(inputs(102));
    layer0_outputs(9474) <= (inputs(40)) xor (inputs(222));
    layer0_outputs(9475) <= not((inputs(74)) or (inputs(226)));
    layer0_outputs(9476) <= (inputs(106)) and not (inputs(10));
    layer0_outputs(9477) <= (inputs(100)) and not (inputs(24));
    layer0_outputs(9478) <= (inputs(105)) and not (inputs(173));
    layer0_outputs(9479) <= not(inputs(31)) or (inputs(76));
    layer0_outputs(9480) <= not(inputs(36)) or (inputs(8));
    layer0_outputs(9481) <= not((inputs(103)) xor (inputs(11)));
    layer0_outputs(9482) <= (inputs(117)) and not (inputs(163));
    layer0_outputs(9483) <= not(inputs(12)) or (inputs(21));
    layer0_outputs(9484) <= (inputs(113)) or (inputs(103));
    layer0_outputs(9485) <= not(inputs(70));
    layer0_outputs(9486) <= (inputs(231)) and not (inputs(3));
    layer0_outputs(9487) <= inputs(151);
    layer0_outputs(9488) <= (inputs(244)) and not (inputs(34));
    layer0_outputs(9489) <= not(inputs(102)) or (inputs(151));
    layer0_outputs(9490) <= (inputs(198)) or (inputs(194));
    layer0_outputs(9491) <= inputs(99);
    layer0_outputs(9492) <= inputs(214);
    layer0_outputs(9493) <= not(inputs(167)) or (inputs(195));
    layer0_outputs(9494) <= not((inputs(20)) or (inputs(25)));
    layer0_outputs(9495) <= not(inputs(198));
    layer0_outputs(9496) <= (inputs(210)) and not (inputs(212));
    layer0_outputs(9497) <= not((inputs(236)) or (inputs(145)));
    layer0_outputs(9498) <= not((inputs(19)) and (inputs(49)));
    layer0_outputs(9499) <= (inputs(120)) and not (inputs(173));
    layer0_outputs(9500) <= not((inputs(196)) or (inputs(255)));
    layer0_outputs(9501) <= (inputs(115)) or (inputs(107));
    layer0_outputs(9502) <= (inputs(24)) and not (inputs(0));
    layer0_outputs(9503) <= (inputs(26)) xor (inputs(156));
    layer0_outputs(9504) <= not((inputs(87)) xor (inputs(14)));
    layer0_outputs(9505) <= (inputs(23)) and not (inputs(111));
    layer0_outputs(9506) <= not(inputs(248));
    layer0_outputs(9507) <= not(inputs(195)) or (inputs(67));
    layer0_outputs(9508) <= not(inputs(228)) or (inputs(206));
    layer0_outputs(9509) <= '1';
    layer0_outputs(9510) <= (inputs(16)) or (inputs(59));
    layer0_outputs(9511) <= (inputs(73)) or (inputs(93));
    layer0_outputs(9512) <= not(inputs(246));
    layer0_outputs(9513) <= (inputs(94)) or (inputs(187));
    layer0_outputs(9514) <= not(inputs(52)) or (inputs(13));
    layer0_outputs(9515) <= not((inputs(7)) and (inputs(161)));
    layer0_outputs(9516) <= not(inputs(105)) or (inputs(143));
    layer0_outputs(9517) <= not((inputs(205)) xor (inputs(224)));
    layer0_outputs(9518) <= not(inputs(190)) or (inputs(149));
    layer0_outputs(9519) <= not((inputs(225)) or (inputs(109)));
    layer0_outputs(9520) <= inputs(86);
    layer0_outputs(9521) <= not((inputs(69)) or (inputs(91)));
    layer0_outputs(9522) <= not(inputs(217)) or (inputs(210));
    layer0_outputs(9523) <= not(inputs(56));
    layer0_outputs(9524) <= (inputs(237)) and not (inputs(106));
    layer0_outputs(9525) <= not(inputs(102)) or (inputs(164));
    layer0_outputs(9526) <= inputs(252);
    layer0_outputs(9527) <= inputs(179);
    layer0_outputs(9528) <= not((inputs(167)) or (inputs(78)));
    layer0_outputs(9529) <= not(inputs(181)) or (inputs(144));
    layer0_outputs(9530) <= (inputs(220)) xor (inputs(52));
    layer0_outputs(9531) <= (inputs(58)) and (inputs(197));
    layer0_outputs(9532) <= not((inputs(79)) or (inputs(61)));
    layer0_outputs(9533) <= not((inputs(203)) xor (inputs(176)));
    layer0_outputs(9534) <= not(inputs(25));
    layer0_outputs(9535) <= not((inputs(212)) or (inputs(39)));
    layer0_outputs(9536) <= inputs(211);
    layer0_outputs(9537) <= (inputs(202)) or (inputs(116));
    layer0_outputs(9538) <= inputs(245);
    layer0_outputs(9539) <= inputs(181);
    layer0_outputs(9540) <= (inputs(102)) and not (inputs(194));
    layer0_outputs(9541) <= not(inputs(119)) or (inputs(141));
    layer0_outputs(9542) <= not(inputs(182));
    layer0_outputs(9543) <= not(inputs(91)) or (inputs(46));
    layer0_outputs(9544) <= (inputs(69)) xor (inputs(138));
    layer0_outputs(9545) <= inputs(124);
    layer0_outputs(9546) <= (inputs(153)) and not (inputs(126));
    layer0_outputs(9547) <= (inputs(242)) xor (inputs(201));
    layer0_outputs(9548) <= (inputs(39)) and not (inputs(243));
    layer0_outputs(9549) <= '0';
    layer0_outputs(9550) <= inputs(121);
    layer0_outputs(9551) <= (inputs(169)) or (inputs(190));
    layer0_outputs(9552) <= not((inputs(120)) xor (inputs(234)));
    layer0_outputs(9553) <= (inputs(110)) and not (inputs(14));
    layer0_outputs(9554) <= (inputs(176)) or (inputs(35));
    layer0_outputs(9555) <= inputs(67);
    layer0_outputs(9556) <= (inputs(53)) or (inputs(131));
    layer0_outputs(9557) <= inputs(83);
    layer0_outputs(9558) <= not((inputs(82)) or (inputs(181)));
    layer0_outputs(9559) <= inputs(34);
    layer0_outputs(9560) <= not((inputs(41)) or (inputs(116)));
    layer0_outputs(9561) <= not(inputs(193)) or (inputs(110));
    layer0_outputs(9562) <= not(inputs(60));
    layer0_outputs(9563) <= (inputs(49)) and (inputs(246));
    layer0_outputs(9564) <= not((inputs(206)) xor (inputs(88)));
    layer0_outputs(9565) <= (inputs(148)) and not (inputs(195));
    layer0_outputs(9566) <= not((inputs(55)) or (inputs(171)));
    layer0_outputs(9567) <= (inputs(197)) and not (inputs(248));
    layer0_outputs(9568) <= (inputs(119)) and not (inputs(87));
    layer0_outputs(9569) <= not((inputs(82)) or (inputs(72)));
    layer0_outputs(9570) <= '1';
    layer0_outputs(9571) <= '1';
    layer0_outputs(9572) <= not((inputs(82)) xor (inputs(226)));
    layer0_outputs(9573) <= (inputs(91)) and not (inputs(38));
    layer0_outputs(9574) <= not(inputs(13)) or (inputs(73));
    layer0_outputs(9575) <= not((inputs(83)) or (inputs(222)));
    layer0_outputs(9576) <= '0';
    layer0_outputs(9577) <= not(inputs(88));
    layer0_outputs(9578) <= not(inputs(40));
    layer0_outputs(9579) <= not((inputs(245)) or (inputs(134)));
    layer0_outputs(9580) <= not((inputs(52)) or (inputs(233)));
    layer0_outputs(9581) <= (inputs(200)) and not (inputs(146));
    layer0_outputs(9582) <= (inputs(73)) or (inputs(109));
    layer0_outputs(9583) <= (inputs(142)) or (inputs(127));
    layer0_outputs(9584) <= not(inputs(144));
    layer0_outputs(9585) <= (inputs(214)) or (inputs(96));
    layer0_outputs(9586) <= not((inputs(92)) xor (inputs(113)));
    layer0_outputs(9587) <= not(inputs(102));
    layer0_outputs(9588) <= (inputs(140)) and not (inputs(16));
    layer0_outputs(9589) <= not(inputs(151));
    layer0_outputs(9590) <= (inputs(131)) or (inputs(194));
    layer0_outputs(9591) <= inputs(178);
    layer0_outputs(9592) <= inputs(76);
    layer0_outputs(9593) <= (inputs(47)) and (inputs(127));
    layer0_outputs(9594) <= inputs(170);
    layer0_outputs(9595) <= '1';
    layer0_outputs(9596) <= not((inputs(187)) and (inputs(74)));
    layer0_outputs(9597) <= inputs(146);
    layer0_outputs(9598) <= not((inputs(209)) or (inputs(214)));
    layer0_outputs(9599) <= (inputs(171)) and not (inputs(220));
    layer0_outputs(9600) <= '1';
    layer0_outputs(9601) <= not(inputs(166)) or (inputs(26));
    layer0_outputs(9602) <= not(inputs(46)) or (inputs(25));
    layer0_outputs(9603) <= (inputs(188)) and (inputs(35));
    layer0_outputs(9604) <= not((inputs(173)) xor (inputs(75)));
    layer0_outputs(9605) <= not(inputs(153)) or (inputs(120));
    layer0_outputs(9606) <= '0';
    layer0_outputs(9607) <= (inputs(93)) or (inputs(87));
    layer0_outputs(9608) <= not((inputs(235)) xor (inputs(217)));
    layer0_outputs(9609) <= (inputs(105)) and (inputs(137));
    layer0_outputs(9610) <= not(inputs(178));
    layer0_outputs(9611) <= not(inputs(25)) or (inputs(211));
    layer0_outputs(9612) <= (inputs(246)) and not (inputs(18));
    layer0_outputs(9613) <= not((inputs(232)) or (inputs(132)));
    layer0_outputs(9614) <= not((inputs(220)) or (inputs(100)));
    layer0_outputs(9615) <= inputs(177);
    layer0_outputs(9616) <= (inputs(188)) or (inputs(241));
    layer0_outputs(9617) <= (inputs(102)) xor (inputs(87));
    layer0_outputs(9618) <= inputs(187);
    layer0_outputs(9619) <= not((inputs(167)) or (inputs(172)));
    layer0_outputs(9620) <= (inputs(173)) xor (inputs(189));
    layer0_outputs(9621) <= not(inputs(181));
    layer0_outputs(9622) <= (inputs(230)) and not (inputs(223));
    layer0_outputs(9623) <= inputs(100);
    layer0_outputs(9624) <= inputs(217);
    layer0_outputs(9625) <= (inputs(61)) or (inputs(133));
    layer0_outputs(9626) <= not((inputs(236)) xor (inputs(87)));
    layer0_outputs(9627) <= (inputs(244)) and (inputs(110));
    layer0_outputs(9628) <= not(inputs(116)) or (inputs(24));
    layer0_outputs(9629) <= not(inputs(198));
    layer0_outputs(9630) <= not(inputs(85)) or (inputs(32));
    layer0_outputs(9631) <= not((inputs(47)) or (inputs(201)));
    layer0_outputs(9632) <= (inputs(210)) and not (inputs(130));
    layer0_outputs(9633) <= inputs(89);
    layer0_outputs(9634) <= (inputs(73)) and not (inputs(201));
    layer0_outputs(9635) <= not(inputs(130)) or (inputs(194));
    layer0_outputs(9636) <= not(inputs(254));
    layer0_outputs(9637) <= inputs(218);
    layer0_outputs(9638) <= (inputs(141)) or (inputs(6));
    layer0_outputs(9639) <= (inputs(236)) and not (inputs(66));
    layer0_outputs(9640) <= not(inputs(154));
    layer0_outputs(9641) <= inputs(131);
    layer0_outputs(9642) <= not((inputs(104)) or (inputs(55)));
    layer0_outputs(9643) <= not((inputs(42)) xor (inputs(69)));
    layer0_outputs(9644) <= inputs(215);
    layer0_outputs(9645) <= not(inputs(8)) or (inputs(166));
    layer0_outputs(9646) <= (inputs(63)) and (inputs(20));
    layer0_outputs(9647) <= not(inputs(223)) or (inputs(144));
    layer0_outputs(9648) <= (inputs(132)) xor (inputs(149));
    layer0_outputs(9649) <= not(inputs(72)) or (inputs(14));
    layer0_outputs(9650) <= not(inputs(118)) or (inputs(205));
    layer0_outputs(9651) <= not((inputs(29)) and (inputs(160)));
    layer0_outputs(9652) <= not((inputs(216)) xor (inputs(103)));
    layer0_outputs(9653) <= not(inputs(26));
    layer0_outputs(9654) <= not((inputs(220)) or (inputs(179)));
    layer0_outputs(9655) <= not(inputs(41));
    layer0_outputs(9656) <= (inputs(17)) or (inputs(77));
    layer0_outputs(9657) <= inputs(113);
    layer0_outputs(9658) <= (inputs(124)) and not (inputs(1));
    layer0_outputs(9659) <= not(inputs(185));
    layer0_outputs(9660) <= not((inputs(157)) or (inputs(42)));
    layer0_outputs(9661) <= (inputs(175)) xor (inputs(28));
    layer0_outputs(9662) <= not(inputs(94));
    layer0_outputs(9663) <= (inputs(200)) and not (inputs(114));
    layer0_outputs(9664) <= '0';
    layer0_outputs(9665) <= inputs(106);
    layer0_outputs(9666) <= (inputs(211)) xor (inputs(196));
    layer0_outputs(9667) <= not(inputs(107)) or (inputs(39));
    layer0_outputs(9668) <= inputs(3);
    layer0_outputs(9669) <= '1';
    layer0_outputs(9670) <= '0';
    layer0_outputs(9671) <= (inputs(32)) xor (inputs(174));
    layer0_outputs(9672) <= not(inputs(162)) or (inputs(160));
    layer0_outputs(9673) <= not(inputs(87));
    layer0_outputs(9674) <= (inputs(44)) and not (inputs(4));
    layer0_outputs(9675) <= not(inputs(186));
    layer0_outputs(9676) <= '1';
    layer0_outputs(9677) <= not((inputs(43)) xor (inputs(6)));
    layer0_outputs(9678) <= (inputs(67)) or (inputs(225));
    layer0_outputs(9679) <= (inputs(14)) and not (inputs(35));
    layer0_outputs(9680) <= not((inputs(99)) xor (inputs(214)));
    layer0_outputs(9681) <= (inputs(33)) and not (inputs(77));
    layer0_outputs(9682) <= (inputs(47)) xor (inputs(230));
    layer0_outputs(9683) <= not(inputs(183));
    layer0_outputs(9684) <= not((inputs(253)) xor (inputs(125)));
    layer0_outputs(9685) <= (inputs(195)) or (inputs(179));
    layer0_outputs(9686) <= (inputs(33)) xor (inputs(252));
    layer0_outputs(9687) <= not(inputs(187)) or (inputs(114));
    layer0_outputs(9688) <= not(inputs(101));
    layer0_outputs(9689) <= not((inputs(91)) or (inputs(228)));
    layer0_outputs(9690) <= not((inputs(116)) or (inputs(106)));
    layer0_outputs(9691) <= (inputs(136)) or (inputs(36));
    layer0_outputs(9692) <= inputs(150);
    layer0_outputs(9693) <= not((inputs(24)) xor (inputs(52)));
    layer0_outputs(9694) <= inputs(199);
    layer0_outputs(9695) <= not((inputs(4)) and (inputs(10)));
    layer0_outputs(9696) <= not(inputs(56));
    layer0_outputs(9697) <= not(inputs(119)) or (inputs(236));
    layer0_outputs(9698) <= (inputs(191)) or (inputs(86));
    layer0_outputs(9699) <= (inputs(98)) xor (inputs(4));
    layer0_outputs(9700) <= inputs(184);
    layer0_outputs(9701) <= not((inputs(120)) or (inputs(127)));
    layer0_outputs(9702) <= not((inputs(175)) and (inputs(159)));
    layer0_outputs(9703) <= not((inputs(15)) xor (inputs(123)));
    layer0_outputs(9704) <= '0';
    layer0_outputs(9705) <= not(inputs(79)) or (inputs(220));
    layer0_outputs(9706) <= (inputs(113)) or (inputs(232));
    layer0_outputs(9707) <= '0';
    layer0_outputs(9708) <= inputs(180);
    layer0_outputs(9709) <= not(inputs(188));
    layer0_outputs(9710) <= not((inputs(53)) or (inputs(24)));
    layer0_outputs(9711) <= not((inputs(136)) xor (inputs(34)));
    layer0_outputs(9712) <= (inputs(193)) xor (inputs(56));
    layer0_outputs(9713) <= (inputs(170)) and not (inputs(61));
    layer0_outputs(9714) <= not((inputs(161)) or (inputs(104)));
    layer0_outputs(9715) <= (inputs(79)) and not (inputs(49));
    layer0_outputs(9716) <= not((inputs(245)) xor (inputs(58)));
    layer0_outputs(9717) <= not((inputs(151)) xor (inputs(152)));
    layer0_outputs(9718) <= not(inputs(199));
    layer0_outputs(9719) <= (inputs(128)) and not (inputs(11));
    layer0_outputs(9720) <= inputs(166);
    layer0_outputs(9721) <= '1';
    layer0_outputs(9722) <= not((inputs(61)) xor (inputs(112)));
    layer0_outputs(9723) <= '0';
    layer0_outputs(9724) <= (inputs(167)) xor (inputs(64));
    layer0_outputs(9725) <= inputs(116);
    layer0_outputs(9726) <= '0';
    layer0_outputs(9727) <= not((inputs(131)) xor (inputs(254)));
    layer0_outputs(9728) <= (inputs(169)) and not (inputs(5));
    layer0_outputs(9729) <= inputs(19);
    layer0_outputs(9730) <= not(inputs(94)) or (inputs(141));
    layer0_outputs(9731) <= not(inputs(140)) or (inputs(146));
    layer0_outputs(9732) <= not(inputs(246));
    layer0_outputs(9733) <= not((inputs(241)) or (inputs(241)));
    layer0_outputs(9734) <= not((inputs(71)) xor (inputs(138)));
    layer0_outputs(9735) <= (inputs(28)) xor (inputs(58));
    layer0_outputs(9736) <= not(inputs(135)) or (inputs(249));
    layer0_outputs(9737) <= not(inputs(127)) or (inputs(31));
    layer0_outputs(9738) <= (inputs(32)) xor (inputs(168));
    layer0_outputs(9739) <= not((inputs(228)) or (inputs(108)));
    layer0_outputs(9740) <= inputs(206);
    layer0_outputs(9741) <= (inputs(39)) or (inputs(67));
    layer0_outputs(9742) <= (inputs(214)) and not (inputs(140));
    layer0_outputs(9743) <= (inputs(176)) or (inputs(75));
    layer0_outputs(9744) <= '1';
    layer0_outputs(9745) <= (inputs(162)) and (inputs(220));
    layer0_outputs(9746) <= (inputs(188)) and not (inputs(82));
    layer0_outputs(9747) <= not((inputs(255)) xor (inputs(138)));
    layer0_outputs(9748) <= not(inputs(135)) or (inputs(95));
    layer0_outputs(9749) <= not(inputs(93)) or (inputs(156));
    layer0_outputs(9750) <= (inputs(247)) and (inputs(61));
    layer0_outputs(9751) <= not(inputs(89)) or (inputs(10));
    layer0_outputs(9752) <= not((inputs(94)) xor (inputs(18)));
    layer0_outputs(9753) <= (inputs(140)) xor (inputs(138));
    layer0_outputs(9754) <= '1';
    layer0_outputs(9755) <= (inputs(181)) and not (inputs(78));
    layer0_outputs(9756) <= not((inputs(5)) or (inputs(227)));
    layer0_outputs(9757) <= '1';
    layer0_outputs(9758) <= inputs(128);
    layer0_outputs(9759) <= not(inputs(216));
    layer0_outputs(9760) <= inputs(58);
    layer0_outputs(9761) <= (inputs(226)) xor (inputs(151));
    layer0_outputs(9762) <= (inputs(11)) and not (inputs(175));
    layer0_outputs(9763) <= (inputs(92)) and not (inputs(99));
    layer0_outputs(9764) <= (inputs(242)) and not (inputs(248));
    layer0_outputs(9765) <= not((inputs(233)) xor (inputs(11)));
    layer0_outputs(9766) <= not((inputs(56)) xor (inputs(55)));
    layer0_outputs(9767) <= (inputs(106)) and not (inputs(246));
    layer0_outputs(9768) <= not((inputs(235)) xor (inputs(10)));
    layer0_outputs(9769) <= not(inputs(126));
    layer0_outputs(9770) <= not(inputs(118));
    layer0_outputs(9771) <= not((inputs(219)) xor (inputs(165)));
    layer0_outputs(9772) <= (inputs(74)) or (inputs(192));
    layer0_outputs(9773) <= (inputs(123)) or (inputs(22));
    layer0_outputs(9774) <= (inputs(67)) xor (inputs(22));
    layer0_outputs(9775) <= inputs(136);
    layer0_outputs(9776) <= not(inputs(148)) or (inputs(242));
    layer0_outputs(9777) <= (inputs(84)) and not (inputs(74));
    layer0_outputs(9778) <= not((inputs(200)) and (inputs(199)));
    layer0_outputs(9779) <= '0';
    layer0_outputs(9780) <= not(inputs(69));
    layer0_outputs(9781) <= (inputs(180)) and not (inputs(254));
    layer0_outputs(9782) <= (inputs(60)) xor (inputs(254));
    layer0_outputs(9783) <= not(inputs(171));
    layer0_outputs(9784) <= not((inputs(147)) or (inputs(39)));
    layer0_outputs(9785) <= (inputs(76)) and not (inputs(129));
    layer0_outputs(9786) <= not(inputs(91));
    layer0_outputs(9787) <= (inputs(235)) and not (inputs(9));
    layer0_outputs(9788) <= not(inputs(97)) or (inputs(251));
    layer0_outputs(9789) <= not(inputs(32)) or (inputs(78));
    layer0_outputs(9790) <= not(inputs(125)) or (inputs(97));
    layer0_outputs(9791) <= not(inputs(85));
    layer0_outputs(9792) <= (inputs(201)) or (inputs(206));
    layer0_outputs(9793) <= not((inputs(201)) or (inputs(18)));
    layer0_outputs(9794) <= not((inputs(98)) or (inputs(148)));
    layer0_outputs(9795) <= not(inputs(127)) or (inputs(48));
    layer0_outputs(9796) <= not((inputs(97)) and (inputs(235)));
    layer0_outputs(9797) <= inputs(242);
    layer0_outputs(9798) <= not((inputs(214)) xor (inputs(185)));
    layer0_outputs(9799) <= (inputs(210)) xor (inputs(240));
    layer0_outputs(9800) <= (inputs(50)) and not (inputs(63));
    layer0_outputs(9801) <= not(inputs(100));
    layer0_outputs(9802) <= not((inputs(13)) xor (inputs(32)));
    layer0_outputs(9803) <= not(inputs(101)) or (inputs(88));
    layer0_outputs(9804) <= not(inputs(58)) or (inputs(109));
    layer0_outputs(9805) <= inputs(230);
    layer0_outputs(9806) <= not(inputs(34));
    layer0_outputs(9807) <= inputs(141);
    layer0_outputs(9808) <= not((inputs(208)) and (inputs(185)));
    layer0_outputs(9809) <= (inputs(98)) or (inputs(202));
    layer0_outputs(9810) <= not(inputs(171)) or (inputs(50));
    layer0_outputs(9811) <= not((inputs(172)) xor (inputs(48)));
    layer0_outputs(9812) <= not((inputs(178)) or (inputs(61)));
    layer0_outputs(9813) <= (inputs(87)) xor (inputs(24));
    layer0_outputs(9814) <= not((inputs(105)) xor (inputs(10)));
    layer0_outputs(9815) <= inputs(106);
    layer0_outputs(9816) <= not(inputs(0)) or (inputs(244));
    layer0_outputs(9817) <= not((inputs(156)) or (inputs(163)));
    layer0_outputs(9818) <= (inputs(216)) xor (inputs(177));
    layer0_outputs(9819) <= not(inputs(133)) or (inputs(69));
    layer0_outputs(9820) <= (inputs(154)) or (inputs(38));
    layer0_outputs(9821) <= '0';
    layer0_outputs(9822) <= not((inputs(92)) or (inputs(60)));
    layer0_outputs(9823) <= (inputs(178)) xor (inputs(232));
    layer0_outputs(9824) <= inputs(181);
    layer0_outputs(9825) <= not((inputs(0)) or (inputs(75)));
    layer0_outputs(9826) <= not(inputs(67));
    layer0_outputs(9827) <= (inputs(161)) and (inputs(142));
    layer0_outputs(9828) <= (inputs(202)) and (inputs(8));
    layer0_outputs(9829) <= (inputs(155)) xor (inputs(96));
    layer0_outputs(9830) <= inputs(184);
    layer0_outputs(9831) <= inputs(118);
    layer0_outputs(9832) <= not(inputs(47)) or (inputs(51));
    layer0_outputs(9833) <= not(inputs(186)) or (inputs(90));
    layer0_outputs(9834) <= (inputs(166)) or (inputs(28));
    layer0_outputs(9835) <= (inputs(141)) or (inputs(83));
    layer0_outputs(9836) <= (inputs(145)) or (inputs(103));
    layer0_outputs(9837) <= not((inputs(128)) xor (inputs(23)));
    layer0_outputs(9838) <= '0';
    layer0_outputs(9839) <= not(inputs(214));
    layer0_outputs(9840) <= '1';
    layer0_outputs(9841) <= not(inputs(27)) or (inputs(35));
    layer0_outputs(9842) <= not(inputs(151));
    layer0_outputs(9843) <= (inputs(189)) or (inputs(147));
    layer0_outputs(9844) <= (inputs(165)) and not (inputs(219));
    layer0_outputs(9845) <= '0';
    layer0_outputs(9846) <= (inputs(121)) and not (inputs(173));
    layer0_outputs(9847) <= inputs(180);
    layer0_outputs(9848) <= (inputs(144)) and not (inputs(25));
    layer0_outputs(9849) <= (inputs(183)) and not (inputs(81));
    layer0_outputs(9850) <= inputs(23);
    layer0_outputs(9851) <= (inputs(152)) and not (inputs(124));
    layer0_outputs(9852) <= '0';
    layer0_outputs(9853) <= (inputs(89)) xor (inputs(175));
    layer0_outputs(9854) <= (inputs(249)) and not (inputs(238));
    layer0_outputs(9855) <= inputs(92);
    layer0_outputs(9856) <= (inputs(124)) xor (inputs(119));
    layer0_outputs(9857) <= (inputs(210)) xor (inputs(110));
    layer0_outputs(9858) <= not(inputs(239)) or (inputs(226));
    layer0_outputs(9859) <= not((inputs(133)) xor (inputs(146)));
    layer0_outputs(9860) <= (inputs(176)) or (inputs(35));
    layer0_outputs(9861) <= not(inputs(139));
    layer0_outputs(9862) <= not(inputs(132));
    layer0_outputs(9863) <= not((inputs(204)) or (inputs(84)));
    layer0_outputs(9864) <= not(inputs(24));
    layer0_outputs(9865) <= inputs(163);
    layer0_outputs(9866) <= not((inputs(211)) xor (inputs(245)));
    layer0_outputs(9867) <= '0';
    layer0_outputs(9868) <= not((inputs(150)) or (inputs(245)));
    layer0_outputs(9869) <= not((inputs(104)) or (inputs(54)));
    layer0_outputs(9870) <= not((inputs(15)) xor (inputs(180)));
    layer0_outputs(9871) <= not((inputs(86)) or (inputs(12)));
    layer0_outputs(9872) <= not(inputs(116));
    layer0_outputs(9873) <= (inputs(230)) xor (inputs(175));
    layer0_outputs(9874) <= inputs(108);
    layer0_outputs(9875) <= (inputs(14)) and (inputs(129));
    layer0_outputs(9876) <= inputs(169);
    layer0_outputs(9877) <= (inputs(127)) xor (inputs(40));
    layer0_outputs(9878) <= not(inputs(50)) or (inputs(146));
    layer0_outputs(9879) <= (inputs(45)) and not (inputs(111));
    layer0_outputs(9880) <= (inputs(78)) or (inputs(179));
    layer0_outputs(9881) <= '1';
    layer0_outputs(9882) <= (inputs(215)) xor (inputs(119));
    layer0_outputs(9883) <= inputs(192);
    layer0_outputs(9884) <= (inputs(47)) or (inputs(178));
    layer0_outputs(9885) <= not(inputs(93));
    layer0_outputs(9886) <= (inputs(97)) or (inputs(186));
    layer0_outputs(9887) <= inputs(181);
    layer0_outputs(9888) <= inputs(49);
    layer0_outputs(9889) <= not(inputs(179));
    layer0_outputs(9890) <= (inputs(255)) and not (inputs(236));
    layer0_outputs(9891) <= (inputs(88)) xor (inputs(14));
    layer0_outputs(9892) <= (inputs(0)) and (inputs(112));
    layer0_outputs(9893) <= (inputs(67)) and not (inputs(233));
    layer0_outputs(9894) <= not((inputs(31)) or (inputs(234)));
    layer0_outputs(9895) <= (inputs(85)) and not (inputs(44));
    layer0_outputs(9896) <= inputs(242);
    layer0_outputs(9897) <= not(inputs(86)) or (inputs(142));
    layer0_outputs(9898) <= (inputs(20)) and not (inputs(200));
    layer0_outputs(9899) <= (inputs(38)) and not (inputs(177));
    layer0_outputs(9900) <= not(inputs(100)) or (inputs(156));
    layer0_outputs(9901) <= not(inputs(88));
    layer0_outputs(9902) <= not(inputs(85)) or (inputs(183));
    layer0_outputs(9903) <= not((inputs(88)) xor (inputs(76)));
    layer0_outputs(9904) <= inputs(41);
    layer0_outputs(9905) <= not(inputs(2)) or (inputs(11));
    layer0_outputs(9906) <= (inputs(157)) or (inputs(45));
    layer0_outputs(9907) <= '1';
    layer0_outputs(9908) <= not(inputs(106));
    layer0_outputs(9909) <= (inputs(68)) and not (inputs(160));
    layer0_outputs(9910) <= not(inputs(213)) or (inputs(160));
    layer0_outputs(9911) <= not(inputs(199)) or (inputs(104));
    layer0_outputs(9912) <= inputs(54);
    layer0_outputs(9913) <= not(inputs(165)) or (inputs(204));
    layer0_outputs(9914) <= inputs(117);
    layer0_outputs(9915) <= not(inputs(220)) or (inputs(46));
    layer0_outputs(9916) <= not(inputs(39)) or (inputs(100));
    layer0_outputs(9917) <= not(inputs(157));
    layer0_outputs(9918) <= inputs(116);
    layer0_outputs(9919) <= (inputs(173)) and not (inputs(9));
    layer0_outputs(9920) <= (inputs(136)) xor (inputs(166));
    layer0_outputs(9921) <= inputs(87);
    layer0_outputs(9922) <= inputs(198);
    layer0_outputs(9923) <= inputs(56);
    layer0_outputs(9924) <= not(inputs(233));
    layer0_outputs(9925) <= (inputs(164)) and not (inputs(248));
    layer0_outputs(9926) <= not(inputs(164));
    layer0_outputs(9927) <= not((inputs(164)) xor (inputs(62)));
    layer0_outputs(9928) <= '1';
    layer0_outputs(9929) <= '1';
    layer0_outputs(9930) <= inputs(206);
    layer0_outputs(9931) <= not((inputs(8)) xor (inputs(91)));
    layer0_outputs(9932) <= not((inputs(21)) xor (inputs(139)));
    layer0_outputs(9933) <= (inputs(111)) or (inputs(151));
    layer0_outputs(9934) <= (inputs(139)) or (inputs(158));
    layer0_outputs(9935) <= (inputs(233)) and (inputs(51));
    layer0_outputs(9936) <= (inputs(188)) or (inputs(78));
    layer0_outputs(9937) <= (inputs(148)) or (inputs(33));
    layer0_outputs(9938) <= not(inputs(29));
    layer0_outputs(9939) <= not((inputs(209)) xor (inputs(1)));
    layer0_outputs(9940) <= not((inputs(220)) or (inputs(52)));
    layer0_outputs(9941) <= inputs(202);
    layer0_outputs(9942) <= not(inputs(218));
    layer0_outputs(9943) <= not(inputs(216));
    layer0_outputs(9944) <= not(inputs(106));
    layer0_outputs(9945) <= (inputs(164)) or (inputs(18));
    layer0_outputs(9946) <= inputs(229);
    layer0_outputs(9947) <= inputs(5);
    layer0_outputs(9948) <= not(inputs(72));
    layer0_outputs(9949) <= inputs(217);
    layer0_outputs(9950) <= not(inputs(126)) or (inputs(238));
    layer0_outputs(9951) <= not(inputs(153));
    layer0_outputs(9952) <= not((inputs(5)) and (inputs(14)));
    layer0_outputs(9953) <= inputs(59);
    layer0_outputs(9954) <= not((inputs(117)) or (inputs(158)));
    layer0_outputs(9955) <= not(inputs(205));
    layer0_outputs(9956) <= not((inputs(168)) or (inputs(245)));
    layer0_outputs(9957) <= (inputs(75)) and not (inputs(66));
    layer0_outputs(9958) <= inputs(149);
    layer0_outputs(9959) <= (inputs(27)) or (inputs(146));
    layer0_outputs(9960) <= not(inputs(239));
    layer0_outputs(9961) <= not((inputs(18)) xor (inputs(90)));
    layer0_outputs(9962) <= (inputs(164)) or (inputs(225));
    layer0_outputs(9963) <= not((inputs(35)) xor (inputs(199)));
    layer0_outputs(9964) <= (inputs(192)) xor (inputs(37));
    layer0_outputs(9965) <= inputs(73);
    layer0_outputs(9966) <= not((inputs(60)) xor (inputs(252)));
    layer0_outputs(9967) <= not(inputs(185));
    layer0_outputs(9968) <= inputs(99);
    layer0_outputs(9969) <= not(inputs(151));
    layer0_outputs(9970) <= not((inputs(57)) or (inputs(32)));
    layer0_outputs(9971) <= not((inputs(41)) xor (inputs(184)));
    layer0_outputs(9972) <= not((inputs(71)) or (inputs(178)));
    layer0_outputs(9973) <= not((inputs(224)) and (inputs(85)));
    layer0_outputs(9974) <= inputs(171);
    layer0_outputs(9975) <= (inputs(118)) and not (inputs(228));
    layer0_outputs(9976) <= (inputs(114)) and (inputs(48));
    layer0_outputs(9977) <= '0';
    layer0_outputs(9978) <= not(inputs(140)) or (inputs(67));
    layer0_outputs(9979) <= '0';
    layer0_outputs(9980) <= (inputs(200)) and not (inputs(52));
    layer0_outputs(9981) <= (inputs(166)) or (inputs(26));
    layer0_outputs(9982) <= (inputs(55)) and not (inputs(14));
    layer0_outputs(9983) <= inputs(93);
    layer0_outputs(9984) <= (inputs(86)) and not (inputs(177));
    layer0_outputs(9985) <= not((inputs(43)) or (inputs(141)));
    layer0_outputs(9986) <= (inputs(33)) xor (inputs(106));
    layer0_outputs(9987) <= not(inputs(118)) or (inputs(163));
    layer0_outputs(9988) <= not(inputs(253)) or (inputs(207));
    layer0_outputs(9989) <= (inputs(94)) and (inputs(82));
    layer0_outputs(9990) <= (inputs(211)) xor (inputs(109));
    layer0_outputs(9991) <= (inputs(47)) xor (inputs(105));
    layer0_outputs(9992) <= not((inputs(122)) xor (inputs(212)));
    layer0_outputs(9993) <= '0';
    layer0_outputs(9994) <= not(inputs(255));
    layer0_outputs(9995) <= not(inputs(61)) or (inputs(13));
    layer0_outputs(9996) <= not((inputs(180)) or (inputs(67)));
    layer0_outputs(9997) <= not((inputs(114)) xor (inputs(142)));
    layer0_outputs(9998) <= not((inputs(187)) xor (inputs(41)));
    layer0_outputs(9999) <= not((inputs(120)) or (inputs(129)));
    layer0_outputs(10000) <= not((inputs(84)) xor (inputs(58)));
    layer0_outputs(10001) <= not(inputs(170)) or (inputs(28));
    layer0_outputs(10002) <= inputs(61);
    layer0_outputs(10003) <= '1';
    layer0_outputs(10004) <= not(inputs(149));
    layer0_outputs(10005) <= not(inputs(106));
    layer0_outputs(10006) <= inputs(165);
    layer0_outputs(10007) <= not((inputs(97)) and (inputs(46)));
    layer0_outputs(10008) <= (inputs(155)) and (inputs(185));
    layer0_outputs(10009) <= (inputs(50)) and not (inputs(226));
    layer0_outputs(10010) <= not(inputs(80)) or (inputs(163));
    layer0_outputs(10011) <= not((inputs(151)) or (inputs(146)));
    layer0_outputs(10012) <= not(inputs(14)) or (inputs(168));
    layer0_outputs(10013) <= not((inputs(180)) or (inputs(153)));
    layer0_outputs(10014) <= inputs(120);
    layer0_outputs(10015) <= not((inputs(92)) xor (inputs(68)));
    layer0_outputs(10016) <= not((inputs(202)) xor (inputs(102)));
    layer0_outputs(10017) <= (inputs(245)) or (inputs(246));
    layer0_outputs(10018) <= not((inputs(107)) xor (inputs(97)));
    layer0_outputs(10019) <= inputs(36);
    layer0_outputs(10020) <= not(inputs(248)) or (inputs(211));
    layer0_outputs(10021) <= inputs(166);
    layer0_outputs(10022) <= not(inputs(206));
    layer0_outputs(10023) <= not((inputs(71)) xor (inputs(229)));
    layer0_outputs(10024) <= not((inputs(237)) or (inputs(18)));
    layer0_outputs(10025) <= not(inputs(146));
    layer0_outputs(10026) <= not(inputs(165)) or (inputs(224));
    layer0_outputs(10027) <= (inputs(5)) xor (inputs(215));
    layer0_outputs(10028) <= (inputs(115)) and not (inputs(5));
    layer0_outputs(10029) <= not(inputs(80));
    layer0_outputs(10030) <= (inputs(54)) or (inputs(140));
    layer0_outputs(10031) <= (inputs(133)) xor (inputs(164));
    layer0_outputs(10032) <= not(inputs(74));
    layer0_outputs(10033) <= (inputs(49)) or (inputs(217));
    layer0_outputs(10034) <= inputs(118);
    layer0_outputs(10035) <= inputs(124);
    layer0_outputs(10036) <= not((inputs(28)) or (inputs(183)));
    layer0_outputs(10037) <= not((inputs(225)) xor (inputs(150)));
    layer0_outputs(10038) <= not(inputs(105)) or (inputs(10));
    layer0_outputs(10039) <= (inputs(181)) and not (inputs(36));
    layer0_outputs(10040) <= not(inputs(113));
    layer0_outputs(10041) <= not(inputs(89)) or (inputs(83));
    layer0_outputs(10042) <= (inputs(78)) or (inputs(92));
    layer0_outputs(10043) <= not(inputs(117));
    layer0_outputs(10044) <= inputs(32);
    layer0_outputs(10045) <= not((inputs(21)) xor (inputs(160)));
    layer0_outputs(10046) <= not(inputs(23));
    layer0_outputs(10047) <= not((inputs(85)) or (inputs(4)));
    layer0_outputs(10048) <= not((inputs(254)) or (inputs(188)));
    layer0_outputs(10049) <= not((inputs(150)) or (inputs(220)));
    layer0_outputs(10050) <= not((inputs(78)) xor (inputs(62)));
    layer0_outputs(10051) <= inputs(195);
    layer0_outputs(10052) <= not(inputs(45));
    layer0_outputs(10053) <= not(inputs(158));
    layer0_outputs(10054) <= not((inputs(212)) xor (inputs(41)));
    layer0_outputs(10055) <= (inputs(115)) or (inputs(249));
    layer0_outputs(10056) <= (inputs(11)) and not (inputs(9));
    layer0_outputs(10057) <= (inputs(88)) xor (inputs(30));
    layer0_outputs(10058) <= (inputs(91)) and not (inputs(9));
    layer0_outputs(10059) <= inputs(104);
    layer0_outputs(10060) <= (inputs(103)) and not (inputs(160));
    layer0_outputs(10061) <= (inputs(71)) xor (inputs(55));
    layer0_outputs(10062) <= not((inputs(209)) xor (inputs(150)));
    layer0_outputs(10063) <= (inputs(85)) or (inputs(122));
    layer0_outputs(10064) <= (inputs(237)) xor (inputs(163));
    layer0_outputs(10065) <= (inputs(175)) xor (inputs(142));
    layer0_outputs(10066) <= not((inputs(101)) or (inputs(205)));
    layer0_outputs(10067) <= (inputs(70)) xor (inputs(122));
    layer0_outputs(10068) <= not((inputs(89)) xor (inputs(115)));
    layer0_outputs(10069) <= not((inputs(249)) and (inputs(74)));
    layer0_outputs(10070) <= not(inputs(33));
    layer0_outputs(10071) <= (inputs(51)) and not (inputs(241));
    layer0_outputs(10072) <= not(inputs(40)) or (inputs(232));
    layer0_outputs(10073) <= not(inputs(232));
    layer0_outputs(10074) <= not(inputs(180)) or (inputs(8));
    layer0_outputs(10075) <= (inputs(72)) and not (inputs(66));
    layer0_outputs(10076) <= inputs(5);
    layer0_outputs(10077) <= inputs(80);
    layer0_outputs(10078) <= not((inputs(106)) xor (inputs(226)));
    layer0_outputs(10079) <= not((inputs(97)) xor (inputs(243)));
    layer0_outputs(10080) <= not((inputs(26)) or (inputs(209)));
    layer0_outputs(10081) <= (inputs(20)) and not (inputs(191));
    layer0_outputs(10082) <= not((inputs(68)) or (inputs(170)));
    layer0_outputs(10083) <= inputs(88);
    layer0_outputs(10084) <= not(inputs(72)) or (inputs(98));
    layer0_outputs(10085) <= not((inputs(56)) xor (inputs(171)));
    layer0_outputs(10086) <= not(inputs(103));
    layer0_outputs(10087) <= not((inputs(204)) or (inputs(148)));
    layer0_outputs(10088) <= not(inputs(103));
    layer0_outputs(10089) <= not((inputs(22)) or (inputs(138)));
    layer0_outputs(10090) <= (inputs(38)) and not (inputs(128));
    layer0_outputs(10091) <= not(inputs(22));
    layer0_outputs(10092) <= not(inputs(22));
    layer0_outputs(10093) <= inputs(120);
    layer0_outputs(10094) <= not(inputs(229));
    layer0_outputs(10095) <= '0';
    layer0_outputs(10096) <= not(inputs(157)) or (inputs(83));
    layer0_outputs(10097) <= inputs(124);
    layer0_outputs(10098) <= (inputs(2)) xor (inputs(168));
    layer0_outputs(10099) <= (inputs(134)) or (inputs(173));
    layer0_outputs(10100) <= not((inputs(111)) or (inputs(85)));
    layer0_outputs(10101) <= not(inputs(207)) or (inputs(32));
    layer0_outputs(10102) <= (inputs(26)) xor (inputs(80));
    layer0_outputs(10103) <= (inputs(19)) xor (inputs(97));
    layer0_outputs(10104) <= not((inputs(130)) xor (inputs(3)));
    layer0_outputs(10105) <= inputs(19);
    layer0_outputs(10106) <= not(inputs(66));
    layer0_outputs(10107) <= not((inputs(194)) xor (inputs(163)));
    layer0_outputs(10108) <= not(inputs(125)) or (inputs(97));
    layer0_outputs(10109) <= not((inputs(164)) xor (inputs(169)));
    layer0_outputs(10110) <= (inputs(92)) or (inputs(65));
    layer0_outputs(10111) <= not(inputs(103)) or (inputs(145));
    layer0_outputs(10112) <= not(inputs(233)) or (inputs(255));
    layer0_outputs(10113) <= (inputs(234)) or (inputs(100));
    layer0_outputs(10114) <= (inputs(70)) and not (inputs(58));
    layer0_outputs(10115) <= (inputs(253)) or (inputs(213));
    layer0_outputs(10116) <= not((inputs(24)) xor (inputs(235)));
    layer0_outputs(10117) <= (inputs(203)) and not (inputs(14));
    layer0_outputs(10118) <= (inputs(152)) and not (inputs(247));
    layer0_outputs(10119) <= not(inputs(130));
    layer0_outputs(10120) <= (inputs(134)) and not (inputs(174));
    layer0_outputs(10121) <= inputs(122);
    layer0_outputs(10122) <= (inputs(183)) and not (inputs(176));
    layer0_outputs(10123) <= not((inputs(11)) xor (inputs(96)));
    layer0_outputs(10124) <= (inputs(148)) or (inputs(39));
    layer0_outputs(10125) <= not((inputs(94)) xor (inputs(74)));
    layer0_outputs(10126) <= not((inputs(56)) xor (inputs(199)));
    layer0_outputs(10127) <= inputs(136);
    layer0_outputs(10128) <= not(inputs(92));
    layer0_outputs(10129) <= not((inputs(2)) or (inputs(253)));
    layer0_outputs(10130) <= inputs(122);
    layer0_outputs(10131) <= not((inputs(112)) or (inputs(152)));
    layer0_outputs(10132) <= '0';
    layer0_outputs(10133) <= not((inputs(111)) or (inputs(87)));
    layer0_outputs(10134) <= not((inputs(63)) and (inputs(158)));
    layer0_outputs(10135) <= (inputs(154)) or (inputs(195));
    layer0_outputs(10136) <= (inputs(172)) or (inputs(83));
    layer0_outputs(10137) <= not((inputs(180)) xor (inputs(253)));
    layer0_outputs(10138) <= (inputs(109)) and not (inputs(11));
    layer0_outputs(10139) <= not((inputs(185)) and (inputs(177)));
    layer0_outputs(10140) <= '0';
    layer0_outputs(10141) <= (inputs(23)) and not (inputs(196));
    layer0_outputs(10142) <= (inputs(186)) and not (inputs(233));
    layer0_outputs(10143) <= (inputs(58)) and not (inputs(24));
    layer0_outputs(10144) <= not((inputs(116)) or (inputs(155)));
    layer0_outputs(10145) <= not(inputs(82));
    layer0_outputs(10146) <= (inputs(97)) xor (inputs(204));
    layer0_outputs(10147) <= not(inputs(61));
    layer0_outputs(10148) <= inputs(168);
    layer0_outputs(10149) <= (inputs(144)) and not (inputs(218));
    layer0_outputs(10150) <= not(inputs(139));
    layer0_outputs(10151) <= not((inputs(164)) or (inputs(142)));
    layer0_outputs(10152) <= inputs(188);
    layer0_outputs(10153) <= (inputs(148)) and not (inputs(202));
    layer0_outputs(10154) <= (inputs(223)) or (inputs(97));
    layer0_outputs(10155) <= (inputs(103)) and (inputs(227));
    layer0_outputs(10156) <= not((inputs(195)) and (inputs(75)));
    layer0_outputs(10157) <= not(inputs(159)) or (inputs(48));
    layer0_outputs(10158) <= not(inputs(88));
    layer0_outputs(10159) <= not(inputs(225));
    layer0_outputs(10160) <= not(inputs(165)) or (inputs(141));
    layer0_outputs(10161) <= (inputs(113)) xor (inputs(84));
    layer0_outputs(10162) <= (inputs(83)) or (inputs(64));
    layer0_outputs(10163) <= not((inputs(252)) or (inputs(72)));
    layer0_outputs(10164) <= not((inputs(126)) xor (inputs(41)));
    layer0_outputs(10165) <= (inputs(191)) xor (inputs(246));
    layer0_outputs(10166) <= '0';
    layer0_outputs(10167) <= (inputs(182)) or (inputs(128));
    layer0_outputs(10168) <= (inputs(109)) xor (inputs(159));
    layer0_outputs(10169) <= not((inputs(251)) or (inputs(195)));
    layer0_outputs(10170) <= not(inputs(4)) or (inputs(164));
    layer0_outputs(10171) <= (inputs(37)) or (inputs(17));
    layer0_outputs(10172) <= not(inputs(163));
    layer0_outputs(10173) <= not(inputs(108));
    layer0_outputs(10174) <= (inputs(216)) and not (inputs(114));
    layer0_outputs(10175) <= not(inputs(28)) or (inputs(197));
    layer0_outputs(10176) <= not(inputs(38));
    layer0_outputs(10177) <= (inputs(235)) or (inputs(130));
    layer0_outputs(10178) <= not(inputs(55));
    layer0_outputs(10179) <= not((inputs(163)) xor (inputs(253)));
    layer0_outputs(10180) <= not((inputs(248)) xor (inputs(235)));
    layer0_outputs(10181) <= (inputs(143)) and not (inputs(127));
    layer0_outputs(10182) <= (inputs(137)) and not (inputs(251));
    layer0_outputs(10183) <= not(inputs(193)) or (inputs(207));
    layer0_outputs(10184) <= inputs(248);
    layer0_outputs(10185) <= (inputs(251)) xor (inputs(72));
    layer0_outputs(10186) <= (inputs(221)) or (inputs(77));
    layer0_outputs(10187) <= '1';
    layer0_outputs(10188) <= inputs(187);
    layer0_outputs(10189) <= (inputs(196)) and (inputs(186));
    layer0_outputs(10190) <= not((inputs(43)) and (inputs(45)));
    layer0_outputs(10191) <= not((inputs(131)) or (inputs(176)));
    layer0_outputs(10192) <= not(inputs(225)) or (inputs(110));
    layer0_outputs(10193) <= not((inputs(179)) or (inputs(27)));
    layer0_outputs(10194) <= (inputs(116)) and not (inputs(4));
    layer0_outputs(10195) <= not((inputs(124)) or (inputs(24)));
    layer0_outputs(10196) <= (inputs(162)) xor (inputs(90));
    layer0_outputs(10197) <= not((inputs(38)) or (inputs(174)));
    layer0_outputs(10198) <= not((inputs(90)) or (inputs(142)));
    layer0_outputs(10199) <= (inputs(132)) and not (inputs(231));
    layer0_outputs(10200) <= (inputs(123)) or (inputs(238));
    layer0_outputs(10201) <= not((inputs(227)) or (inputs(106)));
    layer0_outputs(10202) <= inputs(61);
    layer0_outputs(10203) <= not((inputs(139)) or (inputs(165)));
    layer0_outputs(10204) <= not((inputs(85)) or (inputs(237)));
    layer0_outputs(10205) <= (inputs(96)) or (inputs(233));
    layer0_outputs(10206) <= (inputs(26)) and not (inputs(76));
    layer0_outputs(10207) <= not((inputs(128)) or (inputs(140)));
    layer0_outputs(10208) <= not(inputs(87));
    layer0_outputs(10209) <= (inputs(149)) or (inputs(216));
    layer0_outputs(10210) <= inputs(75);
    layer0_outputs(10211) <= not((inputs(9)) xor (inputs(231)));
    layer0_outputs(10212) <= not((inputs(148)) or (inputs(236)));
    layer0_outputs(10213) <= not((inputs(42)) xor (inputs(123)));
    layer0_outputs(10214) <= not(inputs(199));
    layer0_outputs(10215) <= (inputs(74)) and not (inputs(195));
    layer0_outputs(10216) <= not(inputs(135)) or (inputs(46));
    layer0_outputs(10217) <= not(inputs(14));
    layer0_outputs(10218) <= '1';
    layer0_outputs(10219) <= inputs(26);
    layer0_outputs(10220) <= not(inputs(242));
    layer0_outputs(10221) <= (inputs(81)) and not (inputs(126));
    layer0_outputs(10222) <= (inputs(68)) and not (inputs(125));
    layer0_outputs(10223) <= not(inputs(147));
    layer0_outputs(10224) <= inputs(73);
    layer0_outputs(10225) <= (inputs(105)) xor (inputs(169));
    layer0_outputs(10226) <= (inputs(227)) or (inputs(102));
    layer0_outputs(10227) <= '1';
    layer0_outputs(10228) <= (inputs(171)) and not (inputs(240));
    layer0_outputs(10229) <= inputs(222);
    layer0_outputs(10230) <= (inputs(194)) xor (inputs(203));
    layer0_outputs(10231) <= (inputs(216)) or (inputs(49));
    layer0_outputs(10232) <= '0';
    layer0_outputs(10233) <= (inputs(52)) and not (inputs(191));
    layer0_outputs(10234) <= not((inputs(213)) or (inputs(16)));
    layer0_outputs(10235) <= (inputs(53)) or (inputs(134));
    layer0_outputs(10236) <= '1';
    layer0_outputs(10237) <= not((inputs(81)) or (inputs(171)));
    layer0_outputs(10238) <= not(inputs(206));
    layer0_outputs(10239) <= not(inputs(151)) or (inputs(130));
    layer0_outputs(10240) <= (inputs(32)) and (inputs(87));
    layer0_outputs(10241) <= (inputs(192)) xor (inputs(96));
    layer0_outputs(10242) <= '1';
    layer0_outputs(10243) <= (inputs(196)) or (inputs(213));
    layer0_outputs(10244) <= (inputs(43)) or (inputs(140));
    layer0_outputs(10245) <= (inputs(206)) xor (inputs(135));
    layer0_outputs(10246) <= (inputs(110)) and not (inputs(51));
    layer0_outputs(10247) <= (inputs(247)) xor (inputs(10));
    layer0_outputs(10248) <= (inputs(188)) and not (inputs(132));
    layer0_outputs(10249) <= not(inputs(161)) or (inputs(45));
    layer0_outputs(10250) <= not(inputs(137));
    layer0_outputs(10251) <= (inputs(88)) and not (inputs(179));
    layer0_outputs(10252) <= not(inputs(214));
    layer0_outputs(10253) <= (inputs(104)) and not (inputs(141));
    layer0_outputs(10254) <= inputs(40);
    layer0_outputs(10255) <= not((inputs(138)) or (inputs(227)));
    layer0_outputs(10256) <= not(inputs(214));
    layer0_outputs(10257) <= (inputs(255)) or (inputs(14));
    layer0_outputs(10258) <= (inputs(212)) and not (inputs(47));
    layer0_outputs(10259) <= not(inputs(252)) or (inputs(58));
    layer0_outputs(10260) <= (inputs(80)) or (inputs(136));
    layer0_outputs(10261) <= (inputs(251)) and (inputs(148));
    layer0_outputs(10262) <= not(inputs(42)) or (inputs(250));
    layer0_outputs(10263) <= inputs(231);
    layer0_outputs(10264) <= not(inputs(173)) or (inputs(245));
    layer0_outputs(10265) <= inputs(251);
    layer0_outputs(10266) <= (inputs(231)) or (inputs(248));
    layer0_outputs(10267) <= not((inputs(57)) xor (inputs(137)));
    layer0_outputs(10268) <= inputs(149);
    layer0_outputs(10269) <= '1';
    layer0_outputs(10270) <= not((inputs(163)) xor (inputs(65)));
    layer0_outputs(10271) <= not((inputs(75)) xor (inputs(205)));
    layer0_outputs(10272) <= (inputs(36)) xor (inputs(217));
    layer0_outputs(10273) <= not(inputs(90));
    layer0_outputs(10274) <= (inputs(28)) xor (inputs(232));
    layer0_outputs(10275) <= not(inputs(148)) or (inputs(78));
    layer0_outputs(10276) <= not((inputs(150)) or (inputs(172)));
    layer0_outputs(10277) <= not((inputs(53)) or (inputs(162)));
    layer0_outputs(10278) <= inputs(17);
    layer0_outputs(10279) <= inputs(240);
    layer0_outputs(10280) <= not((inputs(78)) or (inputs(29)));
    layer0_outputs(10281) <= inputs(178);
    layer0_outputs(10282) <= not((inputs(70)) xor (inputs(164)));
    layer0_outputs(10283) <= (inputs(46)) xor (inputs(80));
    layer0_outputs(10284) <= '0';
    layer0_outputs(10285) <= inputs(131);
    layer0_outputs(10286) <= (inputs(215)) xor (inputs(134));
    layer0_outputs(10287) <= inputs(214);
    layer0_outputs(10288) <= not(inputs(37)) or (inputs(235));
    layer0_outputs(10289) <= not((inputs(251)) or (inputs(52)));
    layer0_outputs(10290) <= inputs(147);
    layer0_outputs(10291) <= '1';
    layer0_outputs(10292) <= not((inputs(26)) or (inputs(140)));
    layer0_outputs(10293) <= not(inputs(179));
    layer0_outputs(10294) <= inputs(116);
    layer0_outputs(10295) <= (inputs(95)) xor (inputs(178));
    layer0_outputs(10296) <= not(inputs(71)) or (inputs(16));
    layer0_outputs(10297) <= not(inputs(106)) or (inputs(87));
    layer0_outputs(10298) <= (inputs(235)) xor (inputs(233));
    layer0_outputs(10299) <= (inputs(169)) xor (inputs(185));
    layer0_outputs(10300) <= not(inputs(0));
    layer0_outputs(10301) <= not(inputs(240)) or (inputs(144));
    layer0_outputs(10302) <= not(inputs(214));
    layer0_outputs(10303) <= not(inputs(90)) or (inputs(47));
    layer0_outputs(10304) <= inputs(244);
    layer0_outputs(10305) <= not((inputs(71)) xor (inputs(7)));
    layer0_outputs(10306) <= not((inputs(12)) or (inputs(242)));
    layer0_outputs(10307) <= (inputs(2)) or (inputs(35));
    layer0_outputs(10308) <= '0';
    layer0_outputs(10309) <= (inputs(234)) xor (inputs(241));
    layer0_outputs(10310) <= not(inputs(190)) or (inputs(91));
    layer0_outputs(10311) <= not(inputs(115));
    layer0_outputs(10312) <= not(inputs(59)) or (inputs(1));
    layer0_outputs(10313) <= not((inputs(46)) or (inputs(180)));
    layer0_outputs(10314) <= (inputs(233)) or (inputs(224));
    layer0_outputs(10315) <= inputs(41);
    layer0_outputs(10316) <= not(inputs(90)) or (inputs(45));
    layer0_outputs(10317) <= not(inputs(122)) or (inputs(218));
    layer0_outputs(10318) <= not((inputs(38)) or (inputs(123)));
    layer0_outputs(10319) <= (inputs(132)) and not (inputs(127));
    layer0_outputs(10320) <= '1';
    layer0_outputs(10321) <= inputs(44);
    layer0_outputs(10322) <= not(inputs(74)) or (inputs(149));
    layer0_outputs(10323) <= not((inputs(207)) and (inputs(193)));
    layer0_outputs(10324) <= not((inputs(215)) and (inputs(116)));
    layer0_outputs(10325) <= (inputs(195)) and not (inputs(20));
    layer0_outputs(10326) <= (inputs(194)) and not (inputs(62));
    layer0_outputs(10327) <= not((inputs(199)) xor (inputs(0)));
    layer0_outputs(10328) <= (inputs(50)) and not (inputs(244));
    layer0_outputs(10329) <= (inputs(53)) or (inputs(153));
    layer0_outputs(10330) <= (inputs(7)) xor (inputs(192));
    layer0_outputs(10331) <= not((inputs(234)) xor (inputs(203)));
    layer0_outputs(10332) <= inputs(64);
    layer0_outputs(10333) <= (inputs(40)) xor (inputs(236));
    layer0_outputs(10334) <= not(inputs(230));
    layer0_outputs(10335) <= (inputs(182)) or (inputs(252));
    layer0_outputs(10336) <= inputs(196);
    layer0_outputs(10337) <= (inputs(139)) or (inputs(110));
    layer0_outputs(10338) <= (inputs(153)) and not (inputs(78));
    layer0_outputs(10339) <= not((inputs(185)) xor (inputs(97)));
    layer0_outputs(10340) <= not(inputs(190));
    layer0_outputs(10341) <= not(inputs(136));
    layer0_outputs(10342) <= not((inputs(11)) and (inputs(124)));
    layer0_outputs(10343) <= not((inputs(36)) or (inputs(201)));
    layer0_outputs(10344) <= (inputs(55)) or (inputs(3));
    layer0_outputs(10345) <= (inputs(178)) and not (inputs(208));
    layer0_outputs(10346) <= not((inputs(246)) and (inputs(247)));
    layer0_outputs(10347) <= not(inputs(97)) or (inputs(126));
    layer0_outputs(10348) <= (inputs(103)) or (inputs(156));
    layer0_outputs(10349) <= not(inputs(252)) or (inputs(159));
    layer0_outputs(10350) <= not((inputs(177)) or (inputs(29)));
    layer0_outputs(10351) <= not(inputs(216)) or (inputs(44));
    layer0_outputs(10352) <= (inputs(139)) and not (inputs(249));
    layer0_outputs(10353) <= not((inputs(70)) and (inputs(229)));
    layer0_outputs(10354) <= not(inputs(102)) or (inputs(34));
    layer0_outputs(10355) <= (inputs(9)) xor (inputs(243));
    layer0_outputs(10356) <= not((inputs(148)) and (inputs(9)));
    layer0_outputs(10357) <= not((inputs(58)) xor (inputs(115)));
    layer0_outputs(10358) <= inputs(102);
    layer0_outputs(10359) <= not((inputs(63)) or (inputs(100)));
    layer0_outputs(10360) <= not(inputs(86));
    layer0_outputs(10361) <= '0';
    layer0_outputs(10362) <= inputs(186);
    layer0_outputs(10363) <= (inputs(58)) xor (inputs(93));
    layer0_outputs(10364) <= inputs(80);
    layer0_outputs(10365) <= not(inputs(40));
    layer0_outputs(10366) <= (inputs(143)) or (inputs(229));
    layer0_outputs(10367) <= not(inputs(198));
    layer0_outputs(10368) <= (inputs(191)) xor (inputs(154));
    layer0_outputs(10369) <= not((inputs(71)) xor (inputs(92)));
    layer0_outputs(10370) <= (inputs(80)) xor (inputs(150));
    layer0_outputs(10371) <= not(inputs(156)) or (inputs(16));
    layer0_outputs(10372) <= not((inputs(166)) or (inputs(204)));
    layer0_outputs(10373) <= not(inputs(88)) or (inputs(164));
    layer0_outputs(10374) <= inputs(168);
    layer0_outputs(10375) <= not((inputs(56)) xor (inputs(43)));
    layer0_outputs(10376) <= (inputs(150)) or (inputs(218));
    layer0_outputs(10377) <= not((inputs(96)) xor (inputs(249)));
    layer0_outputs(10378) <= inputs(108);
    layer0_outputs(10379) <= '1';
    layer0_outputs(10380) <= not((inputs(181)) xor (inputs(204)));
    layer0_outputs(10381) <= not(inputs(241)) or (inputs(218));
    layer0_outputs(10382) <= (inputs(105)) and not (inputs(243));
    layer0_outputs(10383) <= inputs(117);
    layer0_outputs(10384) <= not(inputs(253));
    layer0_outputs(10385) <= (inputs(113)) and not (inputs(62));
    layer0_outputs(10386) <= inputs(116);
    layer0_outputs(10387) <= not((inputs(89)) or (inputs(63)));
    layer0_outputs(10388) <= (inputs(47)) and not (inputs(47));
    layer0_outputs(10389) <= (inputs(203)) xor (inputs(151));
    layer0_outputs(10390) <= (inputs(117)) xor (inputs(116));
    layer0_outputs(10391) <= not((inputs(51)) and (inputs(247)));
    layer0_outputs(10392) <= not((inputs(205)) or (inputs(164)));
    layer0_outputs(10393) <= not(inputs(51));
    layer0_outputs(10394) <= (inputs(104)) and not (inputs(15));
    layer0_outputs(10395) <= (inputs(234)) or (inputs(154));
    layer0_outputs(10396) <= (inputs(137)) xor (inputs(67));
    layer0_outputs(10397) <= not((inputs(88)) or (inputs(33)));
    layer0_outputs(10398) <= not(inputs(149));
    layer0_outputs(10399) <= '1';
    layer0_outputs(10400) <= (inputs(150)) or (inputs(167));
    layer0_outputs(10401) <= not((inputs(67)) xor (inputs(154)));
    layer0_outputs(10402) <= not(inputs(235)) or (inputs(253));
    layer0_outputs(10403) <= not(inputs(196));
    layer0_outputs(10404) <= (inputs(52)) and not (inputs(8));
    layer0_outputs(10405) <= not(inputs(199));
    layer0_outputs(10406) <= not(inputs(159)) or (inputs(224));
    layer0_outputs(10407) <= not((inputs(67)) xor (inputs(124)));
    layer0_outputs(10408) <= not(inputs(33)) or (inputs(224));
    layer0_outputs(10409) <= (inputs(195)) xor (inputs(85));
    layer0_outputs(10410) <= (inputs(137)) and not (inputs(180));
    layer0_outputs(10411) <= not((inputs(23)) xor (inputs(70)));
    layer0_outputs(10412) <= not(inputs(108));
    layer0_outputs(10413) <= not((inputs(211)) or (inputs(211)));
    layer0_outputs(10414) <= not(inputs(218));
    layer0_outputs(10415) <= (inputs(222)) and not (inputs(16));
    layer0_outputs(10416) <= (inputs(194)) and (inputs(206));
    layer0_outputs(10417) <= (inputs(195)) xor (inputs(59));
    layer0_outputs(10418) <= (inputs(191)) xor (inputs(252));
    layer0_outputs(10419) <= (inputs(227)) and not (inputs(209));
    layer0_outputs(10420) <= not(inputs(60));
    layer0_outputs(10421) <= not(inputs(44)) or (inputs(8));
    layer0_outputs(10422) <= not(inputs(222)) or (inputs(54));
    layer0_outputs(10423) <= not(inputs(108)) or (inputs(31));
    layer0_outputs(10424) <= (inputs(202)) or (inputs(54));
    layer0_outputs(10425) <= inputs(156);
    layer0_outputs(10426) <= (inputs(229)) xor (inputs(125));
    layer0_outputs(10427) <= not(inputs(206)) or (inputs(39));
    layer0_outputs(10428) <= not(inputs(102));
    layer0_outputs(10429) <= not(inputs(178));
    layer0_outputs(10430) <= (inputs(37)) or (inputs(98));
    layer0_outputs(10431) <= (inputs(2)) or (inputs(160));
    layer0_outputs(10432) <= not((inputs(253)) xor (inputs(189)));
    layer0_outputs(10433) <= (inputs(234)) or (inputs(107));
    layer0_outputs(10434) <= (inputs(179)) xor (inputs(212));
    layer0_outputs(10435) <= (inputs(10)) and (inputs(4));
    layer0_outputs(10436) <= not((inputs(17)) or (inputs(95)));
    layer0_outputs(10437) <= not((inputs(0)) and (inputs(16)));
    layer0_outputs(10438) <= not((inputs(113)) xor (inputs(53)));
    layer0_outputs(10439) <= not(inputs(117));
    layer0_outputs(10440) <= (inputs(25)) and not (inputs(157));
    layer0_outputs(10441) <= not(inputs(155)) or (inputs(16));
    layer0_outputs(10442) <= (inputs(58)) and not (inputs(174));
    layer0_outputs(10443) <= not(inputs(183));
    layer0_outputs(10444) <= (inputs(155)) or (inputs(54));
    layer0_outputs(10445) <= (inputs(170)) and not (inputs(42));
    layer0_outputs(10446) <= (inputs(14)) and (inputs(46));
    layer0_outputs(10447) <= '1';
    layer0_outputs(10448) <= (inputs(250)) or (inputs(119));
    layer0_outputs(10449) <= (inputs(74)) and not (inputs(103));
    layer0_outputs(10450) <= (inputs(182)) xor (inputs(120));
    layer0_outputs(10451) <= (inputs(129)) xor (inputs(29));
    layer0_outputs(10452) <= not((inputs(157)) or (inputs(13)));
    layer0_outputs(10453) <= not((inputs(92)) and (inputs(191)));
    layer0_outputs(10454) <= not((inputs(235)) xor (inputs(249)));
    layer0_outputs(10455) <= (inputs(193)) xor (inputs(233));
    layer0_outputs(10456) <= not(inputs(117));
    layer0_outputs(10457) <= not(inputs(165)) or (inputs(223));
    layer0_outputs(10458) <= not((inputs(213)) or (inputs(179)));
    layer0_outputs(10459) <= (inputs(0)) or (inputs(45));
    layer0_outputs(10460) <= (inputs(42)) xor (inputs(202));
    layer0_outputs(10461) <= not(inputs(15));
    layer0_outputs(10462) <= (inputs(146)) xor (inputs(229));
    layer0_outputs(10463) <= (inputs(221)) and not (inputs(19));
    layer0_outputs(10464) <= not(inputs(39)) or (inputs(28));
    layer0_outputs(10465) <= (inputs(139)) xor (inputs(226));
    layer0_outputs(10466) <= not((inputs(236)) or (inputs(105)));
    layer0_outputs(10467) <= (inputs(12)) or (inputs(31));
    layer0_outputs(10468) <= not(inputs(15)) or (inputs(103));
    layer0_outputs(10469) <= (inputs(140)) xor (inputs(175));
    layer0_outputs(10470) <= (inputs(171)) or (inputs(39));
    layer0_outputs(10471) <= (inputs(72)) or (inputs(16));
    layer0_outputs(10472) <= not(inputs(245));
    layer0_outputs(10473) <= not((inputs(35)) and (inputs(206)));
    layer0_outputs(10474) <= inputs(147);
    layer0_outputs(10475) <= (inputs(74)) and not (inputs(221));
    layer0_outputs(10476) <= not((inputs(254)) xor (inputs(202)));
    layer0_outputs(10477) <= (inputs(141)) and not (inputs(159));
    layer0_outputs(10478) <= (inputs(75)) or (inputs(171));
    layer0_outputs(10479) <= '1';
    layer0_outputs(10480) <= (inputs(213)) or (inputs(61));
    layer0_outputs(10481) <= not((inputs(85)) or (inputs(241)));
    layer0_outputs(10482) <= (inputs(210)) and not (inputs(23));
    layer0_outputs(10483) <= not(inputs(151));
    layer0_outputs(10484) <= (inputs(69)) xor (inputs(187));
    layer0_outputs(10485) <= (inputs(232)) and not (inputs(60));
    layer0_outputs(10486) <= (inputs(200)) and not (inputs(190));
    layer0_outputs(10487) <= not(inputs(221));
    layer0_outputs(10488) <= not((inputs(179)) or (inputs(170)));
    layer0_outputs(10489) <= not((inputs(154)) or (inputs(164)));
    layer0_outputs(10490) <= (inputs(137)) xor (inputs(223));
    layer0_outputs(10491) <= (inputs(125)) and not (inputs(210));
    layer0_outputs(10492) <= (inputs(143)) and (inputs(251));
    layer0_outputs(10493) <= (inputs(250)) xor (inputs(247));
    layer0_outputs(10494) <= (inputs(193)) or (inputs(63));
    layer0_outputs(10495) <= not((inputs(229)) or (inputs(97)));
    layer0_outputs(10496) <= (inputs(142)) xor (inputs(93));
    layer0_outputs(10497) <= not(inputs(67)) or (inputs(65));
    layer0_outputs(10498) <= not(inputs(123));
    layer0_outputs(10499) <= not((inputs(169)) or (inputs(16)));
    layer0_outputs(10500) <= not((inputs(226)) or (inputs(161)));
    layer0_outputs(10501) <= not((inputs(97)) or (inputs(225)));
    layer0_outputs(10502) <= not(inputs(152)) or (inputs(240));
    layer0_outputs(10503) <= (inputs(208)) and not (inputs(160));
    layer0_outputs(10504) <= (inputs(35)) and (inputs(12));
    layer0_outputs(10505) <= (inputs(49)) or (inputs(102));
    layer0_outputs(10506) <= not((inputs(129)) or (inputs(231)));
    layer0_outputs(10507) <= not((inputs(15)) or (inputs(182)));
    layer0_outputs(10508) <= inputs(232);
    layer0_outputs(10509) <= not((inputs(116)) or (inputs(234)));
    layer0_outputs(10510) <= (inputs(217)) and not (inputs(207));
    layer0_outputs(10511) <= (inputs(96)) xor (inputs(167));
    layer0_outputs(10512) <= not((inputs(67)) xor (inputs(91)));
    layer0_outputs(10513) <= (inputs(70)) or (inputs(24));
    layer0_outputs(10514) <= '1';
    layer0_outputs(10515) <= inputs(115);
    layer0_outputs(10516) <= not(inputs(246));
    layer0_outputs(10517) <= '1';
    layer0_outputs(10518) <= not(inputs(153)) or (inputs(120));
    layer0_outputs(10519) <= (inputs(71)) xor (inputs(83));
    layer0_outputs(10520) <= (inputs(38)) and not (inputs(41));
    layer0_outputs(10521) <= not((inputs(61)) or (inputs(134)));
    layer0_outputs(10522) <= not(inputs(50));
    layer0_outputs(10523) <= not((inputs(68)) or (inputs(25)));
    layer0_outputs(10524) <= not(inputs(119)) or (inputs(94));
    layer0_outputs(10525) <= (inputs(245)) xor (inputs(156));
    layer0_outputs(10526) <= (inputs(42)) or (inputs(65));
    layer0_outputs(10527) <= (inputs(87)) xor (inputs(113));
    layer0_outputs(10528) <= (inputs(48)) and not (inputs(165));
    layer0_outputs(10529) <= not((inputs(41)) or (inputs(205)));
    layer0_outputs(10530) <= (inputs(183)) xor (inputs(135));
    layer0_outputs(10531) <= inputs(154);
    layer0_outputs(10532) <= not(inputs(43));
    layer0_outputs(10533) <= inputs(246);
    layer0_outputs(10534) <= not(inputs(100));
    layer0_outputs(10535) <= (inputs(104)) and not (inputs(166));
    layer0_outputs(10536) <= inputs(182);
    layer0_outputs(10537) <= not((inputs(30)) xor (inputs(19)));
    layer0_outputs(10538) <= not((inputs(4)) xor (inputs(140)));
    layer0_outputs(10539) <= (inputs(58)) and not (inputs(67));
    layer0_outputs(10540) <= '0';
    layer0_outputs(10541) <= not(inputs(160)) or (inputs(251));
    layer0_outputs(10542) <= inputs(231);
    layer0_outputs(10543) <= not(inputs(96)) or (inputs(168));
    layer0_outputs(10544) <= (inputs(188)) xor (inputs(48));
    layer0_outputs(10545) <= (inputs(203)) xor (inputs(141));
    layer0_outputs(10546) <= not(inputs(117));
    layer0_outputs(10547) <= '0';
    layer0_outputs(10548) <= (inputs(151)) and not (inputs(5));
    layer0_outputs(10549) <= inputs(132);
    layer0_outputs(10550) <= (inputs(166)) or (inputs(5));
    layer0_outputs(10551) <= (inputs(178)) and not (inputs(235));
    layer0_outputs(10552) <= not(inputs(88));
    layer0_outputs(10553) <= not((inputs(181)) xor (inputs(36)));
    layer0_outputs(10554) <= not((inputs(95)) xor (inputs(216)));
    layer0_outputs(10555) <= not(inputs(33));
    layer0_outputs(10556) <= inputs(246);
    layer0_outputs(10557) <= inputs(105);
    layer0_outputs(10558) <= (inputs(218)) and not (inputs(27));
    layer0_outputs(10559) <= not((inputs(213)) or (inputs(203)));
    layer0_outputs(10560) <= (inputs(221)) or (inputs(31));
    layer0_outputs(10561) <= (inputs(135)) or (inputs(40));
    layer0_outputs(10562) <= not(inputs(68)) or (inputs(146));
    layer0_outputs(10563) <= not((inputs(22)) or (inputs(198)));
    layer0_outputs(10564) <= not(inputs(115)) or (inputs(113));
    layer0_outputs(10565) <= (inputs(181)) and not (inputs(37));
    layer0_outputs(10566) <= not(inputs(84)) or (inputs(71));
    layer0_outputs(10567) <= inputs(65);
    layer0_outputs(10568) <= not((inputs(146)) xor (inputs(70)));
    layer0_outputs(10569) <= not((inputs(253)) xor (inputs(122)));
    layer0_outputs(10570) <= (inputs(150)) or (inputs(147));
    layer0_outputs(10571) <= not(inputs(106));
    layer0_outputs(10572) <= (inputs(122)) and not (inputs(175));
    layer0_outputs(10573) <= (inputs(166)) or (inputs(157));
    layer0_outputs(10574) <= (inputs(223)) xor (inputs(252));
    layer0_outputs(10575) <= (inputs(204)) xor (inputs(156));
    layer0_outputs(10576) <= not(inputs(167)) or (inputs(141));
    layer0_outputs(10577) <= not((inputs(82)) or (inputs(253)));
    layer0_outputs(10578) <= (inputs(135)) and not (inputs(222));
    layer0_outputs(10579) <= not((inputs(109)) or (inputs(185)));
    layer0_outputs(10580) <= '0';
    layer0_outputs(10581) <= not(inputs(77));
    layer0_outputs(10582) <= not(inputs(205));
    layer0_outputs(10583) <= not(inputs(33));
    layer0_outputs(10584) <= not(inputs(223)) or (inputs(140));
    layer0_outputs(10585) <= not((inputs(9)) or (inputs(166)));
    layer0_outputs(10586) <= (inputs(128)) and (inputs(74));
    layer0_outputs(10587) <= (inputs(167)) and not (inputs(90));
    layer0_outputs(10588) <= not((inputs(245)) and (inputs(119)));
    layer0_outputs(10589) <= (inputs(249)) and not (inputs(235));
    layer0_outputs(10590) <= (inputs(7)) or (inputs(28));
    layer0_outputs(10591) <= '1';
    layer0_outputs(10592) <= (inputs(125)) or (inputs(155));
    layer0_outputs(10593) <= '1';
    layer0_outputs(10594) <= (inputs(22)) xor (inputs(161));
    layer0_outputs(10595) <= not(inputs(152)) or (inputs(199));
    layer0_outputs(10596) <= (inputs(42)) xor (inputs(199));
    layer0_outputs(10597) <= (inputs(171)) and not (inputs(45));
    layer0_outputs(10598) <= not((inputs(178)) or (inputs(61)));
    layer0_outputs(10599) <= inputs(65);
    layer0_outputs(10600) <= (inputs(8)) xor (inputs(116));
    layer0_outputs(10601) <= not((inputs(192)) or (inputs(11)));
    layer0_outputs(10602) <= '0';
    layer0_outputs(10603) <= not((inputs(90)) or (inputs(161)));
    layer0_outputs(10604) <= not((inputs(27)) or (inputs(172)));
    layer0_outputs(10605) <= not((inputs(210)) or (inputs(211)));
    layer0_outputs(10606) <= (inputs(33)) xor (inputs(233));
    layer0_outputs(10607) <= inputs(111);
    layer0_outputs(10608) <= '0';
    layer0_outputs(10609) <= (inputs(84)) and (inputs(83));
    layer0_outputs(10610) <= not((inputs(52)) or (inputs(181)));
    layer0_outputs(10611) <= not(inputs(46)) or (inputs(83));
    layer0_outputs(10612) <= not(inputs(72));
    layer0_outputs(10613) <= (inputs(190)) and not (inputs(244));
    layer0_outputs(10614) <= not((inputs(203)) xor (inputs(183)));
    layer0_outputs(10615) <= '1';
    layer0_outputs(10616) <= (inputs(201)) and not (inputs(115));
    layer0_outputs(10617) <= (inputs(207)) xor (inputs(23));
    layer0_outputs(10618) <= inputs(63);
    layer0_outputs(10619) <= (inputs(13)) or (inputs(205));
    layer0_outputs(10620) <= not(inputs(242));
    layer0_outputs(10621) <= inputs(123);
    layer0_outputs(10622) <= not(inputs(150)) or (inputs(211));
    layer0_outputs(10623) <= not(inputs(213)) or (inputs(220));
    layer0_outputs(10624) <= inputs(201);
    layer0_outputs(10625) <= (inputs(82)) or (inputs(34));
    layer0_outputs(10626) <= inputs(118);
    layer0_outputs(10627) <= (inputs(166)) or (inputs(68));
    layer0_outputs(10628) <= not(inputs(42));
    layer0_outputs(10629) <= not(inputs(59)) or (inputs(13));
    layer0_outputs(10630) <= (inputs(229)) or (inputs(69));
    layer0_outputs(10631) <= '1';
    layer0_outputs(10632) <= not(inputs(71));
    layer0_outputs(10633) <= inputs(118);
    layer0_outputs(10634) <= not((inputs(195)) or (inputs(125)));
    layer0_outputs(10635) <= (inputs(140)) and (inputs(183));
    layer0_outputs(10636) <= inputs(119);
    layer0_outputs(10637) <= (inputs(191)) and (inputs(221));
    layer0_outputs(10638) <= not((inputs(146)) and (inputs(68)));
    layer0_outputs(10639) <= (inputs(152)) and (inputs(55));
    layer0_outputs(10640) <= not((inputs(31)) xor (inputs(153)));
    layer0_outputs(10641) <= (inputs(10)) and (inputs(82));
    layer0_outputs(10642) <= not(inputs(137));
    layer0_outputs(10643) <= (inputs(14)) or (inputs(120));
    layer0_outputs(10644) <= not((inputs(245)) xor (inputs(217)));
    layer0_outputs(10645) <= (inputs(47)) or (inputs(184));
    layer0_outputs(10646) <= (inputs(212)) and (inputs(91));
    layer0_outputs(10647) <= not(inputs(201)) or (inputs(18));
    layer0_outputs(10648) <= inputs(125);
    layer0_outputs(10649) <= not(inputs(233)) or (inputs(193));
    layer0_outputs(10650) <= inputs(106);
    layer0_outputs(10651) <= not(inputs(208)) or (inputs(98));
    layer0_outputs(10652) <= not(inputs(144)) or (inputs(227));
    layer0_outputs(10653) <= not((inputs(155)) xor (inputs(79)));
    layer0_outputs(10654) <= (inputs(9)) or (inputs(212));
    layer0_outputs(10655) <= inputs(181);
    layer0_outputs(10656) <= (inputs(169)) and not (inputs(19));
    layer0_outputs(10657) <= (inputs(173)) or (inputs(33));
    layer0_outputs(10658) <= (inputs(157)) or (inputs(179));
    layer0_outputs(10659) <= not(inputs(109));
    layer0_outputs(10660) <= not(inputs(87));
    layer0_outputs(10661) <= not((inputs(42)) or (inputs(197)));
    layer0_outputs(10662) <= (inputs(251)) or (inputs(83));
    layer0_outputs(10663) <= (inputs(228)) or (inputs(186));
    layer0_outputs(10664) <= (inputs(53)) or (inputs(206));
    layer0_outputs(10665) <= not((inputs(111)) xor (inputs(252)));
    layer0_outputs(10666) <= inputs(148);
    layer0_outputs(10667) <= not(inputs(186));
    layer0_outputs(10668) <= inputs(9);
    layer0_outputs(10669) <= inputs(118);
    layer0_outputs(10670) <= not((inputs(137)) xor (inputs(49)));
    layer0_outputs(10671) <= not(inputs(174)) or (inputs(145));
    layer0_outputs(10672) <= not(inputs(62)) or (inputs(7));
    layer0_outputs(10673) <= not((inputs(55)) or (inputs(58)));
    layer0_outputs(10674) <= not((inputs(230)) or (inputs(194)));
    layer0_outputs(10675) <= (inputs(206)) or (inputs(34));
    layer0_outputs(10676) <= not(inputs(165)) or (inputs(195));
    layer0_outputs(10677) <= (inputs(143)) and not (inputs(130));
    layer0_outputs(10678) <= not(inputs(40));
    layer0_outputs(10679) <= not((inputs(14)) xor (inputs(108)));
    layer0_outputs(10680) <= inputs(188);
    layer0_outputs(10681) <= not(inputs(153)) or (inputs(158));
    layer0_outputs(10682) <= not((inputs(157)) xor (inputs(141)));
    layer0_outputs(10683) <= inputs(138);
    layer0_outputs(10684) <= not(inputs(199));
    layer0_outputs(10685) <= (inputs(156)) or (inputs(93));
    layer0_outputs(10686) <= (inputs(176)) or (inputs(177));
    layer0_outputs(10687) <= (inputs(151)) and not (inputs(29));
    layer0_outputs(10688) <= not((inputs(18)) xor (inputs(232)));
    layer0_outputs(10689) <= not((inputs(12)) xor (inputs(109)));
    layer0_outputs(10690) <= (inputs(181)) or (inputs(136));
    layer0_outputs(10691) <= not((inputs(30)) xor (inputs(77)));
    layer0_outputs(10692) <= '1';
    layer0_outputs(10693) <= inputs(201);
    layer0_outputs(10694) <= inputs(120);
    layer0_outputs(10695) <= (inputs(138)) xor (inputs(245));
    layer0_outputs(10696) <= not((inputs(29)) or (inputs(47)));
    layer0_outputs(10697) <= not(inputs(251));
    layer0_outputs(10698) <= (inputs(244)) and not (inputs(78));
    layer0_outputs(10699) <= not(inputs(156));
    layer0_outputs(10700) <= not(inputs(151));
    layer0_outputs(10701) <= not(inputs(103)) or (inputs(190));
    layer0_outputs(10702) <= inputs(238);
    layer0_outputs(10703) <= not((inputs(24)) xor (inputs(29)));
    layer0_outputs(10704) <= (inputs(174)) and not (inputs(223));
    layer0_outputs(10705) <= not((inputs(41)) or (inputs(226)));
    layer0_outputs(10706) <= not((inputs(115)) xor (inputs(112)));
    layer0_outputs(10707) <= not((inputs(20)) xor (inputs(149)));
    layer0_outputs(10708) <= (inputs(41)) and not (inputs(248));
    layer0_outputs(10709) <= (inputs(200)) or (inputs(94));
    layer0_outputs(10710) <= (inputs(188)) or (inputs(9));
    layer0_outputs(10711) <= not((inputs(150)) or (inputs(176)));
    layer0_outputs(10712) <= not((inputs(161)) and (inputs(61)));
    layer0_outputs(10713) <= (inputs(105)) and not (inputs(216));
    layer0_outputs(10714) <= (inputs(152)) xor (inputs(8));
    layer0_outputs(10715) <= not((inputs(59)) and (inputs(59)));
    layer0_outputs(10716) <= (inputs(2)) and (inputs(67));
    layer0_outputs(10717) <= not((inputs(109)) or (inputs(28)));
    layer0_outputs(10718) <= (inputs(90)) and (inputs(108));
    layer0_outputs(10719) <= (inputs(180)) xor (inputs(55));
    layer0_outputs(10720) <= (inputs(38)) or (inputs(193));
    layer0_outputs(10721) <= not(inputs(66));
    layer0_outputs(10722) <= inputs(41);
    layer0_outputs(10723) <= '1';
    layer0_outputs(10724) <= (inputs(95)) and (inputs(92));
    layer0_outputs(10725) <= not((inputs(249)) and (inputs(50)));
    layer0_outputs(10726) <= (inputs(58)) xor (inputs(56));
    layer0_outputs(10727) <= not((inputs(94)) xor (inputs(5)));
    layer0_outputs(10728) <= not((inputs(229)) xor (inputs(53)));
    layer0_outputs(10729) <= (inputs(109)) and not (inputs(25));
    layer0_outputs(10730) <= not(inputs(176)) or (inputs(180));
    layer0_outputs(10731) <= (inputs(236)) and not (inputs(220));
    layer0_outputs(10732) <= not(inputs(44));
    layer0_outputs(10733) <= not((inputs(253)) xor (inputs(240)));
    layer0_outputs(10734) <= (inputs(25)) xor (inputs(30));
    layer0_outputs(10735) <= not((inputs(67)) xor (inputs(61)));
    layer0_outputs(10736) <= (inputs(177)) xor (inputs(56));
    layer0_outputs(10737) <= not((inputs(94)) or (inputs(164)));
    layer0_outputs(10738) <= not((inputs(96)) and (inputs(228)));
    layer0_outputs(10739) <= not((inputs(218)) xor (inputs(214)));
    layer0_outputs(10740) <= not((inputs(21)) or (inputs(196)));
    layer0_outputs(10741) <= (inputs(126)) or (inputs(37));
    layer0_outputs(10742) <= (inputs(198)) and not (inputs(221));
    layer0_outputs(10743) <= (inputs(201)) or (inputs(38));
    layer0_outputs(10744) <= not(inputs(83)) or (inputs(228));
    layer0_outputs(10745) <= not(inputs(222)) or (inputs(35));
    layer0_outputs(10746) <= not(inputs(92));
    layer0_outputs(10747) <= '1';
    layer0_outputs(10748) <= '0';
    layer0_outputs(10749) <= not((inputs(47)) xor (inputs(67)));
    layer0_outputs(10750) <= not(inputs(52)) or (inputs(60));
    layer0_outputs(10751) <= not(inputs(109)) or (inputs(238));
    layer0_outputs(10752) <= not(inputs(72));
    layer0_outputs(10753) <= (inputs(86)) and (inputs(85));
    layer0_outputs(10754) <= not(inputs(220));
    layer0_outputs(10755) <= not((inputs(40)) or (inputs(132)));
    layer0_outputs(10756) <= (inputs(40)) or (inputs(34));
    layer0_outputs(10757) <= (inputs(117)) and not (inputs(254));
    layer0_outputs(10758) <= '0';
    layer0_outputs(10759) <= not((inputs(180)) xor (inputs(53)));
    layer0_outputs(10760) <= not(inputs(23)) or (inputs(238));
    layer0_outputs(10761) <= not(inputs(92)) or (inputs(23));
    layer0_outputs(10762) <= (inputs(14)) and (inputs(222));
    layer0_outputs(10763) <= (inputs(89)) and not (inputs(194));
    layer0_outputs(10764) <= '1';
    layer0_outputs(10765) <= inputs(1);
    layer0_outputs(10766) <= (inputs(85)) or (inputs(162));
    layer0_outputs(10767) <= not(inputs(195));
    layer0_outputs(10768) <= (inputs(23)) or (inputs(147));
    layer0_outputs(10769) <= inputs(132);
    layer0_outputs(10770) <= not(inputs(55));
    layer0_outputs(10771) <= not((inputs(14)) or (inputs(171)));
    layer0_outputs(10772) <= not((inputs(67)) or (inputs(172)));
    layer0_outputs(10773) <= not(inputs(195)) or (inputs(17));
    layer0_outputs(10774) <= not((inputs(123)) or (inputs(230)));
    layer0_outputs(10775) <= (inputs(60)) or (inputs(146));
    layer0_outputs(10776) <= not((inputs(99)) xor (inputs(22)));
    layer0_outputs(10777) <= not((inputs(218)) or (inputs(54)));
    layer0_outputs(10778) <= inputs(131);
    layer0_outputs(10779) <= not(inputs(73));
    layer0_outputs(10780) <= inputs(158);
    layer0_outputs(10781) <= (inputs(150)) and not (inputs(82));
    layer0_outputs(10782) <= (inputs(182)) or (inputs(204));
    layer0_outputs(10783) <= not(inputs(172)) or (inputs(7));
    layer0_outputs(10784) <= not((inputs(156)) xor (inputs(56)));
    layer0_outputs(10785) <= '0';
    layer0_outputs(10786) <= not((inputs(164)) xor (inputs(169)));
    layer0_outputs(10787) <= not((inputs(96)) or (inputs(240)));
    layer0_outputs(10788) <= inputs(58);
    layer0_outputs(10789) <= not(inputs(43)) or (inputs(161));
    layer0_outputs(10790) <= not(inputs(228));
    layer0_outputs(10791) <= not(inputs(143));
    layer0_outputs(10792) <= (inputs(62)) and (inputs(240));
    layer0_outputs(10793) <= (inputs(4)) xor (inputs(154));
    layer0_outputs(10794) <= '0';
    layer0_outputs(10795) <= (inputs(116)) and not (inputs(242));
    layer0_outputs(10796) <= (inputs(163)) or (inputs(49));
    layer0_outputs(10797) <= not((inputs(13)) xor (inputs(52)));
    layer0_outputs(10798) <= (inputs(46)) xor (inputs(41));
    layer0_outputs(10799) <= (inputs(243)) and (inputs(113));
    layer0_outputs(10800) <= (inputs(43)) and not (inputs(225));
    layer0_outputs(10801) <= (inputs(29)) xor (inputs(143));
    layer0_outputs(10802) <= (inputs(169)) xor (inputs(113));
    layer0_outputs(10803) <= not((inputs(22)) xor (inputs(174)));
    layer0_outputs(10804) <= (inputs(159)) or (inputs(100));
    layer0_outputs(10805) <= not(inputs(74)) or (inputs(244));
    layer0_outputs(10806) <= not(inputs(35)) or (inputs(253));
    layer0_outputs(10807) <= (inputs(44)) and not (inputs(177));
    layer0_outputs(10808) <= not(inputs(251));
    layer0_outputs(10809) <= (inputs(52)) or (inputs(110));
    layer0_outputs(10810) <= (inputs(27)) and (inputs(193));
    layer0_outputs(10811) <= (inputs(3)) and not (inputs(130));
    layer0_outputs(10812) <= not(inputs(180)) or (inputs(243));
    layer0_outputs(10813) <= (inputs(161)) or (inputs(246));
    layer0_outputs(10814) <= not(inputs(170)) or (inputs(190));
    layer0_outputs(10815) <= not((inputs(39)) or (inputs(186)));
    layer0_outputs(10816) <= not((inputs(59)) xor (inputs(105)));
    layer0_outputs(10817) <= inputs(42);
    layer0_outputs(10818) <= not((inputs(224)) or (inputs(94)));
    layer0_outputs(10819) <= not((inputs(189)) or (inputs(232)));
    layer0_outputs(10820) <= not((inputs(1)) xor (inputs(137)));
    layer0_outputs(10821) <= inputs(115);
    layer0_outputs(10822) <= (inputs(74)) or (inputs(11));
    layer0_outputs(10823) <= (inputs(1)) or (inputs(163));
    layer0_outputs(10824) <= not((inputs(134)) or (inputs(251)));
    layer0_outputs(10825) <= not((inputs(236)) xor (inputs(152)));
    layer0_outputs(10826) <= not(inputs(200));
    layer0_outputs(10827) <= not((inputs(177)) xor (inputs(235)));
    layer0_outputs(10828) <= inputs(71);
    layer0_outputs(10829) <= not(inputs(152));
    layer0_outputs(10830) <= (inputs(207)) and not (inputs(191));
    layer0_outputs(10831) <= not(inputs(167));
    layer0_outputs(10832) <= not((inputs(165)) xor (inputs(219)));
    layer0_outputs(10833) <= '1';
    layer0_outputs(10834) <= not(inputs(76));
    layer0_outputs(10835) <= not(inputs(115));
    layer0_outputs(10836) <= (inputs(66)) or (inputs(76));
    layer0_outputs(10837) <= inputs(141);
    layer0_outputs(10838) <= not(inputs(99));
    layer0_outputs(10839) <= (inputs(249)) xor (inputs(22));
    layer0_outputs(10840) <= not(inputs(233));
    layer0_outputs(10841) <= (inputs(71)) and not (inputs(42));
    layer0_outputs(10842) <= (inputs(16)) or (inputs(238));
    layer0_outputs(10843) <= '0';
    layer0_outputs(10844) <= not(inputs(234)) or (inputs(234));
    layer0_outputs(10845) <= (inputs(163)) and (inputs(129));
    layer0_outputs(10846) <= (inputs(7)) and (inputs(67));
    layer0_outputs(10847) <= not((inputs(103)) and (inputs(14)));
    layer0_outputs(10848) <= (inputs(92)) and not (inputs(87));
    layer0_outputs(10849) <= (inputs(109)) or (inputs(132));
    layer0_outputs(10850) <= (inputs(86)) and not (inputs(59));
    layer0_outputs(10851) <= (inputs(30)) xor (inputs(106));
    layer0_outputs(10852) <= not((inputs(75)) xor (inputs(130)));
    layer0_outputs(10853) <= not((inputs(198)) xor (inputs(180)));
    layer0_outputs(10854) <= (inputs(231)) xor (inputs(186));
    layer0_outputs(10855) <= (inputs(139)) xor (inputs(142));
    layer0_outputs(10856) <= (inputs(29)) and not (inputs(62));
    layer0_outputs(10857) <= not((inputs(245)) or (inputs(248)));
    layer0_outputs(10858) <= not(inputs(118)) or (inputs(68));
    layer0_outputs(10859) <= (inputs(52)) and not (inputs(242));
    layer0_outputs(10860) <= (inputs(184)) and not (inputs(146));
    layer0_outputs(10861) <= not((inputs(219)) or (inputs(91)));
    layer0_outputs(10862) <= inputs(185);
    layer0_outputs(10863) <= (inputs(177)) or (inputs(22));
    layer0_outputs(10864) <= (inputs(39)) xor (inputs(74));
    layer0_outputs(10865) <= (inputs(93)) xor (inputs(139));
    layer0_outputs(10866) <= (inputs(191)) xor (inputs(74));
    layer0_outputs(10867) <= inputs(108);
    layer0_outputs(10868) <= not(inputs(41)) or (inputs(44));
    layer0_outputs(10869) <= '0';
    layer0_outputs(10870) <= not(inputs(117)) or (inputs(231));
    layer0_outputs(10871) <= (inputs(246)) and (inputs(250));
    layer0_outputs(10872) <= not(inputs(157));
    layer0_outputs(10873) <= not(inputs(69));
    layer0_outputs(10874) <= (inputs(141)) or (inputs(241));
    layer0_outputs(10875) <= not((inputs(243)) xor (inputs(172)));
    layer0_outputs(10876) <= not(inputs(170));
    layer0_outputs(10877) <= not(inputs(150)) or (inputs(78));
    layer0_outputs(10878) <= not((inputs(184)) xor (inputs(3)));
    layer0_outputs(10879) <= not((inputs(108)) or (inputs(40)));
    layer0_outputs(10880) <= inputs(170);
    layer0_outputs(10881) <= (inputs(161)) xor (inputs(130));
    layer0_outputs(10882) <= not(inputs(199));
    layer0_outputs(10883) <= (inputs(242)) and not (inputs(15));
    layer0_outputs(10884) <= not((inputs(142)) xor (inputs(219)));
    layer0_outputs(10885) <= (inputs(90)) and not (inputs(45));
    layer0_outputs(10886) <= (inputs(20)) or (inputs(103));
    layer0_outputs(10887) <= not((inputs(150)) or (inputs(131)));
    layer0_outputs(10888) <= inputs(160);
    layer0_outputs(10889) <= (inputs(169)) and not (inputs(240));
    layer0_outputs(10890) <= inputs(152);
    layer0_outputs(10891) <= not((inputs(180)) or (inputs(175)));
    layer0_outputs(10892) <= not((inputs(89)) or (inputs(185)));
    layer0_outputs(10893) <= '0';
    layer0_outputs(10894) <= not((inputs(180)) xor (inputs(137)));
    layer0_outputs(10895) <= (inputs(154)) or (inputs(77));
    layer0_outputs(10896) <= (inputs(220)) or (inputs(10));
    layer0_outputs(10897) <= not((inputs(147)) or (inputs(101)));
    layer0_outputs(10898) <= not((inputs(54)) or (inputs(175)));
    layer0_outputs(10899) <= (inputs(239)) and not (inputs(241));
    layer0_outputs(10900) <= not(inputs(70)) or (inputs(30));
    layer0_outputs(10901) <= (inputs(83)) xor (inputs(70));
    layer0_outputs(10902) <= (inputs(176)) xor (inputs(132));
    layer0_outputs(10903) <= not(inputs(55)) or (inputs(4));
    layer0_outputs(10904) <= not((inputs(172)) or (inputs(159)));
    layer0_outputs(10905) <= (inputs(253)) xor (inputs(64));
    layer0_outputs(10906) <= not(inputs(130)) or (inputs(157));
    layer0_outputs(10907) <= (inputs(190)) xor (inputs(103));
    layer0_outputs(10908) <= not(inputs(133));
    layer0_outputs(10909) <= inputs(203);
    layer0_outputs(10910) <= (inputs(51)) and not (inputs(225));
    layer0_outputs(10911) <= '0';
    layer0_outputs(10912) <= (inputs(28)) xor (inputs(69));
    layer0_outputs(10913) <= (inputs(202)) and not (inputs(111));
    layer0_outputs(10914) <= inputs(236);
    layer0_outputs(10915) <= (inputs(70)) and (inputs(188));
    layer0_outputs(10916) <= inputs(36);
    layer0_outputs(10917) <= not(inputs(86));
    layer0_outputs(10918) <= not(inputs(234)) or (inputs(78));
    layer0_outputs(10919) <= not((inputs(37)) xor (inputs(84)));
    layer0_outputs(10920) <= inputs(83);
    layer0_outputs(10921) <= not(inputs(72));
    layer0_outputs(10922) <= not(inputs(179));
    layer0_outputs(10923) <= inputs(76);
    layer0_outputs(10924) <= (inputs(81)) xor (inputs(228));
    layer0_outputs(10925) <= (inputs(228)) xor (inputs(143));
    layer0_outputs(10926) <= not((inputs(167)) or (inputs(108)));
    layer0_outputs(10927) <= not(inputs(164)) or (inputs(229));
    layer0_outputs(10928) <= not((inputs(233)) xor (inputs(5)));
    layer0_outputs(10929) <= not((inputs(124)) xor (inputs(50)));
    layer0_outputs(10930) <= (inputs(204)) or (inputs(138));
    layer0_outputs(10931) <= (inputs(227)) xor (inputs(69));
    layer0_outputs(10932) <= not((inputs(154)) xor (inputs(85)));
    layer0_outputs(10933) <= not(inputs(88));
    layer0_outputs(10934) <= (inputs(116)) and (inputs(160));
    layer0_outputs(10935) <= not(inputs(36)) or (inputs(4));
    layer0_outputs(10936) <= (inputs(114)) or (inputs(149));
    layer0_outputs(10937) <= (inputs(235)) and (inputs(53));
    layer0_outputs(10938) <= (inputs(2)) or (inputs(39));
    layer0_outputs(10939) <= not(inputs(55)) or (inputs(248));
    layer0_outputs(10940) <= inputs(112);
    layer0_outputs(10941) <= not((inputs(235)) or (inputs(59)));
    layer0_outputs(10942) <= not((inputs(89)) or (inputs(82)));
    layer0_outputs(10943) <= not(inputs(32)) or (inputs(240));
    layer0_outputs(10944) <= (inputs(121)) and not (inputs(34));
    layer0_outputs(10945) <= inputs(107);
    layer0_outputs(10946) <= inputs(211);
    layer0_outputs(10947) <= (inputs(245)) xor (inputs(206));
    layer0_outputs(10948) <= (inputs(26)) xor (inputs(162));
    layer0_outputs(10949) <= (inputs(13)) or (inputs(100));
    layer0_outputs(10950) <= not((inputs(33)) or (inputs(202)));
    layer0_outputs(10951) <= not(inputs(84));
    layer0_outputs(10952) <= not(inputs(167));
    layer0_outputs(10953) <= (inputs(250)) and not (inputs(237));
    layer0_outputs(10954) <= not((inputs(132)) xor (inputs(101)));
    layer0_outputs(10955) <= not(inputs(59));
    layer0_outputs(10956) <= inputs(177);
    layer0_outputs(10957) <= (inputs(17)) xor (inputs(148));
    layer0_outputs(10958) <= not((inputs(26)) xor (inputs(255)));
    layer0_outputs(10959) <= not(inputs(145));
    layer0_outputs(10960) <= not(inputs(237)) or (inputs(78));
    layer0_outputs(10961) <= (inputs(193)) xor (inputs(53));
    layer0_outputs(10962) <= not(inputs(44)) or (inputs(32));
    layer0_outputs(10963) <= not((inputs(251)) or (inputs(95)));
    layer0_outputs(10964) <= (inputs(143)) and not (inputs(30));
    layer0_outputs(10965) <= not((inputs(200)) xor (inputs(191)));
    layer0_outputs(10966) <= not((inputs(158)) or (inputs(248)));
    layer0_outputs(10967) <= not((inputs(53)) xor (inputs(97)));
    layer0_outputs(10968) <= (inputs(58)) xor (inputs(8));
    layer0_outputs(10969) <= not(inputs(87));
    layer0_outputs(10970) <= not((inputs(138)) or (inputs(83)));
    layer0_outputs(10971) <= not(inputs(181));
    layer0_outputs(10972) <= (inputs(227)) and not (inputs(98));
    layer0_outputs(10973) <= not(inputs(185));
    layer0_outputs(10974) <= not(inputs(41));
    layer0_outputs(10975) <= not(inputs(251)) or (inputs(242));
    layer0_outputs(10976) <= '0';
    layer0_outputs(10977) <= inputs(117);
    layer0_outputs(10978) <= not((inputs(83)) xor (inputs(155)));
    layer0_outputs(10979) <= inputs(187);
    layer0_outputs(10980) <= (inputs(152)) or (inputs(9));
    layer0_outputs(10981) <= not(inputs(177));
    layer0_outputs(10982) <= inputs(37);
    layer0_outputs(10983) <= not((inputs(38)) xor (inputs(209)));
    layer0_outputs(10984) <= not(inputs(107));
    layer0_outputs(10985) <= inputs(52);
    layer0_outputs(10986) <= not(inputs(110));
    layer0_outputs(10987) <= not((inputs(68)) xor (inputs(73)));
    layer0_outputs(10988) <= (inputs(68)) xor (inputs(90));
    layer0_outputs(10989) <= not((inputs(18)) and (inputs(248)));
    layer0_outputs(10990) <= not(inputs(57)) or (inputs(44));
    layer0_outputs(10991) <= inputs(243);
    layer0_outputs(10992) <= (inputs(120)) xor (inputs(187));
    layer0_outputs(10993) <= inputs(88);
    layer0_outputs(10994) <= not(inputs(118));
    layer0_outputs(10995) <= not((inputs(177)) or (inputs(185)));
    layer0_outputs(10996) <= not((inputs(41)) or (inputs(63)));
    layer0_outputs(10997) <= not((inputs(65)) or (inputs(61)));
    layer0_outputs(10998) <= not(inputs(53)) or (inputs(54));
    layer0_outputs(10999) <= not(inputs(92));
    layer0_outputs(11000) <= inputs(76);
    layer0_outputs(11001) <= not(inputs(157)) or (inputs(230));
    layer0_outputs(11002) <= not(inputs(149));
    layer0_outputs(11003) <= not(inputs(252));
    layer0_outputs(11004) <= not(inputs(51));
    layer0_outputs(11005) <= (inputs(253)) xor (inputs(96));
    layer0_outputs(11006) <= (inputs(32)) xor (inputs(30));
    layer0_outputs(11007) <= (inputs(85)) and not (inputs(5));
    layer0_outputs(11008) <= '1';
    layer0_outputs(11009) <= not(inputs(53)) or (inputs(11));
    layer0_outputs(11010) <= not(inputs(171));
    layer0_outputs(11011) <= (inputs(196)) and not (inputs(145));
    layer0_outputs(11012) <= not(inputs(192)) or (inputs(248));
    layer0_outputs(11013) <= (inputs(143)) xor (inputs(169));
    layer0_outputs(11014) <= (inputs(65)) xor (inputs(231));
    layer0_outputs(11015) <= not((inputs(39)) xor (inputs(14)));
    layer0_outputs(11016) <= not(inputs(133));
    layer0_outputs(11017) <= not(inputs(73)) or (inputs(154));
    layer0_outputs(11018) <= not((inputs(234)) or (inputs(140)));
    layer0_outputs(11019) <= inputs(44);
    layer0_outputs(11020) <= '1';
    layer0_outputs(11021) <= not((inputs(51)) xor (inputs(199)));
    layer0_outputs(11022) <= inputs(55);
    layer0_outputs(11023) <= not((inputs(5)) and (inputs(2)));
    layer0_outputs(11024) <= inputs(41);
    layer0_outputs(11025) <= (inputs(194)) xor (inputs(159));
    layer0_outputs(11026) <= (inputs(62)) or (inputs(150));
    layer0_outputs(11027) <= (inputs(14)) xor (inputs(76));
    layer0_outputs(11028) <= not(inputs(169)) or (inputs(125));
    layer0_outputs(11029) <= inputs(220);
    layer0_outputs(11030) <= not(inputs(8)) or (inputs(189));
    layer0_outputs(11031) <= inputs(99);
    layer0_outputs(11032) <= (inputs(23)) and not (inputs(112));
    layer0_outputs(11033) <= inputs(120);
    layer0_outputs(11034) <= (inputs(0)) xor (inputs(224));
    layer0_outputs(11035) <= not(inputs(56)) or (inputs(230));
    layer0_outputs(11036) <= not((inputs(98)) or (inputs(128)));
    layer0_outputs(11037) <= (inputs(252)) and not (inputs(194));
    layer0_outputs(11038) <= not(inputs(247)) or (inputs(10));
    layer0_outputs(11039) <= not(inputs(114)) or (inputs(112));
    layer0_outputs(11040) <= inputs(71);
    layer0_outputs(11041) <= (inputs(12)) and (inputs(211));
    layer0_outputs(11042) <= not(inputs(64)) or (inputs(215));
    layer0_outputs(11043) <= inputs(104);
    layer0_outputs(11044) <= (inputs(75)) xor (inputs(169));
    layer0_outputs(11045) <= inputs(224);
    layer0_outputs(11046) <= (inputs(3)) or (inputs(83));
    layer0_outputs(11047) <= (inputs(173)) and (inputs(223));
    layer0_outputs(11048) <= inputs(120);
    layer0_outputs(11049) <= not(inputs(214)) or (inputs(13));
    layer0_outputs(11050) <= not(inputs(122));
    layer0_outputs(11051) <= not((inputs(250)) xor (inputs(107)));
    layer0_outputs(11052) <= not(inputs(96)) or (inputs(90));
    layer0_outputs(11053) <= not(inputs(31));
    layer0_outputs(11054) <= not((inputs(160)) xor (inputs(247)));
    layer0_outputs(11055) <= not(inputs(149)) or (inputs(36));
    layer0_outputs(11056) <= not((inputs(204)) or (inputs(148)));
    layer0_outputs(11057) <= not((inputs(130)) or (inputs(232)));
    layer0_outputs(11058) <= (inputs(60)) or (inputs(148));
    layer0_outputs(11059) <= not((inputs(73)) xor (inputs(125)));
    layer0_outputs(11060) <= (inputs(79)) xor (inputs(96));
    layer0_outputs(11061) <= (inputs(117)) and not (inputs(129));
    layer0_outputs(11062) <= not(inputs(159));
    layer0_outputs(11063) <= inputs(202);
    layer0_outputs(11064) <= '1';
    layer0_outputs(11065) <= not((inputs(92)) or (inputs(158)));
    layer0_outputs(11066) <= not(inputs(195));
    layer0_outputs(11067) <= not(inputs(132)) or (inputs(196));
    layer0_outputs(11068) <= (inputs(112)) xor (inputs(38));
    layer0_outputs(11069) <= (inputs(23)) or (inputs(125));
    layer0_outputs(11070) <= (inputs(59)) or (inputs(83));
    layer0_outputs(11071) <= not(inputs(133));
    layer0_outputs(11072) <= (inputs(164)) and not (inputs(114));
    layer0_outputs(11073) <= (inputs(241)) and (inputs(44));
    layer0_outputs(11074) <= '1';
    layer0_outputs(11075) <= not(inputs(144));
    layer0_outputs(11076) <= not(inputs(63));
    layer0_outputs(11077) <= (inputs(204)) and not (inputs(64));
    layer0_outputs(11078) <= not(inputs(151));
    layer0_outputs(11079) <= inputs(51);
    layer0_outputs(11080) <= (inputs(57)) xor (inputs(134));
    layer0_outputs(11081) <= (inputs(68)) and not (inputs(247));
    layer0_outputs(11082) <= (inputs(221)) xor (inputs(92));
    layer0_outputs(11083) <= inputs(233);
    layer0_outputs(11084) <= (inputs(102)) and not (inputs(55));
    layer0_outputs(11085) <= (inputs(187)) or (inputs(94));
    layer0_outputs(11086) <= not(inputs(138));
    layer0_outputs(11087) <= not(inputs(233));
    layer0_outputs(11088) <= (inputs(25)) or (inputs(33));
    layer0_outputs(11089) <= not((inputs(25)) or (inputs(227)));
    layer0_outputs(11090) <= not(inputs(139));
    layer0_outputs(11091) <= inputs(87);
    layer0_outputs(11092) <= (inputs(219)) and not (inputs(245));
    layer0_outputs(11093) <= not((inputs(215)) xor (inputs(231)));
    layer0_outputs(11094) <= not((inputs(11)) or (inputs(215)));
    layer0_outputs(11095) <= (inputs(99)) xor (inputs(228));
    layer0_outputs(11096) <= inputs(214);
    layer0_outputs(11097) <= not((inputs(111)) xor (inputs(70)));
    layer0_outputs(11098) <= inputs(237);
    layer0_outputs(11099) <= not(inputs(89)) or (inputs(57));
    layer0_outputs(11100) <= (inputs(25)) or (inputs(137));
    layer0_outputs(11101) <= not(inputs(97)) or (inputs(76));
    layer0_outputs(11102) <= (inputs(78)) and not (inputs(205));
    layer0_outputs(11103) <= (inputs(139)) and not (inputs(21));
    layer0_outputs(11104) <= inputs(148);
    layer0_outputs(11105) <= not(inputs(122)) or (inputs(238));
    layer0_outputs(11106) <= (inputs(192)) and not (inputs(27));
    layer0_outputs(11107) <= not((inputs(240)) xor (inputs(48)));
    layer0_outputs(11108) <= (inputs(134)) and not (inputs(186));
    layer0_outputs(11109) <= (inputs(216)) or (inputs(36));
    layer0_outputs(11110) <= (inputs(232)) xor (inputs(200));
    layer0_outputs(11111) <= not(inputs(81));
    layer0_outputs(11112) <= (inputs(60)) or (inputs(154));
    layer0_outputs(11113) <= inputs(113);
    layer0_outputs(11114) <= (inputs(241)) or (inputs(215));
    layer0_outputs(11115) <= not((inputs(78)) and (inputs(34)));
    layer0_outputs(11116) <= not((inputs(117)) xor (inputs(161)));
    layer0_outputs(11117) <= not((inputs(101)) or (inputs(45)));
    layer0_outputs(11118) <= (inputs(0)) xor (inputs(73));
    layer0_outputs(11119) <= inputs(189);
    layer0_outputs(11120) <= not((inputs(167)) xor (inputs(131)));
    layer0_outputs(11121) <= '1';
    layer0_outputs(11122) <= not((inputs(226)) or (inputs(89)));
    layer0_outputs(11123) <= '1';
    layer0_outputs(11124) <= (inputs(202)) and not (inputs(46));
    layer0_outputs(11125) <= inputs(125);
    layer0_outputs(11126) <= not((inputs(203)) xor (inputs(170)));
    layer0_outputs(11127) <= not((inputs(114)) xor (inputs(180)));
    layer0_outputs(11128) <= inputs(136);
    layer0_outputs(11129) <= not(inputs(116));
    layer0_outputs(11130) <= (inputs(122)) and not (inputs(110));
    layer0_outputs(11131) <= '0';
    layer0_outputs(11132) <= (inputs(170)) or (inputs(235));
    layer0_outputs(11133) <= not((inputs(85)) or (inputs(224)));
    layer0_outputs(11134) <= not((inputs(201)) or (inputs(221)));
    layer0_outputs(11135) <= inputs(173);
    layer0_outputs(11136) <= inputs(214);
    layer0_outputs(11137) <= inputs(179);
    layer0_outputs(11138) <= (inputs(33)) and not (inputs(33));
    layer0_outputs(11139) <= not(inputs(70));
    layer0_outputs(11140) <= (inputs(31)) or (inputs(6));
    layer0_outputs(11141) <= (inputs(136)) and not (inputs(212));
    layer0_outputs(11142) <= not(inputs(130));
    layer0_outputs(11143) <= not(inputs(140)) or (inputs(210));
    layer0_outputs(11144) <= inputs(55);
    layer0_outputs(11145) <= (inputs(34)) and (inputs(247));
    layer0_outputs(11146) <= inputs(95);
    layer0_outputs(11147) <= (inputs(118)) and not (inputs(148));
    layer0_outputs(11148) <= (inputs(168)) or (inputs(231));
    layer0_outputs(11149) <= (inputs(167)) and not (inputs(239));
    layer0_outputs(11150) <= (inputs(89)) or (inputs(233));
    layer0_outputs(11151) <= not((inputs(148)) xor (inputs(48)));
    layer0_outputs(11152) <= (inputs(134)) or (inputs(62));
    layer0_outputs(11153) <= inputs(125);
    layer0_outputs(11154) <= (inputs(254)) and not (inputs(29));
    layer0_outputs(11155) <= not(inputs(135));
    layer0_outputs(11156) <= not(inputs(140)) or (inputs(66));
    layer0_outputs(11157) <= not(inputs(118));
    layer0_outputs(11158) <= inputs(186);
    layer0_outputs(11159) <= not((inputs(2)) or (inputs(136)));
    layer0_outputs(11160) <= (inputs(185)) or (inputs(83));
    layer0_outputs(11161) <= not(inputs(175)) or (inputs(77));
    layer0_outputs(11162) <= not(inputs(88)) or (inputs(202));
    layer0_outputs(11163) <= (inputs(36)) or (inputs(70));
    layer0_outputs(11164) <= inputs(72);
    layer0_outputs(11165) <= (inputs(1)) or (inputs(41));
    layer0_outputs(11166) <= (inputs(69)) and not (inputs(237));
    layer0_outputs(11167) <= inputs(12);
    layer0_outputs(11168) <= not(inputs(219)) or (inputs(209));
    layer0_outputs(11169) <= inputs(57);
    layer0_outputs(11170) <= not(inputs(116)) or (inputs(27));
    layer0_outputs(11171) <= not((inputs(28)) or (inputs(26)));
    layer0_outputs(11172) <= inputs(103);
    layer0_outputs(11173) <= (inputs(93)) xor (inputs(18));
    layer0_outputs(11174) <= (inputs(194)) or (inputs(202));
    layer0_outputs(11175) <= not(inputs(207)) or (inputs(248));
    layer0_outputs(11176) <= not((inputs(150)) or (inputs(31)));
    layer0_outputs(11177) <= not(inputs(17));
    layer0_outputs(11178) <= not((inputs(113)) xor (inputs(30)));
    layer0_outputs(11179) <= (inputs(108)) xor (inputs(177));
    layer0_outputs(11180) <= (inputs(131)) xor (inputs(240));
    layer0_outputs(11181) <= (inputs(205)) or (inputs(71));
    layer0_outputs(11182) <= not((inputs(53)) or (inputs(194)));
    layer0_outputs(11183) <= (inputs(192)) xor (inputs(210));
    layer0_outputs(11184) <= inputs(168);
    layer0_outputs(11185) <= '1';
    layer0_outputs(11186) <= (inputs(43)) or (inputs(5));
    layer0_outputs(11187) <= inputs(193);
    layer0_outputs(11188) <= (inputs(2)) and not (inputs(245));
    layer0_outputs(11189) <= not((inputs(78)) or (inputs(247)));
    layer0_outputs(11190) <= '0';
    layer0_outputs(11191) <= (inputs(207)) xor (inputs(162));
    layer0_outputs(11192) <= not((inputs(161)) or (inputs(25)));
    layer0_outputs(11193) <= not((inputs(135)) xor (inputs(232)));
    layer0_outputs(11194) <= (inputs(55)) and not (inputs(66));
    layer0_outputs(11195) <= (inputs(195)) and not (inputs(16));
    layer0_outputs(11196) <= inputs(56);
    layer0_outputs(11197) <= (inputs(208)) xor (inputs(84));
    layer0_outputs(11198) <= inputs(24);
    layer0_outputs(11199) <= (inputs(222)) and not (inputs(71));
    layer0_outputs(11200) <= (inputs(166)) and not (inputs(250));
    layer0_outputs(11201) <= not(inputs(226)) or (inputs(35));
    layer0_outputs(11202) <= (inputs(223)) or (inputs(135));
    layer0_outputs(11203) <= not(inputs(150)) or (inputs(5));
    layer0_outputs(11204) <= not(inputs(77));
    layer0_outputs(11205) <= not((inputs(107)) or (inputs(194)));
    layer0_outputs(11206) <= inputs(63);
    layer0_outputs(11207) <= (inputs(72)) and not (inputs(177));
    layer0_outputs(11208) <= not((inputs(244)) or (inputs(229)));
    layer0_outputs(11209) <= (inputs(9)) or (inputs(138));
    layer0_outputs(11210) <= inputs(101);
    layer0_outputs(11211) <= not((inputs(3)) xor (inputs(163)));
    layer0_outputs(11212) <= inputs(181);
    layer0_outputs(11213) <= not(inputs(138));
    layer0_outputs(11214) <= not(inputs(116));
    layer0_outputs(11215) <= not(inputs(21));
    layer0_outputs(11216) <= '1';
    layer0_outputs(11217) <= (inputs(168)) xor (inputs(13));
    layer0_outputs(11218) <= inputs(99);
    layer0_outputs(11219) <= '1';
    layer0_outputs(11220) <= not((inputs(237)) xor (inputs(120)));
    layer0_outputs(11221) <= (inputs(142)) and (inputs(15));
    layer0_outputs(11222) <= not((inputs(38)) and (inputs(141)));
    layer0_outputs(11223) <= not(inputs(219)) or (inputs(114));
    layer0_outputs(11224) <= not(inputs(64)) or (inputs(175));
    layer0_outputs(11225) <= (inputs(56)) or (inputs(192));
    layer0_outputs(11226) <= (inputs(67)) xor (inputs(46));
    layer0_outputs(11227) <= (inputs(164)) xor (inputs(18));
    layer0_outputs(11228) <= (inputs(229)) or (inputs(135));
    layer0_outputs(11229) <= (inputs(196)) or (inputs(18));
    layer0_outputs(11230) <= not(inputs(189)) or (inputs(49));
    layer0_outputs(11231) <= (inputs(160)) xor (inputs(16));
    layer0_outputs(11232) <= (inputs(185)) and not (inputs(13));
    layer0_outputs(11233) <= (inputs(98)) or (inputs(226));
    layer0_outputs(11234) <= not((inputs(102)) or (inputs(140)));
    layer0_outputs(11235) <= not((inputs(111)) or (inputs(185)));
    layer0_outputs(11236) <= inputs(136);
    layer0_outputs(11237) <= not((inputs(216)) or (inputs(81)));
    layer0_outputs(11238) <= not(inputs(94)) or (inputs(241));
    layer0_outputs(11239) <= (inputs(99)) xor (inputs(90));
    layer0_outputs(11240) <= not((inputs(120)) xor (inputs(5)));
    layer0_outputs(11241) <= inputs(153);
    layer0_outputs(11242) <= not(inputs(81));
    layer0_outputs(11243) <= inputs(181);
    layer0_outputs(11244) <= inputs(186);
    layer0_outputs(11245) <= inputs(187);
    layer0_outputs(11246) <= (inputs(80)) xor (inputs(155));
    layer0_outputs(11247) <= (inputs(178)) or (inputs(202));
    layer0_outputs(11248) <= not(inputs(102));
    layer0_outputs(11249) <= not((inputs(140)) or (inputs(73)));
    layer0_outputs(11250) <= not((inputs(115)) or (inputs(20)));
    layer0_outputs(11251) <= (inputs(168)) and not (inputs(160));
    layer0_outputs(11252) <= inputs(53);
    layer0_outputs(11253) <= inputs(12);
    layer0_outputs(11254) <= not((inputs(196)) xor (inputs(30)));
    layer0_outputs(11255) <= not((inputs(65)) xor (inputs(68)));
    layer0_outputs(11256) <= (inputs(178)) and not (inputs(223));
    layer0_outputs(11257) <= not((inputs(12)) xor (inputs(207)));
    layer0_outputs(11258) <= not((inputs(170)) or (inputs(149)));
    layer0_outputs(11259) <= not(inputs(96));
    layer0_outputs(11260) <= (inputs(212)) xor (inputs(237));
    layer0_outputs(11261) <= (inputs(144)) and not (inputs(22));
    layer0_outputs(11262) <= not(inputs(120));
    layer0_outputs(11263) <= not((inputs(180)) or (inputs(15)));
    layer0_outputs(11264) <= (inputs(113)) and not (inputs(228));
    layer0_outputs(11265) <= not(inputs(238));
    layer0_outputs(11266) <= not(inputs(130));
    layer0_outputs(11267) <= inputs(115);
    layer0_outputs(11268) <= not((inputs(53)) and (inputs(3)));
    layer0_outputs(11269) <= not(inputs(60));
    layer0_outputs(11270) <= (inputs(14)) and (inputs(0));
    layer0_outputs(11271) <= '1';
    layer0_outputs(11272) <= (inputs(192)) or (inputs(237));
    layer0_outputs(11273) <= not(inputs(62));
    layer0_outputs(11274) <= (inputs(45)) xor (inputs(120));
    layer0_outputs(11275) <= not((inputs(142)) and (inputs(207)));
    layer0_outputs(11276) <= inputs(172);
    layer0_outputs(11277) <= not((inputs(235)) xor (inputs(117)));
    layer0_outputs(11278) <= inputs(58);
    layer0_outputs(11279) <= not(inputs(70)) or (inputs(254));
    layer0_outputs(11280) <= (inputs(166)) and not (inputs(246));
    layer0_outputs(11281) <= (inputs(173)) xor (inputs(107));
    layer0_outputs(11282) <= (inputs(169)) and not (inputs(206));
    layer0_outputs(11283) <= not(inputs(203));
    layer0_outputs(11284) <= inputs(166);
    layer0_outputs(11285) <= inputs(105);
    layer0_outputs(11286) <= not((inputs(147)) and (inputs(246)));
    layer0_outputs(11287) <= not((inputs(155)) and (inputs(102)));
    layer0_outputs(11288) <= inputs(189);
    layer0_outputs(11289) <= not(inputs(41)) or (inputs(244));
    layer0_outputs(11290) <= not(inputs(141)) or (inputs(27));
    layer0_outputs(11291) <= not((inputs(189)) xor (inputs(205)));
    layer0_outputs(11292) <= not(inputs(70));
    layer0_outputs(11293) <= not(inputs(122)) or (inputs(59));
    layer0_outputs(11294) <= (inputs(102)) and not (inputs(98));
    layer0_outputs(11295) <= '0';
    layer0_outputs(11296) <= not((inputs(91)) xor (inputs(6)));
    layer0_outputs(11297) <= not((inputs(209)) xor (inputs(215)));
    layer0_outputs(11298) <= (inputs(230)) or (inputs(192));
    layer0_outputs(11299) <= not((inputs(141)) or (inputs(162)));
    layer0_outputs(11300) <= (inputs(139)) and not (inputs(238));
    layer0_outputs(11301) <= (inputs(50)) and (inputs(95));
    layer0_outputs(11302) <= '1';
    layer0_outputs(11303) <= not(inputs(209)) or (inputs(7));
    layer0_outputs(11304) <= not((inputs(161)) or (inputs(228)));
    layer0_outputs(11305) <= (inputs(192)) xor (inputs(109));
    layer0_outputs(11306) <= not((inputs(35)) or (inputs(42)));
    layer0_outputs(11307) <= (inputs(101)) and not (inputs(208));
    layer0_outputs(11308) <= (inputs(194)) and not (inputs(63));
    layer0_outputs(11309) <= not((inputs(138)) xor (inputs(149)));
    layer0_outputs(11310) <= inputs(89);
    layer0_outputs(11311) <= inputs(168);
    layer0_outputs(11312) <= (inputs(140)) and not (inputs(114));
    layer0_outputs(11313) <= not(inputs(109)) or (inputs(143));
    layer0_outputs(11314) <= (inputs(193)) xor (inputs(122));
    layer0_outputs(11315) <= (inputs(99)) or (inputs(196));
    layer0_outputs(11316) <= (inputs(243)) and not (inputs(244));
    layer0_outputs(11317) <= (inputs(209)) xor (inputs(75));
    layer0_outputs(11318) <= (inputs(23)) or (inputs(195));
    layer0_outputs(11319) <= inputs(76);
    layer0_outputs(11320) <= (inputs(248)) and not (inputs(174));
    layer0_outputs(11321) <= inputs(70);
    layer0_outputs(11322) <= inputs(179);
    layer0_outputs(11323) <= not((inputs(143)) or (inputs(166)));
    layer0_outputs(11324) <= inputs(214);
    layer0_outputs(11325) <= (inputs(93)) xor (inputs(42));
    layer0_outputs(11326) <= (inputs(102)) xor (inputs(153));
    layer0_outputs(11327) <= not((inputs(130)) and (inputs(198)));
    layer0_outputs(11328) <= not((inputs(144)) or (inputs(200)));
    layer0_outputs(11329) <= not(inputs(125));
    layer0_outputs(11330) <= inputs(183);
    layer0_outputs(11331) <= (inputs(201)) or (inputs(65));
    layer0_outputs(11332) <= not(inputs(49));
    layer0_outputs(11333) <= not((inputs(51)) and (inputs(126)));
    layer0_outputs(11334) <= inputs(148);
    layer0_outputs(11335) <= (inputs(110)) xor (inputs(52));
    layer0_outputs(11336) <= (inputs(85)) and not (inputs(203));
    layer0_outputs(11337) <= (inputs(50)) or (inputs(236));
    layer0_outputs(11338) <= (inputs(98)) or (inputs(41));
    layer0_outputs(11339) <= (inputs(87)) and not (inputs(142));
    layer0_outputs(11340) <= (inputs(176)) or (inputs(182));
    layer0_outputs(11341) <= not(inputs(219));
    layer0_outputs(11342) <= not((inputs(54)) xor (inputs(108)));
    layer0_outputs(11343) <= inputs(51);
    layer0_outputs(11344) <= (inputs(54)) or (inputs(162));
    layer0_outputs(11345) <= not(inputs(195));
    layer0_outputs(11346) <= not((inputs(21)) and (inputs(71)));
    layer0_outputs(11347) <= not(inputs(113));
    layer0_outputs(11348) <= not(inputs(67)) or (inputs(249));
    layer0_outputs(11349) <= not((inputs(124)) xor (inputs(242)));
    layer0_outputs(11350) <= (inputs(171)) and (inputs(152));
    layer0_outputs(11351) <= (inputs(102)) xor (inputs(241));
    layer0_outputs(11352) <= (inputs(90)) and not (inputs(232));
    layer0_outputs(11353) <= (inputs(238)) or (inputs(40));
    layer0_outputs(11354) <= (inputs(56)) and not (inputs(192));
    layer0_outputs(11355) <= not((inputs(176)) and (inputs(2)));
    layer0_outputs(11356) <= not((inputs(198)) or (inputs(125)));
    layer0_outputs(11357) <= not(inputs(185)) or (inputs(83));
    layer0_outputs(11358) <= not(inputs(172));
    layer0_outputs(11359) <= not(inputs(153));
    layer0_outputs(11360) <= not(inputs(185));
    layer0_outputs(11361) <= not((inputs(48)) xor (inputs(209)));
    layer0_outputs(11362) <= not(inputs(188)) or (inputs(7));
    layer0_outputs(11363) <= (inputs(117)) and not (inputs(168));
    layer0_outputs(11364) <= (inputs(58)) xor (inputs(43));
    layer0_outputs(11365) <= not(inputs(126));
    layer0_outputs(11366) <= (inputs(0)) or (inputs(199));
    layer0_outputs(11367) <= not(inputs(97)) or (inputs(5));
    layer0_outputs(11368) <= (inputs(174)) xor (inputs(133));
    layer0_outputs(11369) <= (inputs(166)) and not (inputs(21));
    layer0_outputs(11370) <= not(inputs(90));
    layer0_outputs(11371) <= not((inputs(94)) or (inputs(159)));
    layer0_outputs(11372) <= (inputs(178)) xor (inputs(206));
    layer0_outputs(11373) <= inputs(229);
    layer0_outputs(11374) <= not(inputs(109));
    layer0_outputs(11375) <= not(inputs(230)) or (inputs(143));
    layer0_outputs(11376) <= not((inputs(22)) or (inputs(64)));
    layer0_outputs(11377) <= '0';
    layer0_outputs(11378) <= (inputs(75)) and not (inputs(206));
    layer0_outputs(11379) <= not(inputs(39)) or (inputs(177));
    layer0_outputs(11380) <= not(inputs(99));
    layer0_outputs(11381) <= not((inputs(162)) or (inputs(226)));
    layer0_outputs(11382) <= not((inputs(61)) or (inputs(113)));
    layer0_outputs(11383) <= not(inputs(167));
    layer0_outputs(11384) <= (inputs(0)) or (inputs(128));
    layer0_outputs(11385) <= not((inputs(72)) xor (inputs(192)));
    layer0_outputs(11386) <= not((inputs(59)) and (inputs(186)));
    layer0_outputs(11387) <= not(inputs(188));
    layer0_outputs(11388) <= (inputs(53)) xor (inputs(8));
    layer0_outputs(11389) <= inputs(56);
    layer0_outputs(11390) <= (inputs(204)) xor (inputs(186));
    layer0_outputs(11391) <= (inputs(129)) or (inputs(135));
    layer0_outputs(11392) <= not((inputs(159)) or (inputs(152)));
    layer0_outputs(11393) <= not(inputs(89)) or (inputs(236));
    layer0_outputs(11394) <= not(inputs(229));
    layer0_outputs(11395) <= not(inputs(152)) or (inputs(229));
    layer0_outputs(11396) <= not((inputs(136)) xor (inputs(179)));
    layer0_outputs(11397) <= inputs(226);
    layer0_outputs(11398) <= not(inputs(60));
    layer0_outputs(11399) <= (inputs(171)) and not (inputs(84));
    layer0_outputs(11400) <= (inputs(235)) and not (inputs(23));
    layer0_outputs(11401) <= (inputs(179)) and not (inputs(27));
    layer0_outputs(11402) <= (inputs(87)) or (inputs(224));
    layer0_outputs(11403) <= not(inputs(20));
    layer0_outputs(11404) <= (inputs(217)) and not (inputs(45));
    layer0_outputs(11405) <= (inputs(79)) and not (inputs(144));
    layer0_outputs(11406) <= (inputs(101)) xor (inputs(81));
    layer0_outputs(11407) <= inputs(44);
    layer0_outputs(11408) <= not((inputs(149)) xor (inputs(13)));
    layer0_outputs(11409) <= not((inputs(232)) and (inputs(129)));
    layer0_outputs(11410) <= (inputs(22)) xor (inputs(5));
    layer0_outputs(11411) <= inputs(157);
    layer0_outputs(11412) <= (inputs(216)) and not (inputs(247));
    layer0_outputs(11413) <= (inputs(48)) and not (inputs(127));
    layer0_outputs(11414) <= (inputs(238)) xor (inputs(107));
    layer0_outputs(11415) <= not(inputs(77));
    layer0_outputs(11416) <= (inputs(250)) xor (inputs(87));
    layer0_outputs(11417) <= inputs(184);
    layer0_outputs(11418) <= not((inputs(60)) xor (inputs(166)));
    layer0_outputs(11419) <= (inputs(210)) and not (inputs(183));
    layer0_outputs(11420) <= not(inputs(124));
    layer0_outputs(11421) <= not(inputs(127)) or (inputs(227));
    layer0_outputs(11422) <= not((inputs(5)) xor (inputs(157)));
    layer0_outputs(11423) <= (inputs(75)) and (inputs(139));
    layer0_outputs(11424) <= (inputs(168)) and not (inputs(9));
    layer0_outputs(11425) <= (inputs(214)) and not (inputs(192));
    layer0_outputs(11426) <= not(inputs(98));
    layer0_outputs(11427) <= not(inputs(123)) or (inputs(3));
    layer0_outputs(11428) <= inputs(105);
    layer0_outputs(11429) <= inputs(190);
    layer0_outputs(11430) <= inputs(54);
    layer0_outputs(11431) <= (inputs(209)) and not (inputs(14));
    layer0_outputs(11432) <= (inputs(21)) xor (inputs(206));
    layer0_outputs(11433) <= not(inputs(138));
    layer0_outputs(11434) <= not((inputs(67)) xor (inputs(194)));
    layer0_outputs(11435) <= inputs(118);
    layer0_outputs(11436) <= '1';
    layer0_outputs(11437) <= inputs(86);
    layer0_outputs(11438) <= not((inputs(100)) xor (inputs(145)));
    layer0_outputs(11439) <= not(inputs(93));
    layer0_outputs(11440) <= not(inputs(198));
    layer0_outputs(11441) <= not(inputs(187)) or (inputs(37));
    layer0_outputs(11442) <= (inputs(162)) and not (inputs(254));
    layer0_outputs(11443) <= (inputs(120)) xor (inputs(25));
    layer0_outputs(11444) <= not(inputs(68)) or (inputs(251));
    layer0_outputs(11445) <= not(inputs(242)) or (inputs(56));
    layer0_outputs(11446) <= not((inputs(37)) xor (inputs(147)));
    layer0_outputs(11447) <= not(inputs(251));
    layer0_outputs(11448) <= (inputs(10)) and not (inputs(20));
    layer0_outputs(11449) <= not((inputs(183)) xor (inputs(105)));
    layer0_outputs(11450) <= not(inputs(199)) or (inputs(135));
    layer0_outputs(11451) <= not((inputs(77)) or (inputs(10)));
    layer0_outputs(11452) <= (inputs(204)) xor (inputs(44));
    layer0_outputs(11453) <= not(inputs(40)) or (inputs(128));
    layer0_outputs(11454) <= not((inputs(109)) or (inputs(31)));
    layer0_outputs(11455) <= (inputs(199)) xor (inputs(91));
    layer0_outputs(11456) <= (inputs(114)) and (inputs(210));
    layer0_outputs(11457) <= not((inputs(220)) xor (inputs(166)));
    layer0_outputs(11458) <= (inputs(4)) and not (inputs(250));
    layer0_outputs(11459) <= not((inputs(49)) and (inputs(190)));
    layer0_outputs(11460) <= (inputs(137)) and not (inputs(44));
    layer0_outputs(11461) <= inputs(46);
    layer0_outputs(11462) <= not((inputs(10)) or (inputs(178)));
    layer0_outputs(11463) <= (inputs(231)) or (inputs(157));
    layer0_outputs(11464) <= (inputs(221)) or (inputs(23));
    layer0_outputs(11465) <= inputs(13);
    layer0_outputs(11466) <= (inputs(185)) or (inputs(230));
    layer0_outputs(11467) <= (inputs(101)) xor (inputs(229));
    layer0_outputs(11468) <= (inputs(68)) or (inputs(23));
    layer0_outputs(11469) <= not((inputs(144)) or (inputs(203)));
    layer0_outputs(11470) <= not(inputs(192)) or (inputs(253));
    layer0_outputs(11471) <= (inputs(85)) xor (inputs(103));
    layer0_outputs(11472) <= not(inputs(182));
    layer0_outputs(11473) <= (inputs(166)) and not (inputs(102));
    layer0_outputs(11474) <= (inputs(25)) and not (inputs(213));
    layer0_outputs(11475) <= not(inputs(226)) or (inputs(245));
    layer0_outputs(11476) <= inputs(177);
    layer0_outputs(11477) <= not((inputs(134)) or (inputs(224)));
    layer0_outputs(11478) <= not(inputs(167)) or (inputs(80));
    layer0_outputs(11479) <= not((inputs(12)) xor (inputs(86)));
    layer0_outputs(11480) <= (inputs(210)) xor (inputs(69));
    layer0_outputs(11481) <= not(inputs(9));
    layer0_outputs(11482) <= inputs(156);
    layer0_outputs(11483) <= not((inputs(54)) xor (inputs(226)));
    layer0_outputs(11484) <= not((inputs(224)) and (inputs(58)));
    layer0_outputs(11485) <= inputs(102);
    layer0_outputs(11486) <= (inputs(15)) and not (inputs(207));
    layer0_outputs(11487) <= not(inputs(135));
    layer0_outputs(11488) <= not(inputs(147)) or (inputs(235));
    layer0_outputs(11489) <= not(inputs(54));
    layer0_outputs(11490) <= (inputs(40)) xor (inputs(78));
    layer0_outputs(11491) <= not(inputs(140)) or (inputs(35));
    layer0_outputs(11492) <= not(inputs(19)) or (inputs(162));
    layer0_outputs(11493) <= (inputs(5)) and not (inputs(248));
    layer0_outputs(11494) <= not(inputs(86)) or (inputs(43));
    layer0_outputs(11495) <= (inputs(201)) xor (inputs(147));
    layer0_outputs(11496) <= not(inputs(96));
    layer0_outputs(11497) <= inputs(73);
    layer0_outputs(11498) <= not(inputs(215));
    layer0_outputs(11499) <= (inputs(102)) xor (inputs(108));
    layer0_outputs(11500) <= (inputs(87)) and not (inputs(148));
    layer0_outputs(11501) <= (inputs(27)) and not (inputs(63));
    layer0_outputs(11502) <= (inputs(59)) and not (inputs(22));
    layer0_outputs(11503) <= (inputs(106)) and not (inputs(25));
    layer0_outputs(11504) <= (inputs(40)) xor (inputs(127));
    layer0_outputs(11505) <= inputs(150);
    layer0_outputs(11506) <= not(inputs(170)) or (inputs(34));
    layer0_outputs(11507) <= not(inputs(153)) or (inputs(234));
    layer0_outputs(11508) <= inputs(40);
    layer0_outputs(11509) <= (inputs(184)) xor (inputs(170));
    layer0_outputs(11510) <= not(inputs(101));
    layer0_outputs(11511) <= not(inputs(228));
    layer0_outputs(11512) <= '0';
    layer0_outputs(11513) <= not(inputs(103)) or (inputs(241));
    layer0_outputs(11514) <= '0';
    layer0_outputs(11515) <= not((inputs(208)) or (inputs(111)));
    layer0_outputs(11516) <= (inputs(102)) xor (inputs(37));
    layer0_outputs(11517) <= not(inputs(163)) or (inputs(161));
    layer0_outputs(11518) <= not((inputs(246)) and (inputs(47)));
    layer0_outputs(11519) <= inputs(122);
    layer0_outputs(11520) <= (inputs(65)) and (inputs(214));
    layer0_outputs(11521) <= (inputs(205)) xor (inputs(51));
    layer0_outputs(11522) <= inputs(148);
    layer0_outputs(11523) <= (inputs(220)) and not (inputs(54));
    layer0_outputs(11524) <= not(inputs(236));
    layer0_outputs(11525) <= not(inputs(112)) or (inputs(159));
    layer0_outputs(11526) <= not((inputs(70)) or (inputs(12)));
    layer0_outputs(11527) <= (inputs(198)) xor (inputs(185));
    layer0_outputs(11528) <= (inputs(200)) and not (inputs(65));
    layer0_outputs(11529) <= not((inputs(127)) or (inputs(219)));
    layer0_outputs(11530) <= inputs(251);
    layer0_outputs(11531) <= not((inputs(146)) xor (inputs(29)));
    layer0_outputs(11532) <= (inputs(77)) and (inputs(209));
    layer0_outputs(11533) <= inputs(63);
    layer0_outputs(11534) <= not((inputs(144)) xor (inputs(181)));
    layer0_outputs(11535) <= (inputs(23)) xor (inputs(172));
    layer0_outputs(11536) <= not((inputs(29)) xor (inputs(124)));
    layer0_outputs(11537) <= (inputs(17)) xor (inputs(102));
    layer0_outputs(11538) <= not((inputs(220)) or (inputs(86)));
    layer0_outputs(11539) <= not((inputs(103)) or (inputs(186)));
    layer0_outputs(11540) <= (inputs(18)) xor (inputs(157));
    layer0_outputs(11541) <= (inputs(65)) and not (inputs(227));
    layer0_outputs(11542) <= (inputs(223)) and (inputs(9));
    layer0_outputs(11543) <= (inputs(189)) or (inputs(130));
    layer0_outputs(11544) <= not(inputs(234));
    layer0_outputs(11545) <= not((inputs(94)) xor (inputs(254)));
    layer0_outputs(11546) <= inputs(151);
    layer0_outputs(11547) <= (inputs(221)) and not (inputs(67));
    layer0_outputs(11548) <= not(inputs(113)) or (inputs(130));
    layer0_outputs(11549) <= not(inputs(202)) or (inputs(62));
    layer0_outputs(11550) <= not((inputs(166)) xor (inputs(135)));
    layer0_outputs(11551) <= not(inputs(32)) or (inputs(68));
    layer0_outputs(11552) <= (inputs(66)) and (inputs(3));
    layer0_outputs(11553) <= (inputs(105)) and not (inputs(247));
    layer0_outputs(11554) <= not((inputs(126)) or (inputs(219)));
    layer0_outputs(11555) <= (inputs(227)) and not (inputs(157));
    layer0_outputs(11556) <= (inputs(56)) xor (inputs(236));
    layer0_outputs(11557) <= not(inputs(107));
    layer0_outputs(11558) <= not(inputs(37));
    layer0_outputs(11559) <= (inputs(124)) or (inputs(46));
    layer0_outputs(11560) <= '1';
    layer0_outputs(11561) <= '0';
    layer0_outputs(11562) <= not((inputs(218)) xor (inputs(76)));
    layer0_outputs(11563) <= (inputs(0)) or (inputs(135));
    layer0_outputs(11564) <= not((inputs(222)) xor (inputs(170)));
    layer0_outputs(11565) <= (inputs(39)) and not (inputs(225));
    layer0_outputs(11566) <= not((inputs(243)) xor (inputs(8)));
    layer0_outputs(11567) <= (inputs(37)) and not (inputs(33));
    layer0_outputs(11568) <= (inputs(87)) or (inputs(140));
    layer0_outputs(11569) <= (inputs(209)) or (inputs(104));
    layer0_outputs(11570) <= inputs(103);
    layer0_outputs(11571) <= (inputs(163)) and not (inputs(222));
    layer0_outputs(11572) <= not((inputs(84)) or (inputs(64)));
    layer0_outputs(11573) <= not((inputs(156)) or (inputs(63)));
    layer0_outputs(11574) <= not((inputs(212)) and (inputs(70)));
    layer0_outputs(11575) <= not((inputs(193)) xor (inputs(17)));
    layer0_outputs(11576) <= not((inputs(134)) or (inputs(61)));
    layer0_outputs(11577) <= inputs(67);
    layer0_outputs(11578) <= not((inputs(31)) or (inputs(12)));
    layer0_outputs(11579) <= inputs(148);
    layer0_outputs(11580) <= not(inputs(214));
    layer0_outputs(11581) <= not(inputs(138));
    layer0_outputs(11582) <= inputs(86);
    layer0_outputs(11583) <= not((inputs(215)) or (inputs(197)));
    layer0_outputs(11584) <= (inputs(6)) xor (inputs(147));
    layer0_outputs(11585) <= (inputs(77)) or (inputs(179));
    layer0_outputs(11586) <= (inputs(150)) xor (inputs(15));
    layer0_outputs(11587) <= not((inputs(213)) or (inputs(39)));
    layer0_outputs(11588) <= not((inputs(29)) or (inputs(243)));
    layer0_outputs(11589) <= '0';
    layer0_outputs(11590) <= not((inputs(119)) xor (inputs(133)));
    layer0_outputs(11591) <= not((inputs(186)) xor (inputs(90)));
    layer0_outputs(11592) <= not((inputs(21)) xor (inputs(72)));
    layer0_outputs(11593) <= not(inputs(112)) or (inputs(189));
    layer0_outputs(11594) <= (inputs(155)) xor (inputs(95));
    layer0_outputs(11595) <= not((inputs(238)) or (inputs(27)));
    layer0_outputs(11596) <= inputs(5);
    layer0_outputs(11597) <= not(inputs(67)) or (inputs(113));
    layer0_outputs(11598) <= (inputs(198)) xor (inputs(234));
    layer0_outputs(11599) <= inputs(215);
    layer0_outputs(11600) <= inputs(102);
    layer0_outputs(11601) <= (inputs(133)) xor (inputs(74));
    layer0_outputs(11602) <= not((inputs(86)) or (inputs(115)));
    layer0_outputs(11603) <= not((inputs(127)) and (inputs(177)));
    layer0_outputs(11604) <= not((inputs(133)) or (inputs(213)));
    layer0_outputs(11605) <= '1';
    layer0_outputs(11606) <= not(inputs(229));
    layer0_outputs(11607) <= not((inputs(130)) and (inputs(35)));
    layer0_outputs(11608) <= not(inputs(31));
    layer0_outputs(11609) <= not(inputs(131));
    layer0_outputs(11610) <= inputs(63);
    layer0_outputs(11611) <= (inputs(183)) and not (inputs(248));
    layer0_outputs(11612) <= not((inputs(182)) or (inputs(196)));
    layer0_outputs(11613) <= not(inputs(231));
    layer0_outputs(11614) <= not(inputs(20));
    layer0_outputs(11615) <= not((inputs(57)) and (inputs(226)));
    layer0_outputs(11616) <= not((inputs(46)) xor (inputs(235)));
    layer0_outputs(11617) <= not((inputs(177)) xor (inputs(240)));
    layer0_outputs(11618) <= (inputs(87)) and not (inputs(12));
    layer0_outputs(11619) <= (inputs(92)) and not (inputs(194));
    layer0_outputs(11620) <= not((inputs(6)) and (inputs(218)));
    layer0_outputs(11621) <= not((inputs(183)) or (inputs(200)));
    layer0_outputs(11622) <= not(inputs(89)) or (inputs(142));
    layer0_outputs(11623) <= not((inputs(68)) xor (inputs(115)));
    layer0_outputs(11624) <= not(inputs(229));
    layer0_outputs(11625) <= inputs(104);
    layer0_outputs(11626) <= (inputs(159)) and not (inputs(237));
    layer0_outputs(11627) <= '0';
    layer0_outputs(11628) <= not((inputs(150)) or (inputs(125)));
    layer0_outputs(11629) <= inputs(141);
    layer0_outputs(11630) <= not((inputs(126)) xor (inputs(170)));
    layer0_outputs(11631) <= not((inputs(48)) xor (inputs(8)));
    layer0_outputs(11632) <= inputs(225);
    layer0_outputs(11633) <= not((inputs(186)) or (inputs(79)));
    layer0_outputs(11634) <= not(inputs(86)) or (inputs(160));
    layer0_outputs(11635) <= (inputs(116)) and not (inputs(191));
    layer0_outputs(11636) <= inputs(45);
    layer0_outputs(11637) <= not(inputs(204)) or (inputs(115));
    layer0_outputs(11638) <= '1';
    layer0_outputs(11639) <= inputs(70);
    layer0_outputs(11640) <= (inputs(218)) xor (inputs(59));
    layer0_outputs(11641) <= not(inputs(121));
    layer0_outputs(11642) <= not((inputs(132)) xor (inputs(1)));
    layer0_outputs(11643) <= not(inputs(223)) or (inputs(255));
    layer0_outputs(11644) <= inputs(69);
    layer0_outputs(11645) <= not(inputs(38));
    layer0_outputs(11646) <= (inputs(87)) and not (inputs(106));
    layer0_outputs(11647) <= not(inputs(93)) or (inputs(30));
    layer0_outputs(11648) <= not((inputs(238)) or (inputs(61)));
    layer0_outputs(11649) <= not((inputs(239)) xor (inputs(53)));
    layer0_outputs(11650) <= not((inputs(3)) or (inputs(132)));
    layer0_outputs(11651) <= (inputs(71)) or (inputs(21));
    layer0_outputs(11652) <= not((inputs(42)) xor (inputs(88)));
    layer0_outputs(11653) <= inputs(11);
    layer0_outputs(11654) <= (inputs(139)) xor (inputs(216));
    layer0_outputs(11655) <= inputs(168);
    layer0_outputs(11656) <= not(inputs(1)) or (inputs(225));
    layer0_outputs(11657) <= (inputs(210)) and not (inputs(3));
    layer0_outputs(11658) <= (inputs(57)) xor (inputs(225));
    layer0_outputs(11659) <= (inputs(128)) xor (inputs(68));
    layer0_outputs(11660) <= (inputs(158)) xor (inputs(131));
    layer0_outputs(11661) <= not(inputs(165)) or (inputs(207));
    layer0_outputs(11662) <= inputs(117);
    layer0_outputs(11663) <= not((inputs(113)) xor (inputs(245)));
    layer0_outputs(11664) <= (inputs(181)) and not (inputs(138));
    layer0_outputs(11665) <= inputs(118);
    layer0_outputs(11666) <= not(inputs(254));
    layer0_outputs(11667) <= (inputs(222)) xor (inputs(99));
    layer0_outputs(11668) <= not(inputs(95));
    layer0_outputs(11669) <= (inputs(215)) or (inputs(208));
    layer0_outputs(11670) <= (inputs(87)) and not (inputs(23));
    layer0_outputs(11671) <= not(inputs(87)) or (inputs(35));
    layer0_outputs(11672) <= not((inputs(158)) xor (inputs(74)));
    layer0_outputs(11673) <= (inputs(7)) and (inputs(15));
    layer0_outputs(11674) <= (inputs(156)) and not (inputs(251));
    layer0_outputs(11675) <= (inputs(121)) and not (inputs(173));
    layer0_outputs(11676) <= not((inputs(66)) or (inputs(167)));
    layer0_outputs(11677) <= not(inputs(219)) or (inputs(246));
    layer0_outputs(11678) <= (inputs(125)) and (inputs(142));
    layer0_outputs(11679) <= (inputs(173)) xor (inputs(37));
    layer0_outputs(11680) <= not(inputs(26));
    layer0_outputs(11681) <= not(inputs(56));
    layer0_outputs(11682) <= (inputs(150)) and not (inputs(112));
    layer0_outputs(11683) <= (inputs(144)) and not (inputs(123));
    layer0_outputs(11684) <= not(inputs(199)) or (inputs(107));
    layer0_outputs(11685) <= not(inputs(199));
    layer0_outputs(11686) <= inputs(119);
    layer0_outputs(11687) <= not((inputs(103)) or (inputs(113)));
    layer0_outputs(11688) <= (inputs(83)) and not (inputs(16));
    layer0_outputs(11689) <= not(inputs(218));
    layer0_outputs(11690) <= (inputs(111)) xor (inputs(181));
    layer0_outputs(11691) <= (inputs(21)) xor (inputs(120));
    layer0_outputs(11692) <= (inputs(152)) or (inputs(145));
    layer0_outputs(11693) <= not((inputs(234)) xor (inputs(220)));
    layer0_outputs(11694) <= (inputs(140)) or (inputs(230));
    layer0_outputs(11695) <= not(inputs(25)) or (inputs(3));
    layer0_outputs(11696) <= not((inputs(124)) or (inputs(137)));
    layer0_outputs(11697) <= (inputs(109)) and not (inputs(177));
    layer0_outputs(11698) <= not(inputs(107));
    layer0_outputs(11699) <= '1';
    layer0_outputs(11700) <= not((inputs(66)) xor (inputs(172)));
    layer0_outputs(11701) <= (inputs(152)) and not (inputs(72));
    layer0_outputs(11702) <= '0';
    layer0_outputs(11703) <= inputs(84);
    layer0_outputs(11704) <= not(inputs(81)) or (inputs(50));
    layer0_outputs(11705) <= not((inputs(62)) or (inputs(196)));
    layer0_outputs(11706) <= not(inputs(188)) or (inputs(20));
    layer0_outputs(11707) <= not((inputs(17)) xor (inputs(39)));
    layer0_outputs(11708) <= not((inputs(37)) xor (inputs(188)));
    layer0_outputs(11709) <= not((inputs(55)) or (inputs(20)));
    layer0_outputs(11710) <= inputs(126);
    layer0_outputs(11711) <= inputs(239);
    layer0_outputs(11712) <= not((inputs(239)) and (inputs(62)));
    layer0_outputs(11713) <= inputs(175);
    layer0_outputs(11714) <= (inputs(120)) or (inputs(76));
    layer0_outputs(11715) <= not((inputs(97)) xor (inputs(163)));
    layer0_outputs(11716) <= not(inputs(18));
    layer0_outputs(11717) <= not(inputs(156)) or (inputs(142));
    layer0_outputs(11718) <= not(inputs(198)) or (inputs(153));
    layer0_outputs(11719) <= (inputs(100)) or (inputs(120));
    layer0_outputs(11720) <= not(inputs(203));
    layer0_outputs(11721) <= not((inputs(78)) xor (inputs(90)));
    layer0_outputs(11722) <= (inputs(104)) and not (inputs(21));
    layer0_outputs(11723) <= not(inputs(165));
    layer0_outputs(11724) <= (inputs(184)) and not (inputs(65));
    layer0_outputs(11725) <= not(inputs(205));
    layer0_outputs(11726) <= not((inputs(240)) or (inputs(124)));
    layer0_outputs(11727) <= not((inputs(254)) xor (inputs(121)));
    layer0_outputs(11728) <= (inputs(136)) and not (inputs(194));
    layer0_outputs(11729) <= (inputs(175)) and (inputs(170));
    layer0_outputs(11730) <= not((inputs(8)) or (inputs(212)));
    layer0_outputs(11731) <= (inputs(201)) or (inputs(129));
    layer0_outputs(11732) <= not((inputs(201)) or (inputs(141)));
    layer0_outputs(11733) <= (inputs(108)) and not (inputs(20));
    layer0_outputs(11734) <= not(inputs(210)) or (inputs(20));
    layer0_outputs(11735) <= (inputs(57)) or (inputs(242));
    layer0_outputs(11736) <= not(inputs(20)) or (inputs(69));
    layer0_outputs(11737) <= not((inputs(128)) or (inputs(245)));
    layer0_outputs(11738) <= (inputs(35)) or (inputs(69));
    layer0_outputs(11739) <= (inputs(12)) or (inputs(35));
    layer0_outputs(11740) <= inputs(234);
    layer0_outputs(11741) <= '1';
    layer0_outputs(11742) <= not((inputs(77)) or (inputs(215)));
    layer0_outputs(11743) <= (inputs(37)) xor (inputs(99));
    layer0_outputs(11744) <= not(inputs(208)) or (inputs(178));
    layer0_outputs(11745) <= not((inputs(64)) xor (inputs(140)));
    layer0_outputs(11746) <= (inputs(120)) and not (inputs(48));
    layer0_outputs(11747) <= (inputs(8)) xor (inputs(64));
    layer0_outputs(11748) <= inputs(60);
    layer0_outputs(11749) <= not(inputs(134));
    layer0_outputs(11750) <= not((inputs(215)) and (inputs(88)));
    layer0_outputs(11751) <= not(inputs(54)) or (inputs(99));
    layer0_outputs(11752) <= not(inputs(69));
    layer0_outputs(11753) <= inputs(71);
    layer0_outputs(11754) <= inputs(16);
    layer0_outputs(11755) <= (inputs(39)) or (inputs(29));
    layer0_outputs(11756) <= (inputs(15)) and not (inputs(170));
    layer0_outputs(11757) <= not(inputs(158)) or (inputs(233));
    layer0_outputs(11758) <= not(inputs(116));
    layer0_outputs(11759) <= (inputs(44)) or (inputs(27));
    layer0_outputs(11760) <= not((inputs(90)) or (inputs(51)));
    layer0_outputs(11761) <= (inputs(187)) and not (inputs(236));
    layer0_outputs(11762) <= (inputs(255)) xor (inputs(57));
    layer0_outputs(11763) <= (inputs(92)) and not (inputs(122));
    layer0_outputs(11764) <= inputs(200);
    layer0_outputs(11765) <= not((inputs(60)) xor (inputs(19)));
    layer0_outputs(11766) <= (inputs(50)) xor (inputs(169));
    layer0_outputs(11767) <= not((inputs(81)) or (inputs(213)));
    layer0_outputs(11768) <= (inputs(137)) xor (inputs(186));
    layer0_outputs(11769) <= (inputs(242)) or (inputs(80));
    layer0_outputs(11770) <= inputs(16);
    layer0_outputs(11771) <= (inputs(37)) xor (inputs(205));
    layer0_outputs(11772) <= not(inputs(200));
    layer0_outputs(11773) <= (inputs(42)) and not (inputs(21));
    layer0_outputs(11774) <= (inputs(200)) xor (inputs(216));
    layer0_outputs(11775) <= (inputs(78)) or (inputs(167));
    layer0_outputs(11776) <= (inputs(224)) xor (inputs(155));
    layer0_outputs(11777) <= inputs(205);
    layer0_outputs(11778) <= not(inputs(143));
    layer0_outputs(11779) <= (inputs(116)) xor (inputs(117));
    layer0_outputs(11780) <= (inputs(150)) or (inputs(96));
    layer0_outputs(11781) <= (inputs(47)) xor (inputs(10));
    layer0_outputs(11782) <= not((inputs(92)) or (inputs(207)));
    layer0_outputs(11783) <= '1';
    layer0_outputs(11784) <= not(inputs(237)) or (inputs(232));
    layer0_outputs(11785) <= (inputs(246)) and not (inputs(247));
    layer0_outputs(11786) <= not(inputs(131));
    layer0_outputs(11787) <= not(inputs(250));
    layer0_outputs(11788) <= not(inputs(155));
    layer0_outputs(11789) <= not(inputs(40));
    layer0_outputs(11790) <= (inputs(225)) and not (inputs(95));
    layer0_outputs(11791) <= (inputs(195)) xor (inputs(75));
    layer0_outputs(11792) <= not((inputs(60)) xor (inputs(74)));
    layer0_outputs(11793) <= (inputs(48)) or (inputs(87));
    layer0_outputs(11794) <= '1';
    layer0_outputs(11795) <= (inputs(139)) xor (inputs(230));
    layer0_outputs(11796) <= (inputs(93)) or (inputs(230));
    layer0_outputs(11797) <= not(inputs(11)) or (inputs(58));
    layer0_outputs(11798) <= not(inputs(39));
    layer0_outputs(11799) <= (inputs(154)) and not (inputs(125));
    layer0_outputs(11800) <= inputs(253);
    layer0_outputs(11801) <= not((inputs(176)) xor (inputs(224)));
    layer0_outputs(11802) <= inputs(228);
    layer0_outputs(11803) <= (inputs(224)) xor (inputs(49));
    layer0_outputs(11804) <= not(inputs(186));
    layer0_outputs(11805) <= not(inputs(6)) or (inputs(142));
    layer0_outputs(11806) <= not(inputs(220)) or (inputs(212));
    layer0_outputs(11807) <= not(inputs(163));
    layer0_outputs(11808) <= (inputs(82)) and (inputs(220));
    layer0_outputs(11809) <= (inputs(178)) and not (inputs(35));
    layer0_outputs(11810) <= (inputs(85)) xor (inputs(31));
    layer0_outputs(11811) <= (inputs(75)) xor (inputs(69));
    layer0_outputs(11812) <= not((inputs(114)) or (inputs(129)));
    layer0_outputs(11813) <= not((inputs(249)) xor (inputs(148)));
    layer0_outputs(11814) <= (inputs(49)) xor (inputs(206));
    layer0_outputs(11815) <= inputs(146);
    layer0_outputs(11816) <= not((inputs(181)) xor (inputs(161)));
    layer0_outputs(11817) <= not(inputs(201)) or (inputs(252));
    layer0_outputs(11818) <= not(inputs(49));
    layer0_outputs(11819) <= not(inputs(214));
    layer0_outputs(11820) <= not(inputs(158)) or (inputs(243));
    layer0_outputs(11821) <= (inputs(4)) or (inputs(101));
    layer0_outputs(11822) <= not(inputs(147));
    layer0_outputs(11823) <= inputs(182);
    layer0_outputs(11824) <= not(inputs(112)) or (inputs(128));
    layer0_outputs(11825) <= (inputs(31)) or (inputs(195));
    layer0_outputs(11826) <= inputs(107);
    layer0_outputs(11827) <= (inputs(108)) or (inputs(87));
    layer0_outputs(11828) <= not(inputs(102)) or (inputs(254));
    layer0_outputs(11829) <= (inputs(5)) and not (inputs(190));
    layer0_outputs(11830) <= (inputs(155)) xor (inputs(163));
    layer0_outputs(11831) <= '1';
    layer0_outputs(11832) <= not(inputs(115)) or (inputs(48));
    layer0_outputs(11833) <= (inputs(129)) xor (inputs(102));
    layer0_outputs(11834) <= not((inputs(148)) or (inputs(85)));
    layer0_outputs(11835) <= (inputs(175)) and not (inputs(15));
    layer0_outputs(11836) <= (inputs(196)) and not (inputs(220));
    layer0_outputs(11837) <= (inputs(253)) or (inputs(33));
    layer0_outputs(11838) <= (inputs(57)) or (inputs(124));
    layer0_outputs(11839) <= not((inputs(150)) or (inputs(95)));
    layer0_outputs(11840) <= inputs(252);
    layer0_outputs(11841) <= '1';
    layer0_outputs(11842) <= not(inputs(38)) or (inputs(247));
    layer0_outputs(11843) <= not((inputs(195)) xor (inputs(169)));
    layer0_outputs(11844) <= not((inputs(208)) and (inputs(47)));
    layer0_outputs(11845) <= not((inputs(40)) or (inputs(54)));
    layer0_outputs(11846) <= inputs(17);
    layer0_outputs(11847) <= (inputs(33)) xor (inputs(174));
    layer0_outputs(11848) <= inputs(79);
    layer0_outputs(11849) <= (inputs(90)) xor (inputs(208));
    layer0_outputs(11850) <= not(inputs(45));
    layer0_outputs(11851) <= not((inputs(41)) xor (inputs(162)));
    layer0_outputs(11852) <= (inputs(172)) or (inputs(58));
    layer0_outputs(11853) <= not(inputs(84)) or (inputs(227));
    layer0_outputs(11854) <= not(inputs(86)) or (inputs(29));
    layer0_outputs(11855) <= '1';
    layer0_outputs(11856) <= (inputs(234)) and not (inputs(116));
    layer0_outputs(11857) <= (inputs(157)) and not (inputs(226));
    layer0_outputs(11858) <= (inputs(216)) and not (inputs(33));
    layer0_outputs(11859) <= not(inputs(132)) or (inputs(136));
    layer0_outputs(11860) <= not(inputs(89)) or (inputs(160));
    layer0_outputs(11861) <= (inputs(194)) or (inputs(220));
    layer0_outputs(11862) <= not(inputs(196));
    layer0_outputs(11863) <= not(inputs(132));
    layer0_outputs(11864) <= not(inputs(217));
    layer0_outputs(11865) <= not((inputs(247)) or (inputs(216)));
    layer0_outputs(11866) <= not((inputs(1)) or (inputs(113)));
    layer0_outputs(11867) <= inputs(150);
    layer0_outputs(11868) <= (inputs(200)) and not (inputs(129));
    layer0_outputs(11869) <= not(inputs(46)) or (inputs(35));
    layer0_outputs(11870) <= (inputs(94)) or (inputs(97));
    layer0_outputs(11871) <= not(inputs(250));
    layer0_outputs(11872) <= not((inputs(101)) xor (inputs(112)));
    layer0_outputs(11873) <= (inputs(192)) and not (inputs(239));
    layer0_outputs(11874) <= not(inputs(104)) or (inputs(203));
    layer0_outputs(11875) <= (inputs(240)) xor (inputs(73));
    layer0_outputs(11876) <= not((inputs(63)) xor (inputs(231)));
    layer0_outputs(11877) <= (inputs(38)) xor (inputs(53));
    layer0_outputs(11878) <= not((inputs(54)) or (inputs(58)));
    layer0_outputs(11879) <= (inputs(119)) and not (inputs(14));
    layer0_outputs(11880) <= (inputs(252)) and not (inputs(242));
    layer0_outputs(11881) <= not(inputs(116));
    layer0_outputs(11882) <= not(inputs(48));
    layer0_outputs(11883) <= (inputs(193)) xor (inputs(40));
    layer0_outputs(11884) <= not((inputs(207)) xor (inputs(124)));
    layer0_outputs(11885) <= inputs(128);
    layer0_outputs(11886) <= not(inputs(92));
    layer0_outputs(11887) <= (inputs(166)) xor (inputs(44));
    layer0_outputs(11888) <= not(inputs(228)) or (inputs(209));
    layer0_outputs(11889) <= not(inputs(105));
    layer0_outputs(11890) <= (inputs(88)) and (inputs(170));
    layer0_outputs(11891) <= not(inputs(164));
    layer0_outputs(11892) <= not(inputs(83)) or (inputs(2));
    layer0_outputs(11893) <= not(inputs(107));
    layer0_outputs(11894) <= not(inputs(21));
    layer0_outputs(11895) <= (inputs(23)) or (inputs(50));
    layer0_outputs(11896) <= not((inputs(221)) xor (inputs(230)));
    layer0_outputs(11897) <= not(inputs(90));
    layer0_outputs(11898) <= not((inputs(182)) or (inputs(131)));
    layer0_outputs(11899) <= not((inputs(138)) xor (inputs(229)));
    layer0_outputs(11900) <= inputs(123);
    layer0_outputs(11901) <= (inputs(205)) or (inputs(77));
    layer0_outputs(11902) <= inputs(22);
    layer0_outputs(11903) <= not((inputs(250)) xor (inputs(39)));
    layer0_outputs(11904) <= not(inputs(60));
    layer0_outputs(11905) <= not((inputs(217)) or (inputs(124)));
    layer0_outputs(11906) <= not(inputs(150));
    layer0_outputs(11907) <= (inputs(200)) xor (inputs(109));
    layer0_outputs(11908) <= (inputs(147)) xor (inputs(193));
    layer0_outputs(11909) <= not((inputs(69)) and (inputs(104)));
    layer0_outputs(11910) <= (inputs(231)) and (inputs(94));
    layer0_outputs(11911) <= not(inputs(146));
    layer0_outputs(11912) <= not((inputs(24)) or (inputs(152)));
    layer0_outputs(11913) <= inputs(152);
    layer0_outputs(11914) <= (inputs(198)) and (inputs(166));
    layer0_outputs(11915) <= (inputs(207)) and not (inputs(127));
    layer0_outputs(11916) <= (inputs(31)) and not (inputs(244));
    layer0_outputs(11917) <= inputs(118);
    layer0_outputs(11918) <= '0';
    layer0_outputs(11919) <= inputs(178);
    layer0_outputs(11920) <= inputs(156);
    layer0_outputs(11921) <= inputs(98);
    layer0_outputs(11922) <= not((inputs(91)) xor (inputs(95)));
    layer0_outputs(11923) <= (inputs(10)) and not (inputs(244));
    layer0_outputs(11924) <= not(inputs(191));
    layer0_outputs(11925) <= not((inputs(159)) xor (inputs(34)));
    layer0_outputs(11926) <= not(inputs(110)) or (inputs(244));
    layer0_outputs(11927) <= (inputs(173)) xor (inputs(50));
    layer0_outputs(11928) <= (inputs(209)) xor (inputs(72));
    layer0_outputs(11929) <= not(inputs(126)) or (inputs(227));
    layer0_outputs(11930) <= not((inputs(238)) or (inputs(199)));
    layer0_outputs(11931) <= inputs(115);
    layer0_outputs(11932) <= not((inputs(54)) xor (inputs(147)));
    layer0_outputs(11933) <= '1';
    layer0_outputs(11934) <= not(inputs(79)) or (inputs(16));
    layer0_outputs(11935) <= inputs(33);
    layer0_outputs(11936) <= not(inputs(220));
    layer0_outputs(11937) <= (inputs(223)) xor (inputs(221));
    layer0_outputs(11938) <= (inputs(80)) and (inputs(183));
    layer0_outputs(11939) <= '0';
    layer0_outputs(11940) <= (inputs(97)) and not (inputs(123));
    layer0_outputs(11941) <= (inputs(59)) or (inputs(221));
    layer0_outputs(11942) <= not((inputs(248)) xor (inputs(233)));
    layer0_outputs(11943) <= (inputs(112)) or (inputs(235));
    layer0_outputs(11944) <= inputs(180);
    layer0_outputs(11945) <= not((inputs(123)) xor (inputs(60)));
    layer0_outputs(11946) <= not(inputs(53));
    layer0_outputs(11947) <= not(inputs(41)) or (inputs(63));
    layer0_outputs(11948) <= (inputs(32)) and not (inputs(112));
    layer0_outputs(11949) <= not((inputs(57)) xor (inputs(119)));
    layer0_outputs(11950) <= (inputs(165)) or (inputs(128));
    layer0_outputs(11951) <= not((inputs(43)) or (inputs(27)));
    layer0_outputs(11952) <= '1';
    layer0_outputs(11953) <= not((inputs(146)) xor (inputs(126)));
    layer0_outputs(11954) <= (inputs(83)) and not (inputs(227));
    layer0_outputs(11955) <= inputs(118);
    layer0_outputs(11956) <= '0';
    layer0_outputs(11957) <= not(inputs(181));
    layer0_outputs(11958) <= inputs(58);
    layer0_outputs(11959) <= (inputs(231)) xor (inputs(169));
    layer0_outputs(11960) <= (inputs(4)) or (inputs(100));
    layer0_outputs(11961) <= '1';
    layer0_outputs(11962) <= (inputs(109)) or (inputs(217));
    layer0_outputs(11963) <= not((inputs(239)) and (inputs(113)));
    layer0_outputs(11964) <= not((inputs(239)) xor (inputs(166)));
    layer0_outputs(11965) <= '1';
    layer0_outputs(11966) <= (inputs(113)) and not (inputs(226));
    layer0_outputs(11967) <= (inputs(173)) xor (inputs(79));
    layer0_outputs(11968) <= (inputs(246)) xor (inputs(57));
    layer0_outputs(11969) <= not(inputs(155));
    layer0_outputs(11970) <= not(inputs(137));
    layer0_outputs(11971) <= not((inputs(232)) or (inputs(196)));
    layer0_outputs(11972) <= (inputs(247)) xor (inputs(124));
    layer0_outputs(11973) <= (inputs(205)) or (inputs(152));
    layer0_outputs(11974) <= (inputs(247)) xor (inputs(47));
    layer0_outputs(11975) <= not((inputs(240)) or (inputs(215)));
    layer0_outputs(11976) <= not(inputs(91)) or (inputs(218));
    layer0_outputs(11977) <= (inputs(197)) and not (inputs(98));
    layer0_outputs(11978) <= (inputs(111)) or (inputs(154));
    layer0_outputs(11979) <= not((inputs(230)) or (inputs(236)));
    layer0_outputs(11980) <= inputs(141);
    layer0_outputs(11981) <= (inputs(140)) xor (inputs(144));
    layer0_outputs(11982) <= (inputs(55)) or (inputs(99));
    layer0_outputs(11983) <= not(inputs(108));
    layer0_outputs(11984) <= (inputs(45)) or (inputs(95));
    layer0_outputs(11985) <= not(inputs(161));
    layer0_outputs(11986) <= not((inputs(123)) or (inputs(106)));
    layer0_outputs(11987) <= '1';
    layer0_outputs(11988) <= (inputs(14)) or (inputs(206));
    layer0_outputs(11989) <= not(inputs(156));
    layer0_outputs(11990) <= not(inputs(135));
    layer0_outputs(11991) <= not((inputs(115)) or (inputs(28)));
    layer0_outputs(11992) <= not((inputs(252)) and (inputs(113)));
    layer0_outputs(11993) <= not((inputs(44)) xor (inputs(186)));
    layer0_outputs(11994) <= inputs(117);
    layer0_outputs(11995) <= not(inputs(154));
    layer0_outputs(11996) <= (inputs(118)) xor (inputs(21));
    layer0_outputs(11997) <= (inputs(154)) or (inputs(226));
    layer0_outputs(11998) <= inputs(230);
    layer0_outputs(11999) <= (inputs(60)) and (inputs(229));
    layer0_outputs(12000) <= (inputs(224)) xor (inputs(243));
    layer0_outputs(12001) <= (inputs(131)) or (inputs(244));
    layer0_outputs(12002) <= (inputs(76)) xor (inputs(59));
    layer0_outputs(12003) <= not(inputs(197)) or (inputs(77));
    layer0_outputs(12004) <= not(inputs(127)) or (inputs(28));
    layer0_outputs(12005) <= (inputs(17)) xor (inputs(77));
    layer0_outputs(12006) <= inputs(96);
    layer0_outputs(12007) <= not((inputs(215)) xor (inputs(239)));
    layer0_outputs(12008) <= inputs(3);
    layer0_outputs(12009) <= (inputs(208)) and not (inputs(172));
    layer0_outputs(12010) <= (inputs(218)) and not (inputs(125));
    layer0_outputs(12011) <= (inputs(182)) and (inputs(243));
    layer0_outputs(12012) <= not((inputs(252)) or (inputs(134)));
    layer0_outputs(12013) <= not((inputs(8)) or (inputs(166)));
    layer0_outputs(12014) <= (inputs(246)) or (inputs(197));
    layer0_outputs(12015) <= inputs(168);
    layer0_outputs(12016) <= inputs(167);
    layer0_outputs(12017) <= (inputs(138)) and not (inputs(58));
    layer0_outputs(12018) <= not((inputs(88)) or (inputs(194)));
    layer0_outputs(12019) <= not(inputs(167));
    layer0_outputs(12020) <= not(inputs(21));
    layer0_outputs(12021) <= inputs(207);
    layer0_outputs(12022) <= not(inputs(226));
    layer0_outputs(12023) <= not(inputs(77));
    layer0_outputs(12024) <= not((inputs(171)) or (inputs(0)));
    layer0_outputs(12025) <= inputs(103);
    layer0_outputs(12026) <= not((inputs(210)) xor (inputs(7)));
    layer0_outputs(12027) <= (inputs(107)) and not (inputs(161));
    layer0_outputs(12028) <= (inputs(213)) xor (inputs(199));
    layer0_outputs(12029) <= (inputs(112)) and (inputs(207));
    layer0_outputs(12030) <= not((inputs(163)) and (inputs(192)));
    layer0_outputs(12031) <= (inputs(102)) xor (inputs(99));
    layer0_outputs(12032) <= (inputs(140)) xor (inputs(172));
    layer0_outputs(12033) <= not((inputs(249)) or (inputs(153)));
    layer0_outputs(12034) <= not(inputs(33)) or (inputs(187));
    layer0_outputs(12035) <= not((inputs(232)) xor (inputs(26)));
    layer0_outputs(12036) <= inputs(243);
    layer0_outputs(12037) <= (inputs(52)) or (inputs(175));
    layer0_outputs(12038) <= (inputs(131)) xor (inputs(156));
    layer0_outputs(12039) <= (inputs(97)) xor (inputs(95));
    layer0_outputs(12040) <= (inputs(102)) xor (inputs(52));
    layer0_outputs(12041) <= (inputs(154)) and (inputs(190));
    layer0_outputs(12042) <= (inputs(183)) and not (inputs(81));
    layer0_outputs(12043) <= '0';
    layer0_outputs(12044) <= inputs(4);
    layer0_outputs(12045) <= not(inputs(82));
    layer0_outputs(12046) <= (inputs(109)) xor (inputs(205));
    layer0_outputs(12047) <= (inputs(71)) xor (inputs(0));
    layer0_outputs(12048) <= not((inputs(96)) xor (inputs(104)));
    layer0_outputs(12049) <= not((inputs(27)) and (inputs(76)));
    layer0_outputs(12050) <= not((inputs(17)) or (inputs(58)));
    layer0_outputs(12051) <= (inputs(210)) or (inputs(35));
    layer0_outputs(12052) <= not((inputs(20)) or (inputs(8)));
    layer0_outputs(12053) <= inputs(142);
    layer0_outputs(12054) <= '1';
    layer0_outputs(12055) <= (inputs(171)) xor (inputs(112));
    layer0_outputs(12056) <= (inputs(208)) xor (inputs(82));
    layer0_outputs(12057) <= not((inputs(59)) and (inputs(156)));
    layer0_outputs(12058) <= not((inputs(140)) xor (inputs(129)));
    layer0_outputs(12059) <= not(inputs(113)) or (inputs(31));
    layer0_outputs(12060) <= inputs(139);
    layer0_outputs(12061) <= not(inputs(79));
    layer0_outputs(12062) <= (inputs(253)) or (inputs(173));
    layer0_outputs(12063) <= not(inputs(45)) or (inputs(68));
    layer0_outputs(12064) <= not((inputs(220)) xor (inputs(189)));
    layer0_outputs(12065) <= (inputs(162)) xor (inputs(119));
    layer0_outputs(12066) <= (inputs(155)) xor (inputs(156));
    layer0_outputs(12067) <= (inputs(60)) or (inputs(180));
    layer0_outputs(12068) <= not((inputs(180)) xor (inputs(73)));
    layer0_outputs(12069) <= not((inputs(96)) xor (inputs(19)));
    layer0_outputs(12070) <= (inputs(197)) and not (inputs(114));
    layer0_outputs(12071) <= (inputs(161)) xor (inputs(188));
    layer0_outputs(12072) <= not((inputs(105)) xor (inputs(92)));
    layer0_outputs(12073) <= inputs(220);
    layer0_outputs(12074) <= not((inputs(104)) xor (inputs(250)));
    layer0_outputs(12075) <= (inputs(85)) and not (inputs(113));
    layer0_outputs(12076) <= not(inputs(115));
    layer0_outputs(12077) <= inputs(162);
    layer0_outputs(12078) <= (inputs(223)) or (inputs(111));
    layer0_outputs(12079) <= not((inputs(206)) or (inputs(182)));
    layer0_outputs(12080) <= not(inputs(9)) or (inputs(49));
    layer0_outputs(12081) <= (inputs(200)) and not (inputs(210));
    layer0_outputs(12082) <= not(inputs(248)) or (inputs(5));
    layer0_outputs(12083) <= not((inputs(216)) or (inputs(122)));
    layer0_outputs(12084) <= (inputs(23)) xor (inputs(112));
    layer0_outputs(12085) <= not(inputs(136)) or (inputs(141));
    layer0_outputs(12086) <= not(inputs(224));
    layer0_outputs(12087) <= (inputs(161)) xor (inputs(45));
    layer0_outputs(12088) <= (inputs(36)) xor (inputs(243));
    layer0_outputs(12089) <= (inputs(216)) and not (inputs(130));
    layer0_outputs(12090) <= not(inputs(201)) or (inputs(53));
    layer0_outputs(12091) <= (inputs(186)) and not (inputs(144));
    layer0_outputs(12092) <= not(inputs(125));
    layer0_outputs(12093) <= not(inputs(235));
    layer0_outputs(12094) <= (inputs(47)) or (inputs(87));
    layer0_outputs(12095) <= not((inputs(113)) or (inputs(70)));
    layer0_outputs(12096) <= not(inputs(24)) or (inputs(221));
    layer0_outputs(12097) <= not(inputs(107));
    layer0_outputs(12098) <= not((inputs(72)) xor (inputs(177)));
    layer0_outputs(12099) <= not(inputs(218));
    layer0_outputs(12100) <= not((inputs(21)) and (inputs(253)));
    layer0_outputs(12101) <= not((inputs(218)) xor (inputs(202)));
    layer0_outputs(12102) <= inputs(229);
    layer0_outputs(12103) <= not(inputs(251));
    layer0_outputs(12104) <= not(inputs(196));
    layer0_outputs(12105) <= (inputs(95)) xor (inputs(1));
    layer0_outputs(12106) <= not(inputs(75));
    layer0_outputs(12107) <= not(inputs(116));
    layer0_outputs(12108) <= not((inputs(77)) or (inputs(170)));
    layer0_outputs(12109) <= '0';
    layer0_outputs(12110) <= not(inputs(200)) or (inputs(207));
    layer0_outputs(12111) <= not((inputs(92)) xor (inputs(61)));
    layer0_outputs(12112) <= (inputs(129)) and not (inputs(240));
    layer0_outputs(12113) <= not((inputs(164)) xor (inputs(45)));
    layer0_outputs(12114) <= inputs(168);
    layer0_outputs(12115) <= inputs(54);
    layer0_outputs(12116) <= inputs(197);
    layer0_outputs(12117) <= not((inputs(163)) or (inputs(153)));
    layer0_outputs(12118) <= (inputs(232)) or (inputs(241));
    layer0_outputs(12119) <= not(inputs(181));
    layer0_outputs(12120) <= inputs(81);
    layer0_outputs(12121) <= not((inputs(61)) or (inputs(76)));
    layer0_outputs(12122) <= (inputs(183)) or (inputs(101));
    layer0_outputs(12123) <= (inputs(160)) or (inputs(64));
    layer0_outputs(12124) <= not(inputs(40));
    layer0_outputs(12125) <= not(inputs(86));
    layer0_outputs(12126) <= not(inputs(53)) or (inputs(131));
    layer0_outputs(12127) <= not((inputs(88)) xor (inputs(132)));
    layer0_outputs(12128) <= (inputs(65)) and not (inputs(51));
    layer0_outputs(12129) <= (inputs(232)) or (inputs(118));
    layer0_outputs(12130) <= (inputs(11)) or (inputs(59));
    layer0_outputs(12131) <= not((inputs(1)) or (inputs(40)));
    layer0_outputs(12132) <= (inputs(64)) and not (inputs(211));
    layer0_outputs(12133) <= (inputs(252)) xor (inputs(209));
    layer0_outputs(12134) <= not((inputs(217)) xor (inputs(130)));
    layer0_outputs(12135) <= not((inputs(128)) or (inputs(182)));
    layer0_outputs(12136) <= (inputs(89)) or (inputs(246));
    layer0_outputs(12137) <= (inputs(118)) and not (inputs(2));
    layer0_outputs(12138) <= not((inputs(220)) or (inputs(116)));
    layer0_outputs(12139) <= (inputs(211)) or (inputs(143));
    layer0_outputs(12140) <= inputs(121);
    layer0_outputs(12141) <= not(inputs(205)) or (inputs(12));
    layer0_outputs(12142) <= not((inputs(143)) xor (inputs(237)));
    layer0_outputs(12143) <= not(inputs(84));
    layer0_outputs(12144) <= not(inputs(251)) or (inputs(32));
    layer0_outputs(12145) <= not(inputs(72)) or (inputs(51));
    layer0_outputs(12146) <= not(inputs(9));
    layer0_outputs(12147) <= not((inputs(253)) xor (inputs(214)));
    layer0_outputs(12148) <= (inputs(242)) xor (inputs(146));
    layer0_outputs(12149) <= not(inputs(57)) or (inputs(30));
    layer0_outputs(12150) <= not((inputs(47)) and (inputs(33)));
    layer0_outputs(12151) <= (inputs(16)) xor (inputs(71));
    layer0_outputs(12152) <= not(inputs(147)) or (inputs(18));
    layer0_outputs(12153) <= not((inputs(145)) xor (inputs(150)));
    layer0_outputs(12154) <= not(inputs(151));
    layer0_outputs(12155) <= not(inputs(244));
    layer0_outputs(12156) <= not(inputs(193));
    layer0_outputs(12157) <= (inputs(156)) xor (inputs(123));
    layer0_outputs(12158) <= not((inputs(146)) xor (inputs(169)));
    layer0_outputs(12159) <= not(inputs(204)) or (inputs(161));
    layer0_outputs(12160) <= (inputs(30)) xor (inputs(19));
    layer0_outputs(12161) <= not(inputs(201)) or (inputs(124));
    layer0_outputs(12162) <= (inputs(197)) and not (inputs(44));
    layer0_outputs(12163) <= inputs(160);
    layer0_outputs(12164) <= not((inputs(178)) xor (inputs(126)));
    layer0_outputs(12165) <= (inputs(171)) xor (inputs(101));
    layer0_outputs(12166) <= (inputs(135)) xor (inputs(122));
    layer0_outputs(12167) <= (inputs(149)) or (inputs(113));
    layer0_outputs(12168) <= inputs(229);
    layer0_outputs(12169) <= (inputs(56)) xor (inputs(196));
    layer0_outputs(12170) <= inputs(15);
    layer0_outputs(12171) <= not(inputs(148)) or (inputs(174));
    layer0_outputs(12172) <= (inputs(189)) and not (inputs(21));
    layer0_outputs(12173) <= not((inputs(6)) xor (inputs(100)));
    layer0_outputs(12174) <= inputs(101);
    layer0_outputs(12175) <= (inputs(130)) and not (inputs(205));
    layer0_outputs(12176) <= (inputs(194)) xor (inputs(59));
    layer0_outputs(12177) <= (inputs(156)) xor (inputs(48));
    layer0_outputs(12178) <= not((inputs(180)) or (inputs(182)));
    layer0_outputs(12179) <= not((inputs(201)) xor (inputs(185)));
    layer0_outputs(12180) <= not((inputs(242)) or (inputs(250)));
    layer0_outputs(12181) <= (inputs(176)) or (inputs(101));
    layer0_outputs(12182) <= (inputs(184)) xor (inputs(222));
    layer0_outputs(12183) <= (inputs(235)) or (inputs(90));
    layer0_outputs(12184) <= inputs(79);
    layer0_outputs(12185) <= not((inputs(14)) xor (inputs(78)));
    layer0_outputs(12186) <= (inputs(170)) and not (inputs(130));
    layer0_outputs(12187) <= '0';
    layer0_outputs(12188) <= not((inputs(17)) xor (inputs(137)));
    layer0_outputs(12189) <= not(inputs(16));
    layer0_outputs(12190) <= (inputs(239)) or (inputs(14));
    layer0_outputs(12191) <= '0';
    layer0_outputs(12192) <= not((inputs(0)) xor (inputs(74)));
    layer0_outputs(12193) <= '0';
    layer0_outputs(12194) <= (inputs(104)) and not (inputs(172));
    layer0_outputs(12195) <= '1';
    layer0_outputs(12196) <= not(inputs(5)) or (inputs(188));
    layer0_outputs(12197) <= (inputs(110)) or (inputs(103));
    layer0_outputs(12198) <= not(inputs(41));
    layer0_outputs(12199) <= (inputs(235)) xor (inputs(200));
    layer0_outputs(12200) <= not((inputs(178)) xor (inputs(29)));
    layer0_outputs(12201) <= '0';
    layer0_outputs(12202) <= not(inputs(131)) or (inputs(212));
    layer0_outputs(12203) <= not((inputs(197)) xor (inputs(75)));
    layer0_outputs(12204) <= '0';
    layer0_outputs(12205) <= (inputs(138)) xor (inputs(168));
    layer0_outputs(12206) <= not((inputs(136)) or (inputs(22)));
    layer0_outputs(12207) <= not(inputs(70)) or (inputs(21));
    layer0_outputs(12208) <= not((inputs(179)) and (inputs(91)));
    layer0_outputs(12209) <= not(inputs(234)) or (inputs(26));
    layer0_outputs(12210) <= not(inputs(213));
    layer0_outputs(12211) <= (inputs(106)) xor (inputs(105));
    layer0_outputs(12212) <= '1';
    layer0_outputs(12213) <= not((inputs(107)) or (inputs(143)));
    layer0_outputs(12214) <= (inputs(107)) and not (inputs(81));
    layer0_outputs(12215) <= not((inputs(68)) or (inputs(209)));
    layer0_outputs(12216) <= not((inputs(55)) or (inputs(114)));
    layer0_outputs(12217) <= not(inputs(104)) or (inputs(74));
    layer0_outputs(12218) <= not((inputs(224)) or (inputs(115)));
    layer0_outputs(12219) <= not((inputs(93)) xor (inputs(76)));
    layer0_outputs(12220) <= not((inputs(36)) xor (inputs(210)));
    layer0_outputs(12221) <= not(inputs(187)) or (inputs(224));
    layer0_outputs(12222) <= not((inputs(48)) xor (inputs(153)));
    layer0_outputs(12223) <= not((inputs(138)) xor (inputs(34)));
    layer0_outputs(12224) <= not((inputs(121)) or (inputs(138)));
    layer0_outputs(12225) <= not((inputs(126)) xor (inputs(104)));
    layer0_outputs(12226) <= inputs(143);
    layer0_outputs(12227) <= (inputs(230)) xor (inputs(34));
    layer0_outputs(12228) <= not((inputs(253)) or (inputs(34)));
    layer0_outputs(12229) <= not(inputs(178)) or (inputs(4));
    layer0_outputs(12230) <= not(inputs(72)) or (inputs(108));
    layer0_outputs(12231) <= not(inputs(132));
    layer0_outputs(12232) <= not((inputs(44)) or (inputs(42)));
    layer0_outputs(12233) <= not((inputs(255)) xor (inputs(180)));
    layer0_outputs(12234) <= (inputs(165)) and not (inputs(243));
    layer0_outputs(12235) <= (inputs(162)) and not (inputs(79));
    layer0_outputs(12236) <= (inputs(45)) or (inputs(215));
    layer0_outputs(12237) <= (inputs(26)) or (inputs(172));
    layer0_outputs(12238) <= (inputs(200)) or (inputs(66));
    layer0_outputs(12239) <= not((inputs(246)) or (inputs(169)));
    layer0_outputs(12240) <= not((inputs(110)) or (inputs(73)));
    layer0_outputs(12241) <= not((inputs(78)) or (inputs(155)));
    layer0_outputs(12242) <= inputs(236);
    layer0_outputs(12243) <= inputs(45);
    layer0_outputs(12244) <= not((inputs(76)) or (inputs(62)));
    layer0_outputs(12245) <= not((inputs(92)) or (inputs(87)));
    layer0_outputs(12246) <= inputs(148);
    layer0_outputs(12247) <= '0';
    layer0_outputs(12248) <= (inputs(246)) and not (inputs(5));
    layer0_outputs(12249) <= (inputs(173)) and not (inputs(24));
    layer0_outputs(12250) <= (inputs(80)) and (inputs(254));
    layer0_outputs(12251) <= inputs(120);
    layer0_outputs(12252) <= (inputs(1)) xor (inputs(47));
    layer0_outputs(12253) <= not((inputs(30)) xor (inputs(102)));
    layer0_outputs(12254) <= not((inputs(151)) xor (inputs(13)));
    layer0_outputs(12255) <= not((inputs(150)) and (inputs(131)));
    layer0_outputs(12256) <= inputs(165);
    layer0_outputs(12257) <= (inputs(110)) and not (inputs(6));
    layer0_outputs(12258) <= not((inputs(57)) xor (inputs(63)));
    layer0_outputs(12259) <= (inputs(182)) or (inputs(5));
    layer0_outputs(12260) <= (inputs(114)) or (inputs(43));
    layer0_outputs(12261) <= inputs(120);
    layer0_outputs(12262) <= (inputs(56)) and not (inputs(129));
    layer0_outputs(12263) <= not(inputs(122));
    layer0_outputs(12264) <= not(inputs(116));
    layer0_outputs(12265) <= inputs(83);
    layer0_outputs(12266) <= not(inputs(189));
    layer0_outputs(12267) <= (inputs(192)) or (inputs(183));
    layer0_outputs(12268) <= inputs(243);
    layer0_outputs(12269) <= (inputs(185)) and not (inputs(182));
    layer0_outputs(12270) <= not(inputs(195)) or (inputs(127));
    layer0_outputs(12271) <= not(inputs(98)) or (inputs(253));
    layer0_outputs(12272) <= '0';
    layer0_outputs(12273) <= not(inputs(178)) or (inputs(58));
    layer0_outputs(12274) <= inputs(131);
    layer0_outputs(12275) <= not(inputs(39));
    layer0_outputs(12276) <= not((inputs(86)) or (inputs(76)));
    layer0_outputs(12277) <= not((inputs(45)) xor (inputs(210)));
    layer0_outputs(12278) <= (inputs(227)) or (inputs(231));
    layer0_outputs(12279) <= not((inputs(54)) or (inputs(2)));
    layer0_outputs(12280) <= (inputs(156)) or (inputs(54));
    layer0_outputs(12281) <= not(inputs(34)) or (inputs(3));
    layer0_outputs(12282) <= (inputs(42)) xor (inputs(244));
    layer0_outputs(12283) <= not((inputs(159)) xor (inputs(64)));
    layer0_outputs(12284) <= not(inputs(180)) or (inputs(18));
    layer0_outputs(12285) <= (inputs(188)) xor (inputs(107));
    layer0_outputs(12286) <= not(inputs(94)) or (inputs(82));
    layer0_outputs(12287) <= (inputs(71)) or (inputs(231));
    layer0_outputs(12288) <= not((inputs(77)) or (inputs(12)));
    layer0_outputs(12289) <= not((inputs(249)) or (inputs(201)));
    layer0_outputs(12290) <= (inputs(69)) or (inputs(216));
    layer0_outputs(12291) <= not(inputs(101)) or (inputs(178));
    layer0_outputs(12292) <= not(inputs(188)) or (inputs(98));
    layer0_outputs(12293) <= not((inputs(178)) or (inputs(157)));
    layer0_outputs(12294) <= not((inputs(193)) xor (inputs(60)));
    layer0_outputs(12295) <= not(inputs(180));
    layer0_outputs(12296) <= not((inputs(138)) or (inputs(194)));
    layer0_outputs(12297) <= (inputs(13)) or (inputs(224));
    layer0_outputs(12298) <= not(inputs(167)) or (inputs(173));
    layer0_outputs(12299) <= (inputs(23)) xor (inputs(232));
    layer0_outputs(12300) <= (inputs(219)) and not (inputs(185));
    layer0_outputs(12301) <= (inputs(47)) and (inputs(35));
    layer0_outputs(12302) <= not(inputs(151));
    layer0_outputs(12303) <= inputs(24);
    layer0_outputs(12304) <= not(inputs(26));
    layer0_outputs(12305) <= not(inputs(198));
    layer0_outputs(12306) <= (inputs(155)) or (inputs(77));
    layer0_outputs(12307) <= (inputs(166)) xor (inputs(66));
    layer0_outputs(12308) <= not(inputs(101)) or (inputs(81));
    layer0_outputs(12309) <= not((inputs(50)) or (inputs(209)));
    layer0_outputs(12310) <= not(inputs(120)) or (inputs(155));
    layer0_outputs(12311) <= '1';
    layer0_outputs(12312) <= not((inputs(42)) xor (inputs(178)));
    layer0_outputs(12313) <= not((inputs(67)) or (inputs(178)));
    layer0_outputs(12314) <= inputs(106);
    layer0_outputs(12315) <= (inputs(45)) and (inputs(218));
    layer0_outputs(12316) <= (inputs(32)) and (inputs(183));
    layer0_outputs(12317) <= not(inputs(33));
    layer0_outputs(12318) <= not((inputs(201)) xor (inputs(201)));
    layer0_outputs(12319) <= (inputs(199)) and not (inputs(98));
    layer0_outputs(12320) <= not((inputs(219)) xor (inputs(184)));
    layer0_outputs(12321) <= (inputs(245)) xor (inputs(178));
    layer0_outputs(12322) <= not((inputs(57)) and (inputs(57)));
    layer0_outputs(12323) <= not((inputs(119)) and (inputs(224)));
    layer0_outputs(12324) <= (inputs(162)) xor (inputs(183));
    layer0_outputs(12325) <= (inputs(122)) xor (inputs(236));
    layer0_outputs(12326) <= not((inputs(108)) or (inputs(68)));
    layer0_outputs(12327) <= not((inputs(168)) xor (inputs(187)));
    layer0_outputs(12328) <= (inputs(128)) xor (inputs(150));
    layer0_outputs(12329) <= (inputs(19)) and (inputs(13));
    layer0_outputs(12330) <= inputs(118);
    layer0_outputs(12331) <= not((inputs(45)) or (inputs(116)));
    layer0_outputs(12332) <= (inputs(178)) xor (inputs(54));
    layer0_outputs(12333) <= (inputs(67)) or (inputs(189));
    layer0_outputs(12334) <= (inputs(79)) or (inputs(55));
    layer0_outputs(12335) <= not(inputs(188)) or (inputs(62));
    layer0_outputs(12336) <= (inputs(140)) and not (inputs(51));
    layer0_outputs(12337) <= '1';
    layer0_outputs(12338) <= (inputs(83)) or (inputs(155));
    layer0_outputs(12339) <= (inputs(47)) or (inputs(121));
    layer0_outputs(12340) <= inputs(45);
    layer0_outputs(12341) <= inputs(23);
    layer0_outputs(12342) <= (inputs(38)) xor (inputs(46));
    layer0_outputs(12343) <= inputs(49);
    layer0_outputs(12344) <= not((inputs(219)) xor (inputs(158)));
    layer0_outputs(12345) <= not(inputs(86)) or (inputs(250));
    layer0_outputs(12346) <= not(inputs(104));
    layer0_outputs(12347) <= not(inputs(66));
    layer0_outputs(12348) <= (inputs(225)) and not (inputs(190));
    layer0_outputs(12349) <= (inputs(250)) xor (inputs(73));
    layer0_outputs(12350) <= (inputs(154)) and not (inputs(118));
    layer0_outputs(12351) <= (inputs(19)) or (inputs(147));
    layer0_outputs(12352) <= not(inputs(150));
    layer0_outputs(12353) <= not((inputs(161)) and (inputs(220)));
    layer0_outputs(12354) <= (inputs(122)) and not (inputs(150));
    layer0_outputs(12355) <= (inputs(250)) and not (inputs(5));
    layer0_outputs(12356) <= (inputs(232)) and not (inputs(144));
    layer0_outputs(12357) <= not((inputs(11)) and (inputs(20)));
    layer0_outputs(12358) <= not((inputs(92)) xor (inputs(238)));
    layer0_outputs(12359) <= not((inputs(75)) xor (inputs(50)));
    layer0_outputs(12360) <= not((inputs(132)) xor (inputs(30)));
    layer0_outputs(12361) <= not((inputs(160)) and (inputs(59)));
    layer0_outputs(12362) <= '1';
    layer0_outputs(12363) <= inputs(36);
    layer0_outputs(12364) <= (inputs(15)) and not (inputs(17));
    layer0_outputs(12365) <= (inputs(103)) and not (inputs(147));
    layer0_outputs(12366) <= not(inputs(134)) or (inputs(233));
    layer0_outputs(12367) <= (inputs(177)) or (inputs(39));
    layer0_outputs(12368) <= (inputs(37)) and not (inputs(78));
    layer0_outputs(12369) <= (inputs(22)) or (inputs(246));
    layer0_outputs(12370) <= not(inputs(60)) or (inputs(126));
    layer0_outputs(12371) <= not(inputs(72)) or (inputs(40));
    layer0_outputs(12372) <= not(inputs(92)) or (inputs(224));
    layer0_outputs(12373) <= not((inputs(122)) xor (inputs(111)));
    layer0_outputs(12374) <= not(inputs(174));
    layer0_outputs(12375) <= not((inputs(107)) xor (inputs(58)));
    layer0_outputs(12376) <= (inputs(86)) and not (inputs(182));
    layer0_outputs(12377) <= (inputs(163)) and not (inputs(115));
    layer0_outputs(12378) <= not((inputs(109)) or (inputs(92)));
    layer0_outputs(12379) <= '0';
    layer0_outputs(12380) <= (inputs(155)) or (inputs(182));
    layer0_outputs(12381) <= not((inputs(88)) xor (inputs(255)));
    layer0_outputs(12382) <= (inputs(85)) xor (inputs(189));
    layer0_outputs(12383) <= (inputs(214)) xor (inputs(143));
    layer0_outputs(12384) <= '0';
    layer0_outputs(12385) <= (inputs(12)) xor (inputs(232));
    layer0_outputs(12386) <= (inputs(204)) or (inputs(207));
    layer0_outputs(12387) <= (inputs(171)) and not (inputs(239));
    layer0_outputs(12388) <= (inputs(214)) xor (inputs(50));
    layer0_outputs(12389) <= inputs(167);
    layer0_outputs(12390) <= not((inputs(19)) xor (inputs(54)));
    layer0_outputs(12391) <= inputs(96);
    layer0_outputs(12392) <= (inputs(119)) and not (inputs(176));
    layer0_outputs(12393) <= (inputs(62)) or (inputs(194));
    layer0_outputs(12394) <= not((inputs(209)) and (inputs(3)));
    layer0_outputs(12395) <= (inputs(27)) and (inputs(145));
    layer0_outputs(12396) <= (inputs(75)) xor (inputs(56));
    layer0_outputs(12397) <= (inputs(73)) xor (inputs(99));
    layer0_outputs(12398) <= (inputs(100)) and (inputs(116));
    layer0_outputs(12399) <= not(inputs(141));
    layer0_outputs(12400) <= (inputs(127)) or (inputs(53));
    layer0_outputs(12401) <= (inputs(133)) xor (inputs(229));
    layer0_outputs(12402) <= inputs(149);
    layer0_outputs(12403) <= not((inputs(150)) xor (inputs(238)));
    layer0_outputs(12404) <= not((inputs(24)) xor (inputs(234)));
    layer0_outputs(12405) <= not(inputs(231));
    layer0_outputs(12406) <= not(inputs(233)) or (inputs(221));
    layer0_outputs(12407) <= not(inputs(106)) or (inputs(232));
    layer0_outputs(12408) <= (inputs(116)) or (inputs(23));
    layer0_outputs(12409) <= not((inputs(93)) xor (inputs(172)));
    layer0_outputs(12410) <= (inputs(221)) and (inputs(71));
    layer0_outputs(12411) <= not(inputs(167));
    layer0_outputs(12412) <= (inputs(43)) and not (inputs(4));
    layer0_outputs(12413) <= inputs(57);
    layer0_outputs(12414) <= not(inputs(29));
    layer0_outputs(12415) <= not(inputs(87));
    layer0_outputs(12416) <= not(inputs(73));
    layer0_outputs(12417) <= not(inputs(150));
    layer0_outputs(12418) <= '1';
    layer0_outputs(12419) <= not(inputs(62)) or (inputs(248));
    layer0_outputs(12420) <= inputs(243);
    layer0_outputs(12421) <= (inputs(52)) and not (inputs(94));
    layer0_outputs(12422) <= not(inputs(75));
    layer0_outputs(12423) <= (inputs(184)) and not (inputs(143));
    layer0_outputs(12424) <= not((inputs(228)) or (inputs(153)));
    layer0_outputs(12425) <= (inputs(228)) or (inputs(172));
    layer0_outputs(12426) <= inputs(250);
    layer0_outputs(12427) <= (inputs(67)) xor (inputs(195));
    layer0_outputs(12428) <= '0';
    layer0_outputs(12429) <= inputs(94);
    layer0_outputs(12430) <= not(inputs(186));
    layer0_outputs(12431) <= (inputs(26)) and not (inputs(69));
    layer0_outputs(12432) <= inputs(72);
    layer0_outputs(12433) <= inputs(148);
    layer0_outputs(12434) <= (inputs(86)) xor (inputs(193));
    layer0_outputs(12435) <= not(inputs(55)) or (inputs(231));
    layer0_outputs(12436) <= '0';
    layer0_outputs(12437) <= not((inputs(144)) xor (inputs(238)));
    layer0_outputs(12438) <= '0';
    layer0_outputs(12439) <= not(inputs(242)) or (inputs(227));
    layer0_outputs(12440) <= (inputs(117)) xor (inputs(109));
    layer0_outputs(12441) <= '1';
    layer0_outputs(12442) <= (inputs(34)) and (inputs(15));
    layer0_outputs(12443) <= not(inputs(123));
    layer0_outputs(12444) <= (inputs(182)) and (inputs(134));
    layer0_outputs(12445) <= not(inputs(104)) or (inputs(148));
    layer0_outputs(12446) <= not(inputs(101)) or (inputs(244));
    layer0_outputs(12447) <= not(inputs(127)) or (inputs(88));
    layer0_outputs(12448) <= (inputs(229)) xor (inputs(232));
    layer0_outputs(12449) <= not(inputs(212));
    layer0_outputs(12450) <= inputs(202);
    layer0_outputs(12451) <= (inputs(30)) xor (inputs(96));
    layer0_outputs(12452) <= not(inputs(39));
    layer0_outputs(12453) <= inputs(104);
    layer0_outputs(12454) <= (inputs(180)) or (inputs(58));
    layer0_outputs(12455) <= inputs(188);
    layer0_outputs(12456) <= not(inputs(83));
    layer0_outputs(12457) <= (inputs(114)) xor (inputs(5));
    layer0_outputs(12458) <= (inputs(143)) and not (inputs(145));
    layer0_outputs(12459) <= not(inputs(202)) or (inputs(100));
    layer0_outputs(12460) <= inputs(165);
    layer0_outputs(12461) <= (inputs(63)) and not (inputs(227));
    layer0_outputs(12462) <= not((inputs(1)) or (inputs(125)));
    layer0_outputs(12463) <= not((inputs(239)) and (inputs(70)));
    layer0_outputs(12464) <= not(inputs(9)) or (inputs(74));
    layer0_outputs(12465) <= not((inputs(103)) or (inputs(165)));
    layer0_outputs(12466) <= (inputs(125)) or (inputs(228));
    layer0_outputs(12467) <= (inputs(7)) and not (inputs(44));
    layer0_outputs(12468) <= not((inputs(70)) or (inputs(190)));
    layer0_outputs(12469) <= not((inputs(83)) or (inputs(231)));
    layer0_outputs(12470) <= '0';
    layer0_outputs(12471) <= not(inputs(161));
    layer0_outputs(12472) <= (inputs(111)) xor (inputs(51));
    layer0_outputs(12473) <= not((inputs(76)) or (inputs(48)));
    layer0_outputs(12474) <= not(inputs(38));
    layer0_outputs(12475) <= '0';
    layer0_outputs(12476) <= (inputs(193)) or (inputs(201));
    layer0_outputs(12477) <= not((inputs(72)) and (inputs(193)));
    layer0_outputs(12478) <= not((inputs(234)) or (inputs(228)));
    layer0_outputs(12479) <= not((inputs(79)) or (inputs(253)));
    layer0_outputs(12480) <= not((inputs(196)) or (inputs(9)));
    layer0_outputs(12481) <= '1';
    layer0_outputs(12482) <= inputs(10);
    layer0_outputs(12483) <= inputs(22);
    layer0_outputs(12484) <= not(inputs(22));
    layer0_outputs(12485) <= (inputs(56)) or (inputs(109));
    layer0_outputs(12486) <= inputs(95);
    layer0_outputs(12487) <= not(inputs(183)) or (inputs(223));
    layer0_outputs(12488) <= '1';
    layer0_outputs(12489) <= (inputs(103)) and not (inputs(221));
    layer0_outputs(12490) <= (inputs(243)) or (inputs(255));
    layer0_outputs(12491) <= not((inputs(155)) xor (inputs(143)));
    layer0_outputs(12492) <= (inputs(41)) xor (inputs(72));
    layer0_outputs(12493) <= not(inputs(209)) or (inputs(124));
    layer0_outputs(12494) <= not((inputs(83)) xor (inputs(8)));
    layer0_outputs(12495) <= not(inputs(87)) or (inputs(95));
    layer0_outputs(12496) <= not(inputs(27));
    layer0_outputs(12497) <= inputs(181);
    layer0_outputs(12498) <= not(inputs(231)) or (inputs(38));
    layer0_outputs(12499) <= not((inputs(230)) and (inputs(252)));
    layer0_outputs(12500) <= inputs(254);
    layer0_outputs(12501) <= (inputs(74)) or (inputs(192));
    layer0_outputs(12502) <= (inputs(8)) and (inputs(169));
    layer0_outputs(12503) <= not((inputs(168)) xor (inputs(104)));
    layer0_outputs(12504) <= inputs(42);
    layer0_outputs(12505) <= not((inputs(73)) xor (inputs(215)));
    layer0_outputs(12506) <= (inputs(59)) or (inputs(176));
    layer0_outputs(12507) <= inputs(224);
    layer0_outputs(12508) <= not(inputs(130)) or (inputs(96));
    layer0_outputs(12509) <= not(inputs(140)) or (inputs(217));
    layer0_outputs(12510) <= not((inputs(109)) xor (inputs(235)));
    layer0_outputs(12511) <= (inputs(9)) and (inputs(126));
    layer0_outputs(12512) <= not((inputs(106)) xor (inputs(239)));
    layer0_outputs(12513) <= (inputs(59)) and not (inputs(239));
    layer0_outputs(12514) <= not((inputs(82)) or (inputs(196)));
    layer0_outputs(12515) <= (inputs(67)) and not (inputs(157));
    layer0_outputs(12516) <= not((inputs(61)) or (inputs(101)));
    layer0_outputs(12517) <= (inputs(163)) xor (inputs(14));
    layer0_outputs(12518) <= (inputs(175)) and (inputs(25));
    layer0_outputs(12519) <= not(inputs(179)) or (inputs(128));
    layer0_outputs(12520) <= not((inputs(153)) xor (inputs(32)));
    layer0_outputs(12521) <= (inputs(203)) or (inputs(175));
    layer0_outputs(12522) <= (inputs(24)) and not (inputs(78));
    layer0_outputs(12523) <= not((inputs(132)) and (inputs(132)));
    layer0_outputs(12524) <= (inputs(237)) or (inputs(210));
    layer0_outputs(12525) <= (inputs(97)) xor (inputs(78));
    layer0_outputs(12526) <= (inputs(12)) and not (inputs(162));
    layer0_outputs(12527) <= (inputs(4)) xor (inputs(149));
    layer0_outputs(12528) <= inputs(220);
    layer0_outputs(12529) <= not(inputs(127)) or (inputs(242));
    layer0_outputs(12530) <= not((inputs(169)) or (inputs(161)));
    layer0_outputs(12531) <= not((inputs(128)) xor (inputs(72)));
    layer0_outputs(12532) <= not((inputs(4)) and (inputs(238)));
    layer0_outputs(12533) <= not((inputs(96)) and (inputs(53)));
    layer0_outputs(12534) <= not((inputs(13)) xor (inputs(120)));
    layer0_outputs(12535) <= not((inputs(63)) and (inputs(99)));
    layer0_outputs(12536) <= (inputs(144)) or (inputs(119));
    layer0_outputs(12537) <= not((inputs(204)) or (inputs(202)));
    layer0_outputs(12538) <= (inputs(114)) or (inputs(148));
    layer0_outputs(12539) <= not(inputs(151)) or (inputs(174));
    layer0_outputs(12540) <= not(inputs(104)) or (inputs(66));
    layer0_outputs(12541) <= (inputs(198)) or (inputs(74));
    layer0_outputs(12542) <= '1';
    layer0_outputs(12543) <= not(inputs(244));
    layer0_outputs(12544) <= (inputs(213)) or (inputs(98));
    layer0_outputs(12545) <= (inputs(155)) and not (inputs(252));
    layer0_outputs(12546) <= (inputs(163)) xor (inputs(171));
    layer0_outputs(12547) <= (inputs(142)) or (inputs(231));
    layer0_outputs(12548) <= not((inputs(9)) or (inputs(115)));
    layer0_outputs(12549) <= not(inputs(53)) or (inputs(64));
    layer0_outputs(12550) <= (inputs(24)) and (inputs(183));
    layer0_outputs(12551) <= (inputs(49)) or (inputs(213));
    layer0_outputs(12552) <= (inputs(99)) or (inputs(40));
    layer0_outputs(12553) <= (inputs(192)) and not (inputs(82));
    layer0_outputs(12554) <= (inputs(192)) and (inputs(159));
    layer0_outputs(12555) <= not(inputs(241));
    layer0_outputs(12556) <= not(inputs(136));
    layer0_outputs(12557) <= '0';
    layer0_outputs(12558) <= (inputs(229)) xor (inputs(125));
    layer0_outputs(12559) <= not((inputs(247)) or (inputs(254)));
    layer0_outputs(12560) <= not(inputs(10));
    layer0_outputs(12561) <= '0';
    layer0_outputs(12562) <= (inputs(159)) and not (inputs(145));
    layer0_outputs(12563) <= inputs(122);
    layer0_outputs(12564) <= not(inputs(135)) or (inputs(125));
    layer0_outputs(12565) <= inputs(57);
    layer0_outputs(12566) <= not(inputs(169));
    layer0_outputs(12567) <= not((inputs(99)) or (inputs(250)));
    layer0_outputs(12568) <= (inputs(76)) xor (inputs(33));
    layer0_outputs(12569) <= (inputs(93)) or (inputs(190));
    layer0_outputs(12570) <= not(inputs(219)) or (inputs(239));
    layer0_outputs(12571) <= (inputs(14)) and not (inputs(78));
    layer0_outputs(12572) <= (inputs(160)) and not (inputs(191));
    layer0_outputs(12573) <= (inputs(133)) and not (inputs(194));
    layer0_outputs(12574) <= (inputs(10)) xor (inputs(136));
    layer0_outputs(12575) <= not((inputs(48)) xor (inputs(93)));
    layer0_outputs(12576) <= (inputs(88)) and not (inputs(244));
    layer0_outputs(12577) <= not((inputs(229)) and (inputs(178)));
    layer0_outputs(12578) <= (inputs(220)) or (inputs(59));
    layer0_outputs(12579) <= not(inputs(13)) or (inputs(246));
    layer0_outputs(12580) <= inputs(24);
    layer0_outputs(12581) <= not(inputs(38));
    layer0_outputs(12582) <= (inputs(170)) or (inputs(231));
    layer0_outputs(12583) <= inputs(214);
    layer0_outputs(12584) <= not((inputs(98)) or (inputs(133)));
    layer0_outputs(12585) <= (inputs(199)) or (inputs(31));
    layer0_outputs(12586) <= not(inputs(10)) or (inputs(0));
    layer0_outputs(12587) <= (inputs(12)) and not (inputs(30));
    layer0_outputs(12588) <= (inputs(121)) or (inputs(4));
    layer0_outputs(12589) <= (inputs(147)) or (inputs(138));
    layer0_outputs(12590) <= inputs(91);
    layer0_outputs(12591) <= (inputs(69)) or (inputs(207));
    layer0_outputs(12592) <= not((inputs(29)) or (inputs(245)));
    layer0_outputs(12593) <= '1';
    layer0_outputs(12594) <= not((inputs(53)) xor (inputs(181)));
    layer0_outputs(12595) <= not((inputs(114)) xor (inputs(231)));
    layer0_outputs(12596) <= not((inputs(128)) and (inputs(18)));
    layer0_outputs(12597) <= not(inputs(85)) or (inputs(166));
    layer0_outputs(12598) <= (inputs(58)) and not (inputs(35));
    layer0_outputs(12599) <= not((inputs(128)) xor (inputs(67)));
    layer0_outputs(12600) <= not((inputs(104)) or (inputs(246)));
    layer0_outputs(12601) <= (inputs(244)) or (inputs(132));
    layer0_outputs(12602) <= not((inputs(172)) or (inputs(49)));
    layer0_outputs(12603) <= not(inputs(179));
    layer0_outputs(12604) <= (inputs(25)) and not (inputs(15));
    layer0_outputs(12605) <= not(inputs(81));
    layer0_outputs(12606) <= '1';
    layer0_outputs(12607) <= not((inputs(247)) or (inputs(53)));
    layer0_outputs(12608) <= inputs(180);
    layer0_outputs(12609) <= (inputs(67)) and not (inputs(173));
    layer0_outputs(12610) <= inputs(156);
    layer0_outputs(12611) <= not((inputs(139)) xor (inputs(68)));
    layer0_outputs(12612) <= not(inputs(60)) or (inputs(65));
    layer0_outputs(12613) <= (inputs(184)) or (inputs(221));
    layer0_outputs(12614) <= (inputs(172)) and not (inputs(159));
    layer0_outputs(12615) <= (inputs(135)) or (inputs(139));
    layer0_outputs(12616) <= not(inputs(233));
    layer0_outputs(12617) <= not((inputs(203)) xor (inputs(214)));
    layer0_outputs(12618) <= not((inputs(181)) or (inputs(47)));
    layer0_outputs(12619) <= not((inputs(212)) and (inputs(106)));
    layer0_outputs(12620) <= (inputs(149)) and not (inputs(114));
    layer0_outputs(12621) <= not((inputs(255)) xor (inputs(232)));
    layer0_outputs(12622) <= not((inputs(110)) or (inputs(202)));
    layer0_outputs(12623) <= not((inputs(135)) or (inputs(134)));
    layer0_outputs(12624) <= not(inputs(156));
    layer0_outputs(12625) <= (inputs(213)) xor (inputs(158));
    layer0_outputs(12626) <= inputs(223);
    layer0_outputs(12627) <= not((inputs(89)) xor (inputs(233)));
    layer0_outputs(12628) <= not((inputs(233)) or (inputs(93)));
    layer0_outputs(12629) <= not(inputs(209)) or (inputs(81));
    layer0_outputs(12630) <= not((inputs(202)) xor (inputs(225)));
    layer0_outputs(12631) <= (inputs(90)) and not (inputs(203));
    layer0_outputs(12632) <= not((inputs(82)) and (inputs(10)));
    layer0_outputs(12633) <= (inputs(70)) xor (inputs(10));
    layer0_outputs(12634) <= not((inputs(177)) and (inputs(35)));
    layer0_outputs(12635) <= inputs(54);
    layer0_outputs(12636) <= (inputs(21)) or (inputs(89));
    layer0_outputs(12637) <= not(inputs(90));
    layer0_outputs(12638) <= not(inputs(39));
    layer0_outputs(12639) <= (inputs(174)) or (inputs(203));
    layer0_outputs(12640) <= not((inputs(193)) or (inputs(184)));
    layer0_outputs(12641) <= (inputs(213)) xor (inputs(237));
    layer0_outputs(12642) <= (inputs(2)) and not (inputs(4));
    layer0_outputs(12643) <= not((inputs(150)) xor (inputs(97)));
    layer0_outputs(12644) <= (inputs(15)) or (inputs(76));
    layer0_outputs(12645) <= not(inputs(249));
    layer0_outputs(12646) <= (inputs(108)) and not (inputs(124));
    layer0_outputs(12647) <= (inputs(112)) or (inputs(172));
    layer0_outputs(12648) <= not(inputs(129)) or (inputs(39));
    layer0_outputs(12649) <= not(inputs(114));
    layer0_outputs(12650) <= (inputs(91)) and not (inputs(161));
    layer0_outputs(12651) <= not((inputs(246)) xor (inputs(82)));
    layer0_outputs(12652) <= inputs(124);
    layer0_outputs(12653) <= (inputs(237)) or (inputs(34));
    layer0_outputs(12654) <= (inputs(148)) and not (inputs(208));
    layer0_outputs(12655) <= not((inputs(169)) xor (inputs(112)));
    layer0_outputs(12656) <= not((inputs(204)) xor (inputs(173)));
    layer0_outputs(12657) <= not((inputs(179)) xor (inputs(156)));
    layer0_outputs(12658) <= (inputs(225)) and not (inputs(238));
    layer0_outputs(12659) <= not((inputs(200)) xor (inputs(249)));
    layer0_outputs(12660) <= (inputs(129)) xor (inputs(43));
    layer0_outputs(12661) <= not(inputs(136));
    layer0_outputs(12662) <= '0';
    layer0_outputs(12663) <= not((inputs(204)) or (inputs(33)));
    layer0_outputs(12664) <= (inputs(216)) or (inputs(110));
    layer0_outputs(12665) <= not((inputs(111)) xor (inputs(181)));
    layer0_outputs(12666) <= (inputs(5)) xor (inputs(167));
    layer0_outputs(12667) <= (inputs(217)) and not (inputs(65));
    layer0_outputs(12668) <= (inputs(244)) and not (inputs(2));
    layer0_outputs(12669) <= not(inputs(215));
    layer0_outputs(12670) <= inputs(71);
    layer0_outputs(12671) <= inputs(133);
    layer0_outputs(12672) <= (inputs(245)) or (inputs(57));
    layer0_outputs(12673) <= not(inputs(146)) or (inputs(62));
    layer0_outputs(12674) <= not(inputs(74)) or (inputs(240));
    layer0_outputs(12675) <= (inputs(55)) or (inputs(20));
    layer0_outputs(12676) <= (inputs(233)) or (inputs(33));
    layer0_outputs(12677) <= (inputs(238)) xor (inputs(138));
    layer0_outputs(12678) <= not((inputs(86)) or (inputs(26)));
    layer0_outputs(12679) <= '0';
    layer0_outputs(12680) <= not(inputs(149));
    layer0_outputs(12681) <= not(inputs(92)) or (inputs(177));
    layer0_outputs(12682) <= (inputs(101)) xor (inputs(127));
    layer0_outputs(12683) <= (inputs(75)) and not (inputs(18));
    layer0_outputs(12684) <= (inputs(208)) xor (inputs(109));
    layer0_outputs(12685) <= not(inputs(205));
    layer0_outputs(12686) <= not(inputs(96));
    layer0_outputs(12687) <= inputs(246);
    layer0_outputs(12688) <= not(inputs(40));
    layer0_outputs(12689) <= not((inputs(219)) or (inputs(222)));
    layer0_outputs(12690) <= not((inputs(47)) or (inputs(229)));
    layer0_outputs(12691) <= (inputs(94)) and not (inputs(24));
    layer0_outputs(12692) <= not((inputs(223)) xor (inputs(217)));
    layer0_outputs(12693) <= not(inputs(12)) or (inputs(227));
    layer0_outputs(12694) <= (inputs(116)) and not (inputs(110));
    layer0_outputs(12695) <= not((inputs(174)) or (inputs(58)));
    layer0_outputs(12696) <= (inputs(88)) and not (inputs(116));
    layer0_outputs(12697) <= (inputs(57)) and not (inputs(97));
    layer0_outputs(12698) <= (inputs(184)) and not (inputs(37));
    layer0_outputs(12699) <= not((inputs(104)) or (inputs(146)));
    layer0_outputs(12700) <= not(inputs(238));
    layer0_outputs(12701) <= (inputs(188)) or (inputs(117));
    layer0_outputs(12702) <= (inputs(68)) xor (inputs(108));
    layer0_outputs(12703) <= (inputs(225)) and not (inputs(175));
    layer0_outputs(12704) <= not((inputs(194)) or (inputs(57)));
    layer0_outputs(12705) <= not(inputs(137)) or (inputs(162));
    layer0_outputs(12706) <= inputs(67);
    layer0_outputs(12707) <= not((inputs(216)) or (inputs(164)));
    layer0_outputs(12708) <= (inputs(70)) and not (inputs(89));
    layer0_outputs(12709) <= not((inputs(211)) xor (inputs(151)));
    layer0_outputs(12710) <= not(inputs(223));
    layer0_outputs(12711) <= not(inputs(205)) or (inputs(51));
    layer0_outputs(12712) <= not((inputs(147)) or (inputs(172)));
    layer0_outputs(12713) <= not((inputs(199)) xor (inputs(28)));
    layer0_outputs(12714) <= not((inputs(156)) xor (inputs(129)));
    layer0_outputs(12715) <= not(inputs(24));
    layer0_outputs(12716) <= (inputs(219)) and not (inputs(240));
    layer0_outputs(12717) <= (inputs(199)) and not (inputs(230));
    layer0_outputs(12718) <= (inputs(176)) xor (inputs(117));
    layer0_outputs(12719) <= not(inputs(155));
    layer0_outputs(12720) <= not(inputs(119));
    layer0_outputs(12721) <= (inputs(11)) and (inputs(189));
    layer0_outputs(12722) <= not(inputs(196));
    layer0_outputs(12723) <= not(inputs(54)) or (inputs(22));
    layer0_outputs(12724) <= (inputs(4)) and (inputs(145));
    layer0_outputs(12725) <= not(inputs(121)) or (inputs(247));
    layer0_outputs(12726) <= inputs(102);
    layer0_outputs(12727) <= not((inputs(38)) xor (inputs(224)));
    layer0_outputs(12728) <= (inputs(100)) and not (inputs(228));
    layer0_outputs(12729) <= not(inputs(62));
    layer0_outputs(12730) <= (inputs(72)) and not (inputs(26));
    layer0_outputs(12731) <= not((inputs(161)) and (inputs(70)));
    layer0_outputs(12732) <= not((inputs(248)) xor (inputs(8)));
    layer0_outputs(12733) <= not(inputs(187)) or (inputs(93));
    layer0_outputs(12734) <= (inputs(56)) and not (inputs(205));
    layer0_outputs(12735) <= (inputs(36)) or (inputs(89));
    layer0_outputs(12736) <= not((inputs(33)) xor (inputs(110)));
    layer0_outputs(12737) <= not(inputs(59));
    layer0_outputs(12738) <= not((inputs(51)) xor (inputs(233)));
    layer0_outputs(12739) <= (inputs(217)) and not (inputs(251));
    layer0_outputs(12740) <= not((inputs(238)) xor (inputs(149)));
    layer0_outputs(12741) <= (inputs(170)) xor (inputs(107));
    layer0_outputs(12742) <= (inputs(132)) or (inputs(32));
    layer0_outputs(12743) <= not(inputs(181)) or (inputs(112));
    layer0_outputs(12744) <= (inputs(212)) or (inputs(189));
    layer0_outputs(12745) <= (inputs(154)) and not (inputs(219));
    layer0_outputs(12746) <= (inputs(152)) and not (inputs(186));
    layer0_outputs(12747) <= not(inputs(121));
    layer0_outputs(12748) <= not((inputs(75)) or (inputs(114)));
    layer0_outputs(12749) <= (inputs(187)) xor (inputs(64));
    layer0_outputs(12750) <= (inputs(173)) and not (inputs(34));
    layer0_outputs(12751) <= inputs(221);
    layer0_outputs(12752) <= (inputs(69)) xor (inputs(208));
    layer0_outputs(12753) <= not((inputs(222)) and (inputs(110)));
    layer0_outputs(12754) <= not(inputs(202));
    layer0_outputs(12755) <= not((inputs(25)) xor (inputs(10)));
    layer0_outputs(12756) <= not((inputs(41)) xor (inputs(173)));
    layer0_outputs(12757) <= inputs(37);
    layer0_outputs(12758) <= (inputs(135)) and not (inputs(228));
    layer0_outputs(12759) <= inputs(115);
    layer0_outputs(12760) <= (inputs(15)) and not (inputs(98));
    layer0_outputs(12761) <= (inputs(72)) and not (inputs(19));
    layer0_outputs(12762) <= not((inputs(46)) or (inputs(127)));
    layer0_outputs(12763) <= not((inputs(8)) or (inputs(130)));
    layer0_outputs(12764) <= (inputs(119)) xor (inputs(65));
    layer0_outputs(12765) <= not(inputs(179)) or (inputs(79));
    layer0_outputs(12766) <= (inputs(229)) or (inputs(139));
    layer0_outputs(12767) <= not((inputs(158)) xor (inputs(61)));
    layer0_outputs(12768) <= not(inputs(116));
    layer0_outputs(12769) <= (inputs(207)) or (inputs(69));
    layer0_outputs(12770) <= not(inputs(172)) or (inputs(108));
    layer0_outputs(12771) <= not((inputs(26)) and (inputs(178)));
    layer0_outputs(12772) <= (inputs(8)) or (inputs(121));
    layer0_outputs(12773) <= (inputs(127)) and not (inputs(9));
    layer0_outputs(12774) <= (inputs(219)) or (inputs(114));
    layer0_outputs(12775) <= not((inputs(214)) xor (inputs(182)));
    layer0_outputs(12776) <= (inputs(193)) xor (inputs(44));
    layer0_outputs(12777) <= '1';
    layer0_outputs(12778) <= not(inputs(101)) or (inputs(226));
    layer0_outputs(12779) <= not((inputs(240)) xor (inputs(154)));
    layer0_outputs(12780) <= not(inputs(19)) or (inputs(246));
    layer0_outputs(12781) <= (inputs(39)) or (inputs(162));
    layer0_outputs(12782) <= not(inputs(89));
    layer0_outputs(12783) <= '1';
    layer0_outputs(12784) <= not(inputs(29)) or (inputs(162));
    layer0_outputs(12785) <= not(inputs(103));
    layer0_outputs(12786) <= not((inputs(243)) or (inputs(117)));
    layer0_outputs(12787) <= (inputs(40)) and not (inputs(99));
    layer0_outputs(12788) <= not(inputs(62));
    layer0_outputs(12789) <= not(inputs(24)) or (inputs(252));
    layer0_outputs(12790) <= inputs(121);
    layer0_outputs(12791) <= not(inputs(152));
    layer0_outputs(12792) <= not(inputs(4)) or (inputs(48));
    layer0_outputs(12793) <= (inputs(84)) and (inputs(226));
    layer0_outputs(12794) <= not(inputs(46));
    layer0_outputs(12795) <= inputs(68);
    layer0_outputs(12796) <= not(inputs(153));
    layer0_outputs(12797) <= (inputs(51)) and not (inputs(126));
    layer0_outputs(12798) <= not((inputs(176)) and (inputs(47)));
    layer0_outputs(12799) <= (inputs(21)) xor (inputs(30));
    outputs(0) <= layer0_outputs(10097);
    outputs(1) <= (layer0_outputs(8601)) and (layer0_outputs(3347));
    outputs(2) <= layer0_outputs(12485);
    outputs(3) <= layer0_outputs(6084);
    outputs(4) <= layer0_outputs(11800);
    outputs(5) <= not(layer0_outputs(4385)) or (layer0_outputs(838));
    outputs(6) <= not((layer0_outputs(4756)) xor (layer0_outputs(8467)));
    outputs(7) <= (layer0_outputs(12023)) xor (layer0_outputs(5154));
    outputs(8) <= not((layer0_outputs(10298)) or (layer0_outputs(10552)));
    outputs(9) <= not(layer0_outputs(3591));
    outputs(10) <= not(layer0_outputs(4884));
    outputs(11) <= layer0_outputs(5305);
    outputs(12) <= layer0_outputs(2259);
    outputs(13) <= not((layer0_outputs(3839)) or (layer0_outputs(1615)));
    outputs(14) <= layer0_outputs(1237);
    outputs(15) <= not((layer0_outputs(10881)) xor (layer0_outputs(1600)));
    outputs(16) <= not(layer0_outputs(11247)) or (layer0_outputs(5724));
    outputs(17) <= not(layer0_outputs(4638));
    outputs(18) <= not(layer0_outputs(5181));
    outputs(19) <= layer0_outputs(9111);
    outputs(20) <= (layer0_outputs(10050)) and not (layer0_outputs(6428));
    outputs(21) <= not(layer0_outputs(1554));
    outputs(22) <= layer0_outputs(9773);
    outputs(23) <= layer0_outputs(11735);
    outputs(24) <= (layer0_outputs(9037)) xor (layer0_outputs(6714));
    outputs(25) <= layer0_outputs(3379);
    outputs(26) <= not((layer0_outputs(761)) or (layer0_outputs(2111)));
    outputs(27) <= not(layer0_outputs(6348)) or (layer0_outputs(7396));
    outputs(28) <= (layer0_outputs(6550)) and (layer0_outputs(692));
    outputs(29) <= (layer0_outputs(2930)) xor (layer0_outputs(3934));
    outputs(30) <= (layer0_outputs(2859)) and (layer0_outputs(5522));
    outputs(31) <= '1';
    outputs(32) <= not((layer0_outputs(11486)) or (layer0_outputs(12017)));
    outputs(33) <= not(layer0_outputs(4326));
    outputs(34) <= layer0_outputs(3974);
    outputs(35) <= not((layer0_outputs(9309)) xor (layer0_outputs(2423)));
    outputs(36) <= (layer0_outputs(3434)) xor (layer0_outputs(5731));
    outputs(37) <= not((layer0_outputs(6590)) xor (layer0_outputs(4408)));
    outputs(38) <= (layer0_outputs(9503)) and (layer0_outputs(4769));
    outputs(39) <= not((layer0_outputs(6803)) and (layer0_outputs(12543)));
    outputs(40) <= (layer0_outputs(4611)) xor (layer0_outputs(1));
    outputs(41) <= (layer0_outputs(6331)) or (layer0_outputs(9016));
    outputs(42) <= (layer0_outputs(11528)) xor (layer0_outputs(11818));
    outputs(43) <= not(layer0_outputs(2967));
    outputs(44) <= not((layer0_outputs(1799)) or (layer0_outputs(816)));
    outputs(45) <= (layer0_outputs(1493)) or (layer0_outputs(12579));
    outputs(46) <= not(layer0_outputs(866));
    outputs(47) <= (layer0_outputs(7737)) or (layer0_outputs(865));
    outputs(48) <= not((layer0_outputs(3045)) xor (layer0_outputs(3726)));
    outputs(49) <= layer0_outputs(6660);
    outputs(50) <= '1';
    outputs(51) <= not((layer0_outputs(11810)) xor (layer0_outputs(11203)));
    outputs(52) <= not((layer0_outputs(184)) or (layer0_outputs(2319)));
    outputs(53) <= not((layer0_outputs(492)) and (layer0_outputs(7913)));
    outputs(54) <= not(layer0_outputs(1183));
    outputs(55) <= not((layer0_outputs(3658)) xor (layer0_outputs(9081)));
    outputs(56) <= not((layer0_outputs(9230)) and (layer0_outputs(8578)));
    outputs(57) <= not((layer0_outputs(5220)) xor (layer0_outputs(3982)));
    outputs(58) <= (layer0_outputs(11917)) xor (layer0_outputs(7076));
    outputs(59) <= not(layer0_outputs(10755));
    outputs(60) <= not((layer0_outputs(10297)) xor (layer0_outputs(548)));
    outputs(61) <= not(layer0_outputs(5035));
    outputs(62) <= not(layer0_outputs(8184));
    outputs(63) <= not(layer0_outputs(10761));
    outputs(64) <= layer0_outputs(3129);
    outputs(65) <= not(layer0_outputs(11048));
    outputs(66) <= not(layer0_outputs(11313)) or (layer0_outputs(1762));
    outputs(67) <= not(layer0_outputs(8872));
    outputs(68) <= not((layer0_outputs(4961)) or (layer0_outputs(6430)));
    outputs(69) <= layer0_outputs(11811);
    outputs(70) <= (layer0_outputs(12224)) and (layer0_outputs(12600));
    outputs(71) <= (layer0_outputs(11180)) and not (layer0_outputs(9478));
    outputs(72) <= (layer0_outputs(7224)) and (layer0_outputs(11240));
    outputs(73) <= not((layer0_outputs(11832)) or (layer0_outputs(1189)));
    outputs(74) <= layer0_outputs(5438);
    outputs(75) <= not((layer0_outputs(2357)) xor (layer0_outputs(10550)));
    outputs(76) <= not(layer0_outputs(7335));
    outputs(77) <= layer0_outputs(4986);
    outputs(78) <= layer0_outputs(3886);
    outputs(79) <= not(layer0_outputs(9680));
    outputs(80) <= (layer0_outputs(9960)) and (layer0_outputs(829));
    outputs(81) <= (layer0_outputs(7930)) xor (layer0_outputs(9889));
    outputs(82) <= not((layer0_outputs(8059)) xor (layer0_outputs(3630)));
    outputs(83) <= not(layer0_outputs(2075));
    outputs(84) <= (layer0_outputs(3933)) xor (layer0_outputs(11555));
    outputs(85) <= not(layer0_outputs(9058));
    outputs(86) <= (layer0_outputs(8364)) xor (layer0_outputs(10402));
    outputs(87) <= not(layer0_outputs(1685));
    outputs(88) <= not(layer0_outputs(5906));
    outputs(89) <= layer0_outputs(5195);
    outputs(90) <= layer0_outputs(6939);
    outputs(91) <= not(layer0_outputs(8015)) or (layer0_outputs(6528));
    outputs(92) <= not((layer0_outputs(327)) or (layer0_outputs(5758)));
    outputs(93) <= not((layer0_outputs(7815)) and (layer0_outputs(6091)));
    outputs(94) <= layer0_outputs(1067);
    outputs(95) <= not((layer0_outputs(10325)) xor (layer0_outputs(5226)));
    outputs(96) <= (layer0_outputs(773)) and not (layer0_outputs(2466));
    outputs(97) <= layer0_outputs(6762);
    outputs(98) <= (layer0_outputs(3960)) and not (layer0_outputs(8008));
    outputs(99) <= layer0_outputs(10034);
    outputs(100) <= layer0_outputs(5161);
    outputs(101) <= layer0_outputs(12738);
    outputs(102) <= (layer0_outputs(3657)) xor (layer0_outputs(8985));
    outputs(103) <= layer0_outputs(1864);
    outputs(104) <= (layer0_outputs(4174)) and not (layer0_outputs(10520));
    outputs(105) <= layer0_outputs(10726);
    outputs(106) <= (layer0_outputs(8616)) and not (layer0_outputs(2663));
    outputs(107) <= (layer0_outputs(6630)) and not (layer0_outputs(1975));
    outputs(108) <= (layer0_outputs(10972)) and (layer0_outputs(954));
    outputs(109) <= not((layer0_outputs(9976)) xor (layer0_outputs(4667)));
    outputs(110) <= not((layer0_outputs(4075)) or (layer0_outputs(8083)));
    outputs(111) <= layer0_outputs(8780);
    outputs(112) <= layer0_outputs(4393);
    outputs(113) <= layer0_outputs(2932);
    outputs(114) <= not((layer0_outputs(4259)) xor (layer0_outputs(7721)));
    outputs(115) <= not(layer0_outputs(9916)) or (layer0_outputs(580));
    outputs(116) <= not((layer0_outputs(640)) xor (layer0_outputs(8907)));
    outputs(117) <= not(layer0_outputs(9261));
    outputs(118) <= not((layer0_outputs(10799)) and (layer0_outputs(4739)));
    outputs(119) <= not((layer0_outputs(5348)) xor (layer0_outputs(4196)));
    outputs(120) <= '1';
    outputs(121) <= not(layer0_outputs(2080));
    outputs(122) <= not(layer0_outputs(4805));
    outputs(123) <= (layer0_outputs(4125)) and (layer0_outputs(5533));
    outputs(124) <= (layer0_outputs(9026)) and not (layer0_outputs(9012));
    outputs(125) <= (layer0_outputs(10188)) xor (layer0_outputs(4441));
    outputs(126) <= (layer0_outputs(11242)) and not (layer0_outputs(5371));
    outputs(127) <= (layer0_outputs(8310)) and not (layer0_outputs(10202));
    outputs(128) <= layer0_outputs(963);
    outputs(129) <= layer0_outputs(2893);
    outputs(130) <= layer0_outputs(4224);
    outputs(131) <= not(layer0_outputs(4638));
    outputs(132) <= not(layer0_outputs(2693));
    outputs(133) <= layer0_outputs(6493);
    outputs(134) <= (layer0_outputs(3003)) and not (layer0_outputs(6840));
    outputs(135) <= layer0_outputs(5955);
    outputs(136) <= not(layer0_outputs(4655)) or (layer0_outputs(3581));
    outputs(137) <= layer0_outputs(935);
    outputs(138) <= not(layer0_outputs(5824)) or (layer0_outputs(2961));
    outputs(139) <= (layer0_outputs(9865)) and (layer0_outputs(8636));
    outputs(140) <= (layer0_outputs(3191)) and (layer0_outputs(3546));
    outputs(141) <= layer0_outputs(10024);
    outputs(142) <= not((layer0_outputs(4447)) xor (layer0_outputs(6442)));
    outputs(143) <= layer0_outputs(5089);
    outputs(144) <= (layer0_outputs(7616)) or (layer0_outputs(7334));
    outputs(145) <= (layer0_outputs(4203)) xor (layer0_outputs(266));
    outputs(146) <= (layer0_outputs(5215)) and (layer0_outputs(1979));
    outputs(147) <= (layer0_outputs(9607)) xor (layer0_outputs(8873));
    outputs(148) <= not(layer0_outputs(4211)) or (layer0_outputs(2630));
    outputs(149) <= not(layer0_outputs(4289));
    outputs(150) <= not((layer0_outputs(10919)) xor (layer0_outputs(11637)));
    outputs(151) <= (layer0_outputs(218)) and (layer0_outputs(8577));
    outputs(152) <= layer0_outputs(9357);
    outputs(153) <= not((layer0_outputs(3002)) xor (layer0_outputs(6385)));
    outputs(154) <= layer0_outputs(1907);
    outputs(155) <= not(layer0_outputs(6225)) or (layer0_outputs(6139));
    outputs(156) <= (layer0_outputs(8949)) xor (layer0_outputs(5825));
    outputs(157) <= layer0_outputs(4254);
    outputs(158) <= layer0_outputs(1945);
    outputs(159) <= not((layer0_outputs(4560)) and (layer0_outputs(11818)));
    outputs(160) <= (layer0_outputs(12035)) and not (layer0_outputs(11145));
    outputs(161) <= not(layer0_outputs(6570));
    outputs(162) <= not((layer0_outputs(1821)) xor (layer0_outputs(3321)));
    outputs(163) <= layer0_outputs(5204);
    outputs(164) <= not(layer0_outputs(3257));
    outputs(165) <= not(layer0_outputs(4790)) or (layer0_outputs(7803));
    outputs(166) <= layer0_outputs(2595);
    outputs(167) <= (layer0_outputs(2260)) xor (layer0_outputs(5525));
    outputs(168) <= not(layer0_outputs(9118)) or (layer0_outputs(10384));
    outputs(169) <= not(layer0_outputs(7972));
    outputs(170) <= (layer0_outputs(10352)) and not (layer0_outputs(1143));
    outputs(171) <= (layer0_outputs(9967)) xor (layer0_outputs(11505));
    outputs(172) <= not((layer0_outputs(8414)) xor (layer0_outputs(1823)));
    outputs(173) <= not(layer0_outputs(5144));
    outputs(174) <= layer0_outputs(862);
    outputs(175) <= (layer0_outputs(4000)) and not (layer0_outputs(10680));
    outputs(176) <= not((layer0_outputs(1058)) xor (layer0_outputs(10479)));
    outputs(177) <= (layer0_outputs(10163)) xor (layer0_outputs(12029));
    outputs(178) <= (layer0_outputs(6065)) or (layer0_outputs(116));
    outputs(179) <= layer0_outputs(965);
    outputs(180) <= layer0_outputs(3218);
    outputs(181) <= (layer0_outputs(39)) and not (layer0_outputs(6783));
    outputs(182) <= layer0_outputs(12730);
    outputs(183) <= layer0_outputs(2982);
    outputs(184) <= not(layer0_outputs(657));
    outputs(185) <= not(layer0_outputs(10999)) or (layer0_outputs(12036));
    outputs(186) <= layer0_outputs(1026);
    outputs(187) <= (layer0_outputs(3319)) and (layer0_outputs(8303));
    outputs(188) <= not(layer0_outputs(9954));
    outputs(189) <= not(layer0_outputs(5513));
    outputs(190) <= not((layer0_outputs(393)) and (layer0_outputs(1731)));
    outputs(191) <= not((layer0_outputs(12210)) or (layer0_outputs(4189)));
    outputs(192) <= (layer0_outputs(10116)) and not (layer0_outputs(9460));
    outputs(193) <= not((layer0_outputs(8861)) xor (layer0_outputs(1843)));
    outputs(194) <= (layer0_outputs(12207)) xor (layer0_outputs(12247));
    outputs(195) <= not(layer0_outputs(725)) or (layer0_outputs(7511));
    outputs(196) <= not((layer0_outputs(8445)) or (layer0_outputs(4285)));
    outputs(197) <= (layer0_outputs(7520)) and not (layer0_outputs(709));
    outputs(198) <= layer0_outputs(11912);
    outputs(199) <= not(layer0_outputs(1849)) or (layer0_outputs(9625));
    outputs(200) <= not((layer0_outputs(1174)) or (layer0_outputs(4423)));
    outputs(201) <= not(layer0_outputs(1785));
    outputs(202) <= not((layer0_outputs(2898)) xor (layer0_outputs(5703)));
    outputs(203) <= layer0_outputs(8646);
    outputs(204) <= (layer0_outputs(9434)) xor (layer0_outputs(10346));
    outputs(205) <= layer0_outputs(6972);
    outputs(206) <= (layer0_outputs(1784)) and not (layer0_outputs(9015));
    outputs(207) <= not((layer0_outputs(3604)) or (layer0_outputs(54)));
    outputs(208) <= (layer0_outputs(5524)) and not (layer0_outputs(7713));
    outputs(209) <= not((layer0_outputs(9896)) xor (layer0_outputs(9809)));
    outputs(210) <= not((layer0_outputs(5472)) xor (layer0_outputs(5157)));
    outputs(211) <= layer0_outputs(9393);
    outputs(212) <= not(layer0_outputs(6202));
    outputs(213) <= layer0_outputs(146);
    outputs(214) <= not(layer0_outputs(7115));
    outputs(215) <= not(layer0_outputs(11156)) or (layer0_outputs(2518));
    outputs(216) <= not((layer0_outputs(2004)) or (layer0_outputs(4069)));
    outputs(217) <= not(layer0_outputs(6540)) or (layer0_outputs(12334));
    outputs(218) <= (layer0_outputs(4604)) xor (layer0_outputs(8802));
    outputs(219) <= (layer0_outputs(7135)) and not (layer0_outputs(5381));
    outputs(220) <= not(layer0_outputs(9622));
    outputs(221) <= not(layer0_outputs(12179));
    outputs(222) <= (layer0_outputs(11931)) xor (layer0_outputs(8240));
    outputs(223) <= not(layer0_outputs(730));
    outputs(224) <= not((layer0_outputs(531)) and (layer0_outputs(8671)));
    outputs(225) <= not(layer0_outputs(657));
    outputs(226) <= (layer0_outputs(8775)) and not (layer0_outputs(5315));
    outputs(227) <= (layer0_outputs(1778)) and not (layer0_outputs(2342));
    outputs(228) <= not((layer0_outputs(1626)) xor (layer0_outputs(10232)));
    outputs(229) <= (layer0_outputs(9304)) xor (layer0_outputs(11501));
    outputs(230) <= not(layer0_outputs(8258));
    outputs(231) <= layer0_outputs(7066);
    outputs(232) <= not((layer0_outputs(11217)) and (layer0_outputs(11064)));
    outputs(233) <= not(layer0_outputs(1520)) or (layer0_outputs(8560));
    outputs(234) <= layer0_outputs(12791);
    outputs(235) <= (layer0_outputs(2341)) xor (layer0_outputs(10629));
    outputs(236) <= layer0_outputs(1197);
    outputs(237) <= layer0_outputs(4815);
    outputs(238) <= layer0_outputs(7486);
    outputs(239) <= not(layer0_outputs(9293));
    outputs(240) <= (layer0_outputs(11688)) and not (layer0_outputs(6791));
    outputs(241) <= not(layer0_outputs(2510));
    outputs(242) <= layer0_outputs(4295);
    outputs(243) <= not(layer0_outputs(2532));
    outputs(244) <= not((layer0_outputs(12567)) xor (layer0_outputs(965)));
    outputs(245) <= (layer0_outputs(10733)) xor (layer0_outputs(9452));
    outputs(246) <= not(layer0_outputs(5453));
    outputs(247) <= layer0_outputs(4932);
    outputs(248) <= layer0_outputs(10402);
    outputs(249) <= not(layer0_outputs(11143)) or (layer0_outputs(8465));
    outputs(250) <= not((layer0_outputs(7698)) xor (layer0_outputs(5827)));
    outputs(251) <= not(layer0_outputs(8228)) or (layer0_outputs(6885));
    outputs(252) <= (layer0_outputs(8062)) or (layer0_outputs(12727));
    outputs(253) <= (layer0_outputs(8838)) and not (layer0_outputs(3767));
    outputs(254) <= not((layer0_outputs(11790)) xor (layer0_outputs(5783)));
    outputs(255) <= layer0_outputs(5563);
    outputs(256) <= not((layer0_outputs(11895)) xor (layer0_outputs(9524)));
    outputs(257) <= not(layer0_outputs(10455)) or (layer0_outputs(12055));
    outputs(258) <= layer0_outputs(9383);
    outputs(259) <= layer0_outputs(1691);
    outputs(260) <= (layer0_outputs(1228)) xor (layer0_outputs(3126));
    outputs(261) <= not(layer0_outputs(9415));
    outputs(262) <= not((layer0_outputs(8507)) xor (layer0_outputs(7873)));
    outputs(263) <= layer0_outputs(9216);
    outputs(264) <= not(layer0_outputs(11583));
    outputs(265) <= layer0_outputs(8697);
    outputs(266) <= not(layer0_outputs(10490));
    outputs(267) <= not(layer0_outputs(6384));
    outputs(268) <= not(layer0_outputs(7651));
    outputs(269) <= not((layer0_outputs(211)) and (layer0_outputs(11991)));
    outputs(270) <= not((layer0_outputs(12204)) xor (layer0_outputs(7784)));
    outputs(271) <= not((layer0_outputs(2742)) and (layer0_outputs(5265)));
    outputs(272) <= (layer0_outputs(6644)) or (layer0_outputs(9806));
    outputs(273) <= not(layer0_outputs(11856));
    outputs(274) <= layer0_outputs(4107);
    outputs(275) <= layer0_outputs(10797);
    outputs(276) <= (layer0_outputs(11602)) xor (layer0_outputs(5650));
    outputs(277) <= (layer0_outputs(8280)) xor (layer0_outputs(3664));
    outputs(278) <= layer0_outputs(6845);
    outputs(279) <= not((layer0_outputs(11280)) xor (layer0_outputs(10636)));
    outputs(280) <= (layer0_outputs(7309)) and (layer0_outputs(4003));
    outputs(281) <= not(layer0_outputs(9209));
    outputs(282) <= not(layer0_outputs(9460));
    outputs(283) <= (layer0_outputs(7526)) and not (layer0_outputs(9154));
    outputs(284) <= (layer0_outputs(8006)) and not (layer0_outputs(1607));
    outputs(285) <= layer0_outputs(8436);
    outputs(286) <= not((layer0_outputs(6344)) xor (layer0_outputs(2877)));
    outputs(287) <= (layer0_outputs(120)) or (layer0_outputs(74));
    outputs(288) <= (layer0_outputs(10912)) xor (layer0_outputs(2048));
    outputs(289) <= layer0_outputs(2582);
    outputs(290) <= not(layer0_outputs(2814));
    outputs(291) <= not(layer0_outputs(4843)) or (layer0_outputs(2345));
    outputs(292) <= (layer0_outputs(12689)) and not (layer0_outputs(1646));
    outputs(293) <= not(layer0_outputs(5106));
    outputs(294) <= '1';
    outputs(295) <= (layer0_outputs(10101)) xor (layer0_outputs(4187));
    outputs(296) <= not(layer0_outputs(10398));
    outputs(297) <= not(layer0_outputs(1855));
    outputs(298) <= layer0_outputs(2062);
    outputs(299) <= not(layer0_outputs(9984));
    outputs(300) <= not(layer0_outputs(6401));
    outputs(301) <= not((layer0_outputs(5754)) xor (layer0_outputs(10727)));
    outputs(302) <= not((layer0_outputs(1836)) xor (layer0_outputs(3541)));
    outputs(303) <= not((layer0_outputs(4884)) xor (layer0_outputs(10134)));
    outputs(304) <= not(layer0_outputs(5153)) or (layer0_outputs(12590));
    outputs(305) <= layer0_outputs(12206);
    outputs(306) <= layer0_outputs(2892);
    outputs(307) <= not(layer0_outputs(6741));
    outputs(308) <= layer0_outputs(5767);
    outputs(309) <= (layer0_outputs(12463)) xor (layer0_outputs(12604));
    outputs(310) <= layer0_outputs(4479);
    outputs(311) <= not(layer0_outputs(9823));
    outputs(312) <= not(layer0_outputs(8265));
    outputs(313) <= not(layer0_outputs(8551));
    outputs(314) <= not(layer0_outputs(8945));
    outputs(315) <= not(layer0_outputs(6327));
    outputs(316) <= not((layer0_outputs(5004)) and (layer0_outputs(9464)));
    outputs(317) <= not((layer0_outputs(5042)) xor (layer0_outputs(8633)));
    outputs(318) <= not((layer0_outputs(7780)) and (layer0_outputs(11422)));
    outputs(319) <= (layer0_outputs(3758)) or (layer0_outputs(5452));
    outputs(320) <= not(layer0_outputs(1708));
    outputs(321) <= (layer0_outputs(1312)) or (layer0_outputs(7777));
    outputs(322) <= not(layer0_outputs(3352)) or (layer0_outputs(12687));
    outputs(323) <= not((layer0_outputs(2311)) xor (layer0_outputs(7468)));
    outputs(324) <= not(layer0_outputs(10984));
    outputs(325) <= not((layer0_outputs(5527)) or (layer0_outputs(11202)));
    outputs(326) <= not(layer0_outputs(4549));
    outputs(327) <= (layer0_outputs(9465)) and not (layer0_outputs(712));
    outputs(328) <= not((layer0_outputs(11346)) xor (layer0_outputs(7696)));
    outputs(329) <= not((layer0_outputs(1595)) or (layer0_outputs(10370)));
    outputs(330) <= not(layer0_outputs(1496));
    outputs(331) <= (layer0_outputs(3075)) xor (layer0_outputs(6429));
    outputs(332) <= not(layer0_outputs(7817));
    outputs(333) <= layer0_outputs(8544);
    outputs(334) <= layer0_outputs(10349);
    outputs(335) <= layer0_outputs(7345);
    outputs(336) <= not(layer0_outputs(11870)) or (layer0_outputs(11674));
    outputs(337) <= not(layer0_outputs(8290)) or (layer0_outputs(3307));
    outputs(338) <= (layer0_outputs(8975)) xor (layer0_outputs(5360));
    outputs(339) <= layer0_outputs(1902);
    outputs(340) <= layer0_outputs(4976);
    outputs(341) <= layer0_outputs(4922);
    outputs(342) <= (layer0_outputs(3718)) xor (layer0_outputs(6335));
    outputs(343) <= not(layer0_outputs(384));
    outputs(344) <= (layer0_outputs(3009)) and not (layer0_outputs(3715));
    outputs(345) <= not((layer0_outputs(1692)) or (layer0_outputs(6128)));
    outputs(346) <= (layer0_outputs(11433)) and not (layer0_outputs(1761));
    outputs(347) <= not(layer0_outputs(7460)) or (layer0_outputs(12747));
    outputs(348) <= (layer0_outputs(10334)) and (layer0_outputs(3185));
    outputs(349) <= not(layer0_outputs(4527)) or (layer0_outputs(7842));
    outputs(350) <= layer0_outputs(10866);
    outputs(351) <= not(layer0_outputs(2191));
    outputs(352) <= (layer0_outputs(3595)) and not (layer0_outputs(10223));
    outputs(353) <= not((layer0_outputs(7808)) or (layer0_outputs(7684)));
    outputs(354) <= layer0_outputs(5693);
    outputs(355) <= not(layer0_outputs(9577));
    outputs(356) <= not(layer0_outputs(12135)) or (layer0_outputs(10796));
    outputs(357) <= layer0_outputs(9427);
    outputs(358) <= layer0_outputs(3697);
    outputs(359) <= (layer0_outputs(1801)) and not (layer0_outputs(10803));
    outputs(360) <= (layer0_outputs(3941)) and not (layer0_outputs(3521));
    outputs(361) <= not(layer0_outputs(9543)) or (layer0_outputs(11914));
    outputs(362) <= not(layer0_outputs(3551));
    outputs(363) <= not(layer0_outputs(5773));
    outputs(364) <= not((layer0_outputs(10603)) xor (layer0_outputs(5560)));
    outputs(365) <= not(layer0_outputs(10679));
    outputs(366) <= not(layer0_outputs(322)) or (layer0_outputs(1161));
    outputs(367) <= not(layer0_outputs(11184));
    outputs(368) <= (layer0_outputs(8556)) and not (layer0_outputs(11228));
    outputs(369) <= not(layer0_outputs(11879));
    outputs(370) <= not(layer0_outputs(1720));
    outputs(371) <= (layer0_outputs(6289)) xor (layer0_outputs(12550));
    outputs(372) <= (layer0_outputs(253)) or (layer0_outputs(7093));
    outputs(373) <= not(layer0_outputs(6327));
    outputs(374) <= '1';
    outputs(375) <= (layer0_outputs(10)) and not (layer0_outputs(10173));
    outputs(376) <= (layer0_outputs(4030)) and (layer0_outputs(3232));
    outputs(377) <= not(layer0_outputs(5964)) or (layer0_outputs(11980));
    outputs(378) <= layer0_outputs(11423);
    outputs(379) <= not((layer0_outputs(7176)) xor (layer0_outputs(12580)));
    outputs(380) <= not(layer0_outputs(6078));
    outputs(381) <= (layer0_outputs(5482)) or (layer0_outputs(1599));
    outputs(382) <= layer0_outputs(2514);
    outputs(383) <= layer0_outputs(11487);
    outputs(384) <= (layer0_outputs(12789)) and (layer0_outputs(7032));
    outputs(385) <= not(layer0_outputs(11440));
    outputs(386) <= not(layer0_outputs(3812));
    outputs(387) <= (layer0_outputs(2748)) and not (layer0_outputs(2440));
    outputs(388) <= not(layer0_outputs(10927));
    outputs(389) <= (layer0_outputs(707)) and not (layer0_outputs(7715));
    outputs(390) <= not(layer0_outputs(10835));
    outputs(391) <= (layer0_outputs(9504)) xor (layer0_outputs(2547));
    outputs(392) <= not(layer0_outputs(5229));
    outputs(393) <= not(layer0_outputs(7409));
    outputs(394) <= (layer0_outputs(7831)) and (layer0_outputs(6785));
    outputs(395) <= (layer0_outputs(2114)) xor (layer0_outputs(10869));
    outputs(396) <= not(layer0_outputs(759));
    outputs(397) <= not((layer0_outputs(3306)) xor (layer0_outputs(7770)));
    outputs(398) <= layer0_outputs(3395);
    outputs(399) <= not(layer0_outputs(12588));
    outputs(400) <= not((layer0_outputs(1835)) xor (layer0_outputs(813)));
    outputs(401) <= layer0_outputs(4766);
    outputs(402) <= layer0_outputs(10390);
    outputs(403) <= (layer0_outputs(4662)) and not (layer0_outputs(3414));
    outputs(404) <= layer0_outputs(321);
    outputs(405) <= not((layer0_outputs(3990)) or (layer0_outputs(5782)));
    outputs(406) <= not(layer0_outputs(10018));
    outputs(407) <= not(layer0_outputs(583)) or (layer0_outputs(1657));
    outputs(408) <= (layer0_outputs(11101)) xor (layer0_outputs(10630));
    outputs(409) <= not(layer0_outputs(11298));
    outputs(410) <= not((layer0_outputs(224)) xor (layer0_outputs(8005)));
    outputs(411) <= (layer0_outputs(433)) xor (layer0_outputs(2443));
    outputs(412) <= layer0_outputs(1702);
    outputs(413) <= not((layer0_outputs(3925)) xor (layer0_outputs(11720)));
    outputs(414) <= not(layer0_outputs(435)) or (layer0_outputs(3583));
    outputs(415) <= (layer0_outputs(320)) and not (layer0_outputs(5081));
    outputs(416) <= not(layer0_outputs(12171));
    outputs(417) <= not(layer0_outputs(122));
    outputs(418) <= (layer0_outputs(12204)) and not (layer0_outputs(10785));
    outputs(419) <= (layer0_outputs(6004)) and (layer0_outputs(10216));
    outputs(420) <= not(layer0_outputs(7540));
    outputs(421) <= layer0_outputs(4636);
    outputs(422) <= (layer0_outputs(7988)) or (layer0_outputs(8948));
    outputs(423) <= not((layer0_outputs(4104)) xor (layer0_outputs(701)));
    outputs(424) <= not(layer0_outputs(3991));
    outputs(425) <= not(layer0_outputs(3133));
    outputs(426) <= layer0_outputs(11386);
    outputs(427) <= not(layer0_outputs(8496));
    outputs(428) <= layer0_outputs(8807);
    outputs(429) <= not(layer0_outputs(1950));
    outputs(430) <= (layer0_outputs(6837)) and (layer0_outputs(10692));
    outputs(431) <= (layer0_outputs(727)) and (layer0_outputs(11022));
    outputs(432) <= not((layer0_outputs(7809)) xor (layer0_outputs(9990)));
    outputs(433) <= layer0_outputs(401);
    outputs(434) <= not(layer0_outputs(5006));
    outputs(435) <= (layer0_outputs(1520)) xor (layer0_outputs(8626));
    outputs(436) <= not(layer0_outputs(9085));
    outputs(437) <= not(layer0_outputs(9839)) or (layer0_outputs(4162));
    outputs(438) <= not((layer0_outputs(12682)) xor (layer0_outputs(5888)));
    outputs(439) <= (layer0_outputs(337)) xor (layer0_outputs(3762));
    outputs(440) <= layer0_outputs(12401);
    outputs(441) <= layer0_outputs(4067);
    outputs(442) <= not((layer0_outputs(5600)) xor (layer0_outputs(6018)));
    outputs(443) <= layer0_outputs(6305);
    outputs(444) <= (layer0_outputs(370)) xor (layer0_outputs(8104));
    outputs(445) <= not(layer0_outputs(2918));
    outputs(446) <= not((layer0_outputs(10324)) xor (layer0_outputs(2585)));
    outputs(447) <= layer0_outputs(5975);
    outputs(448) <= layer0_outputs(8014);
    outputs(449) <= (layer0_outputs(3210)) xor (layer0_outputs(1795));
    outputs(450) <= not((layer0_outputs(1875)) and (layer0_outputs(9244)));
    outputs(451) <= (layer0_outputs(417)) or (layer0_outputs(6806));
    outputs(452) <= not(layer0_outputs(9278));
    outputs(453) <= (layer0_outputs(8315)) and not (layer0_outputs(5564));
    outputs(454) <= (layer0_outputs(12439)) xor (layer0_outputs(5507));
    outputs(455) <= not((layer0_outputs(11705)) and (layer0_outputs(5901)));
    outputs(456) <= not(layer0_outputs(3095));
    outputs(457) <= (layer0_outputs(2099)) and (layer0_outputs(7284));
    outputs(458) <= layer0_outputs(6150);
    outputs(459) <= layer0_outputs(4052);
    outputs(460) <= not(layer0_outputs(5402));
    outputs(461) <= layer0_outputs(697);
    outputs(462) <= not((layer0_outputs(11459)) xor (layer0_outputs(7594)));
    outputs(463) <= not((layer0_outputs(5461)) or (layer0_outputs(3616)));
    outputs(464) <= (layer0_outputs(10669)) xor (layer0_outputs(3562));
    outputs(465) <= (layer0_outputs(8247)) or (layer0_outputs(44));
    outputs(466) <= layer0_outputs(3069);
    outputs(467) <= not(layer0_outputs(7702));
    outputs(468) <= not((layer0_outputs(9309)) or (layer0_outputs(11498)));
    outputs(469) <= not((layer0_outputs(10077)) xor (layer0_outputs(12141)));
    outputs(470) <= layer0_outputs(2828);
    outputs(471) <= layer0_outputs(1905);
    outputs(472) <= layer0_outputs(9076);
    outputs(473) <= (layer0_outputs(11279)) or (layer0_outputs(12721));
    outputs(474) <= (layer0_outputs(5218)) xor (layer0_outputs(3032));
    outputs(475) <= not(layer0_outputs(9775));
    outputs(476) <= layer0_outputs(7451);
    outputs(477) <= not((layer0_outputs(7989)) or (layer0_outputs(11249)));
    outputs(478) <= not(layer0_outputs(12196));
    outputs(479) <= not(layer0_outputs(8137)) or (layer0_outputs(3657));
    outputs(480) <= not((layer0_outputs(7440)) xor (layer0_outputs(6634)));
    outputs(481) <= (layer0_outputs(3154)) and not (layer0_outputs(8841));
    outputs(482) <= (layer0_outputs(12012)) or (layer0_outputs(2126));
    outputs(483) <= not(layer0_outputs(4861));
    outputs(484) <= layer0_outputs(6526);
    outputs(485) <= not((layer0_outputs(7399)) and (layer0_outputs(3718)));
    outputs(486) <= layer0_outputs(10209);
    outputs(487) <= not(layer0_outputs(446));
    outputs(488) <= (layer0_outputs(7629)) and (layer0_outputs(7361));
    outputs(489) <= (layer0_outputs(7143)) xor (layer0_outputs(4121));
    outputs(490) <= layer0_outputs(185);
    outputs(491) <= '1';
    outputs(492) <= not(layer0_outputs(6703)) or (layer0_outputs(8209));
    outputs(493) <= (layer0_outputs(6746)) and (layer0_outputs(182));
    outputs(494) <= not(layer0_outputs(11691));
    outputs(495) <= layer0_outputs(2617);
    outputs(496) <= layer0_outputs(11629);
    outputs(497) <= not((layer0_outputs(468)) or (layer0_outputs(1015)));
    outputs(498) <= not(layer0_outputs(3588));
    outputs(499) <= not(layer0_outputs(6670));
    outputs(500) <= (layer0_outputs(1519)) xor (layer0_outputs(140));
    outputs(501) <= layer0_outputs(11096);
    outputs(502) <= not((layer0_outputs(12797)) xor (layer0_outputs(1903)));
    outputs(503) <= not((layer0_outputs(3686)) xor (layer0_outputs(9268)));
    outputs(504) <= layer0_outputs(3751);
    outputs(505) <= not(layer0_outputs(6654)) or (layer0_outputs(12745));
    outputs(506) <= not(layer0_outputs(7727));
    outputs(507) <= not((layer0_outputs(10529)) xor (layer0_outputs(5985)));
    outputs(508) <= not(layer0_outputs(10932));
    outputs(509) <= layer0_outputs(7094);
    outputs(510) <= layer0_outputs(6019);
    outputs(511) <= layer0_outputs(2298);
    outputs(512) <= not(layer0_outputs(2708));
    outputs(513) <= layer0_outputs(454);
    outputs(514) <= (layer0_outputs(8999)) and not (layer0_outputs(5933));
    outputs(515) <= (layer0_outputs(6767)) xor (layer0_outputs(10339));
    outputs(516) <= (layer0_outputs(6030)) xor (layer0_outputs(7349));
    outputs(517) <= (layer0_outputs(8975)) xor (layer0_outputs(12654));
    outputs(518) <= not((layer0_outputs(413)) xor (layer0_outputs(4735)));
    outputs(519) <= (layer0_outputs(1688)) or (layer0_outputs(5383));
    outputs(520) <= layer0_outputs(11193);
    outputs(521) <= not((layer0_outputs(5485)) or (layer0_outputs(12111)));
    outputs(522) <= not(layer0_outputs(5646)) or (layer0_outputs(4837));
    outputs(523) <= (layer0_outputs(3936)) and (layer0_outputs(6182));
    outputs(524) <= not(layer0_outputs(2618));
    outputs(525) <= not((layer0_outputs(5464)) xor (layer0_outputs(6074)));
    outputs(526) <= not(layer0_outputs(8262));
    outputs(527) <= not((layer0_outputs(6986)) xor (layer0_outputs(9276)));
    outputs(528) <= not(layer0_outputs(2424)) or (layer0_outputs(6619));
    outputs(529) <= (layer0_outputs(63)) and (layer0_outputs(2287));
    outputs(530) <= not((layer0_outputs(9671)) and (layer0_outputs(9315)));
    outputs(531) <= (layer0_outputs(3222)) xor (layer0_outputs(8826));
    outputs(532) <= (layer0_outputs(2855)) xor (layer0_outputs(4521));
    outputs(533) <= (layer0_outputs(12405)) and not (layer0_outputs(4009));
    outputs(534) <= not((layer0_outputs(1518)) or (layer0_outputs(9703)));
    outputs(535) <= not(layer0_outputs(4523));
    outputs(536) <= (layer0_outputs(1138)) and not (layer0_outputs(11387));
    outputs(537) <= not(layer0_outputs(7865));
    outputs(538) <= layer0_outputs(2150);
    outputs(539) <= layer0_outputs(12217);
    outputs(540) <= layer0_outputs(3769);
    outputs(541) <= not(layer0_outputs(11813));
    outputs(542) <= layer0_outputs(9087);
    outputs(543) <= (layer0_outputs(3756)) and not (layer0_outputs(11228));
    outputs(544) <= not(layer0_outputs(5864));
    outputs(545) <= layer0_outputs(9589);
    outputs(546) <= layer0_outputs(7868);
    outputs(547) <= (layer0_outputs(2553)) xor (layer0_outputs(11541));
    outputs(548) <= (layer0_outputs(6411)) and (layer0_outputs(7071));
    outputs(549) <= (layer0_outputs(11079)) xor (layer0_outputs(12029));
    outputs(550) <= layer0_outputs(10167);
    outputs(551) <= layer0_outputs(519);
    outputs(552) <= not((layer0_outputs(3008)) xor (layer0_outputs(3583)));
    outputs(553) <= (layer0_outputs(7971)) xor (layer0_outputs(10372));
    outputs(554) <= not((layer0_outputs(8491)) xor (layer0_outputs(8771)));
    outputs(555) <= (layer0_outputs(1955)) xor (layer0_outputs(6287));
    outputs(556) <= layer0_outputs(7098);
    outputs(557) <= not((layer0_outputs(6685)) or (layer0_outputs(1053)));
    outputs(558) <= not((layer0_outputs(11077)) and (layer0_outputs(2079)));
    outputs(559) <= not((layer0_outputs(3780)) xor (layer0_outputs(10270)));
    outputs(560) <= not(layer0_outputs(6896));
    outputs(561) <= not((layer0_outputs(12778)) or (layer0_outputs(12430)));
    outputs(562) <= (layer0_outputs(4885)) and not (layer0_outputs(992));
    outputs(563) <= not((layer0_outputs(2753)) and (layer0_outputs(3342)));
    outputs(564) <= (layer0_outputs(7319)) xor (layer0_outputs(11042));
    outputs(565) <= (layer0_outputs(2856)) and (layer0_outputs(10378));
    outputs(566) <= layer0_outputs(12177);
    outputs(567) <= not(layer0_outputs(11048));
    outputs(568) <= not((layer0_outputs(6135)) xor (layer0_outputs(4286)));
    outputs(569) <= (layer0_outputs(11140)) or (layer0_outputs(6192));
    outputs(570) <= not(layer0_outputs(101));
    outputs(571) <= not((layer0_outputs(6882)) xor (layer0_outputs(5051)));
    outputs(572) <= (layer0_outputs(5598)) xor (layer0_outputs(1182));
    outputs(573) <= not((layer0_outputs(5747)) xor (layer0_outputs(3906)));
    outputs(574) <= not((layer0_outputs(3418)) xor (layer0_outputs(8345)));
    outputs(575) <= not(layer0_outputs(2470)) or (layer0_outputs(12526));
    outputs(576) <= not(layer0_outputs(10835)) or (layer0_outputs(5445));
    outputs(577) <= not(layer0_outputs(1428));
    outputs(578) <= (layer0_outputs(4792)) and (layer0_outputs(750));
    outputs(579) <= (layer0_outputs(4574)) xor (layer0_outputs(3404));
    outputs(580) <= (layer0_outputs(3149)) xor (layer0_outputs(2565));
    outputs(581) <= (layer0_outputs(11685)) xor (layer0_outputs(12156));
    outputs(582) <= not(layer0_outputs(8200));
    outputs(583) <= not((layer0_outputs(7559)) or (layer0_outputs(445)));
    outputs(584) <= (layer0_outputs(11784)) xor (layer0_outputs(2216));
    outputs(585) <= layer0_outputs(7108);
    outputs(586) <= (layer0_outputs(16)) or (layer0_outputs(4121));
    outputs(587) <= (layer0_outputs(381)) xor (layer0_outputs(8247));
    outputs(588) <= (layer0_outputs(5908)) and not (layer0_outputs(7177));
    outputs(589) <= not(layer0_outputs(3141));
    outputs(590) <= (layer0_outputs(2362)) and (layer0_outputs(10300));
    outputs(591) <= layer0_outputs(6440);
    outputs(592) <= not(layer0_outputs(11788));
    outputs(593) <= not(layer0_outputs(3055));
    outputs(594) <= not(layer0_outputs(3731));
    outputs(595) <= not((layer0_outputs(6918)) xor (layer0_outputs(6228)));
    outputs(596) <= not(layer0_outputs(7546));
    outputs(597) <= not((layer0_outputs(4192)) or (layer0_outputs(4763)));
    outputs(598) <= layer0_outputs(3152);
    outputs(599) <= not((layer0_outputs(12614)) xor (layer0_outputs(8440)));
    outputs(600) <= not(layer0_outputs(8947));
    outputs(601) <= not(layer0_outputs(5994));
    outputs(602) <= not((layer0_outputs(8814)) xor (layer0_outputs(3249)));
    outputs(603) <= not(layer0_outputs(2700));
    outputs(604) <= not(layer0_outputs(2839));
    outputs(605) <= layer0_outputs(881);
    outputs(606) <= not(layer0_outputs(1370));
    outputs(607) <= (layer0_outputs(1180)) and not (layer0_outputs(398));
    outputs(608) <= (layer0_outputs(1299)) and not (layer0_outputs(7355));
    outputs(609) <= layer0_outputs(11153);
    outputs(610) <= not((layer0_outputs(7086)) xor (layer0_outputs(4532)));
    outputs(611) <= layer0_outputs(8113);
    outputs(612) <= layer0_outputs(2329);
    outputs(613) <= (layer0_outputs(152)) xor (layer0_outputs(4956));
    outputs(614) <= not(layer0_outputs(12278));
    outputs(615) <= layer0_outputs(10565);
    outputs(616) <= not(layer0_outputs(6457)) or (layer0_outputs(4215));
    outputs(617) <= not((layer0_outputs(2073)) xor (layer0_outputs(12239)));
    outputs(618) <= (layer0_outputs(6964)) and (layer0_outputs(12301));
    outputs(619) <= (layer0_outputs(1666)) xor (layer0_outputs(5200));
    outputs(620) <= layer0_outputs(8134);
    outputs(621) <= not(layer0_outputs(5362));
    outputs(622) <= (layer0_outputs(2729)) and not (layer0_outputs(3873));
    outputs(623) <= (layer0_outputs(11072)) and (layer0_outputs(6482));
    outputs(624) <= not((layer0_outputs(1640)) or (layer0_outputs(176)));
    outputs(625) <= (layer0_outputs(1170)) xor (layer0_outputs(12383));
    outputs(626) <= layer0_outputs(11950);
    outputs(627) <= not(layer0_outputs(10293));
    outputs(628) <= (layer0_outputs(9116)) and not (layer0_outputs(3827));
    outputs(629) <= layer0_outputs(7941);
    outputs(630) <= not(layer0_outputs(10564));
    outputs(631) <= (layer0_outputs(125)) xor (layer0_outputs(1780));
    outputs(632) <= layer0_outputs(8100);
    outputs(633) <= (layer0_outputs(7899)) or (layer0_outputs(6087));
    outputs(634) <= not(layer0_outputs(12752));
    outputs(635) <= not(layer0_outputs(3553));
    outputs(636) <= '1';
    outputs(637) <= layer0_outputs(9603);
    outputs(638) <= layer0_outputs(922);
    outputs(639) <= layer0_outputs(10728);
    outputs(640) <= layer0_outputs(4620);
    outputs(641) <= not(layer0_outputs(2449));
    outputs(642) <= (layer0_outputs(858)) xor (layer0_outputs(5795));
    outputs(643) <= (layer0_outputs(8875)) xor (layer0_outputs(11211));
    outputs(644) <= (layer0_outputs(476)) xor (layer0_outputs(639));
    outputs(645) <= not(layer0_outputs(1266));
    outputs(646) <= '1';
    outputs(647) <= not(layer0_outputs(10739));
    outputs(648) <= not(layer0_outputs(7562));
    outputs(649) <= (layer0_outputs(7741)) xor (layer0_outputs(11103));
    outputs(650) <= (layer0_outputs(4748)) and (layer0_outputs(4342));
    outputs(651) <= not(layer0_outputs(9095));
    outputs(652) <= not(layer0_outputs(1619));
    outputs(653) <= layer0_outputs(4209);
    outputs(654) <= (layer0_outputs(225)) xor (layer0_outputs(852));
    outputs(655) <= (layer0_outputs(9093)) and not (layer0_outputs(10912));
    outputs(656) <= not(layer0_outputs(11287)) or (layer0_outputs(7466));
    outputs(657) <= not((layer0_outputs(5175)) and (layer0_outputs(6709)));
    outputs(658) <= layer0_outputs(10917);
    outputs(659) <= not((layer0_outputs(9301)) xor (layer0_outputs(8358)));
    outputs(660) <= not(layer0_outputs(4742)) or (layer0_outputs(10785));
    outputs(661) <= (layer0_outputs(3478)) and not (layer0_outputs(10830));
    outputs(662) <= (layer0_outputs(8092)) xor (layer0_outputs(1440));
    outputs(663) <= not(layer0_outputs(3956));
    outputs(664) <= not((layer0_outputs(12750)) xor (layer0_outputs(6356)));
    outputs(665) <= (layer0_outputs(11392)) and not (layer0_outputs(1746));
    outputs(666) <= (layer0_outputs(11942)) and (layer0_outputs(11945));
    outputs(667) <= layer0_outputs(5411);
    outputs(668) <= not((layer0_outputs(12456)) xor (layer0_outputs(7315)));
    outputs(669) <= (layer0_outputs(7881)) xor (layer0_outputs(3612));
    outputs(670) <= not(layer0_outputs(4782));
    outputs(671) <= not((layer0_outputs(1431)) xor (layer0_outputs(12276)));
    outputs(672) <= (layer0_outputs(11663)) and not (layer0_outputs(882));
    outputs(673) <= not(layer0_outputs(8683)) or (layer0_outputs(5570));
    outputs(674) <= layer0_outputs(3309);
    outputs(675) <= layer0_outputs(4759);
    outputs(676) <= (layer0_outputs(845)) or (layer0_outputs(6128));
    outputs(677) <= layer0_outputs(4076);
    outputs(678) <= (layer0_outputs(7755)) and (layer0_outputs(11568));
    outputs(679) <= not((layer0_outputs(1192)) xor (layer0_outputs(416)));
    outputs(680) <= (layer0_outputs(4151)) or (layer0_outputs(3343));
    outputs(681) <= not(layer0_outputs(6525));
    outputs(682) <= not(layer0_outputs(10653));
    outputs(683) <= not(layer0_outputs(1127));
    outputs(684) <= not((layer0_outputs(9456)) and (layer0_outputs(3885)));
    outputs(685) <= not((layer0_outputs(7008)) and (layer0_outputs(5418)));
    outputs(686) <= not(layer0_outputs(5523));
    outputs(687) <= not((layer0_outputs(8063)) xor (layer0_outputs(4213)));
    outputs(688) <= not(layer0_outputs(4658));
    outputs(689) <= (layer0_outputs(7947)) xor (layer0_outputs(11954));
    outputs(690) <= (layer0_outputs(3441)) or (layer0_outputs(8032));
    outputs(691) <= not((layer0_outputs(1739)) and (layer0_outputs(6127)));
    outputs(692) <= layer0_outputs(1721);
    outputs(693) <= (layer0_outputs(10290)) and (layer0_outputs(12388));
    outputs(694) <= not(layer0_outputs(5178)) or (layer0_outputs(8451));
    outputs(695) <= (layer0_outputs(8282)) xor (layer0_outputs(9581));
    outputs(696) <= not((layer0_outputs(3924)) xor (layer0_outputs(12399)));
    outputs(697) <= not(layer0_outputs(2960));
    outputs(698) <= not(layer0_outputs(12425));
    outputs(699) <= not(layer0_outputs(3964));
    outputs(700) <= layer0_outputs(5441);
    outputs(701) <= not(layer0_outputs(1303)) or (layer0_outputs(8005));
    outputs(702) <= not((layer0_outputs(11948)) xor (layer0_outputs(5605)));
    outputs(703) <= not(layer0_outputs(11329)) or (layer0_outputs(10556));
    outputs(704) <= not(layer0_outputs(7285));
    outputs(705) <= layer0_outputs(4161);
    outputs(706) <= not((layer0_outputs(4411)) or (layer0_outputs(10937)));
    outputs(707) <= not((layer0_outputs(8855)) xor (layer0_outputs(10168)));
    outputs(708) <= not(layer0_outputs(7869));
    outputs(709) <= not(layer0_outputs(10694));
    outputs(710) <= not((layer0_outputs(1475)) xor (layer0_outputs(5674)));
    outputs(711) <= (layer0_outputs(10628)) xor (layer0_outputs(4941));
    outputs(712) <= not((layer0_outputs(12311)) xor (layer0_outputs(7194)));
    outputs(713) <= layer0_outputs(7609);
    outputs(714) <= layer0_outputs(7472);
    outputs(715) <= (layer0_outputs(11291)) and not (layer0_outputs(5345));
    outputs(716) <= (layer0_outputs(2659)) and not (layer0_outputs(10459));
    outputs(717) <= (layer0_outputs(10171)) xor (layer0_outputs(1701));
    outputs(718) <= layer0_outputs(8961);
    outputs(719) <= (layer0_outputs(10719)) and not (layer0_outputs(2240));
    outputs(720) <= (layer0_outputs(12517)) xor (layer0_outputs(11978));
    outputs(721) <= layer0_outputs(5913);
    outputs(722) <= not((layer0_outputs(463)) xor (layer0_outputs(11010)));
    outputs(723) <= layer0_outputs(11843);
    outputs(724) <= layer0_outputs(135);
    outputs(725) <= not((layer0_outputs(2022)) or (layer0_outputs(7344)));
    outputs(726) <= not(layer0_outputs(9550));
    outputs(727) <= not((layer0_outputs(11049)) and (layer0_outputs(6841)));
    outputs(728) <= (layer0_outputs(9534)) xor (layer0_outputs(1766));
    outputs(729) <= (layer0_outputs(1938)) and not (layer0_outputs(11954));
    outputs(730) <= not(layer0_outputs(7693));
    outputs(731) <= not(layer0_outputs(9596));
    outputs(732) <= not((layer0_outputs(11162)) or (layer0_outputs(7190)));
    outputs(733) <= (layer0_outputs(4927)) and (layer0_outputs(10045));
    outputs(734) <= layer0_outputs(7729);
    outputs(735) <= layer0_outputs(8849);
    outputs(736) <= (layer0_outputs(7291)) or (layer0_outputs(7894));
    outputs(737) <= not(layer0_outputs(8163));
    outputs(738) <= layer0_outputs(7557);
    outputs(739) <= layer0_outputs(317);
    outputs(740) <= (layer0_outputs(1834)) xor (layer0_outputs(2338));
    outputs(741) <= not((layer0_outputs(10453)) xor (layer0_outputs(1454)));
    outputs(742) <= not(layer0_outputs(4450));
    outputs(743) <= layer0_outputs(3335);
    outputs(744) <= layer0_outputs(1831);
    outputs(745) <= layer0_outputs(5801);
    outputs(746) <= not((layer0_outputs(6149)) xor (layer0_outputs(11474)));
    outputs(747) <= layer0_outputs(11959);
    outputs(748) <= not(layer0_outputs(8749));
    outputs(749) <= layer0_outputs(10080);
    outputs(750) <= (layer0_outputs(4063)) and not (layer0_outputs(10019));
    outputs(751) <= not(layer0_outputs(9961)) or (layer0_outputs(6219));
    outputs(752) <= not((layer0_outputs(1055)) and (layer0_outputs(6259)));
    outputs(753) <= not(layer0_outputs(9364)) or (layer0_outputs(6970));
    outputs(754) <= not((layer0_outputs(11625)) or (layer0_outputs(7198)));
    outputs(755) <= not((layer0_outputs(2044)) xor (layer0_outputs(11091)));
    outputs(756) <= layer0_outputs(10285);
    outputs(757) <= layer0_outputs(1262);
    outputs(758) <= not((layer0_outputs(8109)) and (layer0_outputs(9302)));
    outputs(759) <= (layer0_outputs(6100)) and not (layer0_outputs(6717));
    outputs(760) <= layer0_outputs(348);
    outputs(761) <= not(layer0_outputs(506));
    outputs(762) <= not(layer0_outputs(11094));
    outputs(763) <= not(layer0_outputs(397)) or (layer0_outputs(1430));
    outputs(764) <= (layer0_outputs(1178)) or (layer0_outputs(7413));
    outputs(765) <= (layer0_outputs(7986)) xor (layer0_outputs(7401));
    outputs(766) <= layer0_outputs(5076);
    outputs(767) <= not(layer0_outputs(4475));
    outputs(768) <= layer0_outputs(12236);
    outputs(769) <= (layer0_outputs(6586)) and not (layer0_outputs(3573));
    outputs(770) <= layer0_outputs(12726);
    outputs(771) <= layer0_outputs(11774);
    outputs(772) <= not(layer0_outputs(3830)) or (layer0_outputs(3893));
    outputs(773) <= not(layer0_outputs(5980)) or (layer0_outputs(7404));
    outputs(774) <= layer0_outputs(9969);
    outputs(775) <= not((layer0_outputs(9913)) or (layer0_outputs(6068)));
    outputs(776) <= not((layer0_outputs(4147)) or (layer0_outputs(2634)));
    outputs(777) <= not(layer0_outputs(11851));
    outputs(778) <= not((layer0_outputs(3031)) xor (layer0_outputs(10907)));
    outputs(779) <= layer0_outputs(11434);
    outputs(780) <= (layer0_outputs(8083)) or (layer0_outputs(6636));
    outputs(781) <= not(layer0_outputs(11217));
    outputs(782) <= (layer0_outputs(12404)) and not (layer0_outputs(4001));
    outputs(783) <= not((layer0_outputs(11762)) xor (layer0_outputs(7849)));
    outputs(784) <= not(layer0_outputs(8238)) or (layer0_outputs(10540));
    outputs(785) <= not(layer0_outputs(4806));
    outputs(786) <= (layer0_outputs(9567)) and not (layer0_outputs(173));
    outputs(787) <= (layer0_outputs(5789)) or (layer0_outputs(12136));
    outputs(788) <= not(layer0_outputs(9397));
    outputs(789) <= not((layer0_outputs(1068)) xor (layer0_outputs(5618)));
    outputs(790) <= (layer0_outputs(9560)) xor (layer0_outputs(4397));
    outputs(791) <= not(layer0_outputs(7052));
    outputs(792) <= not(layer0_outputs(9371)) or (layer0_outputs(10721));
    outputs(793) <= (layer0_outputs(11616)) and (layer0_outputs(3660));
    outputs(794) <= (layer0_outputs(5031)) and not (layer0_outputs(35));
    outputs(795) <= not((layer0_outputs(5894)) xor (layer0_outputs(12281)));
    outputs(796) <= not(layer0_outputs(10313)) or (layer0_outputs(7342));
    outputs(797) <= not(layer0_outputs(5657)) or (layer0_outputs(6529));
    outputs(798) <= (layer0_outputs(6253)) xor (layer0_outputs(359));
    outputs(799) <= not(layer0_outputs(442));
    outputs(800) <= layer0_outputs(10442);
    outputs(801) <= not(layer0_outputs(3610)) or (layer0_outputs(2473));
    outputs(802) <= (layer0_outputs(8023)) and not (layer0_outputs(3535));
    outputs(803) <= not(layer0_outputs(595));
    outputs(804) <= (layer0_outputs(7407)) xor (layer0_outputs(7197));
    outputs(805) <= (layer0_outputs(3742)) xor (layer0_outputs(1579));
    outputs(806) <= not(layer0_outputs(1172));
    outputs(807) <= not(layer0_outputs(6706));
    outputs(808) <= not(layer0_outputs(3879));
    outputs(809) <= not((layer0_outputs(3512)) xor (layer0_outputs(5239)));
    outputs(810) <= (layer0_outputs(10)) and not (layer0_outputs(8682));
    outputs(811) <= not((layer0_outputs(6237)) xor (layer0_outputs(7898)));
    outputs(812) <= not(layer0_outputs(11001));
    outputs(813) <= (layer0_outputs(9806)) and (layer0_outputs(8710));
    outputs(814) <= (layer0_outputs(7968)) xor (layer0_outputs(1248));
    outputs(815) <= layer0_outputs(2377);
    outputs(816) <= not(layer0_outputs(6099));
    outputs(817) <= not(layer0_outputs(11634)) or (layer0_outputs(2575));
    outputs(818) <= not(layer0_outputs(10707));
    outputs(819) <= layer0_outputs(199);
    outputs(820) <= not(layer0_outputs(11025)) or (layer0_outputs(4635));
    outputs(821) <= not(layer0_outputs(1405));
    outputs(822) <= layer0_outputs(2762);
    outputs(823) <= (layer0_outputs(8232)) xor (layer0_outputs(10033));
    outputs(824) <= not(layer0_outputs(10214));
    outputs(825) <= (layer0_outputs(11962)) or (layer0_outputs(3967));
    outputs(826) <= (layer0_outputs(4819)) or (layer0_outputs(7386));
    outputs(827) <= (layer0_outputs(922)) and not (layer0_outputs(9353));
    outputs(828) <= (layer0_outputs(4746)) and not (layer0_outputs(8126));
    outputs(829) <= (layer0_outputs(9552)) and (layer0_outputs(2275));
    outputs(830) <= not(layer0_outputs(12713));
    outputs(831) <= (layer0_outputs(4564)) xor (layer0_outputs(10333));
    outputs(832) <= layer0_outputs(9056);
    outputs(833) <= not(layer0_outputs(842));
    outputs(834) <= (layer0_outputs(11015)) xor (layer0_outputs(6464));
    outputs(835) <= (layer0_outputs(10702)) and (layer0_outputs(12332));
    outputs(836) <= layer0_outputs(6221);
    outputs(837) <= not(layer0_outputs(11680)) or (layer0_outputs(10341));
    outputs(838) <= not(layer0_outputs(9620)) or (layer0_outputs(4150));
    outputs(839) <= not(layer0_outputs(5579));
    outputs(840) <= layer0_outputs(5769);
    outputs(841) <= (layer0_outputs(3869)) and (layer0_outputs(11892));
    outputs(842) <= (layer0_outputs(410)) xor (layer0_outputs(9725));
    outputs(843) <= (layer0_outputs(5760)) xor (layer0_outputs(8073));
    outputs(844) <= not(layer0_outputs(9689));
    outputs(845) <= not(layer0_outputs(5144));
    outputs(846) <= (layer0_outputs(3294)) and not (layer0_outputs(7431));
    outputs(847) <= layer0_outputs(9807);
    outputs(848) <= (layer0_outputs(6877)) xor (layer0_outputs(8183));
    outputs(849) <= layer0_outputs(4591);
    outputs(850) <= not(layer0_outputs(2584));
    outputs(851) <= not((layer0_outputs(3641)) and (layer0_outputs(1632)));
    outputs(852) <= layer0_outputs(1359);
    outputs(853) <= (layer0_outputs(11087)) and (layer0_outputs(9940));
    outputs(854) <= layer0_outputs(7543);
    outputs(855) <= (layer0_outputs(1030)) xor (layer0_outputs(11457));
    outputs(856) <= not(layer0_outputs(7039)) or (layer0_outputs(9234));
    outputs(857) <= layer0_outputs(4832);
    outputs(858) <= (layer0_outputs(4314)) xor (layer0_outputs(3302));
    outputs(859) <= not((layer0_outputs(4953)) or (layer0_outputs(5591)));
    outputs(860) <= not((layer0_outputs(11722)) xor (layer0_outputs(10445)));
    outputs(861) <= (layer0_outputs(8802)) xor (layer0_outputs(4723));
    outputs(862) <= not(layer0_outputs(11878));
    outputs(863) <= (layer0_outputs(2717)) and not (layer0_outputs(12515));
    outputs(864) <= not(layer0_outputs(10270));
    outputs(865) <= layer0_outputs(1412);
    outputs(866) <= not((layer0_outputs(4735)) xor (layer0_outputs(7475)));
    outputs(867) <= (layer0_outputs(11462)) and not (layer0_outputs(10084));
    outputs(868) <= not((layer0_outputs(2944)) xor (layer0_outputs(2196)));
    outputs(869) <= layer0_outputs(4526);
    outputs(870) <= layer0_outputs(1091);
    outputs(871) <= not(layer0_outputs(8716));
    outputs(872) <= not((layer0_outputs(11260)) xor (layer0_outputs(10047)));
    outputs(873) <= not(layer0_outputs(3108));
    outputs(874) <= (layer0_outputs(1630)) xor (layer0_outputs(4217));
    outputs(875) <= (layer0_outputs(6971)) or (layer0_outputs(4923));
    outputs(876) <= not(layer0_outputs(6214));
    outputs(877) <= layer0_outputs(7225);
    outputs(878) <= layer0_outputs(2847);
    outputs(879) <= (layer0_outputs(11125)) xor (layer0_outputs(11895));
    outputs(880) <= (layer0_outputs(10424)) xor (layer0_outputs(6089));
    outputs(881) <= layer0_outputs(12413);
    outputs(882) <= layer0_outputs(9060);
    outputs(883) <= not((layer0_outputs(12360)) and (layer0_outputs(12333)));
    outputs(884) <= layer0_outputs(4938);
    outputs(885) <= not((layer0_outputs(1983)) or (layer0_outputs(2238)));
    outputs(886) <= layer0_outputs(12497);
    outputs(887) <= (layer0_outputs(9254)) xor (layer0_outputs(10650));
    outputs(888) <= layer0_outputs(7580);
    outputs(889) <= not(layer0_outputs(3300));
    outputs(890) <= not((layer0_outputs(7462)) and (layer0_outputs(12627)));
    outputs(891) <= (layer0_outputs(5060)) or (layer0_outputs(9592));
    outputs(892) <= layer0_outputs(847);
    outputs(893) <= (layer0_outputs(3708)) xor (layer0_outputs(4908));
    outputs(894) <= (layer0_outputs(5465)) xor (layer0_outputs(4256));
    outputs(895) <= not(layer0_outputs(9822)) or (layer0_outputs(3415));
    outputs(896) <= (layer0_outputs(466)) and (layer0_outputs(12608));
    outputs(897) <= (layer0_outputs(4174)) and (layer0_outputs(9957));
    outputs(898) <= not(layer0_outputs(1869));
    outputs(899) <= layer0_outputs(11909);
    outputs(900) <= layer0_outputs(11554);
    outputs(901) <= not(layer0_outputs(10253));
    outputs(902) <= (layer0_outputs(6721)) or (layer0_outputs(2317));
    outputs(903) <= not(layer0_outputs(6205)) or (layer0_outputs(6922));
    outputs(904) <= layer0_outputs(402);
    outputs(905) <= layer0_outputs(8989);
    outputs(906) <= (layer0_outputs(1599)) or (layer0_outputs(3135));
    outputs(907) <= (layer0_outputs(8977)) and not (layer0_outputs(8615));
    outputs(908) <= not(layer0_outputs(6708));
    outputs(909) <= layer0_outputs(5871);
    outputs(910) <= not(layer0_outputs(10142)) or (layer0_outputs(10635));
    outputs(911) <= not((layer0_outputs(8300)) or (layer0_outputs(11929)));
    outputs(912) <= not((layer0_outputs(3138)) or (layer0_outputs(6369)));
    outputs(913) <= (layer0_outputs(7924)) and not (layer0_outputs(4285));
    outputs(914) <= (layer0_outputs(11793)) or (layer0_outputs(10289));
    outputs(915) <= not(layer0_outputs(8983));
    outputs(916) <= layer0_outputs(12099);
    outputs(917) <= not(layer0_outputs(2940));
    outputs(918) <= (layer0_outputs(8441)) and not (layer0_outputs(2791));
    outputs(919) <= (layer0_outputs(6671)) xor (layer0_outputs(8714));
    outputs(920) <= not(layer0_outputs(10903));
    outputs(921) <= not(layer0_outputs(9127));
    outputs(922) <= not(layer0_outputs(8205)) or (layer0_outputs(2739));
    outputs(923) <= not(layer0_outputs(3291));
    outputs(924) <= (layer0_outputs(9368)) and not (layer0_outputs(3537));
    outputs(925) <= (layer0_outputs(1488)) xor (layer0_outputs(10409));
    outputs(926) <= layer0_outputs(12583);
    outputs(927) <= not(layer0_outputs(8316));
    outputs(928) <= layer0_outputs(10336);
    outputs(929) <= '1';
    outputs(930) <= not(layer0_outputs(11492)) or (layer0_outputs(2559));
    outputs(931) <= not(layer0_outputs(8586));
    outputs(932) <= layer0_outputs(5561);
    outputs(933) <= (layer0_outputs(2752)) xor (layer0_outputs(1425));
    outputs(934) <= not(layer0_outputs(2695)) or (layer0_outputs(1782));
    outputs(935) <= not(layer0_outputs(10958)) or (layer0_outputs(10073));
    outputs(936) <= (layer0_outputs(6226)) or (layer0_outputs(4034));
    outputs(937) <= not((layer0_outputs(2248)) xor (layer0_outputs(6583)));
    outputs(938) <= not((layer0_outputs(6251)) xor (layer0_outputs(7882)));
    outputs(939) <= not(layer0_outputs(157));
    outputs(940) <= (layer0_outputs(5724)) or (layer0_outputs(9785));
    outputs(941) <= not(layer0_outputs(1077));
    outputs(942) <= not(layer0_outputs(768));
    outputs(943) <= not((layer0_outputs(1190)) and (layer0_outputs(4467)));
    outputs(944) <= not(layer0_outputs(7375));
    outputs(945) <= layer0_outputs(3794);
    outputs(946) <= not((layer0_outputs(12261)) or (layer0_outputs(7450)));
    outputs(947) <= layer0_outputs(3518);
    outputs(948) <= not((layer0_outputs(4509)) xor (layer0_outputs(7027)));
    outputs(949) <= not((layer0_outputs(8055)) xor (layer0_outputs(9496)));
    outputs(950) <= (layer0_outputs(2027)) or (layer0_outputs(732));
    outputs(951) <= (layer0_outputs(6360)) or (layer0_outputs(11755));
    outputs(952) <= (layer0_outputs(678)) and not (layer0_outputs(2793));
    outputs(953) <= not((layer0_outputs(6996)) xor (layer0_outputs(4715)));
    outputs(954) <= (layer0_outputs(11779)) and not (layer0_outputs(1843));
    outputs(955) <= not((layer0_outputs(1607)) xor (layer0_outputs(12211)));
    outputs(956) <= (layer0_outputs(1455)) xor (layer0_outputs(6583));
    outputs(957) <= not(layer0_outputs(6756)) or (layer0_outputs(7576));
    outputs(958) <= (layer0_outputs(6680)) xor (layer0_outputs(5259));
    outputs(959) <= not(layer0_outputs(6240));
    outputs(960) <= not(layer0_outputs(8412));
    outputs(961) <= layer0_outputs(4164);
    outputs(962) <= not(layer0_outputs(8635));
    outputs(963) <= not(layer0_outputs(5301));
    outputs(964) <= not((layer0_outputs(1797)) or (layer0_outputs(614)));
    outputs(965) <= layer0_outputs(5063);
    outputs(966) <= (layer0_outputs(6615)) or (layer0_outputs(10607));
    outputs(967) <= (layer0_outputs(8524)) or (layer0_outputs(5841));
    outputs(968) <= (layer0_outputs(12404)) and not (layer0_outputs(7687));
    outputs(969) <= (layer0_outputs(9151)) xor (layer0_outputs(12195));
    outputs(970) <= not(layer0_outputs(8348));
    outputs(971) <= layer0_outputs(9107);
    outputs(972) <= not((layer0_outputs(12463)) xor (layer0_outputs(3072)));
    outputs(973) <= layer0_outputs(10523);
    outputs(974) <= (layer0_outputs(11375)) and (layer0_outputs(9711));
    outputs(975) <= (layer0_outputs(3816)) and (layer0_outputs(8881));
    outputs(976) <= (layer0_outputs(499)) and not (layer0_outputs(946));
    outputs(977) <= layer0_outputs(7229);
    outputs(978) <= not((layer0_outputs(12115)) xor (layer0_outputs(5607)));
    outputs(979) <= (layer0_outputs(9597)) and not (layer0_outputs(2687));
    outputs(980) <= (layer0_outputs(612)) and (layer0_outputs(5870));
    outputs(981) <= (layer0_outputs(10996)) xor (layer0_outputs(8309));
    outputs(982) <= layer0_outputs(9528);
    outputs(983) <= (layer0_outputs(440)) xor (layer0_outputs(11838));
    outputs(984) <= layer0_outputs(8760);
    outputs(985) <= not(layer0_outputs(10448));
    outputs(986) <= (layer0_outputs(3997)) xor (layer0_outputs(6764));
    outputs(987) <= not((layer0_outputs(3499)) or (layer0_outputs(2359)));
    outputs(988) <= layer0_outputs(1550);
    outputs(989) <= not(layer0_outputs(12392));
    outputs(990) <= (layer0_outputs(7668)) and not (layer0_outputs(4449));
    outputs(991) <= '1';
    outputs(992) <= not(layer0_outputs(10557));
    outputs(993) <= not((layer0_outputs(7308)) xor (layer0_outputs(1974)));
    outputs(994) <= layer0_outputs(6700);
    outputs(995) <= not((layer0_outputs(3087)) and (layer0_outputs(7011)));
    outputs(996) <= not(layer0_outputs(12740));
    outputs(997) <= layer0_outputs(10565);
    outputs(998) <= not((layer0_outputs(9542)) xor (layer0_outputs(12625)));
    outputs(999) <= not((layer0_outputs(5710)) xor (layer0_outputs(11442)));
    outputs(1000) <= not(layer0_outputs(1259));
    outputs(1001) <= not((layer0_outputs(12422)) or (layer0_outputs(7612)));
    outputs(1002) <= (layer0_outputs(8905)) xor (layer0_outputs(1664));
    outputs(1003) <= not(layer0_outputs(4994));
    outputs(1004) <= not(layer0_outputs(3797));
    outputs(1005) <= (layer0_outputs(1310)) xor (layer0_outputs(1410));
    outputs(1006) <= layer0_outputs(10460);
    outputs(1007) <= not((layer0_outputs(1984)) and (layer0_outputs(4037)));
    outputs(1008) <= (layer0_outputs(10514)) xor (layer0_outputs(4086));
    outputs(1009) <= not(layer0_outputs(6277));
    outputs(1010) <= layer0_outputs(12517);
    outputs(1011) <= (layer0_outputs(731)) xor (layer0_outputs(2123));
    outputs(1012) <= not((layer0_outputs(347)) xor (layer0_outputs(7891)));
    outputs(1013) <= (layer0_outputs(9891)) xor (layer0_outputs(7829));
    outputs(1014) <= (layer0_outputs(218)) and not (layer0_outputs(4257));
    outputs(1015) <= layer0_outputs(2502);
    outputs(1016) <= (layer0_outputs(1719)) and (layer0_outputs(5355));
    outputs(1017) <= layer0_outputs(5626);
    outputs(1018) <= not((layer0_outputs(6475)) and (layer0_outputs(6466)));
    outputs(1019) <= (layer0_outputs(11205)) xor (layer0_outputs(9654));
    outputs(1020) <= (layer0_outputs(4129)) or (layer0_outputs(4982));
    outputs(1021) <= not(layer0_outputs(1346));
    outputs(1022) <= (layer0_outputs(12045)) and not (layer0_outputs(107));
    outputs(1023) <= not(layer0_outputs(9201));
    outputs(1024) <= (layer0_outputs(7827)) and not (layer0_outputs(6349));
    outputs(1025) <= not(layer0_outputs(3577));
    outputs(1026) <= layer0_outputs(5360);
    outputs(1027) <= not((layer0_outputs(10938)) xor (layer0_outputs(7323)));
    outputs(1028) <= not(layer0_outputs(4108));
    outputs(1029) <= not(layer0_outputs(10746));
    outputs(1030) <= layer0_outputs(5334);
    outputs(1031) <= not((layer0_outputs(6418)) xor (layer0_outputs(4167)));
    outputs(1032) <= layer0_outputs(4212);
    outputs(1033) <= layer0_outputs(8710);
    outputs(1034) <= layer0_outputs(6050);
    outputs(1035) <= not((layer0_outputs(4050)) or (layer0_outputs(2545)));
    outputs(1036) <= not(layer0_outputs(6354));
    outputs(1037) <= (layer0_outputs(3301)) and not (layer0_outputs(11226));
    outputs(1038) <= (layer0_outputs(10735)) xor (layer0_outputs(83));
    outputs(1039) <= not((layer0_outputs(6422)) xor (layer0_outputs(441)));
    outputs(1040) <= layer0_outputs(3449);
    outputs(1041) <= layer0_outputs(116);
    outputs(1042) <= not(layer0_outputs(3132)) or (layer0_outputs(2123));
    outputs(1043) <= not(layer0_outputs(4113));
    outputs(1044) <= (layer0_outputs(8195)) xor (layer0_outputs(11810));
    outputs(1045) <= not(layer0_outputs(6955));
    outputs(1046) <= layer0_outputs(4161);
    outputs(1047) <= layer0_outputs(1110);
    outputs(1048) <= (layer0_outputs(12155)) and not (layer0_outputs(2350));
    outputs(1049) <= not(layer0_outputs(10329));
    outputs(1050) <= not(layer0_outputs(9873));
    outputs(1051) <= layer0_outputs(989);
    outputs(1052) <= (layer0_outputs(8522)) xor (layer0_outputs(11007));
    outputs(1053) <= not(layer0_outputs(12016));
    outputs(1054) <= (layer0_outputs(4431)) and not (layer0_outputs(404));
    outputs(1055) <= not(layer0_outputs(2651)) or (layer0_outputs(6704));
    outputs(1056) <= (layer0_outputs(6056)) and (layer0_outputs(6054));
    outputs(1057) <= not(layer0_outputs(9243));
    outputs(1058) <= not(layer0_outputs(11998));
    outputs(1059) <= (layer0_outputs(4225)) xor (layer0_outputs(6122));
    outputs(1060) <= (layer0_outputs(6024)) xor (layer0_outputs(4437));
    outputs(1061) <= not((layer0_outputs(10956)) xor (layer0_outputs(9423)));
    outputs(1062) <= not(layer0_outputs(5718)) or (layer0_outputs(12219));
    outputs(1063) <= (layer0_outputs(4378)) and not (layer0_outputs(9211));
    outputs(1064) <= not(layer0_outputs(6140));
    outputs(1065) <= not((layer0_outputs(2573)) xor (layer0_outputs(5671)));
    outputs(1066) <= not((layer0_outputs(12266)) xor (layer0_outputs(1576)));
    outputs(1067) <= layer0_outputs(4716);
    outputs(1068) <= not(layer0_outputs(7604));
    outputs(1069) <= not(layer0_outputs(1850));
    outputs(1070) <= not(layer0_outputs(6622)) or (layer0_outputs(708));
    outputs(1071) <= layer0_outputs(5308);
    outputs(1072) <= not(layer0_outputs(1318));
    outputs(1073) <= not(layer0_outputs(3492));
    outputs(1074) <= (layer0_outputs(508)) xor (layer0_outputs(12549));
    outputs(1075) <= (layer0_outputs(6905)) or (layer0_outputs(11402));
    outputs(1076) <= not((layer0_outputs(9670)) xor (layer0_outputs(9327)));
    outputs(1077) <= (layer0_outputs(2181)) xor (layer0_outputs(2244));
    outputs(1078) <= not((layer0_outputs(11868)) xor (layer0_outputs(8502)));
    outputs(1079) <= (layer0_outputs(5697)) and (layer0_outputs(2896));
    outputs(1080) <= not(layer0_outputs(9629));
    outputs(1081) <= not((layer0_outputs(3238)) xor (layer0_outputs(1021)));
    outputs(1082) <= (layer0_outputs(3250)) xor (layer0_outputs(5931));
    outputs(1083) <= (layer0_outputs(10773)) xor (layer0_outputs(6797));
    outputs(1084) <= layer0_outputs(308);
    outputs(1085) <= (layer0_outputs(11057)) and (layer0_outputs(521));
    outputs(1086) <= (layer0_outputs(4952)) and (layer0_outputs(8263));
    outputs(1087) <= not(layer0_outputs(5231));
    outputs(1088) <= not((layer0_outputs(8075)) xor (layer0_outputs(10727)));
    outputs(1089) <= not(layer0_outputs(4442));
    outputs(1090) <= layer0_outputs(2617);
    outputs(1091) <= (layer0_outputs(1112)) xor (layer0_outputs(5688));
    outputs(1092) <= not(layer0_outputs(2543));
    outputs(1093) <= (layer0_outputs(8097)) and (layer0_outputs(12090));
    outputs(1094) <= layer0_outputs(10268);
    outputs(1095) <= not(layer0_outputs(9518)) or (layer0_outputs(1902));
    outputs(1096) <= not(layer0_outputs(8776));
    outputs(1097) <= (layer0_outputs(2155)) xor (layer0_outputs(4959));
    outputs(1098) <= not(layer0_outputs(2787)) or (layer0_outputs(12767));
    outputs(1099) <= not(layer0_outputs(6377));
    outputs(1100) <= layer0_outputs(3397);
    outputs(1101) <= (layer0_outputs(7609)) and (layer0_outputs(4140));
    outputs(1102) <= (layer0_outputs(9832)) and (layer0_outputs(9836));
    outputs(1103) <= not(layer0_outputs(945)) or (layer0_outputs(11772));
    outputs(1104) <= not(layer0_outputs(4730)) or (layer0_outputs(11984));
    outputs(1105) <= not(layer0_outputs(9972)) or (layer0_outputs(1221));
    outputs(1106) <= not(layer0_outputs(8768));
    outputs(1107) <= (layer0_outputs(11453)) xor (layer0_outputs(3692));
    outputs(1108) <= layer0_outputs(7634);
    outputs(1109) <= not((layer0_outputs(2351)) xor (layer0_outputs(9167)));
    outputs(1110) <= layer0_outputs(8483);
    outputs(1111) <= not(layer0_outputs(11477)) or (layer0_outputs(11640));
    outputs(1112) <= (layer0_outputs(2118)) xor (layer0_outputs(11219));
    outputs(1113) <= not(layer0_outputs(7533));
    outputs(1114) <= not((layer0_outputs(11129)) xor (layer0_outputs(11147)));
    outputs(1115) <= not((layer0_outputs(4401)) xor (layer0_outputs(12249)));
    outputs(1116) <= not(layer0_outputs(3582)) or (layer0_outputs(6669));
    outputs(1117) <= not(layer0_outputs(3491));
    outputs(1118) <= not(layer0_outputs(7091));
    outputs(1119) <= not((layer0_outputs(4176)) xor (layer0_outputs(10399)));
    outputs(1120) <= not(layer0_outputs(8489));
    outputs(1121) <= not((layer0_outputs(7521)) xor (layer0_outputs(5929)));
    outputs(1122) <= not((layer0_outputs(3168)) and (layer0_outputs(2937)));
    outputs(1123) <= (layer0_outputs(516)) and not (layer0_outputs(11400));
    outputs(1124) <= not(layer0_outputs(5472));
    outputs(1125) <= layer0_outputs(11352);
    outputs(1126) <= not((layer0_outputs(7295)) xor (layer0_outputs(11992)));
    outputs(1127) <= layer0_outputs(8468);
    outputs(1128) <= not((layer0_outputs(3817)) or (layer0_outputs(5735)));
    outputs(1129) <= not(layer0_outputs(8241)) or (layer0_outputs(8221));
    outputs(1130) <= not(layer0_outputs(4422));
    outputs(1131) <= (layer0_outputs(6477)) and not (layer0_outputs(1249));
    outputs(1132) <= (layer0_outputs(5116)) or (layer0_outputs(342));
    outputs(1133) <= not(layer0_outputs(10931));
    outputs(1134) <= (layer0_outputs(7236)) xor (layer0_outputs(8772));
    outputs(1135) <= layer0_outputs(154);
    outputs(1136) <= '1';
    outputs(1137) <= (layer0_outputs(2561)) and not (layer0_outputs(9750));
    outputs(1138) <= '1';
    outputs(1139) <= (layer0_outputs(9064)) and (layer0_outputs(2356));
    outputs(1140) <= layer0_outputs(1900);
    outputs(1141) <= (layer0_outputs(10320)) or (layer0_outputs(1133));
    outputs(1142) <= not((layer0_outputs(1105)) and (layer0_outputs(3338)));
    outputs(1143) <= (layer0_outputs(9582)) and not (layer0_outputs(12393));
    outputs(1144) <= (layer0_outputs(4271)) xor (layer0_outputs(8021));
    outputs(1145) <= not(layer0_outputs(5024));
    outputs(1146) <= layer0_outputs(8490);
    outputs(1147) <= not((layer0_outputs(2047)) xor (layer0_outputs(6567)));
    outputs(1148) <= layer0_outputs(6288);
    outputs(1149) <= not((layer0_outputs(2724)) or (layer0_outputs(7434)));
    outputs(1150) <= (layer0_outputs(6494)) xor (layer0_outputs(8568));
    outputs(1151) <= layer0_outputs(7645);
    outputs(1152) <= not(layer0_outputs(3843)) or (layer0_outputs(997));
    outputs(1153) <= not((layer0_outputs(3304)) xor (layer0_outputs(11436)));
    outputs(1154) <= not(layer0_outputs(5289));
    outputs(1155) <= not(layer0_outputs(8662)) or (layer0_outputs(1486));
    outputs(1156) <= not(layer0_outputs(3909));
    outputs(1157) <= not((layer0_outputs(5551)) xor (layer0_outputs(1916)));
    outputs(1158) <= not(layer0_outputs(6770));
    outputs(1159) <= not(layer0_outputs(4626));
    outputs(1160) <= not(layer0_outputs(4442));
    outputs(1161) <= not((layer0_outputs(3560)) or (layer0_outputs(6699)));
    outputs(1162) <= '1';
    outputs(1163) <= not((layer0_outputs(11430)) xor (layer0_outputs(7962)));
    outputs(1164) <= layer0_outputs(8762);
    outputs(1165) <= (layer0_outputs(5846)) xor (layer0_outputs(4980));
    outputs(1166) <= layer0_outputs(3225);
    outputs(1167) <= (layer0_outputs(6015)) and not (layer0_outputs(5776));
    outputs(1168) <= (layer0_outputs(5774)) xor (layer0_outputs(7698));
    outputs(1169) <= not((layer0_outputs(11265)) and (layer0_outputs(11617)));
    outputs(1170) <= (layer0_outputs(1894)) or (layer0_outputs(8037));
    outputs(1171) <= layer0_outputs(299);
    outputs(1172) <= not(layer0_outputs(32));
    outputs(1173) <= not(layer0_outputs(11249)) or (layer0_outputs(12759));
    outputs(1174) <= not((layer0_outputs(7725)) and (layer0_outputs(752)));
    outputs(1175) <= layer0_outputs(11392);
    outputs(1176) <= not(layer0_outputs(6605));
    outputs(1177) <= layer0_outputs(5066);
    outputs(1178) <= not(layer0_outputs(7388));
    outputs(1179) <= not(layer0_outputs(9330));
    outputs(1180) <= layer0_outputs(8173);
    outputs(1181) <= layer0_outputs(12319);
    outputs(1182) <= layer0_outputs(8623);
    outputs(1183) <= (layer0_outputs(3461)) and not (layer0_outputs(1888));
    outputs(1184) <= (layer0_outputs(289)) xor (layer0_outputs(5215));
    outputs(1185) <= (layer0_outputs(5189)) xor (layer0_outputs(12572));
    outputs(1186) <= not(layer0_outputs(123));
    outputs(1187) <= (layer0_outputs(6678)) and (layer0_outputs(3004));
    outputs(1188) <= not((layer0_outputs(10237)) or (layer0_outputs(8810)));
    outputs(1189) <= (layer0_outputs(8572)) xor (layer0_outputs(6273));
    outputs(1190) <= not(layer0_outputs(8877));
    outputs(1191) <= not((layer0_outputs(10574)) and (layer0_outputs(160)));
    outputs(1192) <= not(layer0_outputs(12480));
    outputs(1193) <= not((layer0_outputs(7778)) or (layer0_outputs(283)));
    outputs(1194) <= not(layer0_outputs(5643)) or (layer0_outputs(10153));
    outputs(1195) <= (layer0_outputs(11291)) and (layer0_outputs(4437));
    outputs(1196) <= not((layer0_outputs(3602)) xor (layer0_outputs(12496)));
    outputs(1197) <= not((layer0_outputs(7505)) xor (layer0_outputs(9207)));
    outputs(1198) <= layer0_outputs(8961);
    outputs(1199) <= layer0_outputs(7382);
    outputs(1200) <= layer0_outputs(3344);
    outputs(1201) <= not((layer0_outputs(7639)) xor (layer0_outputs(2321)));
    outputs(1202) <= (layer0_outputs(3737)) and (layer0_outputs(9398));
    outputs(1203) <= not(layer0_outputs(1330));
    outputs(1204) <= not(layer0_outputs(3887));
    outputs(1205) <= layer0_outputs(6242);
    outputs(1206) <= (layer0_outputs(8064)) or (layer0_outputs(2691));
    outputs(1207) <= not(layer0_outputs(960));
    outputs(1208) <= (layer0_outputs(8634)) xor (layer0_outputs(11693));
    outputs(1209) <= (layer0_outputs(2611)) and not (layer0_outputs(10687));
    outputs(1210) <= not(layer0_outputs(7974));
    outputs(1211) <= layer0_outputs(1448);
    outputs(1212) <= not((layer0_outputs(9986)) xor (layer0_outputs(5471)));
    outputs(1213) <= not((layer0_outputs(10783)) and (layer0_outputs(10123)));
    outputs(1214) <= layer0_outputs(11036);
    outputs(1215) <= not((layer0_outputs(7708)) xor (layer0_outputs(2994)));
    outputs(1216) <= not((layer0_outputs(5468)) xor (layer0_outputs(8600)));
    outputs(1217) <= not(layer0_outputs(4448));
    outputs(1218) <= not((layer0_outputs(5328)) xor (layer0_outputs(5412)));
    outputs(1219) <= (layer0_outputs(2418)) xor (layer0_outputs(4413));
    outputs(1220) <= not(layer0_outputs(11913));
    outputs(1221) <= not((layer0_outputs(3082)) and (layer0_outputs(6236)));
    outputs(1222) <= not((layer0_outputs(12742)) xor (layer0_outputs(10970)));
    outputs(1223) <= not((layer0_outputs(124)) or (layer0_outputs(4825)));
    outputs(1224) <= layer0_outputs(9951);
    outputs(1225) <= layer0_outputs(2727);
    outputs(1226) <= not((layer0_outputs(11450)) xor (layer0_outputs(9346)));
    outputs(1227) <= (layer0_outputs(6432)) and not (layer0_outputs(7379));
    outputs(1228) <= not(layer0_outputs(11122));
    outputs(1229) <= not(layer0_outputs(868));
    outputs(1230) <= not(layer0_outputs(2976));
    outputs(1231) <= (layer0_outputs(464)) or (layer0_outputs(5271));
    outputs(1232) <= (layer0_outputs(4586)) or (layer0_outputs(5241));
    outputs(1233) <= (layer0_outputs(3241)) xor (layer0_outputs(4659));
    outputs(1234) <= not((layer0_outputs(4230)) xor (layer0_outputs(12008)));
    outputs(1235) <= layer0_outputs(2334);
    outputs(1236) <= (layer0_outputs(11060)) or (layer0_outputs(1360));
    outputs(1237) <= layer0_outputs(6281);
    outputs(1238) <= not(layer0_outputs(12325));
    outputs(1239) <= layer0_outputs(7979);
    outputs(1240) <= not(layer0_outputs(3511));
    outputs(1241) <= (layer0_outputs(225)) and not (layer0_outputs(2159));
    outputs(1242) <= (layer0_outputs(4380)) and (layer0_outputs(11660));
    outputs(1243) <= (layer0_outputs(941)) xor (layer0_outputs(7958));
    outputs(1244) <= not(layer0_outputs(11625)) or (layer0_outputs(12391));
    outputs(1245) <= '1';
    outputs(1246) <= (layer0_outputs(3874)) and not (layer0_outputs(2886));
    outputs(1247) <= not(layer0_outputs(11055));
    outputs(1248) <= not(layer0_outputs(5273)) or (layer0_outputs(8259));
    outputs(1249) <= not(layer0_outputs(2251));
    outputs(1250) <= not((layer0_outputs(5269)) xor (layer0_outputs(9809)));
    outputs(1251) <= (layer0_outputs(78)) and (layer0_outputs(2564));
    outputs(1252) <= not((layer0_outputs(4626)) or (layer0_outputs(4849)));
    outputs(1253) <= layer0_outputs(683);
    outputs(1254) <= (layer0_outputs(7177)) or (layer0_outputs(4109));
    outputs(1255) <= layer0_outputs(5629);
    outputs(1256) <= (layer0_outputs(8173)) and not (layer0_outputs(9729));
    outputs(1257) <= layer0_outputs(2018);
    outputs(1258) <= not(layer0_outputs(11901)) or (layer0_outputs(7340));
    outputs(1259) <= (layer0_outputs(2248)) and (layer0_outputs(12157));
    outputs(1260) <= not(layer0_outputs(7385));
    outputs(1261) <= not((layer0_outputs(156)) xor (layer0_outputs(10686)));
    outputs(1262) <= (layer0_outputs(6350)) or (layer0_outputs(5099));
    outputs(1263) <= not(layer0_outputs(10081)) or (layer0_outputs(9721));
    outputs(1264) <= not(layer0_outputs(10375));
    outputs(1265) <= not((layer0_outputs(12148)) or (layer0_outputs(3648)));
    outputs(1266) <= (layer0_outputs(6607)) and not (layer0_outputs(4114));
    outputs(1267) <= not((layer0_outputs(1773)) xor (layer0_outputs(2461)));
    outputs(1268) <= (layer0_outputs(2152)) and (layer0_outputs(7130));
    outputs(1269) <= (layer0_outputs(10165)) and not (layer0_outputs(8891));
    outputs(1270) <= not((layer0_outputs(5457)) xor (layer0_outputs(5759)));
    outputs(1271) <= not((layer0_outputs(6944)) and (layer0_outputs(5343)));
    outputs(1272) <= not(layer0_outputs(7518));
    outputs(1273) <= (layer0_outputs(1066)) xor (layer0_outputs(11614));
    outputs(1274) <= not((layer0_outputs(11812)) and (layer0_outputs(6343)));
    outputs(1275) <= (layer0_outputs(7240)) xor (layer0_outputs(5632));
    outputs(1276) <= (layer0_outputs(7899)) xor (layer0_outputs(7730));
    outputs(1277) <= layer0_outputs(4130);
    outputs(1278) <= not(layer0_outputs(5173));
    outputs(1279) <= not(layer0_outputs(6896)) or (layer0_outputs(1411));
    outputs(1280) <= '0';
    outputs(1281) <= not((layer0_outputs(5540)) xor (layer0_outputs(5987)));
    outputs(1282) <= (layer0_outputs(6626)) and (layer0_outputs(10601));
    outputs(1283) <= layer0_outputs(1857);
    outputs(1284) <= (layer0_outputs(11149)) and not (layer0_outputs(4623));
    outputs(1285) <= layer0_outputs(5963);
    outputs(1286) <= (layer0_outputs(2942)) and not (layer0_outputs(6608));
    outputs(1287) <= not((layer0_outputs(6753)) or (layer0_outputs(4044)));
    outputs(1288) <= layer0_outputs(8463);
    outputs(1289) <= not(layer0_outputs(9556));
    outputs(1290) <= layer0_outputs(5925);
    outputs(1291) <= (layer0_outputs(10411)) xor (layer0_outputs(1354));
    outputs(1292) <= (layer0_outputs(10371)) and not (layer0_outputs(455));
    outputs(1293) <= not(layer0_outputs(998));
    outputs(1294) <= layer0_outputs(10144);
    outputs(1295) <= (layer0_outputs(957)) xor (layer0_outputs(3882));
    outputs(1296) <= layer0_outputs(12033);
    outputs(1297) <= layer0_outputs(6624);
    outputs(1298) <= not((layer0_outputs(2723)) xor (layer0_outputs(3777)));
    outputs(1299) <= not(layer0_outputs(9109));
    outputs(1300) <= '0';
    outputs(1301) <= not(layer0_outputs(2198));
    outputs(1302) <= not((layer0_outputs(7993)) xor (layer0_outputs(1279)));
    outputs(1303) <= '0';
    outputs(1304) <= (layer0_outputs(3108)) and not (layer0_outputs(6796));
    outputs(1305) <= (layer0_outputs(4975)) and (layer0_outputs(7787));
    outputs(1306) <= (layer0_outputs(8306)) xor (layer0_outputs(6452));
    outputs(1307) <= (layer0_outputs(2986)) and not (layer0_outputs(10355));
    outputs(1308) <= (layer0_outputs(12596)) and not (layer0_outputs(11601));
    outputs(1309) <= not((layer0_outputs(8727)) or (layer0_outputs(11316)));
    outputs(1310) <= (layer0_outputs(7339)) xor (layer0_outputs(3834));
    outputs(1311) <= layer0_outputs(4541);
    outputs(1312) <= layer0_outputs(9703);
    outputs(1313) <= not(layer0_outputs(7512));
    outputs(1314) <= (layer0_outputs(5866)) xor (layer0_outputs(465));
    outputs(1315) <= layer0_outputs(5412);
    outputs(1316) <= not(layer0_outputs(8324));
    outputs(1317) <= not((layer0_outputs(5390)) or (layer0_outputs(10099)));
    outputs(1318) <= (layer0_outputs(7283)) and not (layer0_outputs(12445));
    outputs(1319) <= not((layer0_outputs(740)) xor (layer0_outputs(632)));
    outputs(1320) <= layer0_outputs(5807);
    outputs(1321) <= not(layer0_outputs(6534));
    outputs(1322) <= not((layer0_outputs(7365)) xor (layer0_outputs(5995)));
    outputs(1323) <= not((layer0_outputs(12136)) xor (layer0_outputs(12790)));
    outputs(1324) <= not((layer0_outputs(10205)) xor (layer0_outputs(1025)));
    outputs(1325) <= not((layer0_outputs(3892)) xor (layer0_outputs(9810)));
    outputs(1326) <= not(layer0_outputs(3435));
    outputs(1327) <= not(layer0_outputs(7200)) or (layer0_outputs(1119));
    outputs(1328) <= (layer0_outputs(12082)) and not (layer0_outputs(6230));
    outputs(1329) <= layer0_outputs(12296);
    outputs(1330) <= layer0_outputs(5705);
    outputs(1331) <= layer0_outputs(1583);
    outputs(1332) <= layer0_outputs(5693);
    outputs(1333) <= not((layer0_outputs(8199)) xor (layer0_outputs(1658)));
    outputs(1334) <= (layer0_outputs(7635)) xor (layer0_outputs(1379));
    outputs(1335) <= not((layer0_outputs(3968)) xor (layer0_outputs(6744)));
    outputs(1336) <= (layer0_outputs(12024)) and not (layer0_outputs(5498));
    outputs(1337) <= not((layer0_outputs(602)) or (layer0_outputs(578)));
    outputs(1338) <= (layer0_outputs(6682)) or (layer0_outputs(11131));
    outputs(1339) <= (layer0_outputs(4198)) and not (layer0_outputs(8148));
    outputs(1340) <= not((layer0_outputs(1610)) xor (layer0_outputs(7520)));
    outputs(1341) <= (layer0_outputs(6069)) xor (layer0_outputs(1498));
    outputs(1342) <= (layer0_outputs(3008)) xor (layer0_outputs(4640));
    outputs(1343) <= (layer0_outputs(1090)) and not (layer0_outputs(10311));
    outputs(1344) <= '0';
    outputs(1345) <= (layer0_outputs(2551)) and not (layer0_outputs(1827));
    outputs(1346) <= (layer0_outputs(830)) and (layer0_outputs(2721));
    outputs(1347) <= not((layer0_outputs(5571)) xor (layer0_outputs(2429)));
    outputs(1348) <= not((layer0_outputs(7955)) xor (layer0_outputs(12467)));
    outputs(1349) <= (layer0_outputs(12255)) and not (layer0_outputs(2869));
    outputs(1350) <= '0';
    outputs(1351) <= (layer0_outputs(10523)) and not (layer0_outputs(1741));
    outputs(1352) <= (layer0_outputs(7414)) xor (layer0_outputs(3313));
    outputs(1353) <= not(layer0_outputs(11585));
    outputs(1354) <= not(layer0_outputs(2278));
    outputs(1355) <= '0';
    outputs(1356) <= not(layer0_outputs(6167));
    outputs(1357) <= not((layer0_outputs(4157)) or (layer0_outputs(1723)));
    outputs(1358) <= not((layer0_outputs(3542)) or (layer0_outputs(4708)));
    outputs(1359) <= layer0_outputs(3118);
    outputs(1360) <= layer0_outputs(5105);
    outputs(1361) <= (layer0_outputs(2671)) and not (layer0_outputs(3802));
    outputs(1362) <= not(layer0_outputs(2703));
    outputs(1363) <= not(layer0_outputs(9223));
    outputs(1364) <= (layer0_outputs(2604)) and not (layer0_outputs(12092));
    outputs(1365) <= (layer0_outputs(3504)) and not (layer0_outputs(5611));
    outputs(1366) <= (layer0_outputs(3761)) and not (layer0_outputs(6689));
    outputs(1367) <= not(layer0_outputs(6081));
    outputs(1368) <= (layer0_outputs(9220)) xor (layer0_outputs(3732));
    outputs(1369) <= (layer0_outputs(5345)) and (layer0_outputs(6984));
    outputs(1370) <= (layer0_outputs(4668)) xor (layer0_outputs(64));
    outputs(1371) <= layer0_outputs(8455);
    outputs(1372) <= layer0_outputs(3093);
    outputs(1373) <= layer0_outputs(6233);
    outputs(1374) <= not(layer0_outputs(5966));
    outputs(1375) <= layer0_outputs(8801);
    outputs(1376) <= (layer0_outputs(10966)) and (layer0_outputs(1489));
    outputs(1377) <= not(layer0_outputs(12));
    outputs(1378) <= (layer0_outputs(9171)) and (layer0_outputs(9808));
    outputs(1379) <= (layer0_outputs(4325)) and not (layer0_outputs(8366));
    outputs(1380) <= not((layer0_outputs(2641)) or (layer0_outputs(7148)));
    outputs(1381) <= not((layer0_outputs(7033)) or (layer0_outputs(1723)));
    outputs(1382) <= (layer0_outputs(11438)) and not (layer0_outputs(11535));
    outputs(1383) <= (layer0_outputs(9861)) and not (layer0_outputs(4208));
    outputs(1384) <= (layer0_outputs(10691)) and not (layer0_outputs(11120));
    outputs(1385) <= (layer0_outputs(2426)) xor (layer0_outputs(10185));
    outputs(1386) <= (layer0_outputs(6853)) and (layer0_outputs(5298));
    outputs(1387) <= (layer0_outputs(11520)) xor (layer0_outputs(8422));
    outputs(1388) <= (layer0_outputs(12462)) and not (layer0_outputs(6713));
    outputs(1389) <= layer0_outputs(10127);
    outputs(1390) <= not((layer0_outputs(10604)) or (layer0_outputs(11462)));
    outputs(1391) <= layer0_outputs(3469);
    outputs(1392) <= (layer0_outputs(4202)) xor (layer0_outputs(6536));
    outputs(1393) <= not(layer0_outputs(1559));
    outputs(1394) <= layer0_outputs(3007);
    outputs(1395) <= (layer0_outputs(9897)) and not (layer0_outputs(4973));
    outputs(1396) <= not(layer0_outputs(545));
    outputs(1397) <= (layer0_outputs(9883)) and not (layer0_outputs(3109));
    outputs(1398) <= not(layer0_outputs(3343));
    outputs(1399) <= '0';
    outputs(1400) <= not((layer0_outputs(5843)) or (layer0_outputs(11095)));
    outputs(1401) <= (layer0_outputs(12783)) and not (layer0_outputs(6385));
    outputs(1402) <= (layer0_outputs(2180)) xor (layer0_outputs(6744));
    outputs(1403) <= '0';
    outputs(1404) <= '0';
    outputs(1405) <= layer0_outputs(10481);
    outputs(1406) <= layer0_outputs(3073);
    outputs(1407) <= not(layer0_outputs(8373));
    outputs(1408) <= not((layer0_outputs(157)) xor (layer0_outputs(8491)));
    outputs(1409) <= layer0_outputs(6765);
    outputs(1410) <= not((layer0_outputs(10911)) or (layer0_outputs(778)));
    outputs(1411) <= (layer0_outputs(9257)) and (layer0_outputs(12379));
    outputs(1412) <= not(layer0_outputs(10575));
    outputs(1413) <= (layer0_outputs(870)) xor (layer0_outputs(3092));
    outputs(1414) <= '0';
    outputs(1415) <= (layer0_outputs(244)) and not (layer0_outputs(7648));
    outputs(1416) <= not(layer0_outputs(12541));
    outputs(1417) <= not((layer0_outputs(8985)) xor (layer0_outputs(7282)));
    outputs(1418) <= layer0_outputs(2774);
    outputs(1419) <= not((layer0_outputs(7628)) or (layer0_outputs(8147)));
    outputs(1420) <= (layer0_outputs(11597)) xor (layer0_outputs(12383));
    outputs(1421) <= (layer0_outputs(11564)) and not (layer0_outputs(9181));
    outputs(1422) <= (layer0_outputs(5297)) and (layer0_outputs(1146));
    outputs(1423) <= not(layer0_outputs(5183));
    outputs(1424) <= (layer0_outputs(12155)) and not (layer0_outputs(880));
    outputs(1425) <= not((layer0_outputs(11654)) or (layer0_outputs(12368)));
    outputs(1426) <= not(layer0_outputs(10885));
    outputs(1427) <= (layer0_outputs(2996)) and (layer0_outputs(8047));
    outputs(1428) <= layer0_outputs(5616);
    outputs(1429) <= not((layer0_outputs(2728)) and (layer0_outputs(8195)));
    outputs(1430) <= not(layer0_outputs(422));
    outputs(1431) <= (layer0_outputs(7341)) and not (layer0_outputs(859));
    outputs(1432) <= layer0_outputs(3101);
    outputs(1433) <= not((layer0_outputs(3652)) xor (layer0_outputs(6793)));
    outputs(1434) <= not((layer0_outputs(7038)) or (layer0_outputs(690)));
    outputs(1435) <= (layer0_outputs(4355)) xor (layer0_outputs(8149));
    outputs(1436) <= not((layer0_outputs(6863)) and (layer0_outputs(6259)));
    outputs(1437) <= layer0_outputs(2970);
    outputs(1438) <= (layer0_outputs(7948)) and (layer0_outputs(12775));
    outputs(1439) <= (layer0_outputs(10649)) and (layer0_outputs(12372));
    outputs(1440) <= (layer0_outputs(12598)) xor (layer0_outputs(1166));
    outputs(1441) <= (layer0_outputs(3607)) and (layer0_outputs(91));
    outputs(1442) <= layer0_outputs(8755);
    outputs(1443) <= (layer0_outputs(8654)) and (layer0_outputs(514));
    outputs(1444) <= layer0_outputs(6367);
    outputs(1445) <= (layer0_outputs(4911)) and not (layer0_outputs(242));
    outputs(1446) <= not(layer0_outputs(8325)) or (layer0_outputs(7769));
    outputs(1447) <= (layer0_outputs(7742)) and not (layer0_outputs(4041));
    outputs(1448) <= not((layer0_outputs(9537)) xor (layer0_outputs(1057)));
    outputs(1449) <= (layer0_outputs(11567)) or (layer0_outputs(11410));
    outputs(1450) <= (layer0_outputs(10263)) xor (layer0_outputs(3457));
    outputs(1451) <= layer0_outputs(5453);
    outputs(1452) <= (layer0_outputs(1920)) and (layer0_outputs(4724));
    outputs(1453) <= not((layer0_outputs(5006)) xor (layer0_outputs(6341)));
    outputs(1454) <= not((layer0_outputs(5330)) xor (layer0_outputs(308)));
    outputs(1455) <= layer0_outputs(11297);
    outputs(1456) <= not((layer0_outputs(6442)) or (layer0_outputs(4856)));
    outputs(1457) <= layer0_outputs(10640);
    outputs(1458) <= (layer0_outputs(1145)) xor (layer0_outputs(11562));
    outputs(1459) <= not((layer0_outputs(6884)) xor (layer0_outputs(4809)));
    outputs(1460) <= layer0_outputs(950);
    outputs(1461) <= (layer0_outputs(3369)) and (layer0_outputs(11592));
    outputs(1462) <= layer0_outputs(10894);
    outputs(1463) <= (layer0_outputs(5762)) and not (layer0_outputs(5235));
    outputs(1464) <= (layer0_outputs(11606)) and not (layer0_outputs(8070));
    outputs(1465) <= (layer0_outputs(6958)) and not (layer0_outputs(7895));
    outputs(1466) <= not((layer0_outputs(1760)) or (layer0_outputs(8031)));
    outputs(1467) <= (layer0_outputs(8105)) and not (layer0_outputs(4119));
    outputs(1468) <= (layer0_outputs(12094)) and not (layer0_outputs(1777));
    outputs(1469) <= (layer0_outputs(3195)) xor (layer0_outputs(12340));
    outputs(1470) <= not((layer0_outputs(2957)) or (layer0_outputs(5139)));
    outputs(1471) <= not((layer0_outputs(9748)) xor (layer0_outputs(12115)));
    outputs(1472) <= not((layer0_outputs(8347)) xor (layer0_outputs(9796)));
    outputs(1473) <= (layer0_outputs(10761)) and (layer0_outputs(1975));
    outputs(1474) <= (layer0_outputs(6295)) xor (layer0_outputs(3215));
    outputs(1475) <= layer0_outputs(9475);
    outputs(1476) <= (layer0_outputs(333)) xor (layer0_outputs(1716));
    outputs(1477) <= (layer0_outputs(6646)) xor (layer0_outputs(11041));
    outputs(1478) <= (layer0_outputs(9765)) and (layer0_outputs(7257));
    outputs(1479) <= (layer0_outputs(3119)) and (layer0_outputs(6644));
    outputs(1480) <= (layer0_outputs(4687)) and not (layer0_outputs(155));
    outputs(1481) <= not(layer0_outputs(4146)) or (layer0_outputs(10002));
    outputs(1482) <= not((layer0_outputs(2110)) or (layer0_outputs(7941)));
    outputs(1483) <= layer0_outputs(11340);
    outputs(1484) <= (layer0_outputs(9894)) and not (layer0_outputs(5108));
    outputs(1485) <= not((layer0_outputs(10053)) xor (layer0_outputs(2405)));
    outputs(1486) <= not(layer0_outputs(828));
    outputs(1487) <= not(layer0_outputs(5690));
    outputs(1488) <= (layer0_outputs(283)) and not (layer0_outputs(4358));
    outputs(1489) <= (layer0_outputs(7488)) xor (layer0_outputs(4689));
    outputs(1490) <= not(layer0_outputs(8284));
    outputs(1491) <= (layer0_outputs(7742)) and not (layer0_outputs(6338));
    outputs(1492) <= layer0_outputs(10374);
    outputs(1493) <= not(layer0_outputs(9934));
    outputs(1494) <= layer0_outputs(2432);
    outputs(1495) <= (layer0_outputs(7151)) and not (layer0_outputs(6215));
    outputs(1496) <= (layer0_outputs(973)) and (layer0_outputs(2505));
    outputs(1497) <= not((layer0_outputs(98)) or (layer0_outputs(3508)));
    outputs(1498) <= (layer0_outputs(2183)) and not (layer0_outputs(798));
    outputs(1499) <= layer0_outputs(2382);
    outputs(1500) <= (layer0_outputs(3271)) xor (layer0_outputs(7884));
    outputs(1501) <= (layer0_outputs(10262)) xor (layer0_outputs(10463));
    outputs(1502) <= (layer0_outputs(5306)) and (layer0_outputs(5995));
    outputs(1503) <= (layer0_outputs(7243)) xor (layer0_outputs(3584));
    outputs(1504) <= (layer0_outputs(1400)) xor (layer0_outputs(10798));
    outputs(1505) <= layer0_outputs(9016);
    outputs(1506) <= (layer0_outputs(7392)) and not (layer0_outputs(7056));
    outputs(1507) <= layer0_outputs(1394);
    outputs(1508) <= (layer0_outputs(10436)) and not (layer0_outputs(2245));
    outputs(1509) <= not((layer0_outputs(3937)) xor (layer0_outputs(7296)));
    outputs(1510) <= (layer0_outputs(8636)) and (layer0_outputs(1643));
    outputs(1511) <= not((layer0_outputs(12169)) xor (layer0_outputs(6629)));
    outputs(1512) <= '1';
    outputs(1513) <= not(layer0_outputs(7228));
    outputs(1514) <= '0';
    outputs(1515) <= (layer0_outputs(2253)) xor (layer0_outputs(5788));
    outputs(1516) <= not((layer0_outputs(3293)) or (layer0_outputs(8539)));
    outputs(1517) <= not((layer0_outputs(4105)) xor (layer0_outputs(2200)));
    outputs(1518) <= (layer0_outputs(11822)) xor (layer0_outputs(5178));
    outputs(1519) <= (layer0_outputs(5216)) and not (layer0_outputs(12129));
    outputs(1520) <= not(layer0_outputs(3040));
    outputs(1521) <= layer0_outputs(11782);
    outputs(1522) <= not(layer0_outputs(6337));
    outputs(1523) <= not(layer0_outputs(11614)) or (layer0_outputs(7791));
    outputs(1524) <= not((layer0_outputs(8812)) xor (layer0_outputs(1707)));
    outputs(1525) <= not(layer0_outputs(250));
    outputs(1526) <= not(layer0_outputs(7133));
    outputs(1527) <= not(layer0_outputs(729));
    outputs(1528) <= layer0_outputs(2534);
    outputs(1529) <= (layer0_outputs(9192)) and not (layer0_outputs(12610));
    outputs(1530) <= (layer0_outputs(10089)) and (layer0_outputs(4337));
    outputs(1531) <= (layer0_outputs(10000)) xor (layer0_outputs(10491));
    outputs(1532) <= '0';
    outputs(1533) <= not(layer0_outputs(6330));
    outputs(1534) <= not((layer0_outputs(7087)) xor (layer0_outputs(6933)));
    outputs(1535) <= layer0_outputs(7825);
    outputs(1536) <= not((layer0_outputs(8268)) xor (layer0_outputs(11321)));
    outputs(1537) <= not((layer0_outputs(12082)) xor (layer0_outputs(4266)));
    outputs(1538) <= not((layer0_outputs(6894)) xor (layer0_outputs(6992)));
    outputs(1539) <= not((layer0_outputs(894)) xor (layer0_outputs(7589)));
    outputs(1540) <= (layer0_outputs(12648)) and (layer0_outputs(1480));
    outputs(1541) <= layer0_outputs(850);
    outputs(1542) <= layer0_outputs(8103);
    outputs(1543) <= layer0_outputs(11479);
    outputs(1544) <= layer0_outputs(3740);
    outputs(1545) <= not((layer0_outputs(859)) or (layer0_outputs(11034)));
    outputs(1546) <= layer0_outputs(481);
    outputs(1547) <= not(layer0_outputs(2652));
    outputs(1548) <= (layer0_outputs(7506)) and not (layer0_outputs(7112));
    outputs(1549) <= layer0_outputs(559);
    outputs(1550) <= layer0_outputs(8413);
    outputs(1551) <= not((layer0_outputs(12596)) or (layer0_outputs(10219)));
    outputs(1552) <= not(layer0_outputs(2312));
    outputs(1553) <= not(layer0_outputs(5194));
    outputs(1554) <= (layer0_outputs(10102)) and (layer0_outputs(2290));
    outputs(1555) <= not((layer0_outputs(12216)) xor (layer0_outputs(6031)));
    outputs(1556) <= (layer0_outputs(5508)) and not (layer0_outputs(7348));
    outputs(1557) <= not((layer0_outputs(7507)) or (layer0_outputs(783)));
    outputs(1558) <= (layer0_outputs(745)) and not (layer0_outputs(12342));
    outputs(1559) <= not((layer0_outputs(630)) xor (layer0_outputs(6647)));
    outputs(1560) <= not((layer0_outputs(12352)) xor (layer0_outputs(6610)));
    outputs(1561) <= (layer0_outputs(12100)) and (layer0_outputs(11946));
    outputs(1562) <= (layer0_outputs(5474)) and (layer0_outputs(9391));
    outputs(1563) <= layer0_outputs(10330);
    outputs(1564) <= not((layer0_outputs(3494)) or (layer0_outputs(10597)));
    outputs(1565) <= not(layer0_outputs(214));
    outputs(1566) <= layer0_outputs(12326);
    outputs(1567) <= not((layer0_outputs(9930)) or (layer0_outputs(8031)));
    outputs(1568) <= not(layer0_outputs(8410));
    outputs(1569) <= not(layer0_outputs(3456));
    outputs(1570) <= (layer0_outputs(10747)) and not (layer0_outputs(9626));
    outputs(1571) <= not((layer0_outputs(4875)) xor (layer0_outputs(10526)));
    outputs(1572) <= not(layer0_outputs(1201));
    outputs(1573) <= (layer0_outputs(7043)) xor (layer0_outputs(6286));
    outputs(1574) <= not(layer0_outputs(6596));
    outputs(1575) <= (layer0_outputs(2966)) and not (layer0_outputs(4220));
    outputs(1576) <= (layer0_outputs(12710)) xor (layer0_outputs(407));
    outputs(1577) <= not(layer0_outputs(6996));
    outputs(1578) <= (layer0_outputs(10489)) and not (layer0_outputs(9694));
    outputs(1579) <= (layer0_outputs(12663)) xor (layer0_outputs(11254));
    outputs(1580) <= (layer0_outputs(7650)) and (layer0_outputs(9178));
    outputs(1581) <= (layer0_outputs(2500)) and (layer0_outputs(12427));
    outputs(1582) <= not((layer0_outputs(3060)) xor (layer0_outputs(3392)));
    outputs(1583) <= not((layer0_outputs(8025)) or (layer0_outputs(6837)));
    outputs(1584) <= layer0_outputs(9626);
    outputs(1585) <= not((layer0_outputs(7428)) or (layer0_outputs(7458)));
    outputs(1586) <= (layer0_outputs(10357)) xor (layer0_outputs(3244));
    outputs(1587) <= (layer0_outputs(9495)) and not (layer0_outputs(6312));
    outputs(1588) <= not(layer0_outputs(6961));
    outputs(1589) <= (layer0_outputs(8554)) xor (layer0_outputs(11004));
    outputs(1590) <= not((layer0_outputs(7912)) or (layer0_outputs(7726)));
    outputs(1591) <= not((layer0_outputs(185)) xor (layer0_outputs(4855)));
    outputs(1592) <= not((layer0_outputs(9021)) or (layer0_outputs(672)));
    outputs(1593) <= not(layer0_outputs(1365));
    outputs(1594) <= '0';
    outputs(1595) <= not(layer0_outputs(4821));
    outputs(1596) <= (layer0_outputs(1285)) and not (layer0_outputs(12619));
    outputs(1597) <= not(layer0_outputs(9501));
    outputs(1598) <= (layer0_outputs(2163)) xor (layer0_outputs(795));
    outputs(1599) <= not((layer0_outputs(1865)) or (layer0_outputs(0)));
    outputs(1600) <= not(layer0_outputs(12003));
    outputs(1601) <= (layer0_outputs(2788)) xor (layer0_outputs(356));
    outputs(1602) <= not((layer0_outputs(6781)) xor (layer0_outputs(1651)));
    outputs(1603) <= not((layer0_outputs(6511)) xor (layer0_outputs(4251)));
    outputs(1604) <= not(layer0_outputs(5653));
    outputs(1605) <= not((layer0_outputs(12594)) xor (layer0_outputs(51)));
    outputs(1606) <= (layer0_outputs(5809)) and not (layer0_outputs(11998));
    outputs(1607) <= not((layer0_outputs(5596)) or (layer0_outputs(11326)));
    outputs(1608) <= (layer0_outputs(8933)) and not (layer0_outputs(434));
    outputs(1609) <= not(layer0_outputs(7484));
    outputs(1610) <= not((layer0_outputs(7935)) or (layer0_outputs(2675)));
    outputs(1611) <= not(layer0_outputs(9476));
    outputs(1612) <= (layer0_outputs(7152)) xor (layer0_outputs(2397));
    outputs(1613) <= not(layer0_outputs(12165));
    outputs(1614) <= not((layer0_outputs(12411)) xor (layer0_outputs(4710)));
    outputs(1615) <= (layer0_outputs(12107)) and not (layer0_outputs(1300));
    outputs(1616) <= not((layer0_outputs(9540)) or (layer0_outputs(5825)));
    outputs(1617) <= layer0_outputs(10254);
    outputs(1618) <= (layer0_outputs(4896)) or (layer0_outputs(3683));
    outputs(1619) <= (layer0_outputs(6783)) xor (layer0_outputs(8429));
    outputs(1620) <= (layer0_outputs(10013)) and (layer0_outputs(1932));
    outputs(1621) <= layer0_outputs(9320);
    outputs(1622) <= (layer0_outputs(1987)) xor (layer0_outputs(9592));
    outputs(1623) <= not((layer0_outputs(1089)) xor (layer0_outputs(10058)));
    outputs(1624) <= '0';
    outputs(1625) <= layer0_outputs(4991);
    outputs(1626) <= not(layer0_outputs(11594));
    outputs(1627) <= not(layer0_outputs(3006));
    outputs(1628) <= not(layer0_outputs(5566));
    outputs(1629) <= (layer0_outputs(1241)) and not (layer0_outputs(9094));
    outputs(1630) <= '0';
    outputs(1631) <= layer0_outputs(8016);
    outputs(1632) <= (layer0_outputs(8289)) and (layer0_outputs(9863));
    outputs(1633) <= layer0_outputs(4937);
    outputs(1634) <= (layer0_outputs(9079)) and (layer0_outputs(7922));
    outputs(1635) <= (layer0_outputs(3164)) and not (layer0_outputs(12210));
    outputs(1636) <= (layer0_outputs(11151)) and (layer0_outputs(7996));
    outputs(1637) <= (layer0_outputs(4954)) and not (layer0_outputs(8781));
    outputs(1638) <= (layer0_outputs(598)) and not (layer0_outputs(3999));
    outputs(1639) <= layer0_outputs(10014);
    outputs(1640) <= not((layer0_outputs(9296)) and (layer0_outputs(748)));
    outputs(1641) <= layer0_outputs(10643);
    outputs(1642) <= (layer0_outputs(139)) xor (layer0_outputs(5252));
    outputs(1643) <= not(layer0_outputs(1163));
    outputs(1644) <= not(layer0_outputs(10582)) or (layer0_outputs(3098));
    outputs(1645) <= not(layer0_outputs(9622));
    outputs(1646) <= (layer0_outputs(4690)) and not (layer0_outputs(1122));
    outputs(1647) <= (layer0_outputs(5761)) and not (layer0_outputs(2982));
    outputs(1648) <= (layer0_outputs(220)) and not (layer0_outputs(10572));
    outputs(1649) <= not(layer0_outputs(5904));
    outputs(1650) <= (layer0_outputs(10499)) and not (layer0_outputs(4645));
    outputs(1651) <= not(layer0_outputs(8849));
    outputs(1652) <= not(layer0_outputs(8349));
    outputs(1653) <= (layer0_outputs(1936)) and not (layer0_outputs(4972));
    outputs(1654) <= (layer0_outputs(8444)) and not (layer0_outputs(11815));
    outputs(1655) <= not((layer0_outputs(8023)) and (layer0_outputs(9561)));
    outputs(1656) <= (layer0_outputs(1512)) or (layer0_outputs(10675));
    outputs(1657) <= not(layer0_outputs(1232));
    outputs(1658) <= not(layer0_outputs(5840));
    outputs(1659) <= (layer0_outputs(10642)) and not (layer0_outputs(11278));
    outputs(1660) <= layer0_outputs(8087);
    outputs(1661) <= (layer0_outputs(3359)) and (layer0_outputs(2904));
    outputs(1662) <= '0';
    outputs(1663) <= (layer0_outputs(888)) and not (layer0_outputs(4854));
    outputs(1664) <= not(layer0_outputs(1472));
    outputs(1665) <= not((layer0_outputs(3134)) or (layer0_outputs(11968)));
    outputs(1666) <= not((layer0_outputs(2135)) or (layer0_outputs(557)));
    outputs(1667) <= '0';
    outputs(1668) <= (layer0_outputs(3415)) and not (layer0_outputs(8456));
    outputs(1669) <= not((layer0_outputs(1559)) or (layer0_outputs(826)));
    outputs(1670) <= '0';
    outputs(1671) <= (layer0_outputs(3148)) xor (layer0_outputs(2289));
    outputs(1672) <= (layer0_outputs(9123)) and not (layer0_outputs(1772));
    outputs(1673) <= not(layer0_outputs(6161));
    outputs(1674) <= not((layer0_outputs(4152)) xor (layer0_outputs(4387)));
    outputs(1675) <= (layer0_outputs(11256)) and not (layer0_outputs(7441));
    outputs(1676) <= layer0_outputs(6438);
    outputs(1677) <= not((layer0_outputs(544)) xor (layer0_outputs(1802)));
    outputs(1678) <= (layer0_outputs(2916)) and (layer0_outputs(10221));
    outputs(1679) <= not(layer0_outputs(2362));
    outputs(1680) <= not(layer0_outputs(6950)) or (layer0_outputs(10334));
    outputs(1681) <= layer0_outputs(1990);
    outputs(1682) <= not(layer0_outputs(12388));
    outputs(1683) <= layer0_outputs(12739);
    outputs(1684) <= (layer0_outputs(1712)) and not (layer0_outputs(7928));
    outputs(1685) <= (layer0_outputs(4456)) and not (layer0_outputs(12315));
    outputs(1686) <= not((layer0_outputs(1698)) xor (layer0_outputs(5053)));
    outputs(1687) <= (layer0_outputs(7416)) and not (layer0_outputs(10822));
    outputs(1688) <= not((layer0_outputs(717)) xor (layer0_outputs(1792)));
    outputs(1689) <= layer0_outputs(12169);
    outputs(1690) <= layer0_outputs(11106);
    outputs(1691) <= (layer0_outputs(6947)) xor (layer0_outputs(11641));
    outputs(1692) <= layer0_outputs(7994);
    outputs(1693) <= layer0_outputs(10578);
    outputs(1694) <= layer0_outputs(6945);
    outputs(1695) <= (layer0_outputs(9643)) and not (layer0_outputs(2239));
    outputs(1696) <= (layer0_outputs(7324)) and not (layer0_outputs(8735));
    outputs(1697) <= layer0_outputs(2146);
    outputs(1698) <= (layer0_outputs(3184)) and (layer0_outputs(10558));
    outputs(1699) <= layer0_outputs(10752);
    outputs(1700) <= layer0_outputs(7039);
    outputs(1701) <= not((layer0_outputs(7873)) xor (layer0_outputs(2446)));
    outputs(1702) <= not((layer0_outputs(12066)) or (layer0_outputs(5335)));
    outputs(1703) <= not((layer0_outputs(67)) xor (layer0_outputs(6314)));
    outputs(1704) <= (layer0_outputs(7961)) or (layer0_outputs(8257));
    outputs(1705) <= (layer0_outputs(113)) and (layer0_outputs(2698));
    outputs(1706) <= (layer0_outputs(905)) and not (layer0_outputs(7889));
    outputs(1707) <= (layer0_outputs(1221)) and not (layer0_outputs(10620));
    outputs(1708) <= not(layer0_outputs(466));
    outputs(1709) <= (layer0_outputs(11532)) and not (layer0_outputs(7806));
    outputs(1710) <= (layer0_outputs(1416)) and not (layer0_outputs(5743));
    outputs(1711) <= not((layer0_outputs(10428)) or (layer0_outputs(12134)));
    outputs(1712) <= layer0_outputs(12245);
    outputs(1713) <= (layer0_outputs(11428)) and not (layer0_outputs(1252));
    outputs(1714) <= (layer0_outputs(896)) and not (layer0_outputs(4927));
    outputs(1715) <= (layer0_outputs(7340)) and (layer0_outputs(3618));
    outputs(1716) <= (layer0_outputs(1134)) and not (layer0_outputs(3240));
    outputs(1717) <= not(layer0_outputs(7437));
    outputs(1718) <= '0';
    outputs(1719) <= not(layer0_outputs(9969));
    outputs(1720) <= not(layer0_outputs(11395));
    outputs(1721) <= (layer0_outputs(8787)) and not (layer0_outputs(5930));
    outputs(1722) <= (layer0_outputs(12176)) and not (layer0_outputs(4857));
    outputs(1723) <= (layer0_outputs(5756)) and not (layer0_outputs(1622));
    outputs(1724) <= '1';
    outputs(1725) <= (layer0_outputs(6566)) xor (layer0_outputs(4499));
    outputs(1726) <= '0';
    outputs(1727) <= (layer0_outputs(1958)) and not (layer0_outputs(10330));
    outputs(1728) <= layer0_outputs(7943);
    outputs(1729) <= not((layer0_outputs(8250)) xor (layer0_outputs(2699)));
    outputs(1730) <= (layer0_outputs(3081)) and (layer0_outputs(3811));
    outputs(1731) <= (layer0_outputs(1081)) xor (layer0_outputs(3061));
    outputs(1732) <= (layer0_outputs(1690)) and not (layer0_outputs(1829));
    outputs(1733) <= (layer0_outputs(11688)) and not (layer0_outputs(4768));
    outputs(1734) <= not((layer0_outputs(6657)) xor (layer0_outputs(770)));
    outputs(1735) <= (layer0_outputs(2674)) xor (layer0_outputs(12531));
    outputs(1736) <= not(layer0_outputs(1149));
    outputs(1737) <= (layer0_outputs(11969)) and not (layer0_outputs(9781));
    outputs(1738) <= not(layer0_outputs(1158));
    outputs(1739) <= not(layer0_outputs(7534));
    outputs(1740) <= not((layer0_outputs(392)) xor (layer0_outputs(8863)));
    outputs(1741) <= not(layer0_outputs(2876));
    outputs(1742) <= not(layer0_outputs(3518));
    outputs(1743) <= (layer0_outputs(8390)) and (layer0_outputs(383));
    outputs(1744) <= not((layer0_outputs(11173)) or (layer0_outputs(8007)));
    outputs(1745) <= layer0_outputs(11418);
    outputs(1746) <= not((layer0_outputs(3418)) or (layer0_outputs(3192)));
    outputs(1747) <= not((layer0_outputs(8304)) or (layer0_outputs(6462)));
    outputs(1748) <= not((layer0_outputs(2613)) xor (layer0_outputs(5632)));
    outputs(1749) <= (layer0_outputs(12357)) xor (layer0_outputs(6808));
    outputs(1750) <= layer0_outputs(430);
    outputs(1751) <= (layer0_outputs(3307)) and not (layer0_outputs(10090));
    outputs(1752) <= layer0_outputs(8763);
    outputs(1753) <= not(layer0_outputs(9461)) or (layer0_outputs(9967));
    outputs(1754) <= not((layer0_outputs(12769)) or (layer0_outputs(11860)));
    outputs(1755) <= layer0_outputs(7132);
    outputs(1756) <= not((layer0_outputs(10076)) or (layer0_outputs(12459)));
    outputs(1757) <= not((layer0_outputs(6552)) and (layer0_outputs(5969)));
    outputs(1758) <= (layer0_outputs(8921)) xor (layer0_outputs(8875));
    outputs(1759) <= not(layer0_outputs(425));
    outputs(1760) <= not(layer0_outputs(10042));
    outputs(1761) <= (layer0_outputs(2891)) and (layer0_outputs(7078));
    outputs(1762) <= (layer0_outputs(3622)) xor (layer0_outputs(10777));
    outputs(1763) <= layer0_outputs(1769);
    outputs(1764) <= not((layer0_outputs(12053)) or (layer0_outputs(5654)));
    outputs(1765) <= (layer0_outputs(3318)) xor (layer0_outputs(8211));
    outputs(1766) <= layer0_outputs(5148);
    outputs(1767) <= not(layer0_outputs(9094));
    outputs(1768) <= (layer0_outputs(24)) and not (layer0_outputs(3506));
    outputs(1769) <= not(layer0_outputs(8811));
    outputs(1770) <= not((layer0_outputs(232)) and (layer0_outputs(10530)));
    outputs(1771) <= not((layer0_outputs(963)) or (layer0_outputs(12550)));
    outputs(1772) <= (layer0_outputs(8514)) xor (layer0_outputs(17));
    outputs(1773) <= not(layer0_outputs(5589));
    outputs(1774) <= (layer0_outputs(12291)) and not (layer0_outputs(8182));
    outputs(1775) <= (layer0_outputs(8345)) and not (layer0_outputs(10965));
    outputs(1776) <= not(layer0_outputs(4155));
    outputs(1777) <= (layer0_outputs(5725)) and not (layer0_outputs(11536));
    outputs(1778) <= not(layer0_outputs(5896)) or (layer0_outputs(374));
    outputs(1779) <= (layer0_outputs(3061)) xor (layer0_outputs(5766));
    outputs(1780) <= not((layer0_outputs(8632)) or (layer0_outputs(2569)));
    outputs(1781) <= layer0_outputs(12224);
    outputs(1782) <= not((layer0_outputs(7401)) and (layer0_outputs(10637)));
    outputs(1783) <= not((layer0_outputs(1291)) and (layer0_outputs(6188)));
    outputs(1784) <= (layer0_outputs(134)) and not (layer0_outputs(5268));
    outputs(1785) <= (layer0_outputs(10022)) and not (layer0_outputs(3790));
    outputs(1786) <= not(layer0_outputs(7781));
    outputs(1787) <= not((layer0_outputs(11701)) xor (layer0_outputs(11797)));
    outputs(1788) <= (layer0_outputs(3612)) xor (layer0_outputs(11579));
    outputs(1789) <= '0';
    outputs(1790) <= layer0_outputs(11995);
    outputs(1791) <= (layer0_outputs(1027)) xor (layer0_outputs(4928));
    outputs(1792) <= not(layer0_outputs(5922)) or (layer0_outputs(8744));
    outputs(1793) <= layer0_outputs(8119);
    outputs(1794) <= (layer0_outputs(8687)) xor (layer0_outputs(11896));
    outputs(1795) <= layer0_outputs(8119);
    outputs(1796) <= not((layer0_outputs(3172)) or (layer0_outputs(2215)));
    outputs(1797) <= layer0_outputs(10589);
    outputs(1798) <= (layer0_outputs(11418)) xor (layer0_outputs(10054));
    outputs(1799) <= (layer0_outputs(12184)) and not (layer0_outputs(46));
    outputs(1800) <= layer0_outputs(6519);
    outputs(1801) <= layer0_outputs(3642);
    outputs(1802) <= (layer0_outputs(10862)) xor (layer0_outputs(9057));
    outputs(1803) <= not((layer0_outputs(9762)) or (layer0_outputs(12387)));
    outputs(1804) <= (layer0_outputs(5774)) and not (layer0_outputs(358));
    outputs(1805) <= layer0_outputs(9445);
    outputs(1806) <= layer0_outputs(7564);
    outputs(1807) <= not((layer0_outputs(3696)) and (layer0_outputs(4377)));
    outputs(1808) <= not((layer0_outputs(2586)) xor (layer0_outputs(12149)));
    outputs(1809) <= (layer0_outputs(12049)) and not (layer0_outputs(5390));
    outputs(1810) <= (layer0_outputs(6549)) and not (layer0_outputs(3628));
    outputs(1811) <= (layer0_outputs(12080)) and not (layer0_outputs(6072));
    outputs(1812) <= not((layer0_outputs(3381)) or (layer0_outputs(11471)));
    outputs(1813) <= layer0_outputs(4370);
    outputs(1814) <= layer0_outputs(9933);
    outputs(1815) <= not((layer0_outputs(12001)) or (layer0_outputs(1207)));
    outputs(1816) <= '0';
    outputs(1817) <= not((layer0_outputs(2969)) xor (layer0_outputs(2595)));
    outputs(1818) <= not((layer0_outputs(11786)) or (layer0_outputs(2131)));
    outputs(1819) <= not((layer0_outputs(1316)) or (layer0_outputs(2190)));
    outputs(1820) <= not((layer0_outputs(2675)) xor (layer0_outputs(2472)));
    outputs(1821) <= not(layer0_outputs(6177));
    outputs(1822) <= not((layer0_outputs(8971)) xor (layer0_outputs(1730)));
    outputs(1823) <= (layer0_outputs(4466)) and not (layer0_outputs(10780));
    outputs(1824) <= (layer0_outputs(1069)) xor (layer0_outputs(679));
    outputs(1825) <= not(layer0_outputs(4647));
    outputs(1826) <= layer0_outputs(6130);
    outputs(1827) <= not((layer0_outputs(953)) or (layer0_outputs(7391)));
    outputs(1828) <= layer0_outputs(5897);
    outputs(1829) <= not((layer0_outputs(1656)) xor (layer0_outputs(11556)));
    outputs(1830) <= (layer0_outputs(3533)) and (layer0_outputs(11293));
    outputs(1831) <= (layer0_outputs(3179)) xor (layer0_outputs(1349));
    outputs(1832) <= '0';
    outputs(1833) <= (layer0_outputs(828)) xor (layer0_outputs(1339));
    outputs(1834) <= not(layer0_outputs(6972));
    outputs(1835) <= not(layer0_outputs(8338));
    outputs(1836) <= '0';
    outputs(1837) <= (layer0_outputs(11043)) and (layer0_outputs(1943));
    outputs(1838) <= not((layer0_outputs(2039)) or (layer0_outputs(7925)));
    outputs(1839) <= (layer0_outputs(3325)) and not (layer0_outputs(8652));
    outputs(1840) <= (layer0_outputs(9453)) and not (layer0_outputs(7195));
    outputs(1841) <= layer0_outputs(2817);
    outputs(1842) <= (layer0_outputs(7052)) xor (layer0_outputs(8829));
    outputs(1843) <= layer0_outputs(8929);
    outputs(1844) <= (layer0_outputs(8294)) and not (layer0_outputs(6036));
    outputs(1845) <= layer0_outputs(2875);
    outputs(1846) <= layer0_outputs(7080);
    outputs(1847) <= not(layer0_outputs(6394));
    outputs(1848) <= (layer0_outputs(5956)) and (layer0_outputs(6853));
    outputs(1849) <= not(layer0_outputs(12237));
    outputs(1850) <= not(layer0_outputs(2388));
    outputs(1851) <= layer0_outputs(11502);
    outputs(1852) <= (layer0_outputs(5725)) and not (layer0_outputs(2898));
    outputs(1853) <= not(layer0_outputs(7354));
    outputs(1854) <= (layer0_outputs(8978)) and (layer0_outputs(2295));
    outputs(1855) <= layer0_outputs(5225);
    outputs(1856) <= (layer0_outputs(11624)) and (layer0_outputs(11196));
    outputs(1857) <= (layer0_outputs(4295)) xor (layer0_outputs(524));
    outputs(1858) <= (layer0_outputs(6010)) and not (layer0_outputs(5636));
    outputs(1859) <= layer0_outputs(4248);
    outputs(1860) <= (layer0_outputs(7478)) and not (layer0_outputs(10129));
    outputs(1861) <= (layer0_outputs(12286)) and (layer0_outputs(1547));
    outputs(1862) <= layer0_outputs(305);
    outputs(1863) <= not((layer0_outputs(8820)) and (layer0_outputs(10827)));
    outputs(1864) <= not((layer0_outputs(280)) xor (layer0_outputs(8785)));
    outputs(1865) <= (layer0_outputs(11456)) and not (layer0_outputs(2540));
    outputs(1866) <= not(layer0_outputs(6499)) or (layer0_outputs(5384));
    outputs(1867) <= (layer0_outputs(8590)) xor (layer0_outputs(7862));
    outputs(1868) <= not((layer0_outputs(5715)) xor (layer0_outputs(9723)));
    outputs(1869) <= not(layer0_outputs(12168));
    outputs(1870) <= not((layer0_outputs(1159)) or (layer0_outputs(12343)));
    outputs(1871) <= (layer0_outputs(5213)) and (layer0_outputs(3534));
    outputs(1872) <= (layer0_outputs(8288)) and not (layer0_outputs(7701));
    outputs(1873) <= not((layer0_outputs(11039)) xor (layer0_outputs(405)));
    outputs(1874) <= not((layer0_outputs(7877)) xor (layer0_outputs(10110)));
    outputs(1875) <= (layer0_outputs(12183)) xor (layer0_outputs(3144));
    outputs(1876) <= not((layer0_outputs(567)) xor (layer0_outputs(10949)));
    outputs(1877) <= (layer0_outputs(1874)) and not (layer0_outputs(3187));
    outputs(1878) <= not((layer0_outputs(6693)) xor (layer0_outputs(7764)));
    outputs(1879) <= (layer0_outputs(10177)) xor (layer0_outputs(10821));
    outputs(1880) <= not((layer0_outputs(2046)) xor (layer0_outputs(2706)));
    outputs(1881) <= (layer0_outputs(4113)) and not (layer0_outputs(11659));
    outputs(1882) <= (layer0_outputs(8085)) and not (layer0_outputs(5793));
    outputs(1883) <= layer0_outputs(5374);
    outputs(1884) <= (layer0_outputs(10154)) and (layer0_outputs(11700));
    outputs(1885) <= not(layer0_outputs(2889));
    outputs(1886) <= layer0_outputs(1335);
    outputs(1887) <= not((layer0_outputs(354)) or (layer0_outputs(12646)));
    outputs(1888) <= '0';
    outputs(1889) <= layer0_outputs(2275);
    outputs(1890) <= not(layer0_outputs(3259));
    outputs(1891) <= (layer0_outputs(1905)) and (layer0_outputs(10325));
    outputs(1892) <= layer0_outputs(11139);
    outputs(1893) <= not(layer0_outputs(9808)) or (layer0_outputs(2112));
    outputs(1894) <= (layer0_outputs(1064)) xor (layer0_outputs(1705));
    outputs(1895) <= not(layer0_outputs(8886));
    outputs(1896) <= (layer0_outputs(5929)) or (layer0_outputs(2841));
    outputs(1897) <= layer0_outputs(4234);
    outputs(1898) <= not(layer0_outputs(3094));
    outputs(1899) <= '0';
    outputs(1900) <= layer0_outputs(6016);
    outputs(1901) <= not(layer0_outputs(10614));
    outputs(1902) <= (layer0_outputs(11763)) and not (layer0_outputs(10306));
    outputs(1903) <= layer0_outputs(10980);
    outputs(1904) <= (layer0_outputs(12038)) xor (layer0_outputs(7100));
    outputs(1905) <= not(layer0_outputs(10625));
    outputs(1906) <= not((layer0_outputs(11767)) xor (layer0_outputs(6426)));
    outputs(1907) <= layer0_outputs(10737);
    outputs(1908) <= (layer0_outputs(2972)) and not (layer0_outputs(11252));
    outputs(1909) <= layer0_outputs(3610);
    outputs(1910) <= (layer0_outputs(6016)) and not (layer0_outputs(7574));
    outputs(1911) <= not((layer0_outputs(4871)) xor (layer0_outputs(1337)));
    outputs(1912) <= (layer0_outputs(3139)) and (layer0_outputs(7137));
    outputs(1913) <= layer0_outputs(7070);
    outputs(1914) <= layer0_outputs(460);
    outputs(1915) <= (layer0_outputs(10694)) xor (layer0_outputs(7178));
    outputs(1916) <= (layer0_outputs(4655)) and (layer0_outputs(2034));
    outputs(1917) <= (layer0_outputs(5494)) xor (layer0_outputs(2613));
    outputs(1918) <= (layer0_outputs(9178)) and not (layer0_outputs(8486));
    outputs(1919) <= '0';
    outputs(1920) <= layer0_outputs(4455);
    outputs(1921) <= (layer0_outputs(6333)) and not (layer0_outputs(12466));
    outputs(1922) <= not((layer0_outputs(12293)) xor (layer0_outputs(7733)));
    outputs(1923) <= (layer0_outputs(609)) and (layer0_outputs(599));
    outputs(1924) <= not(layer0_outputs(6163));
    outputs(1925) <= (layer0_outputs(2755)) xor (layer0_outputs(7762));
    outputs(1926) <= not((layer0_outputs(3905)) or (layer0_outputs(11246)));
    outputs(1927) <= (layer0_outputs(529)) or (layer0_outputs(3538));
    outputs(1928) <= not((layer0_outputs(11593)) xor (layer0_outputs(3256)));
    outputs(1929) <= layer0_outputs(681);
    outputs(1930) <= (layer0_outputs(11649)) and not (layer0_outputs(5490));
    outputs(1931) <= not(layer0_outputs(507));
    outputs(1932) <= (layer0_outputs(2998)) and not (layer0_outputs(11082));
    outputs(1933) <= (layer0_outputs(4116)) and not (layer0_outputs(114));
    outputs(1934) <= not((layer0_outputs(4191)) xor (layer0_outputs(2642)));
    outputs(1935) <= (layer0_outputs(2512)) and (layer0_outputs(12244));
    outputs(1936) <= (layer0_outputs(9602)) xor (layer0_outputs(9824));
    outputs(1937) <= not(layer0_outputs(1913));
    outputs(1938) <= (layer0_outputs(5423)) and (layer0_outputs(771));
    outputs(1939) <= not((layer0_outputs(5089)) xor (layer0_outputs(5199)));
    outputs(1940) <= (layer0_outputs(7676)) xor (layer0_outputs(2611));
    outputs(1941) <= (layer0_outputs(3981)) xor (layer0_outputs(4233));
    outputs(1942) <= not((layer0_outputs(6861)) or (layer0_outputs(8202)));
    outputs(1943) <= (layer0_outputs(344)) xor (layer0_outputs(4733));
    outputs(1944) <= (layer0_outputs(6858)) and (layer0_outputs(10636));
    outputs(1945) <= not(layer0_outputs(9220));
    outputs(1946) <= layer0_outputs(1953);
    outputs(1947) <= not((layer0_outputs(12671)) or (layer0_outputs(10474)));
    outputs(1948) <= layer0_outputs(5114);
    outputs(1949) <= (layer0_outputs(9395)) and not (layer0_outputs(3290));
    outputs(1950) <= (layer0_outputs(4909)) xor (layer0_outputs(8638));
    outputs(1951) <= (layer0_outputs(8158)) xor (layer0_outputs(2026));
    outputs(1952) <= '0';
    outputs(1953) <= (layer0_outputs(6509)) and not (layer0_outputs(9490));
    outputs(1954) <= layer0_outputs(10713);
    outputs(1955) <= layer0_outputs(4684);
    outputs(1956) <= (layer0_outputs(6602)) and not (layer0_outputs(7093));
    outputs(1957) <= (layer0_outputs(4897)) and not (layer0_outputs(12684));
    outputs(1958) <= layer0_outputs(10779);
    outputs(1959) <= (layer0_outputs(5910)) and not (layer0_outputs(6506));
    outputs(1960) <= not(layer0_outputs(6851));
    outputs(1961) <= (layer0_outputs(7364)) and (layer0_outputs(11285));
    outputs(1962) <= (layer0_outputs(9569)) xor (layer0_outputs(1863));
    outputs(1963) <= (layer0_outputs(1379)) and not (layer0_outputs(9317));
    outputs(1964) <= layer0_outputs(8924);
    outputs(1965) <= (layer0_outputs(7522)) xor (layer0_outputs(7551));
    outputs(1966) <= layer0_outputs(8893);
    outputs(1967) <= (layer0_outputs(8721)) xor (layer0_outputs(11642));
    outputs(1968) <= (layer0_outputs(12251)) and (layer0_outputs(7169));
    outputs(1969) <= layer0_outputs(9175);
    outputs(1970) <= (layer0_outputs(8434)) xor (layer0_outputs(10606));
    outputs(1971) <= (layer0_outputs(9281)) and not (layer0_outputs(12040));
    outputs(1972) <= layer0_outputs(12258);
    outputs(1973) <= (layer0_outputs(1891)) and (layer0_outputs(8335));
    outputs(1974) <= (layer0_outputs(4823)) and not (layer0_outputs(3966));
    outputs(1975) <= not((layer0_outputs(11887)) or (layer0_outputs(377)));
    outputs(1976) <= layer0_outputs(1837);
    outputs(1977) <= (layer0_outputs(8618)) and not (layer0_outputs(4878));
    outputs(1978) <= layer0_outputs(2257);
    outputs(1979) <= not((layer0_outputs(5911)) xor (layer0_outputs(5081)));
    outputs(1980) <= layer0_outputs(3157);
    outputs(1981) <= (layer0_outputs(12352)) and not (layer0_outputs(11337));
    outputs(1982) <= (layer0_outputs(1395)) and not (layer0_outputs(1482));
    outputs(1983) <= not((layer0_outputs(5838)) xor (layer0_outputs(5800)));
    outputs(1984) <= not(layer0_outputs(10376));
    outputs(1985) <= (layer0_outputs(6507)) and not (layer0_outputs(3682));
    outputs(1986) <= layer0_outputs(10208);
    outputs(1987) <= (layer0_outputs(4887)) and not (layer0_outputs(11811));
    outputs(1988) <= not(layer0_outputs(4347));
    outputs(1989) <= not((layer0_outputs(2241)) and (layer0_outputs(4183)));
    outputs(1990) <= not(layer0_outputs(759));
    outputs(1991) <= not((layer0_outputs(10284)) or (layer0_outputs(10621)));
    outputs(1992) <= not((layer0_outputs(4084)) or (layer0_outputs(2091)));
    outputs(1993) <= layer0_outputs(10016);
    outputs(1994) <= not(layer0_outputs(9326)) or (layer0_outputs(4646));
    outputs(1995) <= not(layer0_outputs(3653));
    outputs(1996) <= (layer0_outputs(9648)) xor (layer0_outputs(8604));
    outputs(1997) <= (layer0_outputs(2077)) and not (layer0_outputs(11777));
    outputs(1998) <= layer0_outputs(4839);
    outputs(1999) <= not((layer0_outputs(12015)) xor (layer0_outputs(12103)));
    outputs(2000) <= layer0_outputs(11834);
    outputs(2001) <= not((layer0_outputs(7501)) or (layer0_outputs(1995)));
    outputs(2002) <= (layer0_outputs(1396)) and not (layer0_outputs(11516));
    outputs(2003) <= layer0_outputs(8071);
    outputs(2004) <= not((layer0_outputs(12195)) xor (layer0_outputs(4364)));
    outputs(2005) <= not((layer0_outputs(8256)) or (layer0_outputs(6120)));
    outputs(2006) <= layer0_outputs(1951);
    outputs(2007) <= not((layer0_outputs(3606)) xor (layer0_outputs(4446)));
    outputs(2008) <= (layer0_outputs(12670)) xor (layer0_outputs(7311));
    outputs(2009) <= not((layer0_outputs(5884)) or (layer0_outputs(7503)));
    outputs(2010) <= layer0_outputs(5495);
    outputs(2011) <= (layer0_outputs(1863)) and not (layer0_outputs(7193));
    outputs(2012) <= not(layer0_outputs(6328));
    outputs(2013) <= not((layer0_outputs(6332)) xor (layer0_outputs(9802)));
    outputs(2014) <= '0';
    outputs(2015) <= (layer0_outputs(397)) and not (layer0_outputs(9312));
    outputs(2016) <= layer0_outputs(2404);
    outputs(2017) <= (layer0_outputs(1673)) xor (layer0_outputs(9098));
    outputs(2018) <= (layer0_outputs(9875)) and (layer0_outputs(10045));
    outputs(2019) <= not((layer0_outputs(1584)) xor (layer0_outputs(9931)));
    outputs(2020) <= (layer0_outputs(2018)) and not (layer0_outputs(10147));
    outputs(2021) <= (layer0_outputs(5584)) and not (layer0_outputs(9136));
    outputs(2022) <= not((layer0_outputs(7685)) xor (layer0_outputs(4393)));
    outputs(2023) <= (layer0_outputs(4221)) and not (layer0_outputs(6349));
    outputs(2024) <= (layer0_outputs(1265)) and not (layer0_outputs(10269));
    outputs(2025) <= not((layer0_outputs(10288)) and (layer0_outputs(203)));
    outputs(2026) <= not(layer0_outputs(3110));
    outputs(2027) <= not((layer0_outputs(274)) xor (layer0_outputs(4915)));
    outputs(2028) <= layer0_outputs(4567);
    outputs(2029) <= (layer0_outputs(4616)) and not (layer0_outputs(5326));
    outputs(2030) <= not(layer0_outputs(7332));
    outputs(2031) <= (layer0_outputs(4124)) or (layer0_outputs(3702));
    outputs(2032) <= layer0_outputs(11834);
    outputs(2033) <= layer0_outputs(2679);
    outputs(2034) <= (layer0_outputs(6959)) and not (layer0_outputs(6381));
    outputs(2035) <= not((layer0_outputs(4436)) xor (layer0_outputs(153)));
    outputs(2036) <= not(layer0_outputs(9766));
    outputs(2037) <= not((layer0_outputs(6599)) xor (layer0_outputs(11703)));
    outputs(2038) <= not((layer0_outputs(10051)) xor (layer0_outputs(3334)));
    outputs(2039) <= (layer0_outputs(8955)) and (layer0_outputs(6417));
    outputs(2040) <= (layer0_outputs(9628)) and not (layer0_outputs(2141));
    outputs(2041) <= not((layer0_outputs(6141)) or (layer0_outputs(6898)));
    outputs(2042) <= layer0_outputs(1144);
    outputs(2043) <= (layer0_outputs(5177)) and (layer0_outputs(5394));
    outputs(2044) <= (layer0_outputs(11396)) xor (layer0_outputs(12690));
    outputs(2045) <= not(layer0_outputs(8018));
    outputs(2046) <= not((layer0_outputs(7178)) or (layer0_outputs(11724)));
    outputs(2047) <= layer0_outputs(10066);
    outputs(2048) <= not(layer0_outputs(6215));
    outputs(2049) <= not((layer0_outputs(6058)) and (layer0_outputs(5344)));
    outputs(2050) <= (layer0_outputs(8847)) and not (layer0_outputs(11196));
    outputs(2051) <= not((layer0_outputs(11710)) xor (layer0_outputs(2972)));
    outputs(2052) <= (layer0_outputs(11813)) and not (layer0_outputs(12766));
    outputs(2053) <= not(layer0_outputs(4501));
    outputs(2054) <= (layer0_outputs(2409)) xor (layer0_outputs(1309));
    outputs(2055) <= (layer0_outputs(3572)) and not (layer0_outputs(3080));
    outputs(2056) <= (layer0_outputs(1985)) and not (layer0_outputs(8728));
    outputs(2057) <= (layer0_outputs(787)) and not (layer0_outputs(641));
    outputs(2058) <= (layer0_outputs(1283)) and not (layer0_outputs(5413));
    outputs(2059) <= (layer0_outputs(3572)) and (layer0_outputs(6487));
    outputs(2060) <= not(layer0_outputs(7469));
    outputs(2061) <= (layer0_outputs(8084)) and not (layer0_outputs(1321));
    outputs(2062) <= (layer0_outputs(4630)) xor (layer0_outputs(5799));
    outputs(2063) <= (layer0_outputs(3261)) and (layer0_outputs(8846));
    outputs(2064) <= not((layer0_outputs(9055)) or (layer0_outputs(857)));
    outputs(2065) <= layer0_outputs(7187);
    outputs(2066) <= not((layer0_outputs(11540)) or (layer0_outputs(8270)));
    outputs(2067) <= layer0_outputs(10578);
    outputs(2068) <= not((layer0_outputs(2505)) xor (layer0_outputs(11390)));
    outputs(2069) <= not(layer0_outputs(5591));
    outputs(2070) <= layer0_outputs(10954);
    outputs(2071) <= not((layer0_outputs(3001)) xor (layer0_outputs(5745)));
    outputs(2072) <= not((layer0_outputs(11971)) xor (layer0_outputs(11725)));
    outputs(2073) <= (layer0_outputs(8478)) and not (layer0_outputs(7309));
    outputs(2074) <= (layer0_outputs(1756)) and (layer0_outputs(4818));
    outputs(2075) <= not(layer0_outputs(2812));
    outputs(2076) <= (layer0_outputs(7207)) and not (layer0_outputs(10420));
    outputs(2077) <= not(layer0_outputs(6643));
    outputs(2078) <= not((layer0_outputs(12394)) and (layer0_outputs(2367)));
    outputs(2079) <= (layer0_outputs(1344)) and (layer0_outputs(3601));
    outputs(2080) <= (layer0_outputs(12468)) and not (layer0_outputs(12112));
    outputs(2081) <= not((layer0_outputs(10024)) or (layer0_outputs(1621)));
    outputs(2082) <= layer0_outputs(4098);
    outputs(2083) <= not(layer0_outputs(12401));
    outputs(2084) <= layer0_outputs(608);
    outputs(2085) <= (layer0_outputs(6855)) xor (layer0_outputs(2286));
    outputs(2086) <= layer0_outputs(10488);
    outputs(2087) <= (layer0_outputs(4950)) and (layer0_outputs(9927));
    outputs(2088) <= (layer0_outputs(131)) and not (layer0_outputs(12001));
    outputs(2089) <= layer0_outputs(7129);
    outputs(2090) <= not(layer0_outputs(820));
    outputs(2091) <= (layer0_outputs(2796)) xor (layer0_outputs(9426));
    outputs(2092) <= not(layer0_outputs(6695));
    outputs(2093) <= not((layer0_outputs(2094)) xor (layer0_outputs(7946)));
    outputs(2094) <= layer0_outputs(11630);
    outputs(2095) <= (layer0_outputs(2530)) xor (layer0_outputs(9002));
    outputs(2096) <= not((layer0_outputs(12476)) and (layer0_outputs(4094)));
    outputs(2097) <= (layer0_outputs(8130)) and not (layer0_outputs(7549));
    outputs(2098) <= not(layer0_outputs(166));
    outputs(2099) <= (layer0_outputs(11739)) and not (layer0_outputs(4040));
    outputs(2100) <= (layer0_outputs(1764)) and (layer0_outputs(2007));
    outputs(2101) <= (layer0_outputs(11824)) xor (layer0_outputs(10337));
    outputs(2102) <= not((layer0_outputs(6702)) xor (layer0_outputs(5640)));
    outputs(2103) <= layer0_outputs(9992);
    outputs(2104) <= (layer0_outputs(12097)) xor (layer0_outputs(2747));
    outputs(2105) <= layer0_outputs(12584);
    outputs(2106) <= (layer0_outputs(2745)) and not (layer0_outputs(4848));
    outputs(2107) <= layer0_outputs(601);
    outputs(2108) <= '0';
    outputs(2109) <= not(layer0_outputs(2980));
    outputs(2110) <= (layer0_outputs(6345)) and not (layer0_outputs(3216));
    outputs(2111) <= (layer0_outputs(6615)) xor (layer0_outputs(9512));
    outputs(2112) <= (layer0_outputs(10192)) and (layer0_outputs(2934));
    outputs(2113) <= '0';
    outputs(2114) <= layer0_outputs(11725);
    outputs(2115) <= (layer0_outputs(3051)) and (layer0_outputs(343));
    outputs(2116) <= not((layer0_outputs(3575)) xor (layer0_outputs(7246)));
    outputs(2117) <= not((layer0_outputs(10682)) or (layer0_outputs(8927)));
    outputs(2118) <= (layer0_outputs(1537)) and not (layer0_outputs(11322));
    outputs(2119) <= not((layer0_outputs(9843)) xor (layer0_outputs(6204)));
    outputs(2120) <= (layer0_outputs(8774)) and not (layer0_outputs(3939));
    outputs(2121) <= not(layer0_outputs(5036));
    outputs(2122) <= not((layer0_outputs(10916)) or (layer0_outputs(12750)));
    outputs(2123) <= not((layer0_outputs(11563)) xor (layer0_outputs(6858)));
    outputs(2124) <= not((layer0_outputs(10908)) xor (layer0_outputs(6239)));
    outputs(2125) <= (layer0_outputs(8371)) and not (layer0_outputs(12642));
    outputs(2126) <= not((layer0_outputs(146)) or (layer0_outputs(1921)));
    outputs(2127) <= (layer0_outputs(5549)) and not (layer0_outputs(1567));
    outputs(2128) <= not(layer0_outputs(9701));
    outputs(2129) <= layer0_outputs(11248);
    outputs(2130) <= not(layer0_outputs(5266));
    outputs(2131) <= not((layer0_outputs(4667)) and (layer0_outputs(12647)));
    outputs(2132) <= (layer0_outputs(10557)) xor (layer0_outputs(10801));
    outputs(2133) <= (layer0_outputs(5136)) and not (layer0_outputs(10854));
    outputs(2134) <= (layer0_outputs(3377)) xor (layer0_outputs(7452));
    outputs(2135) <= (layer0_outputs(7186)) and not (layer0_outputs(12495));
    outputs(2136) <= (layer0_outputs(1100)) and not (layer0_outputs(1223));
    outputs(2137) <= layer0_outputs(11899);
    outputs(2138) <= (layer0_outputs(1803)) and not (layer0_outputs(8500));
    outputs(2139) <= not(layer0_outputs(4084));
    outputs(2140) <= not(layer0_outputs(9617));
    outputs(2141) <= (layer0_outputs(6077)) and not (layer0_outputs(8131));
    outputs(2142) <= layer0_outputs(10548);
    outputs(2143) <= not((layer0_outputs(5168)) or (layer0_outputs(5407)));
    outputs(2144) <= layer0_outputs(9652);
    outputs(2145) <= not((layer0_outputs(5113)) xor (layer0_outputs(3468)));
    outputs(2146) <= not((layer0_outputs(12686)) or (layer0_outputs(4833)));
    outputs(2147) <= (layer0_outputs(9025)) xor (layer0_outputs(12304));
    outputs(2148) <= (layer0_outputs(5987)) and not (layer0_outputs(9035));
    outputs(2149) <= (layer0_outputs(5726)) and not (layer0_outputs(5341));
    outputs(2150) <= (layer0_outputs(9412)) and not (layer0_outputs(11029));
    outputs(2151) <= not(layer0_outputs(10685));
    outputs(2152) <= not(layer0_outputs(6146));
    outputs(2153) <= (layer0_outputs(6521)) and (layer0_outputs(4538));
    outputs(2154) <= layer0_outputs(3849);
    outputs(2155) <= not(layer0_outputs(12556));
    outputs(2156) <= not((layer0_outputs(2170)) or (layer0_outputs(4859)));
    outputs(2157) <= layer0_outputs(11940);
    outputs(2158) <= '0';
    outputs(2159) <= not(layer0_outputs(8845));
    outputs(2160) <= layer0_outputs(7074);
    outputs(2161) <= layer0_outputs(11752);
    outputs(2162) <= (layer0_outputs(1383)) and (layer0_outputs(1937));
    outputs(2163) <= not((layer0_outputs(9553)) or (layer0_outputs(4034)));
    outputs(2164) <= layer0_outputs(1737);
    outputs(2165) <= (layer0_outputs(9949)) and (layer0_outputs(10929));
    outputs(2166) <= not((layer0_outputs(11852)) xor (layer0_outputs(4596)));
    outputs(2167) <= (layer0_outputs(10273)) and not (layer0_outputs(4268));
    outputs(2168) <= (layer0_outputs(8443)) and (layer0_outputs(9171));
    outputs(2169) <= '0';
    outputs(2170) <= (layer0_outputs(8425)) or (layer0_outputs(1706));
    outputs(2171) <= not((layer0_outputs(9256)) or (layer0_outputs(6475)));
    outputs(2172) <= not((layer0_outputs(4936)) xor (layer0_outputs(1532)));
    outputs(2173) <= (layer0_outputs(9194)) and not (layer0_outputs(8182));
    outputs(2174) <= (layer0_outputs(8566)) xor (layer0_outputs(8630));
    outputs(2175) <= not(layer0_outputs(11499));
    outputs(2176) <= layer0_outputs(405);
    outputs(2177) <= (layer0_outputs(1258)) and not (layer0_outputs(10505));
    outputs(2178) <= layer0_outputs(3961);
    outputs(2179) <= not((layer0_outputs(12741)) xor (layer0_outputs(12694)));
    outputs(2180) <= (layer0_outputs(8048)) xor (layer0_outputs(2165));
    outputs(2181) <= not((layer0_outputs(10875)) xor (layer0_outputs(8658)));
    outputs(2182) <= (layer0_outputs(1067)) xor (layer0_outputs(9258));
    outputs(2183) <= (layer0_outputs(6261)) xor (layer0_outputs(4268));
    outputs(2184) <= (layer0_outputs(2082)) xor (layer0_outputs(445));
    outputs(2185) <= not((layer0_outputs(5654)) or (layer0_outputs(1190)));
    outputs(2186) <= not(layer0_outputs(11152));
    outputs(2187) <= (layer0_outputs(1427)) xor (layer0_outputs(5695));
    outputs(2188) <= not((layer0_outputs(12429)) or (layer0_outputs(9186)));
    outputs(2189) <= not((layer0_outputs(4007)) or (layer0_outputs(6718)));
    outputs(2190) <= not((layer0_outputs(9105)) xor (layer0_outputs(12003)));
    outputs(2191) <= (layer0_outputs(322)) and (layer0_outputs(452));
    outputs(2192) <= not((layer0_outputs(4216)) xor (layer0_outputs(13)));
    outputs(2193) <= not(layer0_outputs(4439));
    outputs(2194) <= layer0_outputs(7147);
    outputs(2195) <= not((layer0_outputs(482)) or (layer0_outputs(4500)));
    outputs(2196) <= not((layer0_outputs(8782)) and (layer0_outputs(12009)));
    outputs(2197) <= (layer0_outputs(12069)) and not (layer0_outputs(47));
    outputs(2198) <= (layer0_outputs(2591)) and (layer0_outputs(5962));
    outputs(2199) <= not((layer0_outputs(12130)) xor (layer0_outputs(9948)));
    outputs(2200) <= layer0_outputs(6354);
    outputs(2201) <= layer0_outputs(2348);
    outputs(2202) <= layer0_outputs(7175);
    outputs(2203) <= not(layer0_outputs(3928));
    outputs(2204) <= not(layer0_outputs(8028));
    outputs(2205) <= layer0_outputs(9715);
    outputs(2206) <= not(layer0_outputs(9962));
    outputs(2207) <= not((layer0_outputs(10527)) xor (layer0_outputs(10148)));
    outputs(2208) <= layer0_outputs(2550);
    outputs(2209) <= '1';
    outputs(2210) <= (layer0_outputs(12039)) and not (layer0_outputs(1422));
    outputs(2211) <= (layer0_outputs(53)) and not (layer0_outputs(12191));
    outputs(2212) <= (layer0_outputs(11058)) xor (layer0_outputs(3798));
    outputs(2213) <= not((layer0_outputs(6619)) or (layer0_outputs(76)));
    outputs(2214) <= (layer0_outputs(2518)) and not (layer0_outputs(4468));
    outputs(2215) <= not((layer0_outputs(297)) and (layer0_outputs(8933)));
    outputs(2216) <= not((layer0_outputs(8484)) xor (layer0_outputs(1553)));
    outputs(2217) <= layer0_outputs(1136);
    outputs(2218) <= not(layer0_outputs(10406));
    outputs(2219) <= (layer0_outputs(3641)) and (layer0_outputs(693));
    outputs(2220) <= not((layer0_outputs(3105)) xor (layer0_outputs(7597)));
    outputs(2221) <= (layer0_outputs(2711)) and not (layer0_outputs(10061));
    outputs(2222) <= (layer0_outputs(6211)) and not (layer0_outputs(129));
    outputs(2223) <= not(layer0_outputs(2780));
    outputs(2224) <= not((layer0_outputs(9874)) or (layer0_outputs(876)));
    outputs(2225) <= layer0_outputs(3498);
    outputs(2226) <= not(layer0_outputs(10041));
    outputs(2227) <= not((layer0_outputs(1585)) xor (layer0_outputs(10582)));
    outputs(2228) <= not((layer0_outputs(9627)) or (layer0_outputs(10404)));
    outputs(2229) <= layer0_outputs(19);
    outputs(2230) <= (layer0_outputs(10315)) and (layer0_outputs(12301));
    outputs(2231) <= not((layer0_outputs(11233)) xor (layer0_outputs(5955)));
    outputs(2232) <= '0';
    outputs(2233) <= not((layer0_outputs(9812)) xor (layer0_outputs(11731)));
    outputs(2234) <= not(layer0_outputs(338));
    outputs(2235) <= not((layer0_outputs(6419)) or (layer0_outputs(10240)));
    outputs(2236) <= not((layer0_outputs(2130)) xor (layer0_outputs(3533)));
    outputs(2237) <= (layer0_outputs(3585)) xor (layer0_outputs(8868));
    outputs(2238) <= not((layer0_outputs(4163)) and (layer0_outputs(10427)));
    outputs(2239) <= (layer0_outputs(10995)) and (layer0_outputs(10598));
    outputs(2240) <= not((layer0_outputs(2800)) xor (layer0_outputs(12790)));
    outputs(2241) <= (layer0_outputs(5620)) and not (layer0_outputs(1635));
    outputs(2242) <= (layer0_outputs(10175)) and not (layer0_outputs(900));
    outputs(2243) <= not(layer0_outputs(251)) or (layer0_outputs(4567));
    outputs(2244) <= not(layer0_outputs(3556));
    outputs(2245) <= layer0_outputs(9020);
    outputs(2246) <= not((layer0_outputs(11302)) xor (layer0_outputs(11195)));
    outputs(2247) <= (layer0_outputs(11098)) xor (layer0_outputs(3412));
    outputs(2248) <= not((layer0_outputs(6846)) xor (layer0_outputs(8540)));
    outputs(2249) <= not((layer0_outputs(2005)) or (layer0_outputs(8234)));
    outputs(2250) <= (layer0_outputs(12724)) and not (layer0_outputs(739));
    outputs(2251) <= layer0_outputs(11065);
    outputs(2252) <= (layer0_outputs(7040)) and (layer0_outputs(4641));
    outputs(2253) <= (layer0_outputs(3553)) and (layer0_outputs(11051));
    outputs(2254) <= not((layer0_outputs(2947)) xor (layer0_outputs(2737)));
    outputs(2255) <= not((layer0_outputs(409)) or (layer0_outputs(3230)));
    outputs(2256) <= (layer0_outputs(8238)) and not (layer0_outputs(12030));
    outputs(2257) <= (layer0_outputs(7446)) xor (layer0_outputs(9939));
    outputs(2258) <= not(layer0_outputs(4612));
    outputs(2259) <= not((layer0_outputs(2795)) or (layer0_outputs(5077)));
    outputs(2260) <= not(layer0_outputs(8317));
    outputs(2261) <= not(layer0_outputs(4628));
    outputs(2262) <= not((layer0_outputs(10951)) xor (layer0_outputs(144)));
    outputs(2263) <= layer0_outputs(4182);
    outputs(2264) <= layer0_outputs(5002);
    outputs(2265) <= not(layer0_outputs(160));
    outputs(2266) <= '0';
    outputs(2267) <= not((layer0_outputs(12302)) or (layer0_outputs(3885)));
    outputs(2268) <= not((layer0_outputs(4195)) or (layer0_outputs(11487)));
    outputs(2269) <= (layer0_outputs(7218)) xor (layer0_outputs(6587));
    outputs(2270) <= (layer0_outputs(7615)) and not (layer0_outputs(9990));
    outputs(2271) <= (layer0_outputs(7791)) and (layer0_outputs(9403));
    outputs(2272) <= layer0_outputs(568);
    outputs(2273) <= (layer0_outputs(8020)) or (layer0_outputs(4349));
    outputs(2274) <= not((layer0_outputs(2339)) xor (layer0_outputs(6907)));
    outputs(2275) <= layer0_outputs(11539);
    outputs(2276) <= not(layer0_outputs(39));
    outputs(2277) <= layer0_outputs(9293);
    outputs(2278) <= (layer0_outputs(1774)) xor (layer0_outputs(9826));
    outputs(2279) <= not((layer0_outputs(11955)) or (layer0_outputs(5836)));
    outputs(2280) <= (layer0_outputs(9203)) and not (layer0_outputs(7555));
    outputs(2281) <= not(layer0_outputs(3420));
    outputs(2282) <= (layer0_outputs(7122)) and not (layer0_outputs(7448));
    outputs(2283) <= (layer0_outputs(12020)) and not (layer0_outputs(1561));
    outputs(2284) <= (layer0_outputs(10052)) and not (layer0_outputs(4919));
    outputs(2285) <= layer0_outputs(9499);
    outputs(2286) <= not(layer0_outputs(5120));
    outputs(2287) <= layer0_outputs(7472);
    outputs(2288) <= not((layer0_outputs(4838)) xor (layer0_outputs(4395)));
    outputs(2289) <= not((layer0_outputs(1770)) xor (layer0_outputs(10012)));
    outputs(2290) <= not(layer0_outputs(6908));
    outputs(2291) <= (layer0_outputs(11323)) xor (layer0_outputs(7296));
    outputs(2292) <= not((layer0_outputs(10768)) or (layer0_outputs(1018)));
    outputs(2293) <= layer0_outputs(804);
    outputs(2294) <= not(layer0_outputs(6150));
    outputs(2295) <= (layer0_outputs(92)) xor (layer0_outputs(8790));
    outputs(2296) <= (layer0_outputs(6595)) and not (layer0_outputs(3234));
    outputs(2297) <= (layer0_outputs(3453)) xor (layer0_outputs(1097));
    outputs(2298) <= not((layer0_outputs(4994)) xor (layer0_outputs(2399)));
    outputs(2299) <= layer0_outputs(311);
    outputs(2300) <= not(layer0_outputs(4147));
    outputs(2301) <= not((layer0_outputs(4047)) xor (layer0_outputs(8608)));
    outputs(2302) <= not(layer0_outputs(3872));
    outputs(2303) <= layer0_outputs(12202);
    outputs(2304) <= layer0_outputs(8157);
    outputs(2305) <= not((layer0_outputs(6138)) or (layer0_outputs(3234)));
    outputs(2306) <= layer0_outputs(9485);
    outputs(2307) <= not((layer0_outputs(8095)) or (layer0_outputs(5520)));
    outputs(2308) <= layer0_outputs(5837);
    outputs(2309) <= not(layer0_outputs(5490));
    outputs(2310) <= layer0_outputs(8880);
    outputs(2311) <= (layer0_outputs(4071)) xor (layer0_outputs(11933));
    outputs(2312) <= layer0_outputs(4968);
    outputs(2313) <= (layer0_outputs(7704)) xor (layer0_outputs(6679));
    outputs(2314) <= layer0_outputs(7657);
    outputs(2315) <= (layer0_outputs(1413)) and (layer0_outputs(4236));
    outputs(2316) <= not(layer0_outputs(10955));
    outputs(2317) <= not(layer0_outputs(9150));
    outputs(2318) <= (layer0_outputs(5775)) xor (layer0_outputs(5766));
    outputs(2319) <= not((layer0_outputs(8777)) or (layer0_outputs(1722)));
    outputs(2320) <= (layer0_outputs(7246)) xor (layer0_outputs(2567));
    outputs(2321) <= not((layer0_outputs(4344)) xor (layer0_outputs(11258)));
    outputs(2322) <= layer0_outputs(6421);
    outputs(2323) <= not(layer0_outputs(10650));
    outputs(2324) <= not((layer0_outputs(11663)) or (layer0_outputs(11224)));
    outputs(2325) <= layer0_outputs(9089);
    outputs(2326) <= (layer0_outputs(4459)) and not (layer0_outputs(807));
    outputs(2327) <= (layer0_outputs(3679)) and (layer0_outputs(5804));
    outputs(2328) <= (layer0_outputs(11719)) and not (layer0_outputs(8257));
    outputs(2329) <= not(layer0_outputs(2689));
    outputs(2330) <= (layer0_outputs(609)) and not (layer0_outputs(7562));
    outputs(2331) <= not(layer0_outputs(1691));
    outputs(2332) <= (layer0_outputs(9211)) and (layer0_outputs(12449));
    outputs(2333) <= (layer0_outputs(10547)) xor (layer0_outputs(4088));
    outputs(2334) <= (layer0_outputs(9327)) xor (layer0_outputs(7301));
    outputs(2335) <= not(layer0_outputs(12601));
    outputs(2336) <= not(layer0_outputs(7722));
    outputs(2337) <= not(layer0_outputs(5528));
    outputs(2338) <= (layer0_outputs(1628)) and (layer0_outputs(3180));
    outputs(2339) <= not(layer0_outputs(5043));
    outputs(2340) <= not((layer0_outputs(1126)) or (layer0_outputs(3597)));
    outputs(2341) <= (layer0_outputs(223)) and not (layer0_outputs(3746));
    outputs(2342) <= not((layer0_outputs(6195)) or (layer0_outputs(9042)));
    outputs(2343) <= (layer0_outputs(10879)) xor (layer0_outputs(9461));
    outputs(2344) <= not(layer0_outputs(61));
    outputs(2345) <= not(layer0_outputs(2730));
    outputs(2346) <= layer0_outputs(10405);
    outputs(2347) <= layer0_outputs(12213);
    outputs(2348) <= not(layer0_outputs(8043));
    outputs(2349) <= (layer0_outputs(4800)) and not (layer0_outputs(4702));
    outputs(2350) <= not((layer0_outputs(3746)) or (layer0_outputs(5777)));
    outputs(2351) <= not((layer0_outputs(10156)) and (layer0_outputs(9272)));
    outputs(2352) <= not((layer0_outputs(4371)) or (layer0_outputs(4265)));
    outputs(2353) <= layer0_outputs(11696);
    outputs(2354) <= (layer0_outputs(10735)) and (layer0_outputs(9758));
    outputs(2355) <= (layer0_outputs(1503)) and not (layer0_outputs(11919));
    outputs(2356) <= not((layer0_outputs(8835)) or (layer0_outputs(6296)));
    outputs(2357) <= not(layer0_outputs(11000));
    outputs(2358) <= not((layer0_outputs(12528)) xor (layer0_outputs(8951)));
    outputs(2359) <= not(layer0_outputs(12433));
    outputs(2360) <= not((layer0_outputs(10236)) and (layer0_outputs(9312)));
    outputs(2361) <= layer0_outputs(4169);
    outputs(2362) <= not((layer0_outputs(12200)) xor (layer0_outputs(10431)));
    outputs(2363) <= layer0_outputs(10596);
    outputs(2364) <= (layer0_outputs(6674)) and not (layer0_outputs(10823));
    outputs(2365) <= '0';
    outputs(2366) <= (layer0_outputs(8594)) and not (layer0_outputs(8110));
    outputs(2367) <= not((layer0_outputs(2911)) xor (layer0_outputs(11345)));
    outputs(2368) <= layer0_outputs(12765);
    outputs(2369) <= not((layer0_outputs(3238)) or (layer0_outputs(5613)));
    outputs(2370) <= (layer0_outputs(3313)) and (layer0_outputs(2614));
    outputs(2371) <= (layer0_outputs(2922)) and (layer0_outputs(588));
    outputs(2372) <= layer0_outputs(5977);
    outputs(2373) <= not(layer0_outputs(10513));
    outputs(2374) <= layer0_outputs(12272);
    outputs(2375) <= (layer0_outputs(5627)) and not (layer0_outputs(3847));
    outputs(2376) <= not((layer0_outputs(10613)) xor (layer0_outputs(1586)));
    outputs(2377) <= (layer0_outputs(2737)) or (layer0_outputs(627));
    outputs(2378) <= not(layer0_outputs(1997));
    outputs(2379) <= layer0_outputs(8067);
    outputs(2380) <= (layer0_outputs(11506)) and not (layer0_outputs(5122));
    outputs(2381) <= (layer0_outputs(4583)) and not (layer0_outputs(7980));
    outputs(2382) <= (layer0_outputs(11567)) xor (layer0_outputs(10407));
    outputs(2383) <= layer0_outputs(9947);
    outputs(2384) <= not(layer0_outputs(144));
    outputs(2385) <= (layer0_outputs(1148)) and not (layer0_outputs(6244));
    outputs(2386) <= not(layer0_outputs(12501));
    outputs(2387) <= (layer0_outputs(6645)) and not (layer0_outputs(10185));
    outputs(2388) <= (layer0_outputs(6633)) and not (layer0_outputs(8567));
    outputs(2389) <= not((layer0_outputs(8362)) or (layer0_outputs(2218)));
    outputs(2390) <= layer0_outputs(1338);
    outputs(2391) <= layer0_outputs(7061);
    outputs(2392) <= (layer0_outputs(7922)) and not (layer0_outputs(7532));
    outputs(2393) <= (layer0_outputs(11235)) xor (layer0_outputs(2785));
    outputs(2394) <= layer0_outputs(1215);
    outputs(2395) <= not((layer0_outputs(5024)) or (layer0_outputs(1666)));
    outputs(2396) <= (layer0_outputs(8475)) xor (layer0_outputs(3052));
    outputs(2397) <= (layer0_outputs(11089)) and not (layer0_outputs(12720));
    outputs(2398) <= not((layer0_outputs(2725)) xor (layer0_outputs(6092)));
    outputs(2399) <= not((layer0_outputs(12060)) or (layer0_outputs(4087)));
    outputs(2400) <= not(layer0_outputs(5198));
    outputs(2401) <= not(layer0_outputs(1179));
    outputs(2402) <= (layer0_outputs(6433)) and not (layer0_outputs(11916));
    outputs(2403) <= layer0_outputs(1083);
    outputs(2404) <= not((layer0_outputs(6235)) and (layer0_outputs(6834)));
    outputs(2405) <= (layer0_outputs(727)) and not (layer0_outputs(11047));
    outputs(2406) <= layer0_outputs(3789);
    outputs(2407) <= (layer0_outputs(10157)) and not (layer0_outputs(9728));
    outputs(2408) <= (layer0_outputs(4207)) xor (layer0_outputs(1406));
    outputs(2409) <= not((layer0_outputs(8932)) or (layer0_outputs(7325)));
    outputs(2410) <= not((layer0_outputs(7766)) or (layer0_outputs(1949)));
    outputs(2411) <= not((layer0_outputs(1181)) or (layer0_outputs(8873)));
    outputs(2412) <= '0';
    outputs(2413) <= layer0_outputs(10488);
    outputs(2414) <= (layer0_outputs(9650)) and not (layer0_outputs(7979));
    outputs(2415) <= (layer0_outputs(2517)) and not (layer0_outputs(4318));
    outputs(2416) <= (layer0_outputs(384)) and not (layer0_outputs(2880));
    outputs(2417) <= not((layer0_outputs(11295)) xor (layer0_outputs(10187)));
    outputs(2418) <= not(layer0_outputs(8747));
    outputs(2419) <= layer0_outputs(3289);
    outputs(2420) <= not((layer0_outputs(3432)) xor (layer0_outputs(1888)));
    outputs(2421) <= layer0_outputs(7572);
    outputs(2422) <= (layer0_outputs(1687)) and (layer0_outputs(7622));
    outputs(2423) <= not((layer0_outputs(7911)) xor (layer0_outputs(11231)));
    outputs(2424) <= (layer0_outputs(11553)) and not (layer0_outputs(7760));
    outputs(2425) <= not(layer0_outputs(4906));
    outputs(2426) <= not((layer0_outputs(11275)) or (layer0_outputs(11712)));
    outputs(2427) <= layer0_outputs(8647);
    outputs(2428) <= (layer0_outputs(314)) and (layer0_outputs(8318));
    outputs(2429) <= not(layer0_outputs(8290)) or (layer0_outputs(9314));
    outputs(2430) <= (layer0_outputs(149)) and not (layer0_outputs(5592));
    outputs(2431) <= (layer0_outputs(5627)) and not (layer0_outputs(10119));
    outputs(2432) <= (layer0_outputs(1980)) and not (layer0_outputs(1526));
    outputs(2433) <= layer0_outputs(5716);
    outputs(2434) <= not((layer0_outputs(1183)) xor (layer0_outputs(6658)));
    outputs(2435) <= (layer0_outputs(4603)) and not (layer0_outputs(284));
    outputs(2436) <= not(layer0_outputs(7158));
    outputs(2437) <= not(layer0_outputs(11437));
    outputs(2438) <= not((layer0_outputs(2705)) or (layer0_outputs(4858)));
    outputs(2439) <= not(layer0_outputs(750));
    outputs(2440) <= not((layer0_outputs(3768)) or (layer0_outputs(8644)));
    outputs(2441) <= (layer0_outputs(436)) and not (layer0_outputs(8185));
    outputs(2442) <= '1';
    outputs(2443) <= layer0_outputs(10225);
    outputs(2444) <= not((layer0_outputs(6372)) xor (layer0_outputs(7320)));
    outputs(2445) <= not((layer0_outputs(12340)) xor (layer0_outputs(497)));
    outputs(2446) <= not(layer0_outputs(3452));
    outputs(2447) <= not((layer0_outputs(8979)) and (layer0_outputs(8028)));
    outputs(2448) <= (layer0_outputs(10632)) and not (layer0_outputs(7908));
    outputs(2449) <= layer0_outputs(12384);
    outputs(2450) <= (layer0_outputs(1247)) and not (layer0_outputs(3251));
    outputs(2451) <= (layer0_outputs(12175)) and not (layer0_outputs(3386));
    outputs(2452) <= not((layer0_outputs(5931)) or (layer0_outputs(5356)));
    outputs(2453) <= not((layer0_outputs(1309)) xor (layer0_outputs(7461)));
    outputs(2454) <= (layer0_outputs(161)) and not (layer0_outputs(6175));
    outputs(2455) <= (layer0_outputs(9609)) and not (layer0_outputs(7021));
    outputs(2456) <= layer0_outputs(2415);
    outputs(2457) <= (layer0_outputs(4490)) xor (layer0_outputs(12613));
    outputs(2458) <= not((layer0_outputs(6464)) or (layer0_outputs(3939)));
    outputs(2459) <= layer0_outputs(12575);
    outputs(2460) <= layer0_outputs(6592);
    outputs(2461) <= (layer0_outputs(10211)) and not (layer0_outputs(259));
    outputs(2462) <= (layer0_outputs(6827)) and not (layer0_outputs(10134));
    outputs(2463) <= '0';
    outputs(2464) <= not(layer0_outputs(12533));
    outputs(2465) <= layer0_outputs(528);
    outputs(2466) <= not(layer0_outputs(576));
    outputs(2467) <= layer0_outputs(2313);
    outputs(2468) <= not((layer0_outputs(1634)) xor (layer0_outputs(5491)));
    outputs(2469) <= (layer0_outputs(11932)) and (layer0_outputs(10100));
    outputs(2470) <= (layer0_outputs(11590)) and not (layer0_outputs(911));
    outputs(2471) <= (layer0_outputs(3796)) and not (layer0_outputs(6939));
    outputs(2472) <= layer0_outputs(2779);
    outputs(2473) <= layer0_outputs(3310);
    outputs(2474) <= (layer0_outputs(12344)) xor (layer0_outputs(7485));
    outputs(2475) <= layer0_outputs(6901);
    outputs(2476) <= not(layer0_outputs(504));
    outputs(2477) <= layer0_outputs(12719);
    outputs(2478) <= not(layer0_outputs(3084));
    outputs(2479) <= not(layer0_outputs(862));
    outputs(2480) <= not((layer0_outputs(2182)) xor (layer0_outputs(2318)));
    outputs(2481) <= not(layer0_outputs(1245));
    outputs(2482) <= (layer0_outputs(699)) and not (layer0_outputs(7036));
    outputs(2483) <= (layer0_outputs(8739)) and (layer0_outputs(12567));
    outputs(2484) <= not(layer0_outputs(5792));
    outputs(2485) <= layer0_outputs(11749);
    outputs(2486) <= layer0_outputs(4293);
    outputs(2487) <= (layer0_outputs(8741)) and not (layer0_outputs(6660));
    outputs(2488) <= not((layer0_outputs(905)) and (layer0_outputs(172)));
    outputs(2489) <= layer0_outputs(4873);
    outputs(2490) <= not((layer0_outputs(11787)) xor (layer0_outputs(8179)));
    outputs(2491) <= layer0_outputs(10632);
    outputs(2492) <= layer0_outputs(11531);
    outputs(2493) <= (layer0_outputs(544)) and (layer0_outputs(6562));
    outputs(2494) <= '0';
    outputs(2495) <= not((layer0_outputs(8966)) xor (layer0_outputs(2871)));
    outputs(2496) <= (layer0_outputs(364)) xor (layer0_outputs(8407));
    outputs(2497) <= '0';
    outputs(2498) <= layer0_outputs(3424);
    outputs(2499) <= layer0_outputs(12009);
    outputs(2500) <= (layer0_outputs(9288)) and (layer0_outputs(9510));
    outputs(2501) <= not(layer0_outputs(9230));
    outputs(2502) <= (layer0_outputs(777)) and not (layer0_outputs(4165));
    outputs(2503) <= not(layer0_outputs(4419));
    outputs(2504) <= (layer0_outputs(5008)) and not (layer0_outputs(9705));
    outputs(2505) <= not(layer0_outputs(12452));
    outputs(2506) <= (layer0_outputs(635)) and (layer0_outputs(10000));
    outputs(2507) <= not((layer0_outputs(4409)) or (layer0_outputs(12782)));
    outputs(2508) <= not((layer0_outputs(1255)) xor (layer0_outputs(6949)));
    outputs(2509) <= layer0_outputs(5000);
    outputs(2510) <= layer0_outputs(6795);
    outputs(2511) <= not(layer0_outputs(10517));
    outputs(2512) <= not((layer0_outputs(11071)) xor (layer0_outputs(9817)));
    outputs(2513) <= not(layer0_outputs(4477));
    outputs(2514) <= layer0_outputs(9069);
    outputs(2515) <= not((layer0_outputs(10051)) xor (layer0_outputs(314)));
    outputs(2516) <= not((layer0_outputs(5498)) or (layer0_outputs(977)));
    outputs(2517) <= not(layer0_outputs(8624));
    outputs(2518) <= not((layer0_outputs(8373)) xor (layer0_outputs(7308)));
    outputs(2519) <= (layer0_outputs(2311)) and not (layer0_outputs(8686));
    outputs(2520) <= not(layer0_outputs(5663));
    outputs(2521) <= (layer0_outputs(5943)) and not (layer0_outputs(12368));
    outputs(2522) <= '0';
    outputs(2523) <= not(layer0_outputs(4795)) or (layer0_outputs(8192));
    outputs(2524) <= not(layer0_outputs(7173));
    outputs(2525) <= layer0_outputs(5679);
    outputs(2526) <= not(layer0_outputs(9479));
    outputs(2527) <= (layer0_outputs(4584)) and (layer0_outputs(10213));
    outputs(2528) <= not(layer0_outputs(174));
    outputs(2529) <= (layer0_outputs(342)) and not (layer0_outputs(3184));
    outputs(2530) <= layer0_outputs(12125);
    outputs(2531) <= not(layer0_outputs(7099));
    outputs(2532) <= not((layer0_outputs(11398)) xor (layer0_outputs(10060)));
    outputs(2533) <= not((layer0_outputs(9506)) xor (layer0_outputs(5974)));
    outputs(2534) <= (layer0_outputs(11113)) and not (layer0_outputs(6267));
    outputs(2535) <= not(layer0_outputs(4957));
    outputs(2536) <= (layer0_outputs(10643)) and (layer0_outputs(10918));
    outputs(2537) <= not((layer0_outputs(652)) or (layer0_outputs(110)));
    outputs(2538) <= not(layer0_outputs(8400));
    outputs(2539) <= (layer0_outputs(6094)) and not (layer0_outputs(2802));
    outputs(2540) <= layer0_outputs(5585);
    outputs(2541) <= (layer0_outputs(8312)) xor (layer0_outputs(12139));
    outputs(2542) <= layer0_outputs(7885);
    outputs(2543) <= not((layer0_outputs(5970)) xor (layer0_outputs(6912)));
    outputs(2544) <= layer0_outputs(5424);
    outputs(2545) <= not((layer0_outputs(8535)) xor (layer0_outputs(9737)));
    outputs(2546) <= layer0_outputs(2273);
    outputs(2547) <= (layer0_outputs(8967)) xor (layer0_outputs(11760));
    outputs(2548) <= layer0_outputs(8246);
    outputs(2549) <= not(layer0_outputs(3854));
    outputs(2550) <= not(layer0_outputs(1006));
    outputs(2551) <= layer0_outputs(11157);
    outputs(2552) <= not((layer0_outputs(8871)) xor (layer0_outputs(450)));
    outputs(2553) <= not((layer0_outputs(7092)) xor (layer0_outputs(12561)));
    outputs(2554) <= layer0_outputs(9633);
    outputs(2555) <= (layer0_outputs(10380)) and (layer0_outputs(1768));
    outputs(2556) <= (layer0_outputs(5608)) and (layer0_outputs(8208));
    outputs(2557) <= (layer0_outputs(2320)) and not (layer0_outputs(4181));
    outputs(2558) <= (layer0_outputs(6276)) and not (layer0_outputs(11326));
    outputs(2559) <= not(layer0_outputs(3837)) or (layer0_outputs(1253));
    outputs(2560) <= not((layer0_outputs(1955)) xor (layer0_outputs(10316)));
    outputs(2561) <= not((layer0_outputs(11464)) xor (layer0_outputs(2577)));
    outputs(2562) <= not((layer0_outputs(7463)) and (layer0_outputs(11693)));
    outputs(2563) <= not(layer0_outputs(9856));
    outputs(2564) <= layer0_outputs(12264);
    outputs(2565) <= (layer0_outputs(6969)) xor (layer0_outputs(3388));
    outputs(2566) <= not(layer0_outputs(11633)) or (layer0_outputs(5274));
    outputs(2567) <= (layer0_outputs(2367)) or (layer0_outputs(6521));
    outputs(2568) <= '1';
    outputs(2569) <= not(layer0_outputs(7838)) or (layer0_outputs(11627));
    outputs(2570) <= layer0_outputs(10207);
    outputs(2571) <= (layer0_outputs(6666)) and not (layer0_outputs(3321));
    outputs(2572) <= layer0_outputs(10329);
    outputs(2573) <= not(layer0_outputs(11035));
    outputs(2574) <= not(layer0_outputs(9601));
    outputs(2575) <= not(layer0_outputs(110)) or (layer0_outputs(12428));
    outputs(2576) <= (layer0_outputs(7773)) xor (layer0_outputs(4590));
    outputs(2577) <= (layer0_outputs(4805)) and (layer0_outputs(1995));
    outputs(2578) <= not(layer0_outputs(9469));
    outputs(2579) <= not((layer0_outputs(9558)) or (layer0_outputs(6542)));
    outputs(2580) <= layer0_outputs(2081);
    outputs(2581) <= not(layer0_outputs(12520));
    outputs(2582) <= (layer0_outputs(7658)) xor (layer0_outputs(12678));
    outputs(2583) <= (layer0_outputs(4199)) or (layer0_outputs(10116));
    outputs(2584) <= (layer0_outputs(12351)) or (layer0_outputs(2143));
    outputs(2585) <= (layer0_outputs(1296)) xor (layer0_outputs(1999));
    outputs(2586) <= layer0_outputs(10506);
    outputs(2587) <= not(layer0_outputs(6403)) or (layer0_outputs(5672));
    outputs(2588) <= (layer0_outputs(6397)) xor (layer0_outputs(12161));
    outputs(2589) <= (layer0_outputs(7004)) xor (layer0_outputs(6410));
    outputs(2590) <= '1';
    outputs(2591) <= '1';
    outputs(2592) <= (layer0_outputs(7797)) xor (layer0_outputs(3469));
    outputs(2593) <= not((layer0_outputs(5456)) xor (layer0_outputs(11773)));
    outputs(2594) <= not((layer0_outputs(9262)) xor (layer0_outputs(1819)));
    outputs(2595) <= not(layer0_outputs(1238));
    outputs(2596) <= not(layer0_outputs(12759));
    outputs(2597) <= not(layer0_outputs(10505));
    outputs(2598) <= not((layer0_outputs(8499)) or (layer0_outputs(8602)));
    outputs(2599) <= not(layer0_outputs(11485));
    outputs(2600) <= not(layer0_outputs(7833)) or (layer0_outputs(6392));
    outputs(2601) <= not((layer0_outputs(2029)) xor (layer0_outputs(11636)));
    outputs(2602) <= not(layer0_outputs(8390)) or (layer0_outputs(10796));
    outputs(2603) <= layer0_outputs(7054);
    outputs(2604) <= not(layer0_outputs(11953)) or (layer0_outputs(9731));
    outputs(2605) <= (layer0_outputs(2396)) xor (layer0_outputs(6422));
    outputs(2606) <= layer0_outputs(4526);
    outputs(2607) <= layer0_outputs(5001);
    outputs(2608) <= (layer0_outputs(6666)) and not (layer0_outputs(4537));
    outputs(2609) <= (layer0_outputs(10098)) and not (layer0_outputs(9125));
    outputs(2610) <= layer0_outputs(11237);
    outputs(2611) <= (layer0_outputs(2913)) xor (layer0_outputs(8743));
    outputs(2612) <= not((layer0_outputs(1043)) xor (layer0_outputs(286)));
    outputs(2613) <= not(layer0_outputs(12025)) or (layer0_outputs(9738));
    outputs(2614) <= (layer0_outputs(1589)) xor (layer0_outputs(764));
    outputs(2615) <= not(layer0_outputs(8225));
    outputs(2616) <= (layer0_outputs(7704)) xor (layer0_outputs(8242));
    outputs(2617) <= layer0_outputs(7385);
    outputs(2618) <= not((layer0_outputs(3813)) xor (layer0_outputs(8882)));
    outputs(2619) <= (layer0_outputs(11511)) and not (layer0_outputs(10055));
    outputs(2620) <= not((layer0_outputs(4615)) xor (layer0_outputs(309)));
    outputs(2621) <= (layer0_outputs(895)) and not (layer0_outputs(7750));
    outputs(2622) <= not((layer0_outputs(7731)) and (layer0_outputs(11348)));
    outputs(2623) <= not((layer0_outputs(1556)) or (layer0_outputs(7191)));
    outputs(2624) <= (layer0_outputs(3419)) xor (layer0_outputs(2415));
    outputs(2625) <= (layer0_outputs(10007)) xor (layer0_outputs(2430));
    outputs(2626) <= not(layer0_outputs(3213));
    outputs(2627) <= layer0_outputs(6301);
    outputs(2628) <= not(layer0_outputs(7880));
    outputs(2629) <= not((layer0_outputs(5087)) xor (layer0_outputs(7196)));
    outputs(2630) <= layer0_outputs(7259);
    outputs(2631) <= not(layer0_outputs(7848));
    outputs(2632) <= layer0_outputs(1117);
    outputs(2633) <= layer0_outputs(5937);
    outputs(2634) <= not((layer0_outputs(5049)) and (layer0_outputs(2453)));
    outputs(2635) <= not((layer0_outputs(10654)) xor (layer0_outputs(6187)));
    outputs(2636) <= not(layer0_outputs(8361));
    outputs(2637) <= not((layer0_outputs(1080)) xor (layer0_outputs(5336)));
    outputs(2638) <= (layer0_outputs(533)) or (layer0_outputs(10655));
    outputs(2639) <= not(layer0_outputs(8190));
    outputs(2640) <= not((layer0_outputs(11524)) and (layer0_outputs(11066)));
    outputs(2641) <= not((layer0_outputs(10168)) xor (layer0_outputs(7432)));
    outputs(2642) <= not((layer0_outputs(11407)) or (layer0_outputs(380)));
    outputs(2643) <= not((layer0_outputs(12705)) xor (layer0_outputs(6825)));
    outputs(2644) <= not((layer0_outputs(3730)) or (layer0_outputs(2068)));
    outputs(2645) <= layer0_outputs(4378);
    outputs(2646) <= not(layer0_outputs(10231));
    outputs(2647) <= (layer0_outputs(966)) xor (layer0_outputs(3839));
    outputs(2648) <= layer0_outputs(5857);
    outputs(2649) <= not(layer0_outputs(1551));
    outputs(2650) <= layer0_outputs(8621);
    outputs(2651) <= layer0_outputs(55);
    outputs(2652) <= (layer0_outputs(10304)) xor (layer0_outputs(4499));
    outputs(2653) <= layer0_outputs(1175);
    outputs(2654) <= not((layer0_outputs(6351)) and (layer0_outputs(4666)));
    outputs(2655) <= not(layer0_outputs(9868));
    outputs(2656) <= (layer0_outputs(4546)) and not (layer0_outputs(4096));
    outputs(2657) <= layer0_outputs(4335);
    outputs(2658) <= not(layer0_outputs(8787)) or (layer0_outputs(1110));
    outputs(2659) <= not(layer0_outputs(8408));
    outputs(2660) <= not(layer0_outputs(2619));
    outputs(2661) <= (layer0_outputs(3366)) and not (layer0_outputs(12040));
    outputs(2662) <= (layer0_outputs(357)) xor (layer0_outputs(1606));
    outputs(2663) <= not(layer0_outputs(3832)) or (layer0_outputs(6413));
    outputs(2664) <= layer0_outputs(5480);
    outputs(2665) <= (layer0_outputs(10281)) and (layer0_outputs(11990));
    outputs(2666) <= (layer0_outputs(9668)) or (layer0_outputs(7206));
    outputs(2667) <= (layer0_outputs(5310)) and (layer0_outputs(5891));
    outputs(2668) <= not(layer0_outputs(3534)) or (layer0_outputs(307));
    outputs(2669) <= not((layer0_outputs(394)) xor (layer0_outputs(9932)));
    outputs(2670) <= not(layer0_outputs(5118));
    outputs(2671) <= not((layer0_outputs(34)) xor (layer0_outputs(9611)));
    outputs(2672) <= layer0_outputs(43);
    outputs(2673) <= not(layer0_outputs(5538)) or (layer0_outputs(1617));
    outputs(2674) <= layer0_outputs(9849);
    outputs(2675) <= not(layer0_outputs(2376)) or (layer0_outputs(7275));
    outputs(2676) <= not((layer0_outputs(3846)) xor (layer0_outputs(1580)));
    outputs(2677) <= not(layer0_outputs(4850));
    outputs(2678) <= (layer0_outputs(7975)) and (layer0_outputs(1124));
    outputs(2679) <= not((layer0_outputs(2801)) xor (layer0_outputs(10452)));
    outputs(2680) <= layer0_outputs(6462);
    outputs(2681) <= (layer0_outputs(10805)) or (layer0_outputs(7916));
    outputs(2682) <= not(layer0_outputs(8625));
    outputs(2683) <= layer0_outputs(9680);
    outputs(2684) <= layer0_outputs(1332);
    outputs(2685) <= (layer0_outputs(5871)) xor (layer0_outputs(4255));
    outputs(2686) <= not(layer0_outputs(11878));
    outputs(2687) <= not(layer0_outputs(7426)) or (layer0_outputs(9340));
    outputs(2688) <= not((layer0_outputs(6524)) or (layer0_outputs(7403)));
    outputs(2689) <= not((layer0_outputs(11003)) xor (layer0_outputs(5012)));
    outputs(2690) <= (layer0_outputs(8046)) or (layer0_outputs(12762));
    outputs(2691) <= not(layer0_outputs(2314));
    outputs(2692) <= layer0_outputs(7910);
    outputs(2693) <= not(layer0_outputs(9438));
    outputs(2694) <= layer0_outputs(3268);
    outputs(2695) <= '1';
    outputs(2696) <= not(layer0_outputs(6999));
    outputs(2697) <= not((layer0_outputs(9733)) xor (layer0_outputs(8056)));
    outputs(2698) <= not(layer0_outputs(8692));
    outputs(2699) <= not((layer0_outputs(7363)) or (layer0_outputs(12770)));
    outputs(2700) <= layer0_outputs(822);
    outputs(2701) <= not(layer0_outputs(10015));
    outputs(2702) <= layer0_outputs(9648);
    outputs(2703) <= layer0_outputs(30);
    outputs(2704) <= not(layer0_outputs(1203));
    outputs(2705) <= not(layer0_outputs(8953));
    outputs(2706) <= layer0_outputs(7671);
    outputs(2707) <= (layer0_outputs(8001)) or (layer0_outputs(4711));
    outputs(2708) <= not(layer0_outputs(9156)) or (layer0_outputs(2616));
    outputs(2709) <= not(layer0_outputs(1246));
    outputs(2710) <= not(layer0_outputs(7395));
    outputs(2711) <= not(layer0_outputs(4675));
    outputs(2712) <= (layer0_outputs(7337)) xor (layer0_outputs(4488));
    outputs(2713) <= layer0_outputs(6917);
    outputs(2714) <= not((layer0_outputs(2568)) xor (layer0_outputs(5095)));
    outputs(2715) <= not(layer0_outputs(9037)) or (layer0_outputs(8918));
    outputs(2716) <= not((layer0_outputs(4542)) xor (layer0_outputs(1982)));
    outputs(2717) <= not((layer0_outputs(9550)) xor (layer0_outputs(7624)));
    outputs(2718) <= layer0_outputs(12327);
    outputs(2719) <= (layer0_outputs(261)) or (layer0_outputs(4038));
    outputs(2720) <= layer0_outputs(12785);
    outputs(2721) <= not(layer0_outputs(8533));
    outputs(2722) <= not(layer0_outputs(6905)) or (layer0_outputs(11530));
    outputs(2723) <= not(layer0_outputs(2402)) or (layer0_outputs(11493));
    outputs(2724) <= not(layer0_outputs(5743));
    outputs(2725) <= not(layer0_outputs(12194));
    outputs(2726) <= (layer0_outputs(7810)) xor (layer0_outputs(9348));
    outputs(2727) <= '1';
    outputs(2728) <= '1';
    outputs(2729) <= not((layer0_outputs(10023)) and (layer0_outputs(12698)));
    outputs(2730) <= not(layer0_outputs(3284)) or (layer0_outputs(2624));
    outputs(2731) <= not((layer0_outputs(9200)) or (layer0_outputs(8102)));
    outputs(2732) <= not((layer0_outputs(10313)) and (layer0_outputs(12722)));
    outputs(2733) <= not(layer0_outputs(8441)) or (layer0_outputs(5478));
    outputs(2734) <= not(layer0_outputs(5260));
    outputs(2735) <= not(layer0_outputs(3773)) or (layer0_outputs(8387));
    outputs(2736) <= (layer0_outputs(278)) and not (layer0_outputs(7272));
    outputs(2737) <= (layer0_outputs(9992)) xor (layer0_outputs(7749));
    outputs(2738) <= (layer0_outputs(1766)) and not (layer0_outputs(133));
    outputs(2739) <= not(layer0_outputs(4131));
    outputs(2740) <= not(layer0_outputs(9514)) or (layer0_outputs(5753));
    outputs(2741) <= layer0_outputs(10311);
    outputs(2742) <= '1';
    outputs(2743) <= layer0_outputs(4950);
    outputs(2744) <= layer0_outputs(11687);
    outputs(2745) <= not((layer0_outputs(863)) xor (layer0_outputs(3850)));
    outputs(2746) <= not(layer0_outputs(6759)) or (layer0_outputs(95));
    outputs(2747) <= (layer0_outputs(6504)) xor (layer0_outputs(8821));
    outputs(2748) <= not(layer0_outputs(2370));
    outputs(2749) <= layer0_outputs(5411);
    outputs(2750) <= not(layer0_outputs(5898)) or (layer0_outputs(11837));
    outputs(2751) <= (layer0_outputs(5005)) and (layer0_outputs(4879));
    outputs(2752) <= layer0_outputs(11157);
    outputs(2753) <= layer0_outputs(3138);
    outputs(2754) <= layer0_outputs(6612);
    outputs(2755) <= not(layer0_outputs(5639));
    outputs(2756) <= layer0_outputs(8293);
    outputs(2757) <= not(layer0_outputs(6318));
    outputs(2758) <= not(layer0_outputs(4478));
    outputs(2759) <= not(layer0_outputs(6997));
    outputs(2760) <= (layer0_outputs(8152)) xor (layer0_outputs(9968));
    outputs(2761) <= not((layer0_outputs(3645)) xor (layer0_outputs(10709)));
    outputs(2762) <= not((layer0_outputs(12748)) xor (layer0_outputs(2524)));
    outputs(2763) <= layer0_outputs(9421);
    outputs(2764) <= not((layer0_outputs(6952)) or (layer0_outputs(1741)));
    outputs(2765) <= layer0_outputs(9328);
    outputs(2766) <= not((layer0_outputs(12031)) or (layer0_outputs(2610)));
    outputs(2767) <= (layer0_outputs(5948)) and not (layer0_outputs(4389));
    outputs(2768) <= (layer0_outputs(6839)) xor (layer0_outputs(8808));
    outputs(2769) <= '1';
    outputs(2770) <= (layer0_outputs(202)) or (layer0_outputs(5459));
    outputs(2771) <= not(layer0_outputs(9621));
    outputs(2772) <= not(layer0_outputs(1480));
    outputs(2773) <= (layer0_outputs(3253)) or (layer0_outputs(11237));
    outputs(2774) <= not(layer0_outputs(2692)) or (layer0_outputs(7697));
    outputs(2775) <= (layer0_outputs(8150)) and (layer0_outputs(11961));
    outputs(2776) <= not((layer0_outputs(6285)) xor (layer0_outputs(6787)));
    outputs(2777) <= not(layer0_outputs(10411));
    outputs(2778) <= not(layer0_outputs(3833));
    outputs(2779) <= (layer0_outputs(1035)) xor (layer0_outputs(5741));
    outputs(2780) <= (layer0_outputs(6794)) xor (layer0_outputs(621));
    outputs(2781) <= layer0_outputs(8584);
    outputs(2782) <= layer0_outputs(525);
    outputs(2783) <= not(layer0_outputs(1250));
    outputs(2784) <= layer0_outputs(3018);
    outputs(2785) <= (layer0_outputs(4838)) xor (layer0_outputs(7200));
    outputs(2786) <= not(layer0_outputs(2463)) or (layer0_outputs(8756));
    outputs(2787) <= layer0_outputs(4901);
    outputs(2788) <= not((layer0_outputs(786)) xor (layer0_outputs(5800)));
    outputs(2789) <= not((layer0_outputs(1989)) and (layer0_outputs(951)));
    outputs(2790) <= (layer0_outputs(6731)) and not (layer0_outputs(1250));
    outputs(2791) <= not(layer0_outputs(1678));
    outputs(2792) <= not(layer0_outputs(8250));
    outputs(2793) <= (layer0_outputs(3814)) and not (layer0_outputs(5406));
    outputs(2794) <= (layer0_outputs(8212)) or (layer0_outputs(4513));
    outputs(2795) <= layer0_outputs(12400);
    outputs(2796) <= (layer0_outputs(11224)) and (layer0_outputs(11991));
    outputs(2797) <= not(layer0_outputs(11996));
    outputs(2798) <= layer0_outputs(10428);
    outputs(2799) <= not(layer0_outputs(6403)) or (layer0_outputs(9305));
    outputs(2800) <= not(layer0_outputs(4538));
    outputs(2801) <= not((layer0_outputs(1029)) xor (layer0_outputs(5781)));
    outputs(2802) <= layer0_outputs(3101);
    outputs(2803) <= not(layer0_outputs(4508));
    outputs(2804) <= not(layer0_outputs(2280));
    outputs(2805) <= (layer0_outputs(738)) xor (layer0_outputs(3963));
    outputs(2806) <= (layer0_outputs(5977)) and (layer0_outputs(6507));
    outputs(2807) <= layer0_outputs(1461);
    outputs(2808) <= (layer0_outputs(11983)) xor (layer0_outputs(12176));
    outputs(2809) <= layer0_outputs(12378);
    outputs(2810) <= layer0_outputs(1058);
    outputs(2811) <= not(layer0_outputs(8544));
    outputs(2812) <= layer0_outputs(9354);
    outputs(2813) <= layer0_outputs(12007);
    outputs(2814) <= (layer0_outputs(6274)) xor (layer0_outputs(8894));
    outputs(2815) <= not(layer0_outputs(2015));
    outputs(2816) <= (layer0_outputs(12014)) and not (layer0_outputs(3322));
    outputs(2817) <= layer0_outputs(6909);
    outputs(2818) <= (layer0_outputs(3243)) xor (layer0_outputs(10115));
    outputs(2819) <= not(layer0_outputs(7917));
    outputs(2820) <= layer0_outputs(2964);
    outputs(2821) <= not((layer0_outputs(6741)) xor (layer0_outputs(7997)));
    outputs(2822) <= (layer0_outputs(4242)) xor (layer0_outputs(10287));
    outputs(2823) <= layer0_outputs(682);
    outputs(2824) <= not(layer0_outputs(3685));
    outputs(2825) <= (layer0_outputs(8269)) or (layer0_outputs(711));
    outputs(2826) <= (layer0_outputs(4416)) xor (layer0_outputs(4609));
    outputs(2827) <= not(layer0_outputs(4548));
    outputs(2828) <= not((layer0_outputs(1496)) and (layer0_outputs(2423)));
    outputs(2829) <= layer0_outputs(5175);
    outputs(2830) <= (layer0_outputs(3287)) xor (layer0_outputs(10808));
    outputs(2831) <= not((layer0_outputs(7224)) xor (layer0_outputs(12540)));
    outputs(2832) <= not(layer0_outputs(10477));
    outputs(2833) <= not(layer0_outputs(8003));
    outputs(2834) <= (layer0_outputs(2916)) xor (layer0_outputs(8786));
    outputs(2835) <= not((layer0_outputs(1698)) and (layer0_outputs(12156)));
    outputs(2836) <= not((layer0_outputs(11610)) or (layer0_outputs(8974)));
    outputs(2837) <= not(layer0_outputs(2777)) or (layer0_outputs(4702));
    outputs(2838) <= (layer0_outputs(12600)) and (layer0_outputs(10200));
    outputs(2839) <= not(layer0_outputs(12279)) or (layer0_outputs(3573));
    outputs(2840) <= (layer0_outputs(3091)) xor (layer0_outputs(6032));
    outputs(2841) <= not((layer0_outputs(8916)) xor (layer0_outputs(10611)));
    outputs(2842) <= not(layer0_outputs(96));
    outputs(2843) <= not((layer0_outputs(6581)) xor (layer0_outputs(12731)));
    outputs(2844) <= layer0_outputs(9851);
    outputs(2845) <= not((layer0_outputs(12006)) xor (layer0_outputs(7568)));
    outputs(2846) <= not(layer0_outputs(9425));
    outputs(2847) <= not(layer0_outputs(10048));
    outputs(2848) <= (layer0_outputs(1825)) and not (layer0_outputs(6819));
    outputs(2849) <= not(layer0_outputs(8213));
    outputs(2850) <= not(layer0_outputs(2600));
    outputs(2851) <= not((layer0_outputs(11241)) xor (layer0_outputs(3417)));
    outputs(2852) <= layer0_outputs(4874);
    outputs(2853) <= not((layer0_outputs(7498)) xor (layer0_outputs(5497)));
    outputs(2854) <= (layer0_outputs(4546)) and not (layer0_outputs(6911));
    outputs(2855) <= not(layer0_outputs(3840));
    outputs(2856) <= not(layer0_outputs(11623)) or (layer0_outputs(2535));
    outputs(2857) <= not((layer0_outputs(9047)) and (layer0_outputs(6631)));
    outputs(2858) <= not((layer0_outputs(6137)) and (layer0_outputs(9973)));
    outputs(2859) <= '1';
    outputs(2860) <= (layer0_outputs(1056)) xor (layer0_outputs(6623));
    outputs(2861) <= not(layer0_outputs(6297));
    outputs(2862) <= not((layer0_outputs(603)) and (layer0_outputs(9084)));
    outputs(2863) <= (layer0_outputs(8344)) xor (layer0_outputs(10115));
    outputs(2864) <= (layer0_outputs(6870)) or (layer0_outputs(11411));
    outputs(2865) <= (layer0_outputs(7168)) xor (layer0_outputs(4944));
    outputs(2866) <= not((layer0_outputs(2126)) and (layer0_outputs(2726)));
    outputs(2867) <= '0';
    outputs(2868) <= not(layer0_outputs(9059));
    outputs(2869) <= layer0_outputs(11240);
    outputs(2870) <= (layer0_outputs(1973)) xor (layer0_outputs(5792));
    outputs(2871) <= not((layer0_outputs(7037)) xor (layer0_outputs(7273)));
    outputs(2872) <= (layer0_outputs(12736)) xor (layer0_outputs(6316));
    outputs(2873) <= layer0_outputs(8850);
    outputs(2874) <= not(layer0_outputs(3336)) or (layer0_outputs(5060));
    outputs(2875) <= (layer0_outputs(9885)) and not (layer0_outputs(2105));
    outputs(2876) <= not((layer0_outputs(3907)) or (layer0_outputs(3386)));
    outputs(2877) <= layer0_outputs(10248);
    outputs(2878) <= layer0_outputs(11137);
    outputs(2879) <= layer0_outputs(7152);
    outputs(2880) <= not(layer0_outputs(6755));
    outputs(2881) <= not(layer0_outputs(319)) or (layer0_outputs(11394));
    outputs(2882) <= not((layer0_outputs(2873)) xor (layer0_outputs(5912)));
    outputs(2883) <= not(layer0_outputs(5392)) or (layer0_outputs(9274));
    outputs(2884) <= layer0_outputs(9902);
    outputs(2885) <= not(layer0_outputs(3068));
    outputs(2886) <= layer0_outputs(2647);
    outputs(2887) <= (layer0_outputs(1750)) xor (layer0_outputs(2990));
    outputs(2888) <= not(layer0_outputs(5192));
    outputs(2889) <= not((layer0_outputs(9905)) xor (layer0_outputs(1950)));
    outputs(2890) <= (layer0_outputs(4235)) xor (layer0_outputs(2743));
    outputs(2891) <= not(layer0_outputs(10816));
    outputs(2892) <= not((layer0_outputs(9360)) and (layer0_outputs(4947)));
    outputs(2893) <= not(layer0_outputs(2697)) or (layer0_outputs(5738));
    outputs(2894) <= '1';
    outputs(2895) <= layer0_outputs(5492);
    outputs(2896) <= layer0_outputs(7180);
    outputs(2897) <= layer0_outputs(8477);
    outputs(2898) <= not(layer0_outputs(9972)) or (layer0_outputs(11542));
    outputs(2899) <= not((layer0_outputs(1756)) or (layer0_outputs(1434)));
    outputs(2900) <= not((layer0_outputs(6404)) and (layer0_outputs(9869)));
    outputs(2901) <= not(layer0_outputs(1115));
    outputs(2902) <= not(layer0_outputs(7011));
    outputs(2903) <= layer0_outputs(9910);
    outputs(2904) <= layer0_outputs(4069);
    outputs(2905) <= not(layer0_outputs(1684)) or (layer0_outputs(2832));
    outputs(2906) <= '1';
    outputs(2907) <= not((layer0_outputs(11286)) xor (layer0_outputs(2998)));
    outputs(2908) <= not(layer0_outputs(49)) or (layer0_outputs(1415));
    outputs(2909) <= layer0_outputs(628);
    outputs(2910) <= layer0_outputs(11369);
    outputs(2911) <= not(layer0_outputs(2682));
    outputs(2912) <= (layer0_outputs(4159)) xor (layer0_outputs(10371));
    outputs(2913) <= not((layer0_outputs(7836)) xor (layer0_outputs(6497)));
    outputs(2914) <= not(layer0_outputs(4440)) or (layer0_outputs(2705));
    outputs(2915) <= not((layer0_outputs(11463)) xor (layer0_outputs(988)));
    outputs(2916) <= (layer0_outputs(8997)) and (layer0_outputs(4563));
    outputs(2917) <= not((layer0_outputs(1603)) or (layer0_outputs(7334)));
    outputs(2918) <= not((layer0_outputs(11518)) xor (layer0_outputs(8051)));
    outputs(2919) <= not((layer0_outputs(2380)) xor (layer0_outputs(10950)));
    outputs(2920) <= not(layer0_outputs(2843));
    outputs(2921) <= not(layer0_outputs(11833));
    outputs(2922) <= not((layer0_outputs(7966)) xor (layer0_outputs(3666)));
    outputs(2923) <= not((layer0_outputs(2481)) and (layer0_outputs(6252)));
    outputs(2924) <= not(layer0_outputs(3665));
    outputs(2925) <= not(layer0_outputs(6082)) or (layer0_outputs(6879));
    outputs(2926) <= not(layer0_outputs(2334));
    outputs(2927) <= (layer0_outputs(8559)) xor (layer0_outputs(12131));
    outputs(2928) <= not((layer0_outputs(10121)) and (layer0_outputs(11519)));
    outputs(2929) <= layer0_outputs(2368);
    outputs(2930) <= not(layer0_outputs(9380)) or (layer0_outputs(10753));
    outputs(2931) <= (layer0_outputs(12013)) xor (layer0_outputs(1196));
    outputs(2932) <= layer0_outputs(6139);
    outputs(2933) <= (layer0_outputs(5271)) xor (layer0_outputs(5316));
    outputs(2934) <= layer0_outputs(2906);
    outputs(2935) <= layer0_outputs(2748);
    outputs(2936) <= not(layer0_outputs(5968));
    outputs(2937) <= not((layer0_outputs(2109)) xor (layer0_outputs(4899)));
    outputs(2938) <= not((layer0_outputs(1123)) and (layer0_outputs(9390)));
    outputs(2939) <= (layer0_outputs(2591)) and not (layer0_outputs(12435));
    outputs(2940) <= not(layer0_outputs(11600));
    outputs(2941) <= not((layer0_outputs(10247)) and (layer0_outputs(11587)));
    outputs(2942) <= not((layer0_outputs(3794)) xor (layer0_outputs(7573)));
    outputs(2943) <= not(layer0_outputs(9578));
    outputs(2944) <= not(layer0_outputs(4938));
    outputs(2945) <= (layer0_outputs(3484)) xor (layer0_outputs(3621));
    outputs(2946) <= not((layer0_outputs(7199)) xor (layer0_outputs(7926)));
    outputs(2947) <= not((layer0_outputs(336)) xor (layer0_outputs(12406)));
    outputs(2948) <= not(layer0_outputs(5211));
    outputs(2949) <= layer0_outputs(11234);
    outputs(2950) <= (layer0_outputs(1833)) xor (layer0_outputs(5068));
    outputs(2951) <= layer0_outputs(6435);
    outputs(2952) <= not((layer0_outputs(1762)) or (layer0_outputs(8168)));
    outputs(2953) <= not((layer0_outputs(2899)) or (layer0_outputs(6984)));
    outputs(2954) <= not((layer0_outputs(6578)) xor (layer0_outputs(4422)));
    outputs(2955) <= not(layer0_outputs(8320));
    outputs(2956) <= not((layer0_outputs(12440)) or (layer0_outputs(724)));
    outputs(2957) <= layer0_outputs(9159);
    outputs(2958) <= layer0_outputs(1495);
    outputs(2959) <= (layer0_outputs(6280)) or (layer0_outputs(2650));
    outputs(2960) <= (layer0_outputs(4409)) xor (layer0_outputs(1292));
    outputs(2961) <= not(layer0_outputs(9698)) or (layer0_outputs(8950));
    outputs(2962) <= layer0_outputs(10086);
    outputs(2963) <= not((layer0_outputs(1479)) and (layer0_outputs(4776)));
    outputs(2964) <= layer0_outputs(6067);
    outputs(2965) <= not(layer0_outputs(9687));
    outputs(2966) <= not((layer0_outputs(9615)) and (layer0_outputs(1826)));
    outputs(2967) <= not(layer0_outputs(3815));
    outputs(2968) <= layer0_outputs(998);
    outputs(2969) <= not((layer0_outputs(8530)) xor (layer0_outputs(6648)));
    outputs(2970) <= not((layer0_outputs(10803)) xor (layer0_outputs(249)));
    outputs(2971) <= not((layer0_outputs(11416)) xor (layer0_outputs(11685)));
    outputs(2972) <= (layer0_outputs(7110)) and (layer0_outputs(9613));
    outputs(2973) <= not(layer0_outputs(11003)) or (layer0_outputs(10715));
    outputs(2974) <= not((layer0_outputs(11636)) xor (layer0_outputs(12075)));
    outputs(2975) <= not((layer0_outputs(7897)) xor (layer0_outputs(9820)));
    outputs(2976) <= layer0_outputs(6511);
    outputs(2977) <= (layer0_outputs(1912)) or (layer0_outputs(1653));
    outputs(2978) <= not(layer0_outputs(2622));
    outputs(2979) <= not(layer0_outputs(4294)) or (layer0_outputs(1467));
    outputs(2980) <= layer0_outputs(12377);
    outputs(2981) <= layer0_outputs(11650);
    outputs(2982) <= (layer0_outputs(6467)) or (layer0_outputs(10108));
    outputs(2983) <= (layer0_outputs(10454)) and not (layer0_outputs(1465));
    outputs(2984) <= not((layer0_outputs(2500)) or (layer0_outputs(5519)));
    outputs(2985) <= (layer0_outputs(2654)) xor (layer0_outputs(8799));
    outputs(2986) <= (layer0_outputs(1981)) and not (layer0_outputs(1254));
    outputs(2987) <= not((layer0_outputs(3554)) xor (layer0_outputs(9034)));
    outputs(2988) <= layer0_outputs(12166);
    outputs(2989) <= (layer0_outputs(3625)) and not (layer0_outputs(11125));
    outputs(2990) <= (layer0_outputs(9574)) and not (layer0_outputs(4804));
    outputs(2991) <= '1';
    outputs(2992) <= not((layer0_outputs(42)) and (layer0_outputs(10365)));
    outputs(2993) <= not(layer0_outputs(12027)) or (layer0_outputs(9708));
    outputs(2994) <= not((layer0_outputs(4639)) xor (layer0_outputs(11738)));
    outputs(2995) <= not(layer0_outputs(1655));
    outputs(2996) <= not((layer0_outputs(6542)) xor (layer0_outputs(11021)));
    outputs(2997) <= not((layer0_outputs(4331)) xor (layer0_outputs(8899)));
    outputs(2998) <= layer0_outputs(5201);
    outputs(2999) <= not(layer0_outputs(12665));
    outputs(3000) <= not(layer0_outputs(11845));
    outputs(3001) <= layer0_outputs(5958);
    outputs(3002) <= layer0_outputs(10614);
    outputs(3003) <= layer0_outputs(7430);
    outputs(3004) <= not(layer0_outputs(10682));
    outputs(3005) <= layer0_outputs(11163);
    outputs(3006) <= not(layer0_outputs(8096));
    outputs(3007) <= not(layer0_outputs(428)) or (layer0_outputs(2363));
    outputs(3008) <= layer0_outputs(9196);
    outputs(3009) <= not(layer0_outputs(4412));
    outputs(3010) <= not(layer0_outputs(11161)) or (layer0_outputs(10148));
    outputs(3011) <= not(layer0_outputs(12770));
    outputs(3012) <= not(layer0_outputs(10992)) or (layer0_outputs(8754));
    outputs(3013) <= (layer0_outputs(10985)) or (layer0_outputs(9886));
    outputs(3014) <= not((layer0_outputs(1510)) xor (layer0_outputs(8832)));
    outputs(3015) <= not(layer0_outputs(2794));
    outputs(3016) <= not((layer0_outputs(5033)) xor (layer0_outputs(10644)));
    outputs(3017) <= (layer0_outputs(2441)) and (layer0_outputs(6037));
    outputs(3018) <= (layer0_outputs(4962)) xor (layer0_outputs(1703));
    outputs(3019) <= (layer0_outputs(6904)) and (layer0_outputs(1775));
    outputs(3020) <= not(layer0_outputs(11469));
    outputs(3021) <= (layer0_outputs(8208)) and not (layer0_outputs(1516));
    outputs(3022) <= layer0_outputs(5133);
    outputs(3023) <= not(layer0_outputs(4758));
    outputs(3024) <= not(layer0_outputs(11176));
    outputs(3025) <= layer0_outputs(1900);
    outputs(3026) <= not(layer0_outputs(7397));
    outputs(3027) <= not(layer0_outputs(11667));
    outputs(3028) <= not((layer0_outputs(7348)) and (layer0_outputs(1587)));
    outputs(3029) <= layer0_outputs(9092);
    outputs(3030) <= layer0_outputs(5129);
    outputs(3031) <= not(layer0_outputs(9298)) or (layer0_outputs(5240));
    outputs(3032) <= layer0_outputs(5181);
    outputs(3033) <= layer0_outputs(9126);
    outputs(3034) <= not((layer0_outputs(1095)) or (layer0_outputs(9346)));
    outputs(3035) <= (layer0_outputs(3537)) or (layer0_outputs(10818));
    outputs(3036) <= not((layer0_outputs(9266)) xor (layer0_outputs(8342)));
    outputs(3037) <= not(layer0_outputs(7363));
    outputs(3038) <= layer0_outputs(11212);
    outputs(3039) <= layer0_outputs(728);
    outputs(3040) <= not(layer0_outputs(10271)) or (layer0_outputs(6676));
    outputs(3041) <= not(layer0_outputs(5798));
    outputs(3042) <= not((layer0_outputs(10677)) xor (layer0_outputs(5324)));
    outputs(3043) <= not(layer0_outputs(9379));
    outputs(3044) <= not((layer0_outputs(6449)) xor (layer0_outputs(1550)));
    outputs(3045) <= (layer0_outputs(2104)) xor (layer0_outputs(9639));
    outputs(3046) <= layer0_outputs(7107);
    outputs(3047) <= not(layer0_outputs(2845)) or (layer0_outputs(12410));
    outputs(3048) <= not(layer0_outputs(4042)) or (layer0_outputs(4514));
    outputs(3049) <= (layer0_outputs(10838)) and (layer0_outputs(8197));
    outputs(3050) <= not(layer0_outputs(7088));
    outputs(3051) <= not((layer0_outputs(8701)) and (layer0_outputs(9596)));
    outputs(3052) <= not(layer0_outputs(6088)) or (layer0_outputs(2893));
    outputs(3053) <= not(layer0_outputs(92));
    outputs(3054) <= not(layer0_outputs(4997));
    outputs(3055) <= not(layer0_outputs(3977));
    outputs(3056) <= not(layer0_outputs(10773));
    outputs(3057) <= not(layer0_outputs(1246)) or (layer0_outputs(825));
    outputs(3058) <= not(layer0_outputs(2084)) or (layer0_outputs(5149));
    outputs(3059) <= layer0_outputs(11016);
    outputs(3060) <= (layer0_outputs(767)) xor (layer0_outputs(11536));
    outputs(3061) <= layer0_outputs(5338);
    outputs(3062) <= not(layer0_outputs(7771)) or (layer0_outputs(8904));
    outputs(3063) <= (layer0_outputs(2)) and (layer0_outputs(12058));
    outputs(3064) <= (layer0_outputs(8358)) xor (layer0_outputs(10641));
    outputs(3065) <= layer0_outputs(8622);
    outputs(3066) <= not((layer0_outputs(7107)) xor (layer0_outputs(9121)));
    outputs(3067) <= layer0_outputs(8309);
    outputs(3068) <= (layer0_outputs(12652)) or (layer0_outputs(6882));
    outputs(3069) <= not((layer0_outputs(9832)) xor (layer0_outputs(2156)));
    outputs(3070) <= (layer0_outputs(1952)) xor (layer0_outputs(855));
    outputs(3071) <= layer0_outputs(8062);
    outputs(3072) <= not((layer0_outputs(12447)) xor (layer0_outputs(1540)));
    outputs(3073) <= not(layer0_outputs(5710));
    outputs(3074) <= (layer0_outputs(11905)) or (layer0_outputs(6171));
    outputs(3075) <= (layer0_outputs(7089)) xor (layer0_outputs(7323));
    outputs(3076) <= not((layer0_outputs(11263)) and (layer0_outputs(7227)));
    outputs(3077) <= layer0_outputs(1964);
    outputs(3078) <= not((layer0_outputs(5222)) xor (layer0_outputs(8066)));
    outputs(3079) <= not(layer0_outputs(516));
    outputs(3080) <= not(layer0_outputs(1913)) or (layer0_outputs(10536));
    outputs(3081) <= not((layer0_outputs(4424)) and (layer0_outputs(9772)));
    outputs(3082) <= not(layer0_outputs(12398));
    outputs(3083) <= not((layer0_outputs(4322)) xor (layer0_outputs(7753)));
    outputs(3084) <= (layer0_outputs(1824)) and (layer0_outputs(3393));
    outputs(3085) <= not((layer0_outputs(3542)) xor (layer0_outputs(2576)));
    outputs(3086) <= layer0_outputs(2397);
    outputs(3087) <= (layer0_outputs(2734)) and not (layer0_outputs(2451));
    outputs(3088) <= not(layer0_outputs(1846)) or (layer0_outputs(12585));
    outputs(3089) <= layer0_outputs(1824);
    outputs(3090) <= (layer0_outputs(2144)) and not (layer0_outputs(3036));
    outputs(3091) <= not(layer0_outputs(1577));
    outputs(3092) <= not(layer0_outputs(3598));
    outputs(3093) <= (layer0_outputs(9730)) and not (layer0_outputs(10025));
    outputs(3094) <= not(layer0_outputs(10529));
    outputs(3095) <= not(layer0_outputs(2150)) or (layer0_outputs(6761));
    outputs(3096) <= layer0_outputs(392);
    outputs(3097) <= not((layer0_outputs(1796)) xor (layer0_outputs(5274)));
    outputs(3098) <= (layer0_outputs(5138)) and not (layer0_outputs(5363));
    outputs(3099) <= (layer0_outputs(10169)) xor (layer0_outputs(2548));
    outputs(3100) <= not((layer0_outputs(2963)) or (layer0_outputs(8574)));
    outputs(3101) <= (layer0_outputs(3360)) xor (layer0_outputs(10904));
    outputs(3102) <= (layer0_outputs(3775)) xor (layer0_outputs(4343));
    outputs(3103) <= layer0_outputs(10006);
    outputs(3104) <= not(layer0_outputs(388));
    outputs(3105) <= not(layer0_outputs(10709)) or (layer0_outputs(6977));
    outputs(3106) <= not(layer0_outputs(10493));
    outputs(3107) <= not((layer0_outputs(12410)) and (layer0_outputs(7756)));
    outputs(3108) <= not(layer0_outputs(7310));
    outputs(3109) <= (layer0_outputs(4948)) xor (layer0_outputs(1948));
    outputs(3110) <= layer0_outputs(5692);
    outputs(3111) <= not((layer0_outputs(9422)) or (layer0_outputs(4535)));
    outputs(3112) <= not(layer0_outputs(4517)) or (layer0_outputs(11190));
    outputs(3113) <= not((layer0_outputs(2372)) and (layer0_outputs(12140)));
    outputs(3114) <= not(layer0_outputs(9132));
    outputs(3115) <= not(layer0_outputs(6169));
    outputs(3116) <= not((layer0_outputs(2000)) and (layer0_outputs(7945)));
    outputs(3117) <= not((layer0_outputs(2938)) or (layer0_outputs(2978)));
    outputs(3118) <= (layer0_outputs(1625)) and not (layer0_outputs(12489));
    outputs(3119) <= (layer0_outputs(4908)) xor (layer0_outputs(1277));
    outputs(3120) <= layer0_outputs(9253);
    outputs(3121) <= (layer0_outputs(1551)) xor (layer0_outputs(3749));
    outputs(3122) <= (layer0_outputs(12409)) xor (layer0_outputs(5532));
    outputs(3123) <= (layer0_outputs(1742)) and not (layer0_outputs(2230));
    outputs(3124) <= not(layer0_outputs(6651));
    outputs(3125) <= not(layer0_outputs(1973));
    outputs(3126) <= (layer0_outputs(2276)) or (layer0_outputs(10136));
    outputs(3127) <= not(layer0_outputs(9572)) or (layer0_outputs(4316));
    outputs(3128) <= (layer0_outputs(12129)) xor (layer0_outputs(6441));
    outputs(3129) <= not((layer0_outputs(6784)) and (layer0_outputs(11362)));
    outputs(3130) <= not(layer0_outputs(3540));
    outputs(3131) <= not(layer0_outputs(8148));
    outputs(3132) <= layer0_outputs(3454);
    outputs(3133) <= not(layer0_outputs(9533));
    outputs(3134) <= not((layer0_outputs(2527)) and (layer0_outputs(6655)));
    outputs(3135) <= not(layer0_outputs(5415));
    outputs(3136) <= not((layer0_outputs(9391)) xor (layer0_outputs(6227)));
    outputs(3137) <= layer0_outputs(10209);
    outputs(3138) <= layer0_outputs(6586);
    outputs(3139) <= not(layer0_outputs(3884)) or (layer0_outputs(3758));
    outputs(3140) <= (layer0_outputs(12349)) xor (layer0_outputs(8401));
    outputs(3141) <= not((layer0_outputs(9306)) xor (layer0_outputs(9606)));
    outputs(3142) <= not((layer0_outputs(4328)) xor (layer0_outputs(2036)));
    outputs(3143) <= not(layer0_outputs(3961));
    outputs(3144) <= (layer0_outputs(4068)) and not (layer0_outputs(6191));
    outputs(3145) <= not((layer0_outputs(11014)) and (layer0_outputs(10139)));
    outputs(3146) <= not(layer0_outputs(5610));
    outputs(3147) <= (layer0_outputs(676)) and not (layer0_outputs(6685));
    outputs(3148) <= (layer0_outputs(8220)) xor (layer0_outputs(3954));
    outputs(3149) <= not((layer0_outputs(559)) or (layer0_outputs(7601)));
    outputs(3150) <= (layer0_outputs(3570)) and not (layer0_outputs(3605));
    outputs(3151) <= not(layer0_outputs(8367));
    outputs(3152) <= (layer0_outputs(10527)) xor (layer0_outputs(2944));
    outputs(3153) <= not(layer0_outputs(11720));
    outputs(3154) <= not(layer0_outputs(3377));
    outputs(3155) <= not((layer0_outputs(5889)) xor (layer0_outputs(8176)));
    outputs(3156) <= layer0_outputs(4779);
    outputs(3157) <= not(layer0_outputs(1922));
    outputs(3158) <= not(layer0_outputs(10011));
    outputs(3159) <= (layer0_outputs(10624)) xor (layer0_outputs(10234));
    outputs(3160) <= not((layer0_outputs(3954)) xor (layer0_outputs(4403)));
    outputs(3161) <= (layer0_outputs(7526)) xor (layer0_outputs(9901));
    outputs(3162) <= layer0_outputs(628);
    outputs(3163) <= not((layer0_outputs(10355)) and (layer0_outputs(8517)));
    outputs(3164) <= (layer0_outputs(11335)) and (layer0_outputs(10860));
    outputs(3165) <= layer0_outputs(9273);
    outputs(3166) <= layer0_outputs(7252);
    outputs(3167) <= not((layer0_outputs(11741)) xor (layer0_outputs(2154)));
    outputs(3168) <= (layer0_outputs(4987)) xor (layer0_outputs(486));
    outputs(3169) <= not(layer0_outputs(8903));
    outputs(3170) <= not(layer0_outputs(5568));
    outputs(3171) <= not((layer0_outputs(9893)) xor (layer0_outputs(2343)));
    outputs(3172) <= layer0_outputs(3363);
    outputs(3173) <= not(layer0_outputs(11147));
    outputs(3174) <= (layer0_outputs(9966)) and not (layer0_outputs(11489));
    outputs(3175) <= layer0_outputs(7080);
    outputs(3176) <= not(layer0_outputs(3025));
    outputs(3177) <= not(layer0_outputs(11792));
    outputs(3178) <= not((layer0_outputs(863)) xor (layer0_outputs(9401)));
    outputs(3179) <= not(layer0_outputs(8488));
    outputs(3180) <= not(layer0_outputs(2122));
    outputs(3181) <= layer0_outputs(270);
    outputs(3182) <= (layer0_outputs(9474)) and not (layer0_outputs(3989));
    outputs(3183) <= not(layer0_outputs(361));
    outputs(3184) <= not(layer0_outputs(3624)) or (layer0_outputs(2558));
    outputs(3185) <= (layer0_outputs(1849)) and not (layer0_outputs(3516));
    outputs(3186) <= (layer0_outputs(6678)) and not (layer0_outputs(4718));
    outputs(3187) <= not(layer0_outputs(4132));
    outputs(3188) <= not(layer0_outputs(12431));
    outputs(3189) <= not(layer0_outputs(3208));
    outputs(3190) <= layer0_outputs(11229);
    outputs(3191) <= not(layer0_outputs(12197));
    outputs(3192) <= (layer0_outputs(5896)) xor (layer0_outputs(2364));
    outputs(3193) <= not(layer0_outputs(6279));
    outputs(3194) <= not(layer0_outputs(5135));
    outputs(3195) <= '1';
    outputs(3196) <= not((layer0_outputs(3767)) xor (layer0_outputs(7607)));
    outputs(3197) <= not(layer0_outputs(12269));
    outputs(3198) <= not(layer0_outputs(8320));
    outputs(3199) <= (layer0_outputs(1724)) xor (layer0_outputs(4439));
    outputs(3200) <= layer0_outputs(11886);
    outputs(3201) <= (layer0_outputs(4332)) or (layer0_outputs(10596));
    outputs(3202) <= (layer0_outputs(48)) and not (layer0_outputs(7447));
    outputs(3203) <= not((layer0_outputs(5162)) xor (layer0_outputs(6129)));
    outputs(3204) <= not(layer0_outputs(4469));
    outputs(3205) <= not((layer0_outputs(11411)) xor (layer0_outputs(2347)));
    outputs(3206) <= not((layer0_outputs(5788)) and (layer0_outputs(11384)));
    outputs(3207) <= not(layer0_outputs(7725)) or (layer0_outputs(2107));
    outputs(3208) <= not((layer0_outputs(9543)) and (layer0_outputs(4688)));
    outputs(3209) <= layer0_outputs(4795);
    outputs(3210) <= not(layer0_outputs(11709));
    outputs(3211) <= not((layer0_outputs(10485)) xor (layer0_outputs(11547)));
    outputs(3212) <= layer0_outputs(11750);
    outputs(3213) <= (layer0_outputs(12559)) and not (layer0_outputs(6124));
    outputs(3214) <= layer0_outputs(12789);
    outputs(3215) <= not((layer0_outputs(9478)) and (layer0_outputs(3820)));
    outputs(3216) <= (layer0_outputs(5938)) xor (layer0_outputs(310));
    outputs(3217) <= (layer0_outputs(5572)) or (layer0_outputs(8375));
    outputs(3218) <= not(layer0_outputs(11661));
    outputs(3219) <= (layer0_outputs(8669)) and (layer0_outputs(6254));
    outputs(3220) <= not((layer0_outputs(7611)) xor (layer0_outputs(12704)));
    outputs(3221) <= (layer0_outputs(11517)) xor (layer0_outputs(9831));
    outputs(3222) <= (layer0_outputs(52)) xor (layer0_outputs(10573));
    outputs(3223) <= not(layer0_outputs(1151));
    outputs(3224) <= not(layer0_outputs(11489));
    outputs(3225) <= (layer0_outputs(10892)) xor (layer0_outputs(10869));
    outputs(3226) <= '1';
    outputs(3227) <= not((layer0_outputs(3532)) and (layer0_outputs(6767)));
    outputs(3228) <= not((layer0_outputs(6843)) xor (layer0_outputs(7203)));
    outputs(3229) <= (layer0_outputs(3031)) and not (layer0_outputs(6849));
    outputs(3230) <= not((layer0_outputs(12162)) xor (layer0_outputs(8307)));
    outputs(3231) <= not(layer0_outputs(1249)) or (layer0_outputs(1389));
    outputs(3232) <= not(layer0_outputs(2040)) or (layer0_outputs(4676));
    outputs(3233) <= (layer0_outputs(199)) and (layer0_outputs(1522));
    outputs(3234) <= (layer0_outputs(12786)) and (layer0_outputs(9765));
    outputs(3235) <= not((layer0_outputs(6055)) and (layer0_outputs(5332)));
    outputs(3236) <= layer0_outputs(12666);
    outputs(3237) <= not(layer0_outputs(3769));
    outputs(3238) <= not(layer0_outputs(2462));
    outputs(3239) <= (layer0_outputs(5559)) xor (layer0_outputs(12556));
    outputs(3240) <= not(layer0_outputs(3913));
    outputs(3241) <= not(layer0_outputs(10865));
    outputs(3242) <= layer0_outputs(2331);
    outputs(3243) <= not((layer0_outputs(5414)) xor (layer0_outputs(3965)));
    outputs(3244) <= (layer0_outputs(12582)) xor (layer0_outputs(10395));
    outputs(3245) <= layer0_outputs(11135);
    outputs(3246) <= not(layer0_outputs(5777));
    outputs(3247) <= (layer0_outputs(6675)) or (layer0_outputs(7902));
    outputs(3248) <= not((layer0_outputs(4242)) xor (layer0_outputs(9114)));
    outputs(3249) <= layer0_outputs(10511);
    outputs(3250) <= not(layer0_outputs(12551)) or (layer0_outputs(10430));
    outputs(3251) <= not((layer0_outputs(1096)) or (layer0_outputs(2803)));
    outputs(3252) <= not((layer0_outputs(3558)) and (layer0_outputs(907)));
    outputs(3253) <= (layer0_outputs(5161)) and not (layer0_outputs(10946));
    outputs(3254) <= layer0_outputs(6304);
    outputs(3255) <= not(layer0_outputs(11706));
    outputs(3256) <= not(layer0_outputs(483)) or (layer0_outputs(9612));
    outputs(3257) <= not(layer0_outputs(4791));
    outputs(3258) <= layer0_outputs(12083);
    outputs(3259) <= layer0_outputs(1008);
    outputs(3260) <= not((layer0_outputs(6159)) xor (layer0_outputs(3779)));
    outputs(3261) <= (layer0_outputs(11108)) or (layer0_outputs(366));
    outputs(3262) <= layer0_outputs(5956);
    outputs(3263) <= (layer0_outputs(7117)) or (layer0_outputs(1704));
    outputs(3264) <= (layer0_outputs(8725)) xor (layer0_outputs(520));
    outputs(3265) <= layer0_outputs(9999);
    outputs(3266) <= layer0_outputs(8899);
    outputs(3267) <= (layer0_outputs(5556)) and (layer0_outputs(9824));
    outputs(3268) <= not((layer0_outputs(5704)) xor (layer0_outputs(4402)));
    outputs(3269) <= layer0_outputs(3019);
    outputs(3270) <= not(layer0_outputs(3479));
    outputs(3271) <= (layer0_outputs(3029)) xor (layer0_outputs(5661));
    outputs(3272) <= (layer0_outputs(11521)) or (layer0_outputs(11364));
    outputs(3273) <= not((layer0_outputs(7643)) xor (layer0_outputs(2004)));
    outputs(3274) <= not(layer0_outputs(2297));
    outputs(3275) <= not((layer0_outputs(10528)) xor (layer0_outputs(2688)));
    outputs(3276) <= not(layer0_outputs(12419)) or (layer0_outputs(9531));
    outputs(3277) <= not(layer0_outputs(5003));
    outputs(3278) <= not((layer0_outputs(8564)) or (layer0_outputs(9427)));
    outputs(3279) <= (layer0_outputs(12346)) and not (layer0_outputs(12300));
    outputs(3280) <= not((layer0_outputs(7439)) xor (layer0_outputs(4282)));
    outputs(3281) <= (layer0_outputs(5633)) and not (layer0_outputs(12011));
    outputs(3282) <= layer0_outputs(3364);
    outputs(3283) <= not(layer0_outputs(9435));
    outputs(3284) <= not(layer0_outputs(6743));
    outputs(3285) <= not(layer0_outputs(58)) or (layer0_outputs(1670));
    outputs(3286) <= not((layer0_outputs(5563)) xor (layer0_outputs(6926)));
    outputs(3287) <= not(layer0_outputs(7997));
    outputs(3288) <= not(layer0_outputs(2653));
    outputs(3289) <= not((layer0_outputs(11308)) xor (layer0_outputs(9467)));
    outputs(3290) <= not(layer0_outputs(11719));
    outputs(3291) <= not((layer0_outputs(9369)) xor (layer0_outputs(11711)));
    outputs(3292) <= (layer0_outputs(2241)) xor (layer0_outputs(10472));
    outputs(3293) <= not(layer0_outputs(1229));
    outputs(3294) <= not((layer0_outputs(7505)) or (layer0_outputs(479)));
    outputs(3295) <= not(layer0_outputs(4281)) or (layer0_outputs(4939));
    outputs(3296) <= (layer0_outputs(9608)) and not (layer0_outputs(12466));
    outputs(3297) <= not(layer0_outputs(10034));
    outputs(3298) <= (layer0_outputs(2535)) or (layer0_outputs(5058));
    outputs(3299) <= layer0_outputs(11119);
    outputs(3300) <= layer0_outputs(2732);
    outputs(3301) <= (layer0_outputs(9816)) and not (layer0_outputs(7412));
    outputs(3302) <= not(layer0_outputs(3680));
    outputs(3303) <= not((layer0_outputs(8656)) and (layer0_outputs(11221)));
    outputs(3304) <= (layer0_outputs(7172)) and not (layer0_outputs(11267));
    outputs(3305) <= not(layer0_outputs(11023)) or (layer0_outputs(11473));
    outputs(3306) <= not(layer0_outputs(3669)) or (layer0_outputs(7504));
    outputs(3307) <= not(layer0_outputs(9523));
    outputs(3308) <= not((layer0_outputs(10298)) xor (layer0_outputs(475)));
    outputs(3309) <= not(layer0_outputs(4494));
    outputs(3310) <= layer0_outputs(3404);
    outputs(3311) <= not((layer0_outputs(7000)) xor (layer0_outputs(1481)));
    outputs(3312) <= not((layer0_outputs(7213)) xor (layer0_outputs(1895)));
    outputs(3313) <= not(layer0_outputs(3276));
    outputs(3314) <= not(layer0_outputs(4671));
    outputs(3315) <= not(layer0_outputs(1674));
    outputs(3316) <= not((layer0_outputs(3324)) and (layer0_outputs(6297)));
    outputs(3317) <= layer0_outputs(1121);
    outputs(3318) <= not(layer0_outputs(8181)) or (layer0_outputs(8800));
    outputs(3319) <= (layer0_outputs(755)) and not (layer0_outputs(8815));
    outputs(3320) <= not((layer0_outputs(934)) and (layer0_outputs(6206)));
    outputs(3321) <= not((layer0_outputs(81)) or (layer0_outputs(8519)));
    outputs(3322) <= (layer0_outputs(4263)) xor (layer0_outputs(9394));
    outputs(3323) <= not((layer0_outputs(10631)) xor (layer0_outputs(2234)));
    outputs(3324) <= not((layer0_outputs(5241)) xor (layer0_outputs(9315)));
    outputs(3325) <= (layer0_outputs(2422)) and not (layer0_outputs(7673));
    outputs(3326) <= (layer0_outputs(7006)) xor (layer0_outputs(7010));
    outputs(3327) <= layer0_outputs(1851);
    outputs(3328) <= (layer0_outputs(8199)) or (layer0_outputs(5292));
    outputs(3329) <= (layer0_outputs(389)) and (layer0_outputs(5794));
    outputs(3330) <= layer0_outputs(9206);
    outputs(3331) <= not(layer0_outputs(8044));
    outputs(3332) <= not(layer0_outputs(11736)) or (layer0_outputs(3946));
    outputs(3333) <= layer0_outputs(9458);
    outputs(3334) <= (layer0_outputs(4400)) xor (layer0_outputs(6838));
    outputs(3335) <= not(layer0_outputs(9026));
    outputs(3336) <= not(layer0_outputs(5709));
    outputs(3337) <= not((layer0_outputs(5128)) xor (layer0_outputs(6499)));
    outputs(3338) <= not(layer0_outputs(6651));
    outputs(3339) <= not(layer0_outputs(12233));
    outputs(3340) <= not((layer0_outputs(4223)) xor (layer0_outputs(7972)));
    outputs(3341) <= not(layer0_outputs(709));
    outputs(3342) <= (layer0_outputs(8526)) or (layer0_outputs(605));
    outputs(3343) <= (layer0_outputs(1654)) and not (layer0_outputs(10542));
    outputs(3344) <= (layer0_outputs(121)) or (layer0_outputs(10800));
    outputs(3345) <= (layer0_outputs(3983)) xor (layer0_outputs(5439));
    outputs(3346) <= layer0_outputs(877);
    outputs(3347) <= not(layer0_outputs(10469)) or (layer0_outputs(5261));
    outputs(3348) <= layer0_outputs(6517);
    outputs(3349) <= layer0_outputs(12690);
    outputs(3350) <= layer0_outputs(8379);
    outputs(3351) <= not(layer0_outputs(7583)) or (layer0_outputs(1893));
    outputs(3352) <= not((layer0_outputs(4892)) xor (layer0_outputs(9934)));
    outputs(3353) <= layer0_outputs(468);
    outputs(3354) <= layer0_outputs(4736);
    outputs(3355) <= not(layer0_outputs(4940));
    outputs(3356) <= not(layer0_outputs(10693)) or (layer0_outputs(10760));
    outputs(3357) <= not(layer0_outputs(312)) or (layer0_outputs(11713));
    outputs(3358) <= not((layer0_outputs(1218)) and (layer0_outputs(10992)));
    outputs(3359) <= (layer0_outputs(3011)) and not (layer0_outputs(4986));
    outputs(3360) <= not(layer0_outputs(12656)) or (layer0_outputs(9820));
    outputs(3361) <= not(layer0_outputs(9529));
    outputs(3362) <= (layer0_outputs(9884)) or (layer0_outputs(2852));
    outputs(3363) <= not(layer0_outputs(4850));
    outputs(3364) <= not((layer0_outputs(3706)) xor (layer0_outputs(3576)));
    outputs(3365) <= layer0_outputs(126);
    outputs(3366) <= (layer0_outputs(5096)) or (layer0_outputs(11251));
    outputs(3367) <= (layer0_outputs(3790)) xor (layer0_outputs(3723));
    outputs(3368) <= (layer0_outputs(1233)) and (layer0_outputs(697));
    outputs(3369) <= (layer0_outputs(6957)) and not (layer0_outputs(8812));
    outputs(3370) <= not(layer0_outputs(1280));
    outputs(3371) <= (layer0_outputs(814)) xor (layer0_outputs(4238));
    outputs(3372) <= not(layer0_outputs(8157)) or (layer0_outputs(12455));
    outputs(3373) <= not(layer0_outputs(11833));
    outputs(3374) <= not((layer0_outputs(7041)) xor (layer0_outputs(2344)));
    outputs(3375) <= not(layer0_outputs(8615));
    outputs(3376) <= layer0_outputs(9587);
    outputs(3377) <= not((layer0_outputs(10750)) and (layer0_outputs(10204)));
    outputs(3378) <= not(layer0_outputs(11911)) or (layer0_outputs(7660));
    outputs(3379) <= not(layer0_outputs(1662)) or (layer0_outputs(6721));
    outputs(3380) <= not((layer0_outputs(3186)) xor (layer0_outputs(6814)));
    outputs(3381) <= not(layer0_outputs(7582));
    outputs(3382) <= not(layer0_outputs(1239)) or (layer0_outputs(2875));
    outputs(3383) <= not(layer0_outputs(7846));
    outputs(3384) <= not((layer0_outputs(1108)) xor (layer0_outputs(824)));
    outputs(3385) <= layer0_outputs(7232);
    outputs(3386) <= (layer0_outputs(5201)) or (layer0_outputs(2789));
    outputs(3387) <= '1';
    outputs(3388) <= not((layer0_outputs(7618)) xor (layer0_outputs(12106)));
    outputs(3389) <= not(layer0_outputs(7648));
    outputs(3390) <= not(layer0_outputs(7289)) or (layer0_outputs(12421));
    outputs(3391) <= (layer0_outputs(8879)) or (layer0_outputs(7076));
    outputs(3392) <= (layer0_outputs(12037)) or (layer0_outputs(12087));
    outputs(3393) <= (layer0_outputs(1967)) or (layer0_outputs(9241));
    outputs(3394) <= not(layer0_outputs(6058));
    outputs(3395) <= not(layer0_outputs(11798));
    outputs(3396) <= (layer0_outputs(2598)) and (layer0_outputs(1647));
    outputs(3397) <= not(layer0_outputs(3228));
    outputs(3398) <= not(layer0_outputs(10910));
    outputs(3399) <= (layer0_outputs(1324)) and (layer0_outputs(13));
    outputs(3400) <= not((layer0_outputs(9581)) or (layer0_outputs(3316)));
    outputs(3401) <= (layer0_outputs(6073)) xor (layer0_outputs(9684));
    outputs(3402) <= not(layer0_outputs(789)) or (layer0_outputs(7794));
    outputs(3403) <= layer0_outputs(1527);
    outputs(3404) <= not((layer0_outputs(9655)) and (layer0_outputs(511)));
    outputs(3405) <= not((layer0_outputs(2087)) or (layer0_outputs(1631)));
    outputs(3406) <= (layer0_outputs(1103)) xor (layer0_outputs(10412));
    outputs(3407) <= not(layer0_outputs(1979));
    outputs(3408) <= not((layer0_outputs(6818)) and (layer0_outputs(6557)));
    outputs(3409) <= (layer0_outputs(7864)) xor (layer0_outputs(12313));
    outputs(3410) <= layer0_outputs(9470);
    outputs(3411) <= not((layer0_outputs(3127)) xor (layer0_outputs(2263)));
    outputs(3412) <= not((layer0_outputs(2234)) xor (layer0_outputs(9248)));
    outputs(3413) <= not((layer0_outputs(10683)) or (layer0_outputs(2822)));
    outputs(3414) <= not(layer0_outputs(8410));
    outputs(3415) <= (layer0_outputs(6580)) and (layer0_outputs(7623));
    outputs(3416) <= not((layer0_outputs(3073)) xor (layer0_outputs(12128)));
    outputs(3417) <= not((layer0_outputs(10594)) and (layer0_outputs(6480)));
    outputs(3418) <= not((layer0_outputs(1739)) xor (layer0_outputs(6790)));
    outputs(3419) <= (layer0_outputs(5496)) xor (layer0_outputs(5876));
    outputs(3420) <= not(layer0_outputs(4579)) or (layer0_outputs(8141));
    outputs(3421) <= (layer0_outputs(7561)) and not (layer0_outputs(10303));
    outputs(3422) <= not((layer0_outputs(6355)) xor (layer0_outputs(10476)));
    outputs(3423) <= layer0_outputs(1002);
    outputs(3424) <= not(layer0_outputs(8582));
    outputs(3425) <= not(layer0_outputs(2958)) or (layer0_outputs(4773));
    outputs(3426) <= not(layer0_outputs(6406));
    outputs(3427) <= (layer0_outputs(7297)) xor (layer0_outputs(1669));
    outputs(3428) <= not(layer0_outputs(6152));
    outputs(3429) <= (layer0_outputs(4532)) xor (layer0_outputs(6617));
    outputs(3430) <= not(layer0_outputs(4771));
    outputs(3431) <= not((layer0_outputs(3908)) xor (layer0_outputs(3503)));
    outputs(3432) <= not(layer0_outputs(4698));
    outputs(3433) <= (layer0_outputs(5240)) or (layer0_outputs(5828));
    outputs(3434) <= not((layer0_outputs(1772)) xor (layer0_outputs(12081)));
    outputs(3435) <= (layer0_outputs(10369)) xor (layer0_outputs(9579));
    outputs(3436) <= (layer0_outputs(3831)) xor (layer0_outputs(10008));
    outputs(3437) <= not((layer0_outputs(10713)) xor (layer0_outputs(5978)));
    outputs(3438) <= layer0_outputs(5478);
    outputs(3439) <= not(layer0_outputs(9446));
    outputs(3440) <= not(layer0_outputs(6019));
    outputs(3441) <= not((layer0_outputs(6805)) xor (layer0_outputs(3433)));
    outputs(3442) <= (layer0_outputs(8639)) xor (layer0_outputs(5814));
    outputs(3443) <= (layer0_outputs(2592)) xor (layer0_outputs(3514));
    outputs(3444) <= not((layer0_outputs(2208)) or (layer0_outputs(8180)));
    outputs(3445) <= (layer0_outputs(806)) and not (layer0_outputs(8293));
    outputs(3446) <= layer0_outputs(4283);
    outputs(3447) <= not(layer0_outputs(12398));
    outputs(3448) <= layer0_outputs(3347);
    outputs(3449) <= layer0_outputs(607);
    outputs(3450) <= not(layer0_outputs(4220));
    outputs(3451) <= (layer0_outputs(7995)) xor (layer0_outputs(10757));
    outputs(3452) <= (layer0_outputs(962)) xor (layer0_outputs(11988));
    outputs(3453) <= not((layer0_outputs(7592)) xor (layer0_outputs(5834)));
    outputs(3454) <= (layer0_outputs(3099)) or (layer0_outputs(1763));
    outputs(3455) <= not(layer0_outputs(11028)) or (layer0_outputs(686));
    outputs(3456) <= layer0_outputs(9303);
    outputs(3457) <= layer0_outputs(5692);
    outputs(3458) <= (layer0_outputs(5150)) xor (layer0_outputs(2769));
    outputs(3459) <= layer0_outputs(6133);
    outputs(3460) <= layer0_outputs(8091);
    outputs(3461) <= layer0_outputs(12565);
    outputs(3462) <= not(layer0_outputs(5082));
    outputs(3463) <= (layer0_outputs(9213)) and (layer0_outputs(12612));
    outputs(3464) <= not(layer0_outputs(2064)) or (layer0_outputs(316));
    outputs(3465) <= not(layer0_outputs(11467));
    outputs(3466) <= layer0_outputs(10191);
    outputs(3467) <= not(layer0_outputs(1879));
    outputs(3468) <= layer0_outputs(9207);
    outputs(3469) <= layer0_outputs(11780);
    outputs(3470) <= (layer0_outputs(10701)) xor (layer0_outputs(4315));
    outputs(3471) <= (layer0_outputs(443)) and not (layer0_outputs(4218));
    outputs(3472) <= not((layer0_outputs(9517)) and (layer0_outputs(12064)));
    outputs(3473) <= not((layer0_outputs(1229)) xor (layer0_outputs(419)));
    outputs(3474) <= not((layer0_outputs(7045)) xor (layer0_outputs(1828)));
    outputs(3475) <= (layer0_outputs(3266)) and not (layer0_outputs(515));
    outputs(3476) <= layer0_outputs(8171);
    outputs(3477) <= not(layer0_outputs(12124));
    outputs(3478) <= layer0_outputs(614);
    outputs(3479) <= not(layer0_outputs(4344)) or (layer0_outputs(6142));
    outputs(3480) <= not((layer0_outputs(5159)) or (layer0_outputs(6157)));
    outputs(3481) <= (layer0_outputs(2090)) xor (layer0_outputs(7027));
    outputs(3482) <= layer0_outputs(10439);
    outputs(3483) <= not(layer0_outputs(4426));
    outputs(3484) <= not(layer0_outputs(7510)) or (layer0_outputs(10811));
    outputs(3485) <= layer0_outputs(8748);
    outputs(3486) <= layer0_outputs(3958);
    outputs(3487) <= layer0_outputs(5190);
    outputs(3488) <= not((layer0_outputs(11868)) and (layer0_outputs(9101)));
    outputs(3489) <= not((layer0_outputs(11330)) xor (layer0_outputs(1049)));
    outputs(3490) <= not(layer0_outputs(12284));
    outputs(3491) <= not(layer0_outputs(5992));
    outputs(3492) <= not((layer0_outputs(1286)) xor (layer0_outputs(10950)));
    outputs(3493) <= not(layer0_outputs(6577));
    outputs(3494) <= not((layer0_outputs(1878)) xor (layer0_outputs(12650)));
    outputs(3495) <= not(layer0_outputs(10784));
    outputs(3496) <= not((layer0_outputs(305)) or (layer0_outputs(9867)));
    outputs(3497) <= (layer0_outputs(6676)) xor (layer0_outputs(11497));
    outputs(3498) <= not(layer0_outputs(10151)) or (layer0_outputs(1858));
    outputs(3499) <= not(layer0_outputs(3791)) or (layer0_outputs(12282));
    outputs(3500) <= not((layer0_outputs(5120)) and (layer0_outputs(5631)));
    outputs(3501) <= (layer0_outputs(4000)) xor (layer0_outputs(9067));
    outputs(3502) <= not(layer0_outputs(5362)) or (layer0_outputs(2242));
    outputs(3503) <= not(layer0_outputs(5391));
    outputs(3504) <= not((layer0_outputs(9580)) xor (layer0_outputs(11999)));
    outputs(3505) <= layer0_outputs(11624);
    outputs(3506) <= (layer0_outputs(1128)) or (layer0_outputs(8000));
    outputs(3507) <= layer0_outputs(10404);
    outputs(3508) <= not((layer0_outputs(5970)) xor (layer0_outputs(8133)));
    outputs(3509) <= layer0_outputs(12127);
    outputs(3510) <= not(layer0_outputs(10172));
    outputs(3511) <= (layer0_outputs(11951)) and (layer0_outputs(11758));
    outputs(3512) <= not(layer0_outputs(12420)) or (layer0_outputs(6510));
    outputs(3513) <= layer0_outputs(7890);
    outputs(3514) <= not(layer0_outputs(2364));
    outputs(3515) <= not(layer0_outputs(7226)) or (layer0_outputs(85));
    outputs(3516) <= not((layer0_outputs(7062)) xor (layer0_outputs(10440)));
    outputs(3517) <= (layer0_outputs(8683)) and (layer0_outputs(2294));
    outputs(3518) <= (layer0_outputs(9843)) or (layer0_outputs(7546));
    outputs(3519) <= (layer0_outputs(1937)) xor (layer0_outputs(9));
    outputs(3520) <= (layer0_outputs(9562)) and not (layer0_outputs(2396));
    outputs(3521) <= not(layer0_outputs(1178));
    outputs(3522) <= layer0_outputs(3490);
    outputs(3523) <= layer0_outputs(8668);
    outputs(3524) <= (layer0_outputs(492)) xor (layer0_outputs(11599));
    outputs(3525) <= not((layer0_outputs(10343)) xor (layer0_outputs(10754)));
    outputs(3526) <= (layer0_outputs(2770)) and not (layer0_outputs(649));
    outputs(3527) <= not(layer0_outputs(6820));
    outputs(3528) <= not((layer0_outputs(1838)) xor (layer0_outputs(1037)));
    outputs(3529) <= (layer0_outputs(8542)) and not (layer0_outputs(2566));
    outputs(3530) <= not((layer0_outputs(7249)) and (layer0_outputs(4290)));
    outputs(3531) <= not((layer0_outputs(3417)) xor (layer0_outputs(3735)));
    outputs(3532) <= not((layer0_outputs(1346)) and (layer0_outputs(11676)));
    outputs(3533) <= not((layer0_outputs(5400)) and (layer0_outputs(2217)));
    outputs(3534) <= layer0_outputs(11881);
    outputs(3535) <= (layer0_outputs(884)) xor (layer0_outputs(4143));
    outputs(3536) <= not((layer0_outputs(4717)) and (layer0_outputs(8684)));
    outputs(3537) <= layer0_outputs(1337);
    outputs(3538) <= not((layer0_outputs(8693)) or (layer0_outputs(6636)));
    outputs(3539) <= not(layer0_outputs(2017));
    outputs(3540) <= not(layer0_outputs(10974));
    outputs(3541) <= layer0_outputs(3252);
    outputs(3542) <= not((layer0_outputs(11210)) xor (layer0_outputs(2335)));
    outputs(3543) <= not(layer0_outputs(12390));
    outputs(3544) <= not((layer0_outputs(5224)) and (layer0_outputs(6368)));
    outputs(3545) <= layer0_outputs(7312);
    outputs(3546) <= not(layer0_outputs(12655));
    outputs(3547) <= layer0_outputs(2974);
    outputs(3548) <= layer0_outputs(2833);
    outputs(3549) <= layer0_outputs(1982);
    outputs(3550) <= layer0_outputs(12450);
    outputs(3551) <= not((layer0_outputs(3260)) and (layer0_outputs(3703)));
    outputs(3552) <= not(layer0_outputs(12607)) or (layer0_outputs(10470));
    outputs(3553) <= not((layer0_outputs(3212)) xor (layer0_outputs(8955)));
    outputs(3554) <= (layer0_outputs(2227)) xor (layer0_outputs(5440));
    outputs(3555) <= layer0_outputs(4680);
    outputs(3556) <= not((layer0_outputs(8440)) and (layer0_outputs(1507)));
    outputs(3557) <= layer0_outputs(2223);
    outputs(3558) <= not(layer0_outputs(6427));
    outputs(3559) <= (layer0_outputs(6794)) xor (layer0_outputs(4971));
    outputs(3560) <= not(layer0_outputs(11637));
    outputs(3561) <= not((layer0_outputs(10446)) xor (layer0_outputs(2035)));
    outputs(3562) <= layer0_outputs(4822);
    outputs(3563) <= not((layer0_outputs(2931)) xor (layer0_outputs(10425)));
    outputs(3564) <= layer0_outputs(12321);
    outputs(3565) <= (layer0_outputs(5062)) xor (layer0_outputs(10945));
    outputs(3566) <= not(layer0_outputs(5529));
    outputs(3567) <= layer0_outputs(11590);
    outputs(3568) <= not((layer0_outputs(774)) and (layer0_outputs(12727)));
    outputs(3569) <= not((layer0_outputs(5910)) and (layer0_outputs(11566)));
    outputs(3570) <= not(layer0_outputs(4961));
    outputs(3571) <= layer0_outputs(8395);
    outputs(3572) <= layer0_outputs(3825);
    outputs(3573) <= layer0_outputs(9122);
    outputs(3574) <= not((layer0_outputs(312)) xor (layer0_outputs(4399)));
    outputs(3575) <= not(layer0_outputs(11383));
    outputs(3576) <= not(layer0_outputs(5032));
    outputs(3577) <= (layer0_outputs(11847)) xor (layer0_outputs(9760));
    outputs(3578) <= (layer0_outputs(11179)) xor (layer0_outputs(558));
    outputs(3579) <= (layer0_outputs(5486)) or (layer0_outputs(2116));
    outputs(3580) <= layer0_outputs(1889);
    outputs(3581) <= (layer0_outputs(6185)) and not (layer0_outputs(6485));
    outputs(3582) <= not(layer0_outputs(489));
    outputs(3583) <= not((layer0_outputs(8479)) or (layer0_outputs(8608)));
    outputs(3584) <= not(layer0_outputs(763)) or (layer0_outputs(8987));
    outputs(3585) <= (layer0_outputs(3471)) and not (layer0_outputs(1631));
    outputs(3586) <= not((layer0_outputs(8888)) or (layer0_outputs(400)));
    outputs(3587) <= not(layer0_outputs(8761));
    outputs(3588) <= not(layer0_outputs(1722));
    outputs(3589) <= not((layer0_outputs(8277)) xor (layer0_outputs(11507)));
    outputs(3590) <= not(layer0_outputs(7366));
    outputs(3591) <= not((layer0_outputs(1562)) xor (layer0_outputs(9640)));
    outputs(3592) <= (layer0_outputs(6878)) and not (layer0_outputs(11254));
    outputs(3593) <= not((layer0_outputs(7872)) xor (layer0_outputs(281)));
    outputs(3594) <= not((layer0_outputs(967)) and (layer0_outputs(10487)));
    outputs(3595) <= (layer0_outputs(11866)) and (layer0_outputs(5824));
    outputs(3596) <= not(layer0_outputs(2538)) or (layer0_outputs(5915));
    outputs(3597) <= not(layer0_outputs(7002)) or (layer0_outputs(6427));
    outputs(3598) <= layer0_outputs(11508);
    outputs(3599) <= not((layer0_outputs(7)) or (layer0_outputs(3303)));
    outputs(3600) <= (layer0_outputs(8319)) and not (layer0_outputs(5152));
    outputs(3601) <= not((layer0_outputs(12108)) xor (layer0_outputs(6942)));
    outputs(3602) <= (layer0_outputs(4179)) xor (layer0_outputs(11019));
    outputs(3603) <= not(layer0_outputs(2733)) or (layer0_outputs(11696));
    outputs(3604) <= (layer0_outputs(3809)) xor (layer0_outputs(9937));
    outputs(3605) <= not(layer0_outputs(6616));
    outputs(3606) <= layer0_outputs(11399);
    outputs(3607) <= not(layer0_outputs(3260));
    outputs(3608) <= not((layer0_outputs(4203)) and (layer0_outputs(5972)));
    outputs(3609) <= not((layer0_outputs(382)) and (layer0_outputs(8854)));
    outputs(3610) <= not(layer0_outputs(746));
    outputs(3611) <= layer0_outputs(8773);
    outputs(3612) <= not((layer0_outputs(2762)) xor (layer0_outputs(9863)));
    outputs(3613) <= (layer0_outputs(1322)) and not (layer0_outputs(4163));
    outputs(3614) <= (layer0_outputs(2457)) xor (layer0_outputs(11985));
    outputs(3615) <= not(layer0_outputs(9499));
    outputs(3616) <= layer0_outputs(2383);
    outputs(3617) <= not((layer0_outputs(1071)) xor (layer0_outputs(1538)));
    outputs(3618) <= layer0_outputs(10094);
    outputs(3619) <= not(layer0_outputs(8106));
    outputs(3620) <= not((layer0_outputs(11751)) and (layer0_outputs(8874)));
    outputs(3621) <= layer0_outputs(7728);
    outputs(3622) <= not((layer0_outputs(8908)) xor (layer0_outputs(2080)));
    outputs(3623) <= layer0_outputs(4895);
    outputs(3624) <= not(layer0_outputs(7410));
    outputs(3625) <= (layer0_outputs(982)) and not (layer0_outputs(12408));
    outputs(3626) <= not((layer0_outputs(7144)) xor (layer0_outputs(1348)));
    outputs(3627) <= (layer0_outputs(4461)) and not (layer0_outputs(7286));
    outputs(3628) <= not(layer0_outputs(10884)) or (layer0_outputs(7646));
    outputs(3629) <= not((layer0_outputs(2179)) xor (layer0_outputs(3830)));
    outputs(3630) <= layer0_outputs(7534);
    outputs(3631) <= layer0_outputs(672);
    outputs(3632) <= not((layer0_outputs(10401)) xor (layer0_outputs(1351)));
    outputs(3633) <= not(layer0_outputs(2649)) or (layer0_outputs(11432));
    outputs(3634) <= not(layer0_outputs(8671));
    outputs(3635) <= not(layer0_outputs(2017));
    outputs(3636) <= (layer0_outputs(6556)) and (layer0_outputs(427));
    outputs(3637) <= layer0_outputs(3592);
    outputs(3638) <= (layer0_outputs(5655)) or (layer0_outputs(12719));
    outputs(3639) <= layer0_outputs(7528);
    outputs(3640) <= not(layer0_outputs(7086)) or (layer0_outputs(1392));
    outputs(3641) <= not(layer0_outputs(12335)) or (layer0_outputs(9974));
    outputs(3642) <= not(layer0_outputs(10059));
    outputs(3643) <= not((layer0_outputs(10399)) and (layer0_outputs(11393)));
    outputs(3644) <= not((layer0_outputs(787)) xor (layer0_outputs(6599)));
    outputs(3645) <= not(layer0_outputs(3434));
    outputs(3646) <= not(layer0_outputs(4996));
    outputs(3647) <= (layer0_outputs(1086)) and not (layer0_outputs(10936));
    outputs(3648) <= not(layer0_outputs(11645));
    outputs(3649) <= layer0_outputs(9487);
    outputs(3650) <= layer0_outputs(6244);
    outputs(3651) <= not((layer0_outputs(2633)) xor (layer0_outputs(7270)));
    outputs(3652) <= not((layer0_outputs(6292)) xor (layer0_outputs(1866)));
    outputs(3653) <= (layer0_outputs(12361)) and not (layer0_outputs(6565));
    outputs(3654) <= not(layer0_outputs(3098)) or (layer0_outputs(5592));
    outputs(3655) <= not((layer0_outputs(4985)) and (layer0_outputs(1146)));
    outputs(3656) <= not(layer0_outputs(5121));
    outputs(3657) <= not(layer0_outputs(3433));
    outputs(3658) <= layer0_outputs(3910);
    outputs(3659) <= not(layer0_outputs(2867)) or (layer0_outputs(10377));
    outputs(3660) <= not(layer0_outputs(3576));
    outputs(3661) <= (layer0_outputs(6580)) and not (layer0_outputs(1947));
    outputs(3662) <= (layer0_outputs(6226)) and not (layer0_outputs(6407));
    outputs(3663) <= not((layer0_outputs(4345)) and (layer0_outputs(9231)));
    outputs(3664) <= (layer0_outputs(11742)) xor (layer0_outputs(2939));
    outputs(3665) <= not(layer0_outputs(2759));
    outputs(3666) <= not((layer0_outputs(6729)) xor (layer0_outputs(9482)));
    outputs(3667) <= (layer0_outputs(11269)) xor (layer0_outputs(10363));
    outputs(3668) <= layer0_outputs(3397);
    outputs(3669) <= layer0_outputs(9228);
    outputs(3670) <= not(layer0_outputs(12390));
    outputs(3671) <= (layer0_outputs(1129)) xor (layer0_outputs(3776));
    outputs(3672) <= (layer0_outputs(12761)) or (layer0_outputs(4014));
    outputs(3673) <= (layer0_outputs(8397)) xor (layer0_outputs(5652));
    outputs(3674) <= (layer0_outputs(1208)) xor (layer0_outputs(9331));
    outputs(3675) <= (layer0_outputs(2582)) or (layer0_outputs(12032));
    outputs(3676) <= not((layer0_outputs(7157)) and (layer0_outputs(10744)));
    outputs(3677) <= not(layer0_outputs(3021));
    outputs(3678) <= layer0_outputs(6933);
    outputs(3679) <= not((layer0_outputs(1042)) xor (layer0_outputs(12507)));
    outputs(3680) <= '1';
    outputs(3681) <= (layer0_outputs(6119)) and not (layer0_outputs(6579));
    outputs(3682) <= layer0_outputs(6736);
    outputs(3683) <= not(layer0_outputs(4561));
    outputs(3684) <= not(layer0_outputs(817));
    outputs(3685) <= layer0_outputs(8766);
    outputs(3686) <= not((layer0_outputs(11621)) xor (layer0_outputs(3705)));
    outputs(3687) <= layer0_outputs(12666);
    outputs(3688) <= not((layer0_outputs(8720)) xor (layer0_outputs(9173)));
    outputs(3689) <= (layer0_outputs(12044)) xor (layer0_outputs(3897));
    outputs(3690) <= not(layer0_outputs(8118));
    outputs(3691) <= layer0_outputs(10687);
    outputs(3692) <= not(layer0_outputs(11483));
    outputs(3693) <= layer0_outputs(5820);
    outputs(3694) <= not(layer0_outputs(5087)) or (layer0_outputs(4111));
    outputs(3695) <= (layer0_outputs(11247)) or (layer0_outputs(1675));
    outputs(3696) <= not(layer0_outputs(10216)) or (layer0_outputs(10098));
    outputs(3697) <= not((layer0_outputs(3782)) xor (layer0_outputs(6989)));
    outputs(3698) <= not(layer0_outputs(1272)) or (layer0_outputs(10165));
    outputs(3699) <= (layer0_outputs(8425)) and not (layer0_outputs(10464));
    outputs(3700) <= not((layer0_outputs(7655)) xor (layer0_outputs(9381)));
    outputs(3701) <= not((layer0_outputs(8133)) xor (layer0_outputs(6635)));
    outputs(3702) <= (layer0_outputs(9161)) xor (layer0_outputs(565));
    outputs(3703) <= (layer0_outputs(2037)) or (layer0_outputs(2554));
    outputs(3704) <= (layer0_outputs(2193)) xor (layer0_outputs(5255));
    outputs(3705) <= (layer0_outputs(4306)) xor (layer0_outputs(2951));
    outputs(3706) <= (layer0_outputs(2139)) xor (layer0_outputs(7075));
    outputs(3707) <= not(layer0_outputs(3832));
    outputs(3708) <= (layer0_outputs(1171)) xor (layer0_outputs(6866));
    outputs(3709) <= not(layer0_outputs(7603));
    outputs(3710) <= (layer0_outputs(7188)) and not (layer0_outputs(12695));
    outputs(3711) <= (layer0_outputs(2392)) and not (layer0_outputs(2597));
    outputs(3712) <= layer0_outputs(11227);
    outputs(3713) <= not(layer0_outputs(9870));
    outputs(3714) <= not((layer0_outputs(4388)) xor (layer0_outputs(1850)));
    outputs(3715) <= not(layer0_outputs(8080));
    outputs(3716) <= (layer0_outputs(5180)) xor (layer0_outputs(3723));
    outputs(3717) <= not(layer0_outputs(3223)) or (layer0_outputs(586));
    outputs(3718) <= layer0_outputs(4741);
    outputs(3719) <= layer0_outputs(11214);
    outputs(3720) <= layer0_outputs(1423);
    outputs(3721) <= (layer0_outputs(9784)) xor (layer0_outputs(8078));
    outputs(3722) <= not(layer0_outputs(9715)) or (layer0_outputs(3181));
    outputs(3723) <= (layer0_outputs(5816)) xor (layer0_outputs(9822));
    outputs(3724) <= (layer0_outputs(8935)) xor (layer0_outputs(3909));
    outputs(3725) <= not((layer0_outputs(106)) and (layer0_outputs(7289)));
    outputs(3726) <= layer0_outputs(4828);
    outputs(3727) <= not((layer0_outputs(2012)) or (layer0_outputs(5028)));
    outputs(3728) <= not(layer0_outputs(9817)) or (layer0_outputs(9650));
    outputs(3729) <= not(layer0_outputs(10848));
    outputs(3730) <= layer0_outputs(4935);
    outputs(3731) <= layer0_outputs(9591);
    outputs(3732) <= (layer0_outputs(12109)) xor (layer0_outputs(3729));
    outputs(3733) <= not(layer0_outputs(10734));
    outputs(3734) <= (layer0_outputs(4383)) xor (layer0_outputs(12252));
    outputs(3735) <= layer0_outputs(6728);
    outputs(3736) <= not(layer0_outputs(742));
    outputs(3737) <= not((layer0_outputs(3408)) xor (layer0_outputs(271)));
    outputs(3738) <= not(layer0_outputs(12663)) or (layer0_outputs(1420));
    outputs(3739) <= (layer0_outputs(8956)) or (layer0_outputs(11859));
    outputs(3740) <= (layer0_outputs(12705)) and not (layer0_outputs(7714));
    outputs(3741) <= not((layer0_outputs(2296)) xor (layer0_outputs(5484)));
    outputs(3742) <= layer0_outputs(3140);
    outputs(3743) <= not(layer0_outputs(5565)) or (layer0_outputs(5662));
    outputs(3744) <= (layer0_outputs(2904)) and (layer0_outputs(12142));
    outputs(3745) <= not((layer0_outputs(4684)) xor (layer0_outputs(8760)));
    outputs(3746) <= not((layer0_outputs(10568)) and (layer0_outputs(7613)));
    outputs(3747) <= not(layer0_outputs(795));
    outputs(3748) <= not((layer0_outputs(7563)) xor (layer0_outputs(7381)));
    outputs(3749) <= not(layer0_outputs(210));
    outputs(3750) <= layer0_outputs(6391);
    outputs(3751) <= layer0_outputs(12749);
    outputs(3752) <= not(layer0_outputs(1397));
    outputs(3753) <= (layer0_outputs(4751)) or (layer0_outputs(6658));
    outputs(3754) <= (layer0_outputs(1332)) and not (layer0_outputs(12002));
    outputs(3755) <= (layer0_outputs(2435)) xor (layer0_outputs(5142));
    outputs(3756) <= layer0_outputs(5401);
    outputs(3757) <= (layer0_outputs(7470)) xor (layer0_outputs(7141));
    outputs(3758) <= not(layer0_outputs(133));
    outputs(3759) <= not(layer0_outputs(11964));
    outputs(3760) <= not((layer0_outputs(6383)) xor (layer0_outputs(4407)));
    outputs(3761) <= (layer0_outputs(12697)) and not (layer0_outputs(9324));
    outputs(3762) <= (layer0_outputs(2138)) or (layer0_outputs(1048));
    outputs(3763) <= not(layer0_outputs(5057)) or (layer0_outputs(4503));
    outputs(3764) <= not(layer0_outputs(4490));
    outputs(3765) <= (layer0_outputs(12110)) and not (layer0_outputs(7952));
    outputs(3766) <= not(layer0_outputs(7936));
    outputs(3767) <= layer0_outputs(14);
    outputs(3768) <= not(layer0_outputs(6362));
    outputs(3769) <= layer0_outputs(7454);
    outputs(3770) <= not((layer0_outputs(11776)) xor (layer0_outputs(6109)));
    outputs(3771) <= not(layer0_outputs(7596));
    outputs(3772) <= not((layer0_outputs(9492)) or (layer0_outputs(10062)));
    outputs(3773) <= not((layer0_outputs(7882)) or (layer0_outputs(10044)));
    outputs(3774) <= not((layer0_outputs(371)) xor (layer0_outputs(9325)));
    outputs(3775) <= (layer0_outputs(12536)) xor (layer0_outputs(5231));
    outputs(3776) <= not((layer0_outputs(7739)) and (layer0_outputs(2432)));
    outputs(3777) <= (layer0_outputs(1207)) and (layer0_outputs(6312));
    outputs(3778) <= not(layer0_outputs(6712));
    outputs(3779) <= not((layer0_outputs(11729)) xor (layer0_outputs(2578)));
    outputs(3780) <= not(layer0_outputs(5046)) or (layer0_outputs(9632));
    outputs(3781) <= layer0_outputs(6748);
    outputs(3782) <= layer0_outputs(1193);
    outputs(3783) <= not(layer0_outputs(1204));
    outputs(3784) <= layer0_outputs(1402);
    outputs(3785) <= (layer0_outputs(9879)) or (layer0_outputs(2444));
    outputs(3786) <= not(layer0_outputs(11964));
    outputs(3787) <= (layer0_outputs(2172)) xor (layer0_outputs(1367));
    outputs(3788) <= not((layer0_outputs(2808)) xor (layer0_outputs(10900)));
    outputs(3789) <= not((layer0_outputs(7981)) and (layer0_outputs(6121)));
    outputs(3790) <= layer0_outputs(7227);
    outputs(3791) <= not(layer0_outputs(1729)) or (layer0_outputs(10449));
    outputs(3792) <= not(layer0_outputs(645)) or (layer0_outputs(2724));
    outputs(3793) <= not((layer0_outputs(1342)) xor (layer0_outputs(4180)));
    outputs(3794) <= not((layer0_outputs(11062)) and (layer0_outputs(11804)));
    outputs(3795) <= not((layer0_outputs(6066)) xor (layer0_outputs(4122)));
    outputs(3796) <= (layer0_outputs(7567)) xor (layer0_outputs(12544));
    outputs(3797) <= not(layer0_outputs(5520));
    outputs(3798) <= not(layer0_outputs(10723)) or (layer0_outputs(7342));
    outputs(3799) <= not((layer0_outputs(877)) and (layer0_outputs(7205)));
    outputs(3800) <= not(layer0_outputs(10277)) or (layer0_outputs(1855));
    outputs(3801) <= (layer0_outputs(12241)) and not (layer0_outputs(6038));
    outputs(3802) <= layer0_outputs(9080);
    outputs(3803) <= not(layer0_outputs(4641));
    outputs(3804) <= (layer0_outputs(6389)) xor (layer0_outputs(11416));
    outputs(3805) <= layer0_outputs(11018);
    outputs(3806) <= layer0_outputs(4386);
    outputs(3807) <= not(layer0_outputs(7486));
    outputs(3808) <= layer0_outputs(6391);
    outputs(3809) <= (layer0_outputs(6114)) xor (layer0_outputs(6779));
    outputs(3810) <= not(layer0_outputs(2815)) or (layer0_outputs(3912));
    outputs(3811) <= not(layer0_outputs(10194));
    outputs(3812) <= layer0_outputs(10534);
    outputs(3813) <= (layer0_outputs(9712)) and (layer0_outputs(5923));
    outputs(3814) <= (layer0_outputs(7496)) or (layer0_outputs(3946));
    outputs(3815) <= not(layer0_outputs(11681));
    outputs(3816) <= (layer0_outputs(10310)) xor (layer0_outputs(12568));
    outputs(3817) <= layer0_outputs(6788);
    outputs(3818) <= not(layer0_outputs(3130));
    outputs(3819) <= not(layer0_outputs(6816));
    outputs(3820) <= layer0_outputs(3564);
    outputs(3821) <= (layer0_outputs(5697)) or (layer0_outputs(7248));
    outputs(3822) <= (layer0_outputs(443)) and (layer0_outputs(11116));
    outputs(3823) <= layer0_outputs(2436);
    outputs(3824) <= not(layer0_outputs(11379));
    outputs(3825) <= not((layer0_outputs(986)) xor (layer0_outputs(346)));
    outputs(3826) <= not(layer0_outputs(7603));
    outputs(3827) <= not(layer0_outputs(1136));
    outputs(3828) <= not(layer0_outputs(754));
    outputs(3829) <= layer0_outputs(10400);
    outputs(3830) <= layer0_outputs(9859);
    outputs(3831) <= not(layer0_outputs(8692));
    outputs(3832) <= (layer0_outputs(5647)) and not (layer0_outputs(6137));
    outputs(3833) <= (layer0_outputs(3608)) and not (layer0_outputs(7190));
    outputs(3834) <= (layer0_outputs(5333)) xor (layer0_outputs(12595));
    outputs(3835) <= not((layer0_outputs(7681)) xor (layer0_outputs(5119)));
    outputs(3836) <= (layer0_outputs(1748)) xor (layer0_outputs(7382));
    outputs(3837) <= not(layer0_outputs(27));
    outputs(3838) <= (layer0_outputs(3411)) xor (layer0_outputs(1836));
    outputs(3839) <= (layer0_outputs(7961)) xor (layer0_outputs(2011));
    outputs(3840) <= layer0_outputs(10885);
    outputs(3841) <= not((layer0_outputs(2145)) and (layer0_outputs(8847)));
    outputs(3842) <= (layer0_outputs(11171)) and not (layer0_outputs(12042));
    outputs(3843) <= (layer0_outputs(1438)) xor (layer0_outputs(7999));
    outputs(3844) <= (layer0_outputs(9121)) xor (layer0_outputs(1820));
    outputs(3845) <= layer0_outputs(11812);
    outputs(3846) <= layer0_outputs(5937);
    outputs(3847) <= not(layer0_outputs(11348)) or (layer0_outputs(1911));
    outputs(3848) <= layer0_outputs(7776);
    outputs(3849) <= (layer0_outputs(11610)) or (layer0_outputs(243));
    outputs(3850) <= (layer0_outputs(8534)) xor (layer0_outputs(2751));
    outputs(3851) <= '1';
    outputs(3852) <= layer0_outputs(11151);
    outputs(3853) <= not((layer0_outputs(10348)) or (layer0_outputs(12431)));
    outputs(3854) <= layer0_outputs(11232);
    outputs(3855) <= not(layer0_outputs(4322));
    outputs(3856) <= not(layer0_outputs(3082)) or (layer0_outputs(11601));
    outputs(3857) <= layer0_outputs(2481);
    outputs(3858) <= not((layer0_outputs(4461)) or (layer0_outputs(1447)));
    outputs(3859) <= not((layer0_outputs(7914)) xor (layer0_outputs(8161)));
    outputs(3860) <= not((layer0_outputs(12797)) xor (layer0_outputs(3358)));
    outputs(3861) <= not(layer0_outputs(10373));
    outputs(3862) <= not(layer0_outputs(7643)) or (layer0_outputs(7408));
    outputs(3863) <= (layer0_outputs(7944)) and (layer0_outputs(7352));
    outputs(3864) <= not((layer0_outputs(11730)) and (layer0_outputs(3663)));
    outputs(3865) <= not(layer0_outputs(5041));
    outputs(3866) <= (layer0_outputs(4582)) and not (layer0_outputs(5975));
    outputs(3867) <= not((layer0_outputs(9584)) and (layer0_outputs(9475)));
    outputs(3868) <= not(layer0_outputs(7973));
    outputs(3869) <= not(layer0_outputs(3943)) or (layer0_outputs(4917));
    outputs(3870) <= not((layer0_outputs(7621)) or (layer0_outputs(8597)));
    outputs(3871) <= (layer0_outputs(4227)) xor (layer0_outputs(6813));
    outputs(3872) <= not(layer0_outputs(8329));
    outputs(3873) <= not(layer0_outputs(9235));
    outputs(3874) <= not(layer0_outputs(11979)) or (layer0_outputs(9776));
    outputs(3875) <= (layer0_outputs(6804)) xor (layer0_outputs(10186));
    outputs(3876) <= (layer0_outputs(6217)) xor (layer0_outputs(5313));
    outputs(3877) <= not(layer0_outputs(8637));
    outputs(3878) <= not(layer0_outputs(1034));
    outputs(3879) <= not(layer0_outputs(1487));
    outputs(3880) <= (layer0_outputs(4462)) and (layer0_outputs(9377));
    outputs(3881) <= layer0_outputs(7699);
    outputs(3882) <= not(layer0_outputs(4928));
    outputs(3883) <= not(layer0_outputs(3942)) or (layer0_outputs(606));
    outputs(3884) <= (layer0_outputs(8444)) xor (layer0_outputs(625));
    outputs(3885) <= not((layer0_outputs(8906)) xor (layer0_outputs(10756)));
    outputs(3886) <= not((layer0_outputs(8288)) xor (layer0_outputs(118)));
    outputs(3887) <= (layer0_outputs(2527)) xor (layer0_outputs(5802));
    outputs(3888) <= not(layer0_outputs(5078)) or (layer0_outputs(994));
    outputs(3889) <= not(layer0_outputs(3948));
    outputs(3890) <= not((layer0_outputs(6256)) or (layer0_outputs(8189)));
    outputs(3891) <= (layer0_outputs(38)) xor (layer0_outputs(9104));
    outputs(3892) <= (layer0_outputs(12502)) xor (layer0_outputs(1694));
    outputs(3893) <= not((layer0_outputs(4137)) xor (layer0_outputs(11877)));
    outputs(3894) <= not(layer0_outputs(2091));
    outputs(3895) <= not(layer0_outputs(10824)) or (layer0_outputs(7419));
    outputs(3896) <= not((layer0_outputs(5213)) xor (layer0_outputs(1361)));
    outputs(3897) <= layer0_outputs(6869);
    outputs(3898) <= not(layer0_outputs(6005));
    outputs(3899) <= not((layer0_outputs(7373)) xor (layer0_outputs(7779)));
    outputs(3900) <= (layer0_outputs(9573)) xor (layer0_outputs(9289));
    outputs(3901) <= layer0_outputs(6106);
    outputs(3902) <= layer0_outputs(4731);
    outputs(3903) <= layer0_outputs(9054);
    outputs(3904) <= '1';
    outputs(3905) <= layer0_outputs(220);
    outputs(3906) <= (layer0_outputs(3250)) xor (layer0_outputs(12726));
    outputs(3907) <= (layer0_outputs(7675)) and not (layer0_outputs(12754));
    outputs(3908) <= layer0_outputs(12641);
    outputs(3909) <= (layer0_outputs(7065)) xor (layer0_outputs(2183));
    outputs(3910) <= (layer0_outputs(2164)) xor (layer0_outputs(3900));
    outputs(3911) <= not(layer0_outputs(2389)) or (layer0_outputs(8406));
    outputs(3912) <= not(layer0_outputs(5491)) or (layer0_outputs(3406));
    outputs(3913) <= (layer0_outputs(11159)) or (layer0_outputs(1672));
    outputs(3914) <= layer0_outputs(720);
    outputs(3915) <= not(layer0_outputs(8066));
    outputs(3916) <= not(layer0_outputs(5370));
    outputs(3917) <= (layer0_outputs(11130)) xor (layer0_outputs(11114));
    outputs(3918) <= (layer0_outputs(9341)) or (layer0_outputs(899));
    outputs(3919) <= not((layer0_outputs(2470)) and (layer0_outputs(2699)));
    outputs(3920) <= (layer0_outputs(7765)) xor (layer0_outputs(1910));
    outputs(3921) <= (layer0_outputs(8429)) and not (layer0_outputs(5844));
    outputs(3922) <= (layer0_outputs(11313)) and not (layer0_outputs(8027));
    outputs(3923) <= (layer0_outputs(7390)) and (layer0_outputs(5630));
    outputs(3924) <= (layer0_outputs(9070)) and (layer0_outputs(3429));
    outputs(3925) <= not((layer0_outputs(12257)) xor (layer0_outputs(5260)));
    outputs(3926) <= (layer0_outputs(10233)) or (layer0_outputs(11875));
    outputs(3927) <= not((layer0_outputs(6222)) and (layer0_outputs(1759)));
    outputs(3928) <= (layer0_outputs(4672)) xor (layer0_outputs(3651));
    outputs(3929) <= not(layer0_outputs(3472));
    outputs(3930) <= not(layer0_outputs(7840));
    outputs(3931) <= not(layer0_outputs(235));
    outputs(3932) <= not(layer0_outputs(10978));
    outputs(3933) <= layer0_outputs(5436);
    outputs(3934) <= layer0_outputs(5595);
    outputs(3935) <= layer0_outputs(8592);
    outputs(3936) <= (layer0_outputs(10866)) and (layer0_outputs(1079));
    outputs(3937) <= not(layer0_outputs(12015));
    outputs(3938) <= (layer0_outputs(6474)) xor (layer0_outputs(12611));
    outputs(3939) <= (layer0_outputs(9247)) xor (layer0_outputs(7959));
    outputs(3940) <= (layer0_outputs(12441)) and not (layer0_outputs(8165));
    outputs(3941) <= (layer0_outputs(4544)) and not (layer0_outputs(8153));
    outputs(3942) <= layer0_outputs(10853);
    outputs(3943) <= (layer0_outputs(417)) or (layer0_outputs(10961));
    outputs(3944) <= not(layer0_outputs(10028));
    outputs(3945) <= layer0_outputs(11359);
    outputs(3946) <= layer0_outputs(2629);
    outputs(3947) <= (layer0_outputs(10326)) and not (layer0_outputs(8399));
    outputs(3948) <= not(layer0_outputs(6448)) or (layer0_outputs(4197));
    outputs(3949) <= (layer0_outputs(8085)) and not (layer0_outputs(1235));
    outputs(3950) <= layer0_outputs(4313);
    outputs(3951) <= (layer0_outputs(12552)) or (layer0_outputs(10825));
    outputs(3952) <= '1';
    outputs(3953) <= not(layer0_outputs(12682));
    outputs(3954) <= (layer0_outputs(5359)) and (layer0_outputs(6206));
    outputs(3955) <= not(layer0_outputs(1705));
    outputs(3956) <= (layer0_outputs(6423)) or (layer0_outputs(4264));
    outputs(3957) <= not((layer0_outputs(6143)) or (layer0_outputs(6342)));
    outputs(3958) <= (layer0_outputs(7368)) xor (layer0_outputs(2108));
    outputs(3959) <= (layer0_outputs(6859)) xor (layer0_outputs(5487));
    outputs(3960) <= not(layer0_outputs(5098));
    outputs(3961) <= not(layer0_outputs(7444));
    outputs(3962) <= (layer0_outputs(8603)) and not (layer0_outputs(4201));
    outputs(3963) <= not(layer0_outputs(9577));
    outputs(3964) <= not(layer0_outputs(10039)) or (layer0_outputs(9280));
    outputs(3965) <= (layer0_outputs(4799)) xor (layer0_outputs(4060));
    outputs(3966) <= not(layer0_outputs(4945));
    outputs(3967) <= layer0_outputs(10672);
    outputs(3968) <= not(layer0_outputs(2178));
    outputs(3969) <= not(layer0_outputs(5263));
    outputs(3970) <= layer0_outputs(1211);
    outputs(3971) <= not(layer0_outputs(9998));
    outputs(3972) <= (layer0_outputs(142)) and (layer0_outputs(6055));
    outputs(3973) <= not(layer0_outputs(11105));
    outputs(3974) <= not(layer0_outputs(3176));
    outputs(3975) <= (layer0_outputs(11109)) and (layer0_outputs(2864));
    outputs(3976) <= not((layer0_outputs(9472)) xor (layer0_outputs(2053)));
    outputs(3977) <= not((layer0_outputs(7038)) xor (layer0_outputs(10343)));
    outputs(3978) <= layer0_outputs(8043);
    outputs(3979) <= '1';
    outputs(3980) <= not((layer0_outputs(3116)) xor (layer0_outputs(4726)));
    outputs(3981) <= layer0_outputs(10585);
    outputs(3982) <= (layer0_outputs(11657)) or (layer0_outputs(10299));
    outputs(3983) <= (layer0_outputs(7678)) and not (layer0_outputs(7089));
    outputs(3984) <= not(layer0_outputs(8159)) or (layer0_outputs(9588));
    outputs(3985) <= (layer0_outputs(11869)) and not (layer0_outputs(5326));
    outputs(3986) <= not(layer0_outputs(10933)) or (layer0_outputs(8214));
    outputs(3987) <= not((layer0_outputs(11986)) or (layer0_outputs(12747)));
    outputs(3988) <= not(layer0_outputs(1500)) or (layer0_outputs(5578));
    outputs(3989) <= '1';
    outputs(3990) <= (layer0_outputs(9695)) xor (layer0_outputs(6754));
    outputs(3991) <= (layer0_outputs(2896)) and not (layer0_outputs(363));
    outputs(3992) <= layer0_outputs(832);
    outputs(3993) <= '1';
    outputs(3994) <= '1';
    outputs(3995) <= (layer0_outputs(944)) xor (layer0_outputs(12209));
    outputs(3996) <= layer0_outputs(7617);
    outputs(3997) <= not((layer0_outputs(10769)) or (layer0_outputs(8487)));
    outputs(3998) <= layer0_outputs(788);
    outputs(3999) <= not(layer0_outputs(1342));
    outputs(4000) <= (layer0_outputs(3350)) xor (layer0_outputs(2276));
    outputs(4001) <= not(layer0_outputs(1333));
    outputs(4002) <= (layer0_outputs(11343)) and not (layer0_outputs(7286));
    outputs(4003) <= (layer0_outputs(2525)) and (layer0_outputs(6458));
    outputs(4004) <= layer0_outputs(12516);
    outputs(4005) <= (layer0_outputs(1506)) xor (layer0_outputs(9853));
    outputs(4006) <= (layer0_outputs(8836)) and not (layer0_outputs(10321));
    outputs(4007) <= not(layer0_outputs(12192));
    outputs(4008) <= not(layer0_outputs(40)) or (layer0_outputs(7158));
    outputs(4009) <= (layer0_outputs(7806)) xor (layer0_outputs(6479));
    outputs(4010) <= not(layer0_outputs(5877));
    outputs(4011) <= (layer0_outputs(2750)) xor (layer0_outputs(2519));
    outputs(4012) <= (layer0_outputs(5214)) xor (layer0_outputs(3333));
    outputs(4013) <= '1';
    outputs(4014) <= layer0_outputs(4501);
    outputs(4015) <= layer0_outputs(9727);
    outputs(4016) <= (layer0_outputs(7540)) xor (layer0_outputs(4477));
    outputs(4017) <= layer0_outputs(10366);
    outputs(4018) <= not(layer0_outputs(12074));
    outputs(4019) <= not((layer0_outputs(2955)) xor (layer0_outputs(12574)));
    outputs(4020) <= (layer0_outputs(367)) and not (layer0_outputs(1212));
    outputs(4021) <= (layer0_outputs(2804)) xor (layer0_outputs(6488));
    outputs(4022) <= not((layer0_outputs(11882)) xor (layer0_outputs(12562)));
    outputs(4023) <= (layer0_outputs(6258)) and not (layer0_outputs(12434));
    outputs(4024) <= (layer0_outputs(7513)) or (layer0_outputs(3125));
    outputs(4025) <= (layer0_outputs(11372)) or (layer0_outputs(8435));
    outputs(4026) <= (layer0_outputs(6980)) xor (layer0_outputs(2034));
    outputs(4027) <= not(layer0_outputs(12733));
    outputs(4028) <= (layer0_outputs(4303)) or (layer0_outputs(2536));
    outputs(4029) <= (layer0_outputs(4250)) xor (layer0_outputs(6350));
    outputs(4030) <= not(layer0_outputs(11292)) or (layer0_outputs(2260));
    outputs(4031) <= not(layer0_outputs(7278));
    outputs(4032) <= not(layer0_outputs(3023));
    outputs(4033) <= (layer0_outputs(9336)) xor (layer0_outputs(560));
    outputs(4034) <= layer0_outputs(10345);
    outputs(4035) <= not((layer0_outputs(7292)) xor (layer0_outputs(8500)));
    outputs(4036) <= not(layer0_outputs(5311));
    outputs(4037) <= layer0_outputs(8690);
    outputs(4038) <= (layer0_outputs(12381)) or (layer0_outputs(5371));
    outputs(4039) <= layer0_outputs(9409);
    outputs(4040) <= (layer0_outputs(2027)) xor (layer0_outputs(8553));
    outputs(4041) <= not((layer0_outputs(8959)) xor (layer0_outputs(7707)));
    outputs(4042) <= (layer0_outputs(7624)) xor (layer0_outputs(7530));
    outputs(4043) <= not(layer0_outputs(10149));
    outputs(4044) <= (layer0_outputs(8175)) and not (layer0_outputs(6720));
    outputs(4045) <= not((layer0_outputs(5737)) xor (layer0_outputs(12043)));
    outputs(4046) <= not(layer0_outputs(7287));
    outputs(4047) <= (layer0_outputs(9439)) xor (layer0_outputs(3466));
    outputs(4048) <= (layer0_outputs(10230)) or (layer0_outputs(2644));
    outputs(4049) <= not(layer0_outputs(1919));
    outputs(4050) <= not((layer0_outputs(2447)) xor (layer0_outputs(3567)));
    outputs(4051) <= (layer0_outputs(4170)) xor (layer0_outputs(9569));
    outputs(4052) <= not(layer0_outputs(1419)) or (layer0_outputs(10135));
    outputs(4053) <= layer0_outputs(8384);
    outputs(4054) <= layer0_outputs(4372);
    outputs(4055) <= not(layer0_outputs(3878));
    outputs(4056) <= (layer0_outputs(8826)) xor (layer0_outputs(11165));
    outputs(4057) <= not(layer0_outputs(4573));
    outputs(4058) <= layer0_outputs(8614);
    outputs(4059) <= not(layer0_outputs(3372));
    outputs(4060) <= not(layer0_outputs(9221));
    outputs(4061) <= (layer0_outputs(11924)) and not (layer0_outputs(11361));
    outputs(4062) <= not(layer0_outputs(12723));
    outputs(4063) <= layer0_outputs(5779);
    outputs(4064) <= not(layer0_outputs(937));
    outputs(4065) <= not(layer0_outputs(10521)) or (layer0_outputs(2428));
    outputs(4066) <= (layer0_outputs(3897)) and (layer0_outputs(6670));
    outputs(4067) <= not(layer0_outputs(7051)) or (layer0_outputs(10956));
    outputs(4068) <= layer0_outputs(9871);
    outputs(4069) <= not(layer0_outputs(12296)) or (layer0_outputs(10695));
    outputs(4070) <= (layer0_outputs(7416)) xor (layer0_outputs(12077));
    outputs(4071) <= layer0_outputs(1135);
    outputs(4072) <= not(layer0_outputs(6898));
    outputs(4073) <= layer0_outputs(10394);
    outputs(4074) <= layer0_outputs(2283);
    outputs(4075) <= (layer0_outputs(12345)) and not (layer0_outputs(3044));
    outputs(4076) <= not((layer0_outputs(4834)) xor (layer0_outputs(3858)));
    outputs(4077) <= layer0_outputs(1647);
    outputs(4078) <= not(layer0_outputs(1998));
    outputs(4079) <= layer0_outputs(6990);
    outputs(4080) <= layer0_outputs(10205);
    outputs(4081) <= (layer0_outputs(10872)) and not (layer0_outputs(7645));
    outputs(4082) <= not(layer0_outputs(9362));
    outputs(4083) <= (layer0_outputs(8304)) or (layer0_outputs(440));
    outputs(4084) <= not(layer0_outputs(6363));
    outputs(4085) <= (layer0_outputs(1130)) or (layer0_outputs(1846));
    outputs(4086) <= layer0_outputs(7259);
    outputs(4087) <= not(layer0_outputs(9629)) or (layer0_outputs(11054));
    outputs(4088) <= (layer0_outputs(3099)) and not (layer0_outputs(3716));
    outputs(4089) <= not(layer0_outputs(5016));
    outputs(4090) <= not(layer0_outputs(7730)) or (layer0_outputs(9555));
    outputs(4091) <= not(layer0_outputs(7056));
    outputs(4092) <= layer0_outputs(7017);
    outputs(4093) <= not((layer0_outputs(215)) and (layer0_outputs(10082)));
    outputs(4094) <= layer0_outputs(6077);
    outputs(4095) <= layer0_outputs(21);
    outputs(4096) <= layer0_outputs(5389);
    outputs(4097) <= not((layer0_outputs(8859)) xor (layer0_outputs(5480)));
    outputs(4098) <= (layer0_outputs(9259)) and (layer0_outputs(11273));
    outputs(4099) <= layer0_outputs(8382);
    outputs(4100) <= not(layer0_outputs(12343)) or (layer0_outputs(10700));
    outputs(4101) <= layer0_outputs(8717);
    outputs(4102) <= not(layer0_outputs(9386));
    outputs(4103) <= not(layer0_outputs(10852));
    outputs(4104) <= not(layer0_outputs(10778));
    outputs(4105) <= (layer0_outputs(9714)) xor (layer0_outputs(7564));
    outputs(4106) <= not(layer0_outputs(7639));
    outputs(4107) <= not(layer0_outputs(5778));
    outputs(4108) <= not(layer0_outputs(12260));
    outputs(4109) <= (layer0_outputs(2547)) and not (layer0_outputs(2210));
    outputs(4110) <= (layer0_outputs(6782)) and not (layer0_outputs(2331));
    outputs(4111) <= layer0_outputs(5506);
    outputs(4112) <= not(layer0_outputs(5141));
    outputs(4113) <= not(layer0_outputs(1558));
    outputs(4114) <= not(layer0_outputs(8376));
    outputs(4115) <= not((layer0_outputs(4309)) or (layer0_outputs(710)));
    outputs(4116) <= (layer0_outputs(9473)) and not (layer0_outputs(2231));
    outputs(4117) <= layer0_outputs(1173);
    outputs(4118) <= layer0_outputs(1411);
    outputs(4119) <= (layer0_outputs(6166)) and not (layer0_outputs(11522));
    outputs(4120) <= (layer0_outputs(8276)) or (layer0_outputs(10711));
    outputs(4121) <= (layer0_outputs(12680)) and not (layer0_outputs(9050));
    outputs(4122) <= (layer0_outputs(8107)) xor (layer0_outputs(2185));
    outputs(4123) <= (layer0_outputs(1193)) and not (layer0_outputs(11167));
    outputs(4124) <= (layer0_outputs(12778)) xor (layer0_outputs(10893));
    outputs(4125) <= not(layer0_outputs(8940)) or (layer0_outputs(3862));
    outputs(4126) <= (layer0_outputs(11628)) or (layer0_outputs(10736));
    outputs(4127) <= layer0_outputs(9727);
    outputs(4128) <= (layer0_outputs(762)) xor (layer0_outputs(12288));
    outputs(4129) <= not(layer0_outputs(10621));
    outputs(4130) <= not((layer0_outputs(5734)) xor (layer0_outputs(4459)));
    outputs(4131) <= not(layer0_outputs(637)) or (layer0_outputs(11085));
    outputs(4132) <= (layer0_outputs(5976)) xor (layer0_outputs(8443));
    outputs(4133) <= layer0_outputs(7346);
    outputs(4134) <= (layer0_outputs(11928)) xor (layer0_outputs(3911));
    outputs(4135) <= not(layer0_outputs(8244));
    outputs(4136) <= not(layer0_outputs(368));
    outputs(4137) <= not((layer0_outputs(1111)) or (layer0_outputs(12525)));
    outputs(4138) <= layer0_outputs(12453);
    outputs(4139) <= layer0_outputs(137);
    outputs(4140) <= not(layer0_outputs(6649));
    outputs(4141) <= not(layer0_outputs(3340));
    outputs(4142) <= layer0_outputs(6686);
    outputs(4143) <= (layer0_outputs(3667)) xor (layer0_outputs(6027));
    outputs(4144) <= not(layer0_outputs(12514)) or (layer0_outputs(6958));
    outputs(4145) <= (layer0_outputs(3416)) and (layer0_outputs(8824));
    outputs(4146) <= layer0_outputs(10792);
    outputs(4147) <= not((layer0_outputs(3531)) or (layer0_outputs(9522)));
    outputs(4148) <= not(layer0_outputs(728));
    outputs(4149) <= not(layer0_outputs(6654)) or (layer0_outputs(10812));
    outputs(4150) <= not(layer0_outputs(3478));
    outputs(4151) <= not(layer0_outputs(5421));
    outputs(4152) <= not((layer0_outputs(4153)) xor (layer0_outputs(2753)));
    outputs(4153) <= not(layer0_outputs(6026)) or (layer0_outputs(2809));
    outputs(4154) <= not(layer0_outputs(3117)) or (layer0_outputs(7984));
    outputs(4155) <= not((layer0_outputs(9317)) or (layer0_outputs(6611)));
    outputs(4156) <= not((layer0_outputs(6771)) or (layer0_outputs(3902)));
    outputs(4157) <= (layer0_outputs(11250)) and (layer0_outputs(7044));
    outputs(4158) <= not(layer0_outputs(8464)) or (layer0_outputs(6954));
    outputs(4159) <= not((layer0_outputs(4945)) xor (layer0_outputs(7322)));
    outputs(4160) <= not(layer0_outputs(11149));
    outputs(4161) <= layer0_outputs(4310);
    outputs(4162) <= layer0_outputs(10121);
    outputs(4163) <= not(layer0_outputs(2483));
    outputs(4164) <= (layer0_outputs(11043)) and not (layer0_outputs(1404));
    outputs(4165) <= not(layer0_outputs(12248)) or (layer0_outputs(7567));
    outputs(4166) <= (layer0_outputs(7087)) or (layer0_outputs(10448));
    outputs(4167) <= not((layer0_outputs(11966)) xor (layer0_outputs(847)));
    outputs(4168) <= not(layer0_outputs(4079));
    outputs(4169) <= not((layer0_outputs(3237)) xor (layer0_outputs(9325)));
    outputs(4170) <= not(layer0_outputs(3381)) or (layer0_outputs(7108));
    outputs(4171) <= layer0_outputs(5363);
    outputs(4172) <= (layer0_outputs(9529)) and (layer0_outputs(2472));
    outputs(4173) <= layer0_outputs(7457);
    outputs(4174) <= not((layer0_outputs(3868)) xor (layer0_outputs(12717)));
    outputs(4175) <= layer0_outputs(12565);
    outputs(4176) <= (layer0_outputs(9554)) or (layer0_outputs(12278));
    outputs(4177) <= (layer0_outputs(10788)) and (layer0_outputs(9504));
    outputs(4178) <= (layer0_outputs(10021)) xor (layer0_outputs(1976));
    outputs(4179) <= not(layer0_outputs(3387)) or (layer0_outputs(3880));
    outputs(4180) <= not((layer0_outputs(7578)) or (layer0_outputs(2235)));
    outputs(4181) <= (layer0_outputs(2330)) xor (layer0_outputs(6439));
    outputs(4182) <= not(layer0_outputs(7192));
    outputs(4183) <= not((layer0_outputs(7335)) and (layer0_outputs(1220)));
    outputs(4184) <= not(layer0_outputs(2107)) or (layer0_outputs(11939));
    outputs(4185) <= not(layer0_outputs(2483));
    outputs(4186) <= (layer0_outputs(5025)) or (layer0_outputs(7140));
    outputs(4187) <= not(layer0_outputs(5470));
    outputs(4188) <= not((layer0_outputs(1317)) and (layer0_outputs(4237)));
    outputs(4189) <= layer0_outputs(11383);
    outputs(4190) <= (layer0_outputs(12173)) and not (layer0_outputs(8355));
    outputs(4191) <= layer0_outputs(1897);
    outputs(4192) <= not(layer0_outputs(1840));
    outputs(4193) <= not(layer0_outputs(3323));
    outputs(4194) <= layer0_outputs(5014);
    outputs(4195) <= (layer0_outputs(11373)) or (layer0_outputs(1042));
    outputs(4196) <= not(layer0_outputs(10084));
    outputs(4197) <= not(layer0_outputs(7126)) or (layer0_outputs(11518));
    outputs(4198) <= (layer0_outputs(9789)) or (layer0_outputs(2571));
    outputs(4199) <= layer0_outputs(12139);
    outputs(4200) <= not(layer0_outputs(3247));
    outputs(4201) <= (layer0_outputs(8273)) and not (layer0_outputs(9279));
    outputs(4202) <= layer0_outputs(5018);
    outputs(4203) <= not((layer0_outputs(5784)) and (layer0_outputs(4261)));
    outputs(4204) <= layer0_outputs(9713);
    outputs(4205) <= layer0_outputs(10681);
    outputs(4206) <= not((layer0_outputs(12593)) xor (layer0_outputs(4670)));
    outputs(4207) <= not((layer0_outputs(6339)) or (layer0_outputs(9051)));
    outputs(4208) <= (layer0_outputs(10697)) xor (layer0_outputs(4581));
    outputs(4209) <= layer0_outputs(3778);
    outputs(4210) <= layer0_outputs(1273);
    outputs(4211) <= not(layer0_outputs(4357)) or (layer0_outputs(11039));
    outputs(4212) <= not((layer0_outputs(1435)) xor (layer0_outputs(4516)));
    outputs(4213) <= not((layer0_outputs(6119)) and (layer0_outputs(4414)));
    outputs(4214) <= (layer0_outputs(3116)) and not (layer0_outputs(4844));
    outputs(4215) <= layer0_outputs(1197);
    outputs(4216) <= layer0_outputs(10535);
    outputs(4217) <= (layer0_outputs(10367)) or (layer0_outputs(256));
    outputs(4218) <= not((layer0_outputs(12442)) xor (layer0_outputs(10396)));
    outputs(4219) <= not(layer0_outputs(11583));
    outputs(4220) <= layer0_outputs(8887);
    outputs(4221) <= not((layer0_outputs(8992)) or (layer0_outputs(96)));
    outputs(4222) <= (layer0_outputs(861)) or (layer0_outputs(2238));
    outputs(4223) <= layer0_outputs(11408);
    outputs(4224) <= (layer0_outputs(257)) xor (layer0_outputs(11468));
    outputs(4225) <= '1';
    outputs(4226) <= (layer0_outputs(553)) and not (layer0_outputs(2740));
    outputs(4227) <= not((layer0_outputs(5076)) or (layer0_outputs(848)));
    outputs(4228) <= layer0_outputs(4356);
    outputs(4229) <= layer0_outputs(12734);
    outputs(4230) <= not(layer0_outputs(2768));
    outputs(4231) <= not(layer0_outputs(4949));
    outputs(4232) <= '1';
    outputs(4233) <= layer0_outputs(9868);
    outputs(4234) <= layer0_outputs(7714);
    outputs(4235) <= (layer0_outputs(9454)) and not (layer0_outputs(2922));
    outputs(4236) <= not((layer0_outputs(9538)) xor (layer0_outputs(7936)));
    outputs(4237) <= layer0_outputs(6516);
    outputs(4238) <= not(layer0_outputs(3626));
    outputs(4239) <= (layer0_outputs(2857)) xor (layer0_outputs(11361));
    outputs(4240) <= not((layer0_outputs(9932)) xor (layer0_outputs(621)));
    outputs(4241) <= not((layer0_outputs(10593)) xor (layer0_outputs(813)));
    outputs(4242) <= (layer0_outputs(1736)) and not (layer0_outputs(4738));
    outputs(4243) <= layer0_outputs(3493);
    outputs(4244) <= not(layer0_outputs(6610));
    outputs(4245) <= not(layer0_outputs(1696));
    outputs(4246) <= (layer0_outputs(7375)) and (layer0_outputs(3365));
    outputs(4247) <= (layer0_outputs(8155)) and not (layer0_outputs(9385));
    outputs(4248) <= not((layer0_outputs(4216)) or (layer0_outputs(380)));
    outputs(4249) <= (layer0_outputs(3817)) xor (layer0_outputs(11865));
    outputs(4250) <= (layer0_outputs(7626)) and not (layer0_outputs(9297));
    outputs(4251) <= layer0_outputs(10475);
    outputs(4252) <= layer0_outputs(6500);
    outputs(4253) <= (layer0_outputs(6638)) or (layer0_outputs(5254));
    outputs(4254) <= not(layer0_outputs(9283));
    outputs(4255) <= layer0_outputs(11854);
    outputs(4256) <= not(layer0_outputs(2945));
    outputs(4257) <= (layer0_outputs(4005)) xor (layer0_outputs(8294));
    outputs(4258) <= (layer0_outputs(3993)) or (layer0_outputs(8830));
    outputs(4259) <= not(layer0_outputs(1106)) or (layer0_outputs(3257));
    outputs(4260) <= not((layer0_outputs(4108)) or (layer0_outputs(2967)));
    outputs(4261) <= layer0_outputs(10414);
    outputs(4262) <= not(layer0_outputs(4202));
    outputs(4263) <= (layer0_outputs(12103)) and (layer0_outputs(2465));
    outputs(4264) <= layer0_outputs(661);
    outputs(4265) <= layer0_outputs(5285);
    outputs(4266) <= layer0_outputs(5140);
    outputs(4267) <= layer0_outputs(558);
    outputs(4268) <= (layer0_outputs(1079)) and (layer0_outputs(1880));
    outputs(4269) <= not((layer0_outputs(7058)) or (layer0_outputs(4691)));
    outputs(4270) <= layer0_outputs(4243);
    outputs(4271) <= layer0_outputs(10420);
    outputs(4272) <= not(layer0_outputs(5379));
    outputs(4273) <= (layer0_outputs(9373)) and not (layer0_outputs(10002));
    outputs(4274) <= layer0_outputs(4313);
    outputs(4275) <= (layer0_outputs(3056)) xor (layer0_outputs(12137));
    outputs(4276) <= layer0_outputs(2914);
    outputs(4277) <= (layer0_outputs(11300)) or (layer0_outputs(707));
    outputs(4278) <= not((layer0_outputs(9124)) and (layer0_outputs(4728)));
    outputs(4279) <= layer0_outputs(5604);
    outputs(4280) <= not((layer0_outputs(113)) or (layer0_outputs(3738)));
    outputs(4281) <= not((layer0_outputs(5243)) xor (layer0_outputs(9718)));
    outputs(4282) <= not((layer0_outputs(9239)) xor (layer0_outputs(9559)));
    outputs(4283) <= not(layer0_outputs(9672)) or (layer0_outputs(4350));
    outputs(4284) <= layer0_outputs(12116);
    outputs(4285) <= not((layer0_outputs(3151)) and (layer0_outputs(8562)));
    outputs(4286) <= not((layer0_outputs(5045)) xor (layer0_outputs(7614)));
    outputs(4287) <= (layer0_outputs(10057)) xor (layer0_outputs(8935));
    outputs(4288) <= (layer0_outputs(254)) and not (layer0_outputs(4901));
    outputs(4289) <= not(layer0_outputs(6357)) or (layer0_outputs(5236));
    outputs(4290) <= layer0_outputs(11256);
    outputs(4291) <= not(layer0_outputs(3973));
    outputs(4292) <= not((layer0_outputs(7239)) and (layer0_outputs(11549)));
    outputs(4293) <= (layer0_outputs(2402)) xor (layer0_outputs(8819));
    outputs(4294) <= layer0_outputs(3947);
    outputs(4295) <= (layer0_outputs(3647)) or (layer0_outputs(4615));
    outputs(4296) <= not(layer0_outputs(10073)) or (layer0_outputs(2664));
    outputs(4297) <= (layer0_outputs(5946)) xor (layer0_outputs(11374));
    outputs(4298) <= not(layer0_outputs(5298));
    outputs(4299) <= not(layer0_outputs(1829)) or (layer0_outputs(10836));
    outputs(4300) <= layer0_outputs(1099);
    outputs(4301) <= (layer0_outputs(4080)) or (layer0_outputs(10077));
    outputs(4302) <= layer0_outputs(11890);
    outputs(4303) <= not((layer0_outputs(10807)) or (layer0_outputs(8665)));
    outputs(4304) <= not(layer0_outputs(11104));
    outputs(4305) <= (layer0_outputs(6942)) or (layer0_outputs(2041));
    outputs(4306) <= not(layer0_outputs(9825));
    outputs(4307) <= layer0_outputs(1695);
    outputs(4308) <= layer0_outputs(2579);
    outputs(4309) <= (layer0_outputs(12064)) and not (layer0_outputs(12274));
    outputs(4310) <= not((layer0_outputs(4540)) or (layer0_outputs(9344)));
    outputs(4311) <= not(layer0_outputs(12045)) or (layer0_outputs(4581));
    outputs(4312) <= layer0_outputs(11726);
    outputs(4313) <= not(layer0_outputs(11775));
    outputs(4314) <= layer0_outputs(4082);
    outputs(4315) <= not((layer0_outputs(11981)) xor (layer0_outputs(586)));
    outputs(4316) <= not(layer0_outputs(2291));
    outputs(4317) <= layer0_outputs(6919);
    outputs(4318) <= not((layer0_outputs(9260)) and (layer0_outputs(3312)));
    outputs(4319) <= (layer0_outputs(4868)) and (layer0_outputs(12218));
    outputs(4320) <= not(layer0_outputs(9326)) or (layer0_outputs(5780));
    outputs(4321) <= not(layer0_outputs(11889)) or (layer0_outputs(7551));
    outputs(4322) <= (layer0_outputs(8378)) xor (layer0_outputs(4736));
    outputs(4323) <= layer0_outputs(6458);
    outputs(4324) <= not((layer0_outputs(12127)) xor (layer0_outputs(11828)));
    outputs(4325) <= not(layer0_outputs(12382));
    outputs(4326) <= not(layer0_outputs(3362)) or (layer0_outputs(10421));
    outputs(4327) <= (layer0_outputs(422)) or (layer0_outputs(10825));
    outputs(4328) <= layer0_outputs(6930);
    outputs(4329) <= not((layer0_outputs(5535)) and (layer0_outputs(1501)));
    outputs(4330) <= not((layer0_outputs(2203)) xor (layer0_outputs(9764)));
    outputs(4331) <= (layer0_outputs(7088)) xor (layer0_outputs(12635));
    outputs(4332) <= layer0_outputs(5681);
    outputs(4333) <= layer0_outputs(5145);
    outputs(4334) <= not(layer0_outputs(8203));
    outputs(4335) <= (layer0_outputs(11061)) xor (layer0_outputs(7293));
    outputs(4336) <= not(layer0_outputs(2113));
    outputs(4337) <= (layer0_outputs(9096)) and (layer0_outputs(9043));
    outputs(4338) <= not((layer0_outputs(7513)) xor (layer0_outputs(11255)));
    outputs(4339) <= not(layer0_outputs(4045));
    outputs(4340) <= (layer0_outputs(4749)) xor (layer0_outputs(8035));
    outputs(4341) <= not((layer0_outputs(1990)) xor (layer0_outputs(6104)));
    outputs(4342) <= not(layer0_outputs(11446)) or (layer0_outputs(1328));
    outputs(4343) <= not(layer0_outputs(10294));
    outputs(4344) <= (layer0_outputs(7644)) and (layer0_outputs(1260));
    outputs(4345) <= (layer0_outputs(2962)) and not (layer0_outputs(7372));
    outputs(4346) <= not((layer0_outputs(5874)) xor (layer0_outputs(7706)));
    outputs(4347) <= (layer0_outputs(9358)) and not (layer0_outputs(4033));
    outputs(4348) <= (layer0_outputs(365)) and not (layer0_outputs(10294));
    outputs(4349) <= not((layer0_outputs(12623)) xor (layer0_outputs(1417)));
    outputs(4350) <= (layer0_outputs(1943)) xor (layer0_outputs(8016));
    outputs(4351) <= not(layer0_outputs(7674));
    outputs(4352) <= layer0_outputs(3412);
    outputs(4353) <= not((layer0_outputs(1003)) or (layer0_outputs(5079)));
    outputs(4354) <= (layer0_outputs(11772)) or (layer0_outputs(8867));
    outputs(4355) <= layer0_outputs(8614);
    outputs(4356) <= not(layer0_outputs(7917));
    outputs(4357) <= not((layer0_outputs(1307)) xor (layer0_outputs(12751)));
    outputs(4358) <= not(layer0_outputs(7610));
    outputs(4359) <= not(layer0_outputs(9514));
    outputs(4360) <= layer0_outputs(6795);
    outputs(4361) <= (layer0_outputs(1408)) and not (layer0_outputs(2865));
    outputs(4362) <= not(layer0_outputs(9048));
    outputs(4363) <= not((layer0_outputs(1385)) xor (layer0_outputs(1409)));
    outputs(4364) <= not(layer0_outputs(7642));
    outputs(4365) <= not(layer0_outputs(9352)) or (layer0_outputs(8829));
    outputs(4366) <= not(layer0_outputs(10387));
    outputs(4367) <= not(layer0_outputs(3143)) or (layer0_outputs(9091));
    outputs(4368) <= layer0_outputs(6230);
    outputs(4369) <= '0';
    outputs(4370) <= layer0_outputs(8341);
    outputs(4371) <= not((layer0_outputs(2993)) xor (layer0_outputs(2884)));
    outputs(4372) <= (layer0_outputs(1671)) xor (layer0_outputs(11673));
    outputs(4373) <= not((layer0_outputs(8303)) and (layer0_outputs(4539)));
    outputs(4374) <= not((layer0_outputs(10777)) and (layer0_outputs(4529)));
    outputs(4375) <= not(layer0_outputs(1957)) or (layer0_outputs(2486));
    outputs(4376) <= (layer0_outputs(626)) and (layer0_outputs(9754));
    outputs(4377) <= not(layer0_outputs(10623));
    outputs(4378) <= not(layer0_outputs(6694));
    outputs(4379) <= layer0_outputs(2190);
    outputs(4380) <= (layer0_outputs(8851)) xor (layer0_outputs(4599));
    outputs(4381) <= (layer0_outputs(10111)) or (layer0_outputs(11835));
    outputs(4382) <= not(layer0_outputs(3870));
    outputs(4383) <= not(layer0_outputs(9262));
    outputs(4384) <= not((layer0_outputs(11012)) xor (layer0_outputs(6172)));
    outputs(4385) <= not(layer0_outputs(7321));
    outputs(4386) <= (layer0_outputs(10661)) or (layer0_outputs(6982));
    outputs(4387) <= not((layer0_outputs(9541)) and (layer0_outputs(10249)));
    outputs(4388) <= (layer0_outputs(7718)) or (layer0_outputs(8644));
    outputs(4389) <= not(layer0_outputs(2524)) or (layer0_outputs(11203));
    outputs(4390) <= (layer0_outputs(8911)) xor (layer0_outputs(11514));
    outputs(4391) <= not(layer0_outputs(2517));
    outputs(4392) <= not(layer0_outputs(5030));
    outputs(4393) <= '1';
    outputs(4394) <= '1';
    outputs(4395) <= layer0_outputs(3210);
    outputs(4396) <= not((layer0_outputs(4120)) xor (layer0_outputs(1195)));
    outputs(4397) <= not(layer0_outputs(9242));
    outputs(4398) <= layer0_outputs(2549);
    outputs(4399) <= not(layer0_outputs(5489)) or (layer0_outputs(12305));
    outputs(4400) <= not(layer0_outputs(279)) or (layer0_outputs(623));
    outputs(4401) <= (layer0_outputs(5221)) xor (layer0_outputs(6355));
    outputs(4402) <= not(layer0_outputs(12728));
    outputs(4403) <= (layer0_outputs(237)) and (layer0_outputs(5283));
    outputs(4404) <= layer0_outputs(11016);
    outputs(4405) <= not(layer0_outputs(3992)) or (layer0_outputs(3530));
    outputs(4406) <= not((layer0_outputs(1941)) xor (layer0_outputs(11448)));
    outputs(4407) <= not(layer0_outputs(5620));
    outputs(4408) <= layer0_outputs(7772);
    outputs(4409) <= not((layer0_outputs(10674)) and (layer0_outputs(12777)));
    outputs(4410) <= (layer0_outputs(11902)) or (layer0_outputs(5805));
    outputs(4411) <= (layer0_outputs(263)) and (layer0_outputs(7269));
    outputs(4412) <= (layer0_outputs(658)) and not (layer0_outputs(1164));
    outputs(4413) <= layer0_outputs(12285);
    outputs(4414) <= not(layer0_outputs(5537));
    outputs(4415) <= not(layer0_outputs(2045));
    outputs(4416) <= layer0_outputs(5593);
    outputs(4417) <= not((layer0_outputs(4346)) xor (layer0_outputs(5981)));
    outputs(4418) <= not((layer0_outputs(11088)) and (layer0_outputs(10353)));
    outputs(4419) <= not(layer0_outputs(4592));
    outputs(4420) <= not((layer0_outputs(4347)) xor (layer0_outputs(442)));
    outputs(4421) <= not(layer0_outputs(7127)) or (layer0_outputs(5738));
    outputs(4422) <= not(layer0_outputs(12275));
    outputs(4423) <= (layer0_outputs(4333)) xor (layer0_outputs(10446));
    outputs(4424) <= layer0_outputs(9492);
    outputs(4425) <= not((layer0_outputs(5652)) xor (layer0_outputs(3181)));
    outputs(4426) <= (layer0_outputs(3920)) xor (layer0_outputs(3619));
    outputs(4427) <= not((layer0_outputs(9408)) and (layer0_outputs(12653)));
    outputs(4428) <= not(layer0_outputs(11138)) or (layer0_outputs(8962));
    outputs(4429) <= (layer0_outputs(4046)) xor (layer0_outputs(10109));
    outputs(4430) <= not(layer0_outputs(663));
    outputs(4431) <= not(layer0_outputs(11971));
    outputs(4432) <= layer0_outputs(3818);
    outputs(4433) <= not(layer0_outputs(7590)) or (layer0_outputs(11037));
    outputs(4434) <= (layer0_outputs(4775)) and not (layer0_outputs(8529));
    outputs(4435) <= not(layer0_outputs(2851)) or (layer0_outputs(4742));
    outputs(4436) <= not((layer0_outputs(6869)) xor (layer0_outputs(12559)));
    outputs(4437) <= layer0_outputs(10309);
    outputs(4438) <= (layer0_outputs(8374)) xor (layer0_outputs(961));
    outputs(4439) <= not(layer0_outputs(5818));
    outputs(4440) <= not(layer0_outputs(9405));
    outputs(4441) <= (layer0_outputs(984)) xor (layer0_outputs(521));
    outputs(4442) <= layer0_outputs(5223);
    outputs(4443) <= (layer0_outputs(1038)) and not (layer0_outputs(5365));
    outputs(4444) <= layer0_outputs(6715);
    outputs(4445) <= not(layer0_outputs(11973));
    outputs(4446) <= not((layer0_outputs(3413)) xor (layer0_outputs(11801)));
    outputs(4447) <= not((layer0_outputs(8677)) and (layer0_outputs(9119)));
    outputs(4448) <= (layer0_outputs(1242)) and (layer0_outputs(5533));
    outputs(4449) <= not((layer0_outputs(345)) xor (layer0_outputs(9440)));
    outputs(4450) <= not(layer0_outputs(789)) or (layer0_outputs(326));
    outputs(4451) <= (layer0_outputs(5921)) and not (layer0_outputs(6078));
    outputs(4452) <= (layer0_outputs(10824)) or (layer0_outputs(10660));
    outputs(4453) <= layer0_outputs(11671);
    outputs(4454) <= not((layer0_outputs(3759)) xor (layer0_outputs(1304)));
    outputs(4455) <= not(layer0_outputs(12754));
    outputs(4456) <= not(layer0_outputs(11979));
    outputs(4457) <= (layer0_outputs(12618)) and not (layer0_outputs(11837));
    outputs(4458) <= layer0_outputs(4761);
    outputs(4459) <= not(layer0_outputs(6734));
    outputs(4460) <= not(layer0_outputs(3273)) or (layer0_outputs(5300));
    outputs(4461) <= not((layer0_outputs(3766)) xor (layer0_outputs(3864)));
    outputs(4462) <= not((layer0_outputs(4971)) or (layer0_outputs(12438)));
    outputs(4463) <= layer0_outputs(4777);
    outputs(4464) <= (layer0_outputs(1719)) xor (layer0_outputs(5999));
    outputs(4465) <= not((layer0_outputs(3183)) xor (layer0_outputs(11651)));
    outputs(4466) <= not(layer0_outputs(7836));
    outputs(4467) <= layer0_outputs(11872);
    outputs(4468) <= not((layer0_outputs(8969)) xor (layer0_outputs(5164)));
    outputs(4469) <= (layer0_outputs(616)) or (layer0_outputs(11575));
    outputs(4470) <= layer0_outputs(10081);
    outputs(4471) <= not(layer0_outputs(12161));
    outputs(4472) <= not((layer0_outputs(82)) xor (layer0_outputs(0)));
    outputs(4473) <= (layer0_outputs(7244)) and (layer0_outputs(7515));
    outputs(4474) <= not((layer0_outputs(892)) or (layer0_outputs(5772)));
    outputs(4475) <= (layer0_outputs(7754)) xor (layer0_outputs(9134));
    outputs(4476) <= not(layer0_outputs(2339)) or (layer0_outputs(6849));
    outputs(4477) <= layer0_outputs(2093);
    outputs(4478) <= not((layer0_outputs(3327)) xor (layer0_outputs(6277)));
    outputs(4479) <= (layer0_outputs(1407)) or (layer0_outputs(3423));
    outputs(4480) <= layer0_outputs(11137);
    outputs(4481) <= layer0_outputs(11466);
    outputs(4482) <= (layer0_outputs(4680)) or (layer0_outputs(1188));
    outputs(4483) <= not((layer0_outputs(5927)) xor (layer0_outputs(7952)));
    outputs(4484) <= layer0_outputs(6421);
    outputs(4485) <= not(layer0_outputs(10815));
    outputs(4486) <= not((layer0_outputs(4433)) xor (layer0_outputs(9249)));
    outputs(4487) <= not(layer0_outputs(810)) or (layer0_outputs(7531));
    outputs(4488) <= (layer0_outputs(11795)) and not (layer0_outputs(10309));
    outputs(4489) <= (layer0_outputs(7003)) and (layer0_outputs(8307));
    outputs(4490) <= (layer0_outputs(4607)) and not (layer0_outputs(4748));
    outputs(4491) <= (layer0_outputs(4493)) xor (layer0_outputs(2327));
    outputs(4492) <= (layer0_outputs(6742)) xor (layer0_outputs(824));
    outputs(4493) <= not((layer0_outputs(11338)) xor (layer0_outputs(10968)));
    outputs(4494) <= '1';
    outputs(4495) <= not(layer0_outputs(8490));
    outputs(4496) <= (layer0_outputs(926)) xor (layer0_outputs(6156));
    outputs(4497) <= layer0_outputs(11120);
    outputs(4498) <= layer0_outputs(3090);
    outputs(4499) <= not(layer0_outputs(8650));
    outputs(4500) <= not((layer0_outputs(2797)) xor (layer0_outputs(11926)));
    outputs(4501) <= not((layer0_outputs(6569)) or (layer0_outputs(7012)));
    outputs(4502) <= layer0_outputs(12186);
    outputs(4503) <= (layer0_outputs(5974)) xor (layer0_outputs(9858));
    outputs(4504) <= not(layer0_outputs(7668));
    outputs(4505) <= not((layer0_outputs(6102)) xor (layer0_outputs(4886)));
    outputs(4506) <= (layer0_outputs(11191)) or (layer0_outputs(6110));
    outputs(4507) <= not((layer0_outputs(8408)) and (layer0_outputs(4291)));
    outputs(4508) <= not(layer0_outputs(9168));
    outputs(4509) <= not(layer0_outputs(3326));
    outputs(4510) <= not(layer0_outputs(8493));
    outputs(4511) <= layer0_outputs(11329);
    outputs(4512) <= not((layer0_outputs(11105)) xor (layer0_outputs(4978)));
    outputs(4513) <= (layer0_outputs(5101)) and not (layer0_outputs(3892));
    outputs(4514) <= (layer0_outputs(6367)) xor (layer0_outputs(933));
    outputs(4515) <= not((layer0_outputs(9484)) xor (layer0_outputs(2799)));
    outputs(4516) <= not(layer0_outputs(7116));
    outputs(4517) <= (layer0_outputs(9355)) xor (layer0_outputs(6470));
    outputs(4518) <= not(layer0_outputs(11328)) or (layer0_outputs(5900));
    outputs(4519) <= (layer0_outputs(10555)) xor (layer0_outputs(9643));
    outputs(4520) <= (layer0_outputs(3976)) xor (layer0_outputs(9323));
    outputs(4521) <= not((layer0_outputs(7857)) xor (layer0_outputs(9595)));
    outputs(4522) <= not((layer0_outputs(12259)) xor (layer0_outputs(4004)));
    outputs(4523) <= layer0_outputs(9258);
    outputs(4524) <= not(layer0_outputs(12494)) or (layer0_outputs(1130));
    outputs(4525) <= not(layer0_outputs(7895));
    outputs(4526) <= (layer0_outputs(4522)) xor (layer0_outputs(12114));
    outputs(4527) <= layer0_outputs(3139);
    outputs(4528) <= not((layer0_outputs(3995)) xor (layer0_outputs(2709)));
    outputs(4529) <= (layer0_outputs(9028)) xor (layer0_outputs(2667));
    outputs(4530) <= not((layer0_outputs(8099)) and (layer0_outputs(2771)));
    outputs(4531) <= not((layer0_outputs(9108)) or (layer0_outputs(5881)));
    outputs(4532) <= (layer0_outputs(5762)) and not (layer0_outputs(10675));
    outputs(4533) <= layer0_outputs(1689);
    outputs(4534) <= not(layer0_outputs(311));
    outputs(4535) <= (layer0_outputs(2427)) and not (layer0_outputs(7574));
    outputs(4536) <= (layer0_outputs(3955)) xor (layer0_outputs(1280));
    outputs(4537) <= not(layer0_outputs(8611));
    outputs(4538) <= (layer0_outputs(11928)) and not (layer0_outputs(10856));
    outputs(4539) <= (layer0_outputs(4384)) or (layer0_outputs(10017));
    outputs(4540) <= layer0_outputs(9630);
    outputs(4541) <= layer0_outputs(2267);
    outputs(4542) <= '1';
    outputs(4543) <= not(layer0_outputs(3180)) or (layer0_outputs(12033));
    outputs(4544) <= (layer0_outputs(3803)) and not (layer0_outputs(7525));
    outputs(4545) <= (layer0_outputs(2630)) or (layer0_outputs(11830));
    outputs(4546) <= not(layer0_outputs(8523));
    outputs(4547) <= not((layer0_outputs(4573)) xor (layer0_outputs(332)));
    outputs(4548) <= not(layer0_outputs(5873));
    outputs(4549) <= (layer0_outputs(7294)) xor (layer0_outputs(8724));
    outputs(4550) <= not((layer0_outputs(4359)) xor (layer0_outputs(5331)));
    outputs(4551) <= (layer0_outputs(4544)) and (layer0_outputs(7024));
    outputs(4552) <= not((layer0_outputs(12464)) xor (layer0_outputs(8459)));
    outputs(4553) <= not((layer0_outputs(1725)) and (layer0_outputs(4116)));
    outputs(4554) <= layer0_outputs(2061);
    outputs(4555) <= (layer0_outputs(10871)) xor (layer0_outputs(7307));
    outputs(4556) <= (layer0_outputs(5713)) xor (layer0_outputs(4937));
    outputs(4557) <= not(layer0_outputs(5145)) or (layer0_outputs(3548));
    outputs(4558) <= not(layer0_outputs(3016)) or (layer0_outputs(12369));
    outputs(4559) <= not(layer0_outputs(1199));
    outputs(4560) <= not(layer0_outputs(6242));
    outputs(4561) <= (layer0_outputs(3953)) and (layer0_outputs(10507));
    outputs(4562) <= not((layer0_outputs(6085)) or (layer0_outputs(2956)));
    outputs(4563) <= not(layer0_outputs(10146));
    outputs(4564) <= not((layer0_outputs(6094)) xor (layer0_outputs(6719)));
    outputs(4565) <= '1';
    outputs(4566) <= (layer0_outputs(4547)) and not (layer0_outputs(10923));
    outputs(4567) <= not(layer0_outputs(360));
    outputs(4568) <= not(layer0_outputs(3676));
    outputs(4569) <= (layer0_outputs(3871)) xor (layer0_outputs(4472));
    outputs(4570) <= (layer0_outputs(3201)) xor (layer0_outputs(7963));
    outputs(4571) <= layer0_outputs(3400);
    outputs(4572) <= layer0_outputs(867);
    outputs(4573) <= (layer0_outputs(8574)) xor (layer0_outputs(2021));
    outputs(4574) <= (layer0_outputs(7665)) and not (layer0_outputs(3219));
    outputs(4575) <= not((layer0_outputs(3841)) xor (layer0_outputs(2666)));
    outputs(4576) <= layer0_outputs(10561);
    outputs(4577) <= (layer0_outputs(11597)) xor (layer0_outputs(12732));
    outputs(4578) <= layer0_outputs(10534);
    outputs(4579) <= not((layer0_outputs(11559)) or (layer0_outputs(9012)));
    outputs(4580) <= not((layer0_outputs(6556)) or (layer0_outputs(3428)));
    outputs(4581) <= (layer0_outputs(12794)) and not (layer0_outputs(671));
    outputs(4582) <= not(layer0_outputs(6582));
    outputs(4583) <= layer0_outputs(10663);
    outputs(4584) <= not(layer0_outputs(6512)) or (layer0_outputs(7474));
    outputs(4585) <= not(layer0_outputs(6550));
    outputs(4586) <= layer0_outputs(1419);
    outputs(4587) <= (layer0_outputs(10984)) xor (layer0_outputs(7666));
    outputs(4588) <= layer0_outputs(5399);
    outputs(4589) <= not((layer0_outputs(4029)) and (layer0_outputs(5290)));
    outputs(4590) <= (layer0_outputs(11682)) xor (layer0_outputs(6897));
    outputs(4591) <= layer0_outputs(10969);
    outputs(4592) <= not(layer0_outputs(12677));
    outputs(4593) <= not(layer0_outputs(2160));
    outputs(4594) <= not(layer0_outputs(7827)) or (layer0_outputs(3905));
    outputs(4595) <= (layer0_outputs(5554)) or (layer0_outputs(9568));
    outputs(4596) <= not((layer0_outputs(7552)) xor (layer0_outputs(1281)));
    outputs(4597) <= (layer0_outputs(12154)) xor (layer0_outputs(4112));
    outputs(4598) <= (layer0_outputs(7568)) and (layer0_outputs(8964));
    outputs(4599) <= not(layer0_outputs(7461));
    outputs(4600) <= not(layer0_outputs(8302));
    outputs(4601) <= (layer0_outputs(9322)) or (layer0_outputs(10425));
    outputs(4602) <= layer0_outputs(1324);
    outputs(4603) <= (layer0_outputs(4963)) and (layer0_outputs(3663));
    outputs(4604) <= (layer0_outputs(8270)) xor (layer0_outputs(7690));
    outputs(4605) <= layer0_outputs(1831);
    outputs(4606) <= not((layer0_outputs(2003)) xor (layer0_outputs(5635)));
    outputs(4607) <= not(layer0_outputs(7590)) or (layer0_outputs(264));
    outputs(4608) <= not(layer0_outputs(10996)) or (layer0_outputs(10943));
    outputs(4609) <= (layer0_outputs(4694)) or (layer0_outputs(7428));
    outputs(4610) <= not(layer0_outputs(624));
    outputs(4611) <= layer0_outputs(9137);
    outputs(4612) <= (layer0_outputs(5806)) xor (layer0_outputs(1061));
    outputs(4613) <= not(layer0_outputs(10492));
    outputs(4614) <= not(layer0_outputs(6306));
    outputs(4615) <= layer0_outputs(7402);
    outputs(4616) <= (layer0_outputs(12314)) xor (layer0_outputs(5723));
    outputs(4617) <= not((layer0_outputs(3728)) or (layer0_outputs(12389)));
    outputs(4618) <= (layer0_outputs(6689)) xor (layer0_outputs(11378));
    outputs(4619) <= '1';
    outputs(4620) <= layer0_outputs(7485);
    outputs(4621) <= (layer0_outputs(9166)) and not (layer0_outputs(3102));
    outputs(4622) <= (layer0_outputs(8045)) xor (layer0_outputs(10227));
    outputs(4623) <= (layer0_outputs(1582)) and not (layer0_outputs(10400));
    outputs(4624) <= layer0_outputs(9162);
    outputs(4625) <= layer0_outputs(11642);
    outputs(4626) <= (layer0_outputs(11754)) or (layer0_outputs(11266));
    outputs(4627) <= not(layer0_outputs(7063)) or (layer0_outputs(1945));
    outputs(4628) <= not(layer0_outputs(6105)) or (layer0_outputs(8514));
    outputs(4629) <= not(layer0_outputs(4540)) or (layer0_outputs(2710));
    outputs(4630) <= not((layer0_outputs(8769)) xor (layer0_outputs(376)));
    outputs(4631) <= (layer0_outputs(1329)) and (layer0_outputs(11117));
    outputs(4632) <= layer0_outputs(10908);
    outputs(4633) <= not((layer0_outputs(6891)) or (layer0_outputs(4949)));
    outputs(4634) <= layer0_outputs(5559);
    outputs(4635) <= layer0_outputs(8887);
    outputs(4636) <= (layer0_outputs(10808)) and (layer0_outputs(9106));
    outputs(4637) <= not((layer0_outputs(6221)) xor (layer0_outputs(9695)));
    outputs(4638) <= (layer0_outputs(10662)) xor (layer0_outputs(2442));
    outputs(4639) <= not((layer0_outputs(9525)) xor (layer0_outputs(4029)));
    outputs(4640) <= (layer0_outputs(1392)) or (layer0_outputs(6068));
    outputs(4641) <= (layer0_outputs(7484)) xor (layer0_outputs(2823));
    outputs(4642) <= (layer0_outputs(10892)) xor (layer0_outputs(12672));
    outputs(4643) <= layer0_outputs(9426);
    outputs(4644) <= not(layer0_outputs(9647)) or (layer0_outputs(4323));
    outputs(4645) <= layer0_outputs(2040);
    outputs(4646) <= not(layer0_outputs(7204)) or (layer0_outputs(11446));
    outputs(4647) <= not((layer0_outputs(3501)) or (layer0_outputs(6210)));
    outputs(4648) <= (layer0_outputs(6992)) xor (layer0_outputs(78));
    outputs(4649) <= not(layer0_outputs(2583));
    outputs(4650) <= not((layer0_outputs(3475)) xor (layer0_outputs(1111)));
    outputs(4651) <= not(layer0_outputs(1769)) or (layer0_outputs(7365));
    outputs(4652) <= (layer0_outputs(5767)) xor (layer0_outputs(7164));
    outputs(4653) <= not(layer0_outputs(11259)) or (layer0_outputs(3803));
    outputs(4654) <= layer0_outputs(7579);
    outputs(4655) <= layer0_outputs(9982);
    outputs(4656) <= (layer0_outputs(7977)) xor (layer0_outputs(11251));
    outputs(4657) <= not(layer0_outputs(9414)) or (layer0_outputs(5431));
    outputs(4658) <= (layer0_outputs(532)) and not (layer0_outputs(7271));
    outputs(4659) <= not(layer0_outputs(6546));
    outputs(4660) <= layer0_outputs(2999);
    outputs(4661) <= (layer0_outputs(2249)) and not (layer0_outputs(266));
    outputs(4662) <= layer0_outputs(11204);
    outputs(4663) <= not(layer0_outputs(11368));
    outputs(4664) <= (layer0_outputs(9281)) and not (layer0_outputs(3244));
    outputs(4665) <= layer0_outputs(1087);
    outputs(4666) <= layer0_outputs(9790);
    outputs(4667) <= layer0_outputs(10299);
    outputs(4668) <= not(layer0_outputs(6022));
    outputs(4669) <= layer0_outputs(12237);
    outputs(4670) <= not(layer0_outputs(3786));
    outputs(4671) <= not(layer0_outputs(195)) or (layer0_outputs(12020));
    outputs(4672) <= layer0_outputs(9073);
    outputs(4673) <= (layer0_outputs(3084)) and not (layer0_outputs(72));
    outputs(4674) <= not(layer0_outputs(9533));
    outputs(4675) <= not(layer0_outputs(9625));
    outputs(4676) <= (layer0_outputs(10026)) and (layer0_outputs(1023));
    outputs(4677) <= not((layer0_outputs(9075)) or (layer0_outputs(6983)));
    outputs(4678) <= not(layer0_outputs(1077)) or (layer0_outputs(1776));
    outputs(4679) <= (layer0_outputs(8619)) and not (layer0_outputs(9437));
    outputs(4680) <= not((layer0_outputs(5747)) xor (layer0_outputs(10840)));
    outputs(4681) <= (layer0_outputs(8427)) xor (layer0_outputs(441));
    outputs(4682) <= not(layer0_outputs(2632)) or (layer0_outputs(536));
    outputs(4683) <= not(layer0_outputs(12048));
    outputs(4684) <= (layer0_outputs(262)) and not (layer0_outputs(5541));
    outputs(4685) <= not(layer0_outputs(2253));
    outputs(4686) <= not(layer0_outputs(6196));
    outputs(4687) <= not((layer0_outputs(6845)) xor (layer0_outputs(6288)));
    outputs(4688) <= layer0_outputs(771);
    outputs(4689) <= layer0_outputs(1331);
    outputs(4690) <= (layer0_outputs(801)) and not (layer0_outputs(849));
    outputs(4691) <= not(layer0_outputs(5091));
    outputs(4692) <= (layer0_outputs(10190)) and (layer0_outputs(4698));
    outputs(4693) <= not((layer0_outputs(10553)) and (layer0_outputs(7701)));
    outputs(4694) <= not((layer0_outputs(6668)) xor (layer0_outputs(7215)));
    outputs(4695) <= not(layer0_outputs(2539));
    outputs(4696) <= not((layer0_outputs(9342)) xor (layer0_outputs(8227)));
    outputs(4697) <= not(layer0_outputs(11911)) or (layer0_outputs(7502));
    outputs(4698) <= not(layer0_outputs(8881));
    outputs(4699) <= not(layer0_outputs(1213));
    outputs(4700) <= (layer0_outputs(105)) and not (layer0_outputs(1637));
    outputs(4701) <= layer0_outputs(12667);
    outputs(4702) <= (layer0_outputs(10312)) and (layer0_outputs(8942));
    outputs(4703) <= not((layer0_outputs(1627)) xor (layer0_outputs(5577)));
    outputs(4704) <= (layer0_outputs(5657)) and (layer0_outputs(9911));
    outputs(4705) <= not(layer0_outputs(421));
    outputs(4706) <= not(layer0_outputs(5954));
    outputs(4707) <= not(layer0_outputs(5822)) or (layer0_outputs(9063));
    outputs(4708) <= not((layer0_outputs(9736)) and (layer0_outputs(5320)));
    outputs(4709) <= (layer0_outputs(6138)) xor (layer0_outputs(237));
    outputs(4710) <= layer0_outputs(11849);
    outputs(4711) <= not((layer0_outputs(1428)) and (layer0_outputs(6432)));
    outputs(4712) <= not(layer0_outputs(6091));
    outputs(4713) <= layer0_outputs(12077);
    outputs(4714) <= not((layer0_outputs(6008)) or (layer0_outputs(4318)));
    outputs(4715) <= (layer0_outputs(2968)) xor (layer0_outputs(11906));
    outputs(4716) <= layer0_outputs(6612);
    outputs(4717) <= (layer0_outputs(4443)) and not (layer0_outputs(9288));
    outputs(4718) <= not(layer0_outputs(2478)) or (layer0_outputs(10462));
    outputs(4719) <= (layer0_outputs(1143)) xor (layer0_outputs(2214));
    outputs(4720) <= layer0_outputs(5444);
    outputs(4721) <= (layer0_outputs(981)) xor (layer0_outputs(642));
    outputs(4722) <= not((layer0_outputs(7696)) xor (layer0_outputs(9146)));
    outputs(4723) <= not(layer0_outputs(2590)) or (layer0_outputs(9883));
    outputs(4724) <= not((layer0_outputs(6722)) or (layer0_outputs(4167)));
    outputs(4725) <= layer0_outputs(6131);
    outputs(4726) <= layer0_outputs(12218);
    outputs(4727) <= not(layer0_outputs(9850)) or (layer0_outputs(12687));
    outputs(4728) <= (layer0_outputs(5531)) and not (layer0_outputs(2403));
    outputs(4729) <= layer0_outputs(7967);
    outputs(4730) <= layer0_outputs(5228);
    outputs(4731) <= layer0_outputs(7618);
    outputs(4732) <= not(layer0_outputs(1275));
    outputs(4733) <= (layer0_outputs(8393)) and not (layer0_outputs(12122));
    outputs(4734) <= (layer0_outputs(10568)) xor (layer0_outputs(3182));
    outputs(4735) <= not(layer0_outputs(10782)) or (layer0_outputs(6601));
    outputs(4736) <= not(layer0_outputs(2970)) or (layer0_outputs(2660));
    outputs(4737) <= not((layer0_outputs(7127)) and (layer0_outputs(164)));
    outputs(4738) <= layer0_outputs(12610);
    outputs(4739) <= not(layer0_outputs(5666)) or (layer0_outputs(8010));
    outputs(4740) <= layer0_outputs(106);
    outputs(4741) <= layer0_outputs(2556);
    outputs(4742) <= (layer0_outputs(12363)) or (layer0_outputs(2736));
    outputs(4743) <= not(layer0_outputs(4621));
    outputs(4744) <= not(layer0_outputs(2085)) or (layer0_outputs(5623));
    outputs(4745) <= not(layer0_outputs(377));
    outputs(4746) <= (layer0_outputs(7329)) or (layer0_outputs(3937));
    outputs(4747) <= (layer0_outputs(7453)) xor (layer0_outputs(12661));
    outputs(4748) <= not(layer0_outputs(6272)) or (layer0_outputs(9053));
    outputs(4749) <= not((layer0_outputs(6886)) and (layer0_outputs(5746)));
    outputs(4750) <= not(layer0_outputs(3990));
    outputs(4751) <= not((layer0_outputs(6456)) xor (layer0_outputs(2497)));
    outputs(4752) <= (layer0_outputs(10302)) xor (layer0_outputs(6025));
    outputs(4753) <= (layer0_outputs(12570)) and not (layer0_outputs(12655));
    outputs(4754) <= (layer0_outputs(11718)) and (layer0_outputs(8563));
    outputs(4755) <= not((layer0_outputs(10113)) or (layer0_outputs(2344)));
    outputs(4756) <= layer0_outputs(1994);
    outputs(4757) <= not((layer0_outputs(2303)) xor (layer0_outputs(4204)));
    outputs(4758) <= not(layer0_outputs(4926)) or (layer0_outputs(9856));
    outputs(4759) <= (layer0_outputs(9651)) and (layer0_outputs(2271));
    outputs(4760) <= not(layer0_outputs(9641));
    outputs(4761) <= not(layer0_outputs(7871));
    outputs(4762) <= not((layer0_outputs(2245)) xor (layer0_outputs(2405)));
    outputs(4763) <= not((layer0_outputs(6663)) and (layer0_outputs(8690)));
    outputs(4764) <= not((layer0_outputs(3904)) or (layer0_outputs(6860)));
    outputs(4765) <= not((layer0_outputs(7303)) xor (layer0_outputs(10518)));
    outputs(4766) <= not(layer0_outputs(7387));
    outputs(4767) <= not((layer0_outputs(10710)) xor (layer0_outputs(2816)));
    outputs(4768) <= layer0_outputs(4482);
    outputs(4769) <= not((layer0_outputs(837)) xor (layer0_outputs(1785)));
    outputs(4770) <= layer0_outputs(3035);
    outputs(4771) <= not(layer0_outputs(11031));
    outputs(4772) <= not((layer0_outputs(5541)) xor (layer0_outputs(5829)));
    outputs(4773) <= not(layer0_outputs(954)) or (layer0_outputs(6985));
    outputs(4774) <= (layer0_outputs(11790)) or (layer0_outputs(11535));
    outputs(4775) <= '1';
    outputs(4776) <= not(layer0_outputs(4899)) or (layer0_outputs(418));
    outputs(4777) <= not((layer0_outputs(11558)) and (layer0_outputs(9804)));
    outputs(4778) <= layer0_outputs(4011);
    outputs(4779) <= layer0_outputs(6959);
    outputs(4780) <= not(layer0_outputs(3973)) or (layer0_outputs(5584));
    outputs(4781) <= not((layer0_outputs(9786)) xor (layer0_outputs(2883)));
    outputs(4782) <= (layer0_outputs(5754)) xor (layer0_outputs(12487));
    outputs(4783) <= not((layer0_outputs(8817)) xor (layer0_outputs(5062)));
    outputs(4784) <= not(layer0_outputs(9711)) or (layer0_outputs(4036));
    outputs(4785) <= layer0_outputs(3263);
    outputs(4786) <= not(layer0_outputs(12504));
    outputs(4787) <= (layer0_outputs(2374)) xor (layer0_outputs(2291));
    outputs(4788) <= layer0_outputs(2549);
    outputs(4789) <= not(layer0_outputs(9196));
    outputs(4790) <= layer0_outputs(11661);
    outputs(4791) <= layer0_outputs(449);
    outputs(4792) <= not((layer0_outputs(7217)) xor (layer0_outputs(2006)));
    outputs(4793) <= (layer0_outputs(5590)) or (layer0_outputs(9989));
    outputs(4794) <= (layer0_outputs(7786)) xor (layer0_outputs(760));
    outputs(4795) <= (layer0_outputs(10990)) xor (layer0_outputs(5569));
    outputs(4796) <= not(layer0_outputs(11474)) or (layer0_outputs(213));
    outputs(4797) <= not((layer0_outputs(1007)) and (layer0_outputs(631)));
    outputs(4798) <= not((layer0_outputs(12005)) or (layer0_outputs(4282)));
    outputs(4799) <= layer0_outputs(1168);
    outputs(4800) <= (layer0_outputs(1521)) xor (layer0_outputs(3664));
    outputs(4801) <= not((layer0_outputs(4141)) xor (layer0_outputs(4958)));
    outputs(4802) <= layer0_outputs(11538);
    outputs(4803) <= not((layer0_outputs(9876)) xor (layer0_outputs(4166)));
    outputs(4804) <= (layer0_outputs(12323)) or (layer0_outputs(3204));
    outputs(4805) <= (layer0_outputs(843)) xor (layer0_outputs(4410));
    outputs(4806) <= layer0_outputs(996);
    outputs(4807) <= (layer0_outputs(10914)) and (layer0_outputs(3986));
    outputs(4808) <= (layer0_outputs(10427)) xor (layer0_outputs(5109));
    outputs(4809) <= (layer0_outputs(10308)) or (layer0_outputs(4241));
    outputs(4810) <= layer0_outputs(3462);
    outputs(4811) <= not((layer0_outputs(11278)) xor (layer0_outputs(5080)));
    outputs(4812) <= layer0_outputs(5417);
    outputs(4813) <= not((layer0_outputs(36)) xor (layer0_outputs(12521)));
    outputs(4814) <= layer0_outputs(12367);
    outputs(4815) <= layer0_outputs(318);
    outputs(4816) <= layer0_outputs(11859);
    outputs(4817) <= (layer0_outputs(8668)) xor (layer0_outputs(3908));
    outputs(4818) <= not(layer0_outputs(399));
    outputs(4819) <= (layer0_outputs(1287)) and not (layer0_outputs(7869));
    outputs(4820) <= (layer0_outputs(3898)) xor (layer0_outputs(11576));
    outputs(4821) <= layer0_outputs(9971);
    outputs(4822) <= layer0_outputs(10133);
    outputs(4823) <= not((layer0_outputs(2219)) xor (layer0_outputs(10784)));
    outputs(4824) <= not(layer0_outputs(4478));
    outputs(4825) <= (layer0_outputs(6205)) xor (layer0_outputs(12309));
    outputs(4826) <= not(layer0_outputs(3147));
    outputs(4827) <= not((layer0_outputs(9345)) xor (layer0_outputs(11679)));
    outputs(4828) <= not((layer0_outputs(11746)) xor (layer0_outputs(10725)));
    outputs(4829) <= not((layer0_outputs(7799)) xor (layer0_outputs(5961)));
    outputs(4830) <= not((layer0_outputs(12477)) and (layer0_outputs(10814)));
    outputs(4831) <= layer0_outputs(9117);
    outputs(4832) <= layer0_outputs(8734);
    outputs(4833) <= not((layer0_outputs(9491)) or (layer0_outputs(4413)));
    outputs(4834) <= not(layer0_outputs(323)) or (layer0_outputs(4657));
    outputs(4835) <= not(layer0_outputs(12532)) or (layer0_outputs(4465));
    outputs(4836) <= not(layer0_outputs(8050));
    outputs(4837) <= not(layer0_outputs(5727));
    outputs(4838) <= not((layer0_outputs(7868)) and (layer0_outputs(8141)));
    outputs(4839) <= not((layer0_outputs(5277)) xor (layer0_outputs(3179)));
    outputs(4840) <= (layer0_outputs(11009)) xor (layer0_outputs(7863));
    outputs(4841) <= not(layer0_outputs(4782));
    outputs(4842) <= not((layer0_outputs(8376)) and (layer0_outputs(5594)));
    outputs(4843) <= (layer0_outputs(9688)) xor (layer0_outputs(9860));
    outputs(4844) <= not((layer0_outputs(12534)) or (layer0_outputs(2491)));
    outputs(4845) <= not(layer0_outputs(11437));
    outputs(4846) <= (layer0_outputs(1287)) and not (layer0_outputs(2115));
    outputs(4847) <= '1';
    outputs(4848) <= not((layer0_outputs(1778)) or (layer0_outputs(1220)));
    outputs(4849) <= (layer0_outputs(8386)) and not (layer0_outputs(8773));
    outputs(4850) <= not(layer0_outputs(12122));
    outputs(4851) <= layer0_outputs(7187);
    outputs(4852) <= (layer0_outputs(10708)) xor (layer0_outputs(10859));
    outputs(4853) <= layer0_outputs(537);
    outputs(4854) <= not((layer0_outputs(3299)) or (layer0_outputs(7754)));
    outputs(4855) <= (layer0_outputs(714)) xor (layer0_outputs(2894));
    outputs(4856) <= layer0_outputs(2680);
    outputs(4857) <= (layer0_outputs(10616)) and not (layer0_outputs(5555));
    outputs(4858) <= not((layer0_outputs(10745)) and (layer0_outputs(2607)));
    outputs(4859) <= (layer0_outputs(3834)) xor (layer0_outputs(7975));
    outputs(4860) <= layer0_outputs(2995);
    outputs(4861) <= not((layer0_outputs(1376)) xor (layer0_outputs(10438)));
    outputs(4862) <= '0';
    outputs(4863) <= (layer0_outputs(4175)) xor (layer0_outputs(1023));
    outputs(4864) <= not((layer0_outputs(8565)) xor (layer0_outputs(11613)));
    outputs(4865) <= not(layer0_outputs(4309));
    outputs(4866) <= not((layer0_outputs(2865)) and (layer0_outputs(10674)));
    outputs(4867) <= (layer0_outputs(2300)) and not (layer0_outputs(2646));
    outputs(4868) <= not(layer0_outputs(11527));
    outputs(4869) <= not(layer0_outputs(5718)) or (layer0_outputs(994));
    outputs(4870) <= not(layer0_outputs(7229));
    outputs(4871) <= not((layer0_outputs(11402)) and (layer0_outputs(6443)));
    outputs(4872) <= not((layer0_outputs(3135)) and (layer0_outputs(11500)));
    outputs(4873) <= not((layer0_outputs(7418)) xor (layer0_outputs(12021)));
    outputs(4874) <= (layer0_outputs(10611)) xor (layer0_outputs(8759));
    outputs(4875) <= not(layer0_outputs(2099));
    outputs(4876) <= not((layer0_outputs(7100)) and (layer0_outputs(2007)));
    outputs(4877) <= not((layer0_outputs(4375)) and (layer0_outputs(10452)));
    outputs(4878) <= not(layer0_outputs(8134));
    outputs(4879) <= not((layer0_outputs(6332)) and (layer0_outputs(7954)));
    outputs(4880) <= not((layer0_outputs(2782)) xor (layer0_outputs(7667)));
    outputs(4881) <= (layer0_outputs(8146)) and not (layer0_outputs(207));
    outputs(4882) <= layer0_outputs(2655);
    outputs(4883) <= layer0_outputs(10580);
    outputs(4884) <= not(layer0_outputs(9779));
    outputs(4885) <= not(layer0_outputs(8591));
    outputs(4886) <= (layer0_outputs(1209)) xor (layer0_outputs(2286));
    outputs(4887) <= layer0_outputs(6437);
    outputs(4888) <= not((layer0_outputs(2999)) xor (layer0_outputs(2786)));
    outputs(4889) <= not((layer0_outputs(7524)) xor (layer0_outputs(12421)));
    outputs(4890) <= not((layer0_outputs(2478)) and (layer0_outputs(12673)));
    outputs(4891) <= layer0_outputs(11390);
    outputs(4892) <= not(layer0_outputs(565)) or (layer0_outputs(36));
    outputs(4893) <= not(layer0_outputs(6062)) or (layer0_outputs(2511));
    outputs(4894) <= layer0_outputs(630);
    outputs(4895) <= layer0_outputs(1203);
    outputs(4896) <= layer0_outputs(7582);
    outputs(4897) <= not((layer0_outputs(8324)) and (layer0_outputs(4452)));
    outputs(4898) <= layer0_outputs(1239);
    outputs(4899) <= (layer0_outputs(6001)) or (layer0_outputs(8651));
    outputs(4900) <= layer0_outputs(2594);
    outputs(4901) <= layer0_outputs(8506);
    outputs(4902) <= (layer0_outputs(9563)) xor (layer0_outputs(1052));
    outputs(4903) <= not((layer0_outputs(10106)) xor (layer0_outputs(5757)));
    outputs(4904) <= not((layer0_outputs(4373)) xor (layer0_outputs(3538)));
    outputs(4905) <= not(layer0_outputs(2639));
    outputs(4906) <= (layer0_outputs(272)) and not (layer0_outputs(990));
    outputs(4907) <= not(layer0_outputs(5386));
    outputs(4908) <= (layer0_outputs(10223)) and (layer0_outputs(12532));
    outputs(4909) <= layer0_outputs(1347);
    outputs(4910) <= not((layer0_outputs(1275)) and (layer0_outputs(8286)));
    outputs(4911) <= not(layer0_outputs(8130)) or (layer0_outputs(845));
    outputs(4912) <= layer0_outputs(8437);
    outputs(4913) <= not(layer0_outputs(1210)) or (layer0_outputs(2330));
    outputs(4914) <= not(layer0_outputs(6116)) or (layer0_outputs(6944));
    outputs(4915) <= layer0_outputs(8389);
    outputs(4916) <= (layer0_outputs(296)) and not (layer0_outputs(4036));
    outputs(4917) <= not(layer0_outputs(1007));
    outputs(4918) <= (layer0_outputs(229)) xor (layer0_outputs(1523));
    outputs(4919) <= not((layer0_outputs(5872)) and (layer0_outputs(6160)));
    outputs(4920) <= (layer0_outputs(3819)) or (layer0_outputs(7406));
    outputs(4921) <= not((layer0_outputs(6194)) xor (layer0_outputs(6771)));
    outputs(4922) <= (layer0_outputs(11775)) xor (layer0_outputs(6118));
    outputs(4923) <= not((layer0_outputs(2043)) and (layer0_outputs(10904)));
    outputs(4924) <= (layer0_outputs(3402)) or (layer0_outputs(4434));
    outputs(4925) <= layer0_outputs(6574);
    outputs(4926) <= not(layer0_outputs(9623));
    outputs(4927) <= not(layer0_outputs(10440));
    outputs(4928) <= (layer0_outputs(10809)) or (layer0_outputs(12446));
    outputs(4929) <= (layer0_outputs(2877)) xor (layer0_outputs(10279));
    outputs(4930) <= layer0_outputs(7986);
    outputs(4931) <= not((layer0_outputs(8991)) and (layer0_outputs(5810)));
    outputs(4932) <= (layer0_outputs(9553)) or (layer0_outputs(1811));
    outputs(4933) <= not(layer0_outputs(9083));
    outputs(4934) <= not((layer0_outputs(198)) or (layer0_outputs(165)));
    outputs(4935) <= (layer0_outputs(8461)) xor (layer0_outputs(256));
    outputs(4936) <= not((layer0_outputs(6831)) xor (layer0_outputs(5434)));
    outputs(4937) <= not(layer0_outputs(3952));
    outputs(4938) <= (layer0_outputs(8109)) and not (layer0_outputs(4896));
    outputs(4939) <= not((layer0_outputs(3043)) or (layer0_outputs(1960)));
    outputs(4940) <= not(layer0_outputs(11727)) or (layer0_outputs(9740));
    outputs(4941) <= not(layer0_outputs(1738)) or (layer0_outputs(7043));
    outputs(4942) <= layer0_outputs(11110);
    outputs(4943) <= not(layer0_outputs(6033));
    outputs(4944) <= (layer0_outputs(8734)) xor (layer0_outputs(5947));
    outputs(4945) <= layer0_outputs(6334);
    outputs(4946) <= (layer0_outputs(3341)) xor (layer0_outputs(2702));
    outputs(4947) <= layer0_outputs(591);
    outputs(4948) <= not(layer0_outputs(10122));
    outputs(4949) <= layer0_outputs(2834);
    outputs(4950) <= not(layer0_outputs(3189));
    outputs(4951) <= not((layer0_outputs(10720)) xor (layer0_outputs(4689)));
    outputs(4952) <= (layer0_outputs(10340)) xor (layer0_outputs(1927));
    outputs(4953) <= layer0_outputs(8658);
    outputs(4954) <= not(layer0_outputs(9903));
    outputs(4955) <= layer0_outputs(854);
    outputs(4956) <= (layer0_outputs(11758)) and (layer0_outputs(7201));
    outputs(4957) <= not(layer0_outputs(7525));
    outputs(4958) <= (layer0_outputs(3032)) and not (layer0_outputs(8281));
    outputs(4959) <= (layer0_outputs(9791)) xor (layer0_outputs(8670));
    outputs(4960) <= not(layer0_outputs(9164)) or (layer0_outputs(4327));
    outputs(4961) <= not(layer0_outputs(11044));
    outputs(4962) <= not((layer0_outputs(5831)) xor (layer0_outputs(6001)));
    outputs(4963) <= layer0_outputs(5665);
    outputs(4964) <= layer0_outputs(7443);
    outputs(4965) <= (layer0_outputs(9464)) or (layer0_outputs(10230));
    outputs(4966) <= layer0_outputs(6876);
    outputs(4967) <= (layer0_outputs(12791)) or (layer0_outputs(8445));
    outputs(4968) <= (layer0_outputs(9291)) and not (layer0_outputs(2111));
    outputs(4969) <= (layer0_outputs(4608)) xor (layer0_outputs(6781));
    outputs(4970) <= (layer0_outputs(2854)) or (layer0_outputs(9062));
    outputs(4971) <= layer0_outputs(8675);
    outputs(4972) <= not(layer0_outputs(7082));
    outputs(4973) <= not((layer0_outputs(6777)) and (layer0_outputs(4851)));
    outputs(4974) <= (layer0_outputs(2368)) xor (layer0_outputs(10069));
    outputs(4975) <= not(layer0_outputs(5));
    outputs(4976) <= (layer0_outputs(5711)) and not (layer0_outputs(4914));
    outputs(4977) <= layer0_outputs(5015);
    outputs(4978) <= not(layer0_outputs(4752));
    outputs(4979) <= not(layer0_outputs(12324));
    outputs(4980) <= (layer0_outputs(5863)) and (layer0_outputs(12488));
    outputs(4981) <= not(layer0_outputs(6873));
    outputs(4982) <= not(layer0_outputs(9138));
    outputs(4983) <= (layer0_outputs(7095)) xor (layer0_outputs(9070));
    outputs(4984) <= (layer0_outputs(9614)) and not (layer0_outputs(2807));
    outputs(4985) <= not((layer0_outputs(11304)) and (layer0_outputs(2174)));
    outputs(4986) <= layer0_outputs(4383);
    outputs(4987) <= layer0_outputs(5244);
    outputs(4988) <= (layer0_outputs(2520)) xor (layer0_outputs(5833));
    outputs(4989) <= not(layer0_outputs(8132));
    outputs(4990) <= not((layer0_outputs(3141)) and (layer0_outputs(7453)));
    outputs(4991) <= (layer0_outputs(11404)) or (layer0_outputs(2621));
    outputs(4992) <= (layer0_outputs(12780)) xor (layer0_outputs(12228));
    outputs(4993) <= (layer0_outputs(10483)) xor (layer0_outputs(10656));
    outputs(4994) <= not(layer0_outputs(10497));
    outputs(4995) <= not((layer0_outputs(6775)) or (layer0_outputs(751)));
    outputs(4996) <= not((layer0_outputs(10262)) xor (layer0_outputs(9161)));
    outputs(4997) <= layer0_outputs(10359);
    outputs(4998) <= layer0_outputs(3226);
    outputs(4999) <= not((layer0_outputs(12320)) xor (layer0_outputs(11405)));
    outputs(5000) <= not((layer0_outputs(9566)) and (layer0_outputs(9337)));
    outputs(5001) <= not((layer0_outputs(5642)) xor (layer0_outputs(1648)));
    outputs(5002) <= not((layer0_outputs(10967)) or (layer0_outputs(5635)));
    outputs(5003) <= not(layer0_outputs(4852));
    outputs(5004) <= not((layer0_outputs(10207)) xor (layer0_outputs(3809)));
    outputs(5005) <= not((layer0_outputs(6549)) and (layer0_outputs(10791)));
    outputs(5006) <= not(layer0_outputs(6856));
    outputs(5007) <= not(layer0_outputs(5082));
    outputs(5008) <= (layer0_outputs(6722)) or (layer0_outputs(7957));
    outputs(5009) <= (layer0_outputs(3526)) and not (layer0_outputs(1640));
    outputs(5010) <= not((layer0_outputs(6241)) xor (layer0_outputs(4269)));
    outputs(5011) <= (layer0_outputs(10870)) and (layer0_outputs(5595));
    outputs(5012) <= layer0_outputs(11399);
    outputs(5013) <= layer0_outputs(8298);
    outputs(5014) <= not(layer0_outputs(4327));
    outputs(5015) <= not(layer0_outputs(634));
    outputs(5016) <= not((layer0_outputs(11571)) xor (layer0_outputs(11615)));
    outputs(5017) <= (layer0_outputs(6749)) and not (layer0_outputs(5176));
    outputs(5018) <= layer0_outputs(11648);
    outputs(5019) <= (layer0_outputs(600)) xor (layer0_outputs(8348));
    outputs(5020) <= (layer0_outputs(7402)) xor (layer0_outputs(551));
    outputs(5021) <= layer0_outputs(9267);
    outputs(5022) <= not(layer0_outputs(3998));
    outputs(5023) <= not((layer0_outputs(12330)) xor (layer0_outputs(10642)));
    outputs(5024) <= (layer0_outputs(8178)) or (layer0_outputs(5049));
    outputs(5025) <= not(layer0_outputs(12336));
    outputs(5026) <= '1';
    outputs(5027) <= (layer0_outputs(8239)) xor (layer0_outputs(7384));
    outputs(5028) <= not(layer0_outputs(477));
    outputs(5029) <= not(layer0_outputs(1311));
    outputs(5030) <= (layer0_outputs(5369)) or (layer0_outputs(10231));
    outputs(5031) <= not((layer0_outputs(1182)) xor (layer0_outputs(9245)));
    outputs(5032) <= not((layer0_outputs(10767)) and (layer0_outputs(10787)));
    outputs(5033) <= not(layer0_outputs(10290));
    outputs(5034) <= not((layer0_outputs(4022)) xor (layer0_outputs(3298)));
    outputs(5035) <= not(layer0_outputs(7822));
    outputs(5036) <= not((layer0_outputs(3452)) and (layer0_outputs(6745)));
    outputs(5037) <= not((layer0_outputs(8457)) xor (layer0_outputs(3810)));
    outputs(5038) <= not(layer0_outputs(4801));
    outputs(5039) <= layer0_outputs(3051);
    outputs(5040) <= (layer0_outputs(10406)) and not (layer0_outputs(8330));
    outputs(5041) <= layer0_outputs(12076);
    outputs(5042) <= not(layer0_outputs(10569)) or (layer0_outputs(2778));
    outputs(5043) <= not(layer0_outputs(12206));
    outputs(5044) <= not(layer0_outputs(7425));
    outputs(5045) <= not((layer0_outputs(500)) and (layer0_outputs(7452)));
    outputs(5046) <= not(layer0_outputs(6248)) or (layer0_outputs(11377));
    outputs(5047) <= not(layer0_outputs(982));
    outputs(5048) <= not((layer0_outputs(1343)) xor (layer0_outputs(1230)));
    outputs(5049) <= not(layer0_outputs(7374));
    outputs(5050) <= not(layer0_outputs(12708));
    outputs(5051) <= layer0_outputs(7677);
    outputs(5052) <= not(layer0_outputs(7846));
    outputs(5053) <= not(layer0_outputs(5377));
    outputs(5054) <= not(layer0_outputs(8353)) or (layer0_outputs(239));
    outputs(5055) <= not((layer0_outputs(8092)) xor (layer0_outputs(1175)));
    outputs(5056) <= layer0_outputs(9871);
    outputs(5057) <= (layer0_outputs(9582)) and (layer0_outputs(7565));
    outputs(5058) <= layer0_outputs(11714);
    outputs(5059) <= not(layer0_outputs(1525));
    outputs(5060) <= not((layer0_outputs(5709)) and (layer0_outputs(1663)));
    outputs(5061) <= (layer0_outputs(6358)) xor (layer0_outputs(241));
    outputs(5062) <= not(layer0_outputs(2464));
    outputs(5063) <= layer0_outputs(2932);
    outputs(5064) <= not((layer0_outputs(5167)) and (layer0_outputs(5770)));
    outputs(5065) <= layer0_outputs(7320);
    outputs(5066) <= (layer0_outputs(9961)) xor (layer0_outputs(3345));
    outputs(5067) <= not(layer0_outputs(7862));
    outputs(5068) <= layer0_outputs(12387);
    outputs(5069) <= layer0_outputs(5128);
    outputs(5070) <= not((layer0_outputs(4554)) and (layer0_outputs(11504)));
    outputs(5071) <= layer0_outputs(1797);
    outputs(5072) <= (layer0_outputs(6856)) xor (layer0_outputs(3331));
    outputs(5073) <= (layer0_outputs(7316)) and (layer0_outputs(4839));
    outputs(5074) <= not(layer0_outputs(5661)) or (layer0_outputs(5463));
    outputs(5075) <= not(layer0_outputs(1743)) or (layer0_outputs(6284));
    outputs(5076) <= (layer0_outputs(7350)) and not (layer0_outputs(6380));
    outputs(5077) <= not(layer0_outputs(2070)) or (layer0_outputs(1230));
    outputs(5078) <= (layer0_outputs(2565)) xor (layer0_outputs(2686));
    outputs(5079) <= (layer0_outputs(1799)) and (layer0_outputs(6271));
    outputs(5080) <= not(layer0_outputs(4401)) or (layer0_outputs(11836));
    outputs(5081) <= layer0_outputs(8860);
    outputs(5082) <= not((layer0_outputs(5918)) xor (layer0_outputs(230)));
    outputs(5083) <= not(layer0_outputs(9714));
    outputs(5084) <= not(layer0_outputs(5515));
    outputs(5085) <= not((layer0_outputs(6118)) xor (layer0_outputs(1969)));
    outputs(5086) <= not(layer0_outputs(1682));
    outputs(5087) <= (layer0_outputs(10552)) xor (layer0_outputs(431));
    outputs(5088) <= not((layer0_outputs(12386)) and (layer0_outputs(12292)));
    outputs(5089) <= (layer0_outputs(9291)) and not (layer0_outputs(2910));
    outputs(5090) <= layer0_outputs(10382);
    outputs(5091) <= not(layer0_outputs(8571)) or (layer0_outputs(9071));
    outputs(5092) <= (layer0_outputs(3420)) xor (layer0_outputs(5612));
    outputs(5093) <= (layer0_outputs(10083)) and not (layer0_outputs(10528));
    outputs(5094) <= (layer0_outputs(9036)) xor (layer0_outputs(6640));
    outputs(5095) <= not(layer0_outputs(12654));
    outputs(5096) <= not((layer0_outputs(10543)) and (layer0_outputs(4915)));
    outputs(5097) <= not((layer0_outputs(3199)) or (layer0_outputs(11367)));
    outputs(5098) <= not((layer0_outputs(9347)) or (layer0_outputs(1251)));
    outputs(5099) <= not((layer0_outputs(6280)) xor (layer0_outputs(3302)));
    outputs(5100) <= not(layer0_outputs(6844)) or (layer0_outputs(6867));
    outputs(5101) <= not(layer0_outputs(2981));
    outputs(5102) <= (layer0_outputs(9881)) and not (layer0_outputs(2448));
    outputs(5103) <= (layer0_outputs(6315)) or (layer0_outputs(6031));
    outputs(5104) <= not((layer0_outputs(8099)) and (layer0_outputs(6979)));
    outputs(5105) <= layer0_outputs(8424);
    outputs(5106) <= not((layer0_outputs(9282)) and (layer0_outputs(8667)));
    outputs(5107) <= not((layer0_outputs(6361)) xor (layer0_outputs(341)));
    outputs(5108) <= not(layer0_outputs(5325));
    outputs(5109) <= (layer0_outputs(4430)) xor (layer0_outputs(12653));
    outputs(5110) <= layer0_outputs(5420);
    outputs(5111) <= (layer0_outputs(12482)) xor (layer0_outputs(11694));
    outputs(5112) <= not(layer0_outputs(11788));
    outputs(5113) <= not(layer0_outputs(4305));
    outputs(5114) <= not((layer0_outputs(2257)) xor (layer0_outputs(7029)));
    outputs(5115) <= not(layer0_outputs(5568));
    outputs(5116) <= layer0_outputs(6528);
    outputs(5117) <= (layer0_outputs(7370)) or (layer0_outputs(8242));
    outputs(5118) <= (layer0_outputs(3122)) and not (layer0_outputs(2946));
    outputs(5119) <= layer0_outputs(3921);
    outputs(5120) <= not(layer0_outputs(7435));
    outputs(5121) <= not((layer0_outputs(11494)) xor (layer0_outputs(4812)));
    outputs(5122) <= '0';
    outputs(5123) <= (layer0_outputs(10197)) and not (layer0_outputs(5991));
    outputs(5124) <= not((layer0_outputs(8339)) or (layer0_outputs(3105)));
    outputs(5125) <= not(layer0_outputs(3496));
    outputs(5126) <= (layer0_outputs(6303)) and not (layer0_outputs(11641));
    outputs(5127) <= not((layer0_outputs(11128)) and (layer0_outputs(8901)));
    outputs(5128) <= not((layer0_outputs(11923)) or (layer0_outputs(4822)));
    outputs(5129) <= not(layer0_outputs(12264));
    outputs(5130) <= not((layer0_outputs(2326)) xor (layer0_outputs(2501)));
    outputs(5131) <= (layer0_outputs(1904)) and not (layer0_outputs(8127));
    outputs(5132) <= not(layer0_outputs(6412)) or (layer0_outputs(5313));
    outputs(5133) <= (layer0_outputs(7314)) xor (layer0_outputs(9973));
    outputs(5134) <= not(layer0_outputs(4382));
    outputs(5135) <= layer0_outputs(7865);
    outputs(5136) <= not((layer0_outputs(4925)) xor (layer0_outputs(5337)));
    outputs(5137) <= not(layer0_outputs(6683)) or (layer0_outputs(5030));
    outputs(5138) <= layer0_outputs(3471);
    outputs(5139) <= layer0_outputs(4394);
    outputs(5140) <= (layer0_outputs(4343)) xor (layer0_outputs(9030));
    outputs(5141) <= not((layer0_outputs(6757)) xor (layer0_outputs(1459)));
    outputs(5142) <= layer0_outputs(4296);
    outputs(5143) <= (layer0_outputs(6257)) xor (layer0_outputs(12522));
    outputs(5144) <= not((layer0_outputs(6761)) xor (layer0_outputs(9821)));
    outputs(5145) <= layer0_outputs(9675);
    outputs(5146) <= not(layer0_outputs(10304));
    outputs(5147) <= not(layer0_outputs(3697));
    outputs(5148) <= (layer0_outputs(7788)) and not (layer0_outputs(10657));
    outputs(5149) <= (layer0_outputs(4891)) and not (layer0_outputs(9498));
    outputs(5150) <= not(layer0_outputs(2270));
    outputs(5151) <= (layer0_outputs(8770)) and not (layer0_outputs(6835));
    outputs(5152) <= (layer0_outputs(11038)) and not (layer0_outputs(5981));
    outputs(5153) <= (layer0_outputs(5728)) and not (layer0_outputs(123));
    outputs(5154) <= not(layer0_outputs(5502)) or (layer0_outputs(3755));
    outputs(5155) <= (layer0_outputs(1335)) and not (layer0_outputs(5318));
    outputs(5156) <= not(layer0_outputs(9640));
    outputs(5157) <= (layer0_outputs(12592)) and not (layer0_outputs(9982));
    outputs(5158) <= layer0_outputs(4993);
    outputs(5159) <= (layer0_outputs(8232)) xor (layer0_outputs(8730));
    outputs(5160) <= not(layer0_outputs(11548));
    outputs(5161) <= not(layer0_outputs(5775));
    outputs(5162) <= not((layer0_outputs(2151)) xor (layer0_outputs(7852)));
    outputs(5163) <= (layer0_outputs(3464)) and not (layer0_outputs(7298));
    outputs(5164) <= not(layer0_outputs(3991));
    outputs(5165) <= (layer0_outputs(6039)) xor (layer0_outputs(1575));
    outputs(5166) <= not((layer0_outputs(10546)) xor (layer0_outputs(4676)));
    outputs(5167) <= not(layer0_outputs(11434));
    outputs(5168) <= not(layer0_outputs(379));
    outputs(5169) <= not(layer0_outputs(4880));
    outputs(5170) <= not(layer0_outputs(6597));
    outputs(5171) <= not(layer0_outputs(3870));
    outputs(5172) <= (layer0_outputs(10392)) and not (layer0_outputs(1046));
    outputs(5173) <= (layer0_outputs(8163)) and (layer0_outputs(403));
    outputs(5174) <= layer0_outputs(12240);
    outputs(5175) <= (layer0_outputs(1150)) and not (layer0_outputs(7324));
    outputs(5176) <= '0';
    outputs(5177) <= (layer0_outputs(11342)) and not (layer0_outputs(11040));
    outputs(5178) <= (layer0_outputs(8920)) and not (layer0_outputs(6470));
    outputs(5179) <= (layer0_outputs(8572)) and not (layer0_outputs(2840));
    outputs(5180) <= layer0_outputs(2031);
    outputs(5181) <= layer0_outputs(2646);
    outputs(5182) <= not(layer0_outputs(1076));
    outputs(5183) <= (layer0_outputs(6966)) and (layer0_outputs(5945));
    outputs(5184) <= not((layer0_outputs(5659)) xor (layer0_outputs(9547)));
    outputs(5185) <= (layer0_outputs(4902)) and not (layer0_outputs(5459));
    outputs(5186) <= (layer0_outputs(7856)) xor (layer0_outputs(6866));
    outputs(5187) <= not(layer0_outputs(9511));
    outputs(5188) <= not((layer0_outputs(7987)) xor (layer0_outputs(8000)));
    outputs(5189) <= (layer0_outputs(3727)) xor (layer0_outputs(4011));
    outputs(5190) <= layer0_outputs(5993);
    outputs(5191) <= '0';
    outputs(5192) <= not((layer0_outputs(7262)) xor (layer0_outputs(4093)));
    outputs(5193) <= not((layer0_outputs(6988)) xor (layer0_outputs(3349)));
    outputs(5194) <= not((layer0_outputs(8624)) or (layer0_outputs(937)));
    outputs(5195) <= not((layer0_outputs(10370)) xor (layer0_outputs(7749)));
    outputs(5196) <= (layer0_outputs(177)) and (layer0_outputs(11428));
    outputs(5197) <= not((layer0_outputs(6416)) xor (layer0_outputs(10822)));
    outputs(5198) <= layer0_outputs(1667);
    outputs(5199) <= not((layer0_outputs(2025)) xor (layer0_outputs(5314)));
    outputs(5200) <= (layer0_outputs(6995)) and not (layer0_outputs(7425));
    outputs(5201) <= layer0_outputs(3896);
    outputs(5202) <= (layer0_outputs(7767)) xor (layer0_outputs(5115));
    outputs(5203) <= not(layer0_outputs(11354));
    outputs(5204) <= not(layer0_outputs(7606));
    outputs(5205) <= (layer0_outputs(8689)) or (layer0_outputs(6821));
    outputs(5206) <= not((layer0_outputs(3926)) or (layer0_outputs(10064)));
    outputs(5207) <= not((layer0_outputs(3678)) or (layer0_outputs(8196)));
    outputs(5208) <= layer0_outputs(6324);
    outputs(5209) <= (layer0_outputs(6494)) and (layer0_outputs(8825));
    outputs(5210) <= not((layer0_outputs(9530)) xor (layer0_outputs(7114)));
    outputs(5211) <= (layer0_outputs(2127)) xor (layer0_outputs(9241));
    outputs(5212) <= not(layer0_outputs(10075));
    outputs(5213) <= '0';
    outputs(5214) <= not(layer0_outputs(12675));
    outputs(5215) <= (layer0_outputs(9630)) and (layer0_outputs(2001));
    outputs(5216) <= not((layer0_outputs(7383)) xor (layer0_outputs(7067)));
    outputs(5217) <= not(layer0_outputs(4048));
    outputs(5218) <= not(layer0_outputs(5510)) or (layer0_outputs(5555));
    outputs(5219) <= (layer0_outputs(8353)) and not (layer0_outputs(419));
    outputs(5220) <= layer0_outputs(8804);
    outputs(5221) <= layer0_outputs(7628);
    outputs(5222) <= not((layer0_outputs(4035)) or (layer0_outputs(756)));
    outputs(5223) <= not(layer0_outputs(2279)) or (layer0_outputs(2757));
    outputs(5224) <= not((layer0_outputs(5862)) xor (layer0_outputs(8944)));
    outputs(5225) <= layer0_outputs(826);
    outputs(5226) <= (layer0_outputs(7429)) and not (layer0_outputs(5667));
    outputs(5227) <= not((layer0_outputs(5329)) xor (layer0_outputs(12613)));
    outputs(5228) <= (layer0_outputs(5645)) and (layer0_outputs(4387));
    outputs(5229) <= not((layer0_outputs(2045)) xor (layer0_outputs(4918)));
    outputs(5230) <= not((layer0_outputs(7277)) xor (layer0_outputs(8898)));
    outputs(5231) <= layer0_outputs(4103);
    outputs(5232) <= not((layer0_outputs(8988)) xor (layer0_outputs(1874)));
    outputs(5233) <= (layer0_outputs(3617)) and not (layer0_outputs(6591));
    outputs(5234) <= not((layer0_outputs(10851)) xor (layer0_outputs(6627)));
    outputs(5235) <= not((layer0_outputs(951)) xor (layer0_outputs(8207)));
    outputs(5236) <= not(layer0_outputs(135));
    outputs(5237) <= not((layer0_outputs(262)) xor (layer0_outputs(8663)));
    outputs(5238) <= layer0_outputs(12498);
    outputs(5239) <= layer0_outputs(876);
    outputs(5240) <= (layer0_outputs(3214)) and not (layer0_outputs(9226));
    outputs(5241) <= layer0_outputs(3339);
    outputs(5242) <= not(layer0_outputs(1936));
    outputs(5243) <= not(layer0_outputs(1925));
    outputs(5244) <= not(layer0_outputs(3978));
    outputs(5245) <= not((layer0_outputs(1713)) xor (layer0_outputs(6257)));
    outputs(5246) <= (layer0_outputs(5406)) and not (layer0_outputs(3017));
    outputs(5247) <= (layer0_outputs(1726)) xor (layer0_outputs(10931));
    outputs(5248) <= (layer0_outputs(1451)) xor (layer0_outputs(9286));
    outputs(5249) <= (layer0_outputs(6401)) and not (layer0_outputs(1839));
    outputs(5250) <= not((layer0_outputs(2849)) and (layer0_outputs(1596)));
    outputs(5251) <= not((layer0_outputs(1717)) xor (layer0_outputs(3188)));
    outputs(5252) <= layer0_outputs(10903);
    outputs(5253) <= not((layer0_outputs(11124)) xor (layer0_outputs(5648)));
    outputs(5254) <= (layer0_outputs(1924)) and (layer0_outputs(1993));
    outputs(5255) <= (layer0_outputs(9377)) and not (layer0_outputs(4601));
    outputs(5256) <= '0';
    outputs(5257) <= layer0_outputs(8938);
    outputs(5258) <= (layer0_outputs(9393)) and not (layer0_outputs(7597));
    outputs(5259) <= not(layer0_outputs(12299));
    outputs(5260) <= layer0_outputs(1683);
    outputs(5261) <= layer0_outputs(6096);
    outputs(5262) <= not((layer0_outputs(4844)) xor (layer0_outputs(101)));
    outputs(5263) <= not((layer0_outputs(1421)) xor (layer0_outputs(2910)));
    outputs(5264) <= not((layer0_outputs(4017)) or (layer0_outputs(1679)));
    outputs(5265) <= layer0_outputs(11509);
    outputs(5266) <= (layer0_outputs(921)) or (layer0_outputs(3985));
    outputs(5267) <= (layer0_outputs(11454)) xor (layer0_outputs(2544));
    outputs(5268) <= (layer0_outputs(6496)) and not (layer0_outputs(1690));
    outputs(5269) <= not(layer0_outputs(12366));
    outputs(5270) <= layer0_outputs(2515);
    outputs(5271) <= (layer0_outputs(10620)) and not (layer0_outputs(1952));
    outputs(5272) <= not((layer0_outputs(9229)) xor (layer0_outputs(10516)));
    outputs(5273) <= not((layer0_outputs(5267)) xor (layer0_outputs(8604)));
    outputs(5274) <= not(layer0_outputs(8180)) or (layer0_outputs(11499));
    outputs(5275) <= not((layer0_outputs(9834)) xor (layer0_outputs(2781)));
    outputs(5276) <= not(layer0_outputs(12107));
    outputs(5277) <= not((layer0_outputs(7305)) xor (layer0_outputs(4629)));
    outputs(5278) <= layer0_outputs(9099);
    outputs(5279) <= (layer0_outputs(10429)) xor (layer0_outputs(1864));
    outputs(5280) <= not((layer0_outputs(6378)) and (layer0_outputs(458)));
    outputs(5281) <= (layer0_outputs(6363)) and (layer0_outputs(1135));
    outputs(5282) <= not(layer0_outputs(2720));
    outputs(5283) <= layer0_outputs(9778);
    outputs(5284) <= not((layer0_outputs(879)) xor (layer0_outputs(10960)));
    outputs(5285) <= not((layer0_outputs(3229)) or (layer0_outputs(4333)));
    outputs(5286) <= not((layer0_outputs(5516)) and (layer0_outputs(8824)));
    outputs(5287) <= layer0_outputs(3807);
    outputs(5288) <= not((layer0_outputs(1073)) and (layer0_outputs(5486)));
    outputs(5289) <= layer0_outputs(581);
    outputs(5290) <= not(layer0_outputs(3510)) or (layer0_outputs(11537));
    outputs(5291) <= (layer0_outputs(447)) and not (layer0_outputs(6547));
    outputs(5292) <= (layer0_outputs(2132)) and not (layer0_outputs(2514));
    outputs(5293) <= not((layer0_outputs(1054)) or (layer0_outputs(5183)));
    outputs(5294) <= (layer0_outputs(10046)) and (layer0_outputs(2462));
    outputs(5295) <= (layer0_outputs(3623)) and not (layer0_outputs(10141));
    outputs(5296) <= (layer0_outputs(8595)) and (layer0_outputs(7420));
    outputs(5297) <= (layer0_outputs(4013)) xor (layer0_outputs(7587));
    outputs(5298) <= (layer0_outputs(9713)) xor (layer0_outputs(3827));
    outputs(5299) <= layer0_outputs(5969);
    outputs(5300) <= not((layer0_outputs(8895)) xor (layer0_outputs(2134)));
    outputs(5301) <= not((layer0_outputs(107)) xor (layer0_outputs(1329)));
    outputs(5302) <= not(layer0_outputs(4444)) or (layer0_outputs(6023));
    outputs(5303) <= not(layer0_outputs(5275));
    outputs(5304) <= not((layer0_outputs(5318)) xor (layer0_outputs(1072)));
    outputs(5305) <= (layer0_outputs(10169)) and not (layer0_outputs(6011));
    outputs(5306) <= not(layer0_outputs(4762)) or (layer0_outputs(6329));
    outputs(5307) <= (layer0_outputs(2006)) and not (layer0_outputs(2193));
    outputs(5308) <= not((layer0_outputs(584)) or (layer0_outputs(9329)));
    outputs(5309) <= layer0_outputs(8129);
    outputs(5310) <= (layer0_outputs(9316)) and not (layer0_outputs(3288));
    outputs(5311) <= (layer0_outputs(3823)) and not (layer0_outputs(5878));
    outputs(5312) <= not(layer0_outputs(9280));
    outputs(5313) <= not(layer0_outputs(7055));
    outputs(5314) <= layer0_outputs(9724);
    outputs(5315) <= not((layer0_outputs(10538)) xor (layer0_outputs(7480)));
    outputs(5316) <= (layer0_outputs(2202)) and not (layer0_outputs(5156));
    outputs(5317) <= (layer0_outputs(1302)) and not (layer0_outputs(68));
    outputs(5318) <= (layer0_outputs(9005)) xor (layer0_outputs(3653));
    outputs(5319) <= not((layer0_outputs(8004)) xor (layer0_outputs(9359)));
    outputs(5320) <= not(layer0_outputs(12407));
    outputs(5321) <= not((layer0_outputs(3774)) or (layer0_outputs(459)));
    outputs(5322) <= (layer0_outputs(11059)) and (layer0_outputs(1117));
    outputs(5323) <= (layer0_outputs(11860)) or (layer0_outputs(3014));
    outputs(5324) <= not(layer0_outputs(11168));
    outputs(5325) <= not(layer0_outputs(1426));
    outputs(5326) <= (layer0_outputs(10233)) and not (layer0_outputs(9900));
    outputs(5327) <= (layer0_outputs(5687)) xor (layer0_outputs(9677));
    outputs(5328) <= not(layer0_outputs(8892));
    outputs(5329) <= not((layer0_outputs(11318)) or (layer0_outputs(2433)));
    outputs(5330) <= not((layer0_outputs(6357)) xor (layer0_outputs(12150)));
    outputs(5331) <= layer0_outputs(9910);
    outputs(5332) <= not((layer0_outputs(9413)) xor (layer0_outputs(2546)));
    outputs(5333) <= not((layer0_outputs(10041)) xor (layer0_outputs(7705)));
    outputs(5334) <= (layer0_outputs(33)) and not (layer0_outputs(5928));
    outputs(5335) <= (layer0_outputs(8402)) xor (layer0_outputs(4876));
    outputs(5336) <= (layer0_outputs(3878)) xor (layer0_outputs(1366));
    outputs(5337) <= (layer0_outputs(9268)) xor (layer0_outputs(12005));
    outputs(5338) <= layer0_outputs(757);
    outputs(5339) <= (layer0_outputs(11751)) and (layer0_outputs(8606));
    outputs(5340) <= not(layer0_outputs(1844));
    outputs(5341) <= (layer0_outputs(20)) and not (layer0_outputs(12546));
    outputs(5342) <= not(layer0_outputs(5397));
    outputs(5343) <= (layer0_outputs(5405)) and (layer0_outputs(941));
    outputs(5344) <= (layer0_outputs(9739)) and not (layer0_outputs(1845));
    outputs(5345) <= not((layer0_outputs(2955)) and (layer0_outputs(519)));
    outputs(5346) <= (layer0_outputs(9031)) xor (layer0_outputs(8462));
    outputs(5347) <= (layer0_outputs(9564)) xor (layer0_outputs(1372));
    outputs(5348) <= (layer0_outputs(9864)) and not (layer0_outputs(4178));
    outputs(5349) <= layer0_outputs(6952);
    outputs(5350) <= layer0_outputs(8928);
    outputs(5351) <= not((layer0_outputs(1074)) xor (layer0_outputs(3295)));
    outputs(5352) <= not((layer0_outputs(10937)) xor (layer0_outputs(6998)));
    outputs(5353) <= (layer0_outputs(10764)) and (layer0_outputs(4796));
    outputs(5354) <= layer0_outputs(3545);
    outputs(5355) <= (layer0_outputs(4571)) and not (layer0_outputs(8758));
    outputs(5356) <= (layer0_outputs(1191)) xor (layer0_outputs(11347));
    outputs(5357) <= not(layer0_outputs(1002));
    outputs(5358) <= (layer0_outputs(1621)) xor (layer0_outputs(8828));
    outputs(5359) <= not((layer0_outputs(9205)) or (layer0_outputs(6002)));
    outputs(5360) <= layer0_outputs(2046);
    outputs(5361) <= not((layer0_outputs(217)) xor (layer0_outputs(11651)));
    outputs(5362) <= not((layer0_outputs(2643)) or (layer0_outputs(9486)));
    outputs(5363) <= (layer0_outputs(5424)) or (layer0_outputs(1278));
    outputs(5364) <= (layer0_outputs(10009)) xor (layer0_outputs(10972));
    outputs(5365) <= not((layer0_outputs(5396)) xor (layer0_outputs(9677)));
    outputs(5366) <= (layer0_outputs(8561)) and not (layer0_outputs(4219));
    outputs(5367) <= layer0_outputs(2756);
    outputs(5368) <= (layer0_outputs(2213)) and (layer0_outputs(4768));
    outputs(5369) <= (layer0_outputs(235)) and not (layer0_outputs(7900));
    outputs(5370) <= not(layer0_outputs(10870));
    outputs(5371) <= layer0_outputs(5358);
    outputs(5372) <= (layer0_outputs(5733)) and not (layer0_outputs(11320));
    outputs(5373) <= '0';
    outputs(5374) <= (layer0_outputs(11963)) and not (layer0_outputs(11694));
    outputs(5375) <= not((layer0_outputs(1214)) xor (layer0_outputs(6121)));
    outputs(5376) <= not((layer0_outputs(1928)) xor (layer0_outputs(4357)));
    outputs(5377) <= not(layer0_outputs(9395));
    outputs(5378) <= (layer0_outputs(3571)) or (layer0_outputs(11267));
    outputs(5379) <= (layer0_outputs(1715)) xor (layer0_outputs(4747));
    outputs(5380) <= not((layer0_outputs(12411)) or (layer0_outputs(3178)));
    outputs(5381) <= layer0_outputs(9565);
    outputs(5382) <= (layer0_outputs(7527)) or (layer0_outputs(6112));
    outputs(5383) <= (layer0_outputs(7341)) and not (layer0_outputs(7230));
    outputs(5384) <= (layer0_outputs(10246)) xor (layer0_outputs(9191));
    outputs(5385) <= (layer0_outputs(10515)) and (layer0_outputs(4139));
    outputs(5386) <= layer0_outputs(9544);
    outputs(5387) <= not((layer0_outputs(5073)) xor (layer0_outputs(12095)));
    outputs(5388) <= not((layer0_outputs(7312)) xor (layer0_outputs(11776)));
    outputs(5389) <= not(layer0_outputs(1394));
    outputs(5390) <= not(layer0_outputs(1412));
    outputs(5391) <= not(layer0_outputs(12171));
    outputs(5392) <= (layer0_outputs(10987)) and not (layer0_outputs(10820));
    outputs(5393) <= (layer0_outputs(4130)) xor (layer0_outputs(260));
    outputs(5394) <= not(layer0_outputs(7185));
    outputs(5395) <= not((layer0_outputs(4985)) or (layer0_outputs(1613)));
    outputs(5396) <= not(layer0_outputs(9335));
    outputs(5397) <= layer0_outputs(689);
    outputs(5398) <= not(layer0_outputs(4023));
    outputs(5399) <= not(layer0_outputs(5521));
    outputs(5400) <= not(layer0_outputs(7888));
    outputs(5401) <= layer0_outputs(3873);
    outputs(5402) <= (layer0_outputs(2618)) and not (layer0_outputs(9208));
    outputs(5403) <= layer0_outputs(3545);
    outputs(5404) <= layer0_outputs(6793);
    outputs(5405) <= not((layer0_outputs(2862)) or (layer0_outputs(3687)));
    outputs(5406) <= not(layer0_outputs(272));
    outputs(5407) <= not(layer0_outputs(2570));
    outputs(5408) <= (layer0_outputs(2043)) and not (layer0_outputs(8813));
    outputs(5409) <= layer0_outputs(2055);
    outputs(5410) <= layer0_outputs(10118);
    outputs(5411) <= layer0_outputs(3683);
    outputs(5412) <= not(layer0_outputs(6309));
    outputs(5413) <= layer0_outputs(3392);
    outputs(5414) <= layer0_outputs(11955);
    outputs(5415) <= not(layer0_outputs(10167)) or (layer0_outputs(4168));
    outputs(5416) <= not(layer0_outputs(12273)) or (layer0_outputs(6181));
    outputs(5417) <= (layer0_outputs(5101)) and not (layer0_outputs(1489));
    outputs(5418) <= layer0_outputs(1663);
    outputs(5419) <= layer0_outputs(2310);
    outputs(5420) <= not((layer0_outputs(9610)) or (layer0_outputs(2340)));
    outputs(5421) <= (layer0_outputs(12711)) and not (layer0_outputs(8910));
    outputs(5422) <= not((layer0_outputs(764)) xor (layer0_outputs(8952)));
    outputs(5423) <= (layer0_outputs(1442)) and (layer0_outputs(8046));
    outputs(5424) <= (layer0_outputs(2927)) and (layer0_outputs(6397));
    outputs(5425) <= (layer0_outputs(194)) and not (layer0_outputs(4418));
    outputs(5426) <= not(layer0_outputs(1017));
    outputs(5427) <= not(layer0_outputs(6487)) or (layer0_outputs(6874));
    outputs(5428) <= not(layer0_outputs(84));
    outputs(5429) <= not(layer0_outputs(4088));
    outputs(5430) <= layer0_outputs(6100);
    outputs(5431) <= layer0_outputs(6402);
    outputs(5432) <= not((layer0_outputs(9764)) xor (layer0_outputs(5656)));
    outputs(5433) <= not((layer0_outputs(1481)) xor (layer0_outputs(6269)));
    outputs(5434) <= not(layer0_outputs(9511));
    outputs(5435) <= not(layer0_outputs(8223));
    outputs(5436) <= layer0_outputs(8366);
    outputs(5437) <= (layer0_outputs(6903)) and not (layer0_outputs(3654));
    outputs(5438) <= not(layer0_outputs(5616));
    outputs(5439) <= (layer0_outputs(6012)) and not (layer0_outputs(11512));
    outputs(5440) <= layer0_outputs(4117);
    outputs(5441) <= not(layer0_outputs(8543));
    outputs(5442) <= (layer0_outputs(12753)) and not (layer0_outputs(9072));
    outputs(5443) <= not((layer0_outputs(8670)) xor (layer0_outputs(5307)));
    outputs(5444) <= not(layer0_outputs(12117));
    outputs(5445) <= not(layer0_outputs(3226));
    outputs(5446) <= layer0_outputs(8973);
    outputs(5447) <= layer0_outputs(12270);
    outputs(5448) <= not((layer0_outputs(2857)) or (layer0_outputs(8962)));
    outputs(5449) <= not(layer0_outputs(6981));
    outputs(5450) <= layer0_outputs(7550);
    outputs(5451) <= not((layer0_outputs(5765)) or (layer0_outputs(5558)));
    outputs(5452) <= not(layer0_outputs(5132));
    outputs(5453) <= (layer0_outputs(4440)) and (layer0_outputs(4835));
    outputs(5454) <= (layer0_outputs(3269)) and not (layer0_outputs(12787));
    outputs(5455) <= (layer0_outputs(7267)) and not (layer0_outputs(5914));
    outputs(5456) <= (layer0_outputs(10349)) and not (layer0_outputs(6575));
    outputs(5457) <= (layer0_outputs(2720)) xor (layer0_outputs(6776));
    outputs(5458) <= (layer0_outputs(9952)) and not (layer0_outputs(3361));
    outputs(5459) <= not(layer0_outputs(3965));
    outputs(5460) <= layer0_outputs(10895);
    outputs(5461) <= not((layer0_outputs(3165)) xor (layer0_outputs(1423)));
    outputs(5462) <= not(layer0_outputs(5890));
    outputs(5463) <= not(layer0_outputs(4042));
    outputs(5464) <= layer0_outputs(7429);
    outputs(5465) <= not(layer0_outputs(5021));
    outputs(5466) <= layer0_outputs(2502);
    outputs(5467) <= not((layer0_outputs(8929)) xor (layer0_outputs(10602)));
    outputs(5468) <= not((layer0_outputs(8943)) and (layer0_outputs(3691)));
    outputs(5469) <= layer0_outputs(757);
    outputs(5470) <= not(layer0_outputs(7030));
    outputs(5471) <= layer0_outputs(1692);
    outputs(5472) <= not(layer0_outputs(12492));
    outputs(5473) <= not((layer0_outputs(5038)) and (layer0_outputs(9226)));
    outputs(5474) <= (layer0_outputs(9443)) and not (layer0_outputs(6454));
    outputs(5475) <= (layer0_outputs(11141)) xor (layer0_outputs(1711));
    outputs(5476) <= (layer0_outputs(627)) xor (layer0_outputs(6043));
    outputs(5477) <= not((layer0_outputs(8909)) and (layer0_outputs(7870)));
    outputs(5478) <= (layer0_outputs(1929)) and (layer0_outputs(7023));
    outputs(5479) <= layer0_outputs(11294);
    outputs(5480) <= layer0_outputs(10977);
    outputs(5481) <= not(layer0_outputs(5283));
    outputs(5482) <= layer0_outputs(3953);
    outputs(5483) <= layer0_outputs(11579);
    outputs(5484) <= not(layer0_outputs(7817)) or (layer0_outputs(6921));
    outputs(5485) <= not(layer0_outputs(12331));
    outputs(5486) <= not((layer0_outputs(1862)) xor (layer0_outputs(8628)));
    outputs(5487) <= not(layer0_outputs(6920));
    outputs(5488) <= not((layer0_outputs(5644)) and (layer0_outputs(11395)));
    outputs(5489) <= (layer0_outputs(6929)) and not (layer0_outputs(6532));
    outputs(5490) <= not(layer0_outputs(552));
    outputs(5491) <= layer0_outputs(226);
    outputs(5492) <= (layer0_outputs(8194)) and not (layer0_outputs(4263));
    outputs(5493) <= not((layer0_outputs(7403)) xor (layer0_outputs(10963)));
    outputs(5494) <= not(layer0_outputs(11244));
    outputs(5495) <= (layer0_outputs(3273)) and not (layer0_outputs(7466));
    outputs(5496) <= not(layer0_outputs(9706));
    outputs(5497) <= not(layer0_outputs(3764));
    outputs(5498) <= (layer0_outputs(6625)) xor (layer0_outputs(6718));
    outputs(5499) <= not(layer0_outputs(6543));
    outputs(5500) <= not((layer0_outputs(10971)) xor (layer0_outputs(2064)));
    outputs(5501) <= layer0_outputs(12628);
    outputs(5502) <= layer0_outputs(1837);
    outputs(5503) <= not((layer0_outputs(7811)) xor (layer0_outputs(3602)));
    outputs(5504) <= layer0_outputs(8781);
    outputs(5505) <= layer0_outputs(7748);
    outputs(5506) <= (layer0_outputs(9521)) and not (layer0_outputs(11078));
    outputs(5507) <= (layer0_outputs(7517)) and not (layer0_outputs(4965));
    outputs(5508) <= (layer0_outputs(10667)) xor (layer0_outputs(5285));
    outputs(5509) <= not(layer0_outputs(1861));
    outputs(5510) <= layer0_outputs(4331);
    outputs(5511) <= layer0_outputs(6642);
    outputs(5512) <= not(layer0_outputs(1200));
    outputs(5513) <= (layer0_outputs(9350)) xor (layer0_outputs(1949));
    outputs(5514) <= layer0_outputs(8665);
    outputs(5515) <= layer0_outputs(1524);
    outputs(5516) <= not(layer0_outputs(12735));
    outputs(5517) <= not(layer0_outputs(2278));
    outputs(5518) <= not(layer0_outputs(3549)) or (layer0_outputs(2161));
    outputs(5519) <= not((layer0_outputs(9819)) xor (layer0_outputs(4449)));
    outputs(5520) <= layer0_outputs(6163);
    outputs(5521) <= layer0_outputs(6740);
    outputs(5522) <= not((layer0_outputs(6787)) xor (layer0_outputs(10608)));
    outputs(5523) <= not(layer0_outputs(11618));
    outputs(5524) <= layer0_outputs(2899);
    outputs(5525) <= not((layer0_outputs(1466)) or (layer0_outputs(10032)));
    outputs(5526) <= (layer0_outputs(12649)) and (layer0_outputs(3353));
    outputs(5527) <= '0';
    outputs(5528) <= layer0_outputs(8794);
    outputs(5529) <= (layer0_outputs(3696)) and not (layer0_outputs(8424));
    outputs(5530) <= (layer0_outputs(2460)) and not (layer0_outputs(1737));
    outputs(5531) <= (layer0_outputs(10125)) and (layer0_outputs(11935));
    outputs(5532) <= not((layer0_outputs(9859)) or (layer0_outputs(9083)));
    outputs(5533) <= not(layer0_outputs(1339));
    outputs(5534) <= '0';
    outputs(5535) <= not((layer0_outputs(12645)) or (layer0_outputs(1569)));
    outputs(5536) <= (layer0_outputs(11827)) xor (layer0_outputs(7445));
    outputs(5537) <= not(layer0_outputs(11786));
    outputs(5538) <= layer0_outputs(12149);
    outputs(5539) <= layer0_outputs(12416);
    outputs(5540) <= not(layer0_outputs(1154));
    outputs(5541) <= not((layer0_outputs(3024)) or (layer0_outputs(6178)));
    outputs(5542) <= (layer0_outputs(4127)) and not (layer0_outputs(6597));
    outputs(5543) <= (layer0_outputs(247)) xor (layer0_outputs(6083));
    outputs(5544) <= (layer0_outputs(5300)) and not (layer0_outputs(8682));
    outputs(5545) <= not(layer0_outputs(12485));
    outputs(5546) <= (layer0_outputs(5771)) xor (layer0_outputs(5976));
    outputs(5547) <= not(layer0_outputs(4661));
    outputs(5548) <= layer0_outputs(5236);
    outputs(5549) <= layer0_outputs(292);
    outputs(5550) <= not((layer0_outputs(10460)) or (layer0_outputs(8375)));
    outputs(5551) <= (layer0_outputs(8607)) and (layer0_outputs(7949));
    outputs(5552) <= layer0_outputs(10054);
    outputs(5553) <= (layer0_outputs(4206)) and not (layer0_outputs(4955));
    outputs(5554) <= layer0_outputs(1736);
    outputs(5555) <= layer0_outputs(6934);
    outputs(5556) <= not(layer0_outputs(1833));
    outputs(5557) <= layer0_outputs(4523);
    outputs(5558) <= layer0_outputs(10158);
    outputs(5559) <= not(layer0_outputs(3069));
    outputs(5560) <= not(layer0_outputs(12202)) or (layer0_outputs(210));
    outputs(5561) <= layer0_outputs(3437);
    outputs(5562) <= not((layer0_outputs(3797)) xor (layer0_outputs(673)));
    outputs(5563) <= layer0_outputs(8190);
    outputs(5564) <= not(layer0_outputs(8418));
    outputs(5565) <= not(layer0_outputs(8846));
    outputs(5566) <= not(layer0_outputs(1191));
    outputs(5567) <= not((layer0_outputs(11331)) or (layer0_outputs(1261)));
    outputs(5568) <= (layer0_outputs(4654)) and not (layer0_outputs(11229));
    outputs(5569) <= (layer0_outputs(7802)) xor (layer0_outputs(2054));
    outputs(5570) <= not(layer0_outputs(11598));
    outputs(5571) <= layer0_outputs(6541);
    outputs(5572) <= layer0_outputs(2122);
    outputs(5573) <= (layer0_outputs(6126)) xor (layer0_outputs(11467));
    outputs(5574) <= layer0_outputs(596);
    outputs(5575) <= not(layer0_outputs(653));
    outputs(5576) <= not(layer0_outputs(10887));
    outputs(5577) <= not(layer0_outputs(12471)) or (layer0_outputs(1554));
    outputs(5578) <= (layer0_outputs(1033)) xor (layer0_outputs(1822));
    outputs(5579) <= not(layer0_outputs(5155));
    outputs(5580) <= not(layer0_outputs(10083));
    outputs(5581) <= not(layer0_outputs(5992));
    outputs(5582) <= not((layer0_outputs(12525)) or (layer0_outputs(9261)));
    outputs(5583) <= (layer0_outputs(10479)) and not (layer0_outputs(7146));
    outputs(5584) <= not((layer0_outputs(81)) xor (layer0_outputs(4720)));
    outputs(5585) <= layer0_outputs(11587);
    outputs(5586) <= not((layer0_outputs(9501)) and (layer0_outputs(2843)));
    outputs(5587) <= (layer0_outputs(7202)) and (layer0_outputs(7732));
    outputs(5588) <= not(layer0_outputs(4338));
    outputs(5589) <= not(layer0_outputs(3639));
    outputs(5590) <= not((layer0_outputs(12703)) xor (layer0_outputs(12664)));
    outputs(5591) <= not((layer0_outputs(10779)) xor (layer0_outputs(12325)));
    outputs(5592) <= (layer0_outputs(8258)) and not (layer0_outputs(8756));
    outputs(5593) <= (layer0_outputs(2783)) and (layer0_outputs(3627));
    outputs(5594) <= (layer0_outputs(5451)) xor (layer0_outputs(9292));
    outputs(5595) <= (layer0_outputs(5256)) and (layer0_outputs(3586));
    outputs(5596) <= (layer0_outputs(5410)) xor (layer0_outputs(10038));
    outputs(5597) <= not(layer0_outputs(12424));
    outputs(5598) <= not((layer0_outputs(1245)) xor (layer0_outputs(8176)));
    outputs(5599) <= not(layer0_outputs(1386));
    outputs(5600) <= not(layer0_outputs(3958));
    outputs(5601) <= (layer0_outputs(6823)) or (layer0_outputs(10846));
    outputs(5602) <= layer0_outputs(3759);
    outputs(5603) <= not(layer0_outputs(1075));
    outputs(5604) <= not(layer0_outputs(1306));
    outputs(5605) <= (layer0_outputs(782)) xor (layer0_outputs(3187));
    outputs(5606) <= (layer0_outputs(6428)) xor (layer0_outputs(11154));
    outputs(5607) <= not(layer0_outputs(12608));
    outputs(5608) <= not(layer0_outputs(9273));
    outputs(5609) <= layer0_outputs(8548);
    outputs(5610) <= not(layer0_outputs(3668));
    outputs(5611) <= layer0_outputs(8793);
    outputs(5612) <= (layer0_outputs(11717)) and not (layer0_outputs(9949));
    outputs(5613) <= not(layer0_outputs(3280));
    outputs(5614) <= (layer0_outputs(860)) and not (layer0_outputs(12672));
    outputs(5615) <= not((layer0_outputs(623)) xor (layer0_outputs(11809)));
    outputs(5616) <= not((layer0_outputs(9068)) xor (layer0_outputs(5199)));
    outputs(5617) <= not(layer0_outputs(11858));
    outputs(5618) <= layer0_outputs(6786);
    outputs(5619) <= not((layer0_outputs(2140)) or (layer0_outputs(34)));
    outputs(5620) <= (layer0_outputs(4376)) xor (layer0_outputs(5619));
    outputs(5621) <= layer0_outputs(11017);
    outputs(5622) <= not((layer0_outputs(599)) xor (layer0_outputs(1800)));
    outputs(5623) <= not((layer0_outputs(793)) and (layer0_outputs(4489)));
    outputs(5624) <= (layer0_outputs(8286)) and not (layer0_outputs(12432));
    outputs(5625) <= not((layer0_outputs(3762)) xor (layer0_outputs(1385)));
    outputs(5626) <= layer0_outputs(2496);
    outputs(5627) <= not((layer0_outputs(10347)) xor (layer0_outputs(9500)));
    outputs(5628) <= not(layer0_outputs(9107));
    outputs(5629) <= (layer0_outputs(12142)) and not (layer0_outputs(8844));
    outputs(5630) <= layer0_outputs(9523);
    outputs(5631) <= (layer0_outputs(735)) and not (layer0_outputs(7339));
    outputs(5632) <= (layer0_outputs(11972)) or (layer0_outputs(1570));
    outputs(5633) <= (layer0_outputs(4115)) and (layer0_outputs(11094));
    outputs(5634) <= (layer0_outputs(12216)) and (layer0_outputs(8946));
    outputs(5635) <= '0';
    outputs(5636) <= layer0_outputs(5327);
    outputs(5637) <= not(layer0_outputs(7184)) or (layer0_outputs(12760));
    outputs(5638) <= not(layer0_outputs(11488)) or (layer0_outputs(1543));
    outputs(5639) <= not(layer0_outputs(11787));
    outputs(5640) <= (layer0_outputs(7400)) and (layer0_outputs(2712));
    outputs(5641) <= (layer0_outputs(11817)) or (layer0_outputs(8605));
    outputs(5642) <= not((layer0_outputs(5585)) xor (layer0_outputs(4330)));
    outputs(5643) <= '0';
    outputs(5644) <= (layer0_outputs(9452)) xor (layer0_outputs(12412));
    outputs(5645) <= not((layer0_outputs(12223)) or (layer0_outputs(137)));
    outputs(5646) <= not((layer0_outputs(9689)) xor (layer0_outputs(2637)));
    outputs(5647) <= '0';
    outputs(5648) <= not((layer0_outputs(10517)) and (layer0_outputs(5058)));
    outputs(5649) <= layer0_outputs(3894);
    outputs(5650) <= (layer0_outputs(2073)) xor (layer0_outputs(6774));
    outputs(5651) <= layer0_outputs(1016);
    outputs(5652) <= (layer0_outputs(3710)) xor (layer0_outputs(8528));
    outputs(5653) <= not(layer0_outputs(12288)) or (layer0_outputs(4817));
    outputs(5654) <= (layer0_outputs(4060)) and not (layer0_outputs(5640));
    outputs(5655) <= not(layer0_outputs(1121));
    outputs(5656) <= not(layer0_outputs(3688));
    outputs(5657) <= not((layer0_outputs(7654)) xor (layer0_outputs(3314)));
    outputs(5658) <= (layer0_outputs(9397)) and (layer0_outputs(1794));
    outputs(5659) <= not(layer0_outputs(8274));
    outputs(5660) <= (layer0_outputs(4913)) and not (layer0_outputs(5296));
    outputs(5661) <= layer0_outputs(904);
    outputs(5662) <= not(layer0_outputs(5275)) or (layer0_outputs(3076));
    outputs(5663) <= not(layer0_outputs(5606));
    outputs(5664) <= not(layer0_outputs(11822));
    outputs(5665) <= not(layer0_outputs(12434)) or (layer0_outputs(4096));
    outputs(5666) <= layer0_outputs(1648);
    outputs(5667) <= not((layer0_outputs(1623)) xor (layer0_outputs(5493)));
    outputs(5668) <= (layer0_outputs(9704)) xor (layer0_outputs(9078));
    outputs(5669) <= not((layer0_outputs(11937)) or (layer0_outputs(705)));
    outputs(5670) <= not(layer0_outputs(2881));
    outputs(5671) <= not((layer0_outputs(3169)) and (layer0_outputs(3389)));
    outputs(5672) <= layer0_outputs(9270);
    outputs(5673) <= not(layer0_outputs(467));
    outputs(5674) <= not((layer0_outputs(8469)) and (layer0_outputs(9816)));
    outputs(5675) <= (layer0_outputs(2160)) xor (layer0_outputs(3152));
    outputs(5676) <= not(layer0_outputs(8065));
    outputs(5677) <= (layer0_outputs(6201)) or (layer0_outputs(11557));
    outputs(5678) <= layer0_outputs(4686);
    outputs(5679) <= not(layer0_outputs(12062)) or (layer0_outputs(9085));
    outputs(5680) <= layer0_outputs(668);
    outputs(5681) <= not((layer0_outputs(8629)) or (layer0_outputs(12259)));
    outputs(5682) <= layer0_outputs(12095);
    outputs(5683) <= not((layer0_outputs(3948)) or (layer0_outputs(8853)));
    outputs(5684) <= layer0_outputs(11358);
    outputs(5685) <= (layer0_outputs(5059)) xor (layer0_outputs(6296));
    outputs(5686) <= (layer0_outputs(3282)) and not (layer0_outputs(1868));
    outputs(5687) <= not(layer0_outputs(12375));
    outputs(5688) <= not((layer0_outputs(6976)) and (layer0_outputs(12375)));
    outputs(5689) <= (layer0_outputs(12330)) and (layer0_outputs(7014));
    outputs(5690) <= (layer0_outputs(11403)) and not (layer0_outputs(9628));
    outputs(5691) <= (layer0_outputs(594)) and (layer0_outputs(6388));
    outputs(5692) <= not(layer0_outputs(4877));
    outputs(5693) <= layer0_outputs(12160);
    outputs(5694) <= not(layer0_outputs(1552)) or (layer0_outputs(1301));
    outputs(5695) <= layer0_outputs(3074);
    outputs(5696) <= not((layer0_outputs(8407)) xor (layer0_outputs(8527)));
    outputs(5697) <= not(layer0_outputs(6411)) or (layer0_outputs(1113));
    outputs(5698) <= (layer0_outputs(3394)) and not (layer0_outputs(5467));
    outputs(5699) <= not(layer0_outputs(10259)) or (layer0_outputs(12205));
    outputs(5700) <= (layer0_outputs(10324)) and (layer0_outputs(718));
    outputs(5701) <= not(layer0_outputs(11433));
    outputs(5702) <= layer0_outputs(469);
    outputs(5703) <= (layer0_outputs(11807)) and not (layer0_outputs(7835));
    outputs(5704) <= (layer0_outputs(10028)) or (layer0_outputs(11205));
    outputs(5705) <= '0';
    outputs(5706) <= layer0_outputs(4898);
    outputs(5707) <= not(layer0_outputs(3015));
    outputs(5708) <= not((layer0_outputs(9017)) or (layer0_outputs(9548)));
    outputs(5709) <= (layer0_outputs(6390)) and not (layer0_outputs(988));
    outputs(5710) <= '1';
    outputs(5711) <= not(layer0_outputs(7279));
    outputs(5712) <= not(layer0_outputs(11902));
    outputs(5713) <= layer0_outputs(4904);
    outputs(5714) <= layer0_outputs(8135);
    outputs(5715) <= (layer0_outputs(9100)) xor (layer0_outputs(5179));
    outputs(5716) <= not(layer0_outputs(3465)) or (layer0_outputs(8605));
    outputs(5717) <= layer0_outputs(11146);
    outputs(5718) <= not(layer0_outputs(7279));
    outputs(5719) <= (layer0_outputs(8848)) and (layer0_outputs(5779));
    outputs(5720) <= layer0_outputs(9133);
    outputs(5721) <= not((layer0_outputs(5783)) xor (layer0_outputs(12227)));
    outputs(5722) <= (layer0_outputs(10447)) xor (layer0_outputs(11129));
    outputs(5723) <= not(layer0_outputs(2661));
    outputs(5724) <= not(layer0_outputs(10539));
    outputs(5725) <= (layer0_outputs(5448)) xor (layer0_outputs(5312));
    outputs(5726) <= not(layer0_outputs(2696));
    outputs(5727) <= not(layer0_outputs(10588)) or (layer0_outputs(340));
    outputs(5728) <= layer0_outputs(11282);
    outputs(5729) <= not(layer0_outputs(7923));
    outputs(5730) <= layer0_outputs(8803);
    outputs(5731) <= (layer0_outputs(2840)) xor (layer0_outputs(2052));
    outputs(5732) <= layer0_outputs(12657);
    outputs(5733) <= not((layer0_outputs(3081)) and (layer0_outputs(2200)));
    outputs(5734) <= not((layer0_outputs(5194)) xor (layer0_outputs(2826)));
    outputs(5735) <= (layer0_outputs(7885)) xor (layer0_outputs(10873));
    outputs(5736) <= layer0_outputs(8841);
    outputs(5737) <= (layer0_outputs(4307)) xor (layer0_outputs(4891));
    outputs(5738) <= layer0_outputs(9420);
    outputs(5739) <= not((layer0_outputs(1527)) and (layer0_outputs(2761)));
    outputs(5740) <= (layer0_outputs(4027)) and not (layer0_outputs(9350));
    outputs(5741) <= (layer0_outputs(6178)) xor (layer0_outputs(4519));
    outputs(5742) <= (layer0_outputs(4898)) and not (layer0_outputs(12386));
    outputs(5743) <= not((layer0_outputs(10888)) or (layer0_outputs(2333)));
    outputs(5744) <= (layer0_outputs(98)) xor (layer0_outputs(9878));
    outputs(5745) <= (layer0_outputs(1508)) xor (layer0_outputs(6268));
    outputs(5746) <= not(layer0_outputs(1264));
    outputs(5747) <= layer0_outputs(12201);
    outputs(5748) <= layer0_outputs(5427);
    outputs(5749) <= not((layer0_outputs(8181)) xor (layer0_outputs(1536)));
    outputs(5750) <= (layer0_outputs(3771)) and not (layer0_outputs(11550));
    outputs(5751) <= not((layer0_outputs(1431)) xor (layer0_outputs(9008)));
    outputs(5752) <= layer0_outputs(2820);
    outputs(5753) <= layer0_outputs(5750);
    outputs(5754) <= (layer0_outputs(3853)) xor (layer0_outputs(11553));
    outputs(5755) <= not(layer0_outputs(9416));
    outputs(5756) <= (layer0_outputs(7032)) and not (layer0_outputs(715));
    outputs(5757) <= (layer0_outputs(5884)) and not (layer0_outputs(9305));
    outputs(5758) <= (layer0_outputs(11732)) and not (layer0_outputs(3829));
    outputs(5759) <= layer0_outputs(1549);
    outputs(5760) <= not((layer0_outputs(1823)) xor (layer0_outputs(8530)));
    outputs(5761) <= (layer0_outputs(1681)) and not (layer0_outputs(6591));
    outputs(5762) <= not(layer0_outputs(10335));
    outputs(5763) <= not(layer0_outputs(7299));
    outputs(5764) <= not((layer0_outputs(11533)) or (layer0_outputs(3020)));
    outputs(5765) <= not(layer0_outputs(10583)) or (layer0_outputs(10351));
    outputs(5766) <= (layer0_outputs(2684)) and not (layer0_outputs(11443));
    outputs(5767) <= not((layer0_outputs(2277)) xor (layer0_outputs(1210)));
    outputs(5768) <= layer0_outputs(4925);
    outputs(5769) <= (layer0_outputs(9888)) xor (layer0_outputs(6393));
    outputs(5770) <= layer0_outputs(10769);
    outputs(5771) <= not(layer0_outputs(7083));
    outputs(5772) <= not(layer0_outputs(6915));
    outputs(5773) <= layer0_outputs(3807);
    outputs(5774) <= (layer0_outputs(10957)) and (layer0_outputs(11362));
    outputs(5775) <= not((layer0_outputs(150)) xor (layer0_outputs(9418)));
    outputs(5776) <= layer0_outputs(12074);
    outputs(5777) <= not(layer0_outputs(5434));
    outputs(5778) <= (layer0_outputs(4783)) and not (layer0_outputs(5760));
    outputs(5779) <= not((layer0_outputs(4195)) xor (layer0_outputs(1636)));
    outputs(5780) <= not(layer0_outputs(6971));
    outputs(5781) <= not(layer0_outputs(3513));
    outputs(5782) <= layer0_outputs(32);
    outputs(5783) <= not(layer0_outputs(7318));
    outputs(5784) <= (layer0_outputs(12132)) and not (layer0_outputs(11265));
    outputs(5785) <= (layer0_outputs(193)) and not (layer0_outputs(8362));
    outputs(5786) <= layer0_outputs(5930);
    outputs(5787) <= (layer0_outputs(12119)) and not (layer0_outputs(12552));
    outputs(5788) <= not(layer0_outputs(10131));
    outputs(5789) <= not(layer0_outputs(9690));
    outputs(5790) <= not((layer0_outputs(9685)) xor (layer0_outputs(7908)));
    outputs(5791) <= not(layer0_outputs(5280));
    outputs(5792) <= not(layer0_outputs(4912)) or (layer0_outputs(898));
    outputs(5793) <= not(layer0_outputs(4572)) or (layer0_outputs(12412));
    outputs(5794) <= (layer0_outputs(10196)) xor (layer0_outputs(1887));
    outputs(5795) <= (layer0_outputs(3812)) and not (layer0_outputs(7414));
    outputs(5796) <= (layer0_outputs(9443)) and not (layer0_outputs(5469));
    outputs(5797) <= (layer0_outputs(8696)) and not (layer0_outputs(154));
    outputs(5798) <= not(layer0_outputs(2870)) or (layer0_outputs(3734));
    outputs(5799) <= (layer0_outputs(6643)) and not (layer0_outputs(10502));
    outputs(5800) <= (layer0_outputs(11074)) and (layer0_outputs(5537));
    outputs(5801) <= layer0_outputs(7001);
    outputs(5802) <= (layer0_outputs(892)) or (layer0_outputs(4142));
    outputs(5803) <= (layer0_outputs(6664)) and not (layer0_outputs(5190));
    outputs(5804) <= (layer0_outputs(5129)) and (layer0_outputs(3221));
    outputs(5805) <= '0';
    outputs(5806) <= (layer0_outputs(12010)) and not (layer0_outputs(4485));
    outputs(5807) <= (layer0_outputs(10234)) and not (layer0_outputs(7769));
    outputs(5808) <= not((layer0_outputs(3496)) xor (layer0_outputs(915)));
    outputs(5809) <= (layer0_outputs(2538)) and not (layer0_outputs(12047));
    outputs(5810) <= (layer0_outputs(10751)) and not (layer0_outputs(4230));
    outputs(5811) <= (layer0_outputs(3357)) and not (layer0_outputs(2808));
    outputs(5812) <= not((layer0_outputs(7831)) xor (layer0_outputs(10001)));
    outputs(5813) <= not(layer0_outputs(8805));
    outputs(5814) <= not(layer0_outputs(11826));
    outputs(5815) <= (layer0_outputs(11371)) and not (layer0_outputs(2541));
    outputs(5816) <= layer0_outputs(7343);
    outputs(5817) <= layer0_outputs(12785);
    outputs(5818) <= not(layer0_outputs(3120));
    outputs(5819) <= not((layer0_outputs(5965)) xor (layer0_outputs(3406)));
    outputs(5820) <= (layer0_outputs(2997)) xor (layer0_outputs(12317));
    outputs(5821) <= not((layer0_outputs(4587)) xor (layer0_outputs(8285)));
    outputs(5822) <= not((layer0_outputs(7069)) xor (layer0_outputs(3994)));
    outputs(5823) <= layer0_outputs(8575);
    outputs(5824) <= (layer0_outputs(10544)) xor (layer0_outputs(4737));
    outputs(5825) <= not((layer0_outputs(276)) or (layer0_outputs(10948)));
    outputs(5826) <= layer0_outputs(2670);
    outputs(5827) <= (layer0_outputs(5048)) and (layer0_outputs(5026));
    outputs(5828) <= not(layer0_outputs(10863));
    outputs(5829) <= not((layer0_outputs(9547)) or (layer0_outputs(8809)));
    outputs(5830) <= not((layer0_outputs(6707)) and (layer0_outputs(2097)));
    outputs(5831) <= not((layer0_outputs(4091)) or (layer0_outputs(7670)));
    outputs(5832) <= (layer0_outputs(5583)) and not (layer0_outputs(1358));
    outputs(5833) <= not((layer0_outputs(3940)) or (layer0_outputs(11337)));
    outputs(5834) <= not((layer0_outputs(7516)) or (layer0_outputs(175)));
    outputs(5835) <= layer0_outputs(415);
    outputs(5836) <= layer0_outputs(9869);
    outputs(5837) <= not(layer0_outputs(4595));
    outputs(5838) <= not(layer0_outputs(1049));
    outputs(5839) <= not(layer0_outputs(899));
    outputs(5840) <= not((layer0_outputs(7598)) xor (layer0_outputs(1591)));
    outputs(5841) <= (layer0_outputs(12295)) and (layer0_outputs(8291));
    outputs(5842) <= not(layer0_outputs(9216));
    outputs(5843) <= not(layer0_outputs(6133));
    outputs(5844) <= (layer0_outputs(2206)) and not (layer0_outputs(6560));
    outputs(5845) <= not(layer0_outputs(10670));
    outputs(5846) <= (layer0_outputs(10378)) xor (layer0_outputs(975));
    outputs(5847) <= (layer0_outputs(8757)) and not (layer0_outputs(2529));
    outputs(5848) <= (layer0_outputs(7950)) and (layer0_outputs(4470));
    outputs(5849) <= layer0_outputs(5580);
    outputs(5850) <= (layer0_outputs(5022)) and (layer0_outputs(6846));
    outputs(5851) <= not(layer0_outputs(11272));
    outputs(5852) <= layer0_outputs(2442);
    outputs(5853) <= not(layer0_outputs(6752));
    outputs(5854) <= (layer0_outputs(2054)) xor (layer0_outputs(9185));
    outputs(5855) <= (layer0_outputs(4156)) xor (layer0_outputs(5707));
    outputs(5856) <= (layer0_outputs(7951)) and not (layer0_outputs(10722));
    outputs(5857) <= layer0_outputs(6051);
    outputs(5858) <= not(layer0_outputs(11067));
    outputs(5859) <= (layer0_outputs(7042)) and not (layer0_outputs(1242));
    outputs(5860) <= not((layer0_outputs(7424)) xor (layer0_outputs(570)));
    outputs(5861) <= not((layer0_outputs(8660)) xor (layer0_outputs(12695)));
    outputs(5862) <= (layer0_outputs(7923)) and (layer0_outputs(4814));
    outputs(5863) <= layer0_outputs(12568);
    outputs(5864) <= not(layer0_outputs(8913)) or (layer0_outputs(6108));
    outputs(5865) <= not(layer0_outputs(3120));
    outputs(5866) <= (layer0_outputs(2727)) xor (layer0_outputs(8475));
    outputs(5867) <= not(layer0_outputs(9394));
    outputs(5868) <= layer0_outputs(6371);
    outputs(5869) <= not((layer0_outputs(10038)) and (layer0_outputs(5314)));
    outputs(5870) <= (layer0_outputs(5234)) or (layer0_outputs(475));
    outputs(5871) <= (layer0_outputs(4981)) xor (layer0_outputs(7245));
    outputs(5872) <= not(layer0_outputs(2576));
    outputs(5873) <= (layer0_outputs(387)) or (layer0_outputs(1922));
    outputs(5874) <= (layer0_outputs(12529)) and not (layer0_outputs(3446));
    outputs(5875) <= (layer0_outputs(3765)) and (layer0_outputs(6168));
    outputs(5876) <= (layer0_outputs(4764)) and not (layer0_outputs(288));
    outputs(5877) <= (layer0_outputs(8868)) and not (layer0_outputs(1915));
    outputs(5878) <= not((layer0_outputs(7090)) and (layer0_outputs(7006)));
    outputs(5879) <= layer0_outputs(11506);
    outputs(5880) <= not(layer0_outputs(691));
    outputs(5881) <= (layer0_outputs(2424)) and not (layer0_outputs(5698));
    outputs(5882) <= layer0_outputs(5772);
    outputs(5883) <= not(layer0_outputs(69));
    outputs(5884) <= layer0_outputs(8889);
    outputs(5885) <= layer0_outputs(3303);
    outputs(5886) <= layer0_outputs(2323);
    outputs(5887) <= (layer0_outputs(4910)) xor (layer0_outputs(2687));
    outputs(5888) <= layer0_outputs(4498);
    outputs(5889) <= (layer0_outputs(4552)) xor (layer0_outputs(200));
    outputs(5890) <= layer0_outputs(6979);
    outputs(5891) <= not(layer0_outputs(3581));
    outputs(5892) <= layer0_outputs(2280);
    outputs(5893) <= (layer0_outputs(10241)) xor (layer0_outputs(11588));
    outputs(5894) <= (layer0_outputs(9783)) and (layer0_outputs(3919));
    outputs(5895) <= not((layer0_outputs(10166)) or (layer0_outputs(9882)));
    outputs(5896) <= not(layer0_outputs(5880));
    outputs(5897) <= (layer0_outputs(8768)) and not (layer0_outputs(1934));
    outputs(5898) <= '0';
    outputs(5899) <= not((layer0_outputs(2144)) xor (layer0_outputs(6900)));
    outputs(5900) <= (layer0_outputs(7096)) and (layer0_outputs(6239));
    outputs(5901) <= layer0_outputs(11058);
    outputs(5902) <= not(layer0_outputs(1086));
    outputs(5903) <= not((layer0_outputs(5859)) or (layer0_outputs(8908)));
    outputs(5904) <= (layer0_outputs(5337)) and (layer0_outputs(6123));
    outputs(5905) <= (layer0_outputs(12119)) and (layer0_outputs(4074));
    outputs(5906) <= not((layer0_outputs(3770)) or (layer0_outputs(5373)));
    outputs(5907) <= (layer0_outputs(1942)) xor (layer0_outputs(8729));
    outputs(5908) <= layer0_outputs(3400);
    outputs(5909) <= (layer0_outputs(10365)) and (layer0_outputs(10819));
    outputs(5910) <= not((layer0_outputs(1954)) xor (layer0_outputs(9286)));
    outputs(5911) <= not((layer0_outputs(4046)) or (layer0_outputs(7916)));
    outputs(5912) <= not((layer0_outputs(3252)) xor (layer0_outputs(6489)));
    outputs(5913) <= layer0_outputs(3182);
    outputs(5914) <= not((layer0_outputs(11766)) xor (layer0_outputs(3743)));
    outputs(5915) <= not((layer0_outputs(12071)) or (layer0_outputs(12486)));
    outputs(5916) <= (layer0_outputs(2262)) xor (layer0_outputs(5421));
    outputs(5917) <= not((layer0_outputs(12429)) or (layer0_outputs(6079)));
    outputs(5918) <= (layer0_outputs(5048)) and not (layer0_outputs(5658));
    outputs(5919) <= (layer0_outputs(983)) and not (layer0_outputs(8340));
    outputs(5920) <= not(layer0_outputs(10576));
    outputs(5921) <= (layer0_outputs(4169)) or (layer0_outputs(5622));
    outputs(5922) <= not(layer0_outputs(6665)) or (layer0_outputs(4664));
    outputs(5923) <= not((layer0_outputs(2643)) xor (layer0_outputs(5828)));
    outputs(5924) <= (layer0_outputs(1425)) and not (layer0_outputs(11792));
    outputs(5925) <= (layer0_outputs(4712)) and not (layer0_outputs(5628));
    outputs(5926) <= not((layer0_outputs(2824)) or (layer0_outputs(10217)));
    outputs(5927) <= layer0_outputs(957);
    outputs(5928) <= (layer0_outputs(1433)) xor (layer0_outputs(8112));
    outputs(5929) <= (layer0_outputs(10971)) and (layer0_outputs(10120));
    outputs(5930) <= (layer0_outputs(3704)) and (layer0_outputs(3185));
    outputs(5931) <= not(layer0_outputs(12796));
    outputs(5932) <= (layer0_outputs(4818)) xor (layer0_outputs(10922));
    outputs(5933) <= not(layer0_outputs(11359));
    outputs(5934) <= layer0_outputs(1293);
    outputs(5935) <= not(layer0_outputs(6090));
    outputs(5936) <= not(layer0_outputs(5542));
    outputs(5937) <= (layer0_outputs(7661)) xor (layer0_outputs(6074));
    outputs(5938) <= (layer0_outputs(10781)) and not (layer0_outputs(3258));
    outputs(5939) <= not(layer0_outputs(2523)) or (layer0_outputs(829));
    outputs(5940) <= layer0_outputs(2953);
    outputs(5941) <= not(layer0_outputs(1861)) or (layer0_outputs(9918));
    outputs(5942) <= (layer0_outputs(7072)) xor (layer0_outputs(11491));
    outputs(5943) <= (layer0_outputs(2237)) xor (layer0_outputs(10392));
    outputs(5944) <= (layer0_outputs(3620)) and (layer0_outputs(1970));
    outputs(5945) <= (layer0_outputs(6581)) and not (layer0_outputs(3645));
    outputs(5946) <= not((layer0_outputs(5944)) or (layer0_outputs(9147)));
    outputs(5947) <= not(layer0_outputs(1959)) or (layer0_outputs(1873));
    outputs(5948) <= not(layer0_outputs(7931));
    outputs(5949) <= not(layer0_outputs(8136));
    outputs(5950) <= layer0_outputs(11947);
    outputs(5951) <= not((layer0_outputs(6719)) and (layer0_outputs(12337)));
    outputs(5952) <= not(layer0_outputs(3365));
    outputs(5953) <= not((layer0_outputs(3085)) xor (layer0_outputs(8068)));
    outputs(5954) <= not((layer0_outputs(7536)) xor (layer0_outputs(2707)));
    outputs(5955) <= (layer0_outputs(8009)) xor (layer0_outputs(11547));
    outputs(5956) <= not(layer0_outputs(5681));
    outputs(5957) <= not(layer0_outputs(10928)) or (layer0_outputs(834));
    outputs(5958) <= not(layer0_outputs(10820));
    outputs(5959) <= not((layer0_outputs(1610)) xor (layer0_outputs(8305)));
    outputs(5960) <= not((layer0_outputs(5570)) xor (layer0_outputs(4266)));
    outputs(5961) <= (layer0_outputs(8740)) and not (layer0_outputs(11920));
    outputs(5962) <= not((layer0_outputs(10154)) or (layer0_outputs(7931)));
    outputs(5963) <= (layer0_outputs(10821)) xor (layer0_outputs(1917));
    outputs(5964) <= (layer0_outputs(5152)) and not (layer0_outputs(1452));
    outputs(5965) <= layer0_outputs(10484);
    outputs(5966) <= not(layer0_outputs(432));
    outputs(5967) <= not(layer0_outputs(8196));
    outputs(5968) <= not((layer0_outputs(2703)) xor (layer0_outputs(749)));
    outputs(5969) <= layer0_outputs(568);
    outputs(5970) <= (layer0_outputs(10511)) and not (layer0_outputs(6951));
    outputs(5971) <= not(layer0_outputs(3110));
    outputs(5972) <= (layer0_outputs(3359)) or (layer0_outputs(6293));
    outputs(5973) <= layer0_outputs(576);
    outputs(5974) <= not((layer0_outputs(11038)) xor (layer0_outputs(10393)));
    outputs(5975) <= not(layer0_outputs(2247));
    outputs(5976) <= (layer0_outputs(10925)) xor (layer0_outputs(6036));
    outputs(5977) <= (layer0_outputs(8582)) and not (layer0_outputs(2348));
    outputs(5978) <= not(layer0_outputs(7733));
    outputs(5979) <= not(layer0_outputs(5391));
    outputs(5980) <= layer0_outputs(10199);
    outputs(5981) <= (layer0_outputs(7647)) and not (layer0_outputs(979));
    outputs(5982) <= not(layer0_outputs(9038));
    outputs(5983) <= not(layer0_outputs(1166));
    outputs(5984) <= (layer0_outputs(3494)) xor (layer0_outputs(62));
    outputs(5985) <= not(layer0_outputs(3680));
    outputs(5986) <= not(layer0_outputs(8287));
    outputs(5987) <= (layer0_outputs(11106)) xor (layer0_outputs(8319));
    outputs(5988) <= not(layer0_outputs(6170));
    outputs(5989) <= (layer0_outputs(8867)) or (layer0_outputs(93));
    outputs(5990) <= not((layer0_outputs(4487)) and (layer0_outputs(3510)));
    outputs(5991) <= not((layer0_outputs(2700)) xor (layer0_outputs(2098)));
    outputs(5992) <= not(layer0_outputs(8400));
    outputs(5993) <= not(layer0_outputs(10521));
    outputs(5994) <= not(layer0_outputs(5603)) or (layer0_outputs(10757));
    outputs(5995) <= not((layer0_outputs(8416)) or (layer0_outputs(4150)));
    outputs(5996) <= not((layer0_outputs(7455)) and (layer0_outputs(6255)));
    outputs(5997) <= (layer0_outputs(8497)) xor (layer0_outputs(10637));
    outputs(5998) <= layer0_outputs(8210);
    outputs(5999) <= layer0_outputs(4772);
    outputs(6000) <= not(layer0_outputs(6056)) or (layer0_outputs(2496));
    outputs(6001) <= layer0_outputs(932);
    outputs(6002) <= (layer0_outputs(810)) and not (layer0_outputs(7875));
    outputs(6003) <= not(layer0_outputs(8179));
    outputs(6004) <= not(layer0_outputs(1343));
    outputs(6005) <= not((layer0_outputs(2167)) xor (layer0_outputs(12016)));
    outputs(6006) <= not((layer0_outputs(12242)) xor (layer0_outputs(9742)));
    outputs(6007) <= (layer0_outputs(6881)) and (layer0_outputs(10585));
    outputs(6008) <= '0';
    outputs(6009) <= (layer0_outputs(7196)) xor (layer0_outputs(10454));
    outputs(6010) <= layer0_outputs(7976);
    outputs(6011) <= (layer0_outputs(4733)) and not (layer0_outputs(3239));
    outputs(6012) <= layer0_outputs(5723);
    outputs(6013) <= not((layer0_outputs(2849)) or (layer0_outputs(9155)));
    outputs(6014) <= layer0_outputs(8724);
    outputs(6015) <= (layer0_outputs(8041)) and (layer0_outputs(5073));
    outputs(6016) <= layer0_outputs(9378);
    outputs(6017) <= not((layer0_outputs(2305)) xor (layer0_outputs(12660)));
    outputs(6018) <= not(layer0_outputs(6530));
    outputs(6019) <= (layer0_outputs(10559)) and not (layer0_outputs(695));
    outputs(6020) <= not((layer0_outputs(2394)) and (layer0_outputs(12294)));
    outputs(6021) <= not(layer0_outputs(10738)) or (layer0_outputs(5870));
    outputs(6022) <= not(layer0_outputs(5542));
    outputs(6023) <= layer0_outputs(10120);
    outputs(6024) <= not((layer0_outputs(1825)) and (layer0_outputs(827)));
    outputs(6025) <= not((layer0_outputs(8780)) or (layer0_outputs(1880)));
    outputs(6026) <= not((layer0_outputs(12349)) or (layer0_outputs(4133)));
    outputs(6027) <= layer0_outputs(11799);
    outputs(6028) <= not(layer0_outputs(7149));
    outputs(6029) <= (layer0_outputs(7575)) and not (layer0_outputs(2818));
    outputs(6030) <= layer0_outputs(12440);
    outputs(6031) <= not(layer0_outputs(65));
    outputs(6032) <= not(layer0_outputs(5536));
    outputs(6033) <= (layer0_outputs(6328)) and not (layer0_outputs(4365));
    outputs(6034) <= not(layer0_outputs(7189));
    outputs(6035) <= not((layer0_outputs(2844)) and (layer0_outputs(5352)));
    outputs(6036) <= (layer0_outputs(11283)) xor (layer0_outputs(2572));
    outputs(6037) <= (layer0_outputs(11589)) or (layer0_outputs(8198));
    outputs(6038) <= not((layer0_outputs(3405)) xor (layer0_outputs(9691)));
    outputs(6039) <= not((layer0_outputs(7415)) xor (layer0_outputs(6301)));
    outputs(6040) <= not((layer0_outputs(9512)) xor (layer0_outputs(9665)));
    outputs(6041) <= not((layer0_outputs(7050)) xor (layer0_outputs(12578)));
    outputs(6042) <= (layer0_outputs(7929)) and (layer0_outputs(5888));
    outputs(6043) <= not(layer0_outputs(7553));
    outputs(6044) <= not((layer0_outputs(7679)) xor (layer0_outputs(10654)));
    outputs(6045) <= not(layer0_outputs(11117));
    outputs(6046) <= layer0_outputs(2266);
    outputs(6047) <= layer0_outputs(12694);
    outputs(6048) <= (layer0_outputs(2837)) and not (layer0_outputs(3923));
    outputs(6049) <= (layer0_outputs(3969)) xor (layer0_outputs(278));
    outputs(6050) <= not(layer0_outputs(7173)) or (layer0_outputs(4817));
    outputs(6051) <= not(layer0_outputs(4973));
    outputs(6052) <= layer0_outputs(8576);
    outputs(6053) <= not((layer0_outputs(7553)) and (layer0_outputs(4126)));
    outputs(6054) <= layer0_outputs(5925);
    outputs(6055) <= not(layer0_outputs(3596));
    outputs(6056) <= layer0_outputs(8976);
    outputs(6057) <= not((layer0_outputs(9176)) xor (layer0_outputs(3450)));
    outputs(6058) <= (layer0_outputs(11202)) or (layer0_outputs(1466));
    outputs(6059) <= '0';
    outputs(6060) <= (layer0_outputs(9006)) and not (layer0_outputs(8435));
    outputs(6061) <= (layer0_outputs(4545)) and not (layer0_outputs(9174));
    outputs(6062) <= (layer0_outputs(1539)) and not (layer0_outputs(3559));
    outputs(6063) <= (layer0_outputs(3091)) xor (layer0_outputs(10554));
    outputs(6064) <= (layer0_outputs(7995)) and (layer0_outputs(5432));
    outputs(6065) <= layer0_outputs(2887);
    outputs(6066) <= layer0_outputs(6874);
    outputs(6067) <= not(layer0_outputs(3212));
    outputs(6068) <= not((layer0_outputs(6052)) xor (layer0_outputs(12399)));
    outputs(6069) <= (layer0_outputs(9732)) and not (layer0_outputs(4708));
    outputs(6070) <= (layer0_outputs(9471)) and (layer0_outputs(5301));
    outputs(6071) <= (layer0_outputs(4014)) xor (layer0_outputs(2464));
    outputs(6072) <= layer0_outputs(4301);
    outputs(6073) <= not(layer0_outputs(5982));
    outputs(6074) <= not(layer0_outputs(7797));
    outputs(6075) <= layer0_outputs(7151);
    outputs(6076) <= layer0_outputs(10695);
    outputs(6077) <= layer0_outputs(4956);
    outputs(6078) <= not(layer0_outputs(70));
    outputs(6079) <= (layer0_outputs(3644)) xor (layer0_outputs(5835));
    outputs(6080) <= not((layer0_outputs(10353)) and (layer0_outputs(3127)));
    outputs(6081) <= (layer0_outputs(9185)) and not (layer0_outputs(2504));
    outputs(6082) <= not(layer0_outputs(2492));
    outputs(6083) <= (layer0_outputs(6052)) and not (layer0_outputs(11344));
    outputs(6084) <= layer0_outputs(1442);
    outputs(6085) <= (layer0_outputs(8300)) and not (layer0_outputs(8685));
    outputs(6086) <= (layer0_outputs(7887)) and (layer0_outputs(7116));
    outputs(6087) <= (layer0_outputs(12181)) and not (layer0_outputs(4586));
    outputs(6088) <= (layer0_outputs(10112)) and not (layer0_outputs(8142));
    outputs(6089) <= not((layer0_outputs(7379)) xor (layer0_outputs(257)));
    outputs(6090) <= (layer0_outputs(4685)) xor (layer0_outputs(5068));
    outputs(6091) <= not(layer0_outputs(11497));
    outputs(6092) <= (layer0_outputs(9999)) and not (layer0_outputs(1387));
    outputs(6093) <= layer0_outputs(8691);
    outputs(6094) <= layer0_outputs(9001);
    outputs(6095) <= (layer0_outputs(5816)) or (layer0_outputs(188));
    outputs(6096) <= not((layer0_outputs(1783)) xor (layer0_outputs(6012)));
    outputs(6097) <= layer0_outputs(4292);
    outputs(6098) <= not((layer0_outputs(11655)) xor (layer0_outputs(4759)));
    outputs(6099) <= (layer0_outputs(11752)) xor (layer0_outputs(2708));
    outputs(6100) <= (layer0_outputs(3934)) xor (layer0_outputs(7504));
    outputs(6101) <= (layer0_outputs(2678)) and not (layer0_outputs(5878));
    outputs(6102) <= (layer0_outputs(6514)) and not (layer0_outputs(4849));
    outputs(6103) <= not(layer0_outputs(12263));
    outputs(6104) <= layer0_outputs(1131);
    outputs(6105) <= (layer0_outputs(10352)) and not (layer0_outputs(2131));
    outputs(6106) <= not(layer0_outputs(4120));
    outputs(6107) <= not(layer0_outputs(321));
    outputs(6108) <= layer0_outputs(2670);
    outputs(6109) <= (layer0_outputs(2152)) xor (layer0_outputs(9189));
    outputs(6110) <= not(layer0_outputs(6913));
    outputs(6111) <= not(layer0_outputs(1202)) or (layer0_outputs(9009));
    outputs(6112) <= not((layer0_outputs(11883)) or (layer0_outputs(4906)));
    outputs(6113) <= not((layer0_outputs(11135)) or (layer0_outputs(11425)));
    outputs(6114) <= not(layer0_outputs(10136));
    outputs(6115) <= (layer0_outputs(487)) xor (layer0_outputs(11181));
    outputs(6116) <= (layer0_outputs(11582)) xor (layer0_outputs(11160));
    outputs(6117) <= (layer0_outputs(11218)) xor (layer0_outputs(8346));
    outputs(6118) <= not(layer0_outputs(10993));
    outputs(6119) <= layer0_outputs(12137);
    outputs(6120) <= (layer0_outputs(12657)) and (layer0_outputs(3399));
    outputs(6121) <= not(layer0_outputs(4613)) or (layer0_outputs(3712));
    outputs(6122) <= (layer0_outputs(11076)) and (layer0_outputs(11103));
    outputs(6123) <= not((layer0_outputs(5279)) and (layer0_outputs(1037)));
    outputs(6124) <= (layer0_outputs(8559)) and not (layer0_outputs(11353));
    outputs(6125) <= not((layer0_outputs(4109)) xor (layer0_outputs(9174)));
    outputs(6126) <= (layer0_outputs(8978)) and not (layer0_outputs(9536));
    outputs(6127) <= not(layer0_outputs(9019));
    outputs(6128) <= not(layer0_outputs(4178));
    outputs(6129) <= layer0_outputs(8037);
    outputs(6130) <= not((layer0_outputs(58)) xor (layer0_outputs(12659)));
    outputs(6131) <= (layer0_outputs(10296)) and (layer0_outputs(702));
    outputs(6132) <= (layer0_outputs(3543)) and not (layer0_outputs(1601));
    outputs(6133) <= not(layer0_outputs(5829)) or (layer0_outputs(4509));
    outputs(6134) <= (layer0_outputs(347)) xor (layer0_outputs(836));
    outputs(6135) <= (layer0_outputs(6611)) and not (layer0_outputs(6006));
    outputs(6136) <= not((layer0_outputs(9605)) or (layer0_outputs(3682)));
    outputs(6137) <= not(layer0_outputs(5254));
    outputs(6138) <= not(layer0_outputs(2924)) or (layer0_outputs(5460));
    outputs(6139) <= not((layer0_outputs(10359)) xor (layer0_outputs(10358)));
    outputs(6140) <= not((layer0_outputs(9263)) or (layer0_outputs(2868)));
    outputs(6141) <= layer0_outputs(11522);
    outputs(6142) <= (layer0_outputs(12090)) and (layer0_outputs(3765));
    outputs(6143) <= not(layer0_outputs(12038));
    outputs(6144) <= (layer0_outputs(12181)) or (layer0_outputs(10459));
    outputs(6145) <= not((layer0_outputs(10801)) xor (layer0_outputs(3209)));
    outputs(6146) <= (layer0_outputs(228)) xor (layer0_outputs(4330));
    outputs(6147) <= not(layer0_outputs(5823));
    outputs(6148) <= not((layer0_outputs(7571)) xor (layer0_outputs(1845)));
    outputs(6149) <= layer0_outputs(8968);
    outputs(6150) <= layer0_outputs(2689);
    outputs(6151) <= layer0_outputs(100);
    outputs(6152) <= not((layer0_outputs(8432)) xor (layer0_outputs(3516)));
    outputs(6153) <= (layer0_outputs(9610)) and not (layer0_outputs(5282));
    outputs(6154) <= not((layer0_outputs(2168)) or (layer0_outputs(7990)));
    outputs(6155) <= not(layer0_outputs(6445));
    outputs(6156) <= not((layer0_outputs(9921)) or (layer0_outputs(3774)));
    outputs(6157) <= (layer0_outputs(5394)) and (layer0_outputs(8966));
    outputs(6158) <= not(layer0_outputs(5918));
    outputs(6159) <= (layer0_outputs(9920)) and not (layer0_outputs(3391));
    outputs(6160) <= (layer0_outputs(4519)) and not (layer0_outputs(12566));
    outputs(6161) <= layer0_outputs(7772);
    outputs(6162) <= not(layer0_outputs(7314));
    outputs(6163) <= (layer0_outputs(6983)) xor (layer0_outputs(9206));
    outputs(6164) <= (layer0_outputs(8765)) xor (layer0_outputs(9602));
    outputs(6165) <= (layer0_outputs(2813)) and (layer0_outputs(7823));
    outputs(6166) <= not((layer0_outputs(11682)) xor (layer0_outputs(11475)));
    outputs(6167) <= not(layer0_outputs(631));
    outputs(6168) <= (layer0_outputs(324)) or (layer0_outputs(11766));
    outputs(6169) <= layer0_outputs(11333);
    outputs(6170) <= not(layer0_outputs(2678));
    outputs(6171) <= not(layer0_outputs(1124));
    outputs(6172) <= not(layer0_outputs(1986)) or (layer0_outputs(11423));
    outputs(6173) <= (layer0_outputs(2579)) xor (layer0_outputs(2175));
    outputs(6174) <= layer0_outputs(10612);
    outputs(6175) <= (layer0_outputs(4871)) and not (layer0_outputs(10499));
    outputs(6176) <= not(layer0_outputs(530)) or (layer0_outputs(2337));
    outputs(6177) <= not(layer0_outputs(5691));
    outputs(6178) <= not(layer0_outputs(5864));
    outputs(6179) <= layer0_outputs(9641);
    outputs(6180) <= layer0_outputs(8864);
    outputs(6181) <= layer0_outputs(1757);
    outputs(6182) <= not((layer0_outputs(791)) and (layer0_outputs(8681)));
    outputs(6183) <= layer0_outputs(1131);
    outputs(6184) <= (layer0_outputs(7132)) and not (layer0_outputs(2416));
    outputs(6185) <= (layer0_outputs(1350)) and not (layer0_outputs(833));
    outputs(6186) <= not(layer0_outputs(1278)) or (layer0_outputs(432));
    outputs(6187) <= (layer0_outputs(3686)) xor (layer0_outputs(6142));
    outputs(6188) <= (layer0_outputs(6008)) and (layer0_outputs(9023));
    outputs(6189) <= (layer0_outputs(814)) xor (layer0_outputs(8160));
    outputs(6190) <= layer0_outputs(6352);
    outputs(6191) <= layer0_outputs(4862);
    outputs(6192) <= (layer0_outputs(9363)) xor (layer0_outputs(9331));
    outputs(6193) <= '0';
    outputs(6194) <= not((layer0_outputs(12633)) or (layer0_outputs(10648)));
    outputs(6195) <= not(layer0_outputs(9562));
    outputs(6196) <= not((layer0_outputs(6209)) or (layer0_outputs(1786)));
    outputs(6197) <= (layer0_outputs(7026)) and not (layer0_outputs(7269));
    outputs(6198) <= not(layer0_outputs(1506));
    outputs(6199) <= (layer0_outputs(3230)) and not (layer0_outputs(561));
    outputs(6200) <= layer0_outputs(11592);
    outputs(6201) <= layer0_outputs(11678);
    outputs(6202) <= not((layer0_outputs(2354)) xor (layer0_outputs(6714)));
    outputs(6203) <= layer0_outputs(5204);
    outputs(6204) <= (layer0_outputs(2353)) and (layer0_outputs(1853));
    outputs(6205) <= layer0_outputs(4902);
    outputs(6206) <= not(layer0_outputs(8997));
    outputs(6207) <= not(layer0_outputs(12199));
    outputs(6208) <= not((layer0_outputs(1733)) xor (layer0_outputs(1152)));
    outputs(6209) <= (layer0_outputs(7188)) and not (layer0_outputs(7252));
    outputs(6210) <= (layer0_outputs(5873)) and (layer0_outputs(4489));
    outputs(6211) <= layer0_outputs(1373);
    outputs(6212) <= not(layer0_outputs(2509));
    outputs(6213) <= (layer0_outputs(7142)) xor (layer0_outputs(11675));
    outputs(6214) <= not(layer0_outputs(5146));
    outputs(6215) <= layer0_outputs(5470);
    outputs(6216) <= layer0_outputs(1357);
    outputs(6217) <= (layer0_outputs(11713)) xor (layer0_outputs(6053));
    outputs(6218) <= layer0_outputs(650);
    outputs(6219) <= not(layer0_outputs(1004));
    outputs(6220) <= not((layer0_outputs(6665)) xor (layer0_outputs(8613)));
    outputs(6221) <= not(layer0_outputs(5257));
    outputs(6222) <= (layer0_outputs(6624)) and not (layer0_outputs(2304));
    outputs(6223) <= (layer0_outputs(9997)) and not (layer0_outputs(11943));
    outputs(6224) <= (layer0_outputs(11080)) and not (layer0_outputs(3850));
    outputs(6225) <= not((layer0_outputs(4366)) or (layer0_outputs(6604)));
    outputs(6226) <= (layer0_outputs(4605)) xor (layer0_outputs(10991));
    outputs(6227) <= (layer0_outputs(6228)) and (layer0_outputs(6232));
    outputs(6228) <= (layer0_outputs(12145)) xor (layer0_outputs(6850));
    outputs(6229) <= (layer0_outputs(4975)) xor (layer0_outputs(2346));
    outputs(6230) <= not((layer0_outputs(9984)) xor (layer0_outputs(3888)));
    outputs(6231) <= (layer0_outputs(10110)) or (layer0_outputs(2136));
    outputs(6232) <= (layer0_outputs(5997)) and (layer0_outputs(10260));
    outputs(6233) <= layer0_outputs(10969);
    outputs(6234) <= (layer0_outputs(7602)) and not (layer0_outputs(7318));
    outputs(6235) <= (layer0_outputs(9480)) and not (layer0_outputs(866));
    outputs(6236) <= layer0_outputs(4428);
    outputs(6237) <= (layer0_outputs(5292)) xor (layer0_outputs(7751));
    outputs(6238) <= layer0_outputs(5065);
    outputs(6239) <= not((layer0_outputs(5055)) xor (layer0_outputs(11987)));
    outputs(6240) <= not(layer0_outputs(1814));
    outputs(6241) <= layer0_outputs(8493);
    outputs(6242) <= not(layer0_outputs(5588));
    outputs(6243) <= not(layer0_outputs(9338));
    outputs(6244) <= (layer0_outputs(2162)) xor (layer0_outputs(4954));
    outputs(6245) <= not(layer0_outputs(5293));
    outputs(6246) <= not((layer0_outputs(2352)) or (layer0_outputs(11185)));
    outputs(6247) <= (layer0_outputs(12128)) xor (layer0_outputs(10882));
    outputs(6248) <= layer0_outputs(12279);
    outputs(6249) <= layer0_outputs(4134);
    outputs(6250) <= not((layer0_outputs(10191)) and (layer0_outputs(4690)));
    outputs(6251) <= layer0_outputs(7049);
    outputs(6252) <= (layer0_outputs(9948)) xor (layer0_outputs(9539));
    outputs(6253) <= not(layer0_outputs(5795));
    outputs(6254) <= not((layer0_outputs(9745)) xor (layer0_outputs(929)));
    outputs(6255) <= not(layer0_outputs(8550));
    outputs(6256) <= (layer0_outputs(12535)) xor (layer0_outputs(887));
    outputs(6257) <= layer0_outputs(4707);
    outputs(6258) <= not((layer0_outputs(8900)) xor (layer0_outputs(10630)));
    outputs(6259) <= layer0_outputs(6166);
    outputs(6260) <= not(layer0_outputs(6517));
    outputs(6261) <= layer0_outputs(8);
    outputs(6262) <= not(layer0_outputs(2050));
    outputs(6263) <= (layer0_outputs(1780)) and (layer0_outputs(6641));
    outputs(6264) <= (layer0_outputs(10092)) and not (layer0_outputs(8718));
    outputs(6265) <= not((layer0_outputs(6107)) xor (layer0_outputs(9693)));
    outputs(6266) <= (layer0_outputs(7844)) and not (layer0_outputs(11069));
    outputs(6267) <= not((layer0_outputs(9465)) or (layer0_outputs(12582)));
    outputs(6268) <= not(layer0_outputs(6707));
    outputs(6269) <= not(layer0_outputs(8858));
    outputs(6270) <= not((layer0_outputs(2448)) xor (layer0_outputs(3684)));
    outputs(6271) <= not((layer0_outputs(9043)) or (layer0_outputs(2184)));
    outputs(6272) <= not(layer0_outputs(9111));
    outputs(6273) <= not(layer0_outputs(3118));
    outputs(6274) <= (layer0_outputs(744)) and not (layer0_outputs(4691));
    outputs(6275) <= (layer0_outputs(2635)) and (layer0_outputs(10878));
    outputs(6276) <= not((layer0_outputs(2851)) xor (layer0_outputs(4794)));
    outputs(6277) <= not(layer0_outputs(6021));
    outputs(6278) <= not(layer0_outputs(7692));
    outputs(6279) <= not((layer0_outputs(12414)) xor (layer0_outputs(3316)));
    outputs(6280) <= layer0_outputs(12355);
    outputs(6281) <= not((layer0_outputs(10967)) xor (layer0_outputs(2013)));
    outputs(6282) <= not((layer0_outputs(2003)) xor (layer0_outputs(11469)));
    outputs(6283) <= not(layer0_outputs(10718));
    outputs(6284) <= not(layer0_outputs(6218));
    outputs(6285) <= (layer0_outputs(5742)) and (layer0_outputs(5017));
    outputs(6286) <= layer0_outputs(574);
    outputs(6287) <= not(layer0_outputs(11417));
    outputs(6288) <= not((layer0_outputs(2225)) or (layer0_outputs(9491)));
    outputs(6289) <= (layer0_outputs(3268)) and (layer0_outputs(2619));
    outputs(6290) <= layer0_outputs(596);
    outputs(6291) <= (layer0_outputs(12518)) xor (layer0_outputs(4314));
    outputs(6292) <= (layer0_outputs(3488)) and not (layer0_outputs(7514));
    outputs(6293) <= not((layer0_outputs(8466)) xor (layer0_outputs(797)));
    outputs(6294) <= not((layer0_outputs(12083)) xor (layer0_outputs(6455)));
    outputs(6295) <= '0';
    outputs(6296) <= (layer0_outputs(8509)) xor (layer0_outputs(9197));
    outputs(6297) <= (layer0_outputs(3855)) xor (layer0_outputs(10422));
    outputs(6298) <= not((layer0_outputs(8930)) xor (layer0_outputs(10189)));
    outputs(6299) <= not((layer0_outputs(7872)) and (layer0_outputs(3285)));
    outputs(6300) <= not((layer0_outputs(10921)) xor (layer0_outputs(3487)));
    outputs(6301) <= not((layer0_outputs(260)) or (layer0_outputs(8507)));
    outputs(6302) <= not(layer0_outputs(7443));
    outputs(6303) <= (layer0_outputs(7357)) and not (layer0_outputs(2623));
    outputs(6304) <= not((layer0_outputs(10471)) or (layer0_outputs(5880)));
    outputs(6305) <= (layer0_outputs(5998)) and not (layer0_outputs(4779));
    outputs(6306) <= (layer0_outputs(8039)) xor (layer0_outputs(1675));
    outputs(6307) <= layer0_outputs(6955);
    outputs(6308) <= not(layer0_outputs(9818));
    outputs(6309) <= not((layer0_outputs(11721)) or (layer0_outputs(8666)));
    outputs(6310) <= not((layer0_outputs(12741)) xor (layer0_outputs(8566)));
    outputs(6311) <= not(layer0_outputs(895));
    outputs(6312) <= layer0_outputs(6640);
    outputs(6313) <= (layer0_outputs(10342)) and (layer0_outputs(7215));
    outputs(6314) <= (layer0_outputs(1031)) and not (layer0_outputs(4589));
    outputs(6315) <= not(layer0_outputs(5874));
    outputs(6316) <= (layer0_outputs(155)) and not (layer0_outputs(5621));
    outputs(6317) <= (layer0_outputs(164)) and not (layer0_outputs(12084));
    outputs(6318) <= (layer0_outputs(7256)) or (layer0_outputs(10874));
    outputs(6319) <= not((layer0_outputs(8036)) xor (layer0_outputs(811)));
    outputs(6320) <= not(layer0_outputs(4013));
    outputs(6321) <= (layer0_outputs(9556)) and (layer0_outputs(11821));
    outputs(6322) <= (layer0_outputs(6584)) and (layer0_outputs(774));
    outputs(6323) <= (layer0_outputs(12164)) xor (layer0_outputs(10720));
    outputs(6324) <= not(layer0_outputs(3781));
    outputs(6325) <= layer0_outputs(11901);
    outputs(6326) <= (layer0_outputs(3956)) and (layer0_outputs(6234));
    outputs(6327) <= not((layer0_outputs(6268)) and (layer0_outputs(10906)));
    outputs(6328) <= not(layer0_outputs(12796));
    outputs(6329) <= not((layer0_outputs(2593)) xor (layer0_outputs(4798)));
    outputs(6330) <= layer0_outputs(11180);
    outputs(6331) <= (layer0_outputs(7938)) and not (layer0_outputs(7747));
    outputs(6332) <= layer0_outputs(556);
    outputs(6333) <= not(layer0_outputs(4355));
    outputs(6334) <= '1';
    outputs(6335) <= (layer0_outputs(886)) and not (layer0_outputs(9777));
    outputs(6336) <= not((layer0_outputs(6910)) or (layer0_outputs(12172)));
    outputs(6337) <= (layer0_outputs(6238)) xor (layer0_outputs(10105));
    outputs(6338) <= (layer0_outputs(6415)) xor (layer0_outputs(8060));
    outputs(6339) <= (layer0_outputs(6780)) and not (layer0_outputs(6889));
    outputs(6340) <= (layer0_outputs(3556)) xor (layer0_outputs(505));
    outputs(6341) <= (layer0_outputs(4214)) or (layer0_outputs(233));
    outputs(6342) <= not((layer0_outputs(11179)) or (layer0_outputs(5238)));
    outputs(6343) <= (layer0_outputs(5291)) and not (layer0_outputs(7491));
    outputs(6344) <= (layer0_outputs(12358)) xor (layer0_outputs(3567));
    outputs(6345) <= not(layer0_outputs(6949));
    outputs(6346) <= not(layer0_outputs(1872));
    outputs(6347) <= (layer0_outputs(11026)) and not (layer0_outputs(18));
    outputs(6348) <= (layer0_outputs(7035)) xor (layer0_outputs(8827));
    outputs(6349) <= not(layer0_outputs(8357));
    outputs(6350) <= not((layer0_outputs(2264)) and (layer0_outputs(3650)));
    outputs(6351) <= not((layer0_outputs(11376)) xor (layer0_outputs(3115)));
    outputs(6352) <= (layer0_outputs(11068)) xor (layer0_outputs(6476));
    outputs(6353) <= layer0_outputs(11701);
    outputs(6354) <= not((layer0_outputs(752)) xor (layer0_outputs(8822)));
    outputs(6355) <= not(layer0_outputs(4310)) or (layer0_outputs(9102));
    outputs(6356) <= not(layer0_outputs(1169));
    outputs(6357) <= (layer0_outputs(2324)) xor (layer0_outputs(9940));
    outputs(6358) <= layer0_outputs(2197);
    outputs(6359) <= (layer0_outputs(2564)) and not (layer0_outputs(10915));
    outputs(6360) <= layer0_outputs(11675);
    outputs(6361) <= layer0_outputs(4784);
    outputs(6362) <= (layer0_outputs(10092)) and not (layer0_outputs(6661));
    outputs(6363) <= (layer0_outputs(9926)) xor (layer0_outputs(7826));
    outputs(6364) <= not((layer0_outputs(8339)) or (layer0_outputs(12443)));
    outputs(6365) <= not((layer0_outputs(12553)) xor (layer0_outputs(3570)));
    outputs(6366) <= layer0_outputs(8625);
    outputs(6367) <= (layer0_outputs(2975)) and not (layer0_outputs(6847));
    outputs(6368) <= layer0_outputs(10891);
    outputs(6369) <= (layer0_outputs(12143)) and not (layer0_outputs(5399));
    outputs(6370) <= not(layer0_outputs(2764));
    outputs(6371) <= not((layer0_outputs(9722)) and (layer0_outputs(1865)));
    outputs(6372) <= layer0_outputs(3810);
    outputs(6373) <= (layer0_outputs(9566)) xor (layer0_outputs(9774));
    outputs(6374) <= (layer0_outputs(10673)) and not (layer0_outputs(7240));
    outputs(6375) <= layer0_outputs(128);
    outputs(6376) <= not(layer0_outputs(1262));
    outputs(6377) <= (layer0_outputs(2149)) and (layer0_outputs(1580));
    outputs(6378) <= (layer0_outputs(11548)) and (layer0_outputs(401));
    outputs(6379) <= not((layer0_outputs(10157)) and (layer0_outputs(132)));
    outputs(6380) <= not((layer0_outputs(1082)) or (layer0_outputs(8531)));
    outputs(6381) <= not(layer0_outputs(12222));
    outputs(6382) <= not(layer0_outputs(6768)) or (layer0_outputs(913));
    outputs(6383) <= (layer0_outputs(9833)) and (layer0_outputs(335));
    outputs(6384) <= not((layer0_outputs(1578)) xor (layer0_outputs(3033)));
    outputs(6385) <= (layer0_outputs(3918)) xor (layer0_outputs(8528));
    outputs(6386) <= (layer0_outputs(11904)) xor (layer0_outputs(5587));
    outputs(6387) <= layer0_outputs(1725);
    outputs(6388) <= not((layer0_outputs(2886)) xor (layer0_outputs(4444)));
    outputs(6389) <= (layer0_outputs(10495)) and (layer0_outputs(11061));
    outputs(6390) <= (layer0_outputs(11918)) and (layer0_outputs(7666));
    outputs(6391) <= not(layer0_outputs(6299));
    outputs(6392) <= not(layer0_outputs(12725));
    outputs(6393) <= '0';
    outputs(6394) <= not(layer0_outputs(9440));
    outputs(6395) <= (layer0_outputs(7300)) and not (layer0_outputs(8627));
    outputs(6396) <= layer0_outputs(5272);
    outputs(6397) <= not((layer0_outputs(4594)) xor (layer0_outputs(5833)));
    outputs(6398) <= not((layer0_outputs(5853)) and (layer0_outputs(3561)));
    outputs(6399) <= (layer0_outputs(8828)) and not (layer0_outputs(8114));
    outputs(6400) <= not(layer0_outputs(4066)) or (layer0_outputs(11480));
    outputs(6401) <= not((layer0_outputs(7734)) xor (layer0_outputs(6659)));
    outputs(6402) <= layer0_outputs(11171);
    outputs(6403) <= not(layer0_outputs(3342)) or (layer0_outputs(1689));
    outputs(6404) <= layer0_outputs(2338);
    outputs(6405) <= not(layer0_outputs(4427));
    outputs(6406) <= (layer0_outputs(10697)) and (layer0_outputs(10634));
    outputs(6407) <= (layer0_outputs(2656)) xor (layer0_outputs(3966));
    outputs(6408) <= layer0_outputs(12544);
    outputs(6409) <= (layer0_outputs(9047)) and not (layer0_outputs(11377));
    outputs(6410) <= (layer0_outputs(10361)) or (layer0_outputs(655));
    outputs(6411) <= not(layer0_outputs(7358)) or (layer0_outputs(753));
    outputs(6412) <= not(layer0_outputs(11248));
    outputs(6413) <= layer0_outputs(8631);
    outputs(6414) <= not(layer0_outputs(9665));
    outputs(6415) <= layer0_outputs(7669);
    outputs(6416) <= not((layer0_outputs(10771)) and (layer0_outputs(3136)));
    outputs(6417) <= not(layer0_outputs(7013));
    outputs(6418) <= not(layer0_outputs(11044));
    outputs(6419) <= not(layer0_outputs(7165));
    outputs(6420) <= not(layer0_outputs(758));
    outputs(6421) <= not(layer0_outputs(5));
    outputs(6422) <= (layer0_outputs(7623)) xor (layer0_outputs(7608));
    outputs(6423) <= layer0_outputs(10670);
    outputs(6424) <= (layer0_outputs(11534)) xor (layer0_outputs(1542));
    outputs(6425) <= (layer0_outputs(12008)) or (layer0_outputs(3451));
    outputs(6426) <= not(layer0_outputs(6490)) or (layer0_outputs(1611));
    outputs(6427) <= (layer0_outputs(5426)) xor (layer0_outputs(6973));
    outputs(6428) <= (layer0_outputs(2410)) xor (layer0_outputs(11274));
    outputs(6429) <= (layer0_outputs(8113)) xor (layer0_outputs(8915));
    outputs(6430) <= layer0_outputs(3227);
    outputs(6431) <= layer0_outputs(10267);
    outputs(6432) <= not((layer0_outputs(10282)) xor (layer0_outputs(10976)));
    outputs(6433) <= (layer0_outputs(5556)) and (layer0_outputs(9944));
    outputs(6434) <= (layer0_outputs(503)) xor (layer0_outputs(5028));
    outputs(6435) <= (layer0_outputs(12518)) xor (layer0_outputs(6786));
    outputs(6436) <= not((layer0_outputs(2580)) xor (layer0_outputs(2879)));
    outputs(6437) <= not((layer0_outputs(9275)) xor (layer0_outputs(12464)));
    outputs(6438) <= layer0_outputs(5134);
    outputs(6439) <= layer0_outputs(12197);
    outputs(6440) <= layer0_outputs(5882);
    outputs(6441) <= layer0_outputs(8529);
    outputs(6442) <= (layer0_outputs(9604)) xor (layer0_outputs(10603));
    outputs(6443) <= layer0_outputs(12510);
    outputs(6444) <= not(layer0_outputs(2558));
    outputs(6445) <= layer0_outputs(5608);
    outputs(6446) <= not(layer0_outputs(7605));
    outputs(6447) <= not(layer0_outputs(1890));
    outputs(6448) <= not((layer0_outputs(3852)) xor (layer0_outputs(2810)));
    outputs(6449) <= layer0_outputs(6300);
    outputs(6450) <= not(layer0_outputs(2780));
    outputs(6451) <= not(layer0_outputs(6326));
    outputs(6452) <= not(layer0_outputs(5409));
    outputs(6453) <= not((layer0_outputs(9770)) xor (layer0_outputs(10542)));
    outputs(6454) <= layer0_outputs(3500);
    outputs(6455) <= not((layer0_outputs(4217)) or (layer0_outputs(2544)));
    outputs(6456) <= (layer0_outputs(9316)) and (layer0_outputs(10466));
    outputs(6457) <= layer0_outputs(1081);
    outputs(6458) <= not((layer0_outputs(11197)) xor (layer0_outputs(8515)));
    outputs(6459) <= layer0_outputs(2252);
    outputs(6460) <= (layer0_outputs(4006)) xor (layer0_outputs(9428));
    outputs(6461) <= (layer0_outputs(9308)) and not (layer0_outputs(5140));
    outputs(6462) <= not((layer0_outputs(5136)) and (layer0_outputs(11257)));
    outputs(6463) <= (layer0_outputs(6337)) or (layer0_outputs(5519));
    outputs(6464) <= layer0_outputs(11889);
    outputs(6465) <= layer0_outputs(1728);
    outputs(6466) <= (layer0_outputs(11449)) and (layer0_outputs(9916));
    outputs(6467) <= (layer0_outputs(10595)) and not (layer0_outputs(5343));
    outputs(6468) <= not((layer0_outputs(6968)) or (layer0_outputs(10855)));
    outputs(6469) <= not((layer0_outputs(4637)) xor (layer0_outputs(4099)));
    outputs(6470) <= not(layer0_outputs(3484));
    outputs(6471) <= (layer0_outputs(6193)) and not (layer0_outputs(6652));
    outputs(6472) <= (layer0_outputs(2632)) or (layer0_outputs(2554));
    outputs(6473) <= (layer0_outputs(8570)) and not (layer0_outputs(4664));
    outputs(6474) <= not((layer0_outputs(2209)) xor (layer0_outputs(3283)));
    outputs(6475) <= not((layer0_outputs(2316)) xor (layer0_outputs(9425)));
    outputs(6476) <= not((layer0_outputs(9405)) xor (layer0_outputs(11449)));
    outputs(6477) <= layer0_outputs(5317);
    outputs(6478) <= not(layer0_outputs(8736)) or (layer0_outputs(11019));
    outputs(6479) <= not(layer0_outputs(6066));
    outputs(6480) <= (layer0_outputs(3901)) xor (layer0_outputs(11664));
    outputs(6481) <= layer0_outputs(5341);
    outputs(6482) <= not((layer0_outputs(7718)) xor (layer0_outputs(11083)));
    outputs(6483) <= not((layer0_outputs(7220)) xor (layer0_outputs(2386)));
    outputs(6484) <= not(layer0_outputs(10664));
    outputs(6485) <= not((layer0_outputs(1289)) or (layer0_outputs(10314)));
    outputs(6486) <= (layer0_outputs(11379)) and not (layer0_outputs(8284));
    outputs(6487) <= layer0_outputs(9693);
    outputs(6488) <= not(layer0_outputs(8688));
    outputs(6489) <= (layer0_outputs(555)) xor (layer0_outputs(7945));
    outputs(6490) <= (layer0_outputs(407)) xor (layer0_outputs(3048));
    outputs(6491) <= not(layer0_outputs(1338));
    outputs(6492) <= not(layer0_outputs(12234)) or (layer0_outputs(1726));
    outputs(6493) <= layer0_outputs(9975);
    outputs(6494) <= (layer0_outputs(7512)) xor (layer0_outputs(1215));
    outputs(6495) <= not(layer0_outputs(12314));
    outputs(6496) <= not(layer0_outputs(818));
    outputs(6497) <= layer0_outputs(1518);
    outputs(6498) <= (layer0_outputs(457)) and not (layer0_outputs(6092));
    outputs(6499) <= not((layer0_outputs(11238)) and (layer0_outputs(8596)));
    outputs(6500) <= not((layer0_outputs(9995)) xor (layer0_outputs(4696)));
    outputs(6501) <= (layer0_outputs(6060)) xor (layer0_outputs(6884));
    outputs(6502) <= (layer0_outputs(12667)) xor (layer0_outputs(7775));
    outputs(6503) <= not((layer0_outputs(253)) xor (layer0_outputs(5973)));
    outputs(6504) <= not(layer0_outputs(8184));
    outputs(6505) <= not((layer0_outputs(4920)) xor (layer0_outputs(651)));
    outputs(6506) <= not((layer0_outputs(7947)) xor (layer0_outputs(662)));
    outputs(6507) <= (layer0_outputs(7261)) xor (layer0_outputs(5821));
    outputs(6508) <= not(layer0_outputs(9773));
    outputs(6509) <= '1';
    outputs(6510) <= layer0_outputs(3278);
    outputs(6511) <= (layer0_outputs(11115)) and not (layer0_outputs(1323));
    outputs(6512) <= '1';
    outputs(6513) <= not(layer0_outputs(4026));
    outputs(6514) <= layer0_outputs(3750);
    outputs(6515) <= layer0_outputs(8394);
    outputs(6516) <= not((layer0_outputs(10413)) xor (layer0_outputs(7389)));
    outputs(6517) <= layer0_outputs(3065);
    outputs(6518) <= layer0_outputs(615);
    outputs(6519) <= not((layer0_outputs(2307)) xor (layer0_outputs(4184)));
    outputs(6520) <= (layer0_outputs(7077)) or (layer0_outputs(2721));
    outputs(6521) <= layer0_outputs(2731);
    outputs(6522) <= layer0_outputs(10117);
    outputs(6523) <= not(layer0_outputs(11828));
    outputs(6524) <= not(layer0_outputs(234));
    outputs(6525) <= not((layer0_outputs(1254)) or (layer0_outputs(10181)));
    outputs(6526) <= layer0_outputs(11122);
    outputs(6527) <= (layer0_outputs(9613)) xor (layer0_outputs(6809));
    outputs(6528) <= not(layer0_outputs(6368)) or (layer0_outputs(10089));
    outputs(6529) <= not((layer0_outputs(2121)) xor (layer0_outputs(8560)));
    outputs(6530) <= not(layer0_outputs(9638));
    outputs(6531) <= not(layer0_outputs(3267)) or (layer0_outputs(10560));
    outputs(6532) <= not((layer0_outputs(2439)) and (layer0_outputs(1257)));
    outputs(6533) <= not((layer0_outputs(5071)) xor (layer0_outputs(1198)));
    outputs(6534) <= not((layer0_outputs(11027)) xor (layer0_outputs(11441)));
    outputs(6535) <= not(layer0_outputs(1695));
    outputs(6536) <= not((layer0_outputs(6630)) xor (layer0_outputs(5689)));
    outputs(6537) <= layer0_outputs(6501);
    outputs(6538) <= not(layer0_outputs(4825));
    outputs(6539) <= not(layer0_outputs(6679));
    outputs(6540) <= (layer0_outputs(5948)) and not (layer0_outputs(8772));
    outputs(6541) <= not(layer0_outputs(8082)) or (layer0_outputs(3739));
    outputs(6542) <= not((layer0_outputs(10494)) xor (layer0_outputs(4245)));
    outputs(6543) <= not((layer0_outputs(1205)) xor (layer0_outputs(4834)));
    outputs(6544) <= (layer0_outputs(7638)) or (layer0_outputs(2192));
    outputs(6545) <= not(layer0_outputs(2744));
    outputs(6546) <= (layer0_outputs(3860)) and not (layer0_outputs(9126));
    outputs(6547) <= not((layer0_outputs(11152)) xor (layer0_outputs(10877)));
    outputs(6548) <= (layer0_outputs(10700)) or (layer0_outputs(2965));
    outputs(6549) <= (layer0_outputs(3368)) xor (layer0_outputs(4868));
    outputs(6550) <= (layer0_outputs(1470)) and not (layer0_outputs(8142));
    outputs(6551) <= (layer0_outputs(3722)) xor (layer0_outputs(3784));
    outputs(6552) <= layer0_outputs(8685);
    outputs(6553) <= not((layer0_outputs(528)) or (layer0_outputs(12256)));
    outputs(6554) <= not((layer0_outputs(3445)) xor (layer0_outputs(4645)));
    outputs(6555) <= layer0_outputs(2806);
    outputs(6556) <= layer0_outputs(3319);
    outputs(6557) <= (layer0_outputs(1881)) and (layer0_outputs(821));
    outputs(6558) <= (layer0_outputs(2395)) xor (layer0_outputs(5861));
    outputs(6559) <= layer0_outputs(5202);
    outputs(6560) <= layer0_outputs(6240);
    outputs(6561) <= not((layer0_outputs(5530)) xor (layer0_outputs(7605)));
    outputs(6562) <= (layer0_outputs(11176)) and not (layer0_outputs(11226));
    outputs(6563) <= (layer0_outputs(11201)) and (layer0_outputs(10577));
    outputs(6564) <= not((layer0_outputs(11785)) xor (layer0_outputs(4329)));
    outputs(6565) <= (layer0_outputs(10977)) or (layer0_outputs(7985));
    outputs(6566) <= (layer0_outputs(4047)) xor (layer0_outputs(2994));
    outputs(6567) <= not(layer0_outputs(4453));
    outputs(6568) <= '0';
    outputs(6569) <= not(layer0_outputs(7554)) or (layer0_outputs(12043));
    outputs(6570) <= layer0_outputs(5467);
    outputs(6571) <= layer0_outputs(10316);
    outputs(6572) <= layer0_outputs(10412);
    outputs(6573) <= layer0_outputs(6646);
    outputs(6574) <= not(layer0_outputs(6017)) or (layer0_outputs(4075));
    outputs(6575) <= (layer0_outputs(5165)) and not (layer0_outputs(1807));
    outputs(6576) <= not(layer0_outputs(7398));
    outputs(6577) <= not(layer0_outputs(5641)) or (layer0_outputs(8417));
    outputs(6578) <= not(layer0_outputs(8754));
    outputs(6579) <= not(layer0_outputs(2669));
    outputs(6580) <= (layer0_outputs(6097)) xor (layer0_outputs(7213));
    outputs(6581) <= not(layer0_outputs(6673));
    outputs(6582) <= layer0_outputs(8501);
    outputs(6583) <= not((layer0_outputs(7920)) xor (layer0_outputs(4377)));
    outputs(6584) <= not(layer0_outputs(3731));
    outputs(6585) <= layer0_outputs(7201);
    outputs(6586) <= layer0_outputs(539);
    outputs(6587) <= layer0_outputs(8631);
    outputs(6588) <= not(layer0_outputs(12634));
    outputs(6589) <= layer0_outputs(2459);
    outputs(6590) <= (layer0_outputs(5867)) xor (layer0_outputs(1424));
    outputs(6591) <= (layer0_outputs(12249)) xor (layer0_outputs(5173));
    outputs(6592) <= (layer0_outputs(6002)) xor (layer0_outputs(7811));
    outputs(6593) <= layer0_outputs(9374);
    outputs(6594) <= layer0_outputs(9462);
    outputs(6595) <= (layer0_outputs(3071)) xor (layer0_outputs(10886));
    outputs(6596) <= not((layer0_outputs(10797)) xor (layer0_outputs(3564)));
    outputs(6597) <= layer0_outputs(6192);
    outputs(6598) <= (layer0_outputs(9985)) and (layer0_outputs(4148));
    outputs(6599) <= (layer0_outputs(7944)) and (layer0_outputs(11455));
    outputs(6600) <= (layer0_outputs(9956)) and not (layer0_outputs(11405));
    outputs(6601) <= not((layer0_outputs(11965)) xor (layer0_outputs(1406)));
    outputs(6602) <= (layer0_outputs(4847)) and not (layer0_outputs(12773));
    outputs(6603) <= not(layer0_outputs(1609));
    outputs(6604) <= layer0_outputs(10070);
    outputs(6605) <= not(layer0_outputs(11398));
    outputs(6606) <= not((layer0_outputs(6688)) xor (layer0_outputs(6742)));
    outputs(6607) <= (layer0_outputs(2347)) and (layer0_outputs(7144));
    outputs(6608) <= not(layer0_outputs(3520)) or (layer0_outputs(3712));
    outputs(6609) <= not((layer0_outputs(3462)) or (layer0_outputs(1044)));
    outputs(6610) <= layer0_outputs(9751);
    outputs(6611) <= layer0_outputs(8014);
    outputs(6612) <= '1';
    outputs(6613) <= layer0_outputs(873);
    outputs(6614) <= not((layer0_outputs(620)) xor (layer0_outputs(6727)));
    outputs(6615) <= not((layer0_outputs(9544)) and (layer0_outputs(171)));
    outputs(6616) <= not((layer0_outputs(7990)) xor (layer0_outputs(10057)));
    outputs(6617) <= not((layer0_outputs(2021)) xor (layer0_outputs(31)));
    outputs(6618) <= (layer0_outputs(5501)) xor (layer0_outputs(5214));
    outputs(6619) <= layer0_outputs(1966);
    outputs(6620) <= (layer0_outputs(5333)) or (layer0_outputs(6868));
    outputs(6621) <= layer0_outputs(9903);
    outputs(6622) <= not(layer0_outputs(10962));
    outputs(6623) <= not(layer0_outputs(1572));
    outputs(6624) <= not((layer0_outputs(7930)) and (layer0_outputs(9962)));
    outputs(6625) <= not((layer0_outputs(3730)) and (layer0_outputs(8645)));
    outputs(6626) <= (layer0_outputs(597)) xor (layer0_outputs(11485));
    outputs(6627) <= not(layer0_outputs(736)) or (layer0_outputs(2284));
    outputs(6628) <= not(layer0_outputs(11126));
    outputs(6629) <= not((layer0_outputs(4448)) xor (layer0_outputs(11097)));
    outputs(6630) <= (layer0_outputs(928)) and not (layer0_outputs(4593));
    outputs(6631) <= layer0_outputs(2239);
    outputs(6632) <= layer0_outputs(178);
    outputs(6633) <= (layer0_outputs(5180)) xor (layer0_outputs(9062));
    outputs(6634) <= layer0_outputs(8926);
    outputs(6635) <= not(layer0_outputs(10982));
    outputs(6636) <= not(layer0_outputs(9092)) or (layer0_outputs(11596));
    outputs(6637) <= (layer0_outputs(8438)) and not (layer0_outputs(10481));
    outputs(6638) <= (layer0_outputs(149)) xor (layer0_outputs(10001));
    outputs(6639) <= layer0_outputs(3282);
    outputs(6640) <= (layer0_outputs(2215)) and not (layer0_outputs(11847));
    outputs(6641) <= not(layer0_outputs(5957));
    outputs(6642) <= (layer0_outputs(9462)) and not (layer0_outputs(10874));
    outputs(6643) <= not((layer0_outputs(6935)) xor (layer0_outputs(4510)));
    outputs(6644) <= not(layer0_outputs(9334));
    outputs(6645) <= (layer0_outputs(8619)) and not (layer0_outputs(4052));
    outputs(6646) <= not((layer0_outputs(6916)) xor (layer0_outputs(12396)));
    outputs(6647) <= (layer0_outputs(6326)) xor (layer0_outputs(4595));
    outputs(6648) <= layer0_outputs(6302);
    outputs(6649) <= layer0_outputs(938);
    outputs(6650) <= not(layer0_outputs(8789)) or (layer0_outputs(3976));
    outputs(6651) <= (layer0_outputs(6836)) and not (layer0_outputs(11908));
    outputs(6652) <= not((layer0_outputs(4451)) xor (layer0_outputs(2672)));
    outputs(6653) <= not(layer0_outputs(5422));
    outputs(6654) <= not((layer0_outputs(10217)) and (layer0_outputs(8516)));
    outputs(6655) <= not(layer0_outputs(4297));
    outputs(6656) <= layer0_outputs(7125);
    outputs(6657) <= not((layer0_outputs(3643)) xor (layer0_outputs(3951)));
    outputs(6658) <= not(layer0_outputs(11778)) or (layer0_outputs(7544));
    outputs(6659) <= (layer0_outputs(8958)) xor (layer0_outputs(4065));
    outputs(6660) <= not(layer0_outputs(6987));
    outputs(6661) <= layer0_outputs(11002);
    outputs(6662) <= layer0_outputs(7331);
    outputs(6663) <= layer0_outputs(4781);
    outputs(6664) <= (layer0_outputs(11647)) xor (layer0_outputs(6044));
    outputs(6665) <= (layer0_outputs(5943)) xor (layer0_outputs(2978));
    outputs(6666) <= layer0_outputs(987);
    outputs(6667) <= not(layer0_outputs(11604)) or (layer0_outputs(11523));
    outputs(6668) <= not((layer0_outputs(10221)) xor (layer0_outputs(3757)));
    outputs(6669) <= not((layer0_outputs(7703)) and (layer0_outputs(1345)));
    outputs(6670) <= (layer0_outputs(3071)) or (layer0_outputs(2827));
    outputs(6671) <= not((layer0_outputs(7338)) xor (layer0_outputs(4480)));
    outputs(6672) <= (layer0_outputs(8264)) and (layer0_outputs(1820));
    outputs(6673) <= (layer0_outputs(5989)) and not (layer0_outputs(2626));
    outputs(6674) <= (layer0_outputs(4209)) xor (layer0_outputs(554));
    outputs(6675) <= (layer0_outputs(12536)) or (layer0_outputs(2903));
    outputs(6676) <= (layer0_outputs(11683)) or (layer0_outputs(11207));
    outputs(6677) <= (layer0_outputs(12578)) xor (layer0_outputs(336));
    outputs(6678) <= not(layer0_outputs(9257)) or (layer0_outputs(6692));
    outputs(6679) <= not(layer0_outputs(5059));
    outputs(6680) <= not(layer0_outputs(2050)) or (layer0_outputs(8805));
    outputs(6681) <= (layer0_outputs(10215)) xor (layer0_outputs(5694));
    outputs(6682) <= not((layer0_outputs(3661)) or (layer0_outputs(9720)));
    outputs(6683) <= not(layer0_outputs(7804));
    outputs(6684) <= not((layer0_outputs(9264)) xor (layer0_outputs(9792)));
    outputs(6685) <= not((layer0_outputs(11544)) xor (layer0_outputs(2734)));
    outputs(6686) <= not(layer0_outputs(10834));
    outputs(6687) <= layer0_outputs(9093);
    outputs(6688) <= layer0_outputs(6366);
    outputs(6689) <= (layer0_outputs(1519)) xor (layer0_outputs(11339));
    outputs(6690) <= (layer0_outputs(5322)) xor (layer0_outputs(6160));
    outputs(6691) <= not(layer0_outputs(9095)) or (layer0_outputs(1653));
    outputs(6692) <= not((layer0_outputs(4582)) xor (layer0_outputs(12700)));
    outputs(6693) <= not((layer0_outputs(1421)) xor (layer0_outputs(10746)));
    outputs(6694) <= not(layer0_outputs(9815)) or (layer0_outputs(10348));
    outputs(6695) <= not(layer0_outputs(8322)) or (layer0_outputs(5037));
    outputs(6696) <= not(layer0_outputs(12678));
    outputs(6697) <= not(layer0_outputs(3170));
    outputs(6698) <= not((layer0_outputs(2194)) xor (layer0_outputs(11032)));
    outputs(6699) <= (layer0_outputs(6740)) xor (layer0_outputs(2269));
    outputs(6700) <= not(layer0_outputs(5306));
    outputs(6701) <= not((layer0_outputs(4087)) and (layer0_outputs(3448)));
    outputs(6702) <= not((layer0_outputs(7456)) xor (layer0_outputs(6500)));
    outputs(6703) <= not(layer0_outputs(5361));
    outputs(6704) <= not((layer0_outputs(7780)) xor (layer0_outputs(9918)));
    outputs(6705) <= layer0_outputs(8791);
    outputs(6706) <= not((layer0_outputs(8917)) xor (layer0_outputs(12261)));
    outputs(6707) <= not((layer0_outputs(908)) and (layer0_outputs(10817)));
    outputs(6708) <= (layer0_outputs(7273)) and not (layer0_outputs(616));
    outputs(6709) <= layer0_outputs(2159);
    outputs(6710) <= not((layer0_outputs(10260)) xor (layer0_outputs(8793)));
    outputs(6711) <= (layer0_outputs(7488)) or (layer0_outputs(543));
    outputs(6712) <= (layer0_outputs(8804)) xor (layer0_outputs(9176));
    outputs(6713) <= (layer0_outputs(3511)) xor (layer0_outputs(6484));
    outputs(6714) <= not(layer0_outputs(1008));
    outputs(6715) <= (layer0_outputs(12146)) xor (layer0_outputs(6763));
    outputs(6716) <= (layer0_outputs(11013)) and not (layer0_outputs(479));
    outputs(6717) <= not(layer0_outputs(7034));
    outputs(6718) <= layer0_outputs(2459);
    outputs(6719) <= not((layer0_outputs(10258)) xor (layer0_outputs(331)));
    outputs(6720) <= layer0_outputs(6278);
    outputs(6721) <= not((layer0_outputs(5454)) xor (layer0_outputs(2292)));
    outputs(6722) <= layer0_outputs(9798);
    outputs(6723) <= (layer0_outputs(1040)) and not (layer0_outputs(3701));
    outputs(6724) <= not((layer0_outputs(6867)) xor (layer0_outputs(8114)));
    outputs(6725) <= (layer0_outputs(931)) and not (layer0_outputs(5851));
    outputs(6726) <= not(layer0_outputs(2556)) or (layer0_outputs(2993));
    outputs(6727) <= (layer0_outputs(286)) and not (layer0_outputs(4652));
    outputs(6728) <= (layer0_outputs(206)) and not (layer0_outputs(8652));
    outputs(6729) <= layer0_outputs(1595);
    outputs(6730) <= not(layer0_outputs(3170));
    outputs(6731) <= not((layer0_outputs(4050)) xor (layer0_outputs(2490)));
    outputs(6732) <= (layer0_outputs(928)) xor (layer0_outputs(11864));
    outputs(6733) <= (layer0_outputs(190)) xor (layer0_outputs(7367));
    outputs(6734) <= not(layer0_outputs(1633));
    outputs(6735) <= layer0_outputs(11884);
    outputs(6736) <= (layer0_outputs(5395)) xor (layer0_outputs(3005));
    outputs(6737) <= layer0_outputs(3698);
    outputs(6738) <= (layer0_outputs(10163)) xor (layer0_outputs(2258));
    outputs(6739) <= layer0_outputs(12774);
    outputs(6740) <= layer0_outputs(11502);
    outputs(6741) <= (layer0_outputs(9955)) xor (layer0_outputs(2205));
    outputs(6742) <= layer0_outputs(10173);
    outputs(6743) <= (layer0_outputs(2529)) xor (layer0_outputs(1021));
    outputs(6744) <= not(layer0_outputs(8717)) or (layer0_outputs(2853));
    outputs(6745) <= (layer0_outputs(8334)) xor (layer0_outputs(11575));
    outputs(6746) <= not((layer0_outputs(4458)) xor (layer0_outputs(4758)));
    outputs(6747) <= (layer0_outputs(10417)) and not (layer0_outputs(10905));
    outputs(6748) <= not(layer0_outputs(844));
    outputs(6749) <= not(layer0_outputs(9404));
    outputs(6750) <= layer0_outputs(733);
    outputs(6751) <= (layer0_outputs(805)) or (layer0_outputs(2309));
    outputs(6752) <= not((layer0_outputs(7197)) xor (layer0_outputs(2605)));
    outputs(6753) <= not(layer0_outputs(9333));
    outputs(6754) <= not((layer0_outputs(394)) and (layer0_outputs(3444)));
    outputs(6755) <= (layer0_outputs(1444)) and not (layer0_outputs(10059));
    outputs(6756) <= not(layer0_outputs(9142));
    outputs(6757) <= not((layer0_outputs(461)) xor (layer0_outputs(1434)));
    outputs(6758) <= not((layer0_outputs(1541)) xor (layer0_outputs(1581)));
    outputs(6759) <= layer0_outputs(7499);
    outputs(6760) <= not(layer0_outputs(8314));
    outputs(6761) <= (layer0_outputs(5419)) and not (layer0_outputs(2166));
    outputs(6762) <= (layer0_outputs(2233)) xor (layer0_outputs(8200));
    outputs(6763) <= (layer0_outputs(940)) and (layer0_outputs(8736));
    outputs(6764) <= not(layer0_outputs(201)) or (layer0_outputs(3290));
    outputs(6765) <= not(layer0_outputs(12234));
    outputs(6766) <= layer0_outputs(7996);
    outputs(6767) <= not((layer0_outputs(5357)) xor (layer0_outputs(12126)));
    outputs(6768) <= layer0_outputs(8034);
    outputs(6769) <= not((layer0_outputs(6253)) xor (layer0_outputs(12000)));
    outputs(6770) <= '0';
    outputs(6771) <= not(layer0_outputs(8327));
    outputs(6772) <= not((layer0_outputs(3348)) xor (layer0_outputs(9222)));
    outputs(6773) <= layer0_outputs(4960);
    outputs(6774) <= not((layer0_outputs(5567)) xor (layer0_outputs(3320)));
    outputs(6775) <= not(layer0_outputs(6123));
    outputs(6776) <= (layer0_outputs(1789)) xor (layer0_outputs(8485));
    outputs(6777) <= not(layer0_outputs(8392)) or (layer0_outputs(472));
    outputs(6778) <= layer0_outputs(3028);
    outputs(6779) <= not((layer0_outputs(3205)) xor (layer0_outputs(282)));
    outputs(6780) <= not((layer0_outputs(583)) and (layer0_outputs(9191)));
    outputs(6781) <= (layer0_outputs(9224)) and not (layer0_outputs(12297));
    outputs(6782) <= not(layer0_outputs(2132));
    outputs(6783) <= layer0_outputs(6434);
    outputs(6784) <= not(layer0_outputs(619)) or (layer0_outputs(7328));
    outputs(6785) <= not(layer0_outputs(10570));
    outputs(6786) <= layer0_outputs(11702);
    outputs(6787) <= '1';
    outputs(6788) <= not(layer0_outputs(6673));
    outputs(6789) <= not((layer0_outputs(555)) xor (layer0_outputs(10826)));
    outputs(6790) <= layer0_outputs(1485);
    outputs(6791) <= not((layer0_outputs(10302)) and (layer0_outputs(11551)));
    outputs(6792) <= not((layer0_outputs(3861)) xor (layer0_outputs(803)));
    outputs(6793) <= not((layer0_outputs(7599)) xor (layer0_outputs(4904)));
    outputs(6794) <= not(layer0_outputs(2768));
    outputs(6795) <= not(layer0_outputs(10006));
    outputs(6796) <= not((layer0_outputs(1711)) xor (layer0_outputs(9172)));
    outputs(6797) <= layer0_outputs(11294);
    outputs(6798) <= not(layer0_outputs(1981));
    outputs(6799) <= (layer0_outputs(4311)) xor (layer0_outputs(8254));
    outputs(6800) <= (layer0_outputs(1033)) and (layer0_outputs(3717));
    outputs(6801) <= (layer0_outputs(12055)) xor (layer0_outputs(11667));
    outputs(6802) <= layer0_outputs(5185);
    outputs(6803) <= layer0_outputs(10201);
    outputs(6804) <= not(layer0_outputs(778)) or (layer0_outputs(1918));
    outputs(6805) <= not(layer0_outputs(3574)) or (layer0_outputs(10181));
    outputs(6806) <= layer0_outputs(6290);
    outputs(6807) <= not(layer0_outputs(6798)) or (layer0_outputs(8245));
    outputs(6808) <= (layer0_outputs(10868)) and not (layer0_outputs(8499));
    outputs(6809) <= not((layer0_outputs(9419)) xor (layer0_outputs(3848)));
    outputs(6810) <= not((layer0_outputs(9164)) xor (layer0_outputs(2201)));
    outputs(6811) <= (layer0_outputs(3391)) xor (layer0_outputs(761));
    outputs(6812) <= not(layer0_outputs(1875));
    outputs(6813) <= not((layer0_outputs(2272)) xor (layer0_outputs(6974)));
    outputs(6814) <= (layer0_outputs(5744)) and not (layer0_outputs(7876));
    outputs(6815) <= not((layer0_outputs(5683)) xor (layer0_outputs(9826)));
    outputs(6816) <= (layer0_outputs(12254)) or (layer0_outputs(5054));
    outputs(6817) <= not((layer0_outputs(8496)) xor (layer0_outputs(8745)));
    outputs(6818) <= (layer0_outputs(3792)) xor (layer0_outputs(550));
    outputs(6819) <= not((layer0_outputs(12111)) and (layer0_outputs(6379)));
    outputs(6820) <= not(layer0_outputs(10946)) or (layer0_outputs(3308));
    outputs(6821) <= (layer0_outputs(6245)) and (layer0_outputs(147));
    outputs(6822) <= layer0_outputs(8089);
    outputs(6823) <= layer0_outputs(7792);
    outputs(6824) <= not(layer0_outputs(12537));
    outputs(6825) <= layer0_outputs(9392);
    outputs(6826) <= layer0_outputs(7991);
    outputs(6827) <= layer0_outputs(8836);
    outputs(6828) <= layer0_outputs(12638);
    outputs(6829) <= not(layer0_outputs(12516));
    outputs(6830) <= layer0_outputs(1386);
    outputs(6831) <= '0';
    outputs(6832) <= not((layer0_outputs(8172)) xor (layer0_outputs(8856)));
    outputs(6833) <= layer0_outputs(5934);
    outputs(6834) <= not((layer0_outputs(610)) xor (layer0_outputs(10369)));
    outputs(6835) <= layer0_outputs(3898);
    outputs(6836) <= not(layer0_outputs(6311));
    outputs(6837) <= not(layer0_outputs(7398));
    outputs(6838) <= (layer0_outputs(10184)) or (layer0_outputs(12205));
    outputs(6839) <= not(layer0_outputs(5464));
    outputs(6840) <= layer0_outputs(11962);
    outputs(6841) <= (layer0_outputs(11919)) xor (layer0_outputs(11427));
    outputs(6842) <= (layer0_outputs(7550)) xor (layer0_outputs(943));
    outputs(6843) <= not((layer0_outputs(6147)) xor (layer0_outputs(9406)));
    outputs(6844) <= not(layer0_outputs(1524)) or (layer0_outputs(10836));
    outputs(6845) <= (layer0_outputs(6158)) xor (layer0_outputs(7999));
    outputs(6846) <= (layer0_outputs(517)) xor (layer0_outputs(11570));
    outputs(6847) <= not((layer0_outputs(3930)) and (layer0_outputs(9434)));
    outputs(6848) <= not((layer0_outputs(10179)) and (layer0_outputs(1344)));
    outputs(6849) <= layer0_outputs(7353);
    outputs(6850) <= not(layer0_outputs(2143));
    outputs(6851) <= not(layer0_outputs(10280)) or (layer0_outputs(2029));
    outputs(6852) <= not(layer0_outputs(3455));
    outputs(6853) <= not(layer0_outputs(12563));
    outputs(6854) <= layer0_outputs(1010);
    outputs(6855) <= not((layer0_outputs(3857)) or (layer0_outputs(1573)));
    outputs(6856) <= '1';
    outputs(6857) <= (layer0_outputs(11669)) or (layer0_outputs(1247));
    outputs(6858) <= (layer0_outputs(9676)) xor (layer0_outputs(11047));
    outputs(6859) <= (layer0_outputs(5433)) or (layer0_outputs(6430));
    outputs(6860) <= (layer0_outputs(962)) or (layer0_outputs(3675));
    outputs(6861) <= not((layer0_outputs(7901)) xor (layer0_outputs(7860)));
    outputs(6862) <= (layer0_outputs(9646)) xor (layer0_outputs(1958));
    outputs(6863) <= (layer0_outputs(4692)) and not (layer0_outputs(6005));
    outputs(6864) <= (layer0_outputs(4420)) and (layer0_outputs(4394));
    outputs(6865) <= not((layer0_outputs(6826)) and (layer0_outputs(7284)));
    outputs(6866) <= (layer0_outputs(5493)) and not (layer0_outputs(6520));
    outputs(6867) <= not(layer0_outputs(12577)) or (layer0_outputs(5063));
    outputs(6868) <= not(layer0_outputs(11872));
    outputs(6869) <= not((layer0_outputs(8525)) xor (layer0_outputs(587)));
    outputs(6870) <= not((layer0_outputs(3218)) xor (layer0_outputs(4340)));
    outputs(6871) <= layer0_outputs(9513);
    outputs(6872) <= not((layer0_outputs(10957)) xor (layer0_outputs(140)));
    outputs(6873) <= not(layer0_outputs(1217)) or (layer0_outputs(523));
    outputs(6874) <= not((layer0_outputs(6716)) or (layer0_outputs(10418)));
    outputs(6875) <= not((layer0_outputs(8620)) xor (layer0_outputs(1128)));
    outputs(6876) <= (layer0_outputs(10669)) or (layer0_outputs(6114));
    outputs(6877) <= (layer0_outputs(8318)) xor (layer0_outputs(11974));
    outputs(6878) <= not(layer0_outputs(2207));
    outputs(6879) <= not(layer0_outputs(8557));
    outputs(6880) <= not(layer0_outputs(511)) or (layer0_outputs(12497));
    outputs(6881) <= not((layer0_outputs(122)) xor (layer0_outputs(10754)));
    outputs(6882) <= (layer0_outputs(10239)) xor (layer0_outputs(6120));
    outputs(6883) <= not((layer0_outputs(1140)) xor (layer0_outputs(3482)));
    outputs(6884) <= not(layer0_outputs(11128));
    outputs(6885) <= layer0_outputs(9682);
    outputs(6886) <= not(layer0_outputs(9793));
    outputs(6887) <= not(layer0_outputs(6752));
    outputs(6888) <= not((layer0_outputs(231)) xor (layer0_outputs(9925)));
    outputs(6889) <= '1';
    outputs(6890) <= (layer0_outputs(2272)) xor (layer0_outputs(5116));
    outputs(6891) <= (layer0_outputs(11774)) or (layer0_outputs(10434));
    outputs(6892) <= not((layer0_outputs(3403)) xor (layer0_outputs(2425)));
    outputs(6893) <= not(layer0_outputs(2399)) or (layer0_outputs(977));
    outputs(6894) <= (layer0_outputs(2391)) and not (layer0_outputs(3603));
    outputs(6895) <= not((layer0_outputs(8448)) or (layer0_outputs(3639)));
    outputs(6896) <= layer0_outputs(5041);
    outputs(6897) <= (layer0_outputs(10696)) xor (layer0_outputs(1069));
    outputs(6898) <= (layer0_outputs(1234)) and not (layer0_outputs(5353));
    outputs(6899) <= layer0_outputs(9657);
    outputs(6900) <= not((layer0_outputs(9489)) or (layer0_outputs(5188)));
    outputs(6901) <= not((layer0_outputs(7728)) xor (layer0_outputs(5209)));
    outputs(6902) <= (layer0_outputs(6902)) xor (layer0_outputs(11132));
    outputs(6903) <= layer0_outputs(2945);
    outputs(6904) <= (layer0_outputs(4644)) and (layer0_outputs(6415));
    outputs(6905) <= not(layer0_outputs(12346)) or (layer0_outputs(1841));
    outputs(6906) <= not(layer0_outputs(11729)) or (layer0_outputs(706));
    outputs(6907) <= layer0_outputs(7413);
    outputs(6908) <= layer0_outputs(1098);
    outputs(6909) <= not((layer0_outputs(12140)) or (layer0_outputs(3421)));
    outputs(6910) <= not(layer0_outputs(2954));
    outputs(6911) <= not(layer0_outputs(4647)) or (layer0_outputs(1827));
    outputs(6912) <= (layer0_outputs(4842)) and not (layer0_outputs(12736));
    outputs(6913) <= (layer0_outputs(10744)) and (layer0_outputs(7820));
    outputs(6914) <= (layer0_outputs(1036)) and not (layer0_outputs(5582));
    outputs(6915) <= layer0_outputs(2631);
    outputs(6916) <= not(layer0_outputs(5351));
    outputs(6917) <= not((layer0_outputs(4045)) xor (layer0_outputs(1852)));
    outputs(6918) <= (layer0_outputs(12615)) and not (layer0_outputs(3630));
    outputs(6919) <= not((layer0_outputs(6107)) xor (layer0_outputs(9854)));
    outputs(6920) <= not(layer0_outputs(6310)) or (layer0_outputs(8044));
    outputs(6921) <= '1';
    outputs(6922) <= (layer0_outputs(9187)) and (layer0_outputs(10926));
    outputs(6923) <= not((layer0_outputs(2428)) xor (layer0_outputs(11886)));
    outputs(6924) <= layer0_outputs(779);
    outputs(6925) <= (layer0_outputs(3739)) xor (layer0_outputs(7221));
    outputs(6926) <= (layer0_outputs(939)) and (layer0_outputs(582));
    outputs(6927) <= layer0_outputs(8766);
    outputs(6928) <= (layer0_outputs(4701)) and not (layer0_outputs(11198));
    outputs(6929) <= (layer0_outputs(12290)) xor (layer0_outputs(11491));
    outputs(6930) <= '0';
    outputs(6931) <= not((layer0_outputs(5548)) xor (layer0_outputs(9639)));
    outputs(6932) <= (layer0_outputs(3223)) and not (layer0_outputs(704));
    outputs(6933) <= layer0_outputs(2602);
    outputs(6934) <= not((layer0_outputs(3078)) or (layer0_outputs(1209)));
    outputs(6935) <= (layer0_outputs(8237)) or (layer0_outputs(12172));
    outputs(6936) <= not(layer0_outputs(7396));
    outputs(6937) <= not(layer0_outputs(4228)) or (layer0_outputs(9710));
    outputs(6938) <= layer0_outputs(9600);
    outputs(6939) <= not(layer0_outputs(10953));
    outputs(6940) <= not(layer0_outputs(5160)) or (layer0_outputs(4031));
    outputs(6941) <= not((layer0_outputs(6159)) xor (layer0_outputs(634)));
    outputs(6942) <= (layer0_outputs(6254)) xor (layer0_outputs(7957));
    outputs(6943) <= not(layer0_outputs(11916));
    outputs(6944) <= layer0_outputs(12220);
    outputs(6945) <= not((layer0_outputs(3460)) xor (layer0_outputs(11085)));
    outputs(6946) <= not(layer0_outputs(11185)) or (layer0_outputs(11829));
    outputs(6947) <= not(layer0_outputs(9084)) or (layer0_outputs(1354));
    outputs(6948) <= not((layer0_outputs(9891)) xor (layer0_outputs(6505)));
    outputs(6949) <= not((layer0_outputs(8707)) and (layer0_outputs(7336)));
    outputs(6950) <= not((layer0_outputs(749)) xor (layer0_outputs(10856)));
    outputs(6951) <= (layer0_outputs(11063)) and not (layer0_outputs(980));
    outputs(6952) <= not((layer0_outputs(11136)) xor (layer0_outputs(8522)));
    outputs(6953) <= not(layer0_outputs(11189));
    outputs(6954) <= (layer0_outputs(7297)) or (layer0_outputs(1697));
    outputs(6955) <= not(layer0_outputs(2384)) or (layer0_outputs(6414));
    outputs(6956) <= layer0_outputs(9467);
    outputs(6957) <= layer0_outputs(7500);
    outputs(6958) <= layer0_outputs(11763);
    outputs(6959) <= not(layer0_outputs(6801));
    outputs(6960) <= not(layer0_outputs(8191)) or (layer0_outputs(5581));
    outputs(6961) <= '1';
    outputs(6962) <= layer0_outputs(12392);
    outputs(6963) <= layer0_outputs(1505);
    outputs(6964) <= '1';
    outputs(6965) <= layer0_outputs(1844);
    outputs(6966) <= not(layer0_outputs(7608)) or (layer0_outputs(4643));
    outputs(6967) <= (layer0_outputs(7122)) xor (layer0_outputs(11380));
    outputs(6968) <= not((layer0_outputs(809)) and (layer0_outputs(10286)));
    outputs(6969) <= (layer0_outputs(10705)) or (layer0_outputs(12500));
    outputs(6970) <= not((layer0_outputs(2648)) xor (layer0_outputs(1286)));
    outputs(6971) <= layer0_outputs(6054);
    outputs(6972) <= not((layer0_outputs(5791)) xor (layer0_outputs(411)));
    outputs(6973) <= not((layer0_outputs(2530)) xor (layer0_outputs(12348)));
    outputs(6974) <= layer0_outputs(5818);
    outputs(6975) <= (layer0_outputs(4774)) and (layer0_outputs(1196));
    outputs(6976) <= not((layer0_outputs(7837)) or (layer0_outputs(2293)));
    outputs(6977) <= layer0_outputs(9411);
    outputs(6978) <= (layer0_outputs(9540)) and (layer0_outputs(7044));
    outputs(6979) <= not((layer0_outputs(9321)) xor (layer0_outputs(4503)));
    outputs(6980) <= not(layer0_outputs(4446));
    outputs(6981) <= not((layer0_outputs(8996)) xor (layer0_outputs(6173)));
    outputs(6982) <= layer0_outputs(11665);
    outputs(6983) <= layer0_outputs(2738);
    outputs(6984) <= not(layer0_outputs(4159));
    outputs(6985) <= (layer0_outputs(8546)) xor (layer0_outputs(10786));
    outputs(6986) <= layer0_outputs(12573);
    outputs(6987) <= not((layer0_outputs(11586)) xor (layer0_outputs(378)));
    outputs(6988) <= layer0_outputs(5716);
    outputs(6989) <= '1';
    outputs(6990) <= not(layer0_outputs(3092));
    outputs(6991) <= not((layer0_outputs(4297)) and (layer0_outputs(7253)));
    outputs(6992) <= not((layer0_outputs(8798)) xor (layer0_outputs(12452)));
    outputs(6993) <= (layer0_outputs(4663)) xor (layer0_outputs(8637));
    outputs(6994) <= not((layer0_outputs(6862)) xor (layer0_outputs(9295)));
    outputs(6995) <= (layer0_outputs(7244)) and (layer0_outputs(10907));
    outputs(6996) <= (layer0_outputs(4403)) xor (layer0_outputs(8999));
    outputs(6997) <= layer0_outputs(7578);
    outputs(6998) <= not((layer0_outputs(11574)) xor (layer0_outputs(10843)));
    outputs(6999) <= (layer0_outputs(446)) or (layer0_outputs(9407));
    outputs(7000) <= (layer0_outputs(1059)) xor (layer0_outputs(7982));
    outputs(7001) <= (layer0_outputs(10601)) and not (layer0_outputs(9237));
    outputs(7002) <= not((layer0_outputs(3278)) xor (layer0_outputs(9213)));
    outputs(7003) <= (layer0_outputs(3528)) and not (layer0_outputs(7903));
    outputs(7004) <= (layer0_outputs(11500)) and not (layer0_outputs(912));
    outputs(7005) <= not(layer0_outputs(8433));
    outputs(7006) <= layer0_outputs(4345);
    outputs(7007) <= layer0_outputs(615);
    outputs(7008) <= not(layer0_outputs(9347));
    outputs(7009) <= not((layer0_outputs(7636)) and (layer0_outputs(2146)));
    outputs(7010) <= not(layer0_outputs(646)) or (layer0_outputs(5016));
    outputs(7011) <= (layer0_outputs(1051)) and not (layer0_outputs(5437));
    outputs(7012) <= (layer0_outputs(5153)) xor (layer0_outputs(8903));
    outputs(7013) <= not((layer0_outputs(7752)) and (layer0_outputs(3276)));
    outputs(7014) <= (layer0_outputs(9430)) xor (layer0_outputs(10533));
    outputs(7015) <= not(layer0_outputs(11862)) or (layer0_outputs(7386));
    outputs(7016) <= not(layer0_outputs(1494)) or (layer0_outputs(5865));
    outputs(7017) <= not(layer0_outputs(3561));
    outputs(7018) <= not(layer0_outputs(10043));
    outputs(7019) <= (layer0_outputs(8745)) and (layer0_outputs(9103));
    outputs(7020) <= layer0_outputs(5230);
    outputs(7021) <= not(layer0_outputs(10124));
    outputs(7022) <= not((layer0_outputs(2477)) xor (layer0_outputs(10338)));
    outputs(7023) <= layer0_outputs(10755);
    outputs(7024) <= not((layer0_outputs(12370)) xor (layer0_outputs(5304)));
    outputs(7025) <= (layer0_outputs(10227)) and (layer0_outputs(5911));
    outputs(7026) <= layer0_outputs(11977);
    outputs(7027) <= (layer0_outputs(5061)) or (layer0_outputs(26));
    outputs(7028) <= layer0_outputs(4160);
    outputs(7029) <= layer0_outputs(11188);
    outputs(7030) <= (layer0_outputs(6294)) xor (layer0_outputs(8239));
    outputs(7031) <= not(layer0_outputs(5354));
    outputs(7032) <= not(layer0_outputs(8769)) or (layer0_outputs(10152));
    outputs(7033) <= layer0_outputs(2698);
    outputs(7034) <= (layer0_outputs(26)) and not (layer0_outputs(675));
    outputs(7035) <= layer0_outputs(6590);
    outputs(7036) <= (layer0_outputs(8753)) xor (layer0_outputs(4780));
    outputs(7037) <= (layer0_outputs(6026)) and not (layer0_outputs(4843));
    outputs(7038) <= (layer0_outputs(7415)) xor (layer0_outputs(7766));
    outputs(7039) <= not(layer0_outputs(8343)) or (layer0_outputs(8744));
    outputs(7040) <= layer0_outputs(4723);
    outputs(7041) <= not(layer0_outputs(1826));
    outputs(7042) <= not(layer0_outputs(6035));
    outputs(7043) <= (layer0_outputs(12096)) and (layer0_outputs(7063));
    outputs(7044) <= layer0_outputs(408);
    outputs(7045) <= not(layer0_outputs(11223)) or (layer0_outputs(4756));
    outputs(7046) <= (layer0_outputs(7333)) xor (layer0_outputs(9710));
    outputs(7047) <= not((layer0_outputs(3339)) and (layer0_outputs(9705)));
    outputs(7048) <= (layer0_outputs(8386)) and not (layer0_outputs(5732));
    outputs(7049) <= not(layer0_outputs(8609));
    outputs(7050) <= not(layer0_outputs(10050)) or (layer0_outputs(6796));
    outputs(7051) <= not((layer0_outputs(1273)) and (layer0_outputs(6448)));
    outputs(7052) <= layer0_outputs(12391);
    outputs(7053) <= not((layer0_outputs(12560)) and (layer0_outputs(11677)));
    outputs(7054) <= (layer0_outputs(4921)) and not (layer0_outputs(3370));
    outputs(7055) <= not(layer0_outputs(8806)) or (layer0_outputs(9936));
    outputs(7056) <= '1';
    outputs(7057) <= (layer0_outputs(7176)) or (layer0_outputs(9593));
    outputs(7058) <= (layer0_outputs(12638)) xor (layer0_outputs(9329));
    outputs(7059) <= (layer0_outputs(7880)) and not (layer0_outputs(4982));
    outputs(7060) <= (layer0_outputs(3593)) xor (layer0_outputs(6207));
    outputs(7061) <= (layer0_outputs(7636)) xor (layer0_outputs(2042));
    outputs(7062) <= layer0_outputs(9535);
    outputs(7063) <= layer0_outputs(7124);
    outputs(7064) <= (layer0_outputs(147)) xor (layer0_outputs(4124));
    outputs(7065) <= not(layer0_outputs(9142));
    outputs(7066) <= not(layer0_outputs(10530));
    outputs(7067) <= (layer0_outputs(7260)) xor (layer0_outputs(3315));
    outputs(7068) <= not(layer0_outputs(12307)) or (layer0_outputs(6868));
    outputs(7069) <= not(layer0_outputs(5734));
    outputs(7070) <= (layer0_outputs(12762)) or (layer0_outputs(7160));
    outputs(7071) <= (layer0_outputs(11588)) xor (layer0_outputs(11607));
    outputs(7072) <= not((layer0_outputs(194)) and (layer0_outputs(935)));
    outputs(7073) <= (layer0_outputs(664)) xor (layer0_outputs(6283));
    outputs(7074) <= (layer0_outputs(80)) xor (layer0_outputs(5094));
    outputs(7075) <= layer0_outputs(1450);
    outputs(7076) <= layer0_outputs(11698);
    outputs(7077) <= not((layer0_outputs(1715)) xor (layer0_outputs(9140)));
    outputs(7078) <= not(layer0_outputs(5084));
    outputs(7079) <= not(layer0_outputs(1164));
    outputs(7080) <= (layer0_outputs(5729)) and not (layer0_outputs(2628));
    outputs(7081) <= not(layer0_outputs(4390));
    outputs(7082) <= (layer0_outputs(10126)) or (layer0_outputs(11662));
    outputs(7083) <= not((layer0_outputs(10419)) xor (layer0_outputs(435)));
    outputs(7084) <= (layer0_outputs(3345)) and not (layer0_outputs(9148));
    outputs(7085) <= layer0_outputs(10099);
    outputs(7086) <= not(layer0_outputs(2765)) or (layer0_outputs(8910));
    outputs(7087) <= not(layer0_outputs(3563));
    outputs(7088) <= (layer0_outputs(4550)) xor (layer0_outputs(6647));
    outputs(7089) <= (layer0_outputs(2349)) xor (layer0_outputs(7174));
    outputs(7090) <= (layer0_outputs(5288)) xor (layer0_outputs(10562));
    outputs(7091) <= layer0_outputs(10417);
    outputs(7092) <= not(layer0_outputs(2744));
    outputs(7093) <= layer0_outputs(1765);
    outputs(7094) <= layer0_outputs(5942);
    outputs(7095) <= (layer0_outputs(5223)) xor (layer0_outputs(12143));
    outputs(7096) <= not(layer0_outputs(12331)) or (layer0_outputs(55));
    outputs(7097) <= not((layer0_outputs(11992)) xor (layer0_outputs(2096)));
    outputs(7098) <= not(layer0_outputs(6724)) or (layer0_outputs(6284));
    outputs(7099) <= not(layer0_outputs(2864));
    outputs(7100) <= not((layer0_outputs(1202)) xor (layer0_outputs(7249)));
    outputs(7101) <= (layer0_outputs(8700)) and not (layer0_outputs(12245));
    outputs(7102) <= layer0_outputs(10004);
    outputs(7103) <= not((layer0_outputs(11029)) xor (layer0_outputs(4778)));
    outputs(7104) <= layer0_outputs(4599);
    outputs(7105) <= not(layer0_outputs(9214)) or (layer0_outputs(10887));
    outputs(7106) <= layer0_outputs(3582);
    outputs(7107) <= (layer0_outputs(7685)) xor (layer0_outputs(1638));
    outputs(7108) <= not((layer0_outputs(12380)) xor (layer0_outputs(6135)));
    outputs(7109) <= (layer0_outputs(6515)) xor (layer0_outputs(9788));
    outputs(7110) <= (layer0_outputs(7265)) xor (layer0_outputs(6924));
    outputs(7111) <= not((layer0_outputs(11804)) xor (layer0_outputs(3931)));
    outputs(7112) <= not((layer0_outputs(9449)) xor (layer0_outputs(9442)));
    outputs(7113) <= not(layer0_outputs(1904)) or (layer0_outputs(2719));
    outputs(7114) <= not(layer0_outputs(2759));
    outputs(7115) <= not(layer0_outputs(2014));
    outputs(7116) <= not(layer0_outputs(3599));
    outputs(7117) <= (layer0_outputs(9589)) xor (layer0_outputs(9970));
    outputs(7118) <= (layer0_outputs(2860)) xor (layer0_outputs(662));
    outputs(7119) <= layer0_outputs(5397);
    outputs(7120) <= not((layer0_outputs(497)) xor (layer0_outputs(5014)));
    outputs(7121) <= not(layer0_outputs(4288));
    outputs(7122) <= (layer0_outputs(12763)) and (layer0_outputs(498));
    outputs(7123) <= not((layer0_outputs(3225)) xor (layer0_outputs(4450)));
    outputs(7124) <= not(layer0_outputs(6916)) or (layer0_outputs(10194));
    outputs(7125) <= not((layer0_outputs(11330)) xor (layer0_outputs(1401)));
    outputs(7126) <= not(layer0_outputs(7800));
    outputs(7127) <= (layer0_outputs(4614)) xor (layer0_outputs(2820));
    outputs(7128) <= (layer0_outputs(10976)) xor (layer0_outputs(1055));
    outputs(7129) <= (layer0_outputs(3514)) or (layer0_outputs(4359));
    outputs(7130) <= layer0_outputs(7729);
    outputs(7131) <= not(layer0_outputs(8433));
    outputs(7132) <= not(layer0_outputs(5701));
    outputs(7133) <= (layer0_outputs(5808)) and (layer0_outputs(1092));
    outputs(7134) <= not(layer0_outputs(6266));
    outputs(7135) <= layer0_outputs(350);
    outputs(7136) <= not((layer0_outputs(7719)) or (layer0_outputs(1004)));
    outputs(7137) <= not((layer0_outputs(6535)) and (layer0_outputs(3736)));
    outputs(7138) <= layer0_outputs(10126);
    outputs(7139) <= (layer0_outputs(3729)) xor (layer0_outputs(10751));
    outputs(7140) <= not((layer0_outputs(4139)) and (layer0_outputs(2588)));
    outputs(7141) <= (layer0_outputs(8222)) or (layer0_outputs(11086));
    outputs(7142) <= (layer0_outputs(2163)) and not (layer0_outputs(12389));
    outputs(7143) <= not(layer0_outputs(7007)) or (layer0_outputs(4556));
    outputs(7144) <= not((layer0_outputs(10495)) and (layer0_outputs(4558)));
    outputs(7145) <= (layer0_outputs(11789)) and not (layer0_outputs(547));
    outputs(7146) <= not((layer0_outputs(911)) xor (layer0_outputs(414)));
    outputs(7147) <= not(layer0_outputs(11957));
    outputs(7148) <= not((layer0_outputs(2385)) xor (layer0_outputs(12658)));
    outputs(7149) <= not(layer0_outputs(3005)) or (layer0_outputs(9419));
    outputs(7150) <= (layer0_outputs(5027)) xor (layer0_outputs(2065));
    outputs(7151) <= layer0_outputs(7586);
    outputs(7152) <= (layer0_outputs(8801)) xor (layer0_outputs(8861));
    outputs(7153) <= (layer0_outputs(1531)) and not (layer0_outputs(12538));
    outputs(7154) <= not(layer0_outputs(3265));
    outputs(7155) <= not(layer0_outputs(6307));
    outputs(7156) <= not((layer0_outputs(10086)) and (layer0_outputs(3930)));
    outputs(7157) <= not(layer0_outputs(6910)) or (layer0_outputs(5430));
    outputs(7158) <= layer0_outputs(12512);
    outputs(7159) <= layer0_outputs(2569);
    outputs(7160) <= not(layer0_outputs(8070));
    outputs(7161) <= (layer0_outputs(7724)) xor (layer0_outputs(6778));
    outputs(7162) <= not(layer0_outputs(10074));
    outputs(7163) <= not((layer0_outputs(710)) and (layer0_outputs(1948)));
    outputs(7164) <= layer0_outputs(1619);
    outputs(7165) <= (layer0_outputs(10184)) xor (layer0_outputs(12605));
    outputs(7166) <= layer0_outputs(12236);
    outputs(7167) <= (layer0_outputs(7128)) xor (layer0_outputs(12576));
    outputs(7168) <= layer0_outputs(8211);
    outputs(7169) <= layer0_outputs(5997);
    outputs(7170) <= not(layer0_outputs(11826));
    outputs(7171) <= not((layer0_outputs(5117)) xor (layer0_outputs(6316)));
    outputs(7172) <= not((layer0_outputs(6738)) xor (layer0_outputs(2401)));
    outputs(7173) <= not(layer0_outputs(7619));
    outputs(7174) <= not(layer0_outputs(40));
    outputs(7175) <= (layer0_outputs(275)) xor (layer0_outputs(128));
    outputs(7176) <= (layer0_outputs(3441)) xor (layer0_outputs(10244));
    outputs(7177) <= (layer0_outputs(7000)) xor (layer0_outputs(3056));
    outputs(7178) <= (layer0_outputs(4058)) or (layer0_outputs(8252));
    outputs(7179) <= not(layer0_outputs(6489));
    outputs(7180) <= not((layer0_outputs(7140)) xor (layer0_outputs(11850)));
    outputs(7181) <= (layer0_outputs(10699)) and (layer0_outputs(2876));
    outputs(7182) <= not(layer0_outputs(6557));
    outputs(7183) <= not(layer0_outputs(9609));
    outputs(7184) <= (layer0_outputs(2385)) and (layer0_outputs(9134));
    outputs(7185) <= not(layer0_outputs(7600)) or (layer0_outputs(11288));
    outputs(7186) <= not(layer0_outputs(12121)) or (layer0_outputs(4382));
    outputs(7187) <= not(layer0_outputs(6321)) or (layer0_outputs(5061));
    outputs(7188) <= layer0_outputs(737);
    outputs(7189) <= layer0_outputs(4704);
    outputs(7190) <= (layer0_outputs(1525)) xor (layer0_outputs(4274));
    outputs(7191) <= (layer0_outputs(5822)) xor (layer0_outputs(7803));
    outputs(7192) <= (layer0_outputs(8943)) xor (layer0_outputs(470));
    outputs(7193) <= not((layer0_outputs(11761)) xor (layer0_outputs(2212)));
    outputs(7194) <= not((layer0_outputs(6041)) xor (layer0_outputs(4688)));
    outputs(7195) <= (layer0_outputs(2761)) xor (layer0_outputs(6314));
    outputs(7196) <= layer0_outputs(3904);
    outputs(7197) <= (layer0_outputs(1165)) xor (layer0_outputs(6017));
    outputs(7198) <= layer0_outputs(6873);
    outputs(7199) <= layer0_outputs(4319);
    outputs(7200) <= '1';
    outputs(7201) <= layer0_outputs(7109);
    outputs(7202) <= layer0_outputs(3944);
    outputs(7203) <= not(layer0_outputs(6014));
    outputs(7204) <= (layer0_outputs(12784)) xor (layer0_outputs(7499));
    outputs(7205) <= not((layer0_outputs(10480)) xor (layer0_outputs(7613)));
    outputs(7206) <= layer0_outputs(11968);
    outputs(7207) <= not(layer0_outputs(148));
    outputs(7208) <= not((layer0_outputs(844)) xor (layer0_outputs(5207)));
    outputs(7209) <= not(layer0_outputs(1495)) or (layer0_outputs(7005));
    outputs(7210) <= not((layer0_outputs(11550)) or (layer0_outputs(5836)));
    outputs(7211) <= not(layer0_outputs(12468));
    outputs(7212) <= not((layer0_outputs(6153)) xor (layer0_outputs(8508)));
    outputs(7213) <= layer0_outputs(838);
    outputs(7214) <= not(layer0_outputs(8215)) or (layer0_outputs(6362));
    outputs(7215) <= not(layer0_outputs(3615)) or (layer0_outputs(8363));
    outputs(7216) <= layer0_outputs(5050);
    outputs(7217) <= (layer0_outputs(8295)) and not (layer0_outputs(6098));
    outputs(7218) <= not(layer0_outputs(7796));
    outputs(7219) <= not((layer0_outputs(7840)) or (layer0_outputs(6723)));
    outputs(7220) <= not((layer0_outputs(10426)) or (layer0_outputs(4696)));
    outputs(7221) <= not((layer0_outputs(11795)) xor (layer0_outputs(5195)));
    outputs(7222) <= not(layer0_outputs(4362));
    outputs(7223) <= (layer0_outputs(6739)) or (layer0_outputs(8737));
    outputs(7224) <= layer0_outputs(9983);
    outputs(7225) <= not((layer0_outputs(10849)) xor (layer0_outputs(8678)));
    outputs(7226) <= not((layer0_outputs(10421)) and (layer0_outputs(11386)));
    outputs(7227) <= not((layer0_outputs(4144)) and (layer0_outputs(4386)));
    outputs(7228) <= (layer0_outputs(3626)) and not (layer0_outputs(9943));
    outputs(7229) <= (layer0_outputs(1961)) xor (layer0_outputs(6652));
    outputs(7230) <= (layer0_outputs(10981)) and not (layer0_outputs(1330));
    outputs(7231) <= not((layer0_outputs(7619)) xor (layer0_outputs(261)));
    outputs(7232) <= (layer0_outputs(12428)) and (layer0_outputs(5650));
    outputs(7233) <= (layer0_outputs(7370)) xor (layer0_outputs(7221));
    outputs(7234) <= (layer0_outputs(4491)) and not (layer0_outputs(11258));
    outputs(7235) <= layer0_outputs(11760);
    outputs(7236) <= (layer0_outputs(7851)) xor (layer0_outputs(4488));
    outputs(7237) <= (layer0_outputs(6041)) and (layer0_outputs(7867));
    outputs(7238) <= not(layer0_outputs(1654)) or (layer0_outputs(5785));
    outputs(7239) <= not(layer0_outputs(11104));
    outputs(7240) <= not(layer0_outputs(4367));
    outputs(7241) <= not(layer0_outputs(3063));
    outputs(7242) <= not(layer0_outputs(2401));
    outputs(7243) <= layer0_outputs(6047);
    outputs(7244) <= (layer0_outputs(11198)) xor (layer0_outputs(335));
    outputs(7245) <= not((layer0_outputs(2806)) xor (layer0_outputs(2129)));
    outputs(7246) <= layer0_outputs(8287);
    outputs(7247) <= layer0_outputs(8842);
    outputs(7248) <= not((layer0_outputs(3150)) xor (layer0_outputs(12590)));
    outputs(7249) <= layer0_outputs(9601);
    outputs(7250) <= not((layer0_outputs(7970)) and (layer0_outputs(167)));
    outputs(7251) <= layer0_outputs(9747);
    outputs(7252) <= (layer0_outputs(9061)) xor (layer0_outputs(9414));
    outputs(7253) <= (layer0_outputs(1168)) xor (layer0_outputs(5281));
    outputs(7254) <= layer0_outputs(12647);
    outputs(7255) <= not(layer0_outputs(5389));
    outputs(7256) <= not(layer0_outputs(3000));
    outputs(7257) <= not(layer0_outputs(2501));
    outputs(7258) <= (layer0_outputs(2984)) and (layer0_outputs(2831));
    outputs(7259) <= (layer0_outputs(12267)) xor (layer0_outputs(6700));
    outputs(7260) <= not((layer0_outputs(9272)) and (layer0_outputs(6359)));
    outputs(7261) <= (layer0_outputs(4294)) xor (layer0_outputs(11109));
    outputs(7262) <= (layer0_outputs(6799)) xor (layer0_outputs(5105));
    outputs(7263) <= not(layer0_outputs(10437)) or (layer0_outputs(4302));
    outputs(7264) <= layer0_outputs(1161);
    outputs(7265) <= (layer0_outputs(10040)) and (layer0_outputs(1629));
    outputs(7266) <= not(layer0_outputs(481)) or (layer0_outputs(6997));
    outputs(7267) <= (layer0_outputs(2793)) xor (layer0_outputs(8707));
    outputs(7268) <= (layer0_outputs(7778)) or (layer0_outputs(9845));
    outputs(7269) <= layer0_outputs(5202);
    outputs(7270) <= (layer0_outputs(5001)) xor (layer0_outputs(4682));
    outputs(7271) <= not((layer0_outputs(8960)) xor (layer0_outputs(3202)));
    outputs(7272) <= layer0_outputs(12509);
    outputs(7273) <= not((layer0_outputs(4693)) xor (layer0_outputs(252)));
    outputs(7274) <= (layer0_outputs(8931)) and not (layer0_outputs(5939));
    outputs(7275) <= layer0_outputs(9041);
    outputs(7276) <= (layer0_outputs(3039)) xor (layer0_outputs(7130));
    outputs(7277) <= (layer0_outputs(1038)) and not (layer0_outputs(22));
    outputs(7278) <= layer0_outputs(11307);
    outputs(7279) <= layer0_outputs(7708);
    outputs(7280) <= not((layer0_outputs(6696)) and (layer0_outputs(11380)));
    outputs(7281) <= not((layer0_outputs(1886)) or (layer0_outputs(8102)));
    outputs(7282) <= not(layer0_outputs(4682));
    outputs(7283) <= not((layer0_outputs(3865)) xor (layer0_outputs(8022)));
    outputs(7284) <= (layer0_outputs(9980)) and not (layer0_outputs(10811));
    outputs(7285) <= (layer0_outputs(8155)) and not (layer0_outputs(1407));
    outputs(7286) <= not((layer0_outputs(9762)) xor (layer0_outputs(5443)));
    outputs(7287) <= not(layer0_outputs(8231));
    outputs(7288) <= (layer0_outputs(6340)) and not (layer0_outputs(12190));
    outputs(7289) <= not((layer0_outputs(60)) xor (layer0_outputs(968)));
    outputs(7290) <= (layer0_outputs(10857)) xor (layer0_outputs(8076));
    outputs(7291) <= not(layer0_outputs(2935)) or (layer0_outputs(1751));
    outputs(7292) <= layer0_outputs(4373);
    outputs(7293) <= not((layer0_outputs(5151)) or (layer0_outputs(12189)));
    outputs(7294) <= '1';
    outputs(7295) <= layer0_outputs(874);
    outputs(7296) <= not((layer0_outputs(3463)) xor (layer0_outputs(470)));
    outputs(7297) <= not((layer0_outputs(10328)) xor (layer0_outputs(1514)));
    outputs(7298) <= layer0_outputs(4784);
    outputs(7299) <= not((layer0_outputs(9674)) xor (layer0_outputs(10445)));
    outputs(7300) <= not((layer0_outputs(821)) xor (layer0_outputs(9336)));
    outputs(7301) <= not(layer0_outputs(8502)) or (layer0_outputs(5029));
    outputs(7302) <= not(layer0_outputs(7278)) or (layer0_outputs(5952));
    outputs(7303) <= not((layer0_outputs(2791)) xor (layer0_outputs(10858)));
    outputs(7304) <= layer0_outputs(11002);
    outputs(7305) <= layer0_outputs(1225);
    outputs(7306) <= (layer0_outputs(1075)) and not (layer0_outputs(3894));
    outputs(7307) <= layer0_outputs(11858);
    outputs(7308) <= not(layer0_outputs(524));
    outputs(7309) <= layer0_outputs(10407);
    outputs(7310) <= not(layer0_outputs(1592));
    outputs(7311) <= (layer0_outputs(130)) xor (layer0_outputs(7662));
    outputs(7312) <= not(layer0_outputs(3026));
    outputs(7313) <= not((layer0_outputs(1430)) xor (layer0_outputs(3286)));
    outputs(7314) <= (layer0_outputs(1517)) xor (layer0_outputs(5281));
    outputs(7315) <= not((layer0_outputs(11309)) and (layer0_outputs(1535)));
    outputs(7316) <= layer0_outputs(4015);
    outputs(7317) <= not(layer0_outputs(11281));
    outputs(7318) <= (layer0_outputs(12338)) and (layer0_outputs(9477));
    outputs(7319) <= (layer0_outputs(8387)) xor (layer0_outputs(4192));
    outputs(7320) <= not((layer0_outputs(4565)) xor (layer0_outputs(12225)));
    outputs(7321) <= not(layer0_outputs(439));
    outputs(7322) <= not(layer0_outputs(2169)) or (layer0_outputs(6603));
    outputs(7323) <= layer0_outputs(6402);
    outputs(7324) <= not(layer0_outputs(6656));
    outputs(7325) <= (layer0_outputs(10987)) xor (layer0_outputs(1095));
    outputs(7326) <= layer0_outputs(5261);
    outputs(7327) <= not((layer0_outputs(8240)) xor (layer0_outputs(7503)));
    outputs(7328) <= (layer0_outputs(11762)) xor (layer0_outputs(2232));
    outputs(7329) <= (layer0_outputs(9376)) xor (layer0_outputs(10104));
    outputs(7330) <= layer0_outputs(4766);
    outputs(7331) <= not((layer0_outputs(12154)) xor (layer0_outputs(5756)));
    outputs(7332) <= (layer0_outputs(1047)) xor (layer0_outputs(1755));
    outputs(7333) <= (layer0_outputs(6409)) and not (layer0_outputs(3270));
    outputs(7334) <= not(layer0_outputs(10182));
    outputs(7335) <= not((layer0_outputs(1334)) xor (layer0_outputs(12319)));
    outputs(7336) <= not((layer0_outputs(7210)) xor (layer0_outputs(3828)));
    outputs(7337) <= not((layer0_outputs(2609)) xor (layer0_outputs(7723)));
    outputs(7338) <= not(layer0_outputs(6614));
    outputs(7339) <= (layer0_outputs(1034)) or (layer0_outputs(8079));
    outputs(7340) <= (layer0_outputs(4363)) or (layer0_outputs(109));
    outputs(7341) <= (layer0_outputs(4798)) xor (layer0_outputs(10220));
    outputs(7342) <= (layer0_outputs(10078)) and not (layer0_outputs(3306));
    outputs(7343) <= not((layer0_outputs(8541)) xor (layer0_outputs(11745)));
    outputs(7344) <= layer0_outputs(12624);
    outputs(7345) <= (layer0_outputs(4530)) xor (layer0_outputs(2829));
    outputs(7346) <= (layer0_outputs(8895)) or (layer0_outputs(245));
    outputs(7347) <= '1';
    outputs(7348) <= layer0_outputs(8436);
    outputs(7349) <= (layer0_outputs(11929)) and not (layer0_outputs(6067));
    outputs(7350) <= layer0_outputs(9880);
    outputs(7351) <= (layer0_outputs(1668)) and not (layer0_outputs(2507));
    outputs(7352) <= not(layer0_outputs(2242));
    outputs(7353) <= not((layer0_outputs(5319)) xor (layer0_outputs(7181)));
    outputs(7354) <= layer0_outputs(4272);
    outputs(7355) <= not(layer0_outputs(6376));
    outputs(7356) <= (layer0_outputs(536)) xor (layer0_outputs(12371));
    outputs(7357) <= layer0_outputs(3975);
    outputs(7358) <= (layer0_outputs(6790)) xor (layer0_outputs(8675));
    outputs(7359) <= not((layer0_outputs(4160)) xor (layer0_outputs(9493)));
    outputs(7360) <= (layer0_outputs(6263)) or (layer0_outputs(1341));
    outputs(7361) <= layer0_outputs(5909);
    outputs(7362) <= (layer0_outputs(5256)) xor (layer0_outputs(3914));
    outputs(7363) <= not(layer0_outputs(8420));
    outputs(7364) <= not((layer0_outputs(10983)) xor (layer0_outputs(1041)));
    outputs(7365) <= layer0_outputs(6161);
    outputs(7366) <= (layer0_outputs(10783)) xor (layer0_outputs(11127));
    outputs(7367) <= not((layer0_outputs(4391)) and (layer0_outputs(11846)));
    outputs(7368) <= not(layer0_outputs(7034));
    outputs(7369) <= (layer0_outputs(9039)) xor (layer0_outputs(12023));
    outputs(7370) <= not(layer0_outputs(9752)) or (layer0_outputs(12075));
    outputs(7371) <= not(layer0_outputs(3876)) or (layer0_outputs(7104));
    outputs(7372) <= not((layer0_outputs(3240)) xor (layer0_outputs(4133)));
    outputs(7373) <= not(layer0_outputs(11692)) or (layer0_outputs(209));
    outputs(7374) <= layer0_outputs(11325);
    outputs(7375) <= layer0_outputs(696);
    outputs(7376) <= (layer0_outputs(10678)) and not (layer0_outputs(2072));
    outputs(7377) <= (layer0_outputs(10923)) xor (layer0_outputs(604));
    outputs(7378) <= (layer0_outputs(4059)) and (layer0_outputs(5196));
    outputs(7379) <= layer0_outputs(1162);
    outputs(7380) <= (layer0_outputs(5309)) xor (layer0_outputs(8679));
    outputs(7381) <= not((layer0_outputs(6488)) xor (layer0_outputs(9379)));
    outputs(7382) <= (layer0_outputs(8154)) and not (layer0_outputs(3297));
    outputs(7383) <= not(layer0_outputs(6951));
    outputs(7384) <= (layer0_outputs(11903)) and not (layer0_outputs(12017));
    outputs(7385) <= layer0_outputs(8832);
    outputs(7386) <= layer0_outputs(1032);
    outputs(7387) <= not((layer0_outputs(9159)) xor (layer0_outputs(9373)));
    outputs(7388) <= not(layer0_outputs(12203)) or (layer0_outputs(10278));
    outputs(7389) <= (layer0_outputs(2124)) xor (layer0_outputs(2878));
    outputs(7390) <= (layer0_outputs(3067)) xor (layer0_outputs(3236));
    outputs(7391) <= layer0_outputs(4145);
    outputs(7392) <= not(layer0_outputs(6134));
    outputs(7393) <= not((layer0_outputs(1271)) xor (layer0_outputs(8884)));
    outputs(7394) <= (layer0_outputs(10176)) xor (layer0_outputs(11861));
    outputs(7395) <= not(layer0_outputs(7223));
    outputs(7396) <= (layer0_outputs(2263)) xor (layer0_outputs(5932));
    outputs(7397) <= not(layer0_outputs(4427));
    outputs(7398) <= not((layer0_outputs(9416)) xor (layer0_outputs(3189)));
    outputs(7399) <= not(layer0_outputs(25)) or (layer0_outputs(5437));
    outputs(7400) <= layer0_outputs(5262);
    outputs(7401) <= (layer0_outputs(4080)) and not (layer0_outputs(751));
    outputs(7402) <= (layer0_outputs(8154)) and (layer0_outputs(3605));
    outputs(7403) <= (layer0_outputs(10004)) and not (layer0_outputs(11657));
    outputs(7404) <= not((layer0_outputs(6459)) or (layer0_outputs(6823)));
    outputs(7405) <= layer0_outputs(10317);
    outputs(7406) <= not((layer0_outputs(11874)) xor (layer0_outputs(4372)));
    outputs(7407) <= not(layer0_outputs(4149)) or (layer0_outputs(3470));
    outputs(7408) <= layer0_outputs(1817);
    outputs(7409) <= not((layer0_outputs(4092)) and (layer0_outputs(6621)));
    outputs(7410) <= not(layer0_outputs(9300)) or (layer0_outputs(3467));
    outputs(7411) <= layer0_outputs(10213);
    outputs(7412) <= (layer0_outputs(7117)) xor (layer0_outputs(9246));
    outputs(7413) <= layer0_outputs(6687);
    outputs(7414) <= layer0_outputs(1060);
    outputs(7415) <= not((layer0_outputs(10410)) or (layer0_outputs(7980)));
    outputs(7416) <= not(layer0_outputs(7939)) or (layer0_outputs(910));
    outputs(7417) <= not((layer0_outputs(8064)) xor (layer0_outputs(1839)));
    outputs(7418) <= not((layer0_outputs(7750)) xor (layer0_outputs(5802)));
    outputs(7419) <= not(layer0_outputs(11458)) or (layer0_outputs(6292));
    outputs(7420) <= not(layer0_outputs(3034)) or (layer0_outputs(6821));
    outputs(7421) <= layer0_outputs(9202);
    outputs(7422) <= '1';
    outputs(7423) <= not(layer0_outputs(11466)) or (layer0_outputs(4566));
    outputs(7424) <= (layer0_outputs(3711)) and not (layer0_outputs(3265));
    outputs(7425) <= layer0_outputs(1391);
    outputs(7426) <= (layer0_outputs(11493)) xor (layer0_outputs(2612));
    outputs(7427) <= (layer0_outputs(6101)) xor (layer0_outputs(5763));
    outputs(7428) <= not(layer0_outputs(4670)) or (layer0_outputs(8917));
    outputs(7429) <= not((layer0_outputs(2377)) xor (layer0_outputs(345)));
    outputs(7430) <= not(layer0_outputs(2049));
    outputs(7431) <= (layer0_outputs(9527)) or (layer0_outputs(8391));
    outputs(7432) <= not(layer0_outputs(6261));
    outputs(7433) <= not(layer0_outputs(3095));
    outputs(7434) <= not(layer0_outputs(12794)) or (layer0_outputs(6947));
    outputs(7435) <= (layer0_outputs(9794)) and not (layer0_outputs(6373));
    outputs(7436) <= not(layer0_outputs(2750)) or (layer0_outputs(4515));
    outputs(7437) <= layer0_outputs(12407);
    outputs(7438) <= not((layer0_outputs(9042)) xor (layer0_outputs(1909)));
    outputs(7439) <= (layer0_outputs(8743)) or (layer0_outputs(8299));
    outputs(7440) <= not(layer0_outputs(3016)) or (layer0_outputs(6890));
    outputs(7441) <= not(layer0_outputs(1380)) or (layer0_outputs(112));
    outputs(7442) <= (layer0_outputs(12643)) and not (layer0_outputs(2662));
    outputs(7443) <= (layer0_outputs(8280)) xor (layer0_outputs(547));
    outputs(7444) <= not(layer0_outputs(10052)) or (layer0_outputs(12035));
    outputs(7445) <= not(layer0_outputs(355)) or (layer0_outputs(8944));
    outputs(7446) <= layer0_outputs(4323);
    outputs(7447) <= '1';
    outputs(7448) <= layer0_outputs(1884);
    outputs(7449) <= (layer0_outputs(7436)) or (layer0_outputs(7003));
    outputs(7450) <= not((layer0_outputs(7015)) xor (layer0_outputs(323)));
    outputs(7451) <= layer0_outputs(8079);
    outputs(7452) <= not(layer0_outputs(4913));
    outputs(7453) <= (layer0_outputs(3173)) xor (layer0_outputs(2648));
    outputs(7454) <= (layer0_outputs(6222)) xor (layer0_outputs(8737));
    outputs(7455) <= layer0_outputs(7783);
    outputs(7456) <= (layer0_outputs(11612)) xor (layer0_outputs(3595));
    outputs(7457) <= not(layer0_outputs(7585)) or (layer0_outputs(5534));
    outputs(7458) <= (layer0_outputs(4890)) xor (layer0_outputs(4452));
    outputs(7459) <= not((layer0_outputs(9110)) xor (layer0_outputs(9278)));
    outputs(7460) <= not((layer0_outputs(6447)) xor (layer0_outputs(7756)));
    outputs(7461) <= (layer0_outputs(2345)) or (layer0_outputs(1303));
    outputs(7462) <= layer0_outputs(1883);
    outputs(7463) <= layer0_outputs(678);
    outputs(7464) <= (layer0_outputs(10679)) xor (layer0_outputs(3694));
    outputs(7465) <= (layer0_outputs(12503)) and not (layer0_outputs(8870));
    outputs(7466) <= (layer0_outputs(2707)) xor (layer0_outputs(2136));
    outputs(7467) <= not(layer0_outputs(11387));
    outputs(7468) <= not(layer0_outputs(9730));
    outputs(7469) <= not(layer0_outputs(4251));
    outputs(7470) <= not(layer0_outputs(6304));
    outputs(7471) <= not(layer0_outputs(5638));
    outputs(7472) <= not(layer0_outputs(1879)) or (layer0_outputs(4916));
    outputs(7473) <= layer0_outputs(5550);
    outputs(7474) <= layer0_outputs(222);
    outputs(7475) <= (layer0_outputs(9193)) and not (layer0_outputs(5232));
    outputs(7476) <= layer0_outputs(205);
    outputs(7477) <= not(layer0_outputs(10997));
    outputs(7478) <= layer0_outputs(8695);
    outputs(7479) <= not((layer0_outputs(59)) and (layer0_outputs(5602)));
    outputs(7480) <= not((layer0_outputs(9451)) and (layer0_outputs(1892)));
    outputs(7481) <= (layer0_outputs(11243)) xor (layer0_outputs(12769));
    outputs(7482) <= not(layer0_outputs(3916));
    outputs(7483) <= not(layer0_outputs(8470));
    outputs(7484) <= (layer0_outputs(2086)) xor (layer0_outputs(11630));
    outputs(7485) <= layer0_outputs(7738);
    outputs(7486) <= layer0_outputs(10210);
    outputs(7487) <= not(layer0_outputs(10285));
    outputs(7488) <= not((layer0_outputs(9653)) xor (layer0_outputs(4627)));
    outputs(7489) <= not((layer0_outputs(130)) xor (layer0_outputs(1552)));
    outputs(7490) <= not((layer0_outputs(4324)) xor (layer0_outputs(6322)));
    outputs(7491) <= not(layer0_outputs(3410));
    outputs(7492) <= layer0_outputs(8788);
    outputs(7493) <= layer0_outputs(2036);
    outputs(7494) <= not(layer0_outputs(3853));
    outputs(7495) <= not((layer0_outputs(1409)) xor (layer0_outputs(9363)));
    outputs(7496) <= not(layer0_outputs(3608)) or (layer0_outputs(5637));
    outputs(7497) <= layer0_outputs(1597);
    outputs(7498) <= not((layer0_outputs(4324)) xor (layer0_outputs(8907)));
    outputs(7499) <= (layer0_outputs(5645)) and not (layer0_outputs(10837));
    outputs(7500) <= not(layer0_outputs(5912));
    outputs(7501) <= not((layer0_outputs(6835)) and (layer0_outputs(3705)));
    outputs(7502) <= not(layer0_outputs(1768)) or (layer0_outputs(6110));
    outputs(7503) <= layer0_outputs(11172);
    outputs(7504) <= not((layer0_outputs(2134)) xor (layer0_outputs(9404)));
    outputs(7505) <= (layer0_outputs(7566)) xor (layer0_outputs(5882));
    outputs(7506) <= not((layer0_outputs(5664)) xor (layer0_outputs(4633)));
    outputs(7507) <= not(layer0_outputs(3380));
    outputs(7508) <= layer0_outputs(9998);
    outputs(7509) <= not(layer0_outputs(1539));
    outputs(7510) <= (layer0_outputs(4555)) and not (layer0_outputs(3436));
    outputs(7511) <= not(layer0_outputs(2757)) or (layer0_outputs(1549));
    outputs(7512) <= layer0_outputs(6807);
    outputs(7513) <= (layer0_outputs(8222)) xor (layer0_outputs(5735));
    outputs(7514) <= layer0_outputs(5749);
    outputs(7515) <= layer0_outputs(10011);
    outputs(7516) <= (layer0_outputs(5346)) and not (layer0_outputs(2562));
    outputs(7517) <= (layer0_outputs(11088)) or (layer0_outputs(480));
    outputs(7518) <= not(layer0_outputs(4097)) or (layer0_outputs(2069));
    outputs(7519) <= (layer0_outputs(11199)) or (layer0_outputs(9507));
    outputs(7520) <= not(layer0_outputs(12575)) or (layer0_outputs(2287));
    outputs(7521) <= not(layer0_outputs(9877));
    outputs(7522) <= (layer0_outputs(12406)) and (layer0_outputs(5150));
    outputs(7523) <= not((layer0_outputs(6197)) and (layer0_outputs(8825)));
    outputs(7524) <= layer0_outputs(12591);
    outputs(7525) <= layer0_outputs(9701);
    outputs(7526) <= not((layer0_outputs(11320)) xor (layer0_outputs(1665)));
    outputs(7527) <= (layer0_outputs(1222)) xor (layer0_outputs(1453));
    outputs(7528) <= (layer0_outputs(1120)) xor (layer0_outputs(10398));
    outputs(7529) <= not(layer0_outputs(633)) or (layer0_outputs(10388));
    outputs(7530) <= not((layer0_outputs(3640)) and (layer0_outputs(1233)));
    outputs(7531) <= not(layer0_outputs(6167));
    outputs(7532) <= not((layer0_outputs(8779)) xor (layer0_outputs(7814)));
    outputs(7533) <= not(layer0_outputs(8931));
    outputs(7534) <= not((layer0_outputs(6930)) xor (layer0_outputs(6214)));
    outputs(7535) <= (layer0_outputs(5847)) and not (layer0_outputs(8901));
    outputs(7536) <= layer0_outputs(10915);
    outputs(7537) <= not(layer0_outputs(303));
    outputs(7538) <= '1';
    outputs(7539) <= not(layer0_outputs(9911)) or (layer0_outputs(11670));
    outputs(7540) <= (layer0_outputs(12317)) and not (layer0_outputs(10613));
    outputs(7541) <= not(layer0_outputs(2713)) or (layer0_outputs(2641));
    outputs(7542) <= (layer0_outputs(12178)) xor (layer0_outputs(3857));
    outputs(7543) <= not((layer0_outputs(873)) and (layer0_outputs(6025)));
    outputs(7544) <= not(layer0_outputs(3423));
    outputs(7545) <= layer0_outputs(12072);
    outputs(7546) <= (layer0_outputs(8937)) and (layer0_outputs(281));
    outputs(7547) <= layer0_outputs(6386);
    outputs(7548) <= not((layer0_outputs(425)) xor (layer0_outputs(12487)));
    outputs(7549) <= not((layer0_outputs(3459)) and (layer0_outputs(7774)));
    outputs(7550) <= not((layer0_outputs(6935)) xor (layer0_outputs(12430)));
    outputs(7551) <= not(layer0_outputs(12397));
    outputs(7552) <= (layer0_outputs(831)) or (layer0_outputs(3158));
    outputs(7553) <= layer0_outputs(6317);
    outputs(7554) <= not(layer0_outputs(5368));
    outputs(7555) <= not(layer0_outputs(10344));
    outputs(7556) <= not((layer0_outputs(11909)) xor (layer0_outputs(3529)));
    outputs(7557) <= not(layer0_outputs(6481)) or (layer0_outputs(8627));
    outputs(7558) <= not((layer0_outputs(4893)) xor (layer0_outputs(575)));
    outputs(7559) <= not((layer0_outputs(11907)) xor (layer0_outputs(7480)));
    outputs(7560) <= layer0_outputs(11453);
    outputs(7561) <= (layer0_outputs(4553)) xor (layer0_outputs(9542));
    outputs(7562) <= layer0_outputs(3901);
    outputs(7563) <= not(layer0_outputs(8009)) or (layer0_outputs(10731));
    outputs(7564) <= layer0_outputs(7695);
    outputs(7565) <= layer0_outputs(1151);
    outputs(7566) <= layer0_outputs(11639);
    outputs(7567) <= not((layer0_outputs(995)) or (layer0_outputs(4816)));
    outputs(7568) <= (layer0_outputs(1547)) xor (layer0_outputs(7688));
    outputs(7569) <= not(layer0_outputs(5603));
    outputs(7570) <= not((layer0_outputs(9351)) xor (layer0_outputs(2660)));
    outputs(7571) <= not(layer0_outputs(9738));
    outputs(7572) <= (layer0_outputs(3131)) xor (layer0_outputs(1446));
    outputs(7573) <= (layer0_outputs(12724)) or (layer0_outputs(3166));
    outputs(7574) <= not(layer0_outputs(9122));
    outputs(7575) <= not((layer0_outputs(6087)) xor (layer0_outputs(879)));
    outputs(7576) <= not(layer0_outputs(1422)) or (layer0_outputs(10363));
    outputs(7577) <= (layer0_outputs(2052)) or (layer0_outputs(2240));
    outputs(7578) <= (layer0_outputs(8393)) xor (layer0_outputs(1099));
    outputs(7579) <= layer0_outputs(6322);
    outputs(7580) <= (layer0_outputs(11349)) and not (layer0_outputs(8125));
    outputs(7581) <= layer0_outputs(10226);
    outputs(7582) <= (layer0_outputs(6151)) xor (layer0_outputs(5691));
    outputs(7583) <= not(layer0_outputs(9958));
    outputs(7584) <= (layer0_outputs(1808)) or (layer0_outputs(11612));
    outputs(7585) <= '1';
    outputs(7586) <= layer0_outputs(3015);
    outputs(7587) <= (layer0_outputs(9103)) and not (layer0_outputs(11756));
    outputs(7588) <= not(layer0_outputs(12771)) or (layer0_outputs(5694));
    outputs(7589) <= not(layer0_outputs(5557));
    outputs(7590) <= layer0_outputs(5967);
    outputs(7591) <= not(layer0_outputs(1274));
    outputs(7592) <= (layer0_outputs(5021)) xor (layer0_outputs(179));
    outputs(7593) <= not((layer0_outputs(1013)) xor (layer0_outputs(6451)));
    outputs(7594) <= layer0_outputs(9181);
    outputs(7595) <= layer0_outputs(4722);
    outputs(7596) <= layer0_outputs(3609);
    outputs(7597) <= not(layer0_outputs(2083)) or (layer0_outputs(9873));
    outputs(7598) <= (layer0_outputs(5376)) xor (layer0_outputs(6553));
    outputs(7599) <= layer0_outputs(7258);
    outputs(7600) <= layer0_outputs(8398);
    outputs(7601) <= (layer0_outputs(8757)) and not (layer0_outputs(12028));
    outputs(7602) <= not(layer0_outputs(9500));
    outputs(7603) <= not((layer0_outputs(792)) xor (layer0_outputs(3160)));
    outputs(7604) <= not((layer0_outputs(10748)) xor (layer0_outputs(554)));
    outputs(7605) <= (layer0_outputs(8451)) or (layer0_outputs(3020));
    outputs(7606) <= (layer0_outputs(3629)) xor (layer0_outputs(351));
    outputs(7607) <= not((layer0_outputs(7963)) or (layer0_outputs(7119)));
    outputs(7608) <= (layer0_outputs(192)) xor (layer0_outputs(7614));
    outputs(7609) <= not(layer0_outputs(3261)) or (layer0_outputs(4277));
    outputs(7610) <= (layer0_outputs(4506)) and not (layer0_outputs(11978));
    outputs(7611) <= not(layer0_outputs(187));
    outputs(7612) <= not((layer0_outputs(8643)) and (layer0_outputs(11327)));
    outputs(7613) <= (layer0_outputs(6423)) and not (layer0_outputs(8835));
    outputs(7614) <= not((layer0_outputs(10868)) xor (layer0_outputs(9980)));
    outputs(7615) <= not((layer0_outputs(9250)) xor (layer0_outputs(12081)));
    outputs(7616) <= (layer0_outputs(527)) xor (layer0_outputs(6227));
    outputs(7617) <= not((layer0_outputs(1625)) and (layer0_outputs(11450)));
    outputs(7618) <= not(layer0_outputs(4151)) or (layer0_outputs(5852));
    outputs(7619) <= (layer0_outputs(3508)) or (layer0_outputs(11531));
    outputs(7620) <= not((layer0_outputs(5806)) xor (layer0_outputs(3987)));
    outputs(7621) <= not(layer0_outputs(9372));
    outputs(7622) <= layer0_outputs(5511);
    outputs(7623) <= not((layer0_outputs(5919)) and (layer0_outputs(1930)));
    outputs(7624) <= (layer0_outputs(4155)) and (layer0_outputs(2892));
    outputs(7625) <= (layer0_outputs(1464)) and not (layer0_outputs(9696));
    outputs(7626) <= layer0_outputs(6746);
    outputs(7627) <= not(layer0_outputs(5662));
    outputs(7628) <= layer0_outputs(8520);
    outputs(7629) <= not((layer0_outputs(12058)) xor (layer0_outputs(10331)));
    outputs(7630) <= not((layer0_outputs(5837)) and (layer0_outputs(2704)));
    outputs(7631) <= (layer0_outputs(12305)) xor (layer0_outputs(8143));
    outputs(7632) <= not((layer0_outputs(6715)) and (layer0_outputs(6148)));
    outputs(7633) <= (layer0_outputs(11222)) xor (layer0_outputs(1345));
    outputs(7634) <= not((layer0_outputs(7333)) or (layer0_outputs(8947)));
    outputs(7635) <= not(layer0_outputs(8378));
    outputs(7636) <= not((layer0_outputs(7156)) xor (layer0_outputs(7998)));
    outputs(7637) <= not((layer0_outputs(8948)) xor (layer0_outputs(12354)));
    outputs(7638) <= (layer0_outputs(9530)) xor (layer0_outputs(1645));
    outputs(7639) <= not((layer0_outputs(114)) xor (layer0_outputs(9691)));
    outputs(7640) <= not(layer0_outputs(4713)) or (layer0_outputs(2852));
    outputs(7641) <= not((layer0_outputs(12246)) xor (layer0_outputs(9664)));
    outputs(7642) <= (layer0_outputs(12569)) or (layer0_outputs(12186));
    outputs(7643) <= layer0_outputs(2028);
    outputs(7644) <= (layer0_outputs(754)) xor (layer0_outputs(7099));
    outputs(7645) <= '1';
    outputs(7646) <= not(layer0_outputs(5938));
    outputs(7647) <= (layer0_outputs(12268)) xor (layer0_outputs(1493));
    outputs(7648) <= (layer0_outputs(10422)) and not (layer0_outputs(12515));
    outputs(7649) <= not((layer0_outputs(1652)) and (layer0_outputs(6872)));
    outputs(7650) <= not((layer0_outputs(7449)) xor (layer0_outputs(11697)));
    outputs(7651) <= layer0_outputs(7094);
    outputs(7652) <= (layer0_outputs(12662)) xor (layer0_outputs(6371));
    outputs(7653) <= not(layer0_outputs(1558));
    outputs(7654) <= (layer0_outputs(2325)) and (layer0_outputs(11192));
    outputs(7655) <= (layer0_outputs(5102)) xor (layer0_outputs(10930));
    outputs(7656) <= not((layer0_outputs(10027)) xor (layer0_outputs(3498)));
    outputs(7657) <= not(layer0_outputs(3034));
    outputs(7658) <= layer0_outputs(3633);
    outputs(7659) <= layer0_outputs(10287);
    outputs(7660) <= not((layer0_outputs(6482)) xor (layer0_outputs(1133)));
    outputs(7661) <= not((layer0_outputs(6525)) xor (layer0_outputs(12684)));
    outputs(7662) <= (layer0_outputs(8747)) or (layer0_outputs(3980));
    outputs(7663) <= layer0_outputs(11050);
    outputs(7664) <= not((layer0_outputs(300)) and (layer0_outputs(7198)));
    outputs(7665) <= (layer0_outputs(1870)) or (layer0_outputs(10901));
    outputs(7666) <= layer0_outputs(11490);
    outputs(7667) <= layer0_outputs(11363);
    outputs(7668) <= not((layer0_outputs(8599)) xor (layer0_outputs(11823)));
    outputs(7669) <= not(layer0_outputs(1548));
    outputs(7670) <= (layer0_outputs(3855)) and (layer0_outputs(5075));
    outputs(7671) <= not(layer0_outputs(9872)) or (layer0_outputs(5553));
    outputs(7672) <= not(layer0_outputs(819)) or (layer0_outputs(2258));
    outputs(7673) <= (layer0_outputs(8217)) xor (layer0_outputs(398));
    outputs(7674) <= not((layer0_outputs(10656)) xor (layer0_outputs(7897)));
    outputs(7675) <= (layer0_outputs(246)) and (layer0_outputs(12651));
    outputs(7676) <= not(layer0_outputs(5084)) or (layer0_outputs(1716));
    outputs(7677) <= layer0_outputs(1248);
    outputs(7678) <= not(layer0_outputs(6987));
    outputs(7679) <= (layer0_outputs(2102)) or (layer0_outputs(11821));
    outputs(7680) <= not(layer0_outputs(9003)) or (layer0_outputs(2369));
    outputs(7681) <= layer0_outputs(8169);
    outputs(7682) <= not((layer0_outputs(5700)) xor (layer0_outputs(366)));
    outputs(7683) <= layer0_outputs(8542);
    outputs(7684) <= layer0_outputs(9445);
    outputs(7685) <= not(layer0_outputs(7356));
    outputs(7686) <= not(layer0_outputs(11310));
    outputs(7687) <= not((layer0_outputs(4674)) xor (layer0_outputs(10723)));
    outputs(7688) <= not((layer0_outputs(6559)) and (layer0_outputs(8412)));
    outputs(7689) <= (layer0_outputs(4827)) or (layer0_outputs(2108));
    outputs(7690) <= layer0_outputs(12425);
    outputs(7691) <= layer0_outputs(12117);
    outputs(7692) <= not((layer0_outputs(7761)) xor (layer0_outputs(981)));
    outputs(7693) <= not(layer0_outputs(1842));
    outputs(7694) <= not(layer0_outputs(5517)) or (layer0_outputs(9828));
    outputs(7695) <= (layer0_outputs(10955)) xor (layer0_outputs(12693));
    outputs(7696) <= not((layer0_outputs(6669)) xor (layer0_outputs(2454)));
    outputs(7697) <= layer0_outputs(8218);
    outputs(7698) <= (layer0_outputs(2608)) and not (layer0_outputs(87));
    outputs(7699) <= not((layer0_outputs(11080)) or (layer0_outputs(2379)));
    outputs(7700) <= not(layer0_outputs(3698));
    outputs(7701) <= not(layer0_outputs(8058)) or (layer0_outputs(7893));
    outputs(7702) <= (layer0_outputs(7866)) and (layer0_outputs(10660));
    outputs(7703) <= not((layer0_outputs(11121)) xor (layer0_outputs(538)));
    outputs(7704) <= not((layer0_outputs(9644)) xor (layer0_outputs(6539)));
    outputs(7705) <= (layer0_outputs(3754)) and not (layer0_outputs(4320));
    outputs(7706) <= (layer0_outputs(7254)) or (layer0_outputs(12622));
    outputs(7707) <= not(layer0_outputs(1101));
    outputs(7708) <= layer0_outputs(11473);
    outputs(7709) <= layer0_outputs(4292);
    outputs(7710) <= not(layer0_outputs(4300));
    outputs(7711) <= not(layer0_outputs(5915));
    outputs(7712) <= not((layer0_outputs(5139)) or (layer0_outputs(2477)));
    outputs(7713) <= layer0_outputs(10739);
    outputs(7714) <= layer0_outputs(679);
    outputs(7715) <= (layer0_outputs(5461)) xor (layer0_outputs(4512));
    outputs(7716) <= (layer0_outputs(134)) and not (layer0_outputs(7378));
    outputs(7717) <= not((layer0_outputs(5839)) xor (layer0_outputs(4943)));
    outputs(7718) <= not((layer0_outputs(7067)) xor (layer0_outputs(6713)));
    outputs(7719) <= (layer0_outputs(11570)) xor (layer0_outputs(11078));
    outputs(7720) <= layer0_outputs(10559);
    outputs(7721) <= (layer0_outputs(9928)) and not (layer0_outputs(5280));
    outputs(7722) <= not(layer0_outputs(6932));
    outputs(7723) <= not(layer0_outputs(1601));
    outputs(7724) <= layer0_outputs(69);
    outputs(7725) <= not(layer0_outputs(4074)) or (layer0_outputs(11045));
    outputs(7726) <= not(layer0_outputs(3760));
    outputs(7727) <= layer0_outputs(10798);
    outputs(7728) <= not((layer0_outputs(3487)) and (layer0_outputs(9360)));
    outputs(7729) <= (layer0_outputs(11250)) xor (layer0_outputs(162));
    outputs(7730) <= layer0_outputs(9099);
    outputs(7731) <= layer0_outputs(4644);
    outputs(7732) <= '1';
    outputs(7733) <= not(layer0_outputs(2185));
    outputs(7734) <= '0';
    outputs(7735) <= layer0_outputs(6814);
    outputs(7736) <= not(layer0_outputs(11333));
    outputs(7737) <= layer0_outputs(8405);
    outputs(7738) <= (layer0_outputs(344)) or (layer0_outputs(12243));
    outputs(7739) <= (layer0_outputs(2303)) and not (layer0_outputs(4725));
    outputs(7740) <= (layer0_outputs(3882)) and not (layer0_outputs(11898));
    outputs(7741) <= not(layer0_outputs(4810)) or (layer0_outputs(8984));
    outputs(7742) <= not((layer0_outputs(890)) or (layer0_outputs(2812)));
    outputs(7743) <= not(layer0_outputs(2187)) or (layer0_outputs(8295));
    outputs(7744) <= layer0_outputs(1376);
    outputs(7745) <= layer0_outputs(1009);
    outputs(7746) <= not((layer0_outputs(6044)) and (layer0_outputs(232)));
    outputs(7747) <= layer0_outputs(3588);
    outputs(7748) <= layer0_outputs(5012);
    outputs(7749) <= not(layer0_outputs(1624));
    outputs(7750) <= not((layer0_outputs(3819)) xor (layer0_outputs(608)));
    outputs(7751) <= not((layer0_outputs(5160)) or (layer0_outputs(11556)));
    outputs(7752) <= (layer0_outputs(878)) and (layer0_outputs(3689));
    outputs(7753) <= not(layer0_outputs(5885));
    outputs(7754) <= not((layer0_outputs(2151)) xor (layer0_outputs(5189)));
    outputs(7755) <= not(layer0_outputs(2300)) or (layer0_outputs(12799));
    outputs(7756) <= (layer0_outputs(2373)) and not (layer0_outputs(4588));
    outputs(7757) <= layer0_outputs(4722);
    outputs(7758) <= not(layer0_outputs(1812));
    outputs(7759) <= layer0_outputs(338);
    outputs(7760) <= layer0_outputs(10387);
    outputs(7761) <= not(layer0_outputs(11951));
    outputs(7762) <= (layer0_outputs(2420)) xor (layer0_outputs(5951));
    outputs(7763) <= not((layer0_outputs(11958)) or (layer0_outputs(4897)));
    outputs(7764) <= not((layer0_outputs(4881)) xor (layer0_outputs(2130)));
    outputs(7765) <= (layer0_outputs(1885)) xor (layer0_outputs(6537));
    outputs(7766) <= (layer0_outputs(7535)) xor (layer0_outputs(12283));
    outputs(7767) <= not((layer0_outputs(9144)) xor (layer0_outputs(2763)));
    outputs(7768) <= (layer0_outputs(11445)) xor (layer0_outputs(10952));
    outputs(7769) <= (layer0_outputs(4031)) and (layer0_outputs(1686));
    outputs(7770) <= not(layer0_outputs(4976));
    outputs(7771) <= not((layer0_outputs(8279)) xor (layer0_outputs(10944)));
    outputs(7772) <= not((layer0_outputs(1413)) xor (layer0_outputs(11672)));
    outputs(7773) <= layer0_outputs(4955);
    outputs(7774) <= not(layer0_outputs(7763));
    outputs(7775) <= not((layer0_outputs(265)) and (layer0_outputs(10844)));
    outputs(7776) <= not((layer0_outputs(2414)) xor (layer0_outputs(7380)));
    outputs(7777) <= not(layer0_outputs(11875));
    outputs(7778) <= not((layer0_outputs(2400)) and (layer0_outputs(3360)));
    outputs(7779) <= layer0_outputs(8476);
    outputs(7780) <= (layer0_outputs(2182)) xor (layer0_outputs(10133));
    outputs(7781) <= layer0_outputs(2012);
    outputs(7782) <= layer0_outputs(11099);
    outputs(7783) <= not(layer0_outputs(3352));
    outputs(7784) <= not(layer0_outputs(7175));
    outputs(7785) <= layer0_outputs(6278);
    outputs(7786) <= (layer0_outputs(507)) and not (layer0_outputs(5122));
    outputs(7787) <= not(layer0_outputs(1940));
    outputs(7788) <= not((layer0_outputs(8282)) xor (layer0_outputs(3671)));
    outputs(7789) <= not(layer0_outputs(3045));
    outputs(7790) <= (layer0_outputs(11409)) and not (layer0_outputs(5250));
    outputs(7791) <= layer0_outputs(9975);
    outputs(7792) <= not(layer0_outputs(12073));
    outputs(7793) <= not(layer0_outputs(8746)) or (layer0_outputs(2526));
    outputs(7794) <= (layer0_outputs(11893)) and (layer0_outputs(6379));
    outputs(7795) <= not(layer0_outputs(8616));
    outputs(7796) <= layer0_outputs(6899);
    outputs(7797) <= (layer0_outputs(10490)) and not (layer0_outputs(11794));
    outputs(7798) <= (layer0_outputs(11853)) xor (layer0_outputs(573));
    outputs(7799) <= not(layer0_outputs(6382));
    outputs(7800) <= layer0_outputs(4865);
    outputs(7801) <= layer0_outputs(4460);
    outputs(7802) <= not(layer0_outputs(2523));
    outputs(7803) <= not(layer0_outputs(5097));
    outputs(7804) <= '1';
    outputs(7805) <= (layer0_outputs(8344)) and not (layer0_outputs(663));
    outputs(7806) <= not((layer0_outputs(5317)) and (layer0_outputs(4198)));
    outputs(7807) <= (layer0_outputs(7860)) xor (layer0_outputs(3662));
    outputs(7808) <= layer0_outputs(10598);
    outputs(7809) <= not((layer0_outputs(5575)) xor (layer0_outputs(7881)));
    outputs(7810) <= (layer0_outputs(11581)) or (layer0_outputs(613));
    outputs(7811) <= not(layer0_outputs(8040));
    outputs(7812) <= not((layer0_outputs(765)) xor (layer0_outputs(2270)));
    outputs(7813) <= (layer0_outputs(89)) and not (layer0_outputs(3233));
    outputs(7814) <= (layer0_outputs(4239)) xor (layer0_outputs(6890));
    outputs(7815) <= not(layer0_outputs(10456));
    outputs(7816) <= (layer0_outputs(12720)) xor (layer0_outputs(7264));
    outputs(7817) <= not((layer0_outputs(11472)) xor (layer0_outputs(7237)));
    outputs(7818) <= not((layer0_outputs(5174)) xor (layer0_outputs(5615)));
    outputs(7819) <= (layer0_outputs(9988)) xor (layer0_outputs(3896));
    outputs(7820) <= layer0_outputs(2933);
    outputs(7821) <= not(layer0_outputs(8788));
    outputs(7822) <= layer0_outputs(2192);
    outputs(7823) <= not(layer0_outputs(8327));
    outputs(7824) <= (layer0_outputs(680)) and not (layer0_outputs(3678));
    outputs(7825) <= not(layer0_outputs(8661));
    outputs(7826) <= layer0_outputs(4223);
    outputs(7827) <= (layer0_outputs(7712)) xor (layer0_outputs(8596));
    outputs(7828) <= not(layer0_outputs(7498)) or (layer0_outputs(6723));
    outputs(7829) <= (layer0_outputs(11208)) and not (layer0_outputs(12356));
    outputs(7830) <= (layer0_outputs(285)) xor (layer0_outputs(570));
    outputs(7831) <= not((layer0_outputs(11070)) xor (layer0_outputs(647)));
    outputs(7832) <= (layer0_outputs(9087)) xor (layer0_outputs(2264));
    outputs(7833) <= not(layer0_outputs(7199));
    outputs(7834) <= layer0_outputs(8981);
    outputs(7835) <= (layer0_outputs(406)) and (layer0_outputs(1148));
    outputs(7836) <= not((layer0_outputs(7894)) xor (layer0_outputs(1781)));
    outputs(7837) <= layer0_outputs(7150);
    outputs(7838) <= layer0_outputs(3693);
    outputs(7839) <= not(layer0_outputs(7500));
    outputs(7840) <= (layer0_outputs(9616)) and not (layer0_outputs(3013));
    outputs(7841) <= not((layer0_outputs(9314)) xor (layer0_outputs(5951)));
    outputs(7842) <= not(layer0_outputs(3066));
    outputs(7843) <= (layer0_outputs(444)) and not (layer0_outputs(6775));
    outputs(7844) <= (layer0_outputs(1758)) and not (layer0_outputs(2375));
    outputs(7845) <= not(layer0_outputs(2408));
    outputs(7846) <= not(layer0_outputs(9803));
    outputs(7847) <= not((layer0_outputs(9441)) xor (layer0_outputs(4699)));
    outputs(7848) <= not(layer0_outputs(9049));
    outputs(7849) <= not((layer0_outputs(7204)) xor (layer0_outputs(11252)));
    outputs(7850) <= not(layer0_outputs(4004));
    outputs(7851) <= layer0_outputs(7298);
    outputs(7852) <= not((layer0_outputs(12059)) xor (layer0_outputs(3768)));
    outputs(7853) <= layer0_outputs(2440);
    outputs(7854) <= not(layer0_outputs(9398));
    outputs(7855) <= (layer0_outputs(12738)) and (layer0_outputs(2057));
    outputs(7856) <= not((layer0_outputs(8234)) xor (layer0_outputs(7976)));
    outputs(7857) <= not(layer0_outputs(7823));
    outputs(7858) <= layer0_outputs(8735);
    outputs(7859) <= layer0_outputs(4017);
    outputs(7860) <= (layer0_outputs(770)) and not (layer0_outputs(4826));
    outputs(7861) <= layer0_outputs(2361);
    outputs(7862) <= (layer0_outputs(402)) xor (layer0_outputs(1752));
    outputs(7863) <= not(layer0_outputs(4714));
    outputs(7864) <= not((layer0_outputs(2492)) or (layer0_outputs(1918)));
    outputs(7865) <= layer0_outputs(2285);
    outputs(7866) <= layer0_outputs(8458);
    outputs(7867) <= layer0_outputs(88);
    outputs(7868) <= layer0_outputs(7681);
    outputs(7869) <= not((layer0_outputs(1798)) xor (layer0_outputs(11917)));
    outputs(7870) <= not(layer0_outputs(5127));
    outputs(7871) <= layer0_outputs(10919);
    outputs(7872) <= not(layer0_outputs(5245)) or (layer0_outputs(7878));
    outputs(7873) <= not(layer0_outputs(11746));
    outputs(7874) <= not(layer0_outputs(10988));
    outputs(7875) <= not(layer0_outputs(2950)) or (layer0_outputs(10780));
    outputs(7876) <= not(layer0_outputs(10553));
    outputs(7877) <= layer0_outputs(9357);
    outputs(7878) <= layer0_outputs(700);
    outputs(7879) <= not(layer0_outputs(7124));
    outputs(7880) <= (layer0_outputs(6724)) and (layer0_outputs(1235));
    outputs(7881) <= layer0_outputs(1014);
    outputs(7882) <= not((layer0_outputs(3881)) and (layer0_outputs(2891)));
    outputs(7883) <= (layer0_outputs(7352)) and not (layer0_outputs(4175));
    outputs(7884) <= not(layer0_outputs(11323));
    outputs(7885) <= not((layer0_outputs(12123)) or (layer0_outputs(10037)));
    outputs(7886) <= not(layer0_outputs(4520));
    outputs(7887) <= (layer0_outputs(4392)) and not (layer0_outputs(7595));
    outputs(7888) <= not(layer0_outputs(5853));
    outputs(7889) <= layer0_outputs(10219);
    outputs(7890) <= not(layer0_outputs(12275));
    outputs(7891) <= not(layer0_outputs(6571));
    outputs(7892) <= not((layer0_outputs(9631)) and (layer0_outputs(4621)));
    outputs(7893) <= (layer0_outputs(9741)) xor (layer0_outputs(11820));
    outputs(7894) <= layer0_outputs(9105);
    outputs(7895) <= (layer0_outputs(3536)) or (layer0_outputs(3563));
    outputs(7896) <= (layer0_outputs(4126)) xor (layer0_outputs(1684));
    outputs(7897) <= not((layer0_outputs(12538)) xor (layer0_outputs(10111)));
    outputs(7898) <= (layer0_outputs(7483)) xor (layer0_outputs(1266));
    outputs(7899) <= not((layer0_outputs(12633)) or (layer0_outputs(1534)));
    outputs(7900) <= not((layer0_outputs(9028)) xor (layer0_outputs(10807)));
    outputs(7901) <= '1';
    outputs(7902) <= not(layer0_outputs(292));
    outputs(7903) <= layer0_outputs(12460);
    outputs(7904) <= not(layer0_outputs(12714));
    outputs(7905) <= not((layer0_outputs(719)) xor (layer0_outputs(8713)));
    outputs(7906) <= layer0_outputs(179);
    outputs(7907) <= (layer0_outputs(9212)) xor (layer0_outputs(4515));
    outputs(7908) <= not((layer0_outputs(11941)) or (layer0_outputs(2154)));
    outputs(7909) <= not((layer0_outputs(9890)) xor (layer0_outputs(5508)));
    outputs(7910) <= not((layer0_outputs(10945)) or (layer0_outputs(11619)));
    outputs(7911) <= layer0_outputs(851);
    outputs(7912) <= not(layer0_outputs(175));
    outputs(7913) <= (layer0_outputs(4948)) and not (layer0_outputs(4535));
    outputs(7914) <= (layer0_outputs(10876)) xor (layer0_outputs(850));
    outputs(7915) <= layer0_outputs(1786);
    outputs(7916) <= (layer0_outputs(12637)) and (layer0_outputs(9131));
    outputs(7917) <= not(layer0_outputs(537));
    outputs(7918) <= layer0_outputs(4622);
    outputs(7919) <= not(layer0_outputs(5812));
    outputs(7920) <= not(layer0_outputs(3468));
    outputs(7921) <= layer0_outputs(10256);
    outputs(7922) <= not(layer0_outputs(8831));
    outputs(7923) <= not(layer0_outputs(8177)) or (layer0_outputs(9266));
    outputs(7924) <= not((layer0_outputs(1899)) xor (layer0_outputs(9995)));
    outputs(7925) <= not(layer0_outputs(7763));
    outputs(7926) <= layer0_outputs(12508);
    outputs(7927) <= not(layer0_outputs(9560));
    outputs(7928) <= not(layer0_outputs(3578));
    outputs(7929) <= not(layer0_outputs(8321));
    outputs(7930) <= (layer0_outputs(2447)) and not (layer0_outputs(3493));
    outputs(7931) <= not(layer0_outputs(4614)) or (layer0_outputs(5832));
    outputs(7932) <= not(layer0_outputs(7267));
    outputs(7933) <= '1';
    outputs(7934) <= layer0_outputs(2679);
    outputs(7935) <= not((layer0_outputs(2266)) or (layer0_outputs(11429)));
    outputs(7936) <= (layer0_outputs(9687)) xor (layer0_outputs(12026));
    outputs(7937) <= (layer0_outputs(1584)) and not (layer0_outputs(7833));
    outputs(7938) <= layer0_outputs(2712);
    outputs(7939) <= (layer0_outputs(6183)) or (layer0_outputs(11985));
    outputs(7940) <= layer0_outputs(1157);
    outputs(7941) <= not(layer0_outputs(6871));
    outputs(7942) <= layer0_outputs(4053);
    outputs(7943) <= layer0_outputs(11819);
    outputs(7944) <= (layer0_outputs(5813)) and not (layer0_outputs(9936));
    outputs(7945) <= not(layer0_outputs(7940));
    outputs(7946) <= not((layer0_outputs(5207)) xor (layer0_outputs(12198)));
    outputs(7947) <= (layer0_outputs(7274)) xor (layer0_outputs(5184));
    outputs(7948) <= layer0_outputs(4697);
    outputs(7949) <= layer0_outputs(11728);
    outputs(7950) <= (layer0_outputs(4131)) xor (layer0_outputs(4707));
    outputs(7951) <= not(layer0_outputs(1734));
    outputs(7952) <= (layer0_outputs(6454)) or (layer0_outputs(11934));
    outputs(7953) <= not(layer0_outputs(4984)) or (layer0_outputs(3555));
    outputs(7954) <= not(layer0_outputs(1593)) or (layer0_outputs(1499));
    outputs(7955) <= (layer0_outputs(12316)) or (layer0_outputs(12718));
    outputs(7956) <= not(layer0_outputs(1881));
    outputs(7957) <= not((layer0_outputs(9810)) xor (layer0_outputs(5433)));
    outputs(7958) <= (layer0_outputs(6824)) xor (layer0_outputs(8120));
    outputs(7959) <= '1';
    outputs(7960) <= not(layer0_outputs(7918));
    outputs(7961) <= (layer0_outputs(7631)) xor (layer0_outputs(1639));
    outputs(7962) <= (layer0_outputs(9840)) and not (layer0_outputs(12490));
    outputs(7963) <= layer0_outputs(3913);
    outputs(7964) <= not(layer0_outputs(6637));
    outputs(7965) <= layer0_outputs(5514);
    outputs(7966) <= (layer0_outputs(6034)) or (layer0_outputs(11283));
    outputs(7967) <= not(layer0_outputs(7376));
    outputs(7968) <= not(layer0_outputs(8731));
    outputs(7969) <= (layer0_outputs(9035)) xor (layer0_outputs(10474));
    outputs(7970) <= not((layer0_outputs(7211)) or (layer0_outputs(5468)));
    outputs(7971) <= not(layer0_outputs(10480));
    outputs(7972) <= not((layer0_outputs(673)) or (layer0_outputs(11429)));
    outputs(7973) <= not(layer0_outputs(9255)) or (layer0_outputs(4711));
    outputs(7974) <= (layer0_outputs(4840)) xor (layer0_outputs(4992));
    outputs(7975) <= (layer0_outputs(9337)) and not (layer0_outputs(10606));
    outputs(7976) <= not((layer0_outputs(1529)) or (layer0_outputs(9731)));
    outputs(7977) <= (layer0_outputs(9694)) and not (layer0_outputs(2811));
    outputs(7978) <= layer0_outputs(3338);
    outputs(7979) <= layer0_outputs(8487);
    outputs(7980) <= not(layer0_outputs(5054));
    outputs(7981) <= not((layer0_outputs(2056)) xor (layer0_outputs(429)));
    outputs(7982) <= (layer0_outputs(8890)) xor (layer0_outputs(7939));
    outputs(7983) <= not(layer0_outputs(9528));
    outputs(7984) <= not(layer0_outputs(248));
    outputs(7985) <= not(layer0_outputs(5614));
    outputs(7986) <= not(layer0_outputs(5590));
    outputs(7987) <= not((layer0_outputs(4700)) xor (layer0_outputs(11632)));
    outputs(7988) <= layer0_outputs(5523);
    outputs(7989) <= (layer0_outputs(8297)) xor (layer0_outputs(1816));
    outputs(7990) <= (layer0_outputs(9708)) or (layer0_outputs(10730));
    outputs(7991) <= not(layer0_outputs(11260));
    outputs(7992) <= not(layer0_outputs(3100));
    outputs(7993) <= (layer0_outputs(1909)) xor (layer0_outputs(10655));
    outputs(7994) <= not((layer0_outputs(811)) xor (layer0_outputs(6810)));
    outputs(7995) <= not(layer0_outputs(4765));
    outputs(7996) <= (layer0_outputs(4966)) or (layer0_outputs(12472));
    outputs(7997) <= layer0_outputs(11312);
    outputs(7998) <= (layer0_outputs(5284)) xor (layer0_outputs(3058));
    outputs(7999) <= not((layer0_outputs(11581)) xor (layer0_outputs(2522)));
    outputs(8000) <= not(layer0_outputs(11573));
    outputs(8001) <= layer0_outputs(10396);
    outputs(8002) <= (layer0_outputs(227)) xor (layer0_outputs(11389));
    outputs(8003) <= not(layer0_outputs(4390));
    outputs(8004) <= not(layer0_outputs(6870));
    outputs(8005) <= not((layer0_outputs(2077)) xor (layer0_outputs(2794)));
    outputs(8006) <= not(layer0_outputs(2659));
    outputs(8007) <= layer0_outputs(3638);
    outputs(8008) <= not((layer0_outputs(10064)) or (layer0_outputs(1996)));
    outputs(8009) <= not((layer0_outputs(11023)) xor (layer0_outputs(1977)));
    outputs(8010) <= layer0_outputs(5597);
    outputs(8011) <= not(layer0_outputs(2764));
    outputs(8012) <= not((layer0_outputs(315)) or (layer0_outputs(12067)));
    outputs(8013) <= layer0_outputs(569);
    outputs(8014) <= not((layer0_outputs(11077)) or (layer0_outputs(7570)));
    outputs(8015) <= layer0_outputs(2033);
    outputs(8016) <= (layer0_outputs(3984)) and not (layer0_outputs(9279));
    outputs(8017) <= not((layer0_outputs(12168)) xor (layer0_outputs(3861)));
    outputs(8018) <= (layer0_outputs(9123)) xor (layer0_outputs(3845));
    outputs(8019) <= not(layer0_outputs(5182)) or (layer0_outputs(2647));
    outputs(8020) <= not(layer0_outputs(5447));
    outputs(8021) <= not((layer0_outputs(6567)) or (layer0_outputs(3114)));
    outputs(8022) <= not(layer0_outputs(12457));
    outputs(8023) <= not(layer0_outputs(5015));
    outputs(8024) <= not(layer0_outputs(4454));
    outputs(8025) <= not((layer0_outputs(4643)) or (layer0_outputs(1700)));
    outputs(8026) <= not(layer0_outputs(10416)) or (layer0_outputs(11155));
    outputs(8027) <= (layer0_outputs(10608)) or (layer0_outputs(10666));
    outputs(8028) <= (layer0_outputs(11634)) xor (layer0_outputs(10717));
    outputs(8029) <= not(layer0_outputs(6600));
    outputs(8030) <= layer0_outputs(10921);
    outputs(8031) <= (layer0_outputs(6606)) and (layer0_outputs(223));
    outputs(8032) <= layer0_outputs(5513);
    outputs(8033) <= (layer0_outputs(2189)) xor (layer0_outputs(6811));
    outputs(8034) <= (layer0_outputs(173)) or (layer0_outputs(11501));
    outputs(8035) <= layer0_outputs(11245);
    outputs(8036) <= layer0_outputs(12373);
    outputs(8037) <= (layer0_outputs(5682)) and not (layer0_outputs(9183));
    outputs(8038) <= (layer0_outputs(12362)) xor (layer0_outputs(5560));
    outputs(8039) <= not((layer0_outputs(3772)) or (layer0_outputs(5321)));
    outputs(8040) <= (layer0_outputs(1816)) xor (layer0_outputs(4629));
    outputs(8041) <= layer0_outputs(10525);
    outputs(8042) <= not((layer0_outputs(2386)) or (layer0_outputs(8778)));
    outputs(8043) <= layer0_outputs(708);
    outputs(8044) <= layer0_outputs(8958);
    outputs(8045) <= not((layer0_outputs(6756)) xor (layer0_outputs(2653)));
    outputs(8046) <= layer0_outputs(7843);
    outputs(8047) <= not(layer0_outputs(8255));
    outputs(8048) <= not(layer0_outputs(2327));
    outputs(8049) <= not(layer0_outputs(733));
    outputs(8050) <= not(layer0_outputs(5413));
    outputs(8051) <= not((layer0_outputs(6029)) or (layer0_outputs(8553)));
    outputs(8052) <= (layer0_outputs(3236)) and not (layer0_outputs(1051));
    outputs(8053) <= not((layer0_outputs(8356)) or (layer0_outputs(161)));
    outputs(8054) <= not(layer0_outputs(1996)) or (layer0_outputs(6765));
    outputs(8055) <= layer0_outputs(3461);
    outputs(8056) <= (layer0_outputs(1426)) and not (layer0_outputs(6366));
    outputs(8057) <= layer0_outputs(88);
    outputs(8058) <= layer0_outputs(1873);
    outputs(8059) <= (layer0_outputs(9474)) and (layer0_outputs(4882));
    outputs(8060) <= not((layer0_outputs(2433)) or (layer0_outputs(6766)));
    outputs(8061) <= not((layer0_outputs(6798)) xor (layer0_outputs(6941)));
    outputs(8062) <= layer0_outputs(5790);
    outputs(8063) <= not((layer0_outputs(5660)) xor (layer0_outputs(10030)));
    outputs(8064) <= not(layer0_outputs(7479)) or (layer0_outputs(8874));
    outputs(8065) <= not(layer0_outputs(4408));
    outputs(8066) <= layer0_outputs(11994);
    outputs(8067) <= not((layer0_outputs(12472)) xor (layer0_outputs(7589)));
    outputs(8068) <= not(layer0_outputs(6608));
    outputs(8069) <= layer0_outputs(5386);
    outputs(8070) <= (layer0_outputs(2493)) or (layer0_outputs(464));
    outputs(8071) <= layer0_outputs(11867);
    outputs(8072) <= not((layer0_outputs(641)) or (layer0_outputs(8077)));
    outputs(8073) <= layer0_outputs(7539);
    outputs(8074) <= not((layer0_outputs(10264)) xor (layer0_outputs(9081)));
    outputs(8075) <= not(layer0_outputs(9783)) or (layer0_outputs(3458));
    outputs(8076) <= not(layer0_outputs(66)) or (layer0_outputs(8600));
    outputs(8077) <= layer0_outputs(11568);
    outputs(8078) <= not(layer0_outputs(10622));
    outputs(8079) <= not(layer0_outputs(7706)) or (layer0_outputs(2119));
    outputs(8080) <= not(layer0_outputs(1025));
    outputs(8081) <= not(layer0_outputs(12374)) or (layer0_outputs(3048));
    outputs(8082) <= layer0_outputs(3871);
    outputs(8083) <= not(layer0_outputs(11723));
    outputs(8084) <= (layer0_outputs(3936)) xor (layer0_outputs(10367));
    outputs(8085) <= not(layer0_outputs(9297));
    outputs(8086) <= (layer0_outputs(10301)) or (layer0_outputs(2166));
    outputs(8087) <= not((layer0_outputs(3448)) xor (layer0_outputs(7559)));
    outputs(8088) <= (layer0_outputs(5978)) xor (layer0_outputs(4065));
    outputs(8089) <= (layer0_outputs(12563)) xor (layer0_outputs(9535));
    outputs(8090) <= not(layer0_outputs(5211));
    outputs(8091) <= (layer0_outputs(6048)) xor (layer0_outputs(10437));
    outputs(8092) <= not((layer0_outputs(334)) and (layer0_outputs(5593)));
    outputs(8093) <= not((layer0_outputs(12065)) xor (layer0_outputs(10288)));
    outputs(8094) <= not(layer0_outputs(7788));
    outputs(8095) <= not(layer0_outputs(2513));
    outputs(8096) <= (layer0_outputs(9755)) and (layer0_outputs(12150));
    outputs(8097) <= layer0_outputs(10663);
    outputs(8098) <= not((layer0_outputs(1702)) xor (layer0_outputs(1930)));
    outputs(8099) <= not(layer0_outputs(997));
    outputs(8100) <= not(layer0_outputs(6927)) or (layer0_outputs(12701));
    outputs(8101) <= layer0_outputs(8816);
    outputs(8102) <= not(layer0_outputs(4283));
    outputs(8103) <= (layer0_outputs(8364)) or (layer0_outputs(2212));
    outputs(8104) <= layer0_outputs(426);
    outputs(8105) <= not((layer0_outputs(3147)) xor (layer0_outputs(2671)));
    outputs(8106) <= layer0_outputs(3149);
    outputs(8107) <= (layer0_outputs(3460)) and (layer0_outputs(1555));
    outputs(8108) <= not(layer0_outputs(10433));
    outputs(8109) <= (layer0_outputs(11069)) or (layer0_outputs(12513));
    outputs(8110) <= layer0_outputs(3816);
    outputs(8111) <= not(layer0_outputs(5127));
    outputs(8112) <= not((layer0_outputs(12555)) and (layer0_outputs(7617)));
    outputs(8113) <= not(layer0_outputs(2819)) or (layer0_outputs(8686));
    outputs(8114) <= not((layer0_outputs(5346)) and (layer0_outputs(1798)));
    outputs(8115) <= (layer0_outputs(5679)) and not (layer0_outputs(8432));
    outputs(8116) <= not((layer0_outputs(7773)) or (layer0_outputs(6117)));
    outputs(8117) <= layer0_outputs(12066);
    outputs(8118) <= (layer0_outputs(9444)) and (layer0_outputs(11907));
    outputs(8119) <= (layer0_outputs(12478)) xor (layer0_outputs(3458));
    outputs(8120) <= layer0_outputs(3262);
    outputs(8121) <= layer0_outputs(12679);
    outputs(8122) <= (layer0_outputs(964)) xor (layer0_outputs(5064));
    outputs(8123) <= not((layer0_outputs(535)) xor (layer0_outputs(9339)));
    outputs(8124) <= not(layer0_outputs(5811)) or (layer0_outputs(8243));
    outputs(8125) <= not(layer0_outputs(11477));
    outputs(8126) <= layer0_outputs(7527);
    outputs(8127) <= not(layer0_outputs(1388)) or (layer0_outputs(7139));
    outputs(8128) <= (layer0_outputs(12698)) and not (layer0_outputs(5143));
    outputs(8129) <= (layer0_outputs(12540)) xor (layer0_outputs(12118));
    outputs(8130) <= not(layer0_outputs(5577));
    outputs(8131) <= not(layer0_outputs(5920)) or (layer0_outputs(8225));
    outputs(8132) <= (layer0_outputs(11483)) and not (layer0_outputs(6932));
    outputs(8133) <= not(layer0_outputs(5456));
    outputs(8134) <= not((layer0_outputs(1141)) xor (layer0_outputs(8372)));
    outputs(8135) <= not(layer0_outputs(10457));
    outputs(8136) <= not(layer0_outputs(772));
    outputs(8137) <= layer0_outputs(575);
    outputs(8138) <= (layer0_outputs(12054)) xor (layer0_outputs(3245));
    outputs(8139) <= (layer0_outputs(12549)) xor (layer0_outputs(10319));
    outputs(8140) <= not(layer0_outputs(5321));
    outputs(8141) <= (layer0_outputs(1784)) and (layer0_outputs(12052));
    outputs(8142) <= (layer0_outputs(9450)) xor (layer0_outputs(972));
    outputs(8143) <= (layer0_outputs(11127)) and (layer0_outputs(4057));
    outputs(8144) <= layer0_outputs(12031);
    outputs(8145) <= layer0_outputs(1807);
    outputs(8146) <= (layer0_outputs(10673)) xor (layer0_outputs(4934));
    outputs(8147) <= not((layer0_outputs(3752)) xor (layer0_outputs(390)));
    outputs(8148) <= (layer0_outputs(9981)) xor (layer0_outputs(9158));
    outputs(8149) <= not(layer0_outputs(1598));
    outputs(8150) <= not(layer0_outputs(11401));
    outputs(8151) <= (layer0_outputs(1604)) xor (layer0_outputs(2332));
    outputs(8152) <= layer0_outputs(3010);
    outputs(8153) <= layer0_outputs(1116);
    outputs(8154) <= (layer0_outputs(5583)) and not (layer0_outputs(4494));
    outputs(8155) <= (layer0_outputs(8144)) and not (layer0_outputs(10875));
    outputs(8156) <= not(layer0_outputs(5890));
    outputs(8157) <= (layer0_outputs(10283)) xor (layer0_outputs(9787));
    outputs(8158) <= not(layer0_outputs(7577));
    outputs(8159) <= (layer0_outputs(12490)) and (layer0_outputs(6519));
    outputs(8160) <= (layer0_outputs(10032)) and (layer0_outputs(6731));
    outputs(8161) <= (layer0_outputs(11264)) xor (layer0_outputs(7161));
    outputs(8162) <= not(layer0_outputs(7828));
    outputs(8163) <= not(layer0_outputs(5496));
    outputs(8164) <= layer0_outputs(7118);
    outputs(8165) <= (layer0_outputs(1141)) xor (layer0_outputs(6627));
    outputs(8166) <= (layer0_outputs(3604)) and not (layer0_outputs(4837));
    outputs(8167) <= (layer0_outputs(9580)) xor (layer0_outputs(5009));
    outputs(8168) <= not(layer0_outputs(6099));
    outputs(8169) <= not(layer0_outputs(11425));
    outputs(8170) <= layer0_outputs(8397);
    outputs(8171) <= not((layer0_outputs(5193)) xor (layer0_outputs(10360)));
    outputs(8172) <= layer0_outputs(9943);
    outputs(8173) <= not((layer0_outputs(6390)) xor (layer0_outputs(3804)));
    outputs(8174) <= not((layer0_outputs(10665)) xor (layer0_outputs(10668)));
    outputs(8175) <= not((layer0_outputs(3079)) and (layer0_outputs(2537)));
    outputs(8176) <= (layer0_outputs(9599)) or (layer0_outputs(3432));
    outputs(8177) <= not(layer0_outputs(10882)) or (layer0_outputs(3589));
    outputs(8178) <= not(layer0_outputs(12541));
    outputs(8179) <= not(layer0_outputs(9790));
    outputs(8180) <= not((layer0_outputs(11815)) xor (layer0_outputs(9145)));
    outputs(8181) <= not(layer0_outputs(4048));
    outputs(8182) <= not(layer0_outputs(7170));
    outputs(8183) <= not((layer0_outputs(9837)) and (layer0_outputs(10789)));
    outputs(8184) <= not(layer0_outputs(12274));
    outputs(8185) <= layer0_outputs(735);
    outputs(8186) <= not((layer0_outputs(9010)) xor (layer0_outputs(6399)));
    outputs(8187) <= (layer0_outputs(238)) and (layer0_outputs(11698));
    outputs(8188) <= (layer0_outputs(6117)) and not (layer0_outputs(2644));
    outputs(8189) <= not((layer0_outputs(10867)) xor (layer0_outputs(2625)));
    outputs(8190) <= not(layer0_outputs(7022));
    outputs(8191) <= layer0_outputs(12166);
    outputs(8192) <= not((layer0_outputs(4093)) xor (layer0_outputs(2407)));
    outputs(8193) <= not((layer0_outputs(10554)) xor (layer0_outputs(3444)));
    outputs(8194) <= not((layer0_outputs(2176)) xor (layer0_outputs(6760)));
    outputs(8195) <= (layer0_outputs(4257)) and (layer0_outputs(2453));
    outputs(8196) <= (layer0_outputs(569)) and not (layer0_outputs(11281));
    outputs(8197) <= not((layer0_outputs(2988)) xor (layer0_outputs(409)));
    outputs(8198) <= layer0_outputs(3253);
    outputs(8199) <= layer0_outputs(1624);
    outputs(8200) <= not(layer0_outputs(11825));
    outputs(8201) <= layer0_outputs(11557);
    outputs(8202) <= not(layer0_outputs(5808));
    outputs(8203) <= not(layer0_outputs(6726));
    outputs(8204) <= layer0_outputs(6570);
    outputs(8205) <= not(layer0_outputs(800));
    outputs(8206) <= layer0_outputs(3167);
    outputs(8207) <= not(layer0_outputs(6690)) or (layer0_outputs(10254));
    outputs(8208) <= (layer0_outputs(2014)) and not (layer0_outputs(2340));
    outputs(8209) <= layer0_outputs(11296);
    outputs(8210) <= layer0_outputs(1293);
    outputs(8211) <= not(layer0_outputs(4611));
    outputs(8212) <= layer0_outputs(1931);
    outputs(8213) <= not(layer0_outputs(12743));
    outputs(8214) <= '1';
    outputs(8215) <= not(layer0_outputs(1926));
    outputs(8216) <= layer0_outputs(4240);
    outputs(8217) <= not((layer0_outputs(11599)) or (layer0_outputs(7600)));
    outputs(8218) <= not(layer0_outputs(4089));
    outputs(8219) <= not(layer0_outputs(1492));
    outputs(8220) <= (layer0_outputs(6431)) xor (layer0_outputs(1093));
    outputs(8221) <= (layer0_outputs(2715)) xor (layer0_outputs(10423));
    outputs(8222) <= not((layer0_outputs(581)) xor (layer0_outputs(4128)));
    outputs(8223) <= not(layer0_outputs(2908));
    outputs(8224) <= not(layer0_outputs(6496)) or (layer0_outputs(12276));
    outputs(8225) <= not((layer0_outputs(3661)) xor (layer0_outputs(8091)));
    outputs(8226) <= (layer0_outputs(12444)) or (layer0_outputs(9664));
    outputs(8227) <= layer0_outputs(5056);
    outputs(8228) <= (layer0_outputs(5460)) xor (layer0_outputs(6029));
    outputs(8229) <= not((layer0_outputs(141)) xor (layer0_outputs(2588)));
    outputs(8230) <= not(layer0_outputs(71));
    outputs(8231) <= layer0_outputs(5761);
    outputs(8232) <= not(layer0_outputs(8494));
    outputs(8233) <= (layer0_outputs(1887)) xor (layer0_outputs(10395));
    outputs(8234) <= not(layer0_outputs(3707)) or (layer0_outputs(8442));
    outputs(8235) <= (layer0_outputs(7832)) xor (layer0_outputs(11873));
    outputs(8236) <= (layer0_outputs(12539)) xor (layer0_outputs(3485));
    outputs(8237) <= not((layer0_outputs(1567)) or (layer0_outputs(7417)));
    outputs(8238) <= (layer0_outputs(11767)) or (layer0_outputs(5430));
    outputs(8239) <= not((layer0_outputs(4841)) xor (layer0_outputs(8727)));
    outputs(8240) <= not(layer0_outputs(10151));
    outputs(8241) <= not(layer0_outputs(5415));
    outputs(8242) <= (layer0_outputs(8170)) xor (layer0_outputs(8100));
    outputs(8243) <= (layer0_outputs(3190)) and (layer0_outputs(1395));
    outputs(8244) <= not(layer0_outputs(3333));
    outputs(8245) <= layer0_outputs(9252);
    outputs(8246) <= not(layer0_outputs(9587)) or (layer0_outputs(5859));
    outputs(8247) <= not(layer0_outputs(5934));
    outputs(8248) <= not((layer0_outputs(8882)) or (layer0_outputs(4833)));
    outputs(8249) <= not(layer0_outputs(5797));
    outputs(8250) <= (layer0_outputs(8664)) xor (layer0_outputs(2315));
    outputs(8251) <= not(layer0_outputs(8146));
    outputs(8252) <= (layer0_outputs(4577)) xor (layer0_outputs(1485));
    outputs(8253) <= (layer0_outputs(8822)) and not (layer0_outputs(9390));
    outputs(8254) <= (layer0_outputs(10507)) xor (layer0_outputs(5206));
    outputs(8255) <= (layer0_outputs(5846)) and not (layer0_outputs(12683));
    outputs(8256) <= not(layer0_outputs(12501));
    outputs(8257) <= not(layer0_outputs(2754));
    outputs(8258) <= layer0_outputs(7313);
    outputs(8259) <= layer0_outputs(9109);
    outputs(8260) <= not(layer0_outputs(1078));
    outputs(8261) <= (layer0_outputs(5500)) and not (layer0_outputs(4570));
    outputs(8262) <= layer0_outputs(2172);
    outputs(8263) <= not(layer0_outputs(9963));
    outputs(8264) <= layer0_outputs(11528);
    outputs(8265) <= layer0_outputs(9759);
    outputs(8266) <= not(layer0_outputs(6398));
    outputs(8267) <= not((layer0_outputs(6657)) and (layer0_outputs(4605)));
    outputs(8268) <= not((layer0_outputs(6855)) xor (layer0_outputs(4671)));
    outputs(8269) <= not((layer0_outputs(367)) xor (layer0_outputs(10899)));
    outputs(8270) <= (layer0_outputs(10690)) and not (layer0_outputs(12696));
    outputs(8271) <= not(layer0_outputs(2787));
    outputs(8272) <= not(layer0_outputs(4073)) or (layer0_outputs(10383));
    outputs(8273) <= not((layer0_outputs(8922)) or (layer0_outputs(891)));
    outputs(8274) <= not((layer0_outputs(2421)) xor (layer0_outputs(2351)));
    outputs(8275) <= (layer0_outputs(7062)) xor (layer0_outputs(6063));
    outputs(8276) <= not(layer0_outputs(6503));
    outputs(8277) <= layer0_outputs(7481);
    outputs(8278) <= layer0_outputs(10805);
    outputs(8279) <= not(layer0_outputs(4482));
    outputs(8280) <= layer0_outputs(5171);
    outputs(8281) <= layer0_outputs(7207);
    outputs(8282) <= layer0_outputs(9594);
    outputs(8283) <= not((layer0_outputs(11447)) xor (layer0_outputs(2426)));
    outputs(8284) <= not(layer0_outputs(2168));
    outputs(8285) <= (layer0_outputs(9219)) and not (layer0_outputs(1194));
    outputs(8286) <= layer0_outputs(9090);
    outputs(8287) <= (layer0_outputs(3474)) and (layer0_outputs(480));
    outputs(8288) <= not(layer0_outputs(3480));
    outputs(8289) <= (layer0_outputs(2324)) xor (layer0_outputs(716));
    outputs(8290) <= layer0_outputs(5276);
    outputs(8291) <= not(layer0_outputs(6151));
    outputs(8292) <= layer0_outputs(8235);
    outputs(8293) <= layer0_outputs(648);
    outputs(8294) <= not((layer0_outputs(4785)) xor (layer0_outputs(4472)));
    outputs(8295) <= not((layer0_outputs(4177)) xor (layer0_outputs(6291)));
    outputs(8296) <= not(layer0_outputs(8110));
    outputs(8297) <= (layer0_outputs(6185)) or (layer0_outputs(11782));
    outputs(8298) <= layer0_outputs(11652);
    outputs(8299) <= (layer0_outputs(11626)) xor (layer0_outputs(12021));
    outputs(8300) <= layer0_outputs(9361);
    outputs(8301) <= not((layer0_outputs(2479)) xor (layer0_outputs(10161)));
    outputs(8302) <= not((layer0_outputs(6038)) xor (layer0_outputs(4992)));
    outputs(8303) <= not(layer0_outputs(10327));
    outputs(8304) <= not(layer0_outputs(7311));
    outputs(8305) <= layer0_outputs(3193);
    outputs(8306) <= not((layer0_outputs(502)) xor (layer0_outputs(12469)));
    outputs(8307) <= (layer0_outputs(7632)) xor (layer0_outputs(1992));
    outputs(8308) <= layer0_outputs(2088);
    outputs(8309) <= not((layer0_outputs(12689)) xor (layer0_outputs(4634)));
    outputs(8310) <= not(layer0_outputs(8643));
    outputs(8311) <= (layer0_outputs(4445)) xor (layer0_outputs(10393));
    outputs(8312) <= (layer0_outputs(7607)) xor (layer0_outputs(5439));
    outputs(8313) <= '0';
    outputs(8314) <= not((layer0_outputs(1062)) xor (layer0_outputs(4931)));
    outputs(8315) <= not((layer0_outputs(8579)) xor (layer0_outputs(9156)));
    outputs(8316) <= layer0_outputs(5630);
    outputs(8317) <= not((layer0_outputs(6650)) and (layer0_outputs(8866)));
    outputs(8318) <= (layer0_outputs(5807)) and not (layer0_outputs(12676));
    outputs(8319) <= (layer0_outputs(2645)) and not (layer0_outputs(7417));
    outputs(8320) <= not(layer0_outputs(6471)) or (layer0_outputs(10855));
    outputs(8321) <= not((layer0_outputs(12699)) xor (layer0_outputs(6991)));
    outputs(8322) <= not(layer0_outputs(8033));
    outputs(8323) <= (layer0_outputs(793)) and not (layer0_outputs(9520));
    outputs(8324) <= (layer0_outputs(7393)) xor (layer0_outputs(7254));
    outputs(8325) <= layer0_outputs(11204);
    outputs(8326) <= not(layer0_outputs(7745));
    outputs(8327) <= layer0_outputs(2722);
    outputs(8328) <= not(layer0_outputs(6498));
    outputs(8329) <= '1';
    outputs(8330) <= layer0_outputs(3883);
    outputs(8331) <= not(layer0_outputs(7345));
    outputs(8332) <= not((layer0_outputs(12602)) xor (layer0_outputs(453)));
    outputs(8333) <= (layer0_outputs(6523)) xor (layer0_outputs(12632));
    outputs(8334) <= (layer0_outputs(11807)) xor (layer0_outputs(7377));
    outputs(8335) <= not(layer0_outputs(9455));
    outputs(8336) <= not((layer0_outputs(3889)) xor (layer0_outputs(5425)));
    outputs(8337) <= not(layer0_outputs(4276));
    outputs(8338) <= layer0_outputs(4579);
    outputs(8339) <= layer0_outputs(2874);
    outputs(8340) <= not((layer0_outputs(10292)) and (layer0_outputs(7640)));
    outputs(8341) <= (layer0_outputs(12480)) and not (layer0_outputs(1446));
    outputs(8342) <= layer0_outputs(7102);
    outputs(8343) <= not(layer0_outputs(2627)) or (layer0_outputs(5700));
    outputs(8344) <= layer0_outputs(3749);
    outputs(8345) <= not((layer0_outputs(1754)) and (layer0_outputs(11921)));
    outputs(8346) <= not(layer0_outputs(1437));
    outputs(8347) <= layer0_outputs(5457);
    outputs(8348) <= not((layer0_outputs(7829)) xor (layer0_outputs(12132)));
    outputs(8349) <= not(layer0_outputs(12092));
    outputs(8350) <= not((layer0_outputs(6760)) xor (layer0_outputs(271)));
    outputs(8351) <= layer0_outputs(4505);
    outputs(8352) <= not((layer0_outputs(7994)) and (layer0_outputs(7558)));
    outputs(8353) <= (layer0_outputs(7242)) or (layer0_outputs(1039));
    outputs(8354) <= not(layer0_outputs(4786));
    outputs(8355) <= layer0_outputs(11182);
    outputs(8356) <= not(layer0_outputs(4760));
    outputs(8357) <= not((layer0_outputs(9879)) or (layer0_outputs(9660)));
    outputs(8358) <= not((layer0_outputs(6879)) xor (layer0_outputs(704)));
    outputs(8359) <= not((layer0_outputs(8934)) xor (layer0_outputs(7542)));
    outputs(8360) <= not((layer0_outputs(9743)) xor (layer0_outputs(1436)));
    outputs(8361) <= layer0_outputs(5239);
    outputs(8362) <= (layer0_outputs(3983)) xor (layer0_outputs(4089));
    outputs(8363) <= not((layer0_outputs(10513)) xor (layer0_outputs(10563)));
    outputs(8364) <= (layer0_outputs(4289)) and (layer0_outputs(9411));
    outputs(8365) <= not(layer0_outputs(9459));
    outputs(8366) <= not(layer0_outputs(12101));
    outputs(8367) <= not((layer0_outputs(8634)) xor (layer0_outputs(7830)));
    outputs(8368) <= not(layer0_outputs(908));
    outputs(8369) <= not(layer0_outputs(3457));
    outputs(8370) <= not((layer0_outputs(7307)) and (layer0_outputs(3027)));
    outputs(8371) <= layer0_outputs(7236);
    outputs(8372) <= layer0_outputs(12782);
    outputs(8373) <= layer0_outputs(3926);
    outputs(8374) <= (layer0_outputs(11363)) and not (layer0_outputs(8513));
    outputs(8375) <= not((layer0_outputs(1076)) xor (layer0_outputs(6747)));
    outputs(8376) <= not((layer0_outputs(6970)) xor (layer0_outputs(3506)));
    outputs(8377) <= not(layer0_outputs(7369));
    outputs(8378) <= not(layer0_outputs(1494));
    outputs(8379) <= not((layer0_outputs(8486)) and (layer0_outputs(5728)));
    outputs(8380) <= layer0_outputs(9844);
    outputs(8381) <= layer0_outputs(4457);
    outputs(8382) <= (layer0_outputs(5085)) and not (layer0_outputs(4379));
    outputs(8383) <= not(layer0_outputs(4143));
    outputs(8384) <= not(layer0_outputs(7785));
    outputs(8385) <= (layer0_outputs(8351)) xor (layer0_outputs(6468));
    outputs(8386) <= layer0_outputs(3054);
    outputs(8387) <= layer0_outputs(2233);
    outputs(8388) <= not(layer0_outputs(1040));
    outputs(8389) <= not(layer0_outputs(3856));
    outputs(8390) <= not((layer0_outputs(6040)) or (layer0_outputs(2900)));
    outputs(8391) <= layer0_outputs(6743);
    outputs(8392) <= (layer0_outputs(12573)) and not (layer0_outputs(12664));
    outputs(8393) <= not((layer0_outputs(2413)) xor (layer0_outputs(4040)));
    outputs(8394) <= layer0_outputs(10512);
    outputs(8395) <= (layer0_outputs(12498)) xor (layer0_outputs(5785));
    outputs(8396) <= layer0_outputs(8126);
    outputs(8397) <= layer0_outputs(9700);
    outputs(8398) <= (layer0_outputs(12263)) xor (layer0_outputs(9963));
    outputs(8399) <= not((layer0_outputs(12761)) and (layer0_outputs(499)));
    outputs(8400) <= layer0_outputs(12627);
    outputs(8401) <= (layer0_outputs(11421)) and not (layer0_outputs(6131));
    outputs(8402) <= not(layer0_outputs(11420));
    outputs(8403) <= not((layer0_outputs(5678)) xor (layer0_outputs(7101)));
    outputs(8404) <= not(layer0_outputs(9767));
    outputs(8405) <= not((layer0_outputs(6802)) and (layer0_outputs(6057)));
    outputs(8406) <= layer0_outputs(5270);
    outputs(8407) <= (layer0_outputs(11655)) or (layer0_outputs(4247));
    outputs(8408) <= layer0_outputs(8274);
    outputs(8409) <= (layer0_outputs(6103)) or (layer0_outputs(5187));
    outputs(8410) <= (layer0_outputs(8218)) xor (layer0_outputs(8928));
    outputs(8411) <= (layer0_outputs(10340)) and not (layer0_outputs(306));
    outputs(8412) <= not((layer0_outputs(10659)) xor (layer0_outputs(181)));
    outputs(8413) <= layer0_outputs(7047);
    outputs(8414) <= (layer0_outputs(1065)) xor (layer0_outputs(5669));
    outputs(8415) <= (layer0_outputs(6514)) and not (layer0_outputs(5952));
    outputs(8416) <= layer0_outputs(8508);
    outputs(8417) <= layer0_outputs(3296);
    outputs(8418) <= (layer0_outputs(7948)) and not (layer0_outputs(1734));
    outputs(8419) <= (layer0_outputs(2979)) and not (layer0_outputs(9782));
    outputs(8420) <= (layer0_outputs(2968)) xor (layer0_outputs(11394));
    outputs(8421) <= (layer0_outputs(4743)) and not (layer0_outputs(8323));
    outputs(8422) <= (layer0_outputs(7764)) xor (layer0_outputs(9965));
    outputs(8423) <= not((layer0_outputs(1603)) or (layer0_outputs(30)));
    outputs(8424) <= (layer0_outputs(6857)) xor (layer0_outputs(2937));
    outputs(8425) <= not((layer0_outputs(8930)) xor (layer0_outputs(2279)));
    outputs(8426) <= not((layer0_outputs(12435)) xor (layer0_outputs(12696)));
    outputs(8427) <= not(layer0_outputs(9985));
    outputs(8428) <= (layer0_outputs(1638)) and (layer0_outputs(8439));
    outputs(8429) <= (layer0_outputs(7171)) xor (layer0_outputs(477));
    outputs(8430) <= not((layer0_outputs(10503)) xor (layer0_outputs(3173)));
    outputs(8431) <= (layer0_outputs(11451)) and (layer0_outputs(12533));
    outputs(8432) <= not(layer0_outputs(11360));
    outputs(8433) <= not((layer0_outputs(8029)) xor (layer0_outputs(9215)));
    outputs(8434) <= not(layer0_outputs(7978));
    outputs(8435) <= not(layer0_outputs(11722)) or (layer0_outputs(5742));
    outputs(8436) <= not((layer0_outputs(458)) and (layer0_outputs(3027)));
    outputs(8437) <= (layer0_outputs(6784)) and (layer0_outputs(4750));
    outputs(8438) <= (layer0_outputs(1886)) xor (layer0_outputs(7841));
    outputs(8439) <= not((layer0_outputs(11412)) xor (layer0_outputs(1154)));
    outputs(8440) <= layer0_outputs(10228);
    outputs(8441) <= not((layer0_outputs(6639)) xor (layer0_outputs(10036)));
    outputs(8442) <= layer0_outputs(5395);
    outputs(8443) <= not((layer0_outputs(1956)) or (layer0_outputs(10222)));
    outputs(8444) <= layer0_outputs(4545);
    outputs(8445) <= not((layer0_outputs(485)) or (layer0_outputs(10344)));
    outputs(8446) <= not((layer0_outputs(8857)) xor (layer0_outputs(1473)));
    outputs(8447) <= not(layer0_outputs(5996));
    outputs(8448) <= not(layer0_outputs(8739));
    outputs(8449) <= layer0_outputs(8505);
    outputs(8450) <= not(layer0_outputs(9798));
    outputs(8451) <= not((layer0_outputs(9901)) xor (layer0_outputs(5047)));
    outputs(8452) <= (layer0_outputs(462)) and not (layer0_outputs(10443));
    outputs(8453) <= layer0_outputs(11505);
    outputs(8454) <= (layer0_outputs(4824)) and not (layer0_outputs(4589));
    outputs(8455) <= not((layer0_outputs(10441)) and (layer0_outputs(7408)));
    outputs(8456) <= (layer0_outputs(1615)) and not (layer0_outputs(5503));
    outputs(8457) <= not((layer0_outputs(4284)) and (layer0_outputs(1871)));
    outputs(8458) <= (layer0_outputs(9830)) and not (layer0_outputs(7966));
    outputs(8459) <= not(layer0_outputs(4905));
    outputs(8460) <= layer0_outputs(505);
    outputs(8461) <= (layer0_outputs(4305)) xor (layer0_outputs(10413));
    outputs(8462) <= not((layer0_outputs(3995)) or (layer0_outputs(8268)));
    outputs(8463) <= (layer0_outputs(4281)) xor (layer0_outputs(9277));
    outputs(8464) <= (layer0_outputs(2178)) xor (layer0_outputs(6381));
    outputs(8465) <= not(layer0_outputs(2173));
    outputs(8466) <= layer0_outputs(8504);
    outputs(8467) <= (layer0_outputs(8335)) and (layer0_outputs(10129));
    outputs(8468) <= not((layer0_outputs(1533)) and (layer0_outputs(10998)));
    outputs(8469) <= not(layer0_outputs(7740));
    outputs(8470) <= not(layer0_outputs(11239));
    outputs(8471) <= not(layer0_outputs(9735));
    outputs(8472) <= layer0_outputs(1537);
    outputs(8473) <= layer0_outputs(6157);
    outputs(8474) <= (layer0_outputs(9791)) and not (layer0_outputs(5123));
    outputs(8475) <= (layer0_outputs(523)) xor (layer0_outputs(4293));
    outputs(8476) <= not((layer0_outputs(10366)) or (layer0_outputs(6667)));
    outputs(8477) <= not((layer0_outputs(5598)) xor (layer0_outputs(9091)));
    outputs(8478) <= not(layer0_outputs(916));
    outputs(8479) <= layer0_outputs(8156);
    outputs(8480) <= (layer0_outputs(7106)) and not (layer0_outputs(11004));
    outputs(8481) <= layer0_outputs(12336);
    outputs(8482) <= not((layer0_outputs(4022)) or (layer0_outputs(12290)));
    outputs(8483) <= not(layer0_outputs(8767));
    outputs(8484) <= (layer0_outputs(1073)) xor (layer0_outputs(6779));
    outputs(8485) <= not((layer0_outputs(2137)) xor (layer0_outputs(8338)));
    outputs(8486) <= not(layer0_outputs(540));
    outputs(8487) <= (layer0_outputs(7665)) xor (layer0_outputs(9912));
    outputs(8488) <= not((layer0_outputs(5659)) xor (layer0_outputs(3137)));
    outputs(8489) <= (layer0_outputs(10458)) and not (layer0_outputs(556));
    outputs(8490) <= (layer0_outputs(6007)) xor (layer0_outputs(618));
    outputs(8491) <= not(layer0_outputs(1362));
    outputs(8492) <= layer0_outputs(7290);
    outputs(8493) <= not((layer0_outputs(9906)) xor (layer0_outputs(6492)));
    outputs(8494) <= not((layer0_outputs(5869)) or (layer0_outputs(2842)));
    outputs(8495) <= not(layer0_outputs(10067));
    outputs(8496) <= not(layer0_outputs(5166)) or (layer0_outputs(10829));
    outputs(8497) <= layer0_outputs(3880);
    outputs(8498) <= layer0_outputs(7442);
    outputs(8499) <= (layer0_outputs(8132)) and (layer0_outputs(10861));
    outputs(8500) <= '0';
    outputs(8501) <= not(layer0_outputs(6577));
    outputs(8502) <= not((layer0_outputs(11172)) xor (layer0_outputs(8821)));
    outputs(8503) <= not((layer0_outputs(5307)) xor (layer0_outputs(10913)));
    outputs(8504) <= not((layer0_outputs(7593)) and (layer0_outputs(2316)));
    outputs(8505) <= (layer0_outputs(3064)) xor (layer0_outputs(8241));
    outputs(8506) <= layer0_outputs(5720);
    outputs(8507) <= (layer0_outputs(566)) and not (layer0_outputs(2574));
    outputs(8508) <= not(layer0_outputs(7181));
    outputs(8509) <= not(layer0_outputs(12403));
    outputs(8510) <= (layer0_outputs(10357)) xor (layer0_outputs(4451));
    outputs(8511) <= layer0_outputs(3755);
    outputs(8512) <= layer0_outputs(76);
    outputs(8513) <= layer0_outputs(9604);
    outputs(8514) <= (layer0_outputs(3281)) and (layer0_outputs(329));
    outputs(8515) <= not(layer0_outputs(8897));
    outputs(8516) <= layer0_outputs(1965);
    outputs(8517) <= (layer0_outputs(3021)) and not (layer0_outputs(1859));
    outputs(8518) <= not(layer0_outputs(1228)) or (layer0_outputs(12073));
    outputs(8519) <= not((layer0_outputs(12606)) xor (layer0_outputs(9463)));
    outputs(8520) <= not(layer0_outputs(11306));
    outputs(8521) <= not(layer0_outputs(11289)) or (layer0_outputs(9036));
    outputs(8522) <= (layer0_outputs(9430)) or (layer0_outputs(3414));
    outputs(8523) <= layer0_outputs(2752);
    outputs(8524) <= not(layer0_outputs(3064));
    outputs(8525) <= layer0_outputs(12192);
    outputs(8526) <= not((layer0_outputs(4432)) or (layer0_outputs(10210)));
    outputs(8527) <= (layer0_outputs(10269)) xor (layer0_outputs(9436));
    outputs(8528) <= not((layer0_outputs(10524)) xor (layer0_outputs(1806)));
    outputs(8529) <= not((layer0_outputs(4188)) xor (layer0_outputs(3838)));
    outputs(8530) <= (layer0_outputs(8792)) xor (layer0_outputs(12051));
    outputs(8531) <= not((layer0_outputs(4609)) xor (layer0_outputs(328)));
    outputs(8532) <= layer0_outputs(2274);
    outputs(8533) <= not((layer0_outputs(9080)) xor (layer0_outputs(7005)));
    outputs(8534) <= not((layer0_outputs(6561)) xor (layer0_outputs(5187)));
    outputs(8535) <= not(layer0_outputs(888));
    outputs(8536) <= not(layer0_outputs(12253));
    outputs(8537) <= not(layer0_outputs(327));
    outputs(8538) <= '1';
    outputs(8539) <= not(layer0_outputs(2988)) or (layer0_outputs(11034));
    outputs(8540) <= not(layer0_outputs(525));
    outputs(8541) <= layer0_outputs(2745);
    outputs(8542) <= layer0_outputs(1977);
    outputs(8543) <= layer0_outputs(10942);
    outputs(8544) <= not(layer0_outputs(7502));
    outputs(8545) <= not(layer0_outputs(2962)) or (layer0_outputs(6945));
    outputs(8546) <= (layer0_outputs(980)) and not (layer0_outputs(1356));
    outputs(8547) <= (layer0_outputs(3068)) xor (layer0_outputs(9555));
    outputs(8548) <= not(layer0_outputs(4946));
    outputs(8549) <= layer0_outputs(5534);
    outputs(8550) <= layer0_outputs(4773);
    outputs(8551) <= (layer0_outputs(7009)) or (layer0_outputs(10035));
    outputs(8552) <= not((layer0_outputs(12298)) or (layer0_outputs(5342)));
    outputs(8553) <= not((layer0_outputs(9493)) or (layer0_outputs(598)));
    outputs(8554) <= (layer0_outputs(12723)) xor (layer0_outputs(5562));
    outputs(8555) <= (layer0_outputs(10728)) xor (layer0_outputs(3530));
    outputs(8556) <= not(layer0_outputs(6043));
    outputs(8557) <= not(layer0_outputs(6339));
    outputs(8558) <= layer0_outputs(10198);
    outputs(8559) <= not(layer0_outputs(2494));
    outputs(8560) <= not(layer0_outputs(1529));
    outputs(8561) <= layer0_outputs(8450);
    outputs(8562) <= not((layer0_outputs(6460)) xor (layer0_outputs(10268)));
    outputs(8563) <= not((layer0_outputs(11609)) xor (layer0_outputs(9836)));
    outputs(8564) <= (layer0_outputs(8082)) xor (layer0_outputs(3047));
    outputs(8565) <= (layer0_outputs(6344)) xor (layer0_outputs(2074));
    outputs(8566) <= not((layer0_outputs(649)) or (layer0_outputs(5983)));
    outputs(8567) <= not(layer0_outputs(6434));
    outputs(8568) <= layer0_outputs(1682);
    outputs(8569) <= not(layer0_outputs(5565)) or (layer0_outputs(8342));
    outputs(8570) <= not((layer0_outputs(10072)) xor (layer0_outputs(10354)));
    outputs(8571) <= (layer0_outputs(4807)) xor (layer0_outputs(10138));
    outputs(8572) <= not((layer0_outputs(11743)) or (layer0_outputs(6164)));
    outputs(8573) <= (layer0_outputs(395)) or (layer0_outputs(11771));
    outputs(8574) <= not((layer0_outputs(12454)) and (layer0_outputs(10218)));
    outputs(8575) <= layer0_outputs(790);
    outputs(8576) <= not((layer0_outputs(7581)) and (layer0_outputs(6706)));
    outputs(8577) <= (layer0_outputs(7915)) xor (layer0_outputs(7731));
    outputs(8578) <= not(layer0_outputs(6626)) or (layer0_outputs(9041));
    outputs(8579) <= not(layer0_outputs(11319));
    outputs(8580) <= (layer0_outputs(2912)) and not (layer0_outputs(2208));
    outputs(8581) <= not(layer0_outputs(4085));
    outputs(8582) <= not((layer0_outputs(2063)) xor (layer0_outputs(9108)));
    outputs(8583) <= not((layer0_outputs(9933)) or (layer0_outputs(7426)));
    outputs(8584) <= not(layer0_outputs(5350));
    outputs(8585) <= not(layer0_outputs(9054));
    outputs(8586) <= (layer0_outputs(10804)) or (layer0_outputs(10800));
    outputs(8587) <= layer0_outputs(11279);
    outputs(8588) <= not((layer0_outputs(6116)) xor (layer0_outputs(1417)));
    outputs(8589) <= layer0_outputs(2587);
    outputs(8590) <= not((layer0_outputs(11259)) xor (layer0_outputs(12329)));
    outputs(8591) <= layer0_outputs(4392);
    outputs(8592) <= (layer0_outputs(349)) and not (layer0_outputs(3539));
    outputs(8593) <= (layer0_outputs(11956)) and not (layer0_outputs(7208));
    outputs(8594) <= not((layer0_outputs(7735)) xor (layer0_outputs(9950)));
    outputs(8595) <= not(layer0_outputs(1282));
    outputs(8596) <= not(layer0_outputs(1646));
    outputs(8597) <= not(layer0_outputs(2825));
    outputs(8598) <= (layer0_outputs(7462)) and not (layer0_outputs(6183));
    outputs(8599) <= (layer0_outputs(11797)) xor (layer0_outputs(8971));
    outputs(8600) <= (layer0_outputs(1458)) or (layer0_outputs(9842));
    outputs(8601) <= layer0_outputs(1294);
    outputs(8602) <= not((layer0_outputs(12677)) or (layer0_outputs(5463)));
    outputs(8603) <= not((layer0_outputs(5043)) xor (layer0_outputs(7166)));
    outputs(8604) <= not((layer0_outputs(8477)) xor (layer0_outputs(251)));
    outputs(8605) <= layer0_outputs(12599);
    outputs(8606) <= not(layer0_outputs(10375));
    outputs(8607) <= (layer0_outputs(10597)) and not (layer0_outputs(7066));
    outputs(8608) <= not(layer0_outputs(11884));
    outputs(8609) <= (layer0_outputs(9449)) and not (layer0_outputs(246));
    outputs(8610) <= not((layer0_outputs(4789)) or (layer0_outputs(4760)));
    outputs(8611) <= not((layer0_outputs(11025)) or (layer0_outputs(9986)));
    outputs(8612) <= (layer0_outputs(462)) xor (layer0_outputs(501));
    outputs(8613) <= layer0_outputs(2597);
    outputs(8614) <= not((layer0_outputs(8789)) and (layer0_outputs(12158)));
    outputs(8615) <= (layer0_outputs(219)) and not (layer0_outputs(1582));
    outputs(8616) <= not((layer0_outputs(5217)) xor (layer0_outputs(9339)));
    outputs(8617) <= (layer0_outputs(9215)) and (layer0_outputs(5594));
    outputs(8618) <= not(layer0_outputs(4886));
    outputs(8619) <= layer0_outputs(339);
    outputs(8620) <= not(layer0_outputs(8578));
    outputs(8621) <= not((layer0_outputs(8115)) and (layer0_outputs(11820)));
    outputs(8622) <= (layer0_outputs(6826)) and not (layer0_outputs(2614));
    outputs(8623) <= layer0_outputs(918);
    outputs(8624) <= layer0_outputs(12240);
    outputs(8625) <= not(layer0_outputs(1882));
    outputs(8626) <= (layer0_outputs(3693)) and (layer0_outputs(11439));
    outputs(8627) <= layer0_outputs(2729);
    outputs(8628) <= layer0_outputs(216);
    outputs(8629) <= (layer0_outputs(3372)) or (layer0_outputs(5008));
    outputs(8630) <= (layer0_outputs(2536)) and not (layer0_outputs(8511));
    outputs(8631) <= '1';
    outputs(8632) <= not(layer0_outputs(3093));
    outputs(8633) <= (layer0_outputs(4491)) xor (layer0_outputs(9598));
    outputs(8634) <= layer0_outputs(2088);
    outputs(8635) <= not((layer0_outputs(3409)) xor (layer0_outputs(8909)));
    outputs(8636) <= layer0_outputs(9069);
    outputs(8637) <= not(layer0_outputs(12285));
    outputs(8638) <= not((layer0_outputs(340)) xor (layer0_outputs(7649)));
    outputs(8639) <= not((layer0_outputs(12680)) or (layer0_outputs(2455)));
    outputs(8640) <= not(layer0_outputs(5495));
    outputs(8641) <= not(layer0_outputs(5414));
    outputs(8642) <= not(layer0_outputs(9585));
    outputs(8643) <= not((layer0_outputs(6342)) xor (layer0_outputs(766)));
    outputs(8644) <= (layer0_outputs(1290)) and not (layer0_outputs(7075));
    outputs(8645) <= (layer0_outputs(1137)) and (layer0_outputs(10220));
    outputs(8646) <= (layer0_outputs(10423)) xor (layer0_outputs(5924));
    outputs(8647) <= layer0_outputs(12160);
    outputs(8648) <= not((layer0_outputs(4740)) xor (layer0_outputs(11504)));
    outputs(8649) <= layer0_outputs(801);
    outputs(8650) <= not((layer0_outputs(3972)) xor (layer0_outputs(3142)));
    outputs(8651) <= not((layer0_outputs(4801)) and (layer0_outputs(3971)));
    outputs(8652) <= not((layer0_outputs(1355)) xor (layer0_outputs(6298)));
    outputs(8653) <= '0';
    outputs(8654) <= not(layer0_outputs(1866));
    outputs(8655) <= layer0_outputs(6447);
    outputs(8656) <= (layer0_outputs(589)) and not (layer0_outputs(2663));
    outputs(8657) <= not(layer0_outputs(717));
    outputs(8658) <= (layer0_outputs(10145)) and not (layer0_outputs(5506));
    outputs(8659) <= layer0_outputs(3070);
    outputs(8660) <= not((layer0_outputs(7552)) xor (layer0_outputs(6871)));
    outputs(8661) <= (layer0_outputs(7629)) and (layer0_outputs(10414));
    outputs(8662) <= not(layer0_outputs(132)) or (layer0_outputs(4332));
    outputs(8663) <= layer0_outputs(2450);
    outputs(8664) <= not((layer0_outputs(1097)) xor (layer0_outputs(10897)));
    outputs(8665) <= not((layer0_outputs(1538)) and (layer0_outputs(10029)));
    outputs(8666) <= not(layer0_outputs(19));
    outputs(8667) <= layer0_outputs(2055);
    outputs(8668) <= not(layer0_outputs(10958));
    outputs(8669) <= '1';
    outputs(8670) <= not(layer0_outputs(9754)) or (layer0_outputs(11611));
    outputs(8671) <= not((layer0_outputs(11042)) xor (layer0_outputs(6915)));
    outputs(8672) <= not((layer0_outputs(2255)) xor (layer0_outputs(6906)));
    outputs(8673) <= (layer0_outputs(5248)) and not (layer0_outputs(6887));
    outputs(8674) <= (layer0_outputs(11665)) and not (layer0_outputs(7620));
    outputs(8675) <= '0';
    outputs(8676) <= (layer0_outputs(12056)) xor (layer0_outputs(10444));
    outputs(8677) <= (layer0_outputs(12688)) xor (layer0_outputs(5106));
    outputs(8678) <= not(layer0_outputs(3049));
    outputs(8679) <= (layer0_outputs(9841)) xor (layer0_outputs(12231));
    outputs(8680) <= layer0_outputs(3067);
    outputs(8681) <= layer0_outputs(8702);
    outputs(8682) <= not((layer0_outputs(12221)) xor (layer0_outputs(7968)));
    outputs(8683) <= not(layer0_outputs(4792));
    outputs(8684) <= (layer0_outputs(6840)) xor (layer0_outputs(10049));
    outputs(8685) <= not(layer0_outputs(5928));
    outputs(8686) <= (layer0_outputs(11580)) and not (layer0_outputs(3229));
    outputs(8687) <= not(layer0_outputs(8298));
    outputs(8688) <= not(layer0_outputs(3763));
    outputs(8689) <= not((layer0_outputs(7025)) or (layer0_outputs(3482)));
    outputs(8690) <= (layer0_outputs(1381)) or (layer0_outputs(9269));
    outputs(8691) <= not(layer0_outputs(1620));
    outputs(8692) <= (layer0_outputs(10501)) xor (layer0_outputs(10924));
    outputs(8693) <= (layer0_outputs(5476)) and (layer0_outputs(8987));
    outputs(8694) <= (layer0_outputs(3090)) xor (layer0_outputs(5080));
    outputs(8695) <= not(layer0_outputs(522)) or (layer0_outputs(12504));
    outputs(8696) <= not(layer0_outputs(9978));
    outputs(8697) <= not(layer0_outputs(5445));
    outputs(8698) <= layer0_outputs(349);
    outputs(8699) <= layer0_outputs(1577);
    outputs(8700) <= layer0_outputs(12344);
    outputs(8701) <= (layer0_outputs(4460)) and not (layer0_outputs(4808));
    outputs(8702) <= (layer0_outputs(5750)) xor (layer0_outputs(3106));
    outputs(8703) <= not(layer0_outputs(8758));
    outputs(8704) <= not((layer0_outputs(3128)) xor (layer0_outputs(12097)));
    outputs(8705) <= not((layer0_outputs(9299)) or (layer0_outputs(2790)));
    outputs(8706) <= layer0_outputs(9332);
    outputs(8707) <= layer0_outputs(10612);
    outputs(8708) <= not(layer0_outputs(9678));
    outputs(8709) <= layer0_outputs(3798);
    outputs(8710) <= (layer0_outputs(9759)) xor (layer0_outputs(1673));
    outputs(8711) <= not((layer0_outputs(1745)) xor (layer0_outputs(7959)));
    outputs(8712) <= not((layer0_outputs(12712)) xor (layer0_outputs(9829)));
    outputs(8713) <= layer0_outputs(3962);
    outputs(8714) <= layer0_outputs(8349);
    outputs(8715) <= layer0_outputs(5296);
    outputs(8716) <= not(layer0_outputs(9735));
    outputs(8717) <= not((layer0_outputs(5299)) xor (layer0_outputs(10150)));
    outputs(8718) <= not(layer0_outputs(5308));
    outputs(8719) <= not(layer0_outputs(3674));
    outputs(8720) <= (layer0_outputs(10900)) or (layer0_outputs(11385));
    outputs(8721) <= not(layer0_outputs(5901));
    outputs(8722) <= layer0_outputs(1441);
    outputs(8723) <= not((layer0_outputs(3408)) and (layer0_outputs(9865)));
    outputs(8724) <= not((layer0_outputs(11783)) and (layer0_outputs(10164)));
    outputs(8725) <= (layer0_outputs(5156)) or (layer0_outputs(7194));
    outputs(8726) <= not((layer0_outputs(10914)) xor (layer0_outputs(5596)));
    outputs(8727) <= layer0_outputs(1504);
    outputs(8728) <= layer0_outputs(1967);
    outputs(8729) <= not(layer0_outputs(8447));
    outputs(8730) <= (layer0_outputs(9056)) xor (layer0_outputs(9996));
    outputs(8731) <= (layer0_outputs(250)) or (layer0_outputs(782));
    outputs(8732) <= not(layer0_outputs(1326)) or (layer0_outputs(1867));
    outputs(8733) <= not(layer0_outputs(5796)) or (layer0_outputs(6520));
    outputs(8734) <= not((layer0_outputs(7839)) or (layer0_outputs(2236)));
    outputs(8735) <= (layer0_outputs(7146)) xor (layer0_outputs(10725));
    outputs(8736) <= layer0_outputs(9906);
    outputs(8737) <= not(layer0_outputs(12162));
    outputs(8738) <= (layer0_outputs(9227)) and not (layer0_outputs(11659));
    outputs(8739) <= (layer0_outputs(9194)) or (layer0_outputs(10350));
    outputs(8740) <= (layer0_outputs(56)) xor (layer0_outputs(4811));
    outputs(8741) <= layer0_outputs(5597);
    outputs(8742) <= layer0_outputs(1683);
    outputs(8743) <= (layer0_outputs(12752)) xor (layer0_outputs(7630));
    outputs(8744) <= layer0_outputs(5840);
    outputs(8745) <= not((layer0_outputs(11169)) xor (layer0_outputs(1911)));
    outputs(8746) <= not(layer0_outputs(9130)) or (layer0_outputs(9588));
    outputs(8747) <= not(layer0_outputs(1224));
    outputs(8748) <= layer0_outputs(6769);
    outputs(8749) <= layer0_outputs(11672);
    outputs(8750) <= (layer0_outputs(5993)) and not (layer0_outputs(493));
    outputs(8751) <= layer0_outputs(10128);
    outputs(8752) <= not((layer0_outputs(10093)) and (layer0_outputs(9954)));
    outputs(8753) <= not(layer0_outputs(284));
    outputs(8754) <= (layer0_outputs(393)) xor (layer0_outputs(6013));
    outputs(8755) <= not(layer0_outputs(3356));
    outputs(8756) <= not(layer0_outputs(9965));
    outputs(8757) <= layer0_outputs(9974);
    outputs(8758) <= not(layer0_outputs(10563));
    outputs(8759) <= not(layer0_outputs(9311));
    outputs(8760) <= layer0_outputs(3831);
    outputs(8761) <= not(layer0_outputs(4182));
    outputs(8762) <= (layer0_outputs(8169)) and (layer0_outputs(2958));
    outputs(8763) <= not(layer0_outputs(388)) or (layer0_outputs(6405));
    outputs(8764) <= not(layer0_outputs(11317));
    outputs(8765) <= not(layer0_outputs(11573));
    outputs(8766) <= layer0_outputs(1274);
    outputs(8767) <= layer0_outputs(11049);
    outputs(8768) <= not(layer0_outputs(1463));
    outputs(8769) <= layer0_outputs(7760);
    outputs(8770) <= not(layer0_outputs(8108)) or (layer0_outputs(10056));
    outputs(8771) <= not(layer0_outputs(6546));
    outputs(8772) <= not(layer0_outputs(3529)) or (layer0_outputs(780));
    outputs(8773) <= (layer0_outputs(8256)) or (layer0_outputs(4683));
    outputs(8774) <= (layer0_outputs(11975)) xor (layer0_outputs(9706));
    outputs(8775) <= not(layer0_outputs(8162));
    outputs(8776) <= not((layer0_outputs(11714)) xor (layer0_outputs(1382)));
    outputs(8777) <= not((layer0_outputs(7871)) xor (layer0_outputs(12628)));
    outputs(8778) <= layer0_outputs(6231);
    outputs(8779) <= (layer0_outputs(12333)) xor (layer0_outputs(9914));
    outputs(8780) <= not(layer0_outputs(5442));
    outputs(8781) <= not(layer0_outputs(7121));
    outputs(8782) <= layer0_outputs(7059);
    outputs(8783) <= layer0_outputs(11471);
    outputs(8784) <= (layer0_outputs(12277)) or (layer0_outputs(7331));
    outputs(8785) <= not(layer0_outputs(11982));
    outputs(8786) <= layer0_outputs(3587);
    outputs(8787) <= not((layer0_outputs(3334)) and (layer0_outputs(5673)));
    outputs(8788) <= layer0_outputs(4983);
    outputs(8789) <= not(layer0_outputs(885));
    outputs(8790) <= not((layer0_outputs(8369)) xor (layer0_outputs(6684)));
    outputs(8791) <= not(layer0_outputs(10532));
    outputs(8792) <= (layer0_outputs(385)) and not (layer0_outputs(6184));
    outputs(8793) <= not((layer0_outputs(5898)) xor (layer0_outputs(11468)));
    outputs(8794) <= not((layer0_outputs(2010)) xor (layer0_outputs(4542)));
    outputs(8795) <= (layer0_outputs(7095)) or (layer0_outputs(3443));
    outputs(8796) <= (layer0_outputs(3987)) xor (layer0_outputs(3465));
    outputs(8797) <= not(layer0_outputs(9116));
    outputs(8798) <= not((layer0_outputs(186)) xor (layer0_outputs(11710)));
    outputs(8799) <= (layer0_outputs(5655)) and not (layer0_outputs(1953));
    outputs(8800) <= (layer0_outputs(1561)) and not (layer0_outputs(2747));
    outputs(8801) <= not(layer0_outputs(6053));
    outputs(8802) <= not(layer0_outputs(4434)) or (layer0_outputs(6963));
    outputs(8803) <= layer0_outputs(8198);
    outputs(8804) <= not((layer0_outputs(10250)) xor (layer0_outputs(9563)));
    outputs(8805) <= layer0_outputs(3375);
    outputs(8806) <= layer0_outputs(9463);
    outputs(8807) <= (layer0_outputs(8311)) or (layer0_outputs(10698));
    outputs(8808) <= layer0_outputs(3527);
    outputs(8809) <= (layer0_outputs(2499)) xor (layer0_outputs(834));
    outputs(8810) <= not(layer0_outputs(7991));
    outputs(8811) <= not((layer0_outputs(473)) xor (layer0_outputs(1181)));
    outputs(8812) <= not(layer0_outputs(8893));
    outputs(8813) <= not((layer0_outputs(11096)) xor (layer0_outputs(4888)));
    outputs(8814) <= layer0_outputs(3875);
    outputs(8815) <= not(layer0_outputs(11235));
    outputs(8816) <= not((layer0_outputs(1546)) xor (layer0_outputs(10766)));
    outputs(8817) <= (layer0_outputs(6953)) xor (layer0_outputs(4306));
    outputs(8818) <= layer0_outputs(1160);
    outputs(8819) <= not(layer0_outputs(12644));
    outputs(8820) <= layer0_outputs(496);
    outputs(8821) <= not(layer0_outputs(10841));
    outputs(8822) <= not((layer0_outputs(11780)) xor (layer0_outputs(8259)));
    outputs(8823) <= (layer0_outputs(9484)) and not (layer0_outputs(4732));
    outputs(8824) <= (layer0_outputs(9271)) or (layer0_outputs(11705));
    outputs(8825) <= not(layer0_outputs(3125)) or (layer0_outputs(3575));
    outputs(8826) <= not((layer0_outputs(3428)) xor (layer0_outputs(6340)));
    outputs(8827) <= (layer0_outputs(10449)) xor (layer0_outputs(10671));
    outputs(8828) <= (layer0_outputs(6815)) xor (layer0_outputs(4095));
    outputs(8829) <= (layer0_outputs(9456)) and not (layer0_outputs(1814));
    outputs(8830) <= layer0_outputs(6909);
    outputs(8831) <= not(layer0_outputs(248));
    outputs(8832) <= not(layer0_outputs(855));
    outputs(8833) <= not((layer0_outputs(268)) xor (layer0_outputs(3413)));
    outputs(8834) <= layer0_outputs(4154);
    outputs(8835) <= not((layer0_outputs(1932)) xor (layer0_outputs(4053)));
    outputs(8836) <= (layer0_outputs(12683)) xor (layer0_outputs(5722));
    outputs(8837) <= not((layer0_outputs(1962)) or (layer0_outputs(2476)));
    outputs(8838) <= not((layer0_outputs(6303)) xor (layer0_outputs(7411)));
    outputs(8839) <= layer0_outputs(12327);
    outputs(8840) <= not(layer0_outputs(5237));
    outputs(8841) <= layer0_outputs(3524);
    outputs(8842) <= not(layer0_outputs(2030));
    outputs(8843) <= layer0_outputs(9275);
    outputs(8844) <= not(layer0_outputs(7538)) or (layer0_outputs(9233));
    outputs(8845) <= not(layer0_outputs(4653));
    outputs(8846) <= not(layer0_outputs(1012));
    outputs(8847) <= not((layer0_outputs(10980)) xor (layer0_outputs(6653)));
    outputs(8848) <= (layer0_outputs(12553)) and (layer0_outputs(12114));
    outputs(8849) <= not((layer0_outputs(183)) xor (layer0_outputs(9177)));
    outputs(8850) <= (layer0_outputs(10858)) xor (layer0_outputs(2521));
    outputs(8851) <= not(layer0_outputs(11618));
    outputs(8852) <= not((layer0_outputs(8850)) xor (layer0_outputs(4417)));
    outputs(8853) <= not((layer0_outputs(3566)) xor (layer0_outputs(3826)));
    outputs(8854) <= not(layer0_outputs(3022));
    outputs(8855) <= layer0_outputs(6631);
    outputs(8856) <= (layer0_outputs(3168)) or (layer0_outputs(5554));
    outputs(8857) <= layer0_outputs(5708);
    outputs(8858) <= layer0_outputs(2445);
    outputs(8859) <= not((layer0_outputs(6318)) xor (layer0_outputs(11215)));
    outputs(8860) <= (layer0_outputs(585)) xor (layer0_outputs(6188));
    outputs(8861) <= (layer0_outputs(5033)) and not (layer0_outputs(8251));
    outputs(8862) <= (layer0_outputs(9654)) and not (layer0_outputs(9763));
    outputs(8863) <= not(layer0_outputs(4893));
    outputs(8864) <= (layer0_outputs(12620)) and not (layer0_outputs(1870));
    outputs(8865) <= not((layer0_outputs(12798)) xor (layer0_outputs(11899)));
    outputs(8866) <= (layer0_outputs(2195)) or (layer0_outputs(1616));
    outputs(8867) <= (layer0_outputs(6090)) and not (layer0_outputs(9162));
    outputs(8868) <= not(layer0_outputs(6990));
    outputs(8869) <= layer0_outputs(9214);
    outputs(8870) <= not(layer0_outputs(4300));
    outputs(8871) <= (layer0_outputs(7004)) xor (layer0_outputs(4738));
    outputs(8872) <= not(layer0_outputs(7702));
    outputs(8873) <= (layer0_outputs(1898)) or (layer0_outputs(10491));
    outputs(8874) <= layer0_outputs(7627);
    outputs(8875) <= layer0_outputs(8213);
    outputs(8876) <= (layer0_outputs(6212)) xor (layer0_outputs(7071));
    outputs(8877) <= (layer0_outputs(6140)) xor (layer0_outputs(7138));
    outputs(8878) <= not(layer0_outputs(3207)) or (layer0_outputs(7205));
    outputs(8879) <= not(layer0_outputs(11638));
    outputs(8880) <= not(layer0_outputs(7427)) or (layer0_outputs(9173));
    outputs(8881) <= not((layer0_outputs(131)) xor (layer0_outputs(9231)));
    outputs(8882) <= layer0_outputs(11334);
    outputs(8883) <= '0';
    outputs(8884) <= (layer0_outputs(9519)) and (layer0_outputs(8485));
    outputs(8885) <= (layer0_outputs(4813)) xor (layer0_outputs(7));
    outputs(8886) <= (layer0_outputs(10910)) xor (layer0_outputs(10451));
    outputs(8887) <= layer0_outputs(9466);
    outputs(8888) <= layer0_outputs(10536);
    outputs(8889) <= (layer0_outputs(2792)) and not (layer0_outputs(1418));
    outputs(8890) <= not(layer0_outputs(2096));
    outputs(8891) <= not(layer0_outputs(1585));
    outputs(8892) <= (layer0_outputs(8858)) or (layer0_outputs(9807));
    outputs(8893) <= not(layer0_outputs(354));
    outputs(8894) <= layer0_outputs(6191);
    outputs(8895) <= layer0_outputs(650);
    outputs(8896) <= not(layer0_outputs(10248)) or (layer0_outputs(1575));
    outputs(8897) <= not(layer0_outputs(9987));
    outputs(8898) <= layer0_outputs(9298);
    outputs(8899) <= layer0_outputs(1098);
    outputs(8900) <= (layer0_outputs(8244)) and not (layer0_outputs(8837));
    outputs(8901) <= (layer0_outputs(3269)) xor (layer0_outputs(3740));
    outputs(8902) <= not(layer0_outputs(11242)) or (layer0_outputs(6757));
    outputs(8903) <= layer0_outputs(790);
    outputs(8904) <= layer0_outputs(10834);
    outputs(8905) <= not((layer0_outputs(8260)) or (layer0_outputs(12569)));
    outputs(8906) <= not(layer0_outputs(4405)) or (layer0_outputs(11704));
    outputs(8907) <= (layer0_outputs(1341)) and not (layer0_outputs(4601));
    outputs(8908) <= layer0_outputs(9097);
    outputs(8909) <= not(layer0_outputs(3802));
    outputs(8910) <= layer0_outputs(12286);
    outputs(8911) <= not((layer0_outputs(518)) xor (layer0_outputs(7105)));
    outputs(8912) <= not(layer0_outputs(8167));
    outputs(8913) <= layer0_outputs(3624);
    outputs(8914) <= layer0_outputs(1213);
    outputs(8915) <= (layer0_outputs(7430)) and not (layer0_outputs(11684));
    outputs(8916) <= layer0_outputs(9830);
    outputs(8917) <= not(layer0_outputs(6672)) or (layer0_outputs(9271));
    outputs(8918) <= (layer0_outputs(2186)) xor (layer0_outputs(3112));
    outputs(8919) <= layer0_outputs(738);
    outputs(8920) <= not(layer0_outputs(8060));
    outputs(8921) <= not(layer0_outputs(9987));
    outputs(8922) <= not((layer0_outputs(11839)) or (layer0_outputs(2701)));
    outputs(8923) <= not(layer0_outputs(9223));
    outputs(8924) <= (layer0_outputs(5757)) xor (layer0_outputs(12771));
    outputs(8925) <= (layer0_outputs(7477)) or (layer0_outputs(1548));
    outputs(8926) <= not(layer0_outputs(6453));
    outputs(8927) <= not(layer0_outputs(1486)) or (layer0_outputs(12345));
    outputs(8928) <= (layer0_outputs(6262)) xor (layer0_outputs(9307));
    outputs(8929) <= (layer0_outputs(6564)) xor (layer0_outputs(9887));
    outputs(8930) <= not((layer0_outputs(7395)) and (layer0_outputs(11306)));
    outputs(8931) <= not((layer0_outputs(2246)) and (layer0_outputs(6536)));
    outputs(8932) <= not(layer0_outputs(10676));
    outputs(8933) <= (layer0_outputs(2446)) and not (layer0_outputs(11021));
    outputs(8934) <= layer0_outputs(187);
    outputs(8935) <= not(layer0_outputs(1477));
    outputs(8936) <= not((layer0_outputs(9269)) xor (layer0_outputs(7927)));
    outputs(8937) <= not(layer0_outputs(6999));
    outputs(8938) <= not(layer0_outputs(4642)) or (layer0_outputs(3982));
    outputs(8939) <= not(layer0_outputs(10738)) or (layer0_outputs(5171));
    outputs(8940) <= (layer0_outputs(9739)) xor (layer0_outputs(10063));
    outputs(8941) <= layer0_outputs(11652);
    outputs(8942) <= (layer0_outputs(7866)) xor (layer0_outputs(1045));
    outputs(8943) <= (layer0_outputs(8326)) and (layer0_outputs(2328));
    outputs(8944) <= not(layer0_outputs(2609));
    outputs(8945) <= not((layer0_outputs(8884)) xor (layer0_outputs(8128)));
    outputs(8946) <= layer0_outputs(7081);
    outputs(8947) <= layer0_outputs(2373);
    outputs(8948) <= (layer0_outputs(9896)) xor (layer0_outputs(625));
    outputs(8949) <= (layer0_outputs(10172)) xor (layer0_outputs(12702));
    outputs(8950) <= not((layer0_outputs(9797)) xor (layer0_outputs(11389)));
    outputs(8951) <= (layer0_outputs(1214)) xor (layer0_outputs(3403));
    outputs(8952) <= not(layer0_outputs(10707)) or (layer0_outputs(8862));
    outputs(8953) <= (layer0_outputs(4259)) xor (layer0_outputs(37));
    outputs(8954) <= layer0_outputs(3078);
    outputs(8955) <= not(layer0_outputs(956));
    outputs(8956) <= not(layer0_outputs(9247));
    outputs(8957) <= (layer0_outputs(7672)) or (layer0_outputs(12514));
    outputs(8958) <= not((layer0_outputs(6981)) and (layer0_outputs(11056)));
    outputs(8959) <= layer0_outputs(500);
    outputs(8960) <= not(layer0_outputs(4551));
    outputs(8961) <= not(layer0_outputs(10840));
    outputs(8962) <= (layer0_outputs(3764)) and not (layer0_outputs(9661));
    outputs(8963) <= (layer0_outputs(8492)) and (layer0_outputs(212));
    outputs(8964) <= (layer0_outputs(11336)) and not (layer0_outputs(8171));
    outputs(8965) <= not(layer0_outputs(2868));
    outputs(8966) <= layer0_outputs(9032);
    outputs(8967) <= (layer0_outputs(9180)) and (layer0_outputs(2800));
    outputs(8968) <= (layer0_outputs(4190)) xor (layer0_outputs(7670));
    outputs(8969) <= (layer0_outputs(4246)) or (layer0_outputs(6229));
    outputs(8970) <= not(layer0_outputs(8322)) or (layer0_outputs(1186));
    outputs(8971) <= (layer0_outputs(921)) xor (layer0_outputs(9634));
    outputs(8972) <= not((layer0_outputs(7360)) xor (layer0_outputs(12505)));
    outputs(8973) <= not(layer0_outputs(5184));
    outputs(8974) <= not((layer0_outputs(11861)) or (layer0_outputs(4425)));
    outputs(8975) <= layer0_outputs(8406);
    outputs(8976) <= layer0_outputs(5736);
    outputs(8977) <= not((layer0_outputs(1708)) xor (layer0_outputs(9958)));
    outputs(8978) <= (layer0_outputs(4123)) or (layer0_outputs(4276));
    outputs(8979) <= (layer0_outputs(9737)) and (layer0_outputs(6245));
    outputs(8980) <= not((layer0_outputs(10574)) or (layer0_outputs(8703)));
    outputs(8981) <= not((layer0_outputs(4102)) xor (layer0_outputs(2343)));
    outputs(8982) <= not((layer0_outputs(1727)) xor (layer0_outputs(325)));
    outputs(8983) <= not((layer0_outputs(955)) or (layer0_outputs(4016)));
    outputs(8984) <= not(layer0_outputs(6957)) or (layer0_outputs(6555));
    outputs(8985) <= not((layer0_outputs(10804)) xor (layer0_outputs(3719)));
    outputs(8986) <= layer0_outputs(7870);
    outputs(8987) <= not(layer0_outputs(3062)) or (layer0_outputs(11534));
    outputs(8988) <= layer0_outputs(8006);
    outputs(8989) <= layer0_outputs(8505);
    outputs(8990) <= not(layer0_outputs(1530));
    outputs(8991) <= not(layer0_outputs(2147));
    outputs(8992) <= not((layer0_outputs(2503)) xor (layer0_outputs(10047)));
    outputs(8993) <= (layer0_outputs(5535)) xor (layer0_outputs(12280));
    outputs(8994) <= not(layer0_outputs(6887));
    outputs(8995) <= layer0_outputs(2859);
    outputs(8996) <= not((layer0_outputs(3593)) or (layer0_outputs(10979)));
    outputs(8997) <= not(layer0_outputs(11942));
    outputs(8998) <= layer0_outputs(3083);
    outputs(8999) <= layer0_outputs(10274);
    outputs(9000) <= layer0_outputs(104);
    outputs(9001) <= not(layer0_outputs(5428));
    outputs(9002) <= (layer0_outputs(2914)) xor (layer0_outputs(7368));
    outputs(9003) <= layer0_outputs(1840);
    outputs(9004) <= layer0_outputs(7800);
    outputs(9005) <= not(layer0_outputs(646)) or (layer0_outputs(12187));
    outputs(9006) <= not((layer0_outputs(10118)) xor (layer0_outputs(12625)));
    outputs(9007) <= '0';
    outputs(9008) <= not(layer0_outputs(5205));
    outputs(9009) <= layer0_outputs(6900);
    outputs(9010) <= not(layer0_outputs(2493));
    outputs(9011) <= (layer0_outputs(8360)) xor (layer0_outputs(10222));
    outputs(9012) <= not(layer0_outputs(11721));
    outputs(9013) <= (layer0_outputs(7771)) xor (layer0_outputs(5628));
    outputs(9014) <= layer0_outputs(8654);
    outputs(9015) <= not(layer0_outputs(956));
    outputs(9016) <= not((layer0_outputs(4350)) xor (layer0_outputs(8417)));
    outputs(9017) <= (layer0_outputs(5005)) and (layer0_outputs(11960));
    outputs(9018) <= not(layer0_outputs(4049));
    outputs(9019) <= not((layer0_outputs(4286)) xor (layer0_outputs(5442)));
    outputs(9020) <= not((layer0_outputs(2959)) xor (layer0_outputs(12767)));
    outputs(9021) <= (layer0_outputs(4177)) and not (layer0_outputs(5191));
    outputs(9022) <= not(layer0_outputs(4864)) or (layer0_outputs(7216));
    outputs(9023) <= (layer0_outputs(12519)) and not (layer0_outputs(7985));
    outputs(9024) <= layer0_outputs(6690);
    outputs(9025) <= (layer0_outputs(4931)) xor (layer0_outputs(5499));
    outputs(9026) <= layer0_outputs(12322);
    outputs(9027) <= not(layer0_outputs(8630));
    outputs(9028) <= not((layer0_outputs(6369)) xor (layer0_outputs(7138)));
    outputs(9029) <= not((layer0_outputs(12013)) xor (layer0_outputs(5458)));
    outputs(9030) <= not(layer0_outputs(11686));
    outputs(9031) <= layer0_outputs(10312);
    outputs(9032) <= (layer0_outputs(6232)) and not (layer0_outputs(2228));
    outputs(9033) <= not((layer0_outputs(8042)) xor (layer0_outputs(3281)));
    outputs(9034) <= (layer0_outputs(6594)) and (layer0_outputs(3565));
    outputs(9035) <= (layer0_outputs(5158)) and not (layer0_outputs(8207));
    outputs(9036) <= not(layer0_outputs(11838));
    outputs(9037) <= not((layer0_outputs(3745)) xor (layer0_outputs(11186)));
    outputs(9038) <= (layer0_outputs(10814)) and not (layer0_outputs(10741));
    outputs(9039) <= (layer0_outputs(6365)) and not (layer0_outputs(1468));
    outputs(9040) <= (layer0_outputs(7059)) and not (layer0_outputs(7667));
    outputs(9041) <= (layer0_outputs(698)) xor (layer0_outputs(4624));
    outputs(9042) <= (layer0_outputs(5382)) xor (layer0_outputs(2525));
    outputs(9043) <= (layer0_outputs(11516)) xor (layer0_outputs(11769));
    outputs(9044) <= layer0_outputs(9793);
    outputs(9045) <= layer0_outputs(11681);
    outputs(9046) <= not(layer0_outputs(788));
    outputs(9047) <= not((layer0_outputs(8543)) xor (layer0_outputs(6994)));
    outputs(9048) <= (layer0_outputs(4051)) xor (layer0_outputs(6633));
    outputs(9049) <= (layer0_outputs(8463)) and not (layer0_outputs(7658));
    outputs(9050) <= layer0_outputs(3174);
    outputs(9051) <= not((layer0_outputs(11970)) xor (layer0_outputs(10531)));
    outputs(9052) <= (layer0_outputs(9160)) and not (layer0_outputs(3650));
    outputs(9053) <= layer0_outputs(8404);
    outputs(9054) <= '0';
    outputs(9055) <= not((layer0_outputs(10706)) xor (layer0_outputs(2438)));
    outputs(9056) <= (layer0_outputs(10579)) and not (layer0_outputs(1974));
    outputs(9057) <= layer0_outputs(2939);
    outputs(9058) <= (layer0_outputs(1006)) and not (layer0_outputs(7909));
    outputs(9059) <= layer0_outputs(6778);
    outputs(9060) <= layer0_outputs(7541);
    outputs(9061) <= (layer0_outputs(3442)) and not (layer0_outputs(2722));
    outputs(9062) <= (layer0_outputs(138)) and not (layer0_outputs(5939));
    outputs(9063) <= (layer0_outputs(11408)) and (layer0_outputs(12775));
    outputs(9064) <= not(layer0_outputs(1896));
    outputs(9065) <= layer0_outputs(4520);
    outputs(9066) <= (layer0_outputs(5469)) and (layer0_outputs(9851));
    outputs(9067) <= (layer0_outputs(3318)) or (layer0_outputs(2743));
    outputs(9068) <= (layer0_outputs(5984)) and (layer0_outputs(3637));
    outputs(9069) <= not(layer0_outputs(11296));
    outputs(9070) <= layer0_outputs(4421);
    outputs(9071) <= not((layer0_outputs(11824)) and (layer0_outputs(3036)));
    outputs(9072) <= layer0_outputs(11527);
    outputs(9073) <= not((layer0_outputs(1963)) or (layer0_outputs(11690)));
    outputs(9074) <= not(layer0_outputs(11976));
    outputs(9075) <= not(layer0_outputs(9931));
    outputs(9076) <= (layer0_outputs(1502)) xor (layer0_outputs(10719));
    outputs(9077) <= not(layer0_outputs(6841));
    outputs(9078) <= layer0_outputs(6102);
    outputs(9079) <= (layer0_outputs(5228)) and not (layer0_outputs(10482));
    outputs(9080) <= not((layer0_outputs(8054)) or (layer0_outputs(8629)));
    outputs(9081) <= layer0_outputs(8321);
    outputs(9082) <= layer0_outputs(1429);
    outputs(9083) <= (layer0_outputs(1123)) or (layer0_outputs(7154));
    outputs(9084) <= layer0_outputs(11209);
    outputs(9085) <= not(layer0_outputs(6913));
    outputs(9086) <= not(layer0_outputs(9831));
    outputs(9087) <= (layer0_outputs(6080)) and not (layer0_outputs(12351));
    outputs(9088) <= not(layer0_outputs(1498));
    outputs(9089) <= not((layer0_outputs(4193)) xor (layer0_outputs(9935)));
    outputs(9090) <= layer0_outputs(8973);
    outputs(9091) <= not(layer0_outputs(10566));
    outputs(9092) <= (layer0_outputs(858)) xor (layer0_outputs(6635));
    outputs(9093) <= layer0_outputs(8314);
    outputs(9094) <= not(layer0_outputs(2628));
    outputs(9095) <= not((layer0_outputs(8738)) xor (layer0_outputs(2668)));
    outputs(9096) <= layer0_outputs(11577);
    outputs(9097) <= not(layer0_outputs(4998));
    outputs(9098) <= not((layer0_outputs(11144)) or (layer0_outputs(9945)));
    outputs(9099) <= not((layer0_outputs(6564)) xor (layer0_outputs(10548)));
    outputs(9100) <= not(layer0_outputs(5960));
    outputs(9101) <= not(layer0_outputs(639));
    outputs(9102) <= not((layer0_outputs(8691)) xor (layer0_outputs(3741)));
    outputs(9103) <= not(layer0_outputs(11162));
    outputs(9104) <= not((layer0_outputs(4920)) xor (layer0_outputs(8641)));
    outputs(9105) <= not((layer0_outputs(731)) xor (layer0_outputs(4399)));
    outputs(9106) <= layer0_outputs(2534);
    outputs(9107) <= not(layer0_outputs(8785));
    outputs(9108) <= (layer0_outputs(1490)) xor (layer0_outputs(4517));
    outputs(9109) <= layer0_outputs(17);
    outputs(9110) <= layer0_outputs(7638);
    outputs(9111) <= (layer0_outputs(3043)) and not (layer0_outputs(126));
    outputs(9112) <= not(layer0_outputs(5826)) or (layer0_outputs(2314));
    outputs(9113) <= not(layer0_outputs(7627));
    outputs(9114) <= '0';
    outputs(9115) <= layer0_outputs(3931);
    outputs(9116) <= not((layer0_outputs(3499)) or (layer0_outputs(4649)));
    outputs(9117) <= layer0_outputs(9383);
    outputs(9118) <= not(layer0_outputs(2283));
    outputs(9119) <= not((layer0_outputs(10208)) and (layer0_outputs(12714)));
    outputs(9120) <= not(layer0_outputs(7652)) or (layer0_outputs(9785));
    outputs(9121) <= (layer0_outputs(10164)) and not (layer0_outputs(6124));
    outputs(9122) <= layer0_outputs(6510);
    outputs(9123) <= layer0_outputs(4642);
    outputs(9124) <= layer0_outputs(4799);
    outputs(9125) <= (layer0_outputs(4100)) xor (layer0_outputs(1353));
    outputs(9126) <= layer0_outputs(7046);
    outputs(9127) <= not((layer0_outputs(11866)) and (layer0_outputs(7765)));
    outputs(9128) <= not(layer0_outputs(8808));
    outputs(9129) <= not(layer0_outputs(10909));
    outputs(9130) <= not(layer0_outputs(3903));
    outputs(9131) <= not((layer0_outputs(4924)) xor (layer0_outputs(5203)));
    outputs(9132) <= layer0_outputs(9459);
    outputs(9133) <= not((layer0_outputs(7179)) xor (layer0_outputs(5013)));
    outputs(9134) <= layer0_outputs(7467);
    outputs(9135) <= layer0_outputs(8273);
    outputs(9136) <= (layer0_outputs(3140)) xor (layer0_outputs(11287));
    outputs(9137) <= (layer0_outputs(11529)) xor (layer0_outputs(8919));
    outputs(9138) <= (layer0_outputs(4171)) and not (layer0_outputs(6535));
    outputs(9139) <= not(layer0_outputs(7787));
    outputs(9140) <= layer0_outputs(6134);
    outputs(9141) <= (layer0_outputs(5458)) xor (layer0_outputs(671));
    outputs(9142) <= layer0_outputs(11644);
    outputs(9143) <= layer0_outputs(4824);
    outputs(9144) <= not(layer0_outputs(3024));
    outputs(9145) <= not((layer0_outputs(9938)) and (layer0_outputs(3962)));
    outputs(9146) <= (layer0_outputs(12164)) and (layer0_outputs(4426));
    outputs(9147) <= layer0_outputs(11926);
    outputs(9148) <= layer0_outputs(5512);
    outputs(9149) <= layer0_outputs(3527);
    outputs(9150) <= layer0_outputs(8047);
    outputs(9151) <= '0';
    outputs(9152) <= not((layer0_outputs(1415)) xor (layer0_outputs(1707)));
    outputs(9153) <= not(layer0_outputs(10690));
    outputs(9154) <= not(layer0_outputs(4136));
    outputs(9155) <= not(layer0_outputs(2856));
    outputs(9156) <= not(layer0_outputs(3665));
    outputs(9157) <= not(layer0_outputs(3500));
    outputs(9158) <= not(layer0_outputs(1968));
    outputs(9159) <= (layer0_outputs(10770)) and not (layer0_outputs(7465));
    outputs(9160) <= not(layer0_outputs(12597));
    outputs(9161) <= layer0_outputs(11765);
    outputs(9162) <= (layer0_outputs(3029)) xor (layer0_outputs(3670));
    outputs(9163) <= not(layer0_outputs(6237));
    outputs(9164) <= (layer0_outputs(10127)) xor (layer0_outputs(923));
    outputs(9165) <= not(layer0_outputs(4369)) or (layer0_outputs(3052));
    outputs(9166) <= (layer0_outputs(5678)) or (layer0_outputs(3818));
    outputs(9167) <= layer0_outputs(10087);
    outputs(9168) <= '0';
    outputs(9169) <= not((layer0_outputs(10525)) xor (layer0_outputs(2961)));
    outputs(9170) <= layer0_outputs(12159);
    outputs(9171) <= (layer0_outputs(7816)) and not (layer0_outputs(1847));
    outputs(9172) <= layer0_outputs(8233);
    outputs(9173) <= (layer0_outputs(8205)) and not (layer0_outputs(5842));
    outputs(9174) <= not(layer0_outputs(7633));
    outputs(9175) <= not(layer0_outputs(1104));
    outputs(9176) <= (layer0_outputs(1011)) and not (layer0_outputs(2020));
    outputs(9177) <= not((layer0_outputs(3443)) or (layer0_outputs(10545)));
    outputs(9178) <= layer0_outputs(10114);
    outputs(9179) <= layer0_outputs(1649);
    outputs(9180) <= (layer0_outputs(9697)) and (layer0_outputs(6555));
    outputs(9181) <= not(layer0_outputs(3700));
    outputs(9182) <= not((layer0_outputs(4787)) xor (layer0_outputs(12076)));
    outputs(9183) <= '0';
    outputs(9184) <= (layer0_outputs(11)) xor (layer0_outputs(8101));
    outputs(9185) <= (layer0_outputs(11975)) and (layer0_outputs(10705));
    outputs(9186) <= (layer0_outputs(8814)) xor (layer0_outputs(82));
    outputs(9187) <= not(layer0_outputs(4788));
    outputs(9188) <= not(layer0_outputs(9021));
    outputs(9189) <= (layer0_outputs(945)) and not (layer0_outputs(6493));
    outputs(9190) <= layer0_outputs(6600);
    outputs(9191) <= (layer0_outputs(1545)) and (layer0_outputs(11639));
    outputs(9192) <= (layer0_outputs(208)) and not (layer0_outputs(4513));
    outputs(9193) <= not((layer0_outputs(3906)) xor (layer0_outputs(7690)));
    outputs(9194) <= layer0_outputs(8007);
    outputs(9195) <= not((layer0_outputs(1906)) xor (layer0_outputs(2491)));
    outputs(9196) <= (layer0_outputs(1699)) xor (layer0_outputs(8532));
    outputs(9197) <= layer0_outputs(192);
    outputs(9198) <= (layer0_outputs(5666)) xor (layer0_outputs(2894));
    outputs(9199) <= (layer0_outputs(9709)) xor (layer0_outputs(9319));
    outputs(9200) <= not((layer0_outputs(6901)) xor (layer0_outputs(1771)));
    outputs(9201) <= (layer0_outputs(9827)) or (layer0_outputs(3647));
    outputs(9202) <= (layer0_outputs(7256)) and not (layer0_outputs(166));
    outputs(9203) <= not((layer0_outputs(12025)) xor (layer0_outputs(8074)));
    outputs(9204) <= (layer0_outputs(1257)) xor (layer0_outputs(12542));
    outputs(9205) <= not((layer0_outputs(5839)) xor (layer0_outputs(5408)));
    outputs(9206) <= not(layer0_outputs(2406)) or (layer0_outputs(12395));
    outputs(9207) <= layer0_outputs(11582);
    outputs(9208) <= (layer0_outputs(8819)) or (layer0_outputs(667));
    outputs(9209) <= '0';
    outputs(9210) <= layer0_outputs(4603);
    outputs(9211) <= not(layer0_outputs(2560));
    outputs(9212) <= layer0_outputs(205);
    outputs(9213) <= not(layer0_outputs(10322));
    outputs(9214) <= layer0_outputs(10276);
    outputs(9215) <= layer0_outputs(4423);
    outputs(9216) <= layer0_outputs(5924);
    outputs(9217) <= (layer0_outputs(6034)) xor (layer0_outputs(2975));
    outputs(9218) <= not((layer0_outputs(10577)) and (layer0_outputs(7560)));
    outputs(9219) <= layer0_outputs(319);
    outputs(9220) <= not((layer0_outputs(11873)) xor (layer0_outputs(4288)));
    outputs(9221) <= layer0_outputs(2062);
    outputs(9222) <= layer0_outputs(4511);
    outputs(9223) <= (layer0_outputs(12306)) and not (layer0_outputs(6569));
    outputs(9224) <= not(layer0_outputs(2511)) or (layer0_outputs(1439));
    outputs(9225) <= not((layer0_outputs(10218)) xor (layer0_outputs(2989)));
    outputs(9226) <= (layer0_outputs(3007)) and not (layer0_outputs(4492));
    outputs(9227) <= not((layer0_outputs(8310)) xor (layer0_outputs(1363)));
    outputs(9228) <= (layer0_outputs(4550)) xor (layer0_outputs(10696));
    outputs(9229) <= (layer0_outputs(4663)) and (layer0_outputs(4015));
    outputs(9230) <= not((layer0_outputs(8428)) or (layer0_outputs(9370)));
    outputs(9231) <= layer0_outputs(7046);
    outputs(9232) <= layer0_outputs(9991);
    outputs(9233) <= not((layer0_outputs(9551)) xor (layer0_outputs(1557)));
    outputs(9234) <= layer0_outputs(2173);
    outputs(9235) <= layer0_outputs(8305);
    outputs(9236) <= '1';
    outputs(9237) <= layer0_outputs(11210);
    outputs(9238) <= layer0_outputs(5670);
    outputs(9239) <= not((layer0_outputs(12283)) xor (layer0_outputs(11594)));
    outputs(9240) <= not((layer0_outputs(3507)) or (layer0_outputs(7853)));
    outputs(9241) <= (layer0_outputs(8934)) xor (layer0_outputs(1894));
    outputs(9242) <= not((layer0_outputs(386)) xor (layer0_outputs(6645)));
    outputs(9243) <= '0';
    outputs(9244) <= not((layer0_outputs(4995)) xor (layer0_outputs(9964)));
    outputs(9245) <= not(layer0_outputs(2927));
    outputs(9246) <= (layer0_outputs(7424)) xor (layer0_outputs(7637));
    outputs(9247) <= (layer0_outputs(6336)) and not (layer0_outputs(11552));
    outputs(9248) <= (layer0_outputs(6498)) xor (layer0_outputs(12019));
    outputs(9249) <= not((layer0_outputs(9254)) xor (layer0_outputs(4537)));
    outputs(9250) <= layer0_outputs(11724);
    outputs(9251) <= layer0_outputs(4919);
    outputs(9252) <= (layer0_outputs(1992)) and not (layer0_outputs(6095));
    outputs(9253) <= not(layer0_outputs(1258)) or (layer0_outputs(3679));
    outputs(9254) <= (layer0_outputs(10724)) xor (layer0_outputs(1053));
    outputs(9255) <= not(layer0_outputs(2917)) or (layer0_outputs(4969));
    outputs(9256) <= layer0_outputs(11699);
    outputs(9257) <= not((layer0_outputs(12405)) and (layer0_outputs(803)));
    outputs(9258) <= not(layer0_outputs(7858));
    outputs(9259) <= not(layer0_outputs(8449));
    outputs(9260) <= layer0_outputs(3788);
    outputs(9261) <= not(layer0_outputs(11286)) or (layer0_outputs(9767));
    outputs(9262) <= not(layer0_outputs(5385));
    outputs(9263) <= (layer0_outputs(7007)) and not (layer0_outputs(4855));
    outputs(9264) <= not(layer0_outputs(6956)) or (layer0_outputs(2821));
    outputs(9265) <= not(layer0_outputs(12675));
    outputs(9266) <= layer0_outputs(9225);
    outputs(9267) <= not((layer0_outputs(5227)) xor (layer0_outputs(180)));
    outputs(9268) <= not((layer0_outputs(10317)) or (layer0_outputs(7432)));
    outputs(9269) <= not(layer0_outputs(4957));
    outputs(9270) <= not(layer0_outputs(3220));
    outputs(9271) <= (layer0_outputs(4400)) and not (layer0_outputs(11967));
    outputs(9272) <= not(layer0_outputs(1988));
    outputs(9273) <= not(layer0_outputs(1710));
    outputs(9274) <= not(layer0_outputs(5069)) or (layer0_outputs(1465));
    outputs(9275) <= not((layer0_outputs(3659)) xor (layer0_outputs(591)));
    outputs(9276) <= not((layer0_outputs(6473)) xor (layer0_outputs(8249)));
    outputs(9277) <= not((layer0_outputs(8476)) or (layer0_outputs(10242)));
    outputs(9278) <= not((layer0_outputs(8795)) xor (layer0_outputs(11683)));
    outputs(9279) <= not((layer0_outputs(8336)) and (layer0_outputs(2606)));
    outputs(9280) <= (layer0_outputs(5540)) xor (layer0_outputs(6588));
    outputs(9281) <= layer0_outputs(10994);
    outputs(9282) <= (layer0_outputs(6566)) and (layer0_outputs(488));
    outputs(9283) <= not(layer0_outputs(8122));
    outputs(9284) <= (layer0_outputs(3791)) xor (layer0_outputs(736));
    outputs(9285) <= (layer0_outputs(11509)) xor (layer0_outputs(5253));
    outputs(9286) <= not(layer0_outputs(6812));
    outputs(9287) <= not((layer0_outputs(6283)) xor (layer0_outputs(12420)));
    outputs(9288) <= layer0_outputs(12650);
    outputs(9289) <= layer0_outputs(5248);
    outputs(9290) <= layer0_outputs(4793);
    outputs(9291) <= not(layer0_outputs(5251));
    outputs(9292) <= layer0_outputs(1925);
    outputs(9293) <= layer0_outputs(10771);
    outputs(9294) <= (layer0_outputs(12365)) xor (layer0_outputs(11046));
    outputs(9295) <= not(layer0_outputs(9431));
    outputs(9296) <= not(layer0_outputs(7542));
    outputs(9297) <= layer0_outputs(1848);
    outputs(9298) <= not(layer0_outputs(3447));
    outputs(9299) <= not((layer0_outputs(7953)) or (layer0_outputs(7438)));
    outputs(9300) <= (layer0_outputs(8392)) or (layer0_outputs(11900));
    outputs(9301) <= not(layer0_outputs(4654));
    outputs(9302) <= not(layer0_outputs(2125));
    outputs(9303) <= not((layer0_outputs(3544)) or (layer0_outputs(9112)));
    outputs(9304) <= (layer0_outputs(7755)) and (layer0_outputs(8996));
    outputs(9305) <= not(layer0_outputs(3196));
    outputs(9306) <= layer0_outputs(7818);
    outputs(9307) <= not((layer0_outputs(2412)) or (layer0_outputs(7712)));
    outputs(9308) <= not((layer0_outputs(7942)) xor (layer0_outputs(11427)));
    outputs(9309) <= (layer0_outputs(12304)) and (layer0_outputs(5000));
    outputs(9310) <= not(layer0_outputs(12616)) or (layer0_outputs(10451));
    outputs(9311) <= (layer0_outputs(2229)) and not (layer0_outputs(12644));
    outputs(9312) <= not(layer0_outputs(3889));
    outputs(9313) <= (layer0_outputs(8750)) and not (layer0_outputs(6317));
    outputs(9314) <= (layer0_outputs(10385)) or (layer0_outputs(3655));
    outputs(9315) <= not(layer0_outputs(4930));
    outputs(9316) <= not(layer0_outputs(6967));
    outputs(9317) <= not(layer0_outputs(8573));
    outputs(9318) <= not(layer0_outputs(2881));
    outputs(9319) <= layer0_outputs(5776);
    outputs(9320) <= layer0_outputs(3311);
    outputs(9321) <= layer0_outputs(1830);
    outputs(9322) <= not(layer0_outputs(3337)) or (layer0_outputs(1241));
    outputs(9323) <= layer0_outputs(3174);
    outputs(9324) <= not((layer0_outputs(2292)) xor (layer0_outputs(9905)));
    outputs(9325) <= not(layer0_outputs(10498));
    outputs(9326) <= not(layer0_outputs(6042)) or (layer0_outputs(4555));
    outputs(9327) <= (layer0_outputs(8071)) and not (layer0_outputs(3753));
    outputs(9328) <= not((layer0_outputs(4665)) or (layer0_outputs(7891)));
    outputs(9329) <= (layer0_outputs(8448)) or (layer0_outputs(2142));
    outputs(9330) <= not((layer0_outputs(12416)) xor (layer0_outputs(10878)));
    outputs(9331) <= layer0_outputs(2885);
    outputs(9332) <= not(layer0_outputs(1898));
    outputs(9333) <= '1';
    outputs(9334) <= not(layer0_outputs(9190));
    outputs(9335) <= not(layer0_outputs(7123)) or (layer0_outputs(1907));
    outputs(9336) <= layer0_outputs(2629);
    outputs(9337) <= not(layer0_outputs(958));
    outputs(9338) <= not((layer0_outputs(6974)) or (layer0_outputs(2772)));
    outputs(9339) <= not(layer0_outputs(12402));
    outputs(9340) <= (layer0_outputs(2872)) xor (layer0_outputs(5966));
    outputs(9341) <= not(layer0_outputs(238));
    outputs(9342) <= not(layer0_outputs(10360)) or (layer0_outputs(5349));
    outputs(9343) <= (layer0_outputs(1479)) and not (layer0_outputs(8798));
    outputs(9344) <= layer0_outputs(1375);
    outputs(9345) <= not(layer0_outputs(9847));
    outputs(9346) <= layer0_outputs(12356);
    outputs(9347) <= not(layer0_outputs(3517));
    outputs(9348) <= not(layer0_outputs(3551));
    outputs(9349) <= not(layer0_outputs(2452));
    outputs(9350) <= not((layer0_outputs(10388)) xor (layer0_outputs(1269)));
    outputs(9351) <= (layer0_outputs(2615)) and (layer0_outputs(6548));
    outputs(9352) <= not(layer0_outputs(9521));
    outputs(9353) <= (layer0_outputs(5676)) and not (layer0_outputs(12065));
    outputs(9354) <= not(layer0_outputs(9584));
    outputs(9355) <= not((layer0_outputs(589)) xor (layer0_outputs(8265)));
    outputs(9356) <= layer0_outputs(8488);
    outputs(9357) <= layer0_outputs(5751);
    outputs(9358) <= layer0_outputs(2980);
    outputs(9359) <= (layer0_outputs(6039)) and not (layer0_outputs(5701));
    outputs(9360) <= not((layer0_outputs(11112)) xor (layer0_outputs(7351)));
    outputs(9361) <= (layer0_outputs(12080)) and not (layer0_outputs(11370));
    outputs(9362) <= not((layer0_outputs(3996)) xor (layer0_outputs(11712)));
    outputs(9363) <= not(layer0_outputs(8706));
    outputs(9364) <= not((layer0_outputs(2254)) and (layer0_outputs(1112)));
    outputs(9365) <= (layer0_outputs(2102)) and not (layer0_outputs(9920));
    outputs(9366) <= not(layer0_outputs(6200));
    outputs(9367) <= not(layer0_outputs(316));
    outputs(9368) <= (layer0_outputs(2674)) and not (layer0_outputs(9615));
    outputs(9369) <= (layer0_outputs(11008)) and (layer0_outputs(6426));
    outputs(9370) <= (layer0_outputs(11520)) xor (layer0_outputs(6629));
    outputs(9371) <= not((layer0_outputs(9386)) xor (layer0_outputs(3272)));
    outputs(9372) <= not((layer0_outputs(12041)) xor (layer0_outputs(1255)));
    outputs(9373) <= not(layer0_outputs(498)) or (layer0_outputs(3824));
    outputs(9374) <= layer0_outputs(9318);
    outputs(9375) <= not(layer0_outputs(9063));
    outputs(9376) <= not(layer0_outputs(1469));
    outputs(9377) <= not(layer0_outputs(10094));
    outputs(9378) <= layer0_outputs(5751);
    outputs(9379) <= layer0_outputs(12603);
    outputs(9380) <= not((layer0_outputs(8221)) xor (layer0_outputs(10677)));
    outputs(9381) <= (layer0_outputs(11351)) xor (layer0_outputs(2515));
    outputs(9382) <= layer0_outputs(11503);
    outputs(9383) <= layer0_outputs(2969);
    outputs(9384) <= not(layer0_outputs(6190));
    outputs(9385) <= not((layer0_outputs(6108)) xor (layer0_outputs(4396)));
    outputs(9386) <= not(layer0_outputs(3289));
    outputs(9387) <= layer0_outputs(6457);
    outputs(9388) <= not(layer0_outputs(1169));
    outputs(9389) <= layer0_outputs(427);
    outputs(9390) <= not((layer0_outputs(4970)) xor (layer0_outputs(10386)));
    outputs(9391) <= (layer0_outputs(9862)) and not (layer0_outputs(1775));
    outputs(9392) <= not(layer0_outputs(7084));
    outputs(9393) <= '0';
    outputs(9394) <= not(layer0_outputs(9487));
    outputs(9395) <= (layer0_outputs(6592)) xor (layer0_outputs(4755));
    outputs(9396) <= not((layer0_outputs(12)) or (layer0_outputs(2179)));
    outputs(9397) <= not(layer0_outputs(227));
    outputs(9398) <= not((layer0_outputs(9902)) and (layer0_outputs(4600)));
    outputs(9399) <= layer0_outputs(12459);
    outputs(9400) <= not((layer0_outputs(10510)) xor (layer0_outputs(8833)));
    outputs(9401) <= layer0_outputs(8833);
    outputs(9402) <= not((layer0_outputs(6018)) xor (layer0_outputs(8331)));
    outputs(9403) <= (layer0_outputs(9519)) and (layer0_outputs(11056));
    outputs(9404) <= (layer0_outputs(3114)) xor (layer0_outputs(915));
    outputs(9405) <= layer0_outputs(8803);
    outputs(9406) <= layer0_outputs(11100);
    outputs(9407) <= (layer0_outputs(8764)) and not (layer0_outputs(6664));
    outputs(9408) <= (layer0_outputs(7212)) and (layer0_outputs(9447));
    outputs(9409) <= not((layer0_outputs(8452)) or (layer0_outputs(9707)));
    outputs(9410) <= layer0_outputs(11285);
    outputs(9411) <= (layer0_outputs(12112)) and not (layer0_outputs(10097));
    outputs(9412) <= (layer0_outputs(1676)) xor (layer0_outputs(7569));
    outputs(9413) <= (layer0_outputs(174)) and not (layer0_outputs(6501));
    outputs(9414) <= not((layer0_outputs(582)) xor (layer0_outputs(7014)));
    outputs(9415) <= not(layer0_outputs(1103));
    outputs(9416) <= not((layer0_outputs(10879)) xor (layer0_outputs(11336)));
    outputs(9417) <= not(layer0_outputs(8541));
    outputs(9418) <= (layer0_outputs(6472)) xor (layer0_outputs(4840));
    outputs(9419) <= not(layer0_outputs(10039));
    outputs(9420) <= (layer0_outputs(1961)) and not (layer0_outputs(6365));
    outputs(9421) <= layer0_outputs(8570);
    outputs(9422) <= layer0_outputs(7821);
    outputs(9423) <= not(layer0_outputs(8660));
    outputs(9424) <= not((layer0_outputs(4267)) or (layer0_outputs(1732)));
    outputs(9425) <= not((layer0_outputs(8703)) or (layer0_outputs(3367)));
    outputs(9426) <= (layer0_outputs(11071)) and not (layer0_outputs(3311));
    outputs(9427) <= not((layer0_outputs(11238)) xor (layer0_outputs(5895)));
    outputs(9428) <= (layer0_outputs(8666)) and not (layer0_outputs(3577));
    outputs(9429) <= (layer0_outputs(6622)) and not (layer0_outputs(2888));
    outputs(9430) <= layer0_outputs(5366);
    outputs(9431) <= (layer0_outputs(8583)) or (layer0_outputs(5916));
    outputs(9432) <= layer0_outputs(10372);
    outputs(9433) <= layer0_outputs(11670);
    outputs(9434) <= not((layer0_outputs(6888)) xor (layer0_outputs(7211)));
    outputs(9435) <= not(layer0_outputs(9564));
    outputs(9436) <= not((layer0_outputs(1712)) or (layer0_outputs(12098)));
    outputs(9437) <= layer0_outputs(5680);
    outputs(9438) <= layer0_outputs(4821);
    outputs(9439) <= (layer0_outputs(8478)) and not (layer0_outputs(6513));
    outputs(9440) <= (layer0_outputs(9172)) and (layer0_outputs(11863));
    outputs(9441) <= not(layer0_outputs(9923));
    outputs(9442) <= (layer0_outputs(12085)) and (layer0_outputs(4326));
    outputs(9443) <= not(layer0_outputs(8807)) or (layer0_outputs(9850));
    outputs(9444) <= not(layer0_outputs(9894)) or (layer0_outputs(4710));
    outputs(9445) <= not((layer0_outputs(3030)) xor (layer0_outputs(8040)));
    outputs(9446) <= not((layer0_outputs(6461)) xor (layer0_outputs(8663)));
    outputs(9447) <= not(layer0_outputs(7673));
    outputs(9448) <= layer0_outputs(11650);
    outputs(9449) <= layer0_outputs(8430);
    outputs(9450) <= (layer0_outputs(8438)) and not (layer0_outputs(5862));
    outputs(9451) <= (layer0_outputs(1063)) and not (layer0_outputs(5921));
    outputs(9452) <= not(layer0_outputs(5763));
    outputs(9453) <= (layer0_outputs(3844)) xor (layer0_outputs(11075));
    outputs(9454) <= layer0_outputs(5339);
    outputs(9455) <= '1';
    outputs(9456) <= layer0_outputs(10251);
    outputs(9457) <= (layer0_outputs(12108)) and not (layer0_outputs(2125));
    outputs(9458) <= not((layer0_outputs(964)) or (layer0_outputs(5349)));
    outputs(9459) <= not(layer0_outputs(3980));
    outputs(9460) <= layer0_outputs(12792);
    outputs(9461) <= layer0_outputs(11007);
    outputs(9462) <= not(layer0_outputs(10497));
    outputs(9463) <= (layer0_outputs(10893)) or (layer0_outputs(3436));
    outputs(9464) <= not(layer0_outputs(11613));
    outputs(9465) <= layer0_outputs(10049);
    outputs(9466) <= (layer0_outputs(21)) and not (layer0_outputs(10991));
    outputs(9467) <= not(layer0_outputs(49));
    outputs(9468) <= layer0_outputs(5451);
    outputs(9469) <= not((layer0_outputs(8495)) or (layer0_outputs(8869)));
    outputs(9470) <= (layer0_outputs(2634)) and (layer0_outputs(4225));
    outputs(9471) <= not((layer0_outputs(11174)) or (layer0_outputs(4633)));
    outputs(9472) <= layer0_outputs(12385);
    outputs(9473) <= layer0_outputs(4585);
    outputs(9474) <= not((layer0_outputs(8946)) xor (layer0_outputs(4062)));
    outputs(9475) <= not((layer0_outputs(11123)) xor (layer0_outputs(3097)));
    outputs(9476) <= layer0_outputs(12153);
    outputs(9477) <= layer0_outputs(1770);
    outputs(9478) <= (layer0_outputs(4918)) and not (layer0_outputs(11206));
    outputs(9479) <= (layer0_outputs(10839)) and not (layer0_outputs(8598));
    outputs(9480) <= not(layer0_outputs(7084));
    outputs(9481) <= not(layer0_outputs(2120)) or (layer0_outputs(2379));
    outputs(9482) <= layer0_outputs(11832);
    outputs(9483) <= (layer0_outputs(6859)) and not (layer0_outputs(387));
    outputs(9484) <= not(layer0_outputs(376));
    outputs(9485) <= not(layer0_outputs(5443));
    outputs(9486) <= not((layer0_outputs(11170)) xor (layer0_outputs(12007)));
    outputs(9487) <= not((layer0_outputs(7028)) and (layer0_outputs(10970)));
    outputs(9488) <= (layer0_outputs(8912)) and not (layer0_outputs(2204));
    outputs(9489) <= layer0_outputs(493);
    outputs(9490) <= not((layer0_outputs(573)) or (layer0_outputs(3134)));
    outputs(9491) <= layer0_outputs(6674);
    outputs(9492) <= not(layer0_outputs(11572)) or (layer0_outputs(6143));
    outputs(9493) <= layer0_outputs(11796);
    outputs(9494) <= '0';
    outputs(9495) <= not(layer0_outputs(7686)) or (layer0_outputs(8584));
    outputs(9496) <= not((layer0_outputs(1759)) or (layer0_outputs(3382)));
    outputs(9497) <= not((layer0_outputs(3410)) xor (layer0_outputs(12592)));
    outputs(9498) <= layer0_outputs(11356);
    outputs(9499) <= layer0_outputs(2063);
    outputs(9500) <= not(layer0_outputs(9814));
    outputs(9501) <= not(layer0_outputs(10774));
    outputs(9502) <= (layer0_outputs(12479)) and (layer0_outputs(7855));
    outputs(9503) <= not((layer0_outputs(7993)) xor (layer0_outputs(12453)));
    outputs(9504) <= not((layer0_outputs(1803)) and (layer0_outputs(12753)));
    outputs(9505) <= layer0_outputs(5448);
    outputs(9506) <= not(layer0_outputs(11510));
    outputs(9507) <= not(layer0_outputs(5950));
    outputs(9508) <= not((layer0_outputs(10909)) or (layer0_outputs(11131)));
    outputs(9509) <= (layer0_outputs(5677)) and (layer0_outputs(871));
    outputs(9510) <= not(layer0_outputs(6313));
    outputs(9511) <= not(layer0_outputs(50));
    outputs(9512) <= (layer0_outputs(7476)) xor (layer0_outputs(9876));
    outputs(9513) <= not((layer0_outputs(1696)) xor (layer0_outputs(9284)));
    outputs(9514) <= (layer0_outputs(7911)) or (layer0_outputs(12776));
    outputs(9515) <= not(layer0_outputs(4640));
    outputs(9516) <= layer0_outputs(3497);
    outputs(9517) <= not((layer0_outputs(9143)) or (layer0_outputs(9976)));
    outputs(9518) <= not(layer0_outputs(2328));
    outputs(9519) <= not(layer0_outputs(11344));
    outputs(9520) <= (layer0_outputs(8261)) xor (layer0_outputs(2673));
    outputs(9521) <= not(layer0_outputs(3571));
    outputs(9522) <= not(layer0_outputs(10819));
    outputs(9523) <= not(layer0_outputs(3207)) or (layer0_outputs(4704));
    outputs(9524) <= not((layer0_outputs(10940)) xor (layer0_outputs(2956)));
    outputs(9525) <= not((layer0_outputs(6198)) xor (layer0_outputs(7877)));
    outputs(9526) <= (layer0_outputs(3620)) and not (layer0_outputs(4298));
    outputs(9527) <= (layer0_outputs(10622)) and not (layer0_outputs(4054));
    outputs(9528) <= (layer0_outputs(12451)) xor (layer0_outputs(10266));
    outputs(9529) <= not((layer0_outputs(6978)) xor (layer0_outputs(1626)));
    outputs(9530) <= not((layer0_outputs(11312)) xor (layer0_outputs(9795)));
    outputs(9531) <= (layer0_outputs(3625)) xor (layer0_outputs(11304));
    outputs(9532) <= not(layer0_outputs(12424));
    outputs(9533) <= (layer0_outputs(6865)) and (layer0_outputs(6836));
    outputs(9534) <= layer0_outputs(7802);
    outputs(9535) <= not(layer0_outputs(3297));
    outputs(9536) <= not((layer0_outputs(11606)) and (layer0_outputs(12059)));
    outputs(9537) <= not(layer0_outputs(5327));
    outputs(9538) <= not((layer0_outputs(2488)) xor (layer0_outputs(8879)));
    outputs(9539) <= not(layer0_outputs(8159));
    outputs(9540) <= layer0_outputs(10087);
    outputs(9541) <= (layer0_outputs(4077)) and (layer0_outputs(10652));
    outputs(9542) <= (layer0_outputs(5690)) and not (layer0_outputs(3237));
    outputs(9543) <= layer0_outputs(10610);
    outputs(9544) <= not((layer0_outputs(3111)) or (layer0_outputs(1174)));
    outputs(9545) <= not(layer0_outputs(10520));
    outputs(9546) <= (layer0_outputs(5093)) xor (layer0_outputs(10848));
    outputs(9547) <= (layer0_outputs(1362)) and not (layer0_outputs(5684));
    outputs(9548) <= layer0_outputs(4239);
    outputs(9549) <= not(layer0_outputs(3329)) or (layer0_outputs(4035));
    outputs(9550) <= layer0_outputs(666);
    outputs(9551) <= (layer0_outputs(3337)) and not (layer0_outputs(2404));
    outputs(9552) <= (layer0_outputs(6617)) or (layer0_outputs(9073));
    outputs(9553) <= not(layer0_outputs(5574));
    outputs(9554) <= (layer0_outputs(12795)) xor (layer0_outputs(6295));
    outputs(9555) <= not((layer0_outputs(239)) xor (layer0_outputs(11161)));
    outputs(9556) <= not(layer0_outputs(5544));
    outputs(9557) <= (layer0_outputs(2749)) and not (layer0_outputs(11309));
    outputs(9558) <= not(layer0_outputs(5967));
    outputs(9559) <= not((layer0_outputs(1295)) xor (layer0_outputs(10386)));
    outputs(9560) <= (layer0_outputs(298)) xor (layer0_outputs(8647));
    outputs(9561) <= (layer0_outputs(1602)) and not (layer0_outputs(12500));
    outputs(9562) <= '0';
    outputs(9563) <= (layer0_outputs(8308)) and not (layer0_outputs(7545));
    outputs(9564) <= layer0_outputs(5210);
    outputs(9565) <= not(layer0_outputs(2038));
    outputs(9566) <= not((layer0_outputs(3796)) xor (layer0_outputs(7905)));
    outputs(9567) <= (layer0_outputs(1087)) and not (layer0_outputs(897));
    outputs(9568) <= layer0_outputs(8411);
    outputs(9569) <= not((layer0_outputs(11324)) xor (layer0_outputs(8078)));
    outputs(9570) <= not(layer0_outputs(12637));
    outputs(9571) <= not((layer0_outputs(4575)) xor (layer0_outputs(6662)));
    outputs(9572) <= not(layer0_outputs(2732));
    outputs(9573) <= (layer0_outputs(6433)) and not (layer0_outputs(3267));
    outputs(9574) <= layer0_outputs(6286);
    outputs(9575) <= layer0_outputs(3783);
    outputs(9576) <= layer0_outputs(1047);
    outputs(9577) <= layer0_outputs(2836);
    outputs(9578) <= (layer0_outputs(11332)) and (layer0_outputs(7793));
    outputs(9579) <= not((layer0_outputs(1218)) and (layer0_outputs(7494)));
    outputs(9580) <= layer0_outputs(7970);
    outputs(9581) <= (layer0_outputs(6695)) and not (layer0_outputs(687));
    outputs(9582) <= not(layer0_outputs(2044));
    outputs(9583) <= not(layer0_outputs(4070));
    outputs(9584) <= (layer0_outputs(20)) and not (layer0_outputs(10265));
    outputs(9585) <= (layer0_outputs(10519)) and not (layer0_outputs(2100));
    outputs(9586) <= not(layer0_outputs(8563));
    outputs(9587) <= not(layer0_outputs(4224));
    outputs(9588) <= (layer0_outputs(10850)) or (layer0_outputs(4086));
    outputs(9589) <= (layer0_outputs(1201)) xor (layer0_outputs(11123));
    outputs(9590) <= not((layer0_outputs(3427)) xor (layer0_outputs(7381)));
    outputs(9591) <= (layer0_outputs(9753)) or (layer0_outputs(8296));
    outputs(9592) <= not(layer0_outputs(5768));
    outputs(9593) <= not(layer0_outputs(2620));
    outputs(9594) <= (layer0_outputs(10161)) xor (layer0_outputs(8374));
    outputs(9595) <= not(layer0_outputs(2676));
    outputs(9596) <= not(layer0_outputs(3058)) or (layer0_outputs(5505));
    outputs(9597) <= not((layer0_outputs(6450)) or (layer0_outputs(4863)));
    outputs(9598) <= not((layer0_outputs(2889)) xor (layer0_outputs(2384)));
    outputs(9599) <= (layer0_outputs(2803)) xor (layer0_outputs(995));
    outputs(9600) <= not(layer0_outputs(1432));
    outputs(9601) <= not(layer0_outputs(2490));
    outputs(9602) <= layer0_outputs(11150);
    outputs(9603) <= (layer0_outputs(4168)) and not (layer0_outputs(8904));
    outputs(9604) <= (layer0_outputs(8770)) and (layer0_outputs(4227));
    outputs(9605) <= (layer0_outputs(12631)) and not (layer0_outputs(3419));
    outputs(9606) <= layer0_outputs(9387);
    outputs(9607) <= not((layer0_outputs(2835)) or (layer0_outputs(11915)));
    outputs(9608) <= not(layer0_outputs(3193));
    outputs(9609) <= (layer0_outputs(7768)) xor (layer0_outputs(5125));
    outputs(9610) <= (layer0_outputs(645)) and not (layer0_outputs(10692));
    outputs(9611) <= not((layer0_outputs(3945)) or (layer0_outputs(8512)));
    outputs(9612) <= layer0_outputs(2421);
    outputs(9613) <= not(layer0_outputs(6129));
    outputs(9614) <= (layer0_outputs(9597)) and not (layer0_outputs(11660));
    outputs(9615) <= not((layer0_outputs(7874)) and (layer0_outputs(10849)));
    outputs(9616) <= not(layer0_outputs(9250));
    outputs(9617) <= not((layer0_outputs(3771)) or (layer0_outputs(6399)));
    outputs(9618) <= not(layer0_outputs(6769));
    outputs(9619) <= not((layer0_outputs(1024)) or (layer0_outputs(2735)));
    outputs(9620) <= not((layer0_outputs(2901)) or (layer0_outputs(8878)));
    outputs(9621) <= layer0_outputs(4436);
    outputs(9622) <= layer0_outputs(10924);
    outputs(9623) <= layer0_outputs(9117);
    outputs(9624) <= not((layer0_outputs(45)) or (layer0_outputs(1641)));
    outputs(9625) <= not(layer0_outputs(5473));
    outputs(9626) <= not((layer0_outputs(11938)) or (layer0_outputs(5295)));
    outputs(9627) <= not(layer0_outputs(10322));
    outputs(9628) <= (layer0_outputs(11976)) xor (layer0_outputs(90));
    outputs(9629) <= not(layer0_outputs(6717));
    outputs(9630) <= not(layer0_outputs(2983));
    outputs(9631) <= (layer0_outputs(10605)) and not (layer0_outputs(4967));
    outputs(9632) <= not((layer0_outputs(9457)) xor (layer0_outputs(4933)));
    outputs(9633) <= not(layer0_outputs(10743));
    outputs(9634) <= (layer0_outputs(7481)) and (layer0_outputs(3981));
    outputs(9635) <= not((layer0_outputs(3915)) xor (layer0_outputs(7905)));
    outputs(9636) <= not((layer0_outputs(655)) or (layer0_outputs(8164)));
    outputs(9637) <= not((layer0_outputs(2288)) xor (layer0_outputs(869)));
    outputs(9638) <= not(layer0_outputs(11133));
    outputs(9639) <= layer0_outputs(2572);
    outputs(9640) <= (layer0_outputs(3814)) and not (layer0_outputs(5050));
    outputs(9641) <= (layer0_outputs(12622)) and (layer0_outputs(9466));
    outputs(9642) <= not(layer0_outputs(687));
    outputs(9643) <= not((layer0_outputs(3691)) xor (layer0_outputs(7752)));
    outputs(9644) <= (layer0_outputs(12203)) and not (layer0_outputs(1924));
    outputs(9645) <= not(layer0_outputs(328));
    outputs(9646) <= not((layer0_outputs(3292)) and (layer0_outputs(1263)));
    outputs(9647) <= not(layer0_outputs(9008)) or (layer0_outputs(5123));
    outputs(9648) <= layer0_outputs(12745);
    outputs(9649) <= not((layer0_outputs(5576)) xor (layer0_outputs(11000)));
    outputs(9650) <= (layer0_outputs(1171)) and not (layer0_outputs(11494));
    outputs(9651) <= (layer0_outputs(9020)) and not (layer0_outputs(6071));
    outputs(9652) <= not(layer0_outputs(5989));
    outputs(9653) <= layer0_outputs(5599);
    outputs(9654) <= not(layer0_outputs(11887));
    outputs(9655) <= not((layer0_outputs(9712)) or (layer0_outputs(9100)));
    outputs(9656) <= not((layer0_outputs(7644)) xor (layer0_outputs(5991)));
    outputs(9657) <= layer0_outputs(2971);
    outputs(9658) <= (layer0_outputs(8554)) xor (layer0_outputs(3550));
    outputs(9659) <= (layer0_outputs(534)) and (layer0_outputs(10974));
    outputs(9660) <= layer0_outputs(1694);
    outputs(9661) <= not((layer0_outputs(7407)) xor (layer0_outputs(11349)));
    outputs(9662) <= (layer0_outputs(5035)) xor (layer0_outputs(11311));
    outputs(9663) <= (layer0_outputs(85)) and not (layer0_outputs(7854));
    outputs(9664) <= not(layer0_outputs(9527));
    outputs(9665) <= not(layer0_outputs(5634)) or (layer0_outputs(3373));
    outputs(9666) <= layer0_outputs(6762);
    outputs(9667) <= not(layer0_outputs(833));
    outputs(9668) <= not(layer0_outputs(8621));
    outputs(9669) <= (layer0_outputs(8072)) xor (layer0_outputs(10602));
    outputs(9670) <= not((layer0_outputs(12787)) xor (layer0_outputs(2858)));
    outputs(9671) <= (layer0_outputs(11677)) and not (layer0_outputs(3674));
    outputs(9672) <= not((layer0_outputs(7218)) xor (layer0_outputs(8537)));
    outputs(9673) <= not(layer0_outputs(683));
    outputs(9674) <= not((layer0_outputs(1234)) xor (layer0_outputs(3513)));
    outputs(9675) <= layer0_outputs(7977);
    outputs(9676) <= layer0_outputs(6903);
    outputs(9677) <= (layer0_outputs(11653)) and not (layer0_outputs(8354));
    outputs(9678) <= not(layer0_outputs(3586));
    outputs(9679) <= (layer0_outputs(1405)) and not (layer0_outputs(5713));
    outputs(9680) <= not((layer0_outputs(4764)) xor (layer0_outputs(11384)));
    outputs(9681) <= not((layer0_outputs(3891)) and (layer0_outputs(5052)));
    outputs(9682) <= layer0_outputs(7493);
    outputs(9683) <= (layer0_outputs(7569)) xor (layer0_outputs(11827));
    outputs(9684) <= layer0_outputs(9748);
    outputs(9685) <= layer0_outputs(9119);
    outputs(9686) <= layer0_outputs(775);
    outputs(9687) <= layer0_outputs(4222);
    outputs(9688) <= (layer0_outputs(7347)) and not (layer0_outputs(7561));
    outputs(9689) <= (layer0_outputs(5699)) or (layer0_outputs(9014));
    outputs(9690) <= layer0_outputs(5104);
    outputs(9691) <= not(layer0_outputs(1899));
    outputs(9692) <= layer0_outputs(2776);
    outputs(9693) <= layer0_outputs(7017);
    outputs(9694) <= (layer0_outputs(8859)) xor (layer0_outputs(502));
    outputs(9695) <= layer0_outputs(8752);
    outputs(9696) <= layer0_outputs(4129);
    outputs(9697) <= not(layer0_outputs(5626));
    outputs(9698) <= not(layer0_outputs(4049));
    outputs(9699) <= not(layer0_outputs(11922));
    outputs(9700) <= not(layer0_outputs(8718));
    outputs(9701) <= (layer0_outputs(3148)) xor (layer0_outputs(5065));
    outputs(9702) <= not(layer0_outputs(6211));
    outputs(9703) <= not((layer0_outputs(8994)) or (layer0_outputs(6158)));
    outputs(9704) <= not(layer0_outputs(9229));
    outputs(9705) <= (layer0_outputs(1988)) and not (layer0_outputs(3808));
    outputs(9706) <= not(layer0_outputs(10232));
    outputs(9707) <= not(layer0_outputs(1179));
    outputs(9708) <= layer0_outputs(5855);
    outputs(9709) <= not(layer0_outputs(429)) or (layer0_outputs(9921));
    outputs(9710) <= not(layer0_outputs(7743));
    outputs(9711) <= layer0_outputs(2992);
    outputs(9712) <= not(layer0_outputs(5526));
    outputs(9713) <= (layer0_outputs(6531)) xor (layer0_outputs(4858));
    outputs(9714) <= not(layer0_outputs(12318));
    outputs(9715) <= not(layer0_outputs(3065)) or (layer0_outputs(8188));
    outputs(9716) <= layer0_outputs(11733);
    outputs(9717) <= not(layer0_outputs(12004)) or (layer0_outputs(5420));
    outputs(9718) <= (layer0_outputs(7351)) xor (layer0_outputs(1198));
    outputs(9719) <= not((layer0_outputs(4959)) xor (layer0_outputs(4091)));
    outputs(9720) <= (layer0_outputs(11297)) xor (layer0_outputs(9848));
    outputs(9721) <= layer0_outputs(2766);
    outputs(9722) <= (layer0_outputs(203)) and not (layer0_outputs(11225));
    outputs(9723) <= not(layer0_outputs(6687));
    outputs(9724) <= not(layer0_outputs(10942));
    outputs(9725) <= (layer0_outputs(8562)) xor (layer0_outputs(5219));
    outputs(9726) <= (layer0_outputs(6345)) or (layer0_outputs(11463));
    outputs(9727) <= not((layer0_outputs(9725)) xor (layer0_outputs(5764)));
    outputs(9728) <= layer0_outputs(2567);
    outputs(9729) <= not((layer0_outputs(11622)) xor (layer0_outputs(3716)));
    outputs(9730) <= not(layer0_outputs(5850));
    outputs(9731) <= not((layer0_outputs(12422)) or (layer0_outputs(11288)));
    outputs(9732) <= not(layer0_outputs(12527));
    outputs(9733) <= (layer0_outputs(42)) and not (layer0_outputs(4480));
    outputs(9734) <= not(layer0_outputs(226));
    outputs(9735) <= not((layer0_outputs(11923)) xor (layer0_outputs(9302)));
    outputs(9736) <= (layer0_outputs(326)) xor (layer0_outputs(2023));
    outputs(9737) <= (layer0_outputs(11862)) and not (layer0_outputs(7491));
    outputs(9738) <= layer0_outputs(8954);
    outputs(9739) <= not((layer0_outputs(7317)) xor (layer0_outputs(4296)));
    outputs(9740) <= not((layer0_outputs(2438)) xor (layer0_outputs(11695)));
    outputs(9741) <= layer0_outputs(5677);
    outputs(9742) <= not((layer0_outputs(11414)) xor (layer0_outputs(11603)));
    outputs(9743) <= not(layer0_outputs(4414));
    outputs(9744) <= (layer0_outputs(3656)) and (layer0_outputs(1951));
    outputs(9745) <= not((layer0_outputs(6513)) xor (layer0_outputs(1334)));
    outputs(9746) <= not((layer0_outputs(7896)) xor (layer0_outputs(12756)));
    outputs(9747) <= not(layer0_outputs(10653));
    outputs(9748) <= not(layer0_outputs(2285));
    outputs(9749) <= not(layer0_outputs(11623));
    outputs(9750) <= not(layer0_outputs(11158));
    outputs(9751) <= not(layer0_outputs(2838)) or (layer0_outputs(4911));
    outputs(9752) <= not(layer0_outputs(4243));
    outputs(9753) <= (layer0_outputs(10634)) and not (layer0_outputs(4900));
    outputs(9754) <= (layer0_outputs(12178)) xor (layer0_outputs(5842));
    outputs(9755) <= not((layer0_outputs(2594)) xor (layer0_outputs(10026)));
    outputs(9756) <= not(layer0_outputs(7153));
    outputs(9757) <= layer0_outputs(3075);
    outputs(9758) <= not((layer0_outputs(9746)) or (layer0_outputs(9616)));
    outputs(9759) <= not((layer0_outputs(8539)) or (layer0_outputs(8094)));
    outputs(9760) <= (layer0_outputs(9707)) or (layer0_outputs(1790));
    outputs(9761) <= not((layer0_outputs(12297)) xor (layer0_outputs(6125)));
    outputs(9762) <= not(layer0_outputs(11092));
    outputs(9763) <= layer0_outputs(8189);
    outputs(9764) <= (layer0_outputs(11301)) xor (layer0_outputs(3279));
    outputs(9765) <= not(layer0_outputs(2521));
    outputs(9766) <= layer0_outputs(4597);
    outputs(9767) <= (layer0_outputs(4619)) xor (layer0_outputs(3635));
    outputs(9768) <= not(layer0_outputs(12341));
    outputs(9769) <= layer0_outputs(5083);
    outputs(9770) <= layer0_outputs(2105);
    outputs(9771) <= layer0_outputs(872);
    outputs(9772) <= not(layer0_outputs(6946));
    outputs(9773) <= (layer0_outputs(7557)) xor (layer0_outputs(4836));
    outputs(9774) <= layer0_outputs(11307);
    outputs(9775) <= (layer0_outputs(12184)) and not (layer0_outputs(11027));
    outputs(9776) <= not((layer0_outputs(5320)) xor (layer0_outputs(2053)));
    outputs(9777) <= layer0_outputs(785);
    outputs(9778) <= (layer0_outputs(3194)) xor (layer0_outputs(2237));
    outputs(9779) <= '0';
    outputs(9780) <= not(layer0_outputs(3867)) or (layer0_outputs(10295));
    outputs(9781) <= not(layer0_outputs(9090));
    outputs(9782) <= not((layer0_outputs(4039)) xor (layer0_outputs(10337)));
    outputs(9783) <= not((layer0_outputs(14)) xor (layer0_outputs(3353)));
    outputs(9784) <= not(layer0_outputs(9310));
    outputs(9785) <= (layer0_outputs(7442)) xor (layer0_outputs(8852));
    outputs(9786) <= not(layer0_outputs(11340));
    outputs(9787) <= not(layer0_outputs(8466));
    outputs(9788) <= layer0_outputs(11644);
    outputs(9789) <= not((layer0_outputs(5369)) xor (layer0_outputs(10981)));
    outputs(9790) <= layer0_outputs(11849);
    outputs(9791) <= not(layer0_outputs(3732)) or (layer0_outputs(2596));
    outputs(9792) <= (layer0_outputs(6811)) and not (layer0_outputs(10351));
    outputs(9793) <= (layer0_outputs(6035)) xor (layer0_outputs(12681));
    outputs(9794) <= (layer0_outputs(9364)) and (layer0_outputs(9994));
    outputs(9795) <= not((layer0_outputs(1810)) xor (layer0_outputs(7713)));
    outputs(9796) <= not(layer0_outputs(7360));
    outputs(9797) <= (layer0_outputs(7790)) xor (layer0_outputs(9396));
    outputs(9798) <= not(layer0_outputs(2826));
    outputs(9799) <= (layer0_outputs(4337)) and (layer0_outputs(3846));
    outputs(9800) <= (layer0_outputs(6694)) and (layer0_outputs(5286));
    outputs(9801) <= not(layer0_outputs(2028));
    outputs(9802) <= (layer0_outputs(6609)) and not (layer0_outputs(1469));
    outputs(9803) <= not((layer0_outputs(5684)) or (layer0_outputs(1102)));
    outputs(9804) <= layer0_outputs(5817);
    outputs(9805) <= (layer0_outputs(10178)) and not (layer0_outputs(11370));
    outputs(9806) <= not(layer0_outputs(776)) or (layer0_outputs(11166));
    outputs(9807) <= (layer0_outputs(119)) xor (layer0_outputs(6250));
    outputs(9808) <= (layer0_outputs(10494)) xor (layer0_outputs(10865));
    outputs(9809) <= not((layer0_outputs(8823)) xor (layer0_outputs(3424)));
    outputs(9810) <= not(layer0_outputs(2520)) or (layer0_outputs(10485));
    outputs(9811) <= (layer0_outputs(4317)) and (layer0_outputs(8722));
    outputs(9812) <= (layer0_outputs(8461)) and not (layer0_outputs(2740));
    outputs(9813) <= (layer0_outputs(7092)) and (layer0_outputs(7337));
    outputs(9814) <= layer0_outputs(10062);
    outputs(9815) <= not(layer0_outputs(4356)) or (layer0_outputs(1628));
    outputs(9816) <= layer0_outputs(11441);
    outputs(9817) <= not((layer0_outputs(4998)) or (layer0_outputs(2833)));
    outputs(9818) <= not(layer0_outputs(2917)) or (layer0_outputs(7459));
    outputs(9819) <= not((layer0_outputs(1509)) and (layer0_outputs(8202)));
    outputs(9820) <= not((layer0_outputs(11342)) xor (layer0_outputs(3829)));
    outputs(9821) <= not(layer0_outputs(4369));
    outputs(9822) <= not(layer0_outputs(11090));
    outputs(9823) <= (layer0_outputs(54)) and (layer0_outputs(2224));
    outputs(9824) <= not(layer0_outputs(1609));
    outputs(9825) <= not(layer0_outputs(6246));
    outputs(9826) <= not((layer0_outputs(584)) or (layer0_outputs(5331)));
    outputs(9827) <= not((layer0_outputs(5168)) xor (layer0_outputs(9686)));
    outputs(9828) <= (layer0_outputs(2458)) and (layer0_outputs(1371));
    outputs(9829) <= not(layer0_outputs(12328));
    outputs(9830) <= (layer0_outputs(2214)) and not (layer0_outputs(3883));
    outputs(9831) <= not(layer0_outputs(5447));
    outputs(9832) <= (layer0_outputs(11496)) xor (layer0_outputs(9515));
    outputs(9833) <= layer0_outputs(5745);
    outputs(9834) <= layer0_outputs(6264);
    outputs(9835) <= (layer0_outputs(10979)) xor (layer0_outputs(938));
    outputs(9836) <= not(layer0_outputs(10600)) or (layer0_outputs(11943));
    outputs(9837) <= not((layer0_outputs(1730)) or (layer0_outputs(5427)));
    outputs(9838) <= not(layer0_outputs(2506));
    outputs(9839) <= (layer0_outputs(1742)) and not (layer0_outputs(7591));
    outputs(9840) <= not((layer0_outputs(9366)) or (layer0_outputs(2189)));
    outputs(9841) <= not((layer0_outputs(1277)) or (layer0_outputs(7394)));
    outputs(9842) <= layer0_outputs(1188);
    outputs(9843) <= (layer0_outputs(3437)) and (layer0_outputs(8597));
    outputs(9844) <= layer0_outputs(12350);
    outputs(9845) <= not(layer0_outputs(8267));
    outputs(9846) <= (layer0_outputs(6320)) xor (layer0_outputs(8328));
    outputs(9847) <= not(layer0_outputs(5428));
    outputs(9848) <= (layer0_outputs(1195)) and not (layer0_outputs(7223));
    outputs(9849) <= not((layer0_outputs(2642)) xor (layer0_outputs(8603)));
    outputs(9850) <= not((layer0_outputs(12257)) or (layer0_outputs(4200)));
    outputs(9851) <= not(layer0_outputs(5137));
    outputs(9852) <= not(layer0_outputs(9877));
    outputs(9853) <= (layer0_outputs(11753)) xor (layer0_outputs(10693));
    outputs(9854) <= (layer0_outputs(5625)) and (layer0_outputs(2863));
    outputs(9855) <= (layer0_outputs(4275)) xor (layer0_outputs(10750));
    outputs(9856) <= not((layer0_outputs(4755)) or (layer0_outputs(2677)));
    outputs(9857) <= layer0_outputs(1614);
    outputs(9858) <= (layer0_outputs(1470)) and not (layer0_outputs(8883));
    outputs(9859) <= (layer0_outputs(4081)) and not (layer0_outputs(2668));
    outputs(9860) <= not((layer0_outputs(3672)) xor (layer0_outputs(3438)));
    outputs(9861) <= layer0_outputs(11806);
    outputs(9862) <= (layer0_outputs(7356)) and not (layer0_outputs(9489));
    outputs(9863) <= not(layer0_outputs(1318));
    outputs(9864) <= layer0_outputs(4617);
    outputs(9865) <= not((layer0_outputs(12373)) xor (layer0_outputs(3652)));
    outputs(9866) <= (layer0_outputs(9642)) xor (layer0_outputs(7374));
    outputs(9867) <= layer0_outputs(11084);
    outputs(9868) <= not(layer0_outputs(9734));
    outputs(9869) <= layer0_outputs(1685);
    outputs(9870) <= layer0_outputs(6541);
    outputs(9871) <= layer0_outputs(2807);
    outputs(9872) <= layer0_outputs(2346);
    outputs(9873) <= not((layer0_outputs(1709)) and (layer0_outputs(7136)));
    outputs(9874) <= (layer0_outputs(1155)) and not (layer0_outputs(11059));
    outputs(9875) <= not((layer0_outputs(9591)) or (layer0_outputs(4721)));
    outputs(9876) <= layer0_outputs(7449);
    outputs(9877) <= not((layer0_outputs(7921)) and (layer0_outputs(3699)));
    outputs(9878) <= (layer0_outputs(6691)) and (layer0_outputs(2085));
    outputs(9879) <= not(layer0_outputs(3227));
    outputs(9880) <= (layer0_outputs(8013)) and not (layer0_outputs(3722));
    outputs(9881) <= not(layer0_outputs(6306));
    outputs(9882) <= (layer0_outputs(2798)) and not (layer0_outputs(9941));
    outputs(9883) <= (layer0_outputs(12308)) xor (layer0_outputs(12529));
    outputs(9884) <= (layer0_outputs(1224)) xor (layer0_outputs(4218));
    outputs(9885) <= layer0_outputs(9675);
    outputs(9886) <= not(layer0_outputs(12681));
    outputs(9887) <= (layer0_outputs(2308)) and (layer0_outputs(12335));
    outputs(9888) <= layer0_outputs(7663);
    outputs(9889) <= not((layer0_outputs(6985)) xor (layer0_outputs(47)));
    outputs(9890) <= '1';
    outputs(9891) <= (layer0_outputs(6348)) and (layer0_outputs(6418));
    outputs(9892) <= (layer0_outputs(12709)) xor (layer0_outputs(3635));
    outputs(9893) <= (layer0_outputs(273)) or (layer0_outputs(191));
    outputs(9894) <= layer0_outputs(2419);
    outputs(9895) <= layer0_outputs(12385);
    outputs(9896) <= not(layer0_outputs(5872));
    outputs(9897) <= (layer0_outputs(2957)) and not (layer0_outputs(4732));
    outputs(9898) <= layer0_outputs(12558);
    outputs(9899) <= (layer0_outputs(11709)) and not (layer0_outputs(2935));
    outputs(9900) <= (layer0_outputs(12669)) xor (layer0_outputs(978));
    outputs(9901) <= layer0_outputs(3242);
    outputs(9902) <= not((layer0_outputs(5378)) xor (layer0_outputs(10812)));
    outputs(9903) <= (layer0_outputs(1771)) and (layer0_outputs(10906));
    outputs(9904) <= not((layer0_outputs(10593)) xor (layer0_outputs(4580)));
    outputs(9905) <= not(layer0_outputs(1176));
    outputs(9906) <= not((layer0_outputs(3383)) xor (layer0_outputs(1212)));
    outputs(9907) <= not(layer0_outputs(9667));
    outputs(9908) <= (layer0_outputs(3923)) xor (layer0_outputs(3158));
    outputs(9909) <= (layer0_outputs(11345)) and not (layer0_outputs(8795));
    outputs(9910) <= not(layer0_outputs(1954));
    outputs(9911) <= not(layer0_outputs(765));
    outputs(9912) <= '1';
    outputs(9913) <= layer0_outputs(6516);
    outputs(9914) <= layer0_outputs(10959);
    outputs(9915) <= layer0_outputs(2686);
    outputs(9916) <= not((layer0_outputs(10063)) xor (layer0_outputs(7933)));
    outputs(9917) <= (layer0_outputs(10717)) and (layer0_outputs(10922));
    outputs(9918) <= layer0_outputs(11451);
    outputs(9919) <= layer0_outputs(10484);
    outputs(9920) <= not(layer0_outputs(2658));
    outputs(9921) <= (layer0_outputs(5722)) and not (layer0_outputs(5064));
    outputs(9922) <= layer0_outputs(2265);
    outputs(9923) <= not((layer0_outputs(3752)) xor (layer0_outputs(6852)));
    outputs(9924) <= not((layer0_outputs(1570)) or (layer0_outputs(8800)));
    outputs(9925) <= layer0_outputs(1926);
    outputs(9926) <= (layer0_outputs(6672)) xor (layer0_outputs(11464));
    outputs(9927) <= not(layer0_outputs(12225)) or (layer0_outputs(2198));
    outputs(9928) <= (layer0_outputs(10048)) and not (layer0_outputs(3324));
    outputs(9929) <= layer0_outputs(3380);
    outputs(9930) <= layer0_outputs(3822);
    outputs(9931) <= not((layer0_outputs(9638)) xor (layer0_outputs(3059)));
    outputs(9932) <= (layer0_outputs(6993)) xor (layer0_outputs(970));
    outputs(9933) <= not((layer0_outputs(12138)) xor (layer0_outputs(12061)));
    outputs(9934) <= not(layer0_outputs(6808));
    outputs(9935) <= not((layer0_outputs(2133)) xor (layer0_outputs(2469)));
    outputs(9936) <= (layer0_outputs(5903)) and not (layer0_outputs(8705));
    outputs(9937) <= not((layer0_outputs(11490)) or (layer0_outputs(4280)));
    outputs(9938) <= not((layer0_outputs(6502)) xor (layer0_outputs(8457)));
    outputs(9939) <= not((layer0_outputs(2755)) or (layer0_outputs(10518)));
    outputs(9940) <= not((layer0_outputs(10187)) xor (layer0_outputs(2599)));
    outputs(9941) <= not(layer0_outputs(10021));
    outputs(9942) <= (layer0_outputs(12419)) and not (layer0_outputs(9559));
    outputs(9943) <= not((layer0_outputs(1635)) or (layer0_outputs(7024)));
    outputs(9944) <= '1';
    outputs(9945) <= not(layer0_outputs(10470));
    outputs(9946) <= (layer0_outputs(12193)) and (layer0_outputs(721));
    outputs(9947) <= not((layer0_outputs(4770)) xor (layer0_outputs(5003)));
    outputs(9948) <= not((layer0_outputs(12744)) xor (layer0_outputs(9981)));
    outputs(9949) <= not(layer0_outputs(11274));
    outputs(9950) <= (layer0_outputs(10627)) xor (layer0_outputs(10341));
    outputs(9951) <= not((layer0_outputs(10703)) xor (layer0_outputs(604)));
    outputs(9952) <= not(layer0_outputs(1896));
    outputs(9953) <= not(layer0_outputs(689));
    outputs(9954) <= layer0_outputs(12312);
    outputs(9955) <= not(layer0_outputs(258));
    outputs(9956) <= layer0_outputs(2489);
    outputs(9957) <= not((layer0_outputs(267)) xor (layer0_outputs(8839)));
    outputs(9958) <= layer0_outputs(12737);
    outputs(9959) <= layer0_outputs(9064);
    outputs(9960) <= (layer0_outputs(3806)) and not (layer0_outputs(955));
    outputs(9961) <= (layer0_outputs(1305)) or (layer0_outputs(3371));
    outputs(9962) <= not(layer0_outputs(659)) or (layer0_outputs(1311));
    outputs(9963) <= (layer0_outputs(4618)) and (layer0_outputs(12152));
    outputs(9964) <= layer0_outputs(1464);
    outputs(9965) <= not((layer0_outputs(4727)) xor (layer0_outputs(9048)));
    outputs(9966) <= (layer0_outputs(2985)) xor (layer0_outputs(8453));
    outputs(9967) <= (layer0_outputs(6865)) and not (layer0_outputs(1226));
    outputs(9968) <= not(layer0_outputs(2920));
    outputs(9969) <= (layer0_outputs(12120)) or (layer0_outputs(10646));
    outputs(9970) <= not(layer0_outputs(10100));
    outputs(9971) <= layer0_outputs(10410);
    outputs(9972) <= not(layer0_outputs(2929));
    outputs(9973) <= not(layer0_outputs(4312));
    outputs(9974) <= not(layer0_outputs(7060));
    outputs(9975) <= not(layer0_outputs(368)) or (layer0_outputs(8799));
    outputs(9976) <= layer0_outputs(7715);
    outputs(9977) <= not((layer0_outputs(7079)) xor (layer0_outputs(6850)));
    outputs(9978) <= (layer0_outputs(11277)) and (layer0_outputs(7736));
    outputs(9979) <= (layer0_outputs(6538)) xor (layer0_outputs(6618));
    outputs(9980) <= (layer0_outputs(8428)) xor (layer0_outputs(762));
    outputs(9981) <= not(layer0_outputs(7992));
    outputs(9982) <= not((layer0_outputs(7439)) or (layer0_outputs(1176)));
    outputs(9983) <= layer0_outputs(870);
    outputs(9984) <= not((layer0_outputs(10860)) xor (layer0_outputs(4193)));
    outputs(9985) <= not(layer0_outputs(7387));
    outputs(9986) <= not(layer0_outputs(9692));
    outputs(9987) <= (layer0_outputs(372)) xor (layer0_outputs(178));
    outputs(9988) <= layer0_outputs(875);
    outputs(9989) <= (layer0_outputs(4493)) and not (layer0_outputs(11977));
    outputs(9990) <= not((layer0_outputs(4066)) and (layer0_outputs(7418)));
    outputs(9991) <= layer0_outputs(5088);
    outputs(9992) <= '0';
    outputs(9993) <= (layer0_outputs(11801)) xor (layer0_outputs(10747));
    outputs(9994) <= not((layer0_outputs(6075)) or (layer0_outputs(11407)));
    outputs(9995) <= not((layer0_outputs(3348)) xor (layer0_outputs(4686)));
    outputs(9996) <= not(layer0_outputs(4560));
    outputs(9997) <= (layer0_outputs(1288)) xor (layer0_outputs(7238));
    outputs(9998) <= not((layer0_outputs(8501)) xor (layer0_outputs(343)));
    outputs(9999) <= (layer0_outputs(7344)) and not (layer0_outputs(6632));
    outputs(10000) <= not((layer0_outputs(7560)) xor (layer0_outputs(5668)));
    outputs(10001) <= layer0_outputs(181);
    outputs(10002) <= layer0_outputs(5044);
    outputs(10003) <= not(layer0_outputs(3274));
    outputs(10004) <= not((layer0_outputs(4576)) xor (layer0_outputs(2850)));
    outputs(10005) <= not(layer0_outputs(9786));
    outputs(10006) <= (layer0_outputs(9966)) and (layer0_outputs(4205));
    outputs(10007) <= not(layer0_outputs(11727));
    outputs(10008) <= layer0_outputs(9573);
    outputs(10009) <= (layer0_outputs(1088)) and not (layer0_outputs(8877));
    outputs(10010) <= not(layer0_outputs(1970));
    outputs(10011) <= not(layer0_outputs(9138));
    outputs(10012) <= not((layer0_outputs(5436)) xor (layer0_outputs(11166)));
    outputs(10013) <= not((layer0_outputs(11835)) xor (layer0_outputs(12291)));
    outputs(10014) <= (layer0_outputs(12495)) xor (layer0_outputs(1396));
    outputs(10015) <= layer0_outputs(9570);
    outputs(10016) <= layer0_outputs(1642);
    outputs(10017) <= not(layer0_outputs(5883));
    outputs(10018) <= not(layer0_outputs(10315));
    outputs(10019) <= not(layer0_outputs(9844));
    outputs(10020) <= layer0_outputs(10662);
    outputs(10021) <= layer0_outputs(1305);
    outputs(10022) <= not(layer0_outputs(11546));
    outputs(10023) <= (layer0_outputs(8123)) xor (layer0_outputs(979));
    outputs(10024) <= not(layer0_outputs(3145));
    outputs(10025) <= layer0_outputs(9621);
    outputs(10026) <= not(layer0_outputs(1217)) or (layer0_outputs(12772));
    outputs(10027) <= not(layer0_outputs(9887));
    outputs(10028) <= not((layer0_outputs(2437)) and (layer0_outputs(2299)));
    outputs(10029) <= not((layer0_outputs(3782)) xor (layer0_outputs(1512)));
    outputs(10030) <= layer0_outputs(4388);
    outputs(10031) <= (layer0_outputs(1535)) and not (layer0_outputs(7903));
    outputs(10032) <= '0';
    outputs(10033) <= (layer0_outputs(8147)) or (layer0_outputs(12316));
    outputs(10034) <= layer0_outputs(8450);
    outputs(10035) <= layer0_outputs(10762);
    outputs(10036) <= layer0_outputs(5670);
    outputs(10037) <= not((layer0_outputs(5291)) xor (layer0_outputs(12589)));
    outputs(10038) <= (layer0_outputs(1664)) xor (layer0_outputs(2773));
    outputs(10039) <= not(layer0_outputs(8002));
    outputs(10040) <= layer0_outputs(9202);
    outputs(10041) <= not((layer0_outputs(6764)) xor (layer0_outputs(11654)));
    outputs(10042) <= layer0_outputs(4140);
    outputs(10043) <= layer0_outputs(11055);
    outputs(10044) <= not(layer0_outputs(592));
    outputs(10045) <= not((layer0_outputs(1312)) xor (layer0_outputs(1456)));
    outputs(10046) <= (layer0_outputs(5847)) and (layer0_outputs(8612));
    outputs(10047) <= layer0_outputs(5885);
    outputs(10048) <= not(layer0_outputs(12512));
    outputs(10049) <= (layer0_outputs(6023)) xor (layer0_outputs(6319));
    outputs(10050) <= (layer0_outputs(5100)) or (layer0_outputs(7111));
    outputs(10051) <= layer0_outputs(10941);
    outputs(10052) <= layer0_outputs(2948);
    outputs(10053) <= layer0_outputs(5302);
    outputs(10054) <= not((layer0_outputs(12530)) xor (layer0_outputs(10020)));
    outputs(10055) <= (layer0_outputs(10145)) xor (layer0_outputs(1662));
    outputs(10056) <= not(layer0_outputs(5282));
    outputs(10057) <= not((layer0_outputs(5639)) xor (layer0_outputs(2209)));
    outputs(10058) <= not(layer0_outputs(6208));
    outputs(10059) <= not(layer0_outputs(6681));
    outputs(10060) <= not(layer0_outputs(3086));
    outputs(10061) <= layer0_outputs(893);
    outputs(10062) <= not((layer0_outputs(2047)) or (layer0_outputs(11245)));
    outputs(10063) <= not((layer0_outputs(204)) xor (layer0_outputs(11067)));
    outputs(10064) <= (layer0_outputs(2845)) and (layer0_outputs(723));
    outputs(10065) <= layer0_outputs(5305);
    outputs(10066) <= layer0_outputs(5732);
    outputs(10067) <= (layer0_outputs(5886)) and not (layer0_outputs(2652));
    outputs(10068) <= (layer0_outputs(10770)) and not (layer0_outputs(3912));
    outputs(10069) <= layer0_outputs(12448);
    outputs(10070) <= not(layer0_outputs(490));
    outputs(10071) <= not((layer0_outputs(1678)) xor (layer0_outputs(5083)));
    outputs(10072) <= not((layer0_outputs(2281)) and (layer0_outputs(6825)));
    outputs(10073) <= not((layer0_outputs(7536)) xor (layer0_outputs(10461)));
    outputs(10074) <= layer0_outputs(6040);
    outputs(10075) <= not(layer0_outputs(3309));
    outputs(10076) <= not(layer0_outputs(389));
    outputs(10077) <= layer0_outputs(1020);
    outputs(10078) <= (layer0_outputs(8385)) or (layer0_outputs(11980));
    outputs(10079) <= (layer0_outputs(10793)) xor (layer0_outputs(11532));
    outputs(10080) <= (layer0_outputs(8248)) xor (layer0_outputs(622));
    outputs(10081) <= (layer0_outputs(7692)) and not (layer0_outputs(3224));
    outputs(10082) <= (layer0_outputs(8797)) xor (layer0_outputs(667));
    outputs(10083) <= (layer0_outputs(12733)) xor (layer0_outputs(5642));
    outputs(10084) <= not((layer0_outputs(9004)) xor (layer0_outputs(823)));
    outputs(10085) <= not(layer0_outputs(6518));
    outputs(10086) <= (layer0_outputs(6698)) xor (layer0_outputs(2471));
    outputs(10087) <= not((layer0_outputs(2119)) xor (layer0_outputs(7659)));
    outputs(10088) <= layer0_outputs(5629);
    outputs(10089) <= not(layer0_outputs(3188)) or (layer0_outputs(7235));
    outputs(10090) <= not(layer0_outputs(3777));
    outputs(10091) <= not(layer0_outputs(11165));
    outputs(10092) <= (layer0_outputs(1056)) xor (layer0_outputs(4008));
    outputs(10093) <= not(layer0_outputs(4438));
    outputs(10094) <= not((layer0_outputs(6194)) xor (layer0_outputs(8206)));
    outputs(10095) <= not((layer0_outputs(10065)) or (layer0_outputs(7336)));
    outputs(10096) <= not((layer0_outputs(5942)) xor (layer0_outputs(12461)));
    outputs(10097) <= not(layer0_outputs(7682));
    outputs(10098) <= not(layer0_outputs(6533));
    outputs(10099) <= not((layer0_outputs(4274)) xor (layer0_outputs(7299)));
    outputs(10100) <= layer0_outputs(7855);
    outputs(10101) <= not(layer0_outputs(2425));
    outputs(10102) <= (layer0_outputs(12693)) and not (layer0_outputs(11664));
    outputs(10103) <= (layer0_outputs(6444)) and not (layer0_outputs(8949));
    outputs(10104) <= not(layer0_outputs(3364));
    outputs(10105) <= not(layer0_outputs(7519));
    outputs(10106) <= (layer0_outputs(7576)) xor (layer0_outputs(8941));
    outputs(10107) <= (layer0_outputs(5696)) and not (layer0_outputs(11565));
    outputs(10108) <= not(layer0_outputs(1686));
    outputs(10109) <= not((layer0_outputs(1253)) or (layer0_outputs(10966)));
    outputs(10110) <= layer0_outputs(12233);
    outputs(10111) <= not(layer0_outputs(10303));
    outputs(10112) <= (layer0_outputs(4917)) xor (layer0_outputs(2042));
    outputs(10113) <= not((layer0_outputs(167)) xor (layer0_outputs(9968)));
    outputs(10114) <= (layer0_outputs(2061)) and not (layer0_outputs(3590));
    outputs(10115) <= (layer0_outputs(11328)) and not (layer0_outputs(7570));
    outputs(10116) <= not(layer0_outputs(4425));
    outputs(10117) <= not(layer0_outputs(5633));
    outputs(10118) <= not(layer0_outputs(5365));
    outputs(10119) <= not((layer0_outputs(3050)) or (layer0_outputs(11153)));
    outputs(10120) <= not((layer0_outputs(1194)) or (layer0_outputs(12511)));
    outputs(10121) <= not((layer0_outputs(12537)) xor (layer0_outputs(6920)));
    outputs(10122) <= layer0_outputs(12258);
    outputs(10123) <= not(layer0_outputs(8399));
    outputs(10124) <= not(layer0_outputs(5316));
    outputs(10125) <= not(layer0_outputs(7328));
    outputs(10126) <= not((layer0_outputs(4078)) xor (layer0_outputs(6272)));
    outputs(10127) <= layer0_outputs(8656);
    outputs(10128) <= not(layer0_outputs(7497));
    outputs(10129) <= not((layer0_outputs(9292)) and (layer0_outputs(6033)));
    outputs(10130) <= (layer0_outputs(1976)) and not (layer0_outputs(9235));
    outputs(10131) <= (layer0_outputs(7234)) and not (layer0_outputs(6589));
    outputs(10132) <= not(layer0_outputs(8484));
    outputs(10133) <= layer0_outputs(4379);
    outputs(10134) <= layer0_outputs(6807);
    outputs(10135) <= not(layer0_outputs(7790));
    outputs(10136) <= not((layer0_outputs(4916)) xor (layer0_outputs(9356)));
    outputs(10137) <= (layer0_outputs(6469)) xor (layer0_outputs(1012));
    outputs(10138) <= (layer0_outputs(1579)) and not (layer0_outputs(472));
    outputs(10139) <= not(layer0_outputs(4021));
    outputs(10140) <= layer0_outputs(2822);
    outputs(10141) <= layer0_outputs(2778);
    outputs(10142) <= not(layer0_outputs(2137));
    outputs(10143) <= not((layer0_outputs(2905)) or (layer0_outputs(932)));
    outputs(10144) <= (layer0_outputs(3552)) xor (layer0_outputs(7955));
    outputs(10145) <= not(layer0_outputs(7388));
    outputs(10146) <= not((layer0_outputs(5270)) or (layer0_outputs(9045)));
    outputs(10147) <= not((layer0_outputs(8974)) xor (layer0_outputs(8702)));
    outputs(10148) <= not((layer0_outputs(8467)) xor (layer0_outputs(7837)));
    outputs(10149) <= (layer0_outputs(2533)) xor (layer0_outputs(4315));
    outputs(10150) <= layer0_outputs(742);
    outputs(10151) <= (layer0_outputs(11638)) xor (layer0_outputs(7555));
    outputs(10152) <= not(layer0_outputs(3632));
    outputs(10153) <= not((layer0_outputs(8681)) xor (layer0_outputs(6266)));
    outputs(10154) <= not(layer0_outputs(8217));
    outputs(10155) <= not(layer0_outputs(1290));
    outputs(10156) <= not((layer0_outputs(10539)) xor (layer0_outputs(2395)));
    outputs(10157) <= not(layer0_outputs(7185));
    outputs(10158) <= (layer0_outputs(10256)) and not (layer0_outputs(5155));
    outputs(10159) <= (layer0_outputs(9546)) or (layer0_outputs(12088));
    outputs(10160) <= (layer0_outputs(289)) and (layer0_outputs(5483));
    outputs(10161) <= (layer0_outputs(4278)) and (layer0_outputs(5286));
    outputs(10162) <= layer0_outputs(11396);
    outputs(10163) <= (layer0_outputs(1109)) and not (layer0_outputs(7162));
    outputs(10164) <= (layer0_outputs(3363)) and not (layer0_outputs(11759));
    outputs(10165) <= not(layer0_outputs(6532));
    outputs(10166) <= not(layer0_outputs(2981)) or (layer0_outputs(7058));
    outputs(10167) <= not(layer0_outputs(9237));
    outputs(10168) <= not(layer0_outputs(5582));
    outputs(10169) <= (layer0_outputs(2097)) and not (layer0_outputs(11585));
    outputs(10170) <= not(layer0_outputs(4757)) or (layer0_outputs(2095));
    outputs(10171) <= (layer0_outputs(12354)) and not (layer0_outputs(6889));
    outputs(10172) <= not((layer0_outputs(8427)) xor (layer0_outputs(7757)));
    outputs(10173) <= not(layer0_outputs(8585));
    outputs(10174) <= (layer0_outputs(9039)) xor (layer0_outputs(7847));
    outputs(10175) <= layer0_outputs(2974);
    outputs(10176) <= '1';
    outputs(10177) <= not((layer0_outputs(2942)) xor (layer0_outputs(4878)));
    outputs(10178) <= not((layer0_outputs(7016)) xor (layer0_outputs(12101)));
    outputs(10179) <= not(layer0_outputs(856));
    outputs(10180) <= not(layer0_outputs(12598));
    outputs(10181) <= (layer0_outputs(6064)) and not (layer0_outputs(10781));
    outputs(10182) <= layer0_outputs(2766);
    outputs(10183) <= not((layer0_outputs(7411)) or (layer0_outputs(11941)));
    outputs(10184) <= not(layer0_outputs(8679));
    outputs(10185) <= not(layer0_outputs(9575));
    outputs(10186) <= layer0_outputs(5404);
    outputs(10187) <= not(layer0_outputs(5739));
    outputs(10188) <= not(layer0_outputs(8924));
    outputs(10189) <= (layer0_outputs(2548)) xor (layer0_outputs(313));
    outputs(10190) <= (layer0_outputs(6616)) and not (layer0_outputs(4061));
    outputs(10191) <= (layer0_outputs(8398)) and (layer0_outputs(10850));
    outputs(10192) <= layer0_outputs(4845);
    outputs(10193) <= not(layer0_outputs(1225));
    outputs(10194) <= not(layer0_outputs(6248)) or (layer0_outputs(9852));
    outputs(10195) <= (layer0_outputs(4500)) and (layer0_outputs(6061));
    outputs(10196) <= not(layer0_outputs(1782));
    outputs(10197) <= (layer0_outputs(990)) and not (layer0_outputs(1490));
    outputs(10198) <= layer0_outputs(4508);
    outputs(10199) <= layer0_outputs(12707);
    outputs(10200) <= not(layer0_outputs(4665));
    outputs(10201) <= not(layer0_outputs(10756));
    outputs(10202) <= not((layer0_outputs(8941)) or (layer0_outputs(7621)));
    outputs(10203) <= not((layer0_outputs(6331)) and (layer0_outputs(8518)));
    outputs(10204) <= (layer0_outputs(8419)) xor (layer0_outputs(12474));
    outputs(10205) <= not(layer0_outputs(3203));
    outputs(10206) <= (layer0_outputs(6720)) xor (layer0_outputs(6554));
    outputs(10207) <= (layer0_outputs(2381)) and not (layer0_outputs(2964));
    outputs(10208) <= '0';
    outputs(10209) <= not((layer0_outputs(9720)) or (layer0_outputs(9344)));
    outputs(10210) <= layer0_outputs(1740);
    outputs(10211) <= (layer0_outputs(9572)) xor (layer0_outputs(2874));
    outputs(10212) <= layer0_outputs(11209);
    outputs(10213) <= not((layer0_outputs(10573)) or (layer0_outputs(12546)));
    outputs(10214) <= (layer0_outputs(2410)) and not (layer0_outputs(9238));
    outputs(10215) <= layer0_outputs(2226);
    outputs(10216) <= (layer0_outputs(7156)) xor (layer0_outputs(6848));
    outputs(10217) <= (layer0_outputs(5142)) and (layer0_outputs(3999));
    outputs(10218) <= not((layer0_outputs(294)) xor (layer0_outputs(3546)));
    outputs(10219) <= (layer0_outputs(3656)) and not (layer0_outputs(2635));
    outputs(10220) <= layer0_outputs(10763);
    outputs(10221) <= (layer0_outputs(11266)) and (layer0_outputs(7825));
    outputs(10222) <= not(layer0_outputs(7031));
    outputs(10223) <= (layer0_outputs(8129)) and not (layer0_outputs(10658));
    outputs(10224) <= layer0_outputs(6290);
    outputs(10225) <= not(layer0_outputs(4457));
    outputs(10226) <= (layer0_outputs(5917)) and (layer0_outputs(2912));
    outputs(10227) <= layer0_outputs(3248);
    outputs(10228) <= (layer0_outputs(11100)) and not (layer0_outputs(38));
    outputs(10229) <= not((layer0_outputs(11731)) xor (layer0_outputs(3852)));
    outputs(10230) <= (layer0_outputs(9454)) xor (layer0_outputs(3992));
    outputs(10231) <= not((layer0_outputs(4115)) xor (layer0_outputs(9585)));
    outputs(10232) <= (layer0_outputs(9112)) xor (layer0_outputs(1462));
    outputs(10233) <= (layer0_outputs(8413)) and not (layer0_outputs(3293));
    outputs(10234) <= (layer0_outputs(11357)) and not (layer0_outputs(6560));
    outputs(10235) <= not((layer0_outputs(9453)) xor (layer0_outputs(12465)));
    outputs(10236) <= not((layer0_outputs(6293)) xor (layer0_outputs(3283)));
    outputs(10237) <= (layer0_outputs(1050)) and not (layer0_outputs(4172));
    outputs(10238) <= layer0_outputs(10737);
    outputs(10239) <= (layer0_outputs(8779)) and (layer0_outputs(6554));
    outputs(10240) <= (layer0_outputs(6833)) xor (layer0_outputs(9672));
    outputs(10241) <= (layer0_outputs(3742)) xor (layer0_outputs(10973));
    outputs(10242) <= not((layer0_outputs(1450)) xor (layer0_outputs(3522)));
    outputs(10243) <= layer0_outputs(12211);
    outputs(10244) <= layer0_outputs(6347);
    outputs(10245) <= (layer0_outputs(9168)) and not (layer0_outputs(10871));
    outputs(10246) <= not(layer0_outputs(9053));
    outputs(10247) <= layer0_outputs(6386);
    outputs(10248) <= not(layer0_outputs(7854)) or (layer0_outputs(52));
    outputs(10249) <= not(layer0_outputs(3783));
    outputs(10250) <= (layer0_outputs(8271)) and not (layer0_outputs(11388));
    outputs(10251) <= layer0_outputs(8673);
    outputs(10252) <= not(layer0_outputs(1677));
    outputs(10253) <= layer0_outputs(168);
    outputs(10254) <= not(layer0_outputs(11906));
    outputs(10255) <= not((layer0_outputs(1237)) or (layer0_outputs(418)));
    outputs(10256) <= not(layer0_outputs(9296));
    outputs(10257) <= not((layer0_outputs(670)) and (layer0_outputs(7906)));
    outputs(10258) <= not(layer0_outputs(9502));
    outputs(10259) <= not((layer0_outputs(590)) xor (layer0_outputs(8061)));
    outputs(10260) <= not((layer0_outputs(3507)) xor (layer0_outputs(11476)));
    outputs(10261) <= not(layer0_outputs(1676));
    outputs(10262) <= (layer0_outputs(1915)) xor (layer0_outputs(11627));
    outputs(10263) <= (layer0_outputs(3296)) xor (layer0_outputs(4341));
    outputs(10264) <= not(layer0_outputs(11922));
    outputs(10265) <= not((layer0_outputs(358)) xor (layer0_outputs(7857)));
    outputs(10266) <= not((layer0_outputs(7238)) xor (layer0_outputs(5656)));
    outputs(10267) <= not(layer0_outputs(10558)) or (layer0_outputs(2355));
    outputs(10268) <= (layer0_outputs(7047)) xor (layer0_outputs(4997));
    outputs(10269) <= not((layer0_outputs(10509)) and (layer0_outputs(8243)));
    outputs(10270) <= not(layer0_outputs(840));
    outputs(10271) <= not(layer0_outputs(8421));
    outputs(10272) <= not(layer0_outputs(11779));
    outputs(10273) <= not((layer0_outputs(5102)) xor (layer0_outputs(3402)));
    outputs(10274) <= (layer0_outputs(6082)) and not (layer0_outputs(1011));
    outputs(10275) <= not(layer0_outputs(5347));
    outputs(10276) <= (layer0_outputs(3644)) xor (layer0_outputs(2665));
    outputs(10277) <= not((layer0_outputs(11148)) xor (layer0_outputs(3600)));
    outputs(10278) <= layer0_outputs(5812);
    outputs(10279) <= not((layer0_outputs(252)) xor (layer0_outputs(11794)));
    outputs(10280) <= layer0_outputs(5466);
    outputs(10281) <= (layer0_outputs(5340)) xor (layer0_outputs(11595));
    outputs(10282) <= not((layer0_outputs(5023)) xor (layer0_outputs(4658)));
    outputs(10283) <= (layer0_outputs(9941)) and not (layer0_outputs(124));
    outputs(10284) <= (layer0_outputs(1361)) xor (layer0_outputs(7495));
    outputs(10285) <= layer0_outputs(12728);
    outputs(10286) <= not(layer0_outputs(3137));
    outputs(10287) <= not(layer0_outputs(7782));
    outputs(10288) <= (layer0_outputs(4256)) and not (layer0_outputs(8521));
    outputs(10289) <= not((layer0_outputs(714)) xor (layer0_outputs(11356)));
    outputs(10290) <= not((layer0_outputs(3327)) xor (layer0_outputs(9284)));
    outputs(10291) <= layer0_outputs(5954);
    outputs(10292) <= not(layer0_outputs(12692));
    outputs(10293) <= (layer0_outputs(3643)) and not (layer0_outputs(5364));
    outputs(10294) <= not((layer0_outputs(483)) and (layer0_outputs(12134)));
    outputs(10295) <= not(layer0_outputs(8552));
    outputs(10296) <= (layer0_outputs(1923)) or (layer0_outputs(10467));
    outputs(10297) <= (layer0_outputs(8024)) and (layer0_outputs(2770));
    outputs(10298) <= not(layer0_outputs(29)) or (layer0_outputs(3949));
    outputs(10299) <= (layer0_outputs(4166)) xor (layer0_outputs(2001));
    outputs(10300) <= layer0_outputs(1747);
    outputs(10301) <= (layer0_outputs(12640)) and (layer0_outputs(2522));
    outputs(10302) <= layer0_outputs(11350);
    outputs(10303) <= (layer0_outputs(121)) xor (layer0_outputs(1571));
    outputs(10304) <= not((layer0_outputs(8409)) and (layer0_outputs(747)));
    outputs(10305) <= not(layer0_outputs(11365));
    outputs(10306) <= not(layer0_outputs(3262)) or (layer0_outputs(4816));
    outputs(10307) <= not((layer0_outputs(11037)) or (layer0_outputs(7528)));
    outputs(10308) <= not(layer0_outputs(9438));
    outputs(10309) <= layer0_outputs(2596);
    outputs(10310) <= not((layer0_outputs(7489)) xor (layer0_outputs(8866)));
    outputs(10311) <= (layer0_outputs(6973)) or (layer0_outputs(5905));
    outputs(10312) <= (layer0_outputs(7751)) xor (layer0_outputs(9402));
    outputs(10313) <= not(layer0_outputs(8751)) or (layer0_outputs(8837));
    outputs(10314) <= (layer0_outputs(5961)) xor (layer0_outputs(2861));
    outputs(10315) <= layer0_outputs(612);
    outputs(10316) <= not(layer0_outputs(7663));
    outputs(10317) <= '1';
    outputs(10318) <= (layer0_outputs(7193)) xor (layer0_outputs(5909));
    outputs(10319) <= (layer0_outputs(10078)) xor (layer0_outputs(5047));
    outputs(10320) <= not((layer0_outputs(8639)) xor (layer0_outputs(2458)));
    outputs(10321) <= (layer0_outputs(2117)) xor (layer0_outputs(8640));
    outputs(10322) <= not((layer0_outputs(10617)) xor (layer0_outputs(11842)));
    outputs(10323) <= (layer0_outputs(9218)) or (layer0_outputs(4521));
    outputs(10324) <= not(layer0_outputs(2802)) or (layer0_outputs(12701));
    outputs(10325) <= (layer0_outputs(2299)) xor (layer0_outputs(991));
    outputs(10326) <= not(layer0_outputs(7801));
    outputs(10327) <= (layer0_outputs(5366)) or (layer0_outputs(2010));
    outputs(10328) <= not(layer0_outputs(5474)) or (layer0_outputs(11684));
    outputs(10329) <= layer0_outputs(8383);
    outputs(10330) <= '1';
    outputs(10331) <= layer0_outputs(9061);
    outputs(10332) <= not(layer0_outputs(2756));
    outputs(10333) <= not((layer0_outputs(383)) xor (layer0_outputs(2398)));
    outputs(10334) <= (layer0_outputs(11524)) and not (layer0_outputs(8923));
    outputs(10335) <= layer0_outputs(1821);
    outputs(10336) <= not(layer0_outputs(2738));
    outputs(10337) <= (layer0_outputs(8156)) xor (layer0_outputs(9110));
    outputs(10338) <= not(layer0_outputs(9749));
    outputs(10339) <= not(layer0_outputs(7950)) or (layer0_outputs(3162));
    outputs(10340) <= not(layer0_outputs(7423));
    outputs(10341) <= not((layer0_outputs(10204)) or (layer0_outputs(9898)));
    outputs(10342) <= not((layer0_outputs(11908)) or (layer0_outputs(4196)));
    outputs(10343) <= not((layer0_outputs(1153)) xor (layer0_outputs(7182)));
    outputs(10344) <= not(layer0_outputs(1160)) or (layer0_outputs(3998));
    outputs(10345) <= not((layer0_outputs(831)) xor (layer0_outputs(2176)));
    outputs(10346) <= not((layer0_outputs(10600)) and (layer0_outputs(10666)));
    outputs(10347) <= '0';
    outputs(10348) <= layer0_outputs(7159);
    outputs(10349) <= not(layer0_outputs(10831)) or (layer0_outputs(3709));
    outputs(10350) <= (layer0_outputs(5791)) xor (layer0_outputs(6739));
    outputs(10351) <= layer0_outputs(799);
    outputs(10352) <= not((layer0_outputs(9212)) xor (layer0_outputs(94)));
    outputs(10353) <= (layer0_outputs(2229)) and (layer0_outputs(10441));
    outputs(10354) <= (layer0_outputs(2282)) xor (layer0_outputs(2775));
    outputs(10355) <= (layer0_outputs(6)) xor (layer0_outputs(3638));
    outputs(10356) <= not(layer0_outputs(5466)) or (layer0_outputs(12646));
    outputs(10357) <= layer0_outputs(1322);
    outputs(10358) <= not((layer0_outputs(2666)) or (layer0_outputs(275)));
    outputs(10359) <= (layer0_outputs(4185)) xor (layer0_outputs(729));
    outputs(10360) <= (layer0_outputs(10676)) xor (layer0_outputs(6046));
    outputs(10361) <= not(layer0_outputs(6045)) or (layer0_outputs(11410));
    outputs(10362) <= not((layer0_outputs(279)) xor (layer0_outputs(6800)));
    outputs(10363) <= not(layer0_outputs(509));
    outputs(10364) <= not((layer0_outputs(5351)) and (layer0_outputs(5538)));
    outputs(10365) <= (layer0_outputs(12581)) xor (layer0_outputs(3613));
    outputs(10366) <= (layer0_outputs(8888)) xor (layer0_outputs(2952));
    outputs(10367) <= (layer0_outputs(9757)) xor (layer0_outputs(791));
    outputs(10368) <= (layer0_outputs(6710)) xor (layer0_outputs(10397));
    outputs(10369) <= layer0_outputs(5958);
    outputs(10370) <= not((layer0_outputs(2693)) xor (layer0_outputs(2555)));
    outputs(10371) <= (layer0_outputs(11900)) or (layer0_outputs(7653));
    outputs(10372) <= (layer0_outputs(5755)) xor (layer0_outputs(8248));
    outputs(10373) <= layer0_outputs(11102);
    outputs(10374) <= layer0_outputs(10633);
    outputs(10375) <= not((layer0_outputs(6162)) and (layer0_outputs(12788)));
    outputs(10376) <= layer0_outputs(10358);
    outputs(10377) <= (layer0_outputs(2155)) and not (layer0_outputs(3748));
    outputs(10378) <= not(layer0_outputs(9552));
    outputs(10379) <= not((layer0_outputs(9153)) xor (layer0_outputs(1296)));
    outputs(10380) <= (layer0_outputs(11068)) xor (layer0_outputs(8775));
    outputs(10381) <= not((layer0_outputs(9503)) or (layer0_outputs(11513)));
    outputs(10382) <= not((layer0_outputs(11289)) or (layer0_outputs(391)));
    outputs(10383) <= layer0_outputs(3040);
    outputs(10384) <= (layer0_outputs(9240)) xor (layer0_outputs(7028));
    outputs(10385) <= (layer0_outputs(8337)) and not (layer0_outputs(9753));
    outputs(10386) <= layer0_outputs(760);
    outputs(10387) <= not((layer0_outputs(7656)) and (layer0_outputs(7448)));
    outputs(10388) <= (layer0_outputs(4273)) and not (layer0_outputs(6030));
    outputs(10389) <= not(layer0_outputs(1856));
    outputs(10390) <= not(layer0_outputs(11510));
    outputs(10391) <= (layer0_outputs(809)) and not (layer0_outputs(11495));
    outputs(10392) <= (layer0_outputs(3579)) xor (layer0_outputs(11246));
    outputs(10393) <= (layer0_outputs(153)) xor (layer0_outputs(1777));
    outputs(10394) <= not((layer0_outputs(5755)) xor (layer0_outputs(827)));
    outputs(10395) <= (layer0_outputs(2730)) or (layer0_outputs(5392));
    outputs(10396) <= layer0_outputs(8852);
    outputs(10397) <= (layer0_outputs(10985)) xor (layer0_outputs(1488));
    outputs(10398) <= layer0_outputs(9169);
    outputs(10399) <= (layer0_outputs(7774)) xor (layer0_outputs(11177));
    outputs(10400) <= layer0_outputs(3902);
    outputs(10401) <= layer0_outputs(1531);
    outputs(10402) <= (layer0_outputs(9647)) or (layer0_outputs(4649));
    outputs(10403) <= layer0_outputs(465);
    outputs(10404) <= not((layer0_outputs(2861)) xor (layer0_outputs(11430)));
    outputs(10405) <= not((layer0_outputs(2586)) and (layer0_outputs(12037)));
    outputs(10406) <= not(layer0_outputs(5352)) or (layer0_outputs(7616));
    outputs(10407) <= not((layer0_outputs(10609)) or (layer0_outputs(6175)));
    outputs(10408) <= (layer0_outputs(2560)) and (layer0_outputs(1313));
    outputs(10409) <= not((layer0_outputs(11965)) xor (layer0_outputs(6558)));
    outputs(10410) <= not(layer0_outputs(8831)) or (layer0_outputs(2581));
    outputs(10411) <= not(layer0_outputs(10831));
    outputs(10412) <= (layer0_outputs(6518)) or (layer0_outputs(6000));
    outputs(10413) <= not(layer0_outputs(3390)) or (layer0_outputs(10182));
    outputs(10414) <= (layer0_outputs(6234)) xor (layer0_outputs(3715));
    outputs(10415) <= not(layer0_outputs(188));
    outputs(10416) <= '1';
    outputs(10417) <= layer0_outputs(10401);
    outputs(10418) <= (layer0_outputs(4353)) xor (layer0_outputs(4361));
    outputs(10419) <= layer0_outputs(2476);
    outputs(10420) <= (layer0_outputs(9204)) xor (layer0_outputs(4681));
    outputs(10421) <= (layer0_outputs(1349)) xor (layer0_outputs(2360));
    outputs(10422) <= layer0_outputs(6229);
    outputs(10423) <= not(layer0_outputs(9780)) or (layer0_outputs(9607));
    outputs(10424) <= (layer0_outputs(12232)) or (layer0_outputs(7170));
    outputs(10425) <= layer0_outputs(10389);
    outputs(10426) <= (layer0_outputs(2124)) xor (layer0_outputs(2435));
    outputs(10427) <= (layer0_outputs(9840)) and not (layer0_outputs(2310));
    outputs(10428) <= not(layer0_outputs(8013));
    outputs(10429) <= layer0_outputs(8472);
    outputs(10430) <= not(layer0_outputs(7103));
    outputs(10431) <= not((layer0_outputs(3384)) xor (layer0_outputs(10123)));
    outputs(10432) <= (layer0_outputs(9044)) and not (layer0_outputs(12087));
    outputs(10433) <= layer0_outputs(1384);
    outputs(10434) <= not(layer0_outputs(11001)) or (layer0_outputs(3124));
    outputs(10435) <= (layer0_outputs(3690)) xor (layer0_outputs(5957));
    outputs(10436) <= '1';
    outputs(10437) <= not((layer0_outputs(5680)) xor (layer0_outputs(1671)));
    outputs(10438) <= not(layer0_outputs(819)) or (layer0_outputs(7053));
    outputs(10439) <= not((layer0_outputs(3190)) and (layer0_outputs(3689)));
    outputs(10440) <= not((layer0_outputs(4081)) and (layer0_outputs(8538)));
    outputs(10441) <= (layer0_outputs(9847)) xor (layer0_outputs(5682));
    outputs(10442) <= not(layer0_outputs(1602));
    outputs(10443) <= not((layer0_outputs(10576)) xor (layer0_outputs(1699)));
    outputs(10444) <= layer0_outputs(2818);
    outputs(10445) <= not(layer0_outputs(3515));
    outputs(10446) <= (layer0_outputs(8193)) xor (layer0_outputs(10476));
    outputs(10447) <= (layer0_outputs(10890)) or (layer0_outputs(11173));
    outputs(10448) <= layer0_outputs(4826);
    outputs(10449) <= layer0_outputs(2322);
    outputs(10450) <= not((layer0_outputs(11880)) xor (layer0_outputs(5617)));
    outputs(10451) <= not(layer0_outputs(10483));
    outputs(10452) <= not(layer0_outputs(6876));
    outputs(10453) <= (layer0_outputs(5990)) xor (layer0_outputs(6452));
    outputs(10454) <= layer0_outputs(1752);
    outputs(10455) <= not(layer0_outputs(3504));
    outputs(10456) <= '1';
    outputs(10457) <= not((layer0_outputs(11877)) or (layer0_outputs(244)));
    outputs(10458) <= not(layer0_outputs(10319));
    outputs(10459) <= (layer0_outputs(7747)) and not (layer0_outputs(6179));
    outputs(10460) <= (layer0_outputs(7511)) and not (layer0_outputs(8764));
    outputs(10461) <= not(layer0_outputs(3491)) or (layer0_outputs(3161));
    outputs(10462) <= (layer0_outputs(4769)) xor (layer0_outputs(5781));
    outputs(10463) <= (layer0_outputs(530)) xor (layer0_outputs(12735));
    outputs(10464) <= layer0_outputs(11989);
    outputs(10465) <= layer0_outputs(3591);
    outputs(10466) <= (layer0_outputs(1092)) and not (layer0_outputs(11374));
    outputs(10467) <= layer0_outputs(3673);
    outputs(10468) <= not((layer0_outputs(143)) xor (layer0_outputs(5663)));
    outputs(10469) <= not(layer0_outputs(11551)) or (layer0_outputs(1066));
    outputs(10470) <= (layer0_outputs(12252)) and not (layer0_outputs(7987));
    outputs(10471) <= not((layer0_outputs(10095)) and (layer0_outputs(2186)));
    outputs(10472) <= layer0_outputs(9724);
    outputs(10473) <= not(layer0_outputs(80));
    outputs(10474) <= not(layer0_outputs(3053)) or (layer0_outputs(3340));
    outputs(10475) <= not(layer0_outputs(5947)) or (layer0_outputs(6587));
    outputs(10476) <= layer0_outputs(4156);
    outputs(10477) <= layer0_outputs(11351);
    outputs(10478) <= (layer0_outputs(9343)) and (layer0_outputs(11413));
    outputs(10479) <= not((layer0_outputs(8569)) or (layer0_outputs(2848)));
    outputs(10480) <= not(layer0_outputs(10645));
    outputs(10481) <= (layer0_outputs(2936)) and not (layer0_outputs(1308));
    outputs(10482) <= layer0_outputs(7222);
    outputs(10483) <= layer0_outputs(3476);
    outputs(10484) <= layer0_outputs(4234);
    outputs(10485) <= (layer0_outputs(822)) xor (layer0_outputs(946));
    outputs(10486) <= layer0_outputs(904);
    outputs(10487) <= not(layer0_outputs(7165));
    outputs(10488) <= not(layer0_outputs(9131));
    outputs(10489) <= not((layer0_outputs(10037)) xor (layer0_outputs(9183)));
    outputs(10490) <= not((layer0_outputs(10595)) xor (layer0_outputs(11275)));
    outputs(10491) <= layer0_outputs(1776);
    outputs(10492) <= (layer0_outputs(816)) xor (layer0_outputs(11819));
    outputs(10493) <= not(layer0_outputs(2100)) or (layer0_outputs(2066));
    outputs(10494) <= (layer0_outputs(6754)) and (layer0_outputs(10742));
    outputs(10495) <= (layer0_outputs(5197)) xor (layer0_outputs(1515));
    outputs(10496) <= not(layer0_outputs(2751)) or (layer0_outputs(7097));
    outputs(10497) <= (layer0_outputs(1868)) and not (layer0_outputs(8732));
    outputs(10498) <= not(layer0_outputs(5266));
    outputs(10499) <= (layer0_outputs(1643)) xor (layer0_outputs(5052));
    outputs(10500) <= (layer0_outputs(4402)) and not (layer0_outputs(8061));
    outputs(10501) <= (layer0_outputs(9855)) or (layer0_outputs(10060));
    outputs(10502) <= (layer0_outputs(4114)) and not (layer0_outputs(976));
    outputs(10503) <= not(layer0_outputs(5875));
    outputs(10504) <= not(layer0_outputs(9151));
    outputs(10505) <= not((layer0_outputs(8678)) and (layer0_outputs(9586)));
    outputs(10506) <= not((layer0_outputs(12269)) and (layer0_outputs(8520)));
    outputs(10507) <= not(layer0_outputs(7937)) or (layer0_outputs(7782));
    outputs(10508) <= not(layer0_outputs(4564));
    outputs(10509) <= not((layer0_outputs(9917)) xor (layer0_outputs(1513)));
    outputs(10510) <= layer0_outputs(6579);
    outputs(10511) <= layer0_outputs(11888);
    outputs(10512) <= layer0_outputs(7020);
    outputs(10513) <= not(layer0_outputs(9371));
    outputs(10514) <= not(layer0_outputs(5914));
    outputs(10515) <= (layer0_outputs(11569)) xor (layer0_outputs(2016));
    outputs(10516) <= '1';
    outputs(10517) <= not(layer0_outputs(7134)) or (layer0_outputs(9348));
    outputs(10518) <= not(layer0_outputs(9276));
    outputs(10519) <= (layer0_outputs(2211)) and (layer0_outputs(9929));
    outputs(10520) <= not(layer0_outputs(8720)) or (layer0_outputs(6323));
    outputs(10521) <= not(layer0_outputs(8464));
    outputs(10522) <= not((layer0_outputs(1808)) xor (layer0_outputs(9166)));
    outputs(10523) <= layer0_outputs(5070);
    outputs(10524) <= not(layer0_outputs(4785)) or (layer0_outputs(11227));
    outputs(10525) <= not(layer0_outputs(7171));
    outputs(10526) <= layer0_outputs(8641);
    outputs(10527) <= (layer0_outputs(7601)) and not (layer0_outputs(3254));
    outputs(10528) <= layer0_outputs(4745);
    outputs(10529) <= not(layer0_outputs(12545));
    outputs(10530) <= layer0_outputs(2823);
    outputs(10531) <= not((layer0_outputs(1709)) and (layer0_outputs(8315)));
    outputs(10532) <= (layer0_outputs(6848)) and not (layer0_outputs(638));
    outputs(10533) <= (layer0_outputs(379)) and (layer0_outputs(4416));
    outputs(10534) <= (layer0_outputs(927)) xor (layer0_outputs(12078));
    outputs(10535) <= not(layer0_outputs(3394));
    outputs(10536) <= not((layer0_outputs(5737)) xor (layer0_outputs(9893)));
    outputs(10537) <= layer0_outputs(3301);
    outputs(10538) <= layer0_outputs(3374);
    outputs(10539) <= (layer0_outputs(486)) or (layer0_outputs(9658));
    outputs(10540) <= (layer0_outputs(1728)) xor (layer0_outputs(3828));
    outputs(10541) <= (layer0_outputs(12594)) xor (layer0_outputs(1268));
    outputs(10542) <= layer0_outputs(1297);
    outputs(10543) <= '1';
    outputs(10544) <= not(layer0_outputs(9267));
    outputs(10545) <= not(layer0_outputs(6324));
    outputs(10546) <= not(layer0_outputs(12085));
    outputs(10547) <= not(layer0_outputs(6220));
    outputs(10548) <= not(layer0_outputs(11723));
    outputs(10549) <= (layer0_outputs(217)) and not (layer0_outputs(12002));
    outputs(10550) <= not((layer0_outputs(2882)) xor (layer0_outputs(5372)));
    outputs(10551) <= layer0_outputs(601);
    outputs(10552) <= layer0_outputs(8540);
    outputs(10553) <= not(layer0_outputs(10380));
    outputs(10554) <= not(layer0_outputs(4797));
    outputs(10555) <= layer0_outputs(4021);
    outputs(10556) <= (layer0_outputs(1753)) xor (layer0_outputs(5103));
    outputs(10557) <= not((layer0_outputs(5843)) xor (layer0_outputs(3438)));
    outputs(10558) <= not((layer0_outputs(4518)) xor (layer0_outputs(4254)));
    outputs(10559) <= not(layer0_outputs(11857));
    outputs(10560) <= (layer0_outputs(4610)) xor (layer0_outputs(4484));
    outputs(10561) <= (layer0_outputs(1478)) and (layer0_outputs(108));
    outputs(10562) <= (layer0_outputs(6250)) xor (layer0_outputs(9076));
    outputs(10563) <= not(layer0_outputs(6287)) or (layer0_outputs(10162));
    outputs(10564) <= layer0_outputs(5066);
    outputs(10565) <= not(layer0_outputs(9780));
    outputs(10566) <= not(layer0_outputs(1563));
    outputs(10567) <= (layer0_outputs(491)) xor (layer0_outputs(9796));
    outputs(10568) <= not((layer0_outputs(3037)) xor (layer0_outputs(1916)));
    outputs(10569) <= not((layer0_outputs(4859)) xor (layer0_outputs(4010)));
    outputs(10570) <= (layer0_outputs(10055)) xor (layer0_outputs(9915));
    outputs(10571) <= layer0_outputs(8458);
    outputs(10572) <= layer0_outputs(1116);
    outputs(10573) <= not((layer0_outputs(6282)) xor (layer0_outputs(12282)));
    outputs(10574) <= not((layer0_outputs(459)) or (layer0_outputs(4068)));
    outputs(10575) <= layer0_outputs(5252);
    outputs(10576) <= (layer0_outputs(7884)) xor (layer0_outputs(4456));
    outputs(10577) <= (layer0_outputs(87)) xor (layer0_outputs(5154));
    outputs(10578) <= '1';
    outputs(10579) <= not((layer0_outputs(10195)) xor (layer0_outputs(10382)));
    outputs(10580) <= layer0_outputs(12382);
    outputs(10581) <= layer0_outputs(7906);
    outputs(10582) <= (layer0_outputs(6291)) xor (layer0_outputs(6235));
    outputs(10583) <= not((layer0_outputs(10197)) xor (layer0_outputs(11753)));
    outputs(10584) <= not(layer0_outputs(11521)) or (layer0_outputs(6747));
    outputs(10585) <= (layer0_outputs(7234)) and not (layer0_outputs(10711));
    outputs(10586) <= (layer0_outputs(10212)) and not (layer0_outputs(9355));
    outputs(10587) <= not((layer0_outputs(2600)) or (layer0_outputs(1613)));
    outputs(10588) <= (layer0_outputs(494)) or (layer0_outputs(12408));
    outputs(10589) <= not((layer0_outputs(2427)) xor (layer0_outputs(7889)));
    outputs(10590) <= layer0_outputs(7915);
    outputs(10591) <= (layer0_outputs(1767)) and not (layer0_outputs(6207));
    outputs(10592) <= layer0_outputs(5517);
    outputs(10593) <= (layer0_outputs(6330)) xor (layer0_outputs(12780));
    outputs(10594) <= (layer0_outputs(6463)) or (layer0_outputs(4860));
    outputs(10595) <= layer0_outputs(4001);
    outputs(10596) <= not((layer0_outputs(4685)) xor (layer0_outputs(5258)));
    outputs(10597) <= not((layer0_outputs(44)) xor (layer0_outputs(8111)));
    outputs(10598) <= not(layer0_outputs(7350));
    outputs(10599) <= (layer0_outputs(8419)) xor (layer0_outputs(942));
    outputs(10600) <= layer0_outputs(10095);
    outputs(10601) <= not(layer0_outputs(334));
    outputs(10602) <= layer0_outputs(1605);
    outputs(10603) <= (layer0_outputs(3714)) xor (layer0_outputs(5823));
    outputs(10604) <= (layer0_outputs(9374)) xor (layer0_outputs(6950));
    outputs(10605) <= not((layer0_outputs(644)) and (layer0_outputs(2020)));
    outputs(10606) <= layer0_outputs(4231);
    outputs(10607) <= layer0_outputs(9683);
    outputs(10608) <= not(layer0_outputs(12742));
    outputs(10609) <= not(layer0_outputs(2210));
    outputs(10610) <= (layer0_outputs(11182)) xor (layer0_outputs(5821));
    outputs(10611) <= not(layer0_outputs(303));
    outputs(10612) <= layer0_outputs(7919);
    outputs(10613) <= (layer0_outputs(11200)) and not (layer0_outputs(7518));
    outputs(10614) <= not((layer0_outputs(8728)) or (layer0_outputs(4861)));
    outputs(10615) <= not(layer0_outputs(5074)) or (layer0_outputs(5769));
    outputs(10616) <= not(layer0_outputs(3041));
    outputs(10617) <= not((layer0_outputs(8885)) and (layer0_outputs(9657)));
    outputs(10618) <= not(layer0_outputs(9481));
    outputs(10619) <= not((layer0_outputs(10347)) xor (layer0_outputs(11236)));
    outputs(10620) <= (layer0_outputs(3485)) xor (layer0_outputs(7907));
    outputs(10621) <= layer0_outputs(3775);
    outputs(10622) <= layer0_outputs(197);
    outputs(10623) <= not((layer0_outputs(1433)) xor (layer0_outputs(457)));
    outputs(10624) <= (layer0_outputs(10174)) or (layer0_outputs(6020));
    outputs(10625) <= not((layer0_outputs(11341)) and (layer0_outputs(5543)));
    outputs(10626) <= (layer0_outputs(1456)) xor (layer0_outputs(2307));
    outputs(10627) <= not(layer0_outputs(215));
    outputs(10628) <= layer0_outputs(6313);
    outputs(10629) <= not(layer0_outputs(9263));
    outputs(10630) <= not((layer0_outputs(3787)) xor (layer0_outputs(10074)));
    outputs(10631) <= not(layer0_outputs(2610)) or (layer0_outputs(8951));
    outputs(10632) <= layer0_outputs(9133);
    outputs(10633) <= not(layer0_outputs(9448));
    outputs(10634) <= (layer0_outputs(10788)) and not (layer0_outputs(5170));
    outputs(10635) <= layer0_outputs(1600);
    outputs(10636) <= (layer0_outputs(6465)) xor (layer0_outputs(9497));
    outputs(10637) <= (layer0_outputs(11334)) xor (layer0_outputs(3970));
    outputs(10638) <= (layer0_outputs(3241)) xor (layer0_outputs(10647));
    outputs(10639) <= not((layer0_outputs(9354)) xor (layer0_outputs(1985)));
    outputs(10640) <= not(layer0_outputs(9219)) or (layer0_outputs(9401));
    outputs(10641) <= not((layer0_outputs(8139)) xor (layer0_outputs(8174)));
    outputs(10642) <= not((layer0_outputs(2640)) and (layer0_outputs(10838)));
    outputs(10643) <= (layer0_outputs(3579)) and not (layer0_outputs(10189));
    outputs(10644) <= layer0_outputs(6963);
    outputs(10645) <= (layer0_outputs(9022)) xor (layer0_outputs(6828));
    outputs(10646) <= layer0_outputs(10510);
    outputs(10647) <= not(layer0_outputs(8998)) or (layer0_outputs(3477));
    outputs(10648) <= not((layer0_outputs(10203)) xor (layer0_outputs(4406)));
    outputs(10649) <= (layer0_outputs(1127)) xor (layer0_outputs(1882));
    outputs(10650) <= (layer0_outputs(12133)) or (layer0_outputs(4336));
    outputs(10651) <= not(layer0_outputs(4405)) or (layer0_outputs(4558));
    outputs(10652) <= not(layer0_outputs(4334)) or (layer0_outputs(4299));
    outputs(10653) <= layer0_outputs(2601);
    outputs(10654) <= not((layer0_outputs(7543)) and (layer0_outputs(4200)));
    outputs(10655) <= not((layer0_outputs(3979)) xor (layer0_outputs(802)));
    outputs(10656) <= not(layer0_outputs(11457));
    outputs(10657) <= (layer0_outputs(3996)) xor (layer0_outputs(2069));
    outputs(10658) <= not(layer0_outputs(12113));
    outputs(10659) <= not(layer0_outputs(5875));
    outputs(10660) <= (layer0_outputs(9011)) and not (layer0_outputs(4486));
    outputs(10661) <= (layer0_outputs(11484)) xor (layer0_outputs(1492));
    outputs(10662) <= not(layer0_outputs(6420)) or (layer0_outputs(11432));
    outputs(10663) <= layer0_outputs(12328);
    outputs(10664) <= not((layer0_outputs(5941)) xor (layer0_outputs(9009)));
    outputs(10665) <= layer0_outputs(4210);
    outputs(10666) <= layer0_outputs(11236);
    outputs(10667) <= (layer0_outputs(6770)) and not (layer0_outputs(6375));
    outputs(10668) <= layer0_outputs(5473);
    outputs(10669) <= layer0_outputs(2809);
    outputs(10670) <= layer0_outputs(1448);
    outputs(10671) <= layer0_outputs(7179);
    outputs(10672) <= (layer0_outputs(5717)) xor (layer0_outputs(7926));
    outputs(10673) <= layer0_outputs(5547);
    outputs(10674) <= (layer0_outputs(5053)) and not (layer0_outputs(1884));
    outputs(10675) <= not(layer0_outputs(4428));
    outputs(10676) <= not(layer0_outputs(656)) or (layer0_outputs(4522));
    outputs(10677) <= layer0_outputs(12158);
    outputs(10678) <= (layer0_outputs(11305)) xor (layer0_outputs(2227));
    outputs(10679) <= (layer0_outputs(5400)) and (layer0_outputs(1231));
    outputs(10680) <= (layer0_outputs(5476)) and not (layer0_outputs(1455));
    outputs(10681) <= not(layer0_outputs(1472));
    outputs(10682) <= not(layer0_outputs(8815)) or (layer0_outputs(2147));
    outputs(10683) <= not((layer0_outputs(1889)) xor (layer0_outputs(4726)));
    outputs(10684) <= not(layer0_outputs(6045));
    outputs(10685) <= layer0_outputs(8762);
    outputs(10686) <= layer0_outputs(11082);
    outputs(10687) <= '1';
    outputs(10688) <= not(layer0_outputs(9522)) or (layer0_outputs(2725));
    outputs(10689) <= not(layer0_outputs(6491));
    outputs(10690) <= not(layer0_outputs(7195));
    outputs(10691) <= (layer0_outputs(6759)) xor (layer0_outputs(10886));
    outputs(10692) <= not((layer0_outputs(6320)) xor (layer0_outputs(8777)));
    outputs(10693) <= layer0_outputs(6538);
    outputs(10694) <= not((layer0_outputs(10368)) or (layer0_outputs(546)));
    outputs(10695) <= layer0_outputs(10633);
    outputs(10696) <= layer0_outputs(8993);
    outputs(10697) <= not((layer0_outputs(10131)) xor (layer0_outputs(12011)));
    outputs(10698) <= layer0_outputs(12089);
    outputs(10699) <= (layer0_outputs(5881)) xor (layer0_outputs(1980));
    outputs(10700) <= (layer0_outputs(6279)) xor (layer0_outputs(1080));
    outputs(10701) <= (layer0_outputs(9025)) or (layer0_outputs(119));
    outputs(10702) <= (layer0_outputs(9304)) and not (layer0_outputs(9024));
    outputs(10703) <= (layer0_outputs(3330)) and not (layer0_outputs(8164));
    outputs(10704) <= not((layer0_outputs(3439)) xor (layer0_outputs(8093)));
    outputs(10705) <= not((layer0_outputs(9051)) xor (layer0_outputs(5086)));
    outputs(10706) <= not((layer0_outputs(6028)) xor (layer0_outputs(1856)));
    outputs(10707) <= not(layer0_outputs(9614));
    outputs(10708) <= not(layer0_outputs(12423));
    outputs(10709) <= (layer0_outputs(4144)) and not (layer0_outputs(701));
    outputs(10710) <= layer0_outputs(12093);
    outputs(10711) <= (layer0_outputs(240)) or (layer0_outputs(4474));
    outputs(10712) <= not((layer0_outputs(8049)) and (layer0_outputs(7154)));
    outputs(10713) <= not((layer0_outputs(6247)) xor (layer0_outputs(7287)));
    outputs(10714) <= not((layer0_outputs(10616)) xor (layer0_outputs(5157)));
    outputs(10715) <= not(layer0_outputs(3472)) or (layer0_outputs(2002));
    outputs(10716) <= layer0_outputs(2971);
    outputs(10717) <= layer0_outputs(8623);
    outputs(10718) <= not(layer0_outputs(3489)) or (layer0_outputs(4831));
    outputs(10719) <= layer0_outputs(4164);
    outputs(10720) <= not(layer0_outputs(12324));
    outputs(10721) <= not((layer0_outputs(6711)) and (layer0_outputs(1735)));
    outputs(10722) <= not(layer0_outputs(3354)) or (layer0_outputs(12609));
    outputs(10723) <= (layer0_outputs(7421)) and not (layer0_outputs(1923));
    outputs(10724) <= (layer0_outputs(5907)) xor (layer0_outputs(12474));
    outputs(10725) <= '0';
    outputs(10726) <= layer0_outputs(2799);
    outputs(10727) <= not(layer0_outputs(12571));
    outputs(10728) <= not((layer0_outputs(5746)) xor (layer0_outputs(7210)));
    outputs(10729) <= layer0_outputs(10872);
    outputs(10730) <= (layer0_outputs(6037)) xor (layer0_outputs(2543));
    outputs(10731) <= (layer0_outputs(4675)) xor (layer0_outputs(3111));
    outputs(10732) <= not((layer0_outputs(6429)) and (layer0_outputs(2503)));
    outputs(10733) <= (layer0_outputs(3813)) xor (layer0_outputs(9741));
    outputs(10734) <= layer0_outputs(3599);
    outputs(10735) <= layer0_outputs(2473);
    outputs(10736) <= (layer0_outputs(4524)) and not (layer0_outputs(9143));
    outputs(10737) <= (layer0_outputs(9508)) and (layer0_outputs(11230));
    outputs(10738) <= not(layer0_outputs(5927));
    outputs(10739) <= (layer0_outputs(1436)) xor (layer0_outputs(4846));
    outputs(10740) <= layer0_outputs(9141);
    outputs(10741) <= not(layer0_outputs(3144));
    outputs(10742) <= not((layer0_outputs(856)) xor (layer0_outputs(7174)));
    outputs(10743) <= (layer0_outputs(11018)) and not (layer0_outputs(5578));
    outputs(10744) <= not(layer0_outputs(4533));
    outputs(10745) <= (layer0_outputs(2127)) and not (layer0_outputs(12315));
    outputs(10746) <= (layer0_outputs(1289)) xor (layer0_outputs(9060));
    outputs(10747) <= not((layer0_outputs(4019)) and (layer0_outputs(11673)));
    outputs(10748) <= not((layer0_outputs(4429)) xor (layer0_outputs(7009)));
    outputs(10749) <= not(layer0_outputs(3522));
    outputs(10750) <= layer0_outputs(11144);
    outputs(10751) <= not(layer0_outputs(6424));
    outputs(10752) <= not((layer0_outputs(9208)) xor (layer0_outputs(5169)));
    outputs(10753) <= layer0_outputs(3440);
    outputs(10754) <= (layer0_outputs(1284)) and (layer0_outputs(7509));
    outputs(10755) <= (layer0_outputs(5621)) xor (layer0_outputs(12144));
    outputs(10756) <= (layer0_outputs(1614)) xor (layer0_outputs(3378));
    outputs(10757) <= not((layer0_outputs(9853)) xor (layer0_outputs(8580)));
    outputs(10758) <= layer0_outputs(5708);
    outputs(10759) <= (layer0_outputs(4857)) or (layer0_outputs(5126));
    outputs(10760) <= (layer0_outputs(6115)) or (layer0_outputs(12760));
    outputs(10761) <= layer0_outputs(11631);
    outputs(10762) <= (layer0_outputs(10377)) and not (layer0_outputs(4321));
    outputs(10763) <= (layer0_outputs(5685)) xor (layer0_outputs(1390));
    outputs(10764) <= (layer0_outputs(5504)) and not (layer0_outputs(10817));
    outputs(10765) <= not(layer0_outputs(7656));
    outputs(10766) <= (layer0_outputs(12208)) and not (layer0_outputs(2557));
    outputs(10767) <= (layer0_outputs(1320)) and not (layer0_outputs(11276));
    outputs(10768) <= (layer0_outputs(11605)) and not (layer0_outputs(9627));
    outputs(10769) <= layer0_outputs(5022);
    outputs(10770) <= not(layer0_outputs(7300));
    outputs(10771) <= not(layer0_outputs(4780)) or (layer0_outputs(7830));
    outputs(10772) <= not((layer0_outputs(7907)) xor (layer0_outputs(6431)));
    outputs(10773) <= not(layer0_outputs(1616));
    outputs(10774) <= (layer0_outputs(9928)) and not (layer0_outputs(7984));
    outputs(10775) <= not(layer0_outputs(6956));
    outputs(10776) <= (layer0_outputs(2829)) xor (layer0_outputs(577));
    outputs(10777) <= not(layer0_outputs(3096));
    outputs(10778) <= layer0_outputs(1105);
    outputs(10779) <= not(layer0_outputs(9380));
    outputs(10780) <= layer0_outputs(5380);
    outputs(10781) <= layer0_outputs(8591);
    outputs(10782) <= not((layer0_outputs(2625)) and (layer0_outputs(2095)));
    outputs(10783) <= layer0_outputs(11686);
    outputs(10784) <= not(layer0_outputs(4876)) or (layer0_outputs(5138));
    outputs(10785) <= (layer0_outputs(8472)) or (layer0_outputs(7577));
    outputs(10786) <= not((layer0_outputs(5790)) xor (layer0_outputs(12462)));
    outputs(10787) <= not(layer0_outputs(11155));
    outputs(10788) <= layer0_outputs(2332);
    outputs(10789) <= (layer0_outputs(9866)) and not (layer0_outputs(11577));
    outputs(10790) <= layer0_outputs(1572);
    outputs(10791) <= (layer0_outputs(197)) and (layer0_outputs(9862));
    outputs(10792) <= not(layer0_outputs(4853));
    outputs(10793) <= (layer0_outputs(297)) xor (layer0_outputs(1677));
    outputs(10794) <= not(layer0_outputs(3369));
    outputs(10795) <= not(layer0_outputs(10160));
    outputs(10796) <= (layer0_outputs(3781)) xor (layer0_outputs(2076));
    outputs(10797) <= not(layer0_outputs(12188));
    outputs(10798) <= (layer0_outputs(5714)) or (layer0_outputs(37));
    outputs(10799) <= not(layer0_outputs(7588)) or (layer0_outputs(6236));
    outputs(10800) <= not(layer0_outputs(9803));
    outputs(10801) <= not((layer0_outputs(11177)) and (layer0_outputs(8840)));
    outputs(10802) <= (layer0_outputs(11480)) or (layer0_outputs(8372));
    outputs(10803) <= not(layer0_outputs(8038)) or (layer0_outputs(4319));
    outputs(10804) <= not((layer0_outputs(8138)) xor (layer0_outputs(1328)));
    outputs(10805) <= layer0_outputs(11669);
    outputs(10806) <= not(layer0_outputs(7105)) or (layer0_outputs(243));
    outputs(10807) <= not((layer0_outputs(9155)) xor (layer0_outputs(9631)));
    outputs(10808) <= not(layer0_outputs(12636)) or (layer0_outputs(8018));
    outputs(10809) <= (layer0_outputs(11052)) and not (layer0_outputs(8991));
    outputs(10810) <= not(layer0_outputs(3467));
    outputs(10811) <= not(layer0_outputs(1064));
    outputs(10812) <= not(layer0_outputs(8278));
    outputs(10813) <= layer0_outputs(846);
    outputs(10814) <= layer0_outputs(1045);
    outputs(10815) <= not(layer0_outputs(1414)) or (layer0_outputs(10876));
    outputs(10816) <= not(layer0_outputs(5070));
    outputs(10817) <= not(layer0_outputs(8316));
    outputs(10818) <= not((layer0_outputs(2838)) or (layer0_outputs(2760)));
    outputs(10819) <= (layer0_outputs(5338)) xor (layer0_outputs(5263));
    outputs(10820) <= not((layer0_outputs(6270)) and (layer0_outputs(12674)));
    outputs(10821) <= not((layer0_outputs(10160)) and (layer0_outputs(3632)));
    outputs(10822) <= not(layer0_outputs(12437));
    outputs(10823) <= layer0_outputs(6325);
    outputs(10824) <= not(layer0_outputs(12545));
    outputs(10825) <= not(layer0_outputs(1399));
    outputs(10826) <= (layer0_outputs(11290)) and not (layer0_outputs(10672));
    outputs(10827) <= (layer0_outputs(7055)) or (layer0_outputs(7012));
    outputs(10828) <= (layer0_outputs(6574)) xor (layer0_outputs(1938));
    outputs(10829) <= not(layer0_outputs(11646)) or (layer0_outputs(7474));
    outputs(10830) <= not((layer0_outputs(9128)) xor (layer0_outputs(9789)));
    outputs(10831) <= not((layer0_outputs(11116)) xor (layer0_outputs(3917)));
    outputs(10832) <= not((layer0_outputs(1617)) xor (layer0_outputs(7085)));
    outputs(10833) <= layer0_outputs(9644);
    outputs(10834) <= (layer0_outputs(1991)) xor (layer0_outputs(5830));
    outputs(10835) <= not(layer0_outputs(6491));
    outputs(10836) <= not(layer0_outputs(6804)) or (layer0_outputs(11005));
    outputs(10837) <= (layer0_outputs(8649)) xor (layer0_outputs(8384));
    outputs(10838) <= layer0_outputs(11690);
    outputs(10839) <= not(layer0_outputs(11584));
    outputs(10840) <= '0';
    outputs(10841) <= (layer0_outputs(1243)) xor (layer0_outputs(12508));
    outputs(10842) <= (layer0_outputs(5455)) or (layer0_outputs(8610));
    outputs(10843) <= not((layer0_outputs(4291)) xor (layer0_outputs(8573)));
    outputs(10844) <= not(layer0_outputs(10832));
    outputs(10845) <= not(layer0_outputs(3744));
    outputs(10846) <= layer0_outputs(12624);
    outputs(10847) <= (layer0_outputs(11932)) xor (layer0_outputs(7965));
    outputs(10848) <= (layer0_outputs(2685)) xor (layer0_outputs(1838));
    outputs(10849) <= not((layer0_outputs(7599)) and (layer0_outputs(7867)));
    outputs(10850) <= (layer0_outputs(12717)) and not (layer0_outputs(9182));
    outputs(10851) <= not((layer0_outputs(6671)) xor (layer0_outputs(10252)));
    outputs(10852) <= (layer0_outputs(385)) and not (layer0_outputs(3136));
    outputs(10853) <= not((layer0_outputs(624)) and (layer0_outputs(5026)));
    outputs(10854) <= not(layer0_outputs(12617));
    outputs(10855) <= not(layer0_outputs(4740)) or (layer0_outputs(8050));
    outputs(10856) <= layer0_outputs(11375);
    outputs(10857) <= not((layer0_outputs(9415)) and (layer0_outputs(5416)));
    outputs(10858) <= layer0_outputs(11619);
    outputs(10859) <= layer0_outputs(3952);
    outputs(10860) <= (layer0_outputs(12018)) and (layer0_outputs(3988));
    outputs(10861) <= not(layer0_outputs(7584));
    outputs(10862) <= not(layer0_outputs(10939)) or (layer0_outputs(11982));
    outputs(10863) <= not((layer0_outputs(8791)) xor (layer0_outputs(6333)));
    outputs(10864) <= not((layer0_outputs(3840)) and (layer0_outputs(6736)));
    outputs(10865) <= not((layer0_outputs(4553)) xor (layer0_outputs(6218)));
    outputs(10866) <= not(layer0_outputs(10684));
    outputs(10867) <= not(layer0_outputs(1167));
    outputs(10868) <= (layer0_outputs(7507)) xor (layer0_outputs(2797));
    outputs(10869) <= not(layer0_outputs(8716)) or (layer0_outputs(1439));
    outputs(10870) <= not(layer0_outputs(6238)) or (layer0_outputs(5020));
    outputs(10871) <= (layer0_outputs(5203)) xor (layer0_outputs(4596));
    outputs(10872) <= not(layer0_outputs(8763)) or (layer0_outputs(4941));
    outputs(10873) <= layer0_outputs(11108);
    outputs(10874) <= not(layer0_outputs(3191));
    outputs(10875) <= layer0_outputs(3795);
    outputs(10876) <= not(layer0_outputs(6573));
    outputs(10877) <= not((layer0_outputs(9970)) or (layer0_outputs(1370)));
    outputs(10878) <= not((layer0_outputs(4334)) xor (layer0_outputs(6838)));
    outputs(10879) <= not((layer0_outputs(7327)) xor (layer0_outputs(562)));
    outputs(10880) <= (layer0_outputs(5965)) xor (layer0_outputs(2378));
    outputs(10881) <= layer0_outputs(1389);
    outputs(10882) <= not((layer0_outputs(4887)) and (layer0_outputs(4531)));
    outputs(10883) <= (layer0_outputs(4557)) and not (layer0_outputs(2832));
    outputs(10884) <= not(layer0_outputs(4339));
    outputs(10885) <= not(layer0_outputs(3264));
    outputs(10886) <= not(layer0_outputs(5980)) or (layer0_outputs(3974));
    outputs(10887) <= layer0_outputs(10561);
    outputs(10888) <= not(layer0_outputs(7326));
    outputs(10889) <= not(layer0_outputs(5304)) or (layer0_outputs(11658));
    outputs(10890) <= (layer0_outputs(12763)) and not (layer0_outputs(3950));
    outputs(10891) <= not((layer0_outputs(11699)) xor (layer0_outputs(8610)));
    outputs(10892) <= '1';
    outputs(10893) <= not(layer0_outputs(2836));
    outputs(10894) <= not(layer0_outputs(6922));
    outputs(10895) <= (layer0_outputs(9477)) xor (layer0_outputs(8994));
    outputs(10896) <= not((layer0_outputs(1369)) and (layer0_outputs(903)));
    outputs(10897) <= (layer0_outputs(12588)) xor (layer0_outputs(832));
    outputs(10898) <= not(layer0_outputs(4965)) or (layer0_outputs(2026));
    outputs(10899) <= layer0_outputs(12779);
    outputs(10900) <= layer0_outputs(5334);
    outputs(10901) <= not((layer0_outputs(4730)) xor (layer0_outputs(2905)));
    outputs(10902) <= (layer0_outputs(9799)) xor (layer0_outputs(9603));
    outputs(10903) <= layer0_outputs(9520);
    outputs(10904) <= not((layer0_outputs(5091)) and (layer0_outputs(5277)));
    outputs(10905) <= not(layer0_outputs(6209));
    outputs(10906) <= layer0_outputs(3760);
    outputs(10907) <= (layer0_outputs(3709)) and (layer0_outputs(7102));
    outputs(10908) <= layer0_outputs(11640);
    outputs(10909) <= not(layer0_outputs(6960));
    outputs(10910) <= (layer0_outputs(11435)) and not (layer0_outputs(9590));
    outputs(10911) <= not((layer0_outputs(12522)) or (layer0_outputs(3206)));
    outputs(10912) <= not(layer0_outputs(1028));
    outputs(10913) <= not(layer0_outputs(4458)) or (layer0_outputs(7145));
    outputs(10914) <= not((layer0_outputs(8105)) xor (layer0_outputs(6164)));
    outputs(10915) <= not(layer0_outputs(6504)) or (layer0_outputs(4367));
    outputs(10916) <= not(layer0_outputs(4376));
    outputs(10917) <= not((layer0_outputs(10861)) and (layer0_outputs(2682)));
    outputs(10918) <= layer0_outputs(7794);
    outputs(10919) <= layer0_outputs(2013);
    outputs(10920) <= layer0_outputs(6446);
    outputs(10921) <= not(layer0_outputs(9541));
    outputs(10922) <= not((layer0_outputs(10566)) and (layer0_outputs(9926)));
    outputs(10923) <= layer0_outputs(12231);
    outputs(10924) <= (layer0_outputs(11603)) and not (layer0_outputs(2009));
    outputs(10925) <= (layer0_outputs(68)) xor (layer0_outputs(6998));
    outputs(10926) <= (layer0_outputs(6702)) and not (layer0_outputs(2259));
    outputs(10927) <= '0';
    outputs(10928) <= not(layer0_outputs(1828));
    outputs(10929) <= (layer0_outputs(12180)) or (layer0_outputs(3143));
    outputs(10930) <= layer0_outputs(7315);
    outputs(10931) <= layer0_outputs(5539);
    outputs(10932) <= layer0_outputs(4607);
    outputs(10933) <= not((layer0_outputs(8330)) xor (layer0_outputs(2083)));
    outputs(10934) <= not(layer0_outputs(5450)) or (layer0_outputs(2148));
    outputs(10935) <= not((layer0_outputs(9239)) xor (layer0_outputs(3501)));
    outputs(10936) <= (layer0_outputs(2760)) xor (layer0_outputs(2654));
    outputs(10937) <= not(layer0_outputs(10954));
    outputs(10938) <= (layer0_outputs(7343)) xor (layer0_outputs(4875));
    outputs(10939) <= (layer0_outputs(9144)) xor (layer0_outputs(2749));
    outputs(10940) <= not(layer0_outputs(8704)) or (layer0_outputs(9526));
    outputs(10941) <= (layer0_outputs(3566)) and not (layer0_outputs(9096));
    outputs(10942) <= not(layer0_outputs(1020));
    outputs(10943) <= not((layer0_outputs(7383)) xor (layer0_outputs(6089)));
    outputs(10944) <= (layer0_outputs(6243)) or (layer0_outputs(11533));
    outputs(10945) <= not((layer0_outputs(11352)) xor (layer0_outputs(11354)));
    outputs(10946) <= layer0_outputs(2531);
    outputs(10947) <= (layer0_outputs(676)) and not (layer0_outputs(4303));
    outputs(10948) <= not(layer0_outputs(7677));
    outputs(10949) <= not((layer0_outputs(10462)) or (layer0_outputs(7266)));
    outputs(10950) <= (layer0_outputs(12697)) or (layer0_outputs(4960));
    outputs(10951) <= layer0_outputs(6697);
    outputs(10952) <= (layer0_outputs(1963)) or (layer0_outputs(6062));
    outputs(10953) <= not((layer0_outputs(560)) xor (layer0_outputs(12376)));
    outputs(10954) <= (layer0_outputs(11140)) xor (layer0_outputs(12732));
    outputs(10955) <= (layer0_outputs(10890)) xor (layer0_outputs(2375));
    outputs(10956) <= not(layer0_outputs(10109));
    outputs(10957) <= not(layer0_outputs(2880));
    outputs(10958) <= (layer0_outputs(333)) xor (layer0_outputs(9384));
    outputs(10959) <= not(layer0_outputs(9938)) or (layer0_outputs(9539));
    outputs(10960) <= not((layer0_outputs(3633)) and (layer0_outputs(11930)));
    outputs(10961) <= layer0_outputs(3949);
    outputs(10962) <= (layer0_outputs(10468)) and not (layer0_outputs(3994));
    outputs(10963) <= (layer0_outputs(6677)) and (layer0_outputs(10730));
    outputs(10964) <= (layer0_outputs(6559)) and not (layer0_outputs(6186));
    outputs(10965) <= not(layer0_outputs(10137));
    outputs(10966) <= layer0_outputs(3220);
    outputs(10967) <= not(layer0_outputs(1)) or (layer0_outputs(10450));
    outputs(10968) <= not((layer0_outputs(8017)) and (layer0_outputs(420)));
    outputs(10969) <= (layer0_outputs(2723)) or (layer0_outputs(4635));
    outputs(10970) <= not((layer0_outputs(10776)) and (layer0_outputs(6530)));
    outputs(10971) <= (layer0_outputs(6101)) xor (layer0_outputs(3466));
    outputs(10972) <= (layer0_outputs(6753)) or (layer0_outputs(3989));
    outputs(10973) <= not(layer0_outputs(2167));
    outputs(10974) <= layer0_outputs(10409);
    outputs(10975) <= layer0_outputs(9163);
    outputs(10976) <= not(layer0_outputs(7789));
    outputs(10977) <= (layer0_outputs(8191)) xor (layer0_outputs(1189));
    outputs(10978) <= (layer0_outputs(11415)) xor (layer0_outputs(12047));
    outputs(10979) <= layer0_outputs(4709);
    outputs(10980) <= layer0_outputs(3335);
    outputs(10981) <= (layer0_outputs(7998)) or (layer0_outputs(12300));
    outputs(10982) <= not((layer0_outputs(8589)) and (layer0_outputs(1834)));
    outputs(10983) <= layer0_outputs(8224);
    outputs(10984) <= (layer0_outputs(2474)) or (layer0_outputs(1036));
    outputs(10985) <= (layer0_outputs(3488)) xor (layer0_outputs(12060));
    outputs(10986) <= layer0_outputs(12551);
    outputs(10987) <= not((layer0_outputs(10665)) and (layer0_outputs(5376)));
    outputs(10988) <= not((layer0_outputs(7687)) and (layer0_outputs(10993)));
    outputs(10989) <= (layer0_outputs(3525)) and (layer0_outputs(4170));
    outputs(10990) <= (layer0_outputs(6027)) and not (layer0_outputs(8813));
    outputs(10991) <= not(layer0_outputs(22)) or (layer0_outputs(6145));
    outputs(10992) <= layer0_outputs(10626);
    outputs(10993) <= not((layer0_outputs(11784)) xor (layer0_outputs(3063)));
    outputs(10994) <= not((layer0_outputs(10072)) and (layer0_outputs(9198)));
    outputs(10995) <= (layer0_outputs(4085)) xor (layer0_outputs(1003));
    outputs(10996) <= not((layer0_outputs(8742)) and (layer0_outputs(4692)));
    outputs(10997) <= (layer0_outputs(11904)) xor (layer0_outputs(4946));
    outputs(10998) <= layer0_outputs(1147);
    outputs(10999) <= (layer0_outputs(3221)) and (layer0_outputs(720));
    outputs(11000) <= (layer0_outputs(7357)) xor (layer0_outputs(4767));
    outputs(11001) <= (layer0_outputs(8059)) and not (layer0_outputs(4146));
    outputs(11002) <= not(layer0_outputs(7807)) or (layer0_outputs(4059));
    outputs(11003) <= not((layer0_outputs(3421)) xor (layer0_outputs(7962)));
    outputs(11004) <= not((layer0_outputs(9017)) xor (layer0_outputs(1134)));
    outputs(11005) <= not((layer0_outputs(820)) xor (layer0_outputs(11481)));
    outputs(11006) <= (layer0_outputs(2526)) xor (layer0_outputs(6246));
    outputs(11007) <= not(layer0_outputs(9368)) or (layer0_outputs(2900));
    outputs(11008) <= not(layer0_outputs(3376));
    outputs(11009) <= not((layer0_outputs(4110)) xor (layer0_outputs(2754)));
    outputs(11010) <= not(layer0_outputs(8796));
    outputs(11011) <= layer0_outputs(2468);
    outputs(11012) <= not((layer0_outputs(1499)) and (layer0_outputs(9032)));
    outputs(11013) <= not((layer0_outputs(3503)) xor (layer0_outputs(7686)));
    outputs(11014) <= not(layer0_outputs(12562));
    outputs(11015) <= (layer0_outputs(4466)) and (layer0_outputs(12441));
    outputs(11016) <= (layer0_outputs(11426)) and not (layer0_outputs(3492));
    outputs(11017) <= not((layer0_outputs(11314)) or (layer0_outputs(6144)));
    outputs(11018) <= layer0_outputs(2383);
    outputs(11019) <= not((layer0_outputs(7082)) xor (layer0_outputs(1441)));
    outputs(11020) <= layer0_outputs(129);
    outputs(11021) <= (layer0_outputs(7470)) and not (layer0_outputs(4554));
    outputs(11022) <= (layer0_outputs(4360)) and not (layer0_outputs(9937));
    outputs(11023) <= (layer0_outputs(8069)) xor (layer0_outputs(4258));
    outputs(11024) <= not((layer0_outputs(7042)) xor (layer0_outputs(8715)));
    outputs(11025) <= not(layer0_outputs(9097));
    outputs(11026) <= (layer0_outputs(6010)) and (layer0_outputs(622));
    outputs(11027) <= not((layer0_outputs(5610)) xor (layer0_outputs(6527)));
    outputs(11028) <= (layer0_outputs(10883)) and not (layer0_outputs(12367));
    outputs(11029) <= not(layer0_outputs(11990));
    outputs(11030) <= layer0_outputs(7724);
    outputs(11031) <= layer0_outputs(5509);
    outputs(11032) <= not((layer0_outputs(8228)) xor (layer0_outputs(11876)));
    outputs(11033) <= not(layer0_outputs(11997));
    outputs(11034) <= layer0_outputs(9074);
    outputs(11035) <= (layer0_outputs(482)) xor (layer0_outputs(391));
    outputs(11036) <= (layer0_outputs(7478)) xor (layer0_outputs(8965));
    outputs(11037) <= not((layer0_outputs(158)) xor (layer0_outputs(12364)));
    outputs(11038) <= layer0_outputs(11643);
    outputs(11039) <= not(layer0_outputs(654));
    outputs(11040) <= (layer0_outputs(9179)) or (layer0_outputs(11523));
    outputs(11041) <= not(layer0_outputs(3163)) or (layer0_outputs(8564));
    outputs(11042) <= layer0_outputs(8706);
    outputs(11043) <= not((layer0_outputs(5257)) xor (layer0_outputs(2349)));
    outputs(11044) <= not((layer0_outputs(263)) xor (layer0_outputs(12268)));
    outputs(11045) <= not(layer0_outputs(6705));
    outputs(11046) <= not(layer0_outputs(6356)) or (layer0_outputs(2983));
    outputs(11047) <= (layer0_outputs(6524)) xor (layer0_outputs(7444));
    outputs(11048) <= (layer0_outputs(10308)) xor (layer0_outputs(5279));
    outputs(11049) <= not(layer0_outputs(5994)) or (layer0_outputs(5637));
    outputs(11050) <= layer0_outputs(5329);
    outputs(11051) <= (layer0_outputs(304)) xor (layer0_outputs(9295));
    outputs(11052) <= layer0_outputs(6733);
    outputs(11053) <= (layer0_outputs(400)) xor (layer0_outputs(8333));
    outputs(11054) <= (layer0_outputs(10025)) xor (layer0_outputs(3387));
    outputs(11055) <= (layer0_outputs(7434)) xor (layer0_outputs(3761));
    outputs(11056) <= not((layer0_outputs(4894)) xor (layer0_outputs(11844)));
    outputs(11057) <= layer0_outputs(12418);
    outputs(11058) <= not((layer0_outputs(9256)) or (layer0_outputs(4232)));
    outputs(11059) <= not(layer0_outputs(7812)) or (layer0_outputs(2884));
    outputs(11060) <= layer0_outputs(8012);
    outputs(11061) <= not(layer0_outputs(11066)) or (layer0_outputs(12230));
    outputs(11062) <= not((layer0_outputs(11052)) xor (layer0_outputs(3684)));
    outputs(11063) <= not((layer0_outputs(4270)) xor (layer0_outputs(9193)));
    outputs(11064) <= not(layer0_outputs(3405)) or (layer0_outputs(4831));
    outputs(11065) <= (layer0_outputs(10639)) or (layer0_outputs(7098));
    outputs(11066) <= layer0_outputs(6726);
    outputs(11067) <= not((layer0_outputs(10307)) or (layer0_outputs(515)));
    outputs(11068) <= layer0_outputs(10591);
    outputs(11069) <= not((layer0_outputs(3010)) xor (layer0_outputs(4561)));
    outputs(11070) <= not((layer0_outputs(504)) and (layer0_outputs(7683)));
    outputs(11071) <= not(layer0_outputs(1018)) or (layer0_outputs(2218));
    outputs(11072) <= (layer0_outputs(3977)) and not (layer0_outputs(11863));
    outputs(11073) <= not((layer0_outputs(5588)) xor (layer0_outputs(11164)));
    outputs(11074) <= (layer0_outputs(8771)) xor (layer0_outputs(8667));
    outputs(11075) <= not((layer0_outputs(6539)) xor (layer0_outputs(3422)));
    outputs(11076) <= (layer0_outputs(11455)) and not (layer0_outputs(10504));
    outputs(11077) <= layer0_outputs(9145);
    outputs(11078) <= layer0_outputs(9747);
    outputs(11079) <= not((layer0_outputs(2992)) or (layer0_outputs(1892)));
    outputs(11080) <= (layer0_outputs(11967)) xor (layer0_outputs(7943));
    outputs(11081) <= not((layer0_outputs(4417)) or (layer0_outputs(11098)));
    outputs(11082) <= not(layer0_outputs(7214));
    outputs(11083) <= (layer0_outputs(7476)) xor (layer0_outputs(5866));
    outputs(11084) <= '1';
    outputs(11085) <= not((layer0_outputs(3351)) and (layer0_outputs(10202)));
    outputs(11086) <= not(layer0_outputs(3214)) or (layer0_outputs(590));
    outputs(11087) <= not(layer0_outputs(10951)) or (layer0_outputs(5860));
    outputs(11088) <= layer0_outputs(4990);
    outputs(11089) <= (layer0_outputs(2128)) xor (layer0_outputs(2157));
    outputs(11090) <= not(layer0_outputs(11874)) or (layer0_outputs(11969));
    outputs(11091) <= not(layer0_outputs(797));
    outputs(11092) <= not(layer0_outputs(2940));
    outputs(11093) <= (layer0_outputs(9436)) xor (layer0_outputs(7495));
    outputs(11094) <= (layer0_outputs(4880)) and not (layer0_outputs(7410));
    outputs(11095) <= layer0_outputs(1410);
    outputs(11096) <= not(layer0_outputs(11543));
    outputs(11097) <= not(layer0_outputs(8632));
    outputs(11098) <= '1';
    outputs(11099) <= layer0_outputs(8588);
    outputs(11100) <= layer0_outputs(7033);
    outputs(11101) <= layer0_outputs(12256);
    outputs(11102) <= not(layer0_outputs(11839));
    outputs(11103) <= not(layer0_outputs(1256));
    outputs(11104) <= not((layer0_outputs(10193)) and (layer0_outputs(9919)));
    outputs(11105) <= not((layer0_outputs(7109)) xor (layer0_outputs(5558)));
    outputs(11106) <= not(layer0_outputs(7680));
    outputs(11107) <= not(layer0_outputs(11220));
    outputs(11108) <= not((layer0_outputs(8365)) or (layer0_outputs(6828)));
    outputs(11109) <= layer0_outputs(2469);
    outputs(11110) <= (layer0_outputs(841)) or (layer0_outputs(7219));
    outputs(11111) <= '1';
    outputs(11112) <= layer0_outputs(5374);
    outputs(11113) <= not(layer0_outputs(10088));
    outputs(11114) <= (layer0_outputs(10291)) and (layer0_outputs(9878));
    outputs(11115) <= not(layer0_outputs(8405));
    outputs(11116) <= not(layer0_outputs(4974));
    outputs(11117) <= not(layer0_outputs(3270));
    outputs(11118) <= (layer0_outputs(2255)) or (layer0_outputs(11796));
    outputs(11119) <= not(layer0_outputs(8965)) or (layer0_outputs(7182));
    outputs(11120) <= layer0_outputs(4438);
    outputs(11121) <= layer0_outputs(1238);
    outputs(11122) <= (layer0_outputs(11461)) xor (layer0_outputs(592));
    outputs(11123) <= not(layer0_outputs(5503));
    outputs(11124) <= not((layer0_outputs(898)) xor (layer0_outputs(1811)));
    outputs(11125) <= not(layer0_outputs(10320)) or (layer0_outputs(11791));
    outputs(11126) <= layer0_outputs(5293);
    outputs(11127) <= not(layer0_outputs(159));
    outputs(11128) <= not((layer0_outputs(12626)) xor (layer0_outputs(5169)));
    outputs(11129) <= (layer0_outputs(2587)) xor (layer0_outputs(5849));
    outputs(11130) <= not(layer0_outputs(1891)) or (layer0_outputs(3239));
    outputs(11131) <= (layer0_outputs(7399)) xor (layer0_outputs(11621));
    outputs(11132) <= not(layer0_outputs(5907));
    outputs(11133) <= layer0_outputs(12307);
    outputs(11134) <= not((layer0_outputs(1644)) xor (layer0_outputs(12527)));
    outputs(11135) <= not((layer0_outputs(12163)) xor (layer0_outputs(9676)));
    outputs(11136) <= layer0_outputs(3055);
    outputs(11137) <= not(layer0_outputs(6014));
    outputs(11138) <= not(layer0_outputs(8004));
    outputs(11139) <= (layer0_outputs(6341)) and (layer0_outputs(10651));
    outputs(11140) <= not((layer0_outputs(4551)) xor (layer0_outputs(3022)));
    outputs(11141) <= layer0_outputs(3756);
    outputs(11142) <= (layer0_outputs(1177)) or (layer0_outputs(8447));
    outputs(11143) <= not((layer0_outputs(11481)) xor (layer0_outputs(11412)));
    outputs(11144) <= not((layer0_outputs(362)) and (layer0_outputs(2813)));
    outputs(11145) <= not(layer0_outputs(8981));
    outputs(11146) <= not(layer0_outputs(5524)) or (layer0_outputs(6113));
    outputs(11147) <= not(layer0_outputs(11562));
    outputs(11148) <= not((layer0_outputs(2590)) xor (layer0_outputs(2669)));
    outputs(11149) <= not((layer0_outputs(10802)) xor (layer0_outputs(9854)));
    outputs(11150) <= not(layer0_outputs(8513));
    outputs(11151) <= layer0_outputs(2250);
    outputs(11152) <= (layer0_outputs(4244)) xor (layer0_outputs(881));
    outputs(11153) <= not((layer0_outputs(8611)) and (layer0_outputs(11646)));
    outputs(11154) <= (layer0_outputs(12022)) and (layer0_outputs(7981));
    outputs(11155) <= not(layer0_outputs(3820));
    outputs(11156) <= (layer0_outputs(2409)) and not (layer0_outputs(8726));
    outputs(11157) <= not((layer0_outputs(8230)) xor (layer0_outputs(1005)));
    outputs(11158) <= not((layer0_outputs(11802)) xor (layer0_outputs(6186)));
    outputs(11159) <= (layer0_outputs(6213)) xor (layer0_outputs(1398));
    outputs(11160) <= not(layer0_outputs(378));
    outputs(11161) <= (layer0_outputs(2194)) or (layer0_outputs(7189));
    outputs(11162) <= layer0_outputs(2156);
    outputs(11163) <= not((layer0_outputs(6319)) and (layer0_outputs(8579)));
    outputs(11164) <= not(layer0_outputs(6461));
    outputs(11165) <= (layer0_outputs(11692)) xor (layer0_outputs(6594));
    outputs(11166) <= (layer0_outputs(12167)) xor (layer0_outputs(9554));
    outputs(11167) <= (layer0_outputs(1487)) and not (layer0_outputs(12191));
    outputs(11168) <= not((layer0_outputs(4979)) xor (layer0_outputs(7477)));
    outputs(11169) <= not((layer0_outputs(8721)) xor (layer0_outputs(5158)));
    outputs(11170) <= not(layer0_outputs(5636));
    outputs(11171) <= not(layer0_outputs(5230));
    outputs(11172) <= not(layer0_outputs(4020));
    outputs(11173) <= not(layer0_outputs(3041));
    outputs(11174) <= not(layer0_outputs(2506)) or (layer0_outputs(1562));
    outputs(11175) <= layer0_outputs(8049);
    outputs(11176) <= not(layer0_outputs(6606)) or (layer0_outputs(1119));
    outputs(11177) <= (layer0_outputs(3169)) and (layer0_outputs(3489));
    outputs(11178) <= not(layer0_outputs(12766));
    outputs(11179) <= (layer0_outputs(9018)) and (layer0_outputs(2354));
    outputs(11180) <= (layer0_outputs(677)) xor (layer0_outputs(11944));
    outputs(11181) <= (layer0_outputs(3217)) xor (layer0_outputs(11848));
    outputs(11182) <= not(layer0_outputs(9829)) or (layer0_outputs(978));
    outputs(11183) <= not(layer0_outputs(12102)) or (layer0_outputs(3666));
    outputs(11184) <= (layer0_outputs(12486)) or (layer0_outputs(1276));
    outputs(11185) <= (layer0_outputs(11006)) or (layer0_outputs(6260));
    outputs(11186) <= (layer0_outputs(6079)) xor (layer0_outputs(4907));
    outputs(11187) <= (layer0_outputs(4832)) and not (layer0_outputs(148));
    outputs(11188) <= (layer0_outputs(4781)) xor (layer0_outputs(10947));
    outputs(11189) <= '0';
    outputs(11190) <= not(layer0_outputs(8618));
    outputs(11191) <= not(layer0_outputs(4877));
    outputs(11192) <= (layer0_outputs(7661)) or (layer0_outputs(12635));
    outputs(11193) <= (layer0_outputs(8503)) xor (layer0_outputs(7451));
    outputs(11194) <= (layer0_outputs(8381)) xor (layer0_outputs(8532));
    outputs(11195) <= (layer0_outputs(7112)) or (layer0_outputs(10901));
    outputs(11196) <= not((layer0_outputs(6725)) xor (layer0_outputs(8726)));
    outputs(11197) <= not((layer0_outputs(1424)) or (layer0_outputs(10961)));
    outputs(11198) <= not((layer0_outputs(5832)) xor (layer0_outputs(2110)));
    outputs(11199) <= not(layer0_outputs(9885)) or (layer0_outputs(10551));
    outputs(11200) <= (layer0_outputs(4141)) xor (layer0_outputs(912));
    outputs(11201) <= (layer0_outputs(11571)) xor (layer0_outputs(10538));
    outputs(11202) <= not(layer0_outputs(8197));
    outputs(11203) <= layer0_outputs(2692);
    outputs(11204) <= not((layer0_outputs(3528)) xor (layer0_outputs(1656)));
    outputs(11205) <= layer0_outputs(2827);
    outputs(11206) <= not(layer0_outputs(5056));
    outputs(11207) <= not((layer0_outputs(8343)) and (layer0_outputs(5704)));
    outputs(11208) <= not(layer0_outputs(202));
    outputs(11209) <= not((layer0_outputs(11896)) xor (layer0_outputs(10792)));
    outputs(11210) <= layer0_outputs(6773);
    outputs(11211) <= not(layer0_outputs(7918));
    outputs(11212) <= layer0_outputs(8473);
    outputs(11213) <= (layer0_outputs(9322)) xor (layer0_outputs(4374));
    outputs(11214) <= not(layer0_outputs(7912));
    outputs(11215) <= not(layer0_outputs(2322));
    outputs(11216) <= (layer0_outputs(11315)) xor (layer0_outputs(9225));
    outputs(11217) <= not(layer0_outputs(890));
    outputs(11218) <= not((layer0_outputs(1921)) and (layer0_outputs(2295)));
    outputs(11219) <= not((layer0_outputs(2103)) xor (layer0_outputs(5780)));
    outputs(11220) <= layer0_outputs(3920);
    outputs(11221) <= not(layer0_outputs(11498));
    outputs(11222) <= not(layer0_outputs(7053));
    outputs(11223) <= (layer0_outputs(12153)) xor (layer0_outputs(10336));
    outputs(11224) <= not((layer0_outputs(6486)) xor (layer0_outputs(6063)));
    outputs(11225) <= not((layer0_outputs(3346)) and (layer0_outputs(3255)));
    outputs(11226) <= layer0_outputs(919);
    outputs(11227) <= layer0_outputs(4774);
    outputs(11228) <= (layer0_outputs(2570)) xor (layer0_outputs(7879));
    outputs(11229) <= (layer0_outputs(9409)) xor (layer0_outputs(9447));
    outputs(11230) <= (layer0_outputs(10379)) xor (layer0_outputs(3089));
    outputs(11231) <= not(layer0_outputs(6801));
    outputs(11232) <= (layer0_outputs(1369)) and not (layer0_outputs(6844));
    outputs(11233) <= not((layer0_outputs(8292)) xor (layer0_outputs(4279)));
    outputs(11234) <= layer0_outputs(9301);
    outputs(11235) <= (layer0_outputs(12454)) or (layer0_outputs(2357));
    outputs(11236) <= not(layer0_outputs(484)) or (layer0_outputs(3517));
    outputs(11237) <= layer0_outputs(4476);
    outputs(11238) <= (layer0_outputs(5539)) or (layer0_outputs(611));
    outputs(11239) <= (layer0_outputs(12577)) xor (layer0_outputs(9027));
    outputs(11240) <= layer0_outputs(10096);
    outputs(11241) <= not(layer0_outputs(8684));
    outputs(11242) <= not((layer0_outputs(10944)) xor (layer0_outputs(5323)));
    outputs(11243) <= (layer0_outputs(9574)) and (layer0_outputs(4107));
    outputs(11244) <= (layer0_outputs(2796)) xor (layer0_outputs(1637));
    outputs(11245) <= not(layer0_outputs(2805));
    outputs(11246) <= not(layer0_outputs(10244));
    outputs(11247) <= not((layer0_outputs(12326)) and (layer0_outputs(12620)));
    outputs(11248) <= not((layer0_outputs(219)) and (layer0_outputs(12159)));
    outputs(11249) <= (layer0_outputs(8075)) and (layer0_outputs(1400));
    outputs(11250) <= not(layer0_outputs(1223));
    outputs(11251) <= not(layer0_outputs(1804)) or (layer0_outputs(947));
    outputs(11252) <= not(layer0_outputs(12102));
    outputs(11253) <= not(layer0_outputs(5299));
    outputs(11254) <= not(layer0_outputs(6408)) or (layer0_outputs(2016));
    outputs(11255) <= not(layer0_outputs(7231));
    outputs(11256) <= not(layer0_outputs(4484));
    outputs(11257) <= not((layer0_outputs(2571)) xor (layer0_outputs(2250)));
    outputs(11258) <= not((layer0_outputs(2650)) xor (layer0_outputs(10925)));
    outputs(11259) <= not((layer0_outputs(6446)) xor (layer0_outputs(6216)));
    outputs(11260) <= layer0_outputs(2512);
    outputs(11261) <= (layer0_outputs(7163)) xor (layer0_outputs(491));
    outputs(11262) <= layer0_outputs(7759);
    outputs(11263) <= not((layer0_outputs(8139)) and (layer0_outputs(3330)));
    outputs(11264) <= layer0_outputs(9);
    outputs(11265) <= not(layer0_outputs(9129));
    outputs(11266) <= not((layer0_outputs(6398)) xor (layer0_outputs(10789)));
    outputs(11267) <= not(layer0_outputs(7367));
    outputs(11268) <= (layer0_outputs(8081)) xor (layer0_outputs(6233));
    outputs(11269) <= (layer0_outputs(6948)) or (layer0_outputs(5278));
    outputs(11270) <= not(layer0_outputs(5379));
    outputs(11271) <= layer0_outputs(11558);
    outputs(11272) <= (layer0_outputs(9154)) and not (layer0_outputs(11584));
    outputs(11273) <= not(layer0_outputs(10212)) or (layer0_outputs(6632));
    outputs(11274) <= (layer0_outputs(540)) xor (layer0_outputs(4371));
    outputs(11275) <= (layer0_outputs(4706)) and not (layer0_outputs(5188));
    outputs(11276) <= not((layer0_outputs(4483)) xor (layer0_outputs(5786)));
    outputs(11277) <= not(layer0_outputs(11482));
    outputs(11278) <= layer0_outputs(4025);
    outputs(11279) <= layer0_outputs(6136);
    outputs(11280) <= not((layer0_outputs(1714)) xor (layer0_outputs(12048)));
    outputs(11281) <= (layer0_outputs(2662)) or (layer0_outputs(4240));
    outputs(11282) <= not(layer0_outputs(7090)) or (layer0_outputs(11));
    outputs(11283) <= layer0_outputs(3368);
    outputs(11284) <= layer0_outputs(3407);
    outputs(11285) <= not((layer0_outputs(7928)) xor (layer0_outputs(2704)));
    outputs(11286) <= (layer0_outputs(1987)) and not (layer0_outputs(12403));
    outputs(11287) <= (layer0_outputs(4568)) or (layer0_outputs(3129));
    outputs(11288) <= not(layer0_outputs(7738));
    outputs(11289) <= not((layer0_outputs(11005)) xor (layer0_outputs(7892)));
    outputs(11290) <= layer0_outputs(12603);
    outputs(11291) <= not(layer0_outputs(9771));
    outputs(11292) <= (layer0_outputs(8151)) and (layer0_outputs(2135));
    outputs(11293) <= layer0_outputs(3673);
    outputs(11294) <= not(layer0_outputs(4208));
    outputs(11295) <= (layer0_outputs(4873)) xor (layer0_outputs(10456));
    outputs(11296) <= layer0_outputs(3860);
    outputs(11297) <= not(layer0_outputs(11232));
    outputs(11298) <= not((layer0_outputs(264)) or (layer0_outputs(5315)));
    outputs(11299) <= not((layer0_outputs(2890)) and (layer0_outputs(6103)));
    outputs(11300) <= not(layer0_outputs(12284)) or (layer0_outputs(6766));
    outputs(11301) <= (layer0_outputs(3054)) xor (layer0_outputs(1592));
    outputs(11302) <= (layer0_outputs(11565)) xor (layer0_outputs(10604));
    outputs(11303) <= not(layer0_outputs(10085)) or (layer0_outputs(10729));
    outputs(11304) <= not((layer0_outputs(506)) xor (layer0_outputs(3104)));
    outputs(11305) <= (layer0_outputs(7736)) xor (layer0_outputs(619));
    outputs(11306) <= not(layer0_outputs(10012)) or (layer0_outputs(11825));
    outputs(11307) <= not((layer0_outputs(4612)) xor (layer0_outputs(302)));
    outputs(11308) <= not((layer0_outputs(7214)) xor (layer0_outputs(4912)));
    outputs(11309) <= (layer0_outputs(6013)) and (layer0_outputs(8534));
    outputs(11310) <= (layer0_outputs(11154)) xor (layer0_outputs(2985));
    outputs(11311) <= layer0_outputs(7710);
    outputs(11312) <= layer0_outputs(1858);
    outputs(11313) <= (layer0_outputs(10766)) xor (layer0_outputs(11169));
    outputs(11314) <= layer0_outputs(1440);
    outputs(11315) <= not((layer0_outputs(330)) and (layer0_outputs(5093)));
    outputs(11316) <= layer0_outputs(4476);
    outputs(11317) <= (layer0_outputs(3890)) and (layer0_outputs(12530));
    outputs(11318) <= not(layer0_outputs(2817));
    outputs(11319) <= layer0_outputs(10143);
    outputs(11320) <= not((layer0_outputs(12053)) or (layer0_outputs(6472)));
    outputs(11321) <= not((layer0_outputs(3246)) xor (layer0_outputs(11277)));
    outputs(11322) <= not(layer0_outputs(8980));
    outputs(11323) <= not(layer0_outputs(9249));
    outputs(11324) <= layer0_outputs(5353);
    outputs(11325) <= '1';
    outputs(11326) <= not(layer0_outputs(7133)) or (layer0_outputs(9362));
    outputs(11327) <= layer0_outputs(3970);
    outputs(11328) <= not(layer0_outputs(1476));
    outputs(11329) <= (layer0_outputs(5727)) xor (layer0_outputs(10397));
    outputs(11330) <= (layer0_outputs(8972)) xor (layer0_outputs(9536));
    outputs(11331) <= (layer0_outputs(10196)) and not (layer0_outputs(5730));
    outputs(11332) <= layer0_outputs(5581);
    outputs(11333) <= layer0_outputs(8575);
    outputs(11334) <= layer0_outputs(10749);
    outputs(11335) <= layer0_outputs(4935);
    outputs(11336) <= not(layer0_outputs(1749));
    outputs(11337) <= layer0_outputs(8536);
    outputs(11338) <= layer0_outputs(12523);
    outputs(11339) <= layer0_outputs(12764);
    outputs(11340) <= not((layer0_outputs(9124)) xor (layer0_outputs(8816)));
    outputs(11341) <= not((layer0_outputs(10652)) and (layer0_outputs(1383)));
    outputs(11342) <= layer0_outputs(3676);
    outputs(11343) <= '0';
    outputs(11344) <= (layer0_outputs(4099)) xor (layer0_outputs(11515));
    outputs(11345) <= not((layer0_outputs(8498)) and (layer0_outputs(11789)));
    outputs(11346) <= layer0_outputs(3215);
    outputs(11347) <= not((layer0_outputs(6305)) xor (layer0_outputs(1729)));
    outputs(11348) <= not((layer0_outputs(11662)) xor (layer0_outputs(6509)));
    outputs(11349) <= not((layer0_outputs(4404)) xor (layer0_outputs(11130)));
    outputs(11350) <= not((layer0_outputs(1789)) xor (layer0_outputs(8090)));
    outputs(11351) <= not((layer0_outputs(8469)) xor (layer0_outputs(2407)));
    outputs(11352) <= layer0_outputs(11707);
    outputs(11353) <= layer0_outputs(7909);
    outputs(11354) <= not(layer0_outputs(9590));
    outputs(11355) <= not(layer0_outputs(8325)) or (layer0_outputs(4429));
    outputs(11356) <= layer0_outputs(12668);
    outputs(11357) <= not(layer0_outputs(8379));
    outputs(11358) <= layer0_outputs(4475);
    outputs(11359) <= layer0_outputs(6816);
    outputs(11360) <= not((layer0_outputs(11883)) xor (layer0_outputs(11711)));
    outputs(11361) <= (layer0_outputs(5815)) and (layer0_outputs(8020));
    outputs(11362) <= (layer0_outputs(455)) xor (layer0_outputs(8271));
    outputs(11363) <= (layer0_outputs(3074)) and not (layer0_outputs(9681));
    outputs(11364) <= layer0_outputs(10245);
    outputs(11365) <= not((layer0_outputs(7789)) and (layer0_outputs(1674)));
    outputs(11366) <= not((layer0_outputs(8894)) xor (layer0_outputs(11679)));
    outputs(11367) <= not((layer0_outputs(476)) xor (layer0_outputs(6407)));
    outputs(11368) <= not(layer0_outputs(12725));
    outputs(11369) <= not(layer0_outputs(11864));
    outputs(11370) <= not((layer0_outputs(6980)) and (layer0_outputs(7354)));
    outputs(11371) <= (layer0_outputs(11083)) xor (layer0_outputs(7637));
    outputs(11372) <= not((layer0_outputs(10743)) and (layer0_outputs(3294)));
    outputs(11373) <= not(layer0_outputs(3201)) or (layer0_outputs(7768));
    outputs(11374) <= (layer0_outputs(3737)) and not (layer0_outputs(1399));
    outputs(11375) <= not(layer0_outputs(11927));
    outputs(11376) <= layer0_outputs(8323);
    outputs(11377) <= not(layer0_outputs(5055)) or (layer0_outputs(12773));
    outputs(11378) <= (layer0_outputs(4453)) xor (layer0_outputs(5856));
    outputs(11379) <= not((layer0_outputs(12397)) xor (layer0_outputs(5011)));
    outputs(11380) <= (layer0_outputs(5614)) or (layer0_outputs(11460));
    outputs(11381) <= layer0_outputs(7235);
    outputs(11382) <= layer0_outputs(5045);
    outputs(11383) <= not((layer0_outputs(12798)) and (layer0_outputs(6223)));
    outputs(11384) <= not((layer0_outputs(11707)) xor (layer0_outputs(145)));
    outputs(11385) <= layer0_outputs(3826);
    outputs(11386) <= not(layer0_outputs(6575));
    outputs(11387) <= (layer0_outputs(2923)) or (layer0_outputs(9855));
    outputs(11388) <= not(layer0_outputs(3754));
    outputs(11389) <= not((layer0_outputs(255)) xor (layer0_outputs(5454)));
    outputs(11390) <= not(layer0_outputs(4741));
    outputs(11391) <= not(layer0_outputs(1966)) or (layer0_outputs(7571));
    outputs(11392) <= (layer0_outputs(7260)) or (layer0_outputs(10068));
    outputs(11393) <= not(layer0_outputs(4172));
    outputs(11394) <= not((layer0_outputs(11063)) xor (layer0_outputs(7721)));
    outputs(11395) <= layer0_outputs(1019);
    outputs(11396) <= layer0_outputs(7064);
    outputs(11397) <= (layer0_outputs(1591)) or (layer0_outputs(8401));
    outputs(11398) <= (layer0_outputs(2058)) and (layer0_outputs(7180));
    outputs(11399) <= not((layer0_outputs(4055)) xor (layer0_outputs(9605)));
    outputs(11400) <= not(layer0_outputs(439));
    outputs(11401) <= not(layer0_outputs(4757)) or (layer0_outputs(3654));
    outputs(11402) <= (layer0_outputs(5869)) and not (layer0_outputs(10948));
    outputs(11403) <= (layer0_outputs(5968)) xor (layer0_outputs(7904));
    outputs(11404) <= '0';
    outputs(11405) <= (layer0_outputs(8959)) xor (layer0_outputs(12004));
    outputs(11406) <= (layer0_outputs(5817)) xor (layer0_outputs(10323));
    outputs(11407) <= not((layer0_outputs(9898)) xor (layer0_outputs(10759)));
    outputs(11408) <= not((layer0_outputs(12488)) xor (layer0_outputs(10461)));
    outputs(11409) <= layer0_outputs(12702);
    outputs(11410) <= not((layer0_outputs(11893)) and (layer0_outputs(5067)));
    outputs(11411) <= layer0_outputs(9163);
    outputs(11412) <= layer0_outputs(12220);
    outputs(11413) <= not((layer0_outputs(12302)) or (layer0_outputs(12044)));
    outputs(11414) <= not(layer0_outputs(1546));
    outputs(11415) <= layer0_outputs(8519);
    outputs(11416) <= not(layer0_outputs(3558)) or (layer0_outputs(11022));
    outputs(11417) <= not((layer0_outputs(11740)) xor (layer0_outputs(12692)));
    outputs(11418) <= (layer0_outputs(11600)) or (layer0_outputs(12174));
    outputs(11419) <= (layer0_outputs(1420)) and not (layer0_outputs(10018));
    outputs(11420) <= '1';
    outputs(11421) <= layer0_outputs(6274);
    outputs(11422) <= (layer0_outputs(4316)) xor (layer0_outputs(5398));
    outputs(11423) <= layer0_outputs(8843);
    outputs(11424) <= not(layer0_outputs(8161)) or (layer0_outputs(3743));
    outputs(11425) <= layer0_outputs(8442);
    outputs(11426) <= not(layer0_outputs(10684));
    outputs(11427) <= not((layer0_outputs(11317)) xor (layer0_outputs(11444)));
    outputs(11428) <= layer0_outputs(3555);
    outputs(11429) <= layer0_outputs(5892);
    outputs(11430) <= (layer0_outputs(216)) or (layer0_outputs(1078));
    outputs(11431) <= (layer0_outputs(9290)) or (layer0_outputs(8844));
    outputs(11432) <= not(layer0_outputs(5820));
    outputs(11433) <= layer0_outputs(3600);
    outputs(11434) <= '1';
    outputs(11435) <= layer0_outputs(490);
    outputs(11436) <= not((layer0_outputs(1687)) or (layer0_outputs(2387)));
    outputs(11437) <= not((layer0_outputs(5222)) xor (layer0_outputs(8033)));
    outputs(11438) <= layer0_outputs(917);
    outputs(11439) <= (layer0_outputs(11470)) xor (layer0_outputs(2633));
    outputs(11440) <= not((layer0_outputs(3988)) xor (layer0_outputs(2281)));
    outputs(11441) <= layer0_outputs(3247);
    outputs(11442) <= (layer0_outputs(8746)) xor (layer0_outputs(9132));
    outputs(11443) <= (layer0_outputs(10135)) xor (layer0_outputs(10772));
    outputs(11444) <= layer0_outputs(5159);
    outputs(11445) <= not(layer0_outputs(3264));
    outputs(11446) <= (layer0_outputs(10863)) and (layer0_outputs(594));
    outputs(11447) <= not((layer0_outputs(176)) xor (layer0_outputs(2430)));
    outputs(11448) <= not(layer0_outputs(10066));
    outputs(11449) <= not(layer0_outputs(4368));
    outputs(11450) <= not(layer0_outputs(4505)) or (layer0_outputs(526));
    outputs(11451) <= (layer0_outputs(10828)) or (layer0_outputs(1800));
    outputs(11452) <= (layer0_outputs(4507)) and not (layer0_outputs(11628));
    outputs(11453) <= not((layer0_outputs(4467)) xor (layer0_outputs(8220)));
    outputs(11454) <= (layer0_outputs(8029)) xor (layer0_outputs(11133));
    outputs(11455) <= (layer0_outputs(4650)) xor (layer0_outputs(7620));
    outputs(11456) <= not(layer0_outputs(644));
    outputs(11457) <= not((layer0_outputs(6412)) xor (layer0_outputs(6198)));
    outputs(11458) <= layer0_outputs(12764);
    outputs(11459) <= not(layer0_outputs(5497));
    outputs(11460) <= not((layer0_outputs(1063)) and (layer0_outputs(2665)));
    outputs(11461) <= not(layer0_outputs(501));
    outputs(11462) <= not(layer0_outputs(4275));
    outputs(11463) <= (layer0_outputs(9583)) xor (layer0_outputs(12528));
    outputs(11464) <= not((layer0_outputs(1016)) xor (layer0_outputs(9006)));
    outputs(11465) <= (layer0_outputs(7688)) xor (layer0_outputs(10619));
    outputs(11466) <= layer0_outputs(12068);
    outputs(11467) <= not((layer0_outputs(1557)) xor (layer0_outputs(7192)));
    outputs(11468) <= not(layer0_outputs(10549));
    outputs(11469) <= not((layer0_outputs(4772)) or (layer0_outputs(3357)));
    outputs(11470) <= not((layer0_outputs(12473)) and (layer0_outputs(11668)));
    outputs(11471) <= not(layer0_outputs(769));
    outputs(11472) <= not(layer0_outputs(1082)) or (layer0_outputs(9814));
    outputs(11473) <= (layer0_outputs(6267)) xor (layer0_outputs(5920));
    outputs(11474) <= not((layer0_outputs(7131)) xor (layer0_outputs(10547)));
    outputs(11475) <= not(layer0_outputs(1718)) or (layer0_outputs(9815));
    outputs(11476) <= (layer0_outputs(5715)) xor (layer0_outputs(9516));
    outputs(11477) <= not(layer0_outputs(6650));
    outputs(11478) <= layer0_outputs(7703);
    outputs(11479) <= (layer0_outputs(2038)) and not (layer0_outputs(8546));
    outputs(11480) <= layer0_outputs(2831);
    outputs(11481) <= (layer0_outputs(10180)) and not (layer0_outputs(12668));
    outputs(11482) <= (layer0_outputs(2475)) xor (layer0_outputs(5573));
    outputs(11483) <= not((layer0_outputs(9468)) xor (layer0_outputs(7167)));
    outputs(11484) <= not((layer0_outputs(10236)) xor (layer0_outputs(9922)));
    outputs(11485) <= not(layer0_outputs(1860)) or (layer0_outputs(1962));
    outputs(11486) <= (layer0_outputs(947)) xor (layer0_outputs(12639));
    outputs(11487) <= (layer0_outputs(5895)) or (layer0_outputs(4214));
    outputs(11488) <= layer0_outputs(10599);
    outputs(11489) <= '0';
    outputs(11490) <= not(layer0_outputs(10252));
    outputs(11491) <= not((layer0_outputs(6810)) or (layer0_outputs(2577)));
    outputs(11492) <= (layer0_outputs(9922)) xor (layer0_outputs(3164));
    outputs(11493) <= not((layer0_outputs(7669)) or (layer0_outputs(12776)));
    outputs(11494) <= not(layer0_outputs(1382));
    outputs(11495) <= layer0_outputs(1375);
    outputs(11496) <= (layer0_outputs(4673)) xor (layer0_outputs(6820));
    outputs(11497) <= layer0_outputs(5242);
    outputs(11498) <= not(layer0_outputs(7767));
    outputs(11499) <= not(layer0_outputs(12503));
    outputs(11500) <= not((layer0_outputs(11616)) xor (layer0_outputs(7580)));
    outputs(11501) <= layer0_outputs(7664);
    outputs(11502) <= not((layer0_outputs(11598)) xor (layer0_outputs(7358)));
    outputs(11503) <= layer0_outputs(5039);
    outputs(11504) <= not((layer0_outputs(11578)) xor (layer0_outputs(7064)));
    outputs(11505) <= layer0_outputs(11733);
    outputs(11506) <= not((layer0_outputs(11315)) xor (layer0_outputs(12179)));
    outputs(11507) <= not(layer0_outputs(1876)) or (layer0_outputs(985));
    outputs(11508) <= not(layer0_outputs(8331));
    outputs(11509) <= not(layer0_outputs(2207));
    outputs(11510) <= not((layer0_outputs(8732)) xor (layer0_outputs(10626)));
    outputs(11511) <= (layer0_outputs(10255)) xor (layer0_outputs(1964));
    outputs(11512) <= (layer0_outputs(2672)) xor (layer0_outputs(12212));
    outputs(11513) <= (layer0_outputs(3933)) and not (layer0_outputs(10683));
    outputs(11514) <= layer0_outputs(10014);
    outputs(11515) <= not((layer0_outputs(629)) and (layer0_outputs(10581)));
    outputs(11516) <= not(layer0_outputs(6886)) or (layer0_outputs(3354));
    outputs(11517) <= not((layer0_outputs(4360)) xor (layer0_outputs(5039)));
    outputs(11518) <= not((layer0_outputs(12070)) xor (layer0_outputs(4395)));
    outputs(11519) <= not((layer0_outputs(8138)) xor (layer0_outputs(9480)));
    outputs(11520) <= (layer0_outputs(10759)) and not (layer0_outputs(11261));
    outputs(11521) <= not(layer0_outputs(3449));
    outputs(11522) <= not(layer0_outputs(7633));
    outputs(11523) <= (layer0_outputs(8633)) and not (layer0_outputs(4958));
    outputs(11524) <= (layer0_outputs(4474)) and not (layer0_outputs(9195));
    outputs(11525) <= not(layer0_outputs(9000));
    outputs(11526) <= layer0_outputs(267);
    outputs(11527) <= (layer0_outputs(2781)) xor (layer0_outputs(2116));
    outputs(11528) <= layer0_outputs(1029);
    outputs(11529) <= (layer0_outputs(5893)) and (layer0_outputs(4714));
    outputs(11530) <= layer0_outputs(12151);
    outputs(11531) <= (layer0_outputs(3580)) and (layer0_outputs(11382));
    outputs(11532) <= not(layer0_outputs(9057));
    outputs(11533) <= not(layer0_outputs(9872)) or (layer0_outputs(8421));
    outputs(11534) <= layer0_outputs(1323);
    outputs(11535) <= not((layer0_outputs(9857)) xor (layer0_outputs(9114)));
    outputs(11536) <= layer0_outputs(6006);
    outputs(11537) <= not(layer0_outputs(6200));
    outputs(11538) <= not(layer0_outputs(6936)) or (layer0_outputs(10149));
    outputs(11539) <= (layer0_outputs(5380)) xor (layer0_outputs(3751));
    outputs(11540) <= not(layer0_outputs(9756)) or (layer0_outputs(4677));
    outputs(11541) <= (layer0_outputs(12094)) xor (layer0_outputs(9356));
    outputs(11542) <= layer0_outputs(4815);
    outputs(11543) <= not((layer0_outputs(8313)) xor (layer0_outputs(3658)));
    outputs(11544) <= (layer0_outputs(799)) xor (layer0_outputs(6424));
    outputs(11545) <= (layer0_outputs(9013)) xor (layer0_outputs(9923));
    outputs(11546) <= not((layer0_outputs(3622)) or (layer0_outputs(2710)));
    outputs(11547) <= layer0_outputs(3366);
    outputs(11548) <= (layer0_outputs(2394)) xor (layer0_outputs(9245));
    outputs(11549) <= (layer0_outputs(11009)) and not (layer0_outputs(9649));
    outputs(11550) <= (layer0_outputs(5407)) xor (layer0_outputs(11452));
    outputs(11551) <= (layer0_outputs(8131)) xor (layer0_outputs(6190));
    outputs(11552) <= (layer0_outputs(4590)) and not (layer0_outputs(5471));
    outputs(11553) <= (layer0_outputs(270)) and not (layer0_outputs(12779));
    outputs(11554) <= not((layer0_outputs(8073)) or (layer0_outputs(7202)));
    outputs(11555) <= not(layer0_outputs(5587));
    outputs(11556) <= not((layer0_outputs(12105)) xor (layer0_outputs(11511)));
    outputs(11557) <= not((layer0_outputs(10710)) xor (layer0_outputs(277)));
    outputs(11558) <= not((layer0_outputs(6196)) xor (layer0_outputs(1414)));
    outputs(11559) <= (layer0_outputs(10936)) and (layer0_outputs(7230));
    outputs(11560) <= (layer0_outputs(1483)) xor (layer0_outputs(4846));
    outputs(11561) <= layer0_outputs(984);
    outputs(11562) <= (layer0_outputs(9685)) xor (layer0_outputs(781));
    outputs(11563) <= layer0_outputs(7166);
    outputs(11564) <= not((layer0_outputs(12539)) xor (layer0_outputs(2158)));
    outputs(11565) <= not(layer0_outputs(10859));
    outputs(11566) <= (layer0_outputs(7875)) xor (layer0_outputs(3854));
    outputs(11567) <= not(layer0_outputs(12267));
    outputs(11568) <= (layer0_outputs(2973)) and not (layer0_outputs(7091));
    outputs(11569) <= layer0_outputs(1307);
    outputs(11570) <= not(layer0_outputs(4041));
    outputs(11571) <= (layer0_outputs(10079)) and not (layer0_outputs(5886));
    outputs(11572) <= not(layer0_outputs(6329));
    outputs(11573) <= not((layer0_outputs(3838)) xor (layer0_outputs(4754)));
    outputs(11574) <= (layer0_outputs(9709)) and (layer0_outputs(7548));
    outputs(11575) <= not(layer0_outputs(7519));
    outputs(11576) <= layer0_outputs(5135);
    outputs(11577) <= not((layer0_outputs(3317)) or (layer0_outputs(11325)));
    outputs(11578) <= layer0_outputs(12665);
    outputs(11579) <= not((layer0_outputs(3837)) xor (layer0_outputs(11816)));
    outputs(11580) <= not((layer0_outputs(12313)) xor (layer0_outputs(5941)));
    outputs(11581) <= not(layer0_outputs(11369));
    outputs(11582) <= (layer0_outputs(6258)) and (layer0_outputs(1935));
    outputs(11583) <= layer0_outputs(11715);
    outputs(11584) <= not(layer0_outputs(254)) or (layer0_outputs(11635));
    outputs(11585) <= not(layer0_outputs(4512));
    outputs(11586) <= layer0_outputs(9370);
    outputs(11587) <= not((layer0_outputs(12437)) xor (layer0_outputs(11090)));
    outputs(11588) <= (layer0_outputs(6311)) and (layer0_outputs(4610));
    outputs(11589) <= (layer0_outputs(1347)) and not (layer0_outputs(4375));
    outputs(11590) <= (layer0_outputs(11475)) and (layer0_outputs(437));
    outputs(11591) <= layer0_outputs(10661);
    outputs(11592) <= (layer0_outputs(603)) xor (layer0_outputs(3986));
    outputs(11593) <= not((layer0_outputs(2540)) xor (layer0_outputs(680)));
    outputs(11594) <= not((layer0_outputs(7662)) xor (layer0_outputs(959)));
    outputs(11595) <= (layer0_outputs(12310)) xor (layer0_outputs(3677));
    outputs(11596) <= (layer0_outputs(2177)) xor (layer0_outputs(7057));
    outputs(11597) <= layer0_outputs(7612);
    outputs(11598) <= not((layer0_outputs(1035)) xor (layer0_outputs(4062)));
    outputs(11599) <= (layer0_outputs(7316)) and not (layer0_outputs(6751));
    outputs(11600) <= (layer0_outputs(4384)) xor (layer0_outputs(753));
    outputs(11601) <= (layer0_outputs(9024)) and not (layer0_outputs(12400));
    outputs(11602) <= not((layer0_outputs(6410)) xor (layer0_outputs(4308)));
    outputs(11603) <= not(layer0_outputs(10373));
    outputs(11604) <= (layer0_outputs(1991)) xor (layer0_outputs(7248));
    outputs(11605) <= not((layer0_outputs(8545)) xor (layer0_outputs(7018)));
    outputs(11606) <= not(layer0_outputs(8964));
    outputs(11607) <= not((layer0_outputs(4073)) xor (layer0_outputs(1706)));
    outputs(11608) <= layer0_outputs(12227);
    outputs(11609) <= (layer0_outputs(339)) xor (layer0_outputs(10318));
    outputs(11610) <= not((layer0_outputs(12439)) xor (layer0_outputs(4721)));
    outputs(11611) <= not((layer0_outputs(5462)) xor (layer0_outputs(9842)));
    outputs(11612) <= (layer0_outputs(10107)) and not (layer0_outputs(5370));
    outputs(11613) <= (layer0_outputs(4903)) and (layer0_outputs(9960));
    outputs(11614) <= layer0_outputs(3872);
    outputs(11615) <= layer0_outputs(10214);
    outputs(11616) <= not(layer0_outputs(4418));
    outputs(11617) <= not(layer0_outputs(7814));
    outputs(11618) <= layer0_outputs(5109);
    outputs(11619) <= not((layer0_outputs(12377)) or (layer0_outputs(2371)));
    outputs(11620) <= not(layer0_outputs(566));
    outputs(11621) <= not((layer0_outputs(2830)) xor (layer0_outputs(8357)));
    outputs(11622) <= (layer0_outputs(9558)) xor (layer0_outputs(6729));
    outputs(11623) <= (layer0_outputs(4744)) xor (layer0_outputs(3456));
    outputs(11624) <= not((layer0_outputs(3356)) xor (layer0_outputs(8053)));
    outputs(11625) <= not(layer0_outputs(3102));
    outputs(11626) <= (layer0_outputs(6072)) xor (layer0_outputs(5432));
    outputs(11627) <= not(layer0_outputs(4005));
    outputs(11628) <= not(layer0_outputs(12781));
    outputs(11629) <= not(layer0_outputs(3968));
    outputs(11630) <= (layer0_outputs(9946)) and not (layer0_outputs(10261));
    outputs(11631) <= layer0_outputs(11817);
    outputs(11632) <= (layer0_outputs(1812)) and (layer0_outputs(4628));
    outputs(11633) <= (layer0_outputs(9971)) xor (layer0_outputs(8474));
    outputs(11634) <= not(layer0_outputs(4030));
    outputs(11635) <= (layer0_outputs(10664)) xor (layer0_outputs(12339));
    outputs(11636) <= layer0_outputs(7822);
    outputs(11637) <= '0';
    outputs(11638) <= not(layer0_outputs(2909)) or (layer0_outputs(4669));
    outputs(11639) <= (layer0_outputs(9857)) xor (layer0_outputs(6692));
    outputs(11640) <= not((layer0_outputs(9352)) or (layer0_outputs(4653)));
    outputs(11641) <= (layer0_outputs(7409)) and not (layer0_outputs(1971));
    outputs(11642) <= layer0_outputs(6168);
    outputs(11643) <= not(layer0_outputs(6210)) or (layer0_outputs(362));
    outputs(11644) <= not((layer0_outputs(2118)) xor (layer0_outputs(5310)));
    outputs(11645) <= (layer0_outputs(10362)) xor (layer0_outputs(5325));
    outputs(11646) <= layer0_outputs(8653);
    outputs(11647) <= not(layer0_outputs(8030)) or (layer0_outputs(6699));
    outputs(11648) <= layer0_outputs(4699);
    outputs(11649) <= layer0_outputs(3943);
    outputs(11650) <= not(layer0_outputs(2325));
    outputs(11651) <= layer0_outputs(5110);
    outputs(11652) <= layer0_outputs(8203);
    outputs(11653) <= (layer0_outputs(1854)) and (layer0_outputs(8607));
    outputs(11654) <= not(layer0_outputs(1397));
    outputs(11655) <= layer0_outputs(817);
    outputs(11656) <= layer0_outputs(2466);
    outputs(11657) <= (layer0_outputs(4364)) xor (layer0_outputs(3086));
    outputs(11658) <= not((layer0_outputs(3525)) xor (layer0_outputs(11115)));
    outputs(11659) <= not((layer0_outputs(10305)) or (layer0_outputs(10477)));
    outputs(11660) <= (layer0_outputs(4342)) and (layer0_outputs(12734));
    outputs(11661) <= not((layer0_outputs(8524)) or (layer0_outputs(7208)));
    outputs(11662) <= not(layer0_outputs(9472));
    outputs(11663) <= not(layer0_outputs(9819));
    outputs(11664) <= layer0_outputs(2883);
    outputs(11665) <= layer0_outputs(7280);
    outputs(11666) <= not(layer0_outputs(4882));
    outputs(11667) <= not((layer0_outputs(4657)) xor (layer0_outputs(6832)));
    outputs(11668) <= not((layer0_outputs(7631)) xor (layer0_outputs(8380)));
    outputs(11669) <= not(layer0_outputs(2455));
    outputs(11670) <= not(layer0_outputs(1912));
    outputs(11671) <= layer0_outputs(3155);
    outputs(11672) <= '1';
    outputs(11673) <= (layer0_outputs(6022)) and not (layer0_outputs(2142));
    outputs(11674) <= not(layer0_outputs(4734));
    outputs(11675) <= not((layer0_outputs(3688)) xor (layer0_outputs(8352)));
    outputs(11676) <= not((layer0_outputs(12189)) xor (layer0_outputs(2897)));
    outputs(11677) <= layer0_outputs(8069);
    outputs(11678) <= layer0_outputs(930);
    outputs(11679) <= not(layer0_outputs(4811));
    outputs(11680) <= layer0_outputs(3165);
    outputs(11681) <= not((layer0_outputs(11738)) xor (layer0_outputs(3726)));
    outputs(11682) <= not(layer0_outputs(4447)) or (layer0_outputs(4587));
    outputs(11683) <= layer0_outputs(8489);
    outputs(11684) <= not((layer0_outputs(1946)) and (layer0_outputs(291)));
    outputs(11685) <= (layer0_outputs(2887)) and not (layer0_outputs(10594));
    outputs(11686) <= not(layer0_outputs(837));
    outputs(11687) <= layer0_outputs(9623);
    outputs(11688) <= (layer0_outputs(2217)) and not (layer0_outputs(9599));
    outputs(11689) <= (layer0_outputs(2414)) xor (layer0_outputs(1813));
    outputs(11690) <= (layer0_outputs(4199)) xor (layer0_outputs(1208));
    outputs(11691) <= layer0_outputs(12287);
    outputs(11692) <= (layer0_outputs(8711)) xor (layer0_outputs(12337));
    outputs(11693) <= not(layer0_outputs(3374));
    outputs(11694) <= layer0_outputs(5838);
    outputs(11695) <= (layer0_outputs(9040)) xor (layer0_outputs(3640));
    outputs(11696) <= '0';
    outputs(11697) <= not(layer0_outputs(8709));
    outputs(11698) <= not(layer0_outputs(3895));
    outputs(11699) <= not((layer0_outputs(2878)) or (layer0_outputs(1162)));
    outputs(11700) <= (layer0_outputs(6172)) xor (layer0_outputs(11284));
    outputs(11701) <= layer0_outputs(5335);
    outputs(11702) <= layer0_outputs(6847);
    outputs(11703) <= not(layer0_outputs(4362));
    outputs(11704) <= not(layer0_outputs(12489));
    outputs(11705) <= (layer0_outputs(999)) xor (layer0_outputs(4435));
    outputs(11706) <= not((layer0_outputs(7431)) xor (layer0_outputs(8468)));
    outputs(11707) <= (layer0_outputs(1650)) and not (layer0_outputs(8275));
    outputs(11708) <= (layer0_outputs(4094)) and (layer0_outputs(1822));
    outputs(11709) <= not(layer0_outputs(1032));
    outputs(11710) <= not((layer0_outputs(5435)) or (layer0_outputs(3454)));
    outputs(11711) <= (layer0_outputs(4210)) xor (layer0_outputs(3060));
    outputs(11712) <= (layer0_outputs(999)) and not (layer0_outputs(8465));
    outputs(11713) <= not(layer0_outputs(5827));
    outputs(11714) <= (layer0_outputs(9055)) xor (layer0_outputs(1320));
    outputs(11715) <= (layer0_outputs(1956)) and not (layer0_outputs(2963));
    outputs(11716) <= not((layer0_outputs(6059)) or (layer0_outputs(11136)));
    outputs(11717) <= not(layer0_outputs(2589));
    outputs(11718) <= (layer0_outputs(1593)) or (layer0_outputs(7953));
    outputs(11719) <= layer0_outputs(8840);
    outputs(11720) <= not(layer0_outputs(2498));
    outputs(11721) <= not(layer0_outputs(2863));
    outputs(11722) <= layer0_outputs(9106);
    outputs(11723) <= not((layer0_outputs(6147)) or (layer0_outputs(163)));
    outputs(11724) <= not(layer0_outputs(5368));
    outputs(11725) <= not(layer0_outputs(10243));
    outputs(11726) <= (layer0_outputs(10716)) or (layer0_outputs(2573));
    outputs(11727) <= (layer0_outputs(768)) and not (layer0_outputs(6529));
    outputs(11728) <= layer0_outputs(9335);
    outputs(11729) <= (layer0_outputs(5759)) and (layer0_outputs(841));
    outputs(11730) <= (layer0_outputs(4872)) and not (layer0_outputs(9432));
    outputs(11731) <= layer0_outputs(12676);
    outputs(11732) <= not((layer0_outputs(74)) and (layer0_outputs(6601)));
    outputs(11733) <= layer0_outputs(4700);
    outputs(11734) <= '1';
    outputs(11735) <= (layer0_outputs(9412)) xor (layer0_outputs(7492));
    outputs(11736) <= (layer0_outputs(1576)) or (layer0_outputs(925));
    outputs(11737) <= (layer0_outputs(9149)) and not (layer0_outputs(1505));
    outputs(11738) <= (layer0_outputs(7748)) and not (layer0_outputs(3211));
    outputs(11739) <= (layer0_outputs(1467)) xor (layer0_outputs(7268));
    outputs(11740) <= (layer0_outputs(3944)) xor (layer0_outputs(3523));
    outputs(11741) <= not((layer0_outputs(6076)) xor (layer0_outputs(7887)));
    outputs(11742) <= not(layer0_outputs(696));
    outputs(11743) <= not((layer0_outputs(4578)) or (layer0_outputs(10071)));
    outputs(11744) <= (layer0_outputs(7893)) or (layer0_outputs(2082));
    outputs(11745) <= layer0_outputs(6180);
    outputs(11746) <= layer0_outputs(2403);
    outputs(11747) <= not((layer0_outputs(7057)) xor (layer0_outputs(2973)));
    outputs(11748) <= not(layer0_outputs(7965));
    outputs(11749) <= not((layer0_outputs(10586)) or (layer0_outputs(11914)));
    outputs(11750) <= not(layer0_outputs(12740));
    outputs(11751) <= (layer0_outputs(7421)) and (layer0_outputs(5922));
    outputs(11752) <= layer0_outputs(3806);
    outputs(11753) <= not(layer0_outputs(986));
    outputs(11754) <= not((layer0_outputs(1463)) xor (layer0_outputs(3748)));
    outputs(11755) <= (layer0_outputs(4411)) and not (layer0_outputs(12363));
    outputs(11756) <= not((layer0_outputs(8036)) xor (layer0_outputs(9244)));
    outputs(11757) <= (layer0_outputs(2184)) and not (layer0_outputs(10742));
    outputs(11758) <= '1';
    outputs(11759) <= (layer0_outputs(8784)) xor (layer0_outputs(11993));
    outputs(11760) <= not(layer0_outputs(7468));
    outputs(11761) <= (layer0_outputs(5601)) and not (layer0_outputs(5615));
    outputs(11762) <= layer0_outputs(8459);
    outputs(11763) <= not((layer0_outputs(228)) or (layer0_outputs(6495)));
    outputs(11764) <= not((layer0_outputs(3694)) xor (layer0_outputs(9801)));
    outputs(11765) <= layer0_outputs(2885);
    outputs(11766) <= layer0_outputs(2495);
    outputs(11767) <= (layer0_outputs(5625)) and not (layer0_outputs(4142));
    outputs(11768) <= layer0_outputs(3915);
    outputs(11769) <= (layer0_outputs(4481)) xor (layer0_outputs(1555));
    outputs(11770) <= (layer0_outputs(2274)) and (layer0_outputs(9428));
    outputs(11771) <= layer0_outputs(8774);
    outputs(11772) <= layer0_outputs(3172);
    outputs(11773) <= (layer0_outputs(8783)) and not (layer0_outputs(4695));
    outputs(11774) <= not(layer0_outputs(6634));
    outputs(11775) <= layer0_outputs(3993);
    outputs(11776) <= layer0_outputs(6088);
    outputs(11777) <= not(layer0_outputs(8231));
    outputs(11778) <= not(layer0_outputs(5092)) or (layer0_outputs(10810));
    outputs(11779) <= (layer0_outputs(11542)) xor (layer0_outputs(1199));
    outputs(11780) <= not((layer0_outputs(6878)) xor (layer0_outputs(7142)));
    outputs(11781) <= not(layer0_outputs(471));
    outputs(11782) <= layer0_outputs(5324);
    outputs(11783) <= not(layer0_outputs(3574));
    outputs(11784) <= not((layer0_outputs(776)) xor (layer0_outputs(12039)));
    outputs(11785) <= layer0_outputs(3379);
    outputs(11786) <= not((layer0_outputs(7147)) or (layer0_outputs(593)));
    outputs(11787) <= not((layer0_outputs(8759)) or (layer0_outputs(11212)));
    outputs(11788) <= not((layer0_outputs(8269)) xor (layer0_outputs(3231)));
    outputs(11789) <= not((layer0_outputs(12413)) xor (layer0_outputs(414)));
    outputs(11790) <= not((layer0_outputs(4984)) xor (layer0_outputs(8796)));
    outputs(11791) <= layer0_outputs(1560);
    outputs(11792) <= (layer0_outputs(5019)) and not (layer0_outputs(8439));
    outputs(11793) <= (layer0_outputs(7598)) xor (layer0_outputs(7241));
    outputs(11794) <= layer0_outputs(10492);
    outputs(11795) <= not((layer0_outputs(11262)) xor (layer0_outputs(1325)));
    outputs(11796) <= not((layer0_outputs(8012)) xor (layer0_outputs(8919)));
    outputs(11797) <= not(layer0_outputs(1429)) or (layer0_outputs(7460));
    outputs(11798) <= not(layer0_outputs(5526)) or (layer0_outputs(8688));
    outputs(11799) <= (layer0_outputs(4152)) xor (layer0_outputs(10809));
    outputs(11800) <= not(layer0_outputs(6904)) or (layer0_outputs(11972));
    outputs(11801) <= not(layer0_outputs(7397));
    outputs(11802) <= (layer0_outputs(120)) and not (layer0_outputs(3103));
    outputs(11803) <= layer0_outputs(8042);
    outputs(11804) <= (layer0_outputs(5018)) and not (layer0_outputs(8));
    outputs(11805) <= layer0_outputs(9255);
    outputs(11806) <= not(layer0_outputs(3787)) or (layer0_outputs(1057));
    outputs(11807) <= (layer0_outputs(7405)) xor (layer0_outputs(9895));
    outputs(11808) <= not(layer0_outputs(7737));
    outputs(11809) <= '0';
    outputs(11810) <= (layer0_outputs(10031)) and not (layer0_outputs(7761));
    outputs(11811) <= layer0_outputs(3042);
    outputs(11812) <= not(layer0_outputs(8460));
    outputs(11813) <= layer0_outputs(12730);
    outputs(11814) <= not(layer0_outputs(11973));
    outputs(11815) <= not(layer0_outputs(5741)) or (layer0_outputs(1184));
    outputs(11816) <= (layer0_outputs(4651)) xor (layer0_outputs(2948));
    outputs(11817) <= not(layer0_outputs(12584));
    outputs(11818) <= '0';
    outputs(11819) <= not((layer0_outputs(7001)) or (layer0_outputs(2467)));
    outputs(11820) <= not(layer0_outputs(611));
    outputs(11821) <= layer0_outputs(7310);
    outputs(11822) <= not((layer0_outputs(10278)) or (layer0_outputs(7422)));
    outputs(11823) <= not((layer0_outputs(3924)) xor (layer0_outputs(4802)));
    outputs(11824) <= layer0_outputs(4231);
    outputs(11825) <= layer0_outputs(10610);
    outputs(11826) <= not(layer0_outputs(329));
    outputs(11827) <= layer0_outputs(5857);
    outputs(11828) <= layer0_outputs(3393);
    outputs(11829) <= not(layer0_outputs(3044));
    outputs(11830) <= layer0_outputs(7393);
    outputs(11831) <= layer0_outputs(3887);
    outputs(11832) <= layer0_outputs(2578);
    outputs(11833) <= not((layer0_outputs(4753)) and (layer0_outputs(3918)));
    outputs(11834) <= layer0_outputs(8549);
    outputs(11835) <= (layer0_outputs(8446)) and (layer0_outputs(6558));
    outputs(11836) <= not((layer0_outputs(2684)) and (layer0_outputs(9186)));
    outputs(11837) <= layer0_outputs(10224);
    outputs(11838) <= not(layer0_outputs(2112));
    outputs(11839) <= not((layer0_outputs(11170)) xor (layer0_outputs(12109)));
    outputs(11840) <= (layer0_outputs(3792)) xor (layer0_outputs(5752));
    outputs(11841) <= layer0_outputs(6451);
    outputs(11842) <= (layer0_outputs(8025)) xor (layer0_outputs(10008));
    outputs(11843) <= layer0_outputs(1297);
    outputs(11844) <= not(layer0_outputs(12415));
    outputs(11845) <= layer0_outputs(4471);
    outputs(11846) <= (layer0_outputs(12484)) xor (layer0_outputs(4455));
    outputs(11847) <= layer0_outputs(7835);
    outputs(11848) <= layer0_outputs(6199);
    outputs(11849) <= (layer0_outputs(10516)) and (layer0_outputs(9023));
    outputs(11850) <= not(layer0_outputs(7136));
    outputs(11851) <= (layer0_outputs(11845)) and not (layer0_outputs(12478));
    outputs(11852) <= not((layer0_outputs(3171)) or (layer0_outputs(4681)));
    outputs(11853) <= (layer0_outputs(8547)) and not (layer0_outputs(1360));
    outputs(11854) <= layer0_outputs(2023);
    outputs(11855) <= not(layer0_outputs(5229));
    outputs(11856) <= not((layer0_outputs(7149)) xor (layer0_outputs(11168)));
    outputs(11857) <= layer0_outputs(11406);
    outputs(11858) <= not((layer0_outputs(12758)) xor (layer0_outputs(10929)));
    outputs(11859) <= layer0_outputs(950);
    outputs(11860) <= layer0_outputs(6003);
    outputs(11861) <= not(layer0_outputs(180));
    outputs(11862) <= (layer0_outputs(1644)) xor (layer0_outputs(3858));
    outputs(11863) <= not((layer0_outputs(4907)) and (layer0_outputs(8915)));
    outputs(11864) <= layer0_outputs(6011);
    outputs(11865) <= (layer0_outputs(10198)) xor (layer0_outputs(7798));
    outputs(11866) <= not(layer0_outputs(4803)) or (layer0_outputs(4565));
    outputs(11867) <= layer0_outputs(11539);
    outputs(11868) <= (layer0_outputs(4194)) and (layer0_outputs(6609));
    outputs(11869) <= (layer0_outputs(11800)) and (layer0_outputs(5378));
    outputs(11870) <= not(layer0_outputs(10990));
    outputs(11871) <= not(layer0_outputs(7492));
    outputs(11872) <= not(layer0_outputs(12098));
    outputs(11873) <= not(layer0_outputs(12125));
    outputs(11874) <= not((layer0_outputs(8306)) xor (layer0_outputs(9127)));
    outputs(11875) <= not(layer0_outputs(11213));
    outputs(11876) <= (layer0_outputs(12617)) xor (layer0_outputs(9679));
    outputs(11877) <= (layer0_outputs(7611)) xor (layer0_outputs(10794));
    outputs(11878) <= not((layer0_outputs(3329)) and (layer0_outputs(3151)));
    outputs(11879) <= not(layer0_outputs(1172));
    outputs(11880) <= not(layer0_outputs(529)) or (layer0_outputs(2562));
    outputs(11881) <= (layer0_outputs(10259)) and (layer0_outputs(12131));
    outputs(11882) <= (layer0_outputs(6928)) xor (layer0_outputs(478));
    outputs(11883) <= layer0_outputs(4222);
    outputs(11884) <= (layer0_outputs(3744)) xor (layer0_outputs(9684));
    outputs(11885) <= not(layer0_outputs(5586));
    outputs(11886) <= (layer0_outputs(11417)) xor (layer0_outputs(7163));
    outputs(11887) <= not(layer0_outputs(2456));
    outputs(11888) <= (layer0_outputs(10496)) xor (layer0_outputs(5782));
    outputs(11889) <= not(layer0_outputs(3217));
    outputs(11890) <= layer0_outputs(2356);
    outputs(11891) <= not(layer0_outputs(2989));
    outputs(11892) <= layer0_outputs(12079);
    outputs(11893) <= not(layer0_outputs(4556));
    outputs(11894) <= not((layer0_outputs(471)) and (layer0_outputs(3851)));
    outputs(11895) <= not(layer0_outputs(269));
    outputs(11896) <= not(layer0_outputs(10310));
    outputs(11897) <= not((layer0_outputs(2273)) xor (layer0_outputs(11142)));
    outputs(11898) <= (layer0_outputs(8236)) xor (layer0_outputs(11438));
    outputs(11899) <= not((layer0_outputs(7420)) xor (layer0_outputs(10245)));
    outputs(11900) <= (layer0_outputs(5009)) and not (layer0_outputs(4280));
    outputs(11901) <= not(layer0_outputs(8937));
    outputs(11902) <= not((layer0_outputs(4185)) or (layer0_outputs(8152)));
    outputs(11903) <= (layer0_outputs(8783)) xor (layer0_outputs(526));
    outputs(11904) <= not((layer0_outputs(50)) xor (layer0_outputs(11454)));
    outputs(11905) <= layer0_outputs(7457);
    outputs(11906) <= (layer0_outputs(7232)) xor (layer0_outputs(4236));
    outputs(11907) <= not(layer0_outputs(3972));
    outputs(11908) <= (layer0_outputs(7020)) xor (layer0_outputs(12706));
    outputs(11909) <= (layer0_outputs(10772)) and not (layer0_outputs(918));
    outputs(11910) <= not(layer0_outputs(564));
    outputs(11911) <= '0';
    outputs(11912) <= (layer0_outputs(1733)) and not (layer0_outputs(12520));
    outputs(11913) <= not((layer0_outputs(1652)) xor (layer0_outputs(8970)));
    outputs(11914) <= (layer0_outputs(1749)) and (layer0_outputs(1871));
    outputs(11915) <= (layer0_outputs(2546)) and (layer0_outputs(6573));
    outputs(11916) <= not(layer0_outputs(5631));
    outputs(11917) <= not((layer0_outputs(5114)) xor (layer0_outputs(5619)));
    outputs(11918) <= (layer0_outputs(5071)) and not (layer0_outputs(7859));
    outputs(11919) <= not(layer0_outputs(531)) or (layer0_outputs(11564));
    outputs(11920) <= (layer0_outputs(5226)) and (layer0_outputs(7183));
    outputs(11921) <= not((layer0_outputs(518)) xor (layer0_outputs(9118)));
    outputs(11922) <= not(layer0_outputs(2467));
    outputs(11923) <= layer0_outputs(1265);
    outputs(11924) <= (layer0_outputs(234)) xor (layer0_outputs(12289));
    outputs(11925) <= not((layer0_outputs(8512)) or (layer0_outputs(835)));
    outputs(11926) <= (layer0_outputs(11308)) xor (layer0_outputs(3274));
    outputs(11927) <= not((layer0_outputs(6460)) xor (layer0_outputs(10419)));
    outputs(11928) <= (layer0_outputs(9046)) xor (layer0_outputs(4600));
    outputs(11929) <= not((layer0_outputs(6965)) xor (layer0_outputs(2051)));
    outputs(11930) <= (layer0_outputs(186)) xor (layer0_outputs(891));
    outputs(11931) <= (layer0_outputs(10889)) and not (layer0_outputs(12564));
    outputs(11932) <= (layer0_outputs(11444)) and (layer0_outputs(5224));
    outputs(11933) <= (layer0_outputs(914)) and not (layer0_outputs(6372));
    outputs(11934) <= layer0_outputs(1259);
    outputs(11935) <= layer0_outputs(6456);
    outputs(11936) <= (layer0_outputs(12548)) xor (layer0_outputs(2389));
    outputs(11937) <= layer0_outputs(11241);
    outputs(11938) <= not(layer0_outputs(4479));
    outputs(11939) <= layer0_outputs(3407);
    outputs(11940) <= (layer0_outputs(613)) xor (layer0_outputs(6892));
    outputs(11941) <= layer0_outputs(9058);
    outputs(11942) <= (layer0_outputs(9578)) and (layer0_outputs(4002));
    outputs(11943) <= not(layer0_outputs(2717));
    outputs(11944) <= layer0_outputs(6588);
    outputs(11945) <= layer0_outputs(1363);
    outputs(11946) <= layer0_outputs(4623);
    outputs(11947) <= not((layer0_outputs(3677)) and (layer0_outputs(5848)));
    outputs(11948) <= layer0_outputs(6180);
    outputs(11949) <= layer0_outputs(2249);
    outputs(11950) <= layer0_outputs(8740);
    outputs(11951) <= not((layer0_outputs(6620)) xor (layer0_outputs(3772)));
    outputs(11952) <= not((layer0_outputs(2092)) xor (layer0_outputs(4525)));
    outputs(11953) <= not(layer0_outputs(1009)) or (layer0_outputs(7377));
    outputs(11954) <= (layer0_outputs(6308)) xor (layer0_outputs(1315));
    outputs(11955) <= (layer0_outputs(3699)) and not (layer0_outputs(9150));
    outputs(11956) <= layer0_outputs(2181);
    outputs(11957) <= not(layer0_outputs(5085));
    outputs(11958) <= not((layer0_outputs(4660)) xor (layer0_outputs(301)));
    outputs(11959) <= not(layer0_outputs(7306));
    outputs(11960) <= (layer0_outputs(1533)) xor (layer0_outputs(1155));
    outputs(11961) <= layer0_outputs(4007);
    outputs(11962) <= layer0_outputs(5935);
    outputs(11963) <= not((layer0_outputs(2758)) or (layer0_outputs(4813)));
    outputs(11964) <= not(layer0_outputs(3128));
    outputs(11965) <= (layer0_outputs(6396)) xor (layer0_outputs(2361));
    outputs(11966) <= not(layer0_outputs(10286));
    outputs(11967) <= not(layer0_outputs(7566));
    outputs(11968) <= not((layer0_outputs(8704)) xor (layer0_outputs(4032)));
    outputs(11969) <= not((layer0_outputs(7441)) xor (layer0_outputs(2931)));
    outputs(11970) <= (layer0_outputs(5384)) xor (layer0_outputs(10926));
    outputs(11971) <= not((layer0_outputs(8592)) xor (layer0_outputs(7641)));
    outputs(11972) <= layer0_outputs(4111);
    outputs(11973) <= layer0_outputs(8065);
    outputs(11974) <= not(layer0_outputs(10913)) or (layer0_outputs(10618));
    outputs(11975) <= not(layer0_outputs(1267));
    outputs(11976) <= layer0_outputs(4618);
    outputs(11977) <= layer0_outputs(8993);
    outputs(11978) <= not((layer0_outputs(4712)) xor (layer0_outputs(1832)));
    outputs(11979) <= not((layer0_outputs(3713)) xor (layer0_outputs(3554)));
    outputs(11980) <= (layer0_outputs(2533)) xor (layer0_outputs(11950));
    outputs(11981) <= not((layer0_outputs(3960)) and (layer0_outputs(10877)));
    outputs(11982) <= not((layer0_outputs(209)) xor (layer0_outputs(11231)));
    outputs(11983) <= not((layer0_outputs(2057)) xor (layer0_outputs(4793)));
    outputs(11984) <= not(layer0_outputs(3589));
    outputs(11985) <= layer0_outputs(8272);
    outputs(11986) <= not(layer0_outputs(10186));
    outputs(11987) <= not(layer0_outputs(41));
    outputs(11988) <= (layer0_outputs(4552)) and not (layer0_outputs(10575));
    outputs(11989) <= not(layer0_outputs(3320));
    outputs(11990) <= (layer0_outputs(3057)) xor (layer0_outputs(2306));
    outputs(11991) <= (layer0_outputs(1244)) xor (layer0_outputs(4189));
    outputs(11992) <= not((layer0_outputs(8719)) and (layer0_outputs(6830)));
    outputs(11993) <= layer0_outputs(916);
    outputs(11994) <= not(layer0_outputs(800));
    outputs(11995) <= (layer0_outputs(2979)) and (layer0_outputs(636));
    outputs(11996) <= not(layer0_outputs(939));
    outputs(11997) <= layer0_outputs(4576);
    outputs(11998) <= (layer0_outputs(2694)) and (layer0_outputs(5893));
    outputs(11999) <= not(layer0_outputs(2907));
    outputs(12000) <= (layer0_outputs(1993)) xor (layer0_outputs(9502));
    outputs(12001) <= not((layer0_outputs(4098)) xor (layer0_outputs(11138)));
    outputs(12002) <= not((layer0_outputs(11643)) xor (layer0_outputs(9187)));
    outputs(12003) <= (layer0_outputs(682)) xor (layer0_outputs(4238));
    outputs(12004) <= '0';
    outputs(12005) <= (layer0_outputs(1805)) xor (layer0_outputs(11404));
    outputs(12006) <= (layer0_outputs(2141)) xor (layer0_outputs(11830));
    outputs(12007) <= '0';
    outputs(12008) <= not(layer0_outputs(1530));
    outputs(12009) <= (layer0_outputs(8090)) and (layer0_outputs(4389));
    outputs(12010) <= layer0_outputs(8865);
    outputs(12011) <= (layer0_outputs(6872)) xor (layer0_outputs(11853));
    outputs(12012) <= layer0_outputs(8533);
    outputs(12013) <= layer0_outputs(10508);
    outputs(12014) <= layer0_outputs(8661);
    outputs(12015) <= not((layer0_outputs(6625)) xor (layer0_outputs(2930)));
    outputs(12016) <= not((layer0_outputs(9989)) xor (layer0_outputs(355)));
    outputs(12017) <= (layer0_outputs(6931)) and (layer0_outputs(8856));
    outputs(12018) <= (layer0_outputs(2294)) and not (layer0_outputs(6668));
    outputs(12019) <= not((layer0_outputs(10142)) xor (layer0_outputs(10837)));
    outputs(12020) <= not(layer0_outputs(7366));
    outputs(12021) <= not((layer0_outputs(2735)) xor (layer0_outputs(11995)));
    outputs(12022) <= not(layer0_outputs(2033));
    outputs(12023) <= not(layer0_outputs(7593)) or (layer0_outputs(9149));
    outputs(12024) <= layer0_outputs(5208);
    outputs(12025) <= layer0_outputs(10999);
    outputs(12026) <= layer0_outputs(9387);
    outputs(12027) <= not(layer0_outputs(6009));
    outputs(12028) <= not(layer0_outputs(8642));
    outputs(12029) <= (layer0_outputs(718)) or (layer0_outputs(11093));
    outputs(12030) <= (layer0_outputs(10927)) xor (layer0_outputs(4632));
    outputs(12031) <= layer0_outputs(9071);
    outputs(12032) <= '0';
    outputs(12033) <= not((layer0_outputs(11898)) xor (layer0_outputs(1015)));
    outputs(12034) <= not(layer0_outputs(8482));
    outputs(12035) <= (layer0_outputs(12601)) and (layer0_outputs(8297));
    outputs(12036) <= not(layer0_outputs(11949));
    outputs(12037) <= not(layer0_outputs(8388));
    outputs(12038) <= not((layer0_outputs(33)) xor (layer0_outputs(6260)));
    outputs(12039) <= not(layer0_outputs(7228));
    outputs(12040) <= not(layer0_outputs(1391));
    outputs(12041) <= layer0_outputs(48);
    outputs(12042) <= not(layer0_outputs(6263));
    outputs(12043) <= layer0_outputs(5536);
    outputs(12044) <= layer0_outputs(2977);
    outputs(12045) <= not(layer0_outputs(10267));
    outputs(12046) <= (layer0_outputs(8498)) and not (layer0_outputs(8506));
    outputs(12047) <= not((layer0_outputs(12342)) xor (layer0_outputs(11963)));
    outputs(12048) <= not(layer0_outputs(7288)) or (layer0_outputs(10261));
    outputs(12049) <= not(layer0_outputs(117));
    outputs(12050) <= not((layer0_outputs(3299)) xor (layer0_outputs(987)));
    outputs(12051) <= not(layer0_outputs(12380));
    outputs(12052) <= not((layer0_outputs(1074)) xor (layer0_outputs(8117)));
    outputs(12053) <= layer0_outputs(6809);
    outputs(12054) <= (layer0_outputs(9776)) xor (layer0_outputs(8752));
    outputs(12055) <= not((layer0_outputs(9345)) xor (layer0_outputs(2434)));
    outputs(12056) <= (layer0_outputs(4598)) and not (layer0_outputs(3103));
    outputs(12057) <= layer0_outputs(12027);
    outputs(12058) <= layer0_outputs(7155);
    outputs(12059) <= not((layer0_outputs(12615)) xor (layer0_outputs(2776)));
    outputs(12060) <= (layer0_outputs(7302)) and not (layer0_outputs(2417));
    outputs(12061) <= not(layer0_outputs(1986)) or (layer0_outputs(7118));
    outputs(12062) <= layer0_outputs(3440);
    outputs(12063) <= layer0_outputs(11460);
    outputs(12064) <= (layer0_outputs(10806)) and not (layer0_outputs(4990));
    outputs(12065) <= not(layer0_outputs(2067));
    outputs(12066) <= layer0_outputs(10826);
    outputs(12067) <= not((layer0_outputs(12099)) and (layer0_outputs(786)));
    outputs(12068) <= not((layer0_outputs(1096)) xor (layer0_outputs(4020)));
    outputs(12069) <= not(layer0_outputs(7809)) or (layer0_outputs(2113));
    outputs(12070) <= layer0_outputs(9308);
    outputs(12071) <= not((layer0_outputs(6145)) xor (layer0_outputs(10467)));
    outputs(12072) <= layer0_outputs(2677);
    outputs(12073) <= layer0_outputs(12157);
    outputs(12074) <= (layer0_outputs(1200)) xor (layer0_outputs(3845));
    outputs(12075) <= (layer0_outputs(10188)) or (layer0_outputs(7719));
    outputs(12076) <= not(layer0_outputs(2318));
    outputs(12077) <= not(layer0_outputs(9897));
    outputs(12078) <= not(layer0_outputs(5562));
    outputs(12079) <= not(layer0_outputs(7482));
    outputs(12080) <= not(layer0_outputs(2288));
    outputs(12081) <= not(layer0_outputs(2746));
    outputs(12082) <= not((layer0_outputs(6780)) xor (layer0_outputs(6479)));
    outputs(12083) <= (layer0_outputs(11814)) or (layer0_outputs(12235));
    outputs(12084) <= (layer0_outputs(10873)) and not (layer0_outputs(1070));
    outputs(12085) <= layer0_outputs(11691);
    outputs(12086) <= (layer0_outputs(11358)) and (layer0_outputs(2960));
    outputs(12087) <= not(layer0_outputs(510));
    outputs(12088) <= not((layer0_outputs(11572)) xor (layer0_outputs(9812)));
    outputs(12089) <= not(layer0_outputs(5653)) or (layer0_outputs(732));
    outputs(12090) <= (layer0_outputs(8034)) xor (layer0_outputs(9251));
    outputs(12091) <= not((layer0_outputs(1668)) xor (layer0_outputs(11732)));
    outputs(12092) <= (layer0_outputs(4674)) and not (layer0_outputs(10144));
    outputs(12093) <= (layer0_outputs(5688)) xor (layer0_outputs(7584));
    outputs(12094) <= (layer0_outputs(2104)) and not (layer0_outputs(5164));
    outputs(12095) <= not((layer0_outputs(5354)) or (layer0_outputs(1068)));
    outputs(12096) <= not((layer0_outputs(3940)) xor (layer0_outputs(9674)));
    outputs(12097) <= '0';
    outputs(12098) <= layer0_outputs(11118);
    outputs(12099) <= layer0_outputs(2265);
    outputs(12100) <= (layer0_outputs(452)) and not (layer0_outputs(6881));
    outputs(12101) <= (layer0_outputs(9996)) and not (layer0_outputs(12250));
    outputs(12102) <= (layer0_outputs(5604)) xor (layer0_outputs(10478));
    outputs(12103) <= layer0_outputs(12611);
    outputs(12104) <= layer0_outputs(11095);
    outputs(12105) <= layer0_outputs(9846);
    outputs(12106) <= (layer0_outputs(10239)) or (layer0_outputs(11124));
    outputs(12107) <= not((layer0_outputs(9632)) xor (layer0_outputs(10332)));
    outputs(12108) <= (layer0_outputs(8794)) xor (layer0_outputs(10618));
    outputs(12109) <= not((layer0_outputs(6772)) or (layer0_outputs(5042)));
    outputs(12110) <= not((layer0_outputs(1511)) xor (layer0_outputs(4770)));
    outputs(12111) <= not(layer0_outputs(10569));
    outputs(12112) <= (layer0_outputs(919)) xor (layer0_outputs(1147));
    outputs(12113) <= (layer0_outputs(410)) xor (layer0_outputs(10265));
    outputs(12114) <= not((layer0_outputs(11615)) xor (layer0_outputs(9367)));
    outputs(12115) <= layer0_outputs(214);
    outputs(12116) <= layer0_outputs(5425);
    outputs(12117) <= (layer0_outputs(3687)) xor (layer0_outputs(7819));
    outputs(12118) <= not(layer0_outputs(1101));
    outputs(12119) <= (layer0_outputs(9633)) xor (layer0_outputs(6883));
    outputs(12120) <= not(layer0_outputs(12086)) or (layer0_outputs(8525));
    outputs(12121) <= not((layer0_outputs(12523)) xor (layer0_outputs(4132)));
    outputs(12122) <= not((layer0_outputs(11629)) or (layer0_outputs(3801)));
    outputs(12123) <= not(layer0_outputs(11748)) or (layer0_outputs(3919));
    outputs(12124) <= not((layer0_outputs(7743)) xor (layer0_outputs(3784)));
    outputs(12125) <= not(layer0_outputs(5130));
    outputs(12126) <= not(layer0_outputs(6576));
    outputs(12127) <= not((layer0_outputs(12353)) xor (layer0_outputs(4464)));
    outputs(12128) <= not(layer0_outputs(5404));
    outputs(12129) <= not(layer0_outputs(7162));
    outputs(12130) <= not((layer0_outputs(11338)) or (layer0_outputs(6130)));
    outputs(12131) <= (layer0_outputs(1219)) xor (layer0_outputs(4365));
    outputs(12132) <= (layer0_outputs(10079)) xor (layer0_outputs(4562));
    outputs(12133) <= not((layer0_outputs(3778)) or (layer0_outputs(11829)));
    outputs(12134) <= not(layer0_outputs(12028)) or (layer0_outputs(4771));
    outputs(12135) <= (layer0_outputs(3670)) xor (layer0_outputs(9429));
    outputs(12136) <= not(layer0_outputs(2205)) or (layer0_outputs(8301));
    outputs(12137) <= layer0_outputs(9545);
    outputs(12138) <= layer0_outputs(10930);
    outputs(12139) <= not(layer0_outputs(7675));
    outputs(12140) <= not(layer0_outputs(1026));
    outputs(12141) <= not((layer0_outputs(10432)) xor (layer0_outputs(9209)));
    outputs(12142) <= layer0_outputs(9299);
    outputs(12143) <= not((layer0_outputs(1014)) xor (layer0_outputs(852)));
    outputs(12144) <= (layer0_outputs(11318)) xor (layer0_outputs(1126));
    outputs(12145) <= (layer0_outputs(2645)) and not (layer0_outputs(11086));
    outputs(12146) <= not(layer0_outputs(6382));
    outputs(12147) <= not(layer0_outputs(10389));
    outputs(12148) <= (layer0_outputs(4597)) and (layer0_outputs(143));
    outputs(12149) <= not(layer0_outputs(1449));
    outputs(12150) <= (layer0_outputs(206)) xor (layer0_outputs(9950));
    outputs(12151) <= not((layer0_outputs(7851)) xor (layer0_outputs(3371)));
    outputs(12152) <= (layer0_outputs(4810)) xor (layer0_outputs(572));
    outputs(12153) <= not(layer0_outputs(8938));
    outputs(12154) <= not((layer0_outputs(127)) xor (layer0_outputs(7610)));
    outputs(12155) <= (layer0_outputs(11591)) xor (layer0_outputs(4237));
    outputs(12156) <= layer0_outputs(10159);
    outputs(12157) <= not((layer0_outputs(4933)) xor (layer0_outputs(11257)));
    outputs(12158) <= not((layer0_outputs(9490)) xor (layer0_outputs(8311)));
    outputs(12159) <= (layer0_outputs(4090)) xor (layer0_outputs(4656));
    outputs(12160) <= (layer0_outputs(2701)) and (layer0_outputs(8219));
    outputs(12161) <= not((layer0_outputs(9320)) xor (layer0_outputs(9699)));
    outputs(12162) <= layer0_outputs(12483);
    outputs(12163) <= (layer0_outputs(4534)) and not (layer0_outputs(9497));
    outputs(12164) <= layer0_outputs(10075);
    outputs(12165) <= (layer0_outputs(9889)) xor (layer0_outputs(1267));
    outputs(12166) <= (layer0_outputs(9655)) and (layer0_outputs(11164));
    outputs(12167) <= layer0_outputs(545);
    outputs(12168) <= (layer0_outputs(10765)) or (layer0_outputs(5010));
    outputs(12169) <= not((layer0_outputs(12470)) xor (layer0_outputs(3445)));
    outputs(12170) <= not(layer0_outputs(665));
    outputs(12171) <= not((layer0_outputs(12130)) xor (layer0_outputs(4201)));
    outputs(12172) <= not((layer0_outputs(9253)) xor (layer0_outputs(11113)));
    outputs(12173) <= not((layer0_outputs(10323)) xor (layer0_outputs(4936)));
    outputs(12174) <= (layer0_outputs(4929)) xor (layer0_outputs(6360));
    outputs(12175) <= not(layer0_outputs(11051));
    outputs(12176) <= not((layer0_outputs(1291)) xor (layer0_outputs(8267)));
    outputs(12177) <= layer0_outputs(2608);
    outputs(12178) <= (layer0_outputs(10466)) xor (layer0_outputs(5112));
    outputs(12179) <= not(layer0_outputs(3344));
    outputs(12180) <= not((layer0_outputs(3483)) xor (layer0_outputs(8088)));
    outputs(12181) <= (layer0_outputs(4148)) and (layer0_outputs(3450));
    outputs(12182) <= layer0_outputs(7391);
    outputs(12183) <= layer0_outputs(8651);
    outputs(12184) <= not((layer0_outputs(1243)) xor (layer0_outputs(8531)));
    outputs(12185) <= not((layer0_outputs(2566)) or (layer0_outputs(5904)));
    outputs(12186) <= layer0_outputs(1901);
    outputs(12187) <= not(layer0_outputs(7606));
    outputs(12188) <= layer0_outputs(10338);
    outputs(12189) <= not(layer0_outputs(10509));
    outputs(12190) <= (layer0_outputs(10339)) xor (layer0_outputs(541));
    outputs(12191) <= layer0_outputs(5219);
    outputs(12192) <= not(layer0_outputs(6264));
    outputs(12193) <= (layer0_outputs(4363)) and not (layer0_outputs(6435));
    outputs(12194) <= layer0_outputs(10815);
    outputs(12195) <= (layer0_outputs(9283)) and not (layer0_outputs(11350));
    outputs(12196) <= '1';
    outputs(12197) <= (layer0_outputs(5079)) xor (layer0_outputs(12244));
    outputs(12198) <= layer0_outputs(5403);
    outputs(12199) <= not(layer0_outputs(2261));
    outputs(12200) <= (layer0_outputs(6923)) xor (layer0_outputs(9457));
    outputs(12201) <= not((layer0_outputs(11482)) or (layer0_outputs(7679)));
    outputs(12202) <= not((layer0_outputs(7026)) xor (layer0_outputs(4968)));
    outputs(12203) <= not((layer0_outputs(6466)) xor (layer0_outputs(5455)));
    outputs(12204) <= (layer0_outputs(9232)) and not (layer0_outputs(12427));
    outputs(12205) <= (layer0_outputs(7313)) and not (layer0_outputs(313));
    outputs(12206) <= (layer0_outputs(4930)) xor (layer0_outputs(9307));
    outputs(12207) <= not(layer0_outputs(10112));
    outputs(12208) <= (layer0_outputs(620)) and (layer0_outputs(8470));
    outputs(12209) <= not((layer0_outputs(10177)) xor (layer0_outputs(12534)));
    outputs(12210) <= layer0_outputs(3785);
    outputs(12211) <= not((layer0_outputs(5210)) xor (layer0_outputs(5249)));
    outputs(12212) <= not((layer0_outputs(8571)) xor (layer0_outputs(7853)));
    outputs(12213) <= not(layer0_outputs(669));
    outputs(12214) <= not(layer0_outputs(423)) or (layer0_outputs(2313));
    outputs(12215) <= not(layer0_outputs(11243));
    outputs(12216) <= layer0_outputs(9813);
    outputs(12217) <= (layer0_outputs(4473)) xor (layer0_outputs(3945));
    outputs(12218) <= not((layer0_outputs(9659)) xor (layer0_outputs(2262)));
    outputs(12219) <= not(layer0_outputs(2866));
    outputs(12220) <= not((layer0_outputs(7506)) or (layer0_outputs(3719)));
    outputs(12221) <= not((layer0_outputs(127)) xor (layer0_outputs(10862)));
    outputs(12222) <= not((layer0_outputs(9717)) and (layer0_outputs(12643)));
    outputs(12223) <= layer0_outputs(12774);
    outputs(12224) <= not(layer0_outputs(5172));
    outputs(12225) <= not((layer0_outputs(3077)) and (layer0_outputs(7321)));
    outputs(12226) <= layer0_outputs(10935);
    outputs(12227) <= not((layer0_outputs(2487)) xor (layer0_outputs(3256)));
    outputs(12228) <= not(layer0_outputs(5576));
    outputs(12229) <= (layer0_outputs(6926)) and not (layer0_outputs(6688));
    outputs(12230) <= not((layer0_outputs(10897)) xor (layer0_outputs(5883)));
    outputs(12231) <= not(layer0_outputs(9761));
    outputs(12232) <= (layer0_outputs(12010)) and (layer0_outputs(3531));
    outputs(12233) <= not(layer0_outputs(4207));
    outputs(12234) <= not((layer0_outputs(6851)) and (layer0_outputs(6081)));
    outputs(12235) <= not(layer0_outputs(5705));
    outputs(12236) <= layer0_outputs(6453);
    outputs(12237) <= layer0_outputs(588);
    outputs(12238) <= layer0_outputs(1013);
    outputs(12239) <= (layer0_outputs(4659)) xor (layer0_outputs(2771));
    outputs(12240) <= layer0_outputs(7647);
    outputs(12241) <= layer0_outputs(6315);
    outputs(12242) <= not(layer0_outputs(7372)) or (layer0_outputs(10155));
    outputs(12243) <= layer0_outputs(7290);
    outputs(12244) <= layer0_outputs(3714);
    outputs(12245) <= not(layer0_outputs(9525));
    outputs(12246) <= (layer0_outputs(10117)) xor (layer0_outputs(10376));
    outputs(12247) <= not(layer0_outputs(1302)) or (layer0_outputs(11148));
    outputs(12248) <= (layer0_outputs(4617)) and not (layer0_outputs(6842));
    outputs(12249) <= not((layer0_outputs(11298)) xor (layer0_outputs(6891)));
    outputs(12250) <= layer0_outputs(1588);
    outputs(12251) <= (layer0_outputs(8587)) xor (layer0_outputs(11791));
    outputs(12252) <= layer0_outputs(2509);
    outputs(12253) <= not((layer0_outputs(3675)) xor (layer0_outputs(4669)));
    outputs(12254) <= (layer0_outputs(10137)) xor (layer0_outputs(7465));
    outputs(12255) <= (layer0_outputs(7282)) and not (layer0_outputs(8599));
    outputs(12256) <= not(layer0_outputs(61));
    outputs(12257) <= not((layer0_outputs(9396)) and (layer0_outputs(7524)));
    outputs(12258) <= not((layer0_outputs(746)) or (layer0_outputs(3893)));
    outputs(12259) <= not((layer0_outputs(7716)) or (layer0_outputs(6827)));
    outputs(12260) <= (layer0_outputs(12185)) xor (layer0_outputs(11310));
    outputs(12261) <= (layer0_outputs(318)) and (layer0_outputs(902));
    outputs(12262) <= not(layer0_outputs(7016)) or (layer0_outputs(12214));
    outputs(12263) <= not((layer0_outputs(3280)) xor (layer0_outputs(247)));
    outputs(12264) <= not((layer0_outputs(2488)) xor (layer0_outputs(6015)));
    outputs(12265) <= not((layer0_outputs(740)) xor (layer0_outputs(4158)));
    outputs(12266) <= layer0_outputs(12126);
    outputs(12267) <= (layer0_outputs(5573)) and (layer0_outputs(3166));
    outputs(12268) <= layer0_outputs(433);
    outputs(12269) <= (layer0_outputs(3598)) and (layer0_outputs(3721));
    outputs(12270) <= not((layer0_outputs(9805)) xor (layer0_outputs(11327)));
    outputs(12271) <= (layer0_outputs(936)) xor (layer0_outputs(1791));
    outputs(12272) <= layer0_outputs(10572);
    outputs(12273) <= layer0_outputs(4003);
    outputs(12274) <= not(layer0_outputs(10486));
    outputs(12275) <= layer0_outputs(3459);
    outputs(12276) <= (layer0_outputs(10532)) and not (layer0_outputs(1165));
    outputs(12277) <= not((layer0_outputs(2959)) xor (layer0_outputs(8165)));
    outputs(12278) <= not((layer0_outputs(4118)) xor (layer0_outputs(4514)));
    outputs(12279) <= (layer0_outputs(3875)) xor (layer0_outputs(2199));
    outputs(12280) <= not(layer0_outputs(8936));
    outputs(12281) <= not((layer0_outputs(10712)) xor (layer0_outputs(7134)));
    outputs(12282) <= (layer0_outputs(1368)) and (layer0_outputs(6471));
    outputs(12283) <= (layer0_outputs(3157)) or (layer0_outputs(2087));
    outputs(12284) <= (layer0_outputs(11041)) xor (layer0_outputs(7070));
    outputs(12285) <= not(layer0_outputs(11024));
    outputs(12286) <= (layer0_outputs(2342)) xor (layer0_outputs(849));
    outputs(12287) <= not((layer0_outputs(9334)) xor (layer0_outputs(287)));
    outputs(12288) <= not((layer0_outputs(2928)) xor (layer0_outputs(8588)));
    outputs(12289) <= not(layer0_outputs(512));
    outputs(12290) <= not(layer0_outputs(12308));
    outputs(12291) <= not((layer0_outputs(8414)) xor (layer0_outputs(2847)));
    outputs(12292) <= (layer0_outputs(6132)) and (layer0_outputs(8705));
    outputs(12293) <= not((layer0_outputs(12262)) xor (layer0_outputs(2289)));
    outputs(12294) <= not(layer0_outputs(11324));
    outputs(12295) <= layer0_outputs(3028);
    outputs(12296) <= not(layer0_outputs(370)) or (layer0_outputs(6154));
    outputs(12297) <= not(layer0_outputs(8210));
    outputs(12298) <= not(layer0_outputs(108));
    outputs(12299) <= layer0_outputs(7709);
    outputs(12300) <= not(layer0_outputs(10627));
    outputs(12301) <= (layer0_outputs(3216)) and (layer0_outputs(5849));
    outputs(12302) <= (layer0_outputs(840)) xor (layer0_outputs(9784));
    outputs(12303) <= (layer0_outputs(10898)) and not (layer0_outputs(3355));
    outputs(12304) <= (layer0_outputs(7604)) and (layer0_outputs(10786));
    outputs(12305) <= not(layer0_outputs(9046)) or (layer0_outputs(11414));
    outputs(12306) <= not((layer0_outputs(808)) xor (layer0_outputs(1216)));
    outputs(12307) <= (layer0_outputs(1604)) and not (layer0_outputs(3033));
    outputs(12308) <= layer0_outputs(11519);
    outputs(12309) <= (layer0_outputs(8552)) xor (layer0_outputs(5544));
    outputs(12310) <= layer0_outputs(1560);
    outputs(12311) <= not((layer0_outputs(3122)) xor (layer0_outputs(3552)));
    outputs(12312) <= (layer0_outputs(4888)) xor (layer0_outputs(1460));
    outputs(12313) <= (layer0_outputs(3601)) xor (layer0_outputs(2391));
    outputs(12314) <= not((layer0_outputs(3388)) or (layer0_outputs(426)));
    outputs(12315) <= not(layer0_outputs(10816));
    outputs(12316) <= (layer0_outputs(9825)) and not (layer0_outputs(5477));
    outputs(12317) <= not((layer0_outputs(5858)) xor (layer0_outputs(4320)));
    outputs(12318) <= not((layer0_outputs(2378)) xor (layer0_outputs(10502)));
    outputs(12319) <= (layer0_outputs(12712)) and not (layer0_outputs(3018));
    outputs(12320) <= layer0_outputs(4883);
    outputs(12321) <= not((layer0_outputs(11778)) xor (layer0_outputs(11632)));
    outputs(12322) <= not((layer0_outputs(11781)) or (layer0_outputs(4212)));
    outputs(12323) <= (layer0_outputs(5232)) xor (layer0_outputs(12768));
    outputs(12324) <= not((layer0_outputs(12744)) xor (layer0_outputs(2943)));
    outputs(12325) <= (layer0_outputs(7956)) or (layer0_outputs(10416));
    outputs(12326) <= (layer0_outputs(2231)) and not (layer0_outputs(3050));
    outputs(12327) <= layer0_outputs(5347);
    outputs(12328) <= not(layer0_outputs(6568));
    outputs(12329) <= (layer0_outputs(6527)) xor (layer0_outputs(2769));
    outputs(12330) <= layer0_outputs(9734);
    outputs(12331) <= (layer0_outputs(8150)) xor (layer0_outputs(5132));
    outputs(12332) <= not(layer0_outputs(7901));
    outputs(12333) <= not(layer0_outputs(6141));
    outputs(12334) <= not((layer0_outputs(6923)) or (layer0_outputs(9618)));
    outputs(12335) <= not((layer0_outputs(10496)) or (layer0_outputs(8550)));
    outputs(12336) <= (layer0_outputs(3476)) and (layer0_outputs(10806));
    outputs(12337) <= not(layer0_outputs(1445));
    outputs(12338) <= (layer0_outputs(4)) xor (layer0_outputs(11806));
    outputs(12339) <= (layer0_outputs(5647)) and (layer0_outputs(7355));
    outputs(12340) <= (layer0_outputs(2742)) xor (layer0_outputs(12215));
    outputs(12341) <= (layer0_outputs(8010)) and not (layer0_outputs(5731));
    outputs(12342) <= layer0_outputs(9265);
    outputs(12343) <= not((layer0_outputs(4070)) xor (layer0_outputs(11937)));
    outputs(12344) <= not(layer0_outputs(2508));
    outputs(12345) <= layer0_outputs(4765);
    outputs(12346) <= not(layer0_outputs(8283));
    outputs(12347) <= not((layer0_outputs(12792)) xor (layer0_outputs(428)));
    outputs(12348) <= (layer0_outputs(8039)) xor (layer0_outputs(5242));
    outputs(12349) <= not((layer0_outputs(5855)) or (layer0_outputs(11388)));
    outputs(12350) <= (layer0_outputs(8992)) xor (layer0_outputs(302));
    outputs(12351) <= (layer0_outputs(3483)) xor (layer0_outputs(3747));
    outputs(12352) <= (layer0_outputs(10271)) and not (layer0_outputs(11920));
    outputs(12353) <= layer0_outputs(6710);
    outputs(12354) <= (layer0_outputs(158)) and not (layer0_outputs(2691));
    outputs(12355) <= (layer0_outputs(1000)) xor (layer0_outputs(2128));
    outputs(12356) <= layer0_outputs(2032);
    outputs(12357) <= not((layer0_outputs(6281)) xor (layer0_outputs(6231)));
    outputs(12358) <= not((layer0_outputs(896)) xor (layer0_outputs(3668)));
    outputs(12359) <= not((layer0_outputs(6751)) or (layer0_outputs(700)));
    outputs(12360) <= not((layer0_outputs(12521)) xor (layer0_outputs(5979)));
    outputs(12361) <= not((layer0_outputs(5350)) or (layer0_outputs(2489)));
    outputs(12362) <= layer0_outputs(2805);
    outputs(12363) <= not(layer0_outputs(9104));
    outputs(12364) <= not(layer0_outputs(10201));
    outputs(12365) <= not(layer0_outputs(1735)) or (layer0_outputs(10854));
    outputs(12366) <= (layer0_outputs(721)) and (layer0_outputs(7501));
    outputs(12367) <= not(layer0_outputs(2528));
    outputs(12368) <= (layer0_outputs(9953)) xor (layer0_outputs(12640));
    outputs(12369) <= (layer0_outputs(3121)) xor (layer0_outputs(9136));
    outputs(12370) <= not(layer0_outputs(4106));
    outputs(12371) <= not(layer0_outputs(9074));
    outputs(12372) <= (layer0_outputs(10986)) and (layer0_outputs(9619));
    outputs(12373) <= layer0_outputs(9642);
    outputs(12374) <= (layer0_outputs(11118)) or (layer0_outputs(5440));
    outputs(12375) <= layer0_outputs(9988);
    outputs(12376) <= not(layer0_outputs(221));
    outputs(12377) <= layer0_outputs(509);
    outputs(12378) <= not((layer0_outputs(5805)) xor (layer0_outputs(11270)));
    outputs(12379) <= (layer0_outputs(3603)) xor (layer0_outputs(10238));
    outputs(12380) <= not(layer0_outputs(10235));
    outputs(12381) <= not(layer0_outputs(9697)) or (layer0_outputs(11918));
    outputs(12382) <= (layer0_outputs(3865)) and (layer0_outputs(12602));
    outputs(12383) <= (layer0_outputs(10537)) and (layer0_outputs(1402));
    outputs(12384) <= not((layer0_outputs(5854)) xor (layer0_outputs(4695)));
    outputs(12385) <= not(layer0_outputs(9369)) or (layer0_outputs(8411));
    outputs(12386) <= not((layer0_outputs(2552)) xor (layer0_outputs(4679)));
    outputs(12387) <= (layer0_outputs(3)) and not (layer0_outputs(8096));
    outputs(12388) <= (layer0_outputs(5740)) and not (layer0_outputs(1848));
    outputs(12389) <= not(layer0_outputs(5707));
    outputs(12390) <= not(layer0_outputs(4592));
    outputs(12391) <= (layer0_outputs(688)) xor (layer0_outputs(11211));
    outputs(12392) <= not((layer0_outputs(12147)) xor (layer0_outputs(12460)));
    outputs(12393) <= (layer0_outputs(12332)) xor (layer0_outputs(1596));
    outputs(12394) <= layer0_outputs(6184);
    outputs(12395) <= not((layer0_outputs(9311)) xor (layer0_outputs(9915)));
    outputs(12396) <= (layer0_outputs(3821)) xor (layer0_outputs(3271));
    outputs(12397) <= not(layer0_outputs(602)) or (layer0_outputs(1044));
    outputs(12398) <= not((layer0_outputs(11986)) and (layer0_outputs(8820)));
    outputs(12399) <= (layer0_outputs(508)) xor (layer0_outputs(4835));
    outputs(12400) <= layer0_outputs(557);
    outputs(12401) <= (layer0_outputs(7285)) and not (layer0_outputs(10793));
    outputs(12402) <= not(layer0_outputs(8590));
    outputs(12403) <= not((layer0_outputs(5258)) xor (layer0_outputs(6093)));
    outputs(12404) <= layer0_outputs(1790);
    outputs(12405) <= (layer0_outputs(10226)) and not (layer0_outputs(9432));
    outputs(12406) <= not(layer0_outputs(12306));
    outputs(12407) <= (layer0_outputs(5092)) xor (layer0_outputs(9788));
    outputs(12408) <= not((layer0_outputs(9979)) or (layer0_outputs(12072)));
    outputs(12409) <= not(layer0_outputs(2541));
    outputs(12410) <= (layer0_outputs(5233)) and not (layer0_outputs(2416));
    outputs(12411) <= not(layer0_outputs(10609));
    outputs(12412) <= not((layer0_outputs(629)) xor (layer0_outputs(11112)));
    outputs(12413) <= (layer0_outputs(12746)) and not (layer0_outputs(6533));
    outputs(12414) <= layer0_outputs(4165);
    outputs(12415) <= '0';
    outputs(12416) <= layer0_outputs(10891);
    outputs(12417) <= not((layer0_outputs(1545)) xor (layer0_outputs(9942)));
    outputs(12418) <= not(layer0_outputs(9516));
    outputs(12419) <= layer0_outputs(2895);
    outputs(12420) <= not((layer0_outputs(12121)) xor (layer0_outputs(12019)));
    outputs(12421) <= (layer0_outputs(12743)) and not (layer0_outputs(9886));
    outputs(12422) <= not((layer0_outputs(4025)) xor (layer0_outputs(4134)));
    outputs(12423) <= (layer0_outputs(10275)) xor (layer0_outputs(1710));
    outputs(12424) <= (layer0_outputs(3735)) and not (layer0_outputs(390));
    outputs(12425) <= not(layer0_outputs(2636));
    outputs(12426) <= not(layer0_outputs(3649));
    outputs(12427) <= not((layer0_outputs(8370)) xor (layer0_outputs(3631)));
    outputs(12428) <= not(layer0_outputs(8359));
    outputs(12429) <= layer0_outputs(10715);
    outputs(12430) <= layer0_outputs(6755);
    outputs(12431) <= not((layer0_outputs(878)) xor (layer0_outputs(12376)));
    outputs(12432) <= (layer0_outputs(585)) and (layer0_outputs(10541));
    outputs(12433) <= layer0_outputs(1292);
    outputs(12434) <= not((layer0_outputs(7863)) xor (layer0_outputs(3248)));
    outputs(12435) <= not((layer0_outputs(169)) or (layer0_outputs(7841)));
    outputs(12436) <= not(layer0_outputs(8954));
    outputs(12437) <= layer0_outputs(28);
    outputs(12438) <= not((layer0_outputs(11046)) or (layer0_outputs(1104)));
    outputs(12439) <= not((layer0_outputs(9818)) xor (layer0_outputs(11195)));
    outputs(12440) <= not((layer0_outputs(8939)) or (layer0_outputs(9082)));
    outputs(12441) <= not(layer0_outputs(12371));
    outputs(12442) <= not(layer0_outputs(2798)) or (layer0_outputs(1282));
    outputs(12443) <= (layer0_outputs(7937)) xor (layer0_outputs(1461));
    outputs(12444) <= layer0_outputs(3447);
    outputs(12445) <= not(layer0_outputs(535));
    outputs(12446) <= not((layer0_outputs(8106)) or (layer0_outputs(11110)));
    outputs(12447) <= layer0_outputs(2308);
    outputs(12448) <= (layer0_outputs(10567)) xor (layer0_outputs(1139));
    outputs(12449) <= layer0_outputs(10009);
    outputs(12450) <= not(layer0_outputs(12238));
    outputs(12451) <= layer0_outputs(5671);
    outputs(12452) <= not((layer0_outputs(9913)) xor (layer0_outputs(11912)));
    outputs(12453) <= (layer0_outputs(3963)) and not (layer0_outputs(7711));
    outputs(12454) <= not((layer0_outputs(8385)) xor (layer0_outputs(3629)));
    outputs(12455) <= not(layer0_outputs(8650));
    outputs(12456) <= (layer0_outputs(3442)) xor (layer0_outputs(11331));
    outputs(12457) <= not((layer0_outputs(3609)) xor (layer0_outputs(10590)));
    outputs(12458) <= not(layer0_outputs(4502));
    outputs(12459) <= layer0_outputs(5667);
    outputs(12460) <= not((layer0_outputs(1457)) and (layer0_outputs(9768)));
    outputs(12461) <= (layer0_outputs(2936)) and not (layer0_outputs(3921));
    outputs(12462) <= layer0_outputs(4910);
    outputs(12463) <= (layer0_outputs(3146)) xor (layer0_outputs(5387));
    outputs(12464) <= not((layer0_outputs(9881)) xor (layer0_outputs(8646)));
    outputs(12465) <= not((layer0_outputs(7237)) xor (layer0_outputs(3925)));
    outputs(12466) <= layer0_outputs(10932);
    outputs(12467) <= not((layer0_outputs(5618)) xor (layer0_outputs(8645)));
    outputs(12468) <= not(layer0_outputs(10424));
    outputs(12469) <= not(layer0_outputs(7933));
    outputs(12470) <= not((layer0_outputs(3745)) xor (layer0_outputs(685)));
    outputs(12471) <= not(layer0_outputs(4469));
    outputs(12472) <= (layer0_outputs(12524)) xor (layer0_outputs(2071));
    outputs(12473) <= not(layer0_outputs(3957));
    outputs(12474) <= not((layer0_outputs(6064)) and (layer0_outputs(8388)));
    outputs(12475) <= not(layer0_outputs(7030));
    outputs(12476) <= not((layer0_outputs(5748)) and (layer0_outputs(89)));
    outputs(12477) <= layer0_outputs(6929);
    outputs(12478) <= (layer0_outputs(4934)) xor (layer0_outputs(2834));
    outputs(12479) <= not(layer0_outputs(5295));
    outputs(12480) <= (layer0_outputs(7585)) xor (layer0_outputs(5170));
    outputs(12481) <= not(layer0_outputs(10827));
    outputs(12482) <= not((layer0_outputs(549)) and (layer0_outputs(9455)));
    outputs(12483) <= not((layer0_outputs(3162)) xor (layer0_outputs(2943)));
    outputs(12484) <= (layer0_outputs(7798)) xor (layer0_outputs(8715));
    outputs(12485) <= not((layer0_outputs(11910)) xor (layer0_outputs(10122)));
    outputs(12486) <= not(layer0_outputs(12173));
    outputs(12487) <= layer0_outputs(7160);
    outputs(12488) <= not((layer0_outputs(2954)) or (layer0_outputs(11284)));
    outputs(12489) <= (layer0_outputs(5905)) xor (layer0_outputs(10607));
    outputs(12490) <= (layer0_outputs(8864)) and (layer0_outputs(6883));
    outputs(12491) <= (layer0_outputs(9378)) and not (layer0_outputs(4351));
    outputs(12492) <= (layer0_outputs(1158)) xor (layer0_outputs(4978));
    outputs(12493) <= not((layer0_outputs(12394)) and (layer0_outputs(10847)));
    outputs(12494) <= not(layer0_outputs(7148));
    outputs(12495) <= '0';
    outputs(12496) <= not((layer0_outputs(10381)) xor (layer0_outputs(6282)));
    outputs(12497) <= (layer0_outputs(6938)) or (layer0_outputs(737));
    outputs(12498) <= layer0_outputs(12492);
    outputs(12499) <= not((layer0_outputs(12201)) or (layer0_outputs(6854)));
    outputs(12500) <= not((layer0_outputs(2372)) xor (layer0_outputs(2398)));
    outputs(12501) <= not((layer0_outputs(4622)) xor (layer0_outputs(1767)));
    outputs(12502) <= not(layer0_outputs(6824));
    outputs(12503) <= not((layer0_outputs(12482)) or (layer0_outputs(9781)));
    outputs(12504) <= layer0_outputs(6593);
    outputs(12505) <= not(layer0_outputs(3350));
    outputs(12506) <= not(layer0_outputs(1142));
    outputs(12507) <= (layer0_outputs(9636)) and not (layer0_outputs(10272));
    outputs(12508) <= not((layer0_outputs(7330)) xor (layer0_outputs(10224)));
    outputs(12509) <= not(layer0_outputs(10211)) or (layer0_outputs(12721));
    outputs(12510) <= (layer0_outputs(9557)) xor (layer0_outputs(6046));
    outputs(12511) <= not(layer0_outputs(4812)) or (layer0_outputs(7723));
    outputs(12512) <= layer0_outputs(8276);
    outputs(12513) <= not(layer0_outputs(7689));
    outputs(12514) <= not(layer0_outputs(1227));
    outputs(12515) <= not((layer0_outputs(5402)) xor (layer0_outputs(3199)));
    outputs(12516) <= layer0_outputs(8403);
    outputs(12517) <= not(layer0_outputs(6508));
    outputs(12518) <= (layer0_outputs(1649)) and (layer0_outputs(2996));
    outputs(12519) <= (layer0_outputs(3634)) and not (layer0_outputs(306));
    outputs(12520) <= (layer0_outputs(3323)) xor (layer0_outputs(6842));
    outputs(12521) <= (layer0_outputs(5982)) xor (layer0_outputs(10680));
    outputs(12522) <= not((layer0_outputs(2365)) xor (layer0_outputs(8655)));
    outputs(12523) <= (layer0_outputs(12251)) xor (layer0_outputs(11479));
    outputs(12524) <= not((layer0_outputs(1316)) xor (layer0_outputs(9203)));
    outputs(12525) <= not((layer0_outputs(474)) xor (layer0_outputs(685)));
    outputs(12526) <= layer0_outputs(4719);
    outputs(12527) <= (layer0_outputs(12049)) and (layer0_outputs(2220));
    outputs(12528) <= not(layer0_outputs(1994));
    outputs(12529) <= not((layer0_outputs(9013)) xor (layer0_outputs(1681)));
    outputs(12530) <= (layer0_outputs(3700)) and (layer0_outputs(10058));
    outputs(12531) <= not(layer0_outputs(9656));
    outputs(12532) <= not((layer0_outputs(8263)) xor (layer0_outputs(10266)));
    outputs(12533) <= (layer0_outputs(11957)) and not (layer0_outputs(9618));
    outputs(12534) <= not(layer0_outputs(3163)) or (layer0_outputs(4380));
    outputs(12535) <= not((layer0_outputs(1295)) xor (layer0_outputs(5996)));
    outputs(12536) <= not(layer0_outputs(11823)) or (layer0_outputs(4890));
    outputs(12537) <= layer0_outputs(2695);
    outputs(12538) <= not((layer0_outputs(10732)) xor (layer0_outputs(4298)));
    outputs(12539) <= layer0_outputs(3547);
    outputs(12540) <= (layer0_outputs(12484)) and not (layer0_outputs(10170));
    outputs(12541) <= not(layer0_outputs(7539));
    outputs(12542) <= not(layer0_outputs(4102));
    outputs(12543) <= (layer0_outputs(854)) and not (layer0_outputs(2175));
    outputs(12544) <= not((layer0_outputs(4504)) or (layer0_outputs(8456)));
    outputs(12545) <= not((layer0_outputs(836)) xor (layer0_outputs(12783)));
    outputs(12546) <= layer0_outputs(2305);
    outputs(12547) <= not(layer0_outputs(8395));
    outputs(12548) <= (layer0_outputs(7594)) and not (layer0_outputs(11032));
    outputs(12549) <= not(layer0_outputs(7129));
    outputs(12550) <= (layer0_outputs(725)) xor (layer0_outputs(6334));
    outputs(12551) <= not((layer0_outputs(8923)) or (layer0_outputs(10023)));
    outputs(12552) <= layer0_outputs(5361);
    outputs(12553) <= not((layer0_outputs(11366)) xor (layer0_outputs(5530)));
    outputs(12554) <= not(layer0_outputs(9924));
    outputs(12555) <= not((layer0_outputs(6620)) xor (layer0_outputs(8076)));
    outputs(12556) <= (layer0_outputs(10581)) and not (layer0_outputs(6265));
    outputs(12557) <= not(layer0_outputs(9408));
    outputs(12558) <= layer0_outputs(10390);
    outputs(12559) <= (layer0_outputs(9811)) and not (layer0_outputs(4803));
    outputs(12560) <= (layer0_outputs(10880)) xor (layer0_outputs(6042));
    outputs(12561) <= (layer0_outputs(5949)) xor (layer0_outputs(11435));
    outputs(12562) <= (layer0_outputs(5029)) xor (layer0_outputs(4043));
    outputs(12563) <= not(layer0_outputs(6476));
    outputs(12564) <= (layer0_outputs(8862)) and not (layer0_outputs(7051));
    outputs(12565) <= not(layer0_outputs(5561));
    outputs(12566) <= (layer0_outputs(8391)) xor (layer0_outputs(5512));
    outputs(12567) <= layer0_outputs(6966);
    outputs(12568) <= not((layer0_outputs(9040)) or (layer0_outputs(4485)));
    outputs(12569) <= '1';
    outputs(12570) <= layer0_outputs(3947);
    outputs(12571) <= (layer0_outputs(1819)) and (layer0_outputs(3375));
    outputs(12572) <= not(layer0_outputs(3886));
    outputs(12573) <= layer0_outputs(7795);
    outputs(12574) <= not((layer0_outputs(1571)) xor (layer0_outputs(4797)));
    outputs(12575) <= layer0_outputs(8693);
    outputs(12576) <= layer0_outputs(11742);
    outputs(12577) <= (layer0_outputs(1504)) and (layer0_outputs(71));
    outputs(12578) <= not(layer0_outputs(1478));
    outputs(12579) <= (layer0_outputs(4947)) and (layer0_outputs(7641));
    outputs(12580) <= not((layer0_outputs(4267)) or (layer0_outputs(9388)));
    outputs(12581) <= (layer0_outputs(1765)) and not (layer0_outputs(5383));
    outputs(12582) <= (layer0_outputs(12524)) xor (layer0_outputs(3159));
    outputs(12583) <= (layer0_outputs(9192)) xor (layer0_outputs(12287));
    outputs(12584) <= layer0_outputs(9341);
    outputs(12585) <= layer0_outputs(8224);
    outputs(12586) <= not((layer0_outputs(993)) xor (layer0_outputs(11057)));
    outputs(12587) <= not(layer0_outputs(2388));
    outputs(12588) <= (layer0_outputs(12358)) and not (layer0_outputs(10550));
    outputs(12589) <= not((layer0_outputs(7934)) xor (layer0_outputs(2486)));
    outputs(12590) <= (layer0_outputs(10741)) and not (layer0_outputs(4963));
    outputs(12591) <= not(layer0_outputs(3928));
    outputs(12592) <= (layer0_outputs(3899)) and not (layer0_outputs(1449));
    outputs(12593) <= layer0_outputs(2923);
    outputs(12594) <= layer0_outputs(10383);
    outputs(12595) <= not(layer0_outputs(9382));
    outputs(12596) <= layer0_outputs(1608);
    outputs(12597) <= not(layer0_outputs(695));
    outputs(12598) <= layer0_outputs(6663);
    outputs(12599) <= not(layer0_outputs(1326)) or (layer0_outputs(1264));
    outputs(12600) <= not(layer0_outputs(11220));
    outputs(12601) <= (layer0_outputs(6364)) and not (layer0_outputs(1670));
    outputs(12602) <= not((layer0_outputs(4591)) xor (layer0_outputs(3704)));
    outputs(12603) <= (layer0_outputs(2056)) and not (layer0_outputs(3929));
    outputs(12604) <= not((layer0_outputs(4847)) xor (layer0_outputs(3642)));
    outputs(12605) <= layer0_outputs(11093);
    outputs(12606) <= not(layer0_outputs(4867));
    outputs(12607) <= (layer0_outputs(10085)) and not (layer0_outputs(5940));
    outputs(12608) <= not((layer0_outputs(5589)) xor (layer0_outputs(11183)));
    outputs(12609) <= not(layer0_outputs(12093));
    outputs(12610) <= (layer0_outputs(10385)) or (layer0_outputs(6485));
    outputs(12611) <= (layer0_outputs(6738)) xor (layer0_outputs(5149));
    outputs(12612) <= not((layer0_outputs(9956)) or (layer0_outputs(9794)));
    outputs(12613) <= (layer0_outputs(11744)) xor (layer0_outputs(9222));
    outputs(12614) <= (layer0_outputs(8699)) and not (layer0_outputs(1997));
    outputs(12615) <= not(layer0_outputs(7288));
    outputs(12616) <= not((layer0_outputs(265)) xor (layer0_outputs(3757)));
    outputs(12617) <= not((layer0_outputs(6994)) xor (layer0_outputs(9184)));
    outputs(12618) <= (layer0_outputs(9422)) xor (layer0_outputs(11431));
    outputs(12619) <= (layer0_outputs(10844)) and not (layer0_outputs(11836));
    outputs(12620) <= not(layer0_outputs(12067));
    outputs(12621) <= not(layer0_outputs(2585));
    outputs(12622) <= not((layer0_outputs(8041)) or (layer0_outputs(7657)));
    outputs(12623) <= not(layer0_outputs(10658));
    outputs(12624) <= (layer0_outputs(3046)) xor (layer0_outputs(942));
    outputs(12625) <= not(layer0_outputs(12443));
    outputs(12626) <= (layer0_outputs(8712)) xor (layer0_outputs(6782));
    outputs(12627) <= not(layer0_outputs(8328));
    outputs(12628) <= (layer0_outputs(4135)) xor (layer0_outputs(1301));
    outputs(12629) <= not((layer0_outputs(2256)) xor (layer0_outputs(4583)));
    outputs(12630) <= not(layer0_outputs(7317)) or (layer0_outputs(5894));
    outputs(12631) <= not(layer0_outputs(9690));
    outputs(12632) <= (layer0_outputs(2434)) and (layer0_outputs(7433));
    outputs(12633) <= not((layer0_outputs(8127)) xor (layer0_outputs(6774)));
    outputs(12634) <= not((layer0_outputs(12165)) xor (layer0_outputs(7141)));
    outputs(12635) <= not((layer0_outputs(2507)) xor (layer0_outputs(11952)));
    outputs(12636) <= (layer0_outputs(9066)) and not (layer0_outputs(1170));
    outputs(12637) <= layer0_outputs(5040);
    outputs(12638) <= layer0_outputs(12630);
    outputs(12639) <= not(layer0_outputs(693));
    outputs(12640) <= not(layer0_outputs(4625)) or (layer0_outputs(11397));
    outputs(12641) <= not((layer0_outputs(7746)) or (layer0_outputs(4287)));
    outputs(12642) <= not(layer0_outputs(3012)) or (layer0_outputs(10113));
    outputs(12643) <= (layer0_outputs(6748)) xor (layer0_outputs(6641));
    outputs(12644) <= not(layer0_outputs(11841)) or (layer0_outputs(9078));
    outputs(12645) <= layer0_outputs(104);
    outputs(12646) <= not(layer0_outputs(7479));
    outputs(12647) <= not(layer0_outputs(10255));
    outputs(12648) <= not(layer0_outputs(1167)) or (layer0_outputs(5388));
    outputs(12649) <= layer0_outputs(851);
    outputs(12650) <= not(layer0_outputs(1978));
    outputs(12651) <= not((layer0_outputs(597)) xor (layer0_outputs(6907)));
    outputs(12652) <= layer0_outputs(11586);
    outputs(12653) <= layer0_outputs(12409);
    outputs(12654) <= not(layer0_outputs(9147));
    outputs(12655) <= layer0_outputs(2926);
    outputs(12656) <= (layer0_outputs(10902)) and (layer0_outputs(6271));
    outputs(12657) <= (layer0_outputs(4304)) and not (layer0_outputs(11697));
    outputs(12658) <= (layer0_outputs(2148)) xor (layer0_outputs(496));
    outputs(12659) <= not((layer0_outputs(7674)) xor (layer0_outputs(640)));
    outputs(12660) <= not((layer0_outputs(7626)) and (layer0_outputs(423)));
    outputs(12661) <= not((layer0_outputs(10498)) and (layer0_outputs(9000)));
    outputs(12662) <= not(layer0_outputs(6437));
    outputs(12663) <= layer0_outputs(10403);
    outputs(12664) <= (layer0_outputs(5916)) and (layer0_outputs(11851));
    outputs(12665) <= not(layer0_outputs(10439));
    outputs(12666) <= layer0_outputs(2676);
    outputs(12667) <= not(layer0_outputs(6338)) or (layer0_outputs(656));
    outputs(12668) <= not(layer0_outputs(6370));
    outputs(12669) <= not((layer0_outputs(996)) xor (layer0_outputs(9835)));
    outputs(12670) <= not(layer0_outputs(10016)) or (layer0_outputs(5494));
    outputs(12671) <= layer0_outputs(4250);
    outputs(12672) <= not(layer0_outputs(931));
    outputs(12673) <= not((layer0_outputs(5963)) xor (layer0_outputs(2232)));
    outputs(12674) <= layer0_outputs(6976);
    outputs(12675) <= (layer0_outputs(6309)) xor (layer0_outputs(4211));
    outputs(12676) <= not((layer0_outputs(8626)) xor (layer0_outputs(9417)));
    outputs(12677) <= (layer0_outputs(8913)) and not (layer0_outputs(11602));
    outputs(12678) <= (layer0_outputs(4661)) xor (layer0_outputs(539));
    outputs(12679) <= layer0_outputs(11415);
    outputs(12680) <= not(layer0_outputs(11355)) or (layer0_outputs(3776));
    outputs(12681) <= layer0_outputs(12079);
    outputs(12682) <= not(layer0_outputs(4856));
    outputs(12683) <= (layer0_outputs(7697)) or (layer0_outputs(4194));
    outputs(12684) <= (layer0_outputs(403)) and not (layer0_outputs(11335));
    outputs(12685) <= not((layer0_outputs(8003)) xor (layer0_outputs(9702)));
    outputs(12686) <= not(layer0_outputs(8192));
    outputs(12687) <= layer0_outputs(7220);
    outputs(12688) <= layer0_outputs(1474);
    outputs(12689) <= layer0_outputs(1758);
    outputs(12690) <= not((layer0_outputs(1374)) xor (layer0_outputs(10605)));
    outputs(12691) <= (layer0_outputs(8536)) and not (layer0_outputs(8178));
    outputs(12692) <= not((layer0_outputs(5339)) xor (layer0_outputs(10625)));
    outputs(12693) <= (layer0_outputs(2031)) and (layer0_outputs(10760));
    outputs(12694) <= not((layer0_outputs(7281)) xor (layer0_outputs(11936)));
    outputs(12695) <= layer0_outputs(5272);
    outputs(12696) <= not((layer0_outputs(6730)) xor (layer0_outputs(12576)));
    outputs(12697) <= not(layer0_outputs(848));
    outputs(12698) <= layer0_outputs(7159);
    outputs(12699) <= layer0_outputs(10982);
    outputs(12700) <= not(layer0_outputs(4023));
    outputs(12701) <= (layer0_outputs(1403)) and (layer0_outputs(7128));
    outputs(12702) <= layer0_outputs(11768);
    outputs(12703) <= not(layer0_outputs(10685));
    outputs(12704) <= (layer0_outputs(9285)) xor (layer0_outputs(4718));
    outputs(12705) <= not((layer0_outputs(1978)) or (layer0_outputs(4398)));
    outputs(12706) <= layer0_outputs(5611);
    outputs(12707) <= not(layer0_outputs(1211));
    outputs(12708) <= layer0_outputs(11440);
    outputs(12709) <= (layer0_outputs(1787)) xor (layer0_outputs(4987));
    outputs(12710) <= (layer0_outputs(8990)) xor (layer0_outputs(2484));
    outputs(12711) <= (layer0_outputs(3355)) and not (layer0_outputs(2335));
    outputs(12712) <= layer0_outputs(5141);
    outputs(12713) <= not(layer0_outputs(10938));
    outputs(12714) <= layer0_outputs(10978);
    outputs(12715) <= (layer0_outputs(2990)) xor (layer0_outputs(2620));
    outputs(12716) <= (layer0_outputs(10546)) xor (layer0_outputs(11617));
    outputs(12717) <= not((layer0_outputs(2915)) and (layer0_outputs(7131)));
    outputs(12718) <= (layer0_outputs(348)) xor (layer0_outputs(1906));
    outputs(12719) <= layer0_outputs(6051);
    outputs(12720) <= not(layer0_outputs(1897));
    outputs(12721) <= layer0_outputs(4173);
    outputs(12722) <= not(layer0_outputs(2902));
    outputs(12723) <= (layer0_outputs(10053)) and not (layer0_outputs(705));
    outputs(12724) <= not(layer0_outputs(11385));
    outputs(12725) <= layer0_outputs(1738);
    outputs(12726) <= (layer0_outputs(7821)) and not (layer0_outputs(5841));
    outputs(12727) <= not(layer0_outputs(1019));
    outputs(12728) <= layer0_outputs(9129);
    outputs(12729) <= layer0_outputs(10902);
    outputs(12730) <= (layer0_outputs(3133)) xor (layer0_outputs(7615));
    outputs(12731) <= not(layer0_outputs(360)) or (layer0_outputs(2934));
    outputs(12732) <= not(layer0_outputs(2022));
    outputs(12733) <= (layer0_outputs(2078)) and (layer0_outputs(293));
    outputs(12734) <= not((layer0_outputs(10918)) and (layer0_outputs(4398)));
    outputs(12735) <= layer0_outputs(661);
    outputs(12736) <= not(layer0_outputs(5244));
    outputs(12737) <= layer0_outputs(8080);
    outputs(12738) <= layer0_outputs(12295);
    outputs(12739) <= (layer0_outputs(8098)) xor (layer0_outputs(10623));
    outputs(12740) <= not((layer0_outputs(2869)) xor (layer0_outputs(2816)));
    outputs(12741) <= not((layer0_outputs(8402)) xor (layer0_outputs(7992)));
    outputs(12742) <= not((layer0_outputs(818)) xor (layer0_outputs(10841)));
    outputs(12743) <= (layer0_outputs(8473)) and not (layer0_outputs(1590));
    outputs(12744) <= not(layer0_outputs(3520));
    outputs(12745) <= not((layer0_outputs(5854)) xor (layer0_outputs(83)));
    outputs(12746) <= (layer0_outputs(2871)) or (layer0_outputs(8299));
    outputs(12747) <= not(layer0_outputs(2862));
    outputs(12748) <= (layer0_outputs(9189)) xor (layer0_outputs(5385));
    outputs(12749) <= (layer0_outputs(4778)) xor (layer0_outputs(4009));
    outputs(12750) <= (layer0_outputs(8889)) xor (layer0_outputs(6543));
    outputs(12751) <= (layer0_outputs(3305)) xor (layer0_outputs(9197));
    outputs(12752) <= not((layer0_outputs(424)) xor (layer0_outputs(7371)));
    outputs(12753) <= (layer0_outputs(6112)) xor (layer0_outputs(4608));
    outputs(12754) <= not(layer0_outputs(6481)) or (layer0_outputs(11541));
    outputs(12755) <= not((layer0_outputs(9652)) xor (layer0_outputs(1321)));
    outputs(12756) <= not((layer0_outputs(7883)) or (layer0_outputs(9157)));
    outputs(12757) <= not((layer0_outputs(9424)) xor (layer0_outputs(10842)));
    outputs(12758) <= (layer0_outputs(371)) and (layer0_outputs(10015));
    outputs(12759) <= not(layer0_outputs(10681));
    outputs(12760) <= not(layer0_outputs(1718));
    outputs(12761) <= not(layer0_outputs(7547));
    outputs(12762) <= not((layer0_outputs(11060)) xor (layer0_outputs(7649)));
    outputs(12763) <= not((layer0_outputs(10030)) or (layer0_outputs(9182)));
    outputs(12764) <= not(layer0_outputs(3596)) or (layer0_outputs(4575));
    outputs(12765) <= layer0_outputs(3464);
    outputs(12766) <= not((layer0_outputs(7842)) xor (layer0_outputs(10257)));
    outputs(12767) <= not((layer0_outputs(9306)) xor (layer0_outputs(11855)));
    outputs(12768) <= (layer0_outputs(10853)) and (layer0_outputs(1934));
    outputs(12769) <= not((layer0_outputs(3006)) xor (layer0_outputs(2101)));
    outputs(12770) <= not((layer0_outputs(2411)) xor (layer0_outputs(9007)));
    outputs(12771) <= (layer0_outputs(6438)) xor (layer0_outputs(4463));
    outputs(12772) <= (layer0_outputs(222)) xor (layer0_outputs(309));
    outputs(12773) <= not(layer0_outputs(1157));
    outputs(12774) <= (layer0_outputs(5899)) xor (layer0_outputs(6776));
    outputs(12775) <= layer0_outputs(1805);
    outputs(12776) <= layer0_outputs(3383);
    outputs(12777) <= not((layer0_outputs(1010)) or (layer0_outputs(11850)));
    outputs(12778) <= not((layer0_outputs(6136)) xor (layer0_outputs(10952)));
    outputs(12779) <= layer0_outputs(11263);
    outputs(12780) <= (layer0_outputs(7805)) and not (layer0_outputs(1294));
    outputs(12781) <= not(layer0_outputs(10356)) or (layer0_outputs(5418));
    outputs(12782) <= not((layer0_outputs(6642)) or (layer0_outputs(5848)));
    outputs(12783) <= (layer0_outputs(6893)) and not (layer0_outputs(8567));
    outputs(12784) <= (layer0_outputs(1444)) and not (layer0_outputs(8168));
    outputs(12785) <= (layer0_outputs(617)) xor (layer0_outputs(3292));
    outputs(12786) <= (layer0_outputs(2197)) and not (layer0_outputs(9945));
    outputs(12787) <= (layer0_outputs(2460)) and not (layer0_outputs(7435));
    outputs(12788) <= not((layer0_outputs(6585)) xor (layer0_outputs(10813)));
    outputs(12789) <= '1';
    outputs(12790) <= not(layer0_outputs(4673));
    outputs(12791) <= (layer0_outputs(5518)) xor (layer0_outputs(864));
    outputs(12792) <= layer0_outputs(907);
    outputs(12793) <= not(layer0_outputs(11158));
    outputs(12794) <= layer0_outputs(361);
    outputs(12795) <= (layer0_outputs(5553)) xor (layer0_outputs(3685));
    outputs(12796) <= not(layer0_outputs(9113));
    outputs(12797) <= layer0_outputs(5902);
    outputs(12798) <= not((layer0_outputs(4746)) xor (layer0_outputs(885)));
    outputs(12799) <= not((layer0_outputs(9908)) xor (layer0_outputs(5381)));

end Behavioral;
