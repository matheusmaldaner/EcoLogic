library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(10239 downto 0);

begin

    layer0_outputs(0) <= not((inputs(100)) or (inputs(42)));
    layer0_outputs(1) <= not(inputs(235));
    layer0_outputs(2) <= not(inputs(246)) or (inputs(241));
    layer0_outputs(3) <= not(inputs(184)) or (inputs(146));
    layer0_outputs(4) <= not((inputs(162)) or (inputs(216)));
    layer0_outputs(5) <= not(inputs(94)) or (inputs(161));
    layer0_outputs(6) <= (inputs(133)) or (inputs(1));
    layer0_outputs(7) <= not((inputs(53)) xor (inputs(160)));
    layer0_outputs(8) <= not((inputs(189)) and (inputs(254)));
    layer0_outputs(9) <= (inputs(65)) or (inputs(227));
    layer0_outputs(10) <= not(inputs(168)) or (inputs(33));
    layer0_outputs(11) <= (inputs(75)) xor (inputs(18));
    layer0_outputs(12) <= not(inputs(58)) or (inputs(243));
    layer0_outputs(13) <= not((inputs(104)) or (inputs(253)));
    layer0_outputs(14) <= (inputs(213)) and not (inputs(103));
    layer0_outputs(15) <= not((inputs(160)) or (inputs(214)));
    layer0_outputs(16) <= not(inputs(46));
    layer0_outputs(17) <= inputs(0);
    layer0_outputs(18) <= not((inputs(109)) or (inputs(50)));
    layer0_outputs(19) <= (inputs(175)) and not (inputs(141));
    layer0_outputs(20) <= (inputs(229)) and not (inputs(130));
    layer0_outputs(21) <= not(inputs(212)) or (inputs(46));
    layer0_outputs(22) <= not((inputs(100)) and (inputs(135)));
    layer0_outputs(23) <= (inputs(115)) and (inputs(112));
    layer0_outputs(24) <= (inputs(227)) and not (inputs(113));
    layer0_outputs(25) <= not(inputs(236)) or (inputs(15));
    layer0_outputs(26) <= (inputs(123)) and (inputs(48));
    layer0_outputs(27) <= (inputs(187)) or (inputs(62));
    layer0_outputs(28) <= (inputs(10)) and not (inputs(192));
    layer0_outputs(29) <= (inputs(220)) xor (inputs(64));
    layer0_outputs(30) <= inputs(215);
    layer0_outputs(31) <= not((inputs(63)) or (inputs(83)));
    layer0_outputs(32) <= (inputs(200)) or (inputs(155));
    layer0_outputs(33) <= inputs(94);
    layer0_outputs(34) <= (inputs(57)) or (inputs(34));
    layer0_outputs(35) <= not((inputs(60)) or (inputs(15)));
    layer0_outputs(36) <= not(inputs(74)) or (inputs(96));
    layer0_outputs(37) <= not((inputs(116)) or (inputs(188)));
    layer0_outputs(38) <= '0';
    layer0_outputs(39) <= inputs(119);
    layer0_outputs(40) <= (inputs(180)) and not (inputs(66));
    layer0_outputs(41) <= (inputs(41)) or (inputs(247));
    layer0_outputs(42) <= not(inputs(164));
    layer0_outputs(43) <= (inputs(171)) or (inputs(140));
    layer0_outputs(44) <= not(inputs(179));
    layer0_outputs(45) <= not((inputs(139)) or (inputs(188)));
    layer0_outputs(46) <= not(inputs(228));
    layer0_outputs(47) <= not(inputs(14));
    layer0_outputs(48) <= not(inputs(16)) or (inputs(242));
    layer0_outputs(49) <= not(inputs(28)) or (inputs(206));
    layer0_outputs(50) <= not(inputs(14)) or (inputs(171));
    layer0_outputs(51) <= not(inputs(152)) or (inputs(203));
    layer0_outputs(52) <= (inputs(170)) and not (inputs(213));
    layer0_outputs(53) <= (inputs(196)) or (inputs(203));
    layer0_outputs(54) <= not((inputs(98)) or (inputs(137)));
    layer0_outputs(55) <= not(inputs(17));
    layer0_outputs(56) <= not(inputs(228));
    layer0_outputs(57) <= not(inputs(23)) or (inputs(125));
    layer0_outputs(58) <= not(inputs(159));
    layer0_outputs(59) <= not((inputs(237)) xor (inputs(181)));
    layer0_outputs(60) <= not((inputs(8)) or (inputs(107)));
    layer0_outputs(61) <= not((inputs(182)) xor (inputs(152)));
    layer0_outputs(62) <= (inputs(105)) and not (inputs(176));
    layer0_outputs(63) <= (inputs(221)) or (inputs(160));
    layer0_outputs(64) <= not(inputs(32)) or (inputs(244));
    layer0_outputs(65) <= (inputs(244)) and not (inputs(158));
    layer0_outputs(66) <= inputs(197);
    layer0_outputs(67) <= not(inputs(3));
    layer0_outputs(68) <= not((inputs(165)) or (inputs(145)));
    layer0_outputs(69) <= (inputs(21)) or (inputs(84));
    layer0_outputs(70) <= not(inputs(72));
    layer0_outputs(71) <= not((inputs(54)) or (inputs(140)));
    layer0_outputs(72) <= not((inputs(233)) and (inputs(174)));
    layer0_outputs(73) <= inputs(98);
    layer0_outputs(74) <= not((inputs(155)) xor (inputs(178)));
    layer0_outputs(75) <= inputs(119);
    layer0_outputs(76) <= inputs(193);
    layer0_outputs(77) <= inputs(92);
    layer0_outputs(78) <= not(inputs(248)) or (inputs(235));
    layer0_outputs(79) <= (inputs(228)) or (inputs(128));
    layer0_outputs(80) <= not(inputs(11));
    layer0_outputs(81) <= not(inputs(95));
    layer0_outputs(82) <= inputs(153);
    layer0_outputs(83) <= not((inputs(108)) xor (inputs(103)));
    layer0_outputs(84) <= not((inputs(155)) xor (inputs(124)));
    layer0_outputs(85) <= not((inputs(19)) or (inputs(33)));
    layer0_outputs(86) <= not(inputs(109));
    layer0_outputs(87) <= (inputs(251)) and not (inputs(72));
    layer0_outputs(88) <= (inputs(61)) or (inputs(89));
    layer0_outputs(89) <= (inputs(62)) or (inputs(54));
    layer0_outputs(90) <= (inputs(139)) or (inputs(252));
    layer0_outputs(91) <= '1';
    layer0_outputs(92) <= not(inputs(49));
    layer0_outputs(93) <= not((inputs(210)) or (inputs(0)));
    layer0_outputs(94) <= (inputs(165)) xor (inputs(177));
    layer0_outputs(95) <= not((inputs(209)) or (inputs(21)));
    layer0_outputs(96) <= (inputs(89)) xor (inputs(153));
    layer0_outputs(97) <= (inputs(27)) and not (inputs(191));
    layer0_outputs(98) <= not(inputs(108));
    layer0_outputs(99) <= not((inputs(99)) or (inputs(15)));
    layer0_outputs(100) <= (inputs(116)) and (inputs(93));
    layer0_outputs(101) <= not((inputs(39)) or (inputs(9)));
    layer0_outputs(102) <= (inputs(26)) xor (inputs(207));
    layer0_outputs(103) <= inputs(247);
    layer0_outputs(104) <= not((inputs(52)) xor (inputs(114)));
    layer0_outputs(105) <= not((inputs(111)) or (inputs(50)));
    layer0_outputs(106) <= not((inputs(238)) or (inputs(72)));
    layer0_outputs(107) <= not(inputs(97));
    layer0_outputs(108) <= (inputs(12)) xor (inputs(141));
    layer0_outputs(109) <= not(inputs(170)) or (inputs(151));
    layer0_outputs(110) <= inputs(217);
    layer0_outputs(111) <= inputs(230);
    layer0_outputs(112) <= inputs(166);
    layer0_outputs(113) <= not(inputs(245)) or (inputs(153));
    layer0_outputs(114) <= (inputs(28)) or (inputs(73));
    layer0_outputs(115) <= (inputs(137)) and not (inputs(158));
    layer0_outputs(116) <= inputs(44);
    layer0_outputs(117) <= not(inputs(99)) or (inputs(27));
    layer0_outputs(118) <= inputs(114);
    layer0_outputs(119) <= not((inputs(165)) or (inputs(253)));
    layer0_outputs(120) <= (inputs(21)) xor (inputs(85));
    layer0_outputs(121) <= (inputs(51)) and not (inputs(191));
    layer0_outputs(122) <= not(inputs(42)) or (inputs(157));
    layer0_outputs(123) <= (inputs(120)) and not (inputs(95));
    layer0_outputs(124) <= not((inputs(125)) xor (inputs(122)));
    layer0_outputs(125) <= inputs(224);
    layer0_outputs(126) <= not(inputs(98)) or (inputs(190));
    layer0_outputs(127) <= not((inputs(207)) xor (inputs(60)));
    layer0_outputs(128) <= (inputs(235)) xor (inputs(124));
    layer0_outputs(129) <= (inputs(3)) or (inputs(136));
    layer0_outputs(130) <= '0';
    layer0_outputs(131) <= not(inputs(125));
    layer0_outputs(132) <= not((inputs(42)) or (inputs(4)));
    layer0_outputs(133) <= not((inputs(66)) or (inputs(204)));
    layer0_outputs(134) <= not((inputs(51)) and (inputs(102)));
    layer0_outputs(135) <= not(inputs(152)) or (inputs(159));
    layer0_outputs(136) <= not(inputs(179));
    layer0_outputs(137) <= (inputs(62)) and not (inputs(117));
    layer0_outputs(138) <= inputs(132);
    layer0_outputs(139) <= not((inputs(204)) xor (inputs(124)));
    layer0_outputs(140) <= not((inputs(48)) or (inputs(167)));
    layer0_outputs(141) <= not((inputs(42)) xor (inputs(102)));
    layer0_outputs(142) <= not((inputs(244)) xor (inputs(250)));
    layer0_outputs(143) <= not(inputs(166));
    layer0_outputs(144) <= (inputs(38)) and not (inputs(235));
    layer0_outputs(145) <= not((inputs(129)) xor (inputs(39)));
    layer0_outputs(146) <= inputs(73);
    layer0_outputs(147) <= (inputs(213)) xor (inputs(38));
    layer0_outputs(148) <= inputs(185);
    layer0_outputs(149) <= inputs(140);
    layer0_outputs(150) <= not(inputs(175));
    layer0_outputs(151) <= not((inputs(25)) or (inputs(49)));
    layer0_outputs(152) <= not(inputs(43)) or (inputs(46));
    layer0_outputs(153) <= not(inputs(138));
    layer0_outputs(154) <= not(inputs(206)) or (inputs(174));
    layer0_outputs(155) <= (inputs(248)) or (inputs(144));
    layer0_outputs(156) <= not((inputs(85)) xor (inputs(145)));
    layer0_outputs(157) <= not(inputs(170)) or (inputs(44));
    layer0_outputs(158) <= '0';
    layer0_outputs(159) <= (inputs(180)) and (inputs(70));
    layer0_outputs(160) <= not(inputs(245)) or (inputs(150));
    layer0_outputs(161) <= inputs(21);
    layer0_outputs(162) <= (inputs(153)) and not (inputs(193));
    layer0_outputs(163) <= inputs(67);
    layer0_outputs(164) <= not((inputs(147)) or (inputs(152)));
    layer0_outputs(165) <= not((inputs(242)) xor (inputs(179)));
    layer0_outputs(166) <= not((inputs(212)) or (inputs(60)));
    layer0_outputs(167) <= inputs(213);
    layer0_outputs(168) <= (inputs(60)) or (inputs(192));
    layer0_outputs(169) <= not(inputs(106));
    layer0_outputs(170) <= not((inputs(16)) or (inputs(40)));
    layer0_outputs(171) <= (inputs(125)) and (inputs(123));
    layer0_outputs(172) <= (inputs(237)) or (inputs(160));
    layer0_outputs(173) <= inputs(128);
    layer0_outputs(174) <= (inputs(225)) and not (inputs(79));
    layer0_outputs(175) <= (inputs(130)) or (inputs(237));
    layer0_outputs(176) <= inputs(41);
    layer0_outputs(177) <= not((inputs(185)) or (inputs(144)));
    layer0_outputs(178) <= '0';
    layer0_outputs(179) <= (inputs(104)) and (inputs(33));
    layer0_outputs(180) <= not(inputs(254)) or (inputs(156));
    layer0_outputs(181) <= (inputs(155)) xor (inputs(148));
    layer0_outputs(182) <= inputs(132);
    layer0_outputs(183) <= (inputs(214)) or (inputs(129));
    layer0_outputs(184) <= not((inputs(64)) or (inputs(180)));
    layer0_outputs(185) <= not(inputs(178));
    layer0_outputs(186) <= not((inputs(145)) or (inputs(80)));
    layer0_outputs(187) <= inputs(120);
    layer0_outputs(188) <= (inputs(213)) and not (inputs(53));
    layer0_outputs(189) <= inputs(122);
    layer0_outputs(190) <= (inputs(90)) or (inputs(21));
    layer0_outputs(191) <= (inputs(222)) and not (inputs(206));
    layer0_outputs(192) <= (inputs(102)) or (inputs(43));
    layer0_outputs(193) <= inputs(117);
    layer0_outputs(194) <= not((inputs(158)) or (inputs(47)));
    layer0_outputs(195) <= not((inputs(45)) or (inputs(110)));
    layer0_outputs(196) <= (inputs(37)) or (inputs(22));
    layer0_outputs(197) <= not((inputs(66)) or (inputs(14)));
    layer0_outputs(198) <= not((inputs(50)) xor (inputs(221)));
    layer0_outputs(199) <= not(inputs(84));
    layer0_outputs(200) <= not(inputs(8)) or (inputs(39));
    layer0_outputs(201) <= inputs(214);
    layer0_outputs(202) <= not((inputs(199)) xor (inputs(200)));
    layer0_outputs(203) <= inputs(152);
    layer0_outputs(204) <= inputs(214);
    layer0_outputs(205) <= not(inputs(56)) or (inputs(81));
    layer0_outputs(206) <= not((inputs(152)) xor (inputs(201)));
    layer0_outputs(207) <= (inputs(179)) xor (inputs(35));
    layer0_outputs(208) <= not((inputs(134)) or (inputs(122)));
    layer0_outputs(209) <= not((inputs(121)) or (inputs(192)));
    layer0_outputs(210) <= (inputs(231)) xor (inputs(152));
    layer0_outputs(211) <= '0';
    layer0_outputs(212) <= (inputs(146)) or (inputs(196));
    layer0_outputs(213) <= not(inputs(242));
    layer0_outputs(214) <= (inputs(231)) and not (inputs(64));
    layer0_outputs(215) <= (inputs(125)) and not (inputs(198));
    layer0_outputs(216) <= not(inputs(237));
    layer0_outputs(217) <= '1';
    layer0_outputs(218) <= (inputs(154)) and (inputs(160));
    layer0_outputs(219) <= not((inputs(49)) or (inputs(254)));
    layer0_outputs(220) <= '0';
    layer0_outputs(221) <= not(inputs(92));
    layer0_outputs(222) <= not((inputs(44)) xor (inputs(231)));
    layer0_outputs(223) <= not((inputs(129)) xor (inputs(185)));
    layer0_outputs(224) <= (inputs(42)) or (inputs(208));
    layer0_outputs(225) <= (inputs(13)) or (inputs(237));
    layer0_outputs(226) <= (inputs(182)) xor (inputs(138));
    layer0_outputs(227) <= not(inputs(218)) or (inputs(31));
    layer0_outputs(228) <= (inputs(220)) and not (inputs(97));
    layer0_outputs(229) <= (inputs(143)) or (inputs(223));
    layer0_outputs(230) <= inputs(213);
    layer0_outputs(231) <= (inputs(62)) and not (inputs(139));
    layer0_outputs(232) <= (inputs(167)) and not (inputs(211));
    layer0_outputs(233) <= (inputs(121)) and (inputs(153));
    layer0_outputs(234) <= not((inputs(59)) or (inputs(4)));
    layer0_outputs(235) <= not(inputs(244)) or (inputs(168));
    layer0_outputs(236) <= (inputs(163)) or (inputs(206));
    layer0_outputs(237) <= not(inputs(56)) or (inputs(50));
    layer0_outputs(238) <= not((inputs(117)) xor (inputs(174)));
    layer0_outputs(239) <= '1';
    layer0_outputs(240) <= not(inputs(3));
    layer0_outputs(241) <= inputs(72);
    layer0_outputs(242) <= inputs(174);
    layer0_outputs(243) <= (inputs(94)) xor (inputs(187));
    layer0_outputs(244) <= not((inputs(213)) or (inputs(229)));
    layer0_outputs(245) <= not((inputs(161)) xor (inputs(130)));
    layer0_outputs(246) <= (inputs(193)) or (inputs(210));
    layer0_outputs(247) <= not((inputs(144)) or (inputs(220)));
    layer0_outputs(248) <= not((inputs(36)) or (inputs(167)));
    layer0_outputs(249) <= inputs(21);
    layer0_outputs(250) <= (inputs(70)) xor (inputs(90));
    layer0_outputs(251) <= not(inputs(40)) or (inputs(217));
    layer0_outputs(252) <= not(inputs(224)) or (inputs(19));
    layer0_outputs(253) <= not((inputs(124)) or (inputs(96)));
    layer0_outputs(254) <= not((inputs(216)) xor (inputs(148)));
    layer0_outputs(255) <= (inputs(226)) or (inputs(233));
    layer0_outputs(256) <= (inputs(215)) and not (inputs(46));
    layer0_outputs(257) <= not((inputs(65)) xor (inputs(204)));
    layer0_outputs(258) <= inputs(84);
    layer0_outputs(259) <= (inputs(230)) and not (inputs(121));
    layer0_outputs(260) <= (inputs(159)) xor (inputs(218));
    layer0_outputs(261) <= inputs(200);
    layer0_outputs(262) <= inputs(122);
    layer0_outputs(263) <= (inputs(69)) xor (inputs(81));
    layer0_outputs(264) <= not(inputs(114)) or (inputs(233));
    layer0_outputs(265) <= inputs(18);
    layer0_outputs(266) <= not((inputs(31)) or (inputs(234)));
    layer0_outputs(267) <= (inputs(141)) xor (inputs(29));
    layer0_outputs(268) <= inputs(252);
    layer0_outputs(269) <= inputs(90);
    layer0_outputs(270) <= not(inputs(60));
    layer0_outputs(271) <= not(inputs(226));
    layer0_outputs(272) <= not((inputs(111)) xor (inputs(88)));
    layer0_outputs(273) <= inputs(194);
    layer0_outputs(274) <= not(inputs(90));
    layer0_outputs(275) <= not(inputs(233));
    layer0_outputs(276) <= not(inputs(17)) or (inputs(175));
    layer0_outputs(277) <= not((inputs(3)) or (inputs(3)));
    layer0_outputs(278) <= inputs(50);
    layer0_outputs(279) <= '0';
    layer0_outputs(280) <= not(inputs(22)) or (inputs(161));
    layer0_outputs(281) <= inputs(27);
    layer0_outputs(282) <= inputs(8);
    layer0_outputs(283) <= not((inputs(55)) xor (inputs(8)));
    layer0_outputs(284) <= not(inputs(118));
    layer0_outputs(285) <= (inputs(238)) and (inputs(140));
    layer0_outputs(286) <= (inputs(4)) or (inputs(188));
    layer0_outputs(287) <= not(inputs(193)) or (inputs(71));
    layer0_outputs(288) <= '0';
    layer0_outputs(289) <= not(inputs(250)) or (inputs(185));
    layer0_outputs(290) <= not(inputs(126)) or (inputs(93));
    layer0_outputs(291) <= not(inputs(187)) or (inputs(134));
    layer0_outputs(292) <= inputs(40);
    layer0_outputs(293) <= not(inputs(38));
    layer0_outputs(294) <= (inputs(102)) xor (inputs(52));
    layer0_outputs(295) <= not(inputs(14));
    layer0_outputs(296) <= not((inputs(158)) xor (inputs(218)));
    layer0_outputs(297) <= (inputs(144)) xor (inputs(198));
    layer0_outputs(298) <= not(inputs(36));
    layer0_outputs(299) <= not((inputs(99)) xor (inputs(82)));
    layer0_outputs(300) <= not((inputs(24)) or (inputs(211)));
    layer0_outputs(301) <= (inputs(226)) or (inputs(207));
    layer0_outputs(302) <= not((inputs(221)) or (inputs(212)));
    layer0_outputs(303) <= inputs(31);
    layer0_outputs(304) <= not((inputs(172)) or (inputs(215)));
    layer0_outputs(305) <= not(inputs(202));
    layer0_outputs(306) <= not(inputs(167)) or (inputs(79));
    layer0_outputs(307) <= not((inputs(244)) or (inputs(172)));
    layer0_outputs(308) <= inputs(241);
    layer0_outputs(309) <= inputs(121);
    layer0_outputs(310) <= (inputs(5)) or (inputs(78));
    layer0_outputs(311) <= (inputs(231)) and not (inputs(31));
    layer0_outputs(312) <= (inputs(88)) and not (inputs(224));
    layer0_outputs(313) <= inputs(15);
    layer0_outputs(314) <= (inputs(191)) xor (inputs(183));
    layer0_outputs(315) <= (inputs(102)) and not (inputs(125));
    layer0_outputs(316) <= not(inputs(153));
    layer0_outputs(317) <= (inputs(111)) or (inputs(94));
    layer0_outputs(318) <= (inputs(29)) or (inputs(16));
    layer0_outputs(319) <= not(inputs(116));
    layer0_outputs(320) <= (inputs(124)) or (inputs(4));
    layer0_outputs(321) <= not(inputs(178));
    layer0_outputs(322) <= not(inputs(177));
    layer0_outputs(323) <= inputs(33);
    layer0_outputs(324) <= inputs(105);
    layer0_outputs(325) <= not((inputs(39)) or (inputs(48)));
    layer0_outputs(326) <= inputs(213);
    layer0_outputs(327) <= not(inputs(86)) or (inputs(188));
    layer0_outputs(328) <= not(inputs(21));
    layer0_outputs(329) <= (inputs(117)) xor (inputs(221));
    layer0_outputs(330) <= (inputs(5)) xor (inputs(70));
    layer0_outputs(331) <= not((inputs(1)) or (inputs(120)));
    layer0_outputs(332) <= not((inputs(143)) or (inputs(243)));
    layer0_outputs(333) <= (inputs(71)) and not (inputs(18));
    layer0_outputs(334) <= not((inputs(98)) xor (inputs(81)));
    layer0_outputs(335) <= (inputs(74)) or (inputs(129));
    layer0_outputs(336) <= (inputs(168)) or (inputs(253));
    layer0_outputs(337) <= (inputs(18)) or (inputs(34));
    layer0_outputs(338) <= (inputs(132)) and not (inputs(227));
    layer0_outputs(339) <= (inputs(144)) xor (inputs(181));
    layer0_outputs(340) <= '0';
    layer0_outputs(341) <= inputs(128);
    layer0_outputs(342) <= not(inputs(202));
    layer0_outputs(343) <= inputs(100);
    layer0_outputs(344) <= not((inputs(119)) and (inputs(9)));
    layer0_outputs(345) <= (inputs(217)) and not (inputs(235));
    layer0_outputs(346) <= not(inputs(85));
    layer0_outputs(347) <= (inputs(239)) or (inputs(238));
    layer0_outputs(348) <= inputs(49);
    layer0_outputs(349) <= (inputs(84)) or (inputs(45));
    layer0_outputs(350) <= inputs(105);
    layer0_outputs(351) <= not(inputs(254)) or (inputs(252));
    layer0_outputs(352) <= (inputs(105)) and not (inputs(34));
    layer0_outputs(353) <= (inputs(8)) and not (inputs(244));
    layer0_outputs(354) <= not((inputs(59)) xor (inputs(33)));
    layer0_outputs(355) <= not((inputs(137)) or (inputs(153)));
    layer0_outputs(356) <= not(inputs(129)) or (inputs(102));
    layer0_outputs(357) <= not((inputs(122)) xor (inputs(157)));
    layer0_outputs(358) <= (inputs(225)) or (inputs(197));
    layer0_outputs(359) <= inputs(132);
    layer0_outputs(360) <= not((inputs(24)) and (inputs(72)));
    layer0_outputs(361) <= not(inputs(57));
    layer0_outputs(362) <= not((inputs(211)) or (inputs(188)));
    layer0_outputs(363) <= not(inputs(58));
    layer0_outputs(364) <= not((inputs(68)) xor (inputs(80)));
    layer0_outputs(365) <= not(inputs(84));
    layer0_outputs(366) <= not((inputs(234)) xor (inputs(206)));
    layer0_outputs(367) <= not(inputs(73));
    layer0_outputs(368) <= inputs(192);
    layer0_outputs(369) <= not(inputs(82));
    layer0_outputs(370) <= not(inputs(227));
    layer0_outputs(371) <= (inputs(206)) or (inputs(109));
    layer0_outputs(372) <= inputs(50);
    layer0_outputs(373) <= not((inputs(193)) xor (inputs(58)));
    layer0_outputs(374) <= (inputs(156)) and not (inputs(252));
    layer0_outputs(375) <= not((inputs(197)) or (inputs(82)));
    layer0_outputs(376) <= (inputs(182)) or (inputs(34));
    layer0_outputs(377) <= not(inputs(174));
    layer0_outputs(378) <= not((inputs(24)) xor (inputs(191)));
    layer0_outputs(379) <= not(inputs(83)) or (inputs(65));
    layer0_outputs(380) <= (inputs(61)) and not (inputs(113));
    layer0_outputs(381) <= not((inputs(21)) xor (inputs(142)));
    layer0_outputs(382) <= (inputs(136)) and not (inputs(202));
    layer0_outputs(383) <= inputs(110);
    layer0_outputs(384) <= not(inputs(77));
    layer0_outputs(385) <= inputs(150);
    layer0_outputs(386) <= not(inputs(26)) or (inputs(216));
    layer0_outputs(387) <= not((inputs(108)) xor (inputs(111)));
    layer0_outputs(388) <= not((inputs(18)) or (inputs(152)));
    layer0_outputs(389) <= not((inputs(255)) or (inputs(192)));
    layer0_outputs(390) <= not(inputs(210));
    layer0_outputs(391) <= (inputs(31)) and (inputs(211));
    layer0_outputs(392) <= not(inputs(155)) or (inputs(131));
    layer0_outputs(393) <= not((inputs(133)) and (inputs(68)));
    layer0_outputs(394) <= (inputs(39)) and not (inputs(161));
    layer0_outputs(395) <= not(inputs(111)) or (inputs(253));
    layer0_outputs(396) <= not((inputs(126)) or (inputs(179)));
    layer0_outputs(397) <= not((inputs(20)) xor (inputs(159)));
    layer0_outputs(398) <= inputs(189);
    layer0_outputs(399) <= inputs(165);
    layer0_outputs(400) <= not((inputs(99)) or (inputs(3)));
    layer0_outputs(401) <= not(inputs(53));
    layer0_outputs(402) <= (inputs(38)) and (inputs(69));
    layer0_outputs(403) <= not((inputs(87)) xor (inputs(60)));
    layer0_outputs(404) <= (inputs(136)) or (inputs(43));
    layer0_outputs(405) <= (inputs(234)) and not (inputs(126));
    layer0_outputs(406) <= not(inputs(104));
    layer0_outputs(407) <= not(inputs(132));
    layer0_outputs(408) <= not((inputs(168)) or (inputs(236)));
    layer0_outputs(409) <= not((inputs(8)) and (inputs(133)));
    layer0_outputs(410) <= not((inputs(183)) or (inputs(63)));
    layer0_outputs(411) <= not(inputs(116));
    layer0_outputs(412) <= '0';
    layer0_outputs(413) <= '1';
    layer0_outputs(414) <= (inputs(160)) or (inputs(179));
    layer0_outputs(415) <= not((inputs(251)) or (inputs(185)));
    layer0_outputs(416) <= (inputs(40)) or (inputs(109));
    layer0_outputs(417) <= not((inputs(113)) xor (inputs(16)));
    layer0_outputs(418) <= not((inputs(174)) and (inputs(159)));
    layer0_outputs(419) <= not(inputs(150));
    layer0_outputs(420) <= (inputs(209)) and not (inputs(205));
    layer0_outputs(421) <= not((inputs(104)) or (inputs(208)));
    layer0_outputs(422) <= not(inputs(53)) or (inputs(190));
    layer0_outputs(423) <= not((inputs(135)) xor (inputs(194)));
    layer0_outputs(424) <= (inputs(70)) xor (inputs(33));
    layer0_outputs(425) <= not((inputs(198)) or (inputs(185)));
    layer0_outputs(426) <= not(inputs(120));
    layer0_outputs(427) <= (inputs(183)) and (inputs(108));
    layer0_outputs(428) <= (inputs(180)) and not (inputs(74));
    layer0_outputs(429) <= not((inputs(187)) xor (inputs(241)));
    layer0_outputs(430) <= (inputs(178)) and not (inputs(43));
    layer0_outputs(431) <= (inputs(165)) xor (inputs(146));
    layer0_outputs(432) <= not(inputs(83)) or (inputs(72));
    layer0_outputs(433) <= (inputs(44)) and not (inputs(15));
    layer0_outputs(434) <= (inputs(140)) and (inputs(139));
    layer0_outputs(435) <= not((inputs(131)) xor (inputs(100)));
    layer0_outputs(436) <= not((inputs(216)) and (inputs(187)));
    layer0_outputs(437) <= (inputs(214)) and not (inputs(96));
    layer0_outputs(438) <= not(inputs(252));
    layer0_outputs(439) <= not(inputs(245)) or (inputs(15));
    layer0_outputs(440) <= (inputs(72)) and (inputs(44));
    layer0_outputs(441) <= not((inputs(60)) or (inputs(130)));
    layer0_outputs(442) <= (inputs(173)) or (inputs(80));
    layer0_outputs(443) <= inputs(154);
    layer0_outputs(444) <= not((inputs(143)) or (inputs(225)));
    layer0_outputs(445) <= not((inputs(213)) or (inputs(37)));
    layer0_outputs(446) <= not((inputs(184)) and (inputs(201)));
    layer0_outputs(447) <= not(inputs(188));
    layer0_outputs(448) <= not((inputs(2)) and (inputs(175)));
    layer0_outputs(449) <= (inputs(10)) or (inputs(0));
    layer0_outputs(450) <= not(inputs(93));
    layer0_outputs(451) <= '1';
    layer0_outputs(452) <= (inputs(61)) and (inputs(20));
    layer0_outputs(453) <= not((inputs(132)) or (inputs(186)));
    layer0_outputs(454) <= inputs(171);
    layer0_outputs(455) <= not((inputs(177)) or (inputs(194)));
    layer0_outputs(456) <= not(inputs(145)) or (inputs(57));
    layer0_outputs(457) <= not(inputs(228));
    layer0_outputs(458) <= inputs(30);
    layer0_outputs(459) <= not(inputs(120));
    layer0_outputs(460) <= inputs(180);
    layer0_outputs(461) <= not((inputs(133)) or (inputs(101)));
    layer0_outputs(462) <= not((inputs(207)) or (inputs(220)));
    layer0_outputs(463) <= not((inputs(142)) or (inputs(79)));
    layer0_outputs(464) <= (inputs(106)) xor (inputs(232));
    layer0_outputs(465) <= inputs(100);
    layer0_outputs(466) <= inputs(25);
    layer0_outputs(467) <= (inputs(70)) xor (inputs(65));
    layer0_outputs(468) <= not((inputs(223)) or (inputs(5)));
    layer0_outputs(469) <= inputs(215);
    layer0_outputs(470) <= inputs(22);
    layer0_outputs(471) <= not(inputs(221));
    layer0_outputs(472) <= not((inputs(191)) or (inputs(176)));
    layer0_outputs(473) <= inputs(34);
    layer0_outputs(474) <= not(inputs(213));
    layer0_outputs(475) <= not(inputs(132)) or (inputs(48));
    layer0_outputs(476) <= not((inputs(82)) or (inputs(111)));
    layer0_outputs(477) <= not(inputs(217));
    layer0_outputs(478) <= inputs(233);
    layer0_outputs(479) <= not((inputs(9)) xor (inputs(4)));
    layer0_outputs(480) <= not((inputs(161)) xor (inputs(245)));
    layer0_outputs(481) <= (inputs(244)) and (inputs(55));
    layer0_outputs(482) <= (inputs(245)) and not (inputs(48));
    layer0_outputs(483) <= not((inputs(225)) or (inputs(64)));
    layer0_outputs(484) <= (inputs(227)) and not (inputs(20));
    layer0_outputs(485) <= inputs(89);
    layer0_outputs(486) <= (inputs(22)) or (inputs(123));
    layer0_outputs(487) <= not(inputs(153));
    layer0_outputs(488) <= not(inputs(152));
    layer0_outputs(489) <= '1';
    layer0_outputs(490) <= not((inputs(147)) or (inputs(232)));
    layer0_outputs(491) <= inputs(68);
    layer0_outputs(492) <= not((inputs(230)) or (inputs(228)));
    layer0_outputs(493) <= not((inputs(144)) xor (inputs(81)));
    layer0_outputs(494) <= (inputs(103)) and not (inputs(199));
    layer0_outputs(495) <= (inputs(245)) and (inputs(11));
    layer0_outputs(496) <= not(inputs(123));
    layer0_outputs(497) <= (inputs(107)) and not (inputs(235));
    layer0_outputs(498) <= not(inputs(210)) or (inputs(48));
    layer0_outputs(499) <= inputs(24);
    layer0_outputs(500) <= not((inputs(47)) xor (inputs(238)));
    layer0_outputs(501) <= not((inputs(87)) xor (inputs(115)));
    layer0_outputs(502) <= not((inputs(135)) xor (inputs(36)));
    layer0_outputs(503) <= inputs(165);
    layer0_outputs(504) <= inputs(215);
    layer0_outputs(505) <= not(inputs(6)) or (inputs(214));
    layer0_outputs(506) <= not(inputs(89));
    layer0_outputs(507) <= '1';
    layer0_outputs(508) <= (inputs(176)) xor (inputs(144));
    layer0_outputs(509) <= inputs(152);
    layer0_outputs(510) <= (inputs(170)) and not (inputs(249));
    layer0_outputs(511) <= (inputs(112)) xor (inputs(219));
    layer0_outputs(512) <= not(inputs(19));
    layer0_outputs(513) <= inputs(90);
    layer0_outputs(514) <= (inputs(252)) and (inputs(159));
    layer0_outputs(515) <= not(inputs(242));
    layer0_outputs(516) <= (inputs(17)) and not (inputs(175));
    layer0_outputs(517) <= (inputs(249)) or (inputs(94));
    layer0_outputs(518) <= not(inputs(70)) or (inputs(173));
    layer0_outputs(519) <= not(inputs(163));
    layer0_outputs(520) <= not(inputs(231));
    layer0_outputs(521) <= (inputs(145)) or (inputs(91));
    layer0_outputs(522) <= (inputs(76)) and not (inputs(30));
    layer0_outputs(523) <= not((inputs(233)) xor (inputs(168)));
    layer0_outputs(524) <= (inputs(170)) xor (inputs(122));
    layer0_outputs(525) <= not(inputs(3)) or (inputs(161));
    layer0_outputs(526) <= (inputs(136)) and not (inputs(64));
    layer0_outputs(527) <= not((inputs(79)) xor (inputs(91)));
    layer0_outputs(528) <= (inputs(189)) or (inputs(130));
    layer0_outputs(529) <= (inputs(148)) and not (inputs(202));
    layer0_outputs(530) <= not((inputs(147)) xor (inputs(67)));
    layer0_outputs(531) <= not(inputs(73));
    layer0_outputs(532) <= not(inputs(125));
    layer0_outputs(533) <= not(inputs(0));
    layer0_outputs(534) <= inputs(215);
    layer0_outputs(535) <= inputs(130);
    layer0_outputs(536) <= (inputs(154)) or (inputs(45));
    layer0_outputs(537) <= not((inputs(178)) or (inputs(207)));
    layer0_outputs(538) <= (inputs(40)) or (inputs(116));
    layer0_outputs(539) <= not(inputs(31));
    layer0_outputs(540) <= not((inputs(141)) or (inputs(26)));
    layer0_outputs(541) <= not((inputs(210)) or (inputs(95)));
    layer0_outputs(542) <= (inputs(78)) and not (inputs(2));
    layer0_outputs(543) <= not((inputs(167)) or (inputs(151)));
    layer0_outputs(544) <= inputs(200);
    layer0_outputs(545) <= not((inputs(237)) or (inputs(29)));
    layer0_outputs(546) <= (inputs(150)) and not (inputs(99));
    layer0_outputs(547) <= inputs(141);
    layer0_outputs(548) <= not(inputs(200));
    layer0_outputs(549) <= not(inputs(20));
    layer0_outputs(550) <= not(inputs(187));
    layer0_outputs(551) <= (inputs(129)) xor (inputs(83));
    layer0_outputs(552) <= not((inputs(155)) or (inputs(84)));
    layer0_outputs(553) <= (inputs(186)) and not (inputs(3));
    layer0_outputs(554) <= (inputs(216)) and not (inputs(105));
    layer0_outputs(555) <= (inputs(167)) and not (inputs(5));
    layer0_outputs(556) <= (inputs(1)) and not (inputs(4));
    layer0_outputs(557) <= '0';
    layer0_outputs(558) <= (inputs(25)) and not (inputs(225));
    layer0_outputs(559) <= (inputs(8)) xor (inputs(47));
    layer0_outputs(560) <= not((inputs(216)) or (inputs(171)));
    layer0_outputs(561) <= inputs(131);
    layer0_outputs(562) <= (inputs(176)) or (inputs(60));
    layer0_outputs(563) <= inputs(42);
    layer0_outputs(564) <= not(inputs(182));
    layer0_outputs(565) <= (inputs(80)) or (inputs(172));
    layer0_outputs(566) <= not(inputs(122));
    layer0_outputs(567) <= inputs(47);
    layer0_outputs(568) <= not(inputs(198)) or (inputs(192));
    layer0_outputs(569) <= not(inputs(153)) or (inputs(118));
    layer0_outputs(570) <= not((inputs(50)) and (inputs(89)));
    layer0_outputs(571) <= inputs(38);
    layer0_outputs(572) <= (inputs(239)) xor (inputs(132));
    layer0_outputs(573) <= not(inputs(21)) or (inputs(29));
    layer0_outputs(574) <= not((inputs(100)) xor (inputs(147)));
    layer0_outputs(575) <= not(inputs(37));
    layer0_outputs(576) <= (inputs(177)) or (inputs(165));
    layer0_outputs(577) <= inputs(85);
    layer0_outputs(578) <= (inputs(84)) and not (inputs(109));
    layer0_outputs(579) <= inputs(205);
    layer0_outputs(580) <= not(inputs(100));
    layer0_outputs(581) <= not(inputs(104)) or (inputs(176));
    layer0_outputs(582) <= not((inputs(65)) or (inputs(87)));
    layer0_outputs(583) <= not(inputs(21));
    layer0_outputs(584) <= inputs(113);
    layer0_outputs(585) <= (inputs(247)) xor (inputs(58));
    layer0_outputs(586) <= not((inputs(0)) or (inputs(215)));
    layer0_outputs(587) <= (inputs(15)) and not (inputs(137));
    layer0_outputs(588) <= not((inputs(171)) and (inputs(195)));
    layer0_outputs(589) <= (inputs(44)) or (inputs(6));
    layer0_outputs(590) <= inputs(16);
    layer0_outputs(591) <= not(inputs(74)) or (inputs(236));
    layer0_outputs(592) <= (inputs(59)) and not (inputs(71));
    layer0_outputs(593) <= not(inputs(247));
    layer0_outputs(594) <= inputs(53);
    layer0_outputs(595) <= inputs(6);
    layer0_outputs(596) <= inputs(168);
    layer0_outputs(597) <= not(inputs(78));
    layer0_outputs(598) <= not((inputs(249)) or (inputs(18)));
    layer0_outputs(599) <= inputs(145);
    layer0_outputs(600) <= (inputs(140)) and not (inputs(50));
    layer0_outputs(601) <= (inputs(230)) and not (inputs(75));
    layer0_outputs(602) <= not(inputs(118));
    layer0_outputs(603) <= inputs(163);
    layer0_outputs(604) <= not(inputs(218));
    layer0_outputs(605) <= inputs(31);
    layer0_outputs(606) <= inputs(161);
    layer0_outputs(607) <= inputs(139);
    layer0_outputs(608) <= (inputs(128)) and not (inputs(143));
    layer0_outputs(609) <= (inputs(243)) xor (inputs(216));
    layer0_outputs(610) <= not(inputs(25));
    layer0_outputs(611) <= not((inputs(72)) xor (inputs(108)));
    layer0_outputs(612) <= not(inputs(131));
    layer0_outputs(613) <= inputs(114);
    layer0_outputs(614) <= not((inputs(129)) xor (inputs(116)));
    layer0_outputs(615) <= not(inputs(87));
    layer0_outputs(616) <= (inputs(76)) or (inputs(192));
    layer0_outputs(617) <= inputs(108);
    layer0_outputs(618) <= (inputs(191)) xor (inputs(165));
    layer0_outputs(619) <= (inputs(169)) or (inputs(18));
    layer0_outputs(620) <= not(inputs(195));
    layer0_outputs(621) <= not(inputs(88));
    layer0_outputs(622) <= inputs(165);
    layer0_outputs(623) <= (inputs(96)) or (inputs(95));
    layer0_outputs(624) <= not(inputs(105));
    layer0_outputs(625) <= inputs(184);
    layer0_outputs(626) <= (inputs(113)) or (inputs(111));
    layer0_outputs(627) <= not((inputs(37)) or (inputs(52)));
    layer0_outputs(628) <= (inputs(186)) and not (inputs(97));
    layer0_outputs(629) <= inputs(128);
    layer0_outputs(630) <= not((inputs(51)) or (inputs(108)));
    layer0_outputs(631) <= inputs(56);
    layer0_outputs(632) <= not((inputs(126)) xor (inputs(199)));
    layer0_outputs(633) <= (inputs(152)) and not (inputs(211));
    layer0_outputs(634) <= not(inputs(61));
    layer0_outputs(635) <= (inputs(166)) and not (inputs(81));
    layer0_outputs(636) <= not(inputs(86));
    layer0_outputs(637) <= (inputs(87)) xor (inputs(43));
    layer0_outputs(638) <= (inputs(140)) xor (inputs(204));
    layer0_outputs(639) <= not((inputs(203)) xor (inputs(104)));
    layer0_outputs(640) <= not(inputs(103)) or (inputs(125));
    layer0_outputs(641) <= (inputs(205)) and (inputs(185));
    layer0_outputs(642) <= (inputs(210)) xor (inputs(92));
    layer0_outputs(643) <= (inputs(73)) or (inputs(140));
    layer0_outputs(644) <= not(inputs(146));
    layer0_outputs(645) <= not((inputs(64)) or (inputs(232)));
    layer0_outputs(646) <= not(inputs(218));
    layer0_outputs(647) <= inputs(98);
    layer0_outputs(648) <= not((inputs(28)) or (inputs(238)));
    layer0_outputs(649) <= not((inputs(57)) or (inputs(241)));
    layer0_outputs(650) <= '0';
    layer0_outputs(651) <= inputs(6);
    layer0_outputs(652) <= not((inputs(222)) xor (inputs(60)));
    layer0_outputs(653) <= not(inputs(91));
    layer0_outputs(654) <= not((inputs(0)) or (inputs(40)));
    layer0_outputs(655) <= (inputs(170)) xor (inputs(191));
    layer0_outputs(656) <= not(inputs(214)) or (inputs(131));
    layer0_outputs(657) <= not((inputs(33)) or (inputs(187)));
    layer0_outputs(658) <= not((inputs(172)) or (inputs(222)));
    layer0_outputs(659) <= not((inputs(244)) xor (inputs(36)));
    layer0_outputs(660) <= not(inputs(207)) or (inputs(81));
    layer0_outputs(661) <= (inputs(38)) or (inputs(255));
    layer0_outputs(662) <= (inputs(61)) or (inputs(58));
    layer0_outputs(663) <= not(inputs(180));
    layer0_outputs(664) <= not(inputs(146));
    layer0_outputs(665) <= inputs(162);
    layer0_outputs(666) <= not((inputs(177)) xor (inputs(220)));
    layer0_outputs(667) <= inputs(124);
    layer0_outputs(668) <= inputs(164);
    layer0_outputs(669) <= '1';
    layer0_outputs(670) <= (inputs(17)) xor (inputs(135));
    layer0_outputs(671) <= (inputs(19)) xor (inputs(253));
    layer0_outputs(672) <= (inputs(199)) or (inputs(184));
    layer0_outputs(673) <= not((inputs(28)) or (inputs(95)));
    layer0_outputs(674) <= (inputs(210)) or (inputs(247));
    layer0_outputs(675) <= (inputs(126)) and not (inputs(246));
    layer0_outputs(676) <= inputs(51);
    layer0_outputs(677) <= not(inputs(151));
    layer0_outputs(678) <= (inputs(254)) xor (inputs(99));
    layer0_outputs(679) <= not(inputs(73));
    layer0_outputs(680) <= (inputs(75)) and not (inputs(163));
    layer0_outputs(681) <= (inputs(106)) and not (inputs(229));
    layer0_outputs(682) <= not(inputs(18));
    layer0_outputs(683) <= not((inputs(141)) or (inputs(157)));
    layer0_outputs(684) <= not((inputs(150)) xor (inputs(80)));
    layer0_outputs(685) <= inputs(228);
    layer0_outputs(686) <= inputs(22);
    layer0_outputs(687) <= (inputs(9)) or (inputs(116));
    layer0_outputs(688) <= (inputs(111)) or (inputs(97));
    layer0_outputs(689) <= (inputs(233)) and not (inputs(64));
    layer0_outputs(690) <= inputs(128);
    layer0_outputs(691) <= (inputs(183)) and not (inputs(42));
    layer0_outputs(692) <= (inputs(112)) xor (inputs(170));
    layer0_outputs(693) <= (inputs(52)) xor (inputs(54));
    layer0_outputs(694) <= inputs(189);
    layer0_outputs(695) <= not(inputs(219));
    layer0_outputs(696) <= '0';
    layer0_outputs(697) <= not((inputs(97)) xor (inputs(159)));
    layer0_outputs(698) <= (inputs(112)) and not (inputs(32));
    layer0_outputs(699) <= (inputs(134)) and (inputs(94));
    layer0_outputs(700) <= (inputs(104)) xor (inputs(3));
    layer0_outputs(701) <= (inputs(144)) xor (inputs(168));
    layer0_outputs(702) <= (inputs(158)) or (inputs(73));
    layer0_outputs(703) <= (inputs(64)) and not (inputs(59));
    layer0_outputs(704) <= inputs(133);
    layer0_outputs(705) <= inputs(106);
    layer0_outputs(706) <= (inputs(93)) xor (inputs(153));
    layer0_outputs(707) <= (inputs(38)) or (inputs(54));
    layer0_outputs(708) <= (inputs(0)) or (inputs(63));
    layer0_outputs(709) <= not((inputs(41)) xor (inputs(160)));
    layer0_outputs(710) <= not((inputs(217)) xor (inputs(41)));
    layer0_outputs(711) <= (inputs(134)) and not (inputs(72));
    layer0_outputs(712) <= (inputs(120)) and not (inputs(219));
    layer0_outputs(713) <= not((inputs(242)) or (inputs(103)));
    layer0_outputs(714) <= (inputs(139)) and (inputs(75));
    layer0_outputs(715) <= not(inputs(84)) or (inputs(157));
    layer0_outputs(716) <= inputs(44);
    layer0_outputs(717) <= (inputs(127)) or (inputs(66));
    layer0_outputs(718) <= not((inputs(110)) or (inputs(145)));
    layer0_outputs(719) <= not((inputs(156)) or (inputs(1)));
    layer0_outputs(720) <= (inputs(226)) and not (inputs(131));
    layer0_outputs(721) <= (inputs(145)) or (inputs(48));
    layer0_outputs(722) <= (inputs(237)) xor (inputs(52));
    layer0_outputs(723) <= (inputs(65)) and (inputs(179));
    layer0_outputs(724) <= (inputs(25)) xor (inputs(110));
    layer0_outputs(725) <= (inputs(45)) xor (inputs(81));
    layer0_outputs(726) <= not((inputs(191)) or (inputs(36)));
    layer0_outputs(727) <= (inputs(3)) or (inputs(212));
    layer0_outputs(728) <= not(inputs(64));
    layer0_outputs(729) <= (inputs(230)) or (inputs(4));
    layer0_outputs(730) <= not((inputs(4)) xor (inputs(102)));
    layer0_outputs(731) <= not((inputs(229)) or (inputs(175)));
    layer0_outputs(732) <= not((inputs(253)) and (inputs(236)));
    layer0_outputs(733) <= (inputs(49)) or (inputs(124));
    layer0_outputs(734) <= (inputs(63)) or (inputs(8));
    layer0_outputs(735) <= inputs(164);
    layer0_outputs(736) <= not((inputs(66)) or (inputs(67)));
    layer0_outputs(737) <= (inputs(207)) and not (inputs(241));
    layer0_outputs(738) <= not((inputs(197)) xor (inputs(14)));
    layer0_outputs(739) <= not(inputs(252)) or (inputs(197));
    layer0_outputs(740) <= not((inputs(165)) and (inputs(151)));
    layer0_outputs(741) <= not((inputs(85)) or (inputs(35)));
    layer0_outputs(742) <= not(inputs(226)) or (inputs(141));
    layer0_outputs(743) <= not((inputs(183)) xor (inputs(149)));
    layer0_outputs(744) <= (inputs(222)) and not (inputs(155));
    layer0_outputs(745) <= (inputs(57)) or (inputs(120));
    layer0_outputs(746) <= not((inputs(240)) and (inputs(147)));
    layer0_outputs(747) <= not((inputs(106)) and (inputs(10)));
    layer0_outputs(748) <= not(inputs(85));
    layer0_outputs(749) <= not(inputs(104));
    layer0_outputs(750) <= (inputs(183)) and not (inputs(144));
    layer0_outputs(751) <= inputs(166);
    layer0_outputs(752) <= not((inputs(200)) and (inputs(228)));
    layer0_outputs(753) <= (inputs(178)) or (inputs(146));
    layer0_outputs(754) <= (inputs(192)) and not (inputs(241));
    layer0_outputs(755) <= not((inputs(188)) or (inputs(34)));
    layer0_outputs(756) <= (inputs(221)) and (inputs(202));
    layer0_outputs(757) <= (inputs(146)) xor (inputs(215));
    layer0_outputs(758) <= not((inputs(8)) xor (inputs(217)));
    layer0_outputs(759) <= '1';
    layer0_outputs(760) <= inputs(226);
    layer0_outputs(761) <= (inputs(71)) xor (inputs(83));
    layer0_outputs(762) <= (inputs(159)) or (inputs(126));
    layer0_outputs(763) <= (inputs(127)) or (inputs(148));
    layer0_outputs(764) <= not((inputs(57)) or (inputs(49)));
    layer0_outputs(765) <= inputs(198);
    layer0_outputs(766) <= not(inputs(67)) or (inputs(221));
    layer0_outputs(767) <= not((inputs(92)) or (inputs(49)));
    layer0_outputs(768) <= inputs(78);
    layer0_outputs(769) <= not((inputs(39)) and (inputs(115)));
    layer0_outputs(770) <= (inputs(243)) xor (inputs(13));
    layer0_outputs(771) <= not(inputs(120));
    layer0_outputs(772) <= (inputs(146)) or (inputs(162));
    layer0_outputs(773) <= (inputs(246)) and not (inputs(161));
    layer0_outputs(774) <= (inputs(68)) and not (inputs(247));
    layer0_outputs(775) <= (inputs(213)) and not (inputs(164));
    layer0_outputs(776) <= not((inputs(199)) or (inputs(104)));
    layer0_outputs(777) <= (inputs(222)) or (inputs(36));
    layer0_outputs(778) <= not(inputs(81));
    layer0_outputs(779) <= inputs(173);
    layer0_outputs(780) <= not(inputs(98));
    layer0_outputs(781) <= (inputs(104)) xor (inputs(42));
    layer0_outputs(782) <= not(inputs(150));
    layer0_outputs(783) <= not((inputs(170)) xor (inputs(233)));
    layer0_outputs(784) <= not(inputs(39)) or (inputs(124));
    layer0_outputs(785) <= not(inputs(177));
    layer0_outputs(786) <= inputs(225);
    layer0_outputs(787) <= (inputs(66)) or (inputs(43));
    layer0_outputs(788) <= (inputs(125)) or (inputs(3));
    layer0_outputs(789) <= not((inputs(162)) or (inputs(251)));
    layer0_outputs(790) <= inputs(26);
    layer0_outputs(791) <= (inputs(193)) or (inputs(68));
    layer0_outputs(792) <= '0';
    layer0_outputs(793) <= not((inputs(134)) xor (inputs(167)));
    layer0_outputs(794) <= (inputs(117)) xor (inputs(129));
    layer0_outputs(795) <= not(inputs(99));
    layer0_outputs(796) <= not((inputs(53)) or (inputs(47)));
    layer0_outputs(797) <= (inputs(98)) and not (inputs(250));
    layer0_outputs(798) <= not(inputs(83));
    layer0_outputs(799) <= inputs(203);
    layer0_outputs(800) <= not(inputs(173)) or (inputs(128));
    layer0_outputs(801) <= not(inputs(202));
    layer0_outputs(802) <= (inputs(135)) or (inputs(245));
    layer0_outputs(803) <= not(inputs(200)) or (inputs(228));
    layer0_outputs(804) <= not(inputs(21));
    layer0_outputs(805) <= not(inputs(11));
    layer0_outputs(806) <= (inputs(242)) xor (inputs(74));
    layer0_outputs(807) <= inputs(184);
    layer0_outputs(808) <= (inputs(140)) xor (inputs(170));
    layer0_outputs(809) <= (inputs(88)) xor (inputs(93));
    layer0_outputs(810) <= inputs(195);
    layer0_outputs(811) <= inputs(179);
    layer0_outputs(812) <= (inputs(191)) and (inputs(151));
    layer0_outputs(813) <= not(inputs(108));
    layer0_outputs(814) <= not((inputs(148)) and (inputs(159)));
    layer0_outputs(815) <= inputs(157);
    layer0_outputs(816) <= (inputs(140)) xor (inputs(27));
    layer0_outputs(817) <= (inputs(154)) and not (inputs(167));
    layer0_outputs(818) <= inputs(200);
    layer0_outputs(819) <= (inputs(136)) and not (inputs(4));
    layer0_outputs(820) <= inputs(128);
    layer0_outputs(821) <= not(inputs(212)) or (inputs(83));
    layer0_outputs(822) <= not(inputs(71));
    layer0_outputs(823) <= not(inputs(56));
    layer0_outputs(824) <= inputs(61);
    layer0_outputs(825) <= (inputs(5)) or (inputs(241));
    layer0_outputs(826) <= (inputs(50)) or (inputs(76));
    layer0_outputs(827) <= not((inputs(75)) or (inputs(10)));
    layer0_outputs(828) <= not(inputs(136));
    layer0_outputs(829) <= (inputs(49)) and not (inputs(46));
    layer0_outputs(830) <= inputs(88);
    layer0_outputs(831) <= not((inputs(241)) xor (inputs(1)));
    layer0_outputs(832) <= (inputs(108)) and not (inputs(83));
    layer0_outputs(833) <= (inputs(61)) or (inputs(98));
    layer0_outputs(834) <= not((inputs(220)) or (inputs(174)));
    layer0_outputs(835) <= not(inputs(33)) or (inputs(127));
    layer0_outputs(836) <= not((inputs(206)) xor (inputs(110)));
    layer0_outputs(837) <= (inputs(233)) or (inputs(202));
    layer0_outputs(838) <= (inputs(14)) or (inputs(100));
    layer0_outputs(839) <= not((inputs(6)) or (inputs(33)));
    layer0_outputs(840) <= inputs(169);
    layer0_outputs(841) <= '1';
    layer0_outputs(842) <= inputs(148);
    layer0_outputs(843) <= not(inputs(8));
    layer0_outputs(844) <= not((inputs(110)) or (inputs(75)));
    layer0_outputs(845) <= (inputs(74)) and not (inputs(35));
    layer0_outputs(846) <= inputs(133);
    layer0_outputs(847) <= (inputs(126)) or (inputs(12));
    layer0_outputs(848) <= (inputs(79)) xor (inputs(21));
    layer0_outputs(849) <= inputs(134);
    layer0_outputs(850) <= (inputs(73)) and not (inputs(193));
    layer0_outputs(851) <= not(inputs(233)) or (inputs(253));
    layer0_outputs(852) <= not(inputs(20));
    layer0_outputs(853) <= not(inputs(113)) or (inputs(55));
    layer0_outputs(854) <= not((inputs(46)) xor (inputs(133)));
    layer0_outputs(855) <= not((inputs(238)) or (inputs(40)));
    layer0_outputs(856) <= not(inputs(142)) or (inputs(121));
    layer0_outputs(857) <= not(inputs(244)) or (inputs(103));
    layer0_outputs(858) <= not(inputs(99)) or (inputs(15));
    layer0_outputs(859) <= not(inputs(108)) or (inputs(207));
    layer0_outputs(860) <= not((inputs(251)) or (inputs(159)));
    layer0_outputs(861) <= inputs(68);
    layer0_outputs(862) <= inputs(195);
    layer0_outputs(863) <= (inputs(208)) or (inputs(217));
    layer0_outputs(864) <= not(inputs(190));
    layer0_outputs(865) <= (inputs(252)) or (inputs(230));
    layer0_outputs(866) <= not(inputs(203)) or (inputs(118));
    layer0_outputs(867) <= not((inputs(41)) and (inputs(44)));
    layer0_outputs(868) <= inputs(201);
    layer0_outputs(869) <= (inputs(9)) and not (inputs(65));
    layer0_outputs(870) <= not((inputs(251)) or (inputs(133)));
    layer0_outputs(871) <= (inputs(153)) or (inputs(17));
    layer0_outputs(872) <= not(inputs(117)) or (inputs(62));
    layer0_outputs(873) <= inputs(89);
    layer0_outputs(874) <= not((inputs(38)) or (inputs(193)));
    layer0_outputs(875) <= not(inputs(123));
    layer0_outputs(876) <= not(inputs(244));
    layer0_outputs(877) <= (inputs(81)) or (inputs(103));
    layer0_outputs(878) <= not((inputs(67)) xor (inputs(84)));
    layer0_outputs(879) <= not(inputs(143));
    layer0_outputs(880) <= not((inputs(245)) xor (inputs(214)));
    layer0_outputs(881) <= inputs(236);
    layer0_outputs(882) <= (inputs(218)) xor (inputs(209));
    layer0_outputs(883) <= not(inputs(122));
    layer0_outputs(884) <= not(inputs(98));
    layer0_outputs(885) <= inputs(196);
    layer0_outputs(886) <= '1';
    layer0_outputs(887) <= (inputs(104)) and not (inputs(152));
    layer0_outputs(888) <= inputs(162);
    layer0_outputs(889) <= (inputs(87)) and not (inputs(16));
    layer0_outputs(890) <= not((inputs(15)) xor (inputs(150)));
    layer0_outputs(891) <= not(inputs(43));
    layer0_outputs(892) <= not((inputs(44)) and (inputs(12)));
    layer0_outputs(893) <= not(inputs(242));
    layer0_outputs(894) <= (inputs(28)) and (inputs(9));
    layer0_outputs(895) <= inputs(159);
    layer0_outputs(896) <= not(inputs(118)) or (inputs(160));
    layer0_outputs(897) <= not((inputs(134)) xor (inputs(163)));
    layer0_outputs(898) <= not((inputs(203)) and (inputs(224)));
    layer0_outputs(899) <= not((inputs(143)) xor (inputs(233)));
    layer0_outputs(900) <= inputs(67);
    layer0_outputs(901) <= not(inputs(116));
    layer0_outputs(902) <= inputs(56);
    layer0_outputs(903) <= (inputs(180)) or (inputs(209));
    layer0_outputs(904) <= not(inputs(203));
    layer0_outputs(905) <= (inputs(23)) xor (inputs(211));
    layer0_outputs(906) <= inputs(112);
    layer0_outputs(907) <= (inputs(149)) and not (inputs(20));
    layer0_outputs(908) <= (inputs(45)) or (inputs(244));
    layer0_outputs(909) <= (inputs(163)) and (inputs(227));
    layer0_outputs(910) <= inputs(14);
    layer0_outputs(911) <= (inputs(223)) or (inputs(212));
    layer0_outputs(912) <= not((inputs(116)) xor (inputs(122)));
    layer0_outputs(913) <= not((inputs(183)) or (inputs(62)));
    layer0_outputs(914) <= not(inputs(132));
    layer0_outputs(915) <= not(inputs(20)) or (inputs(69));
    layer0_outputs(916) <= inputs(228);
    layer0_outputs(917) <= (inputs(60)) and not (inputs(214));
    layer0_outputs(918) <= (inputs(150)) and not (inputs(113));
    layer0_outputs(919) <= not(inputs(133));
    layer0_outputs(920) <= not((inputs(201)) or (inputs(190)));
    layer0_outputs(921) <= not(inputs(51)) or (inputs(110));
    layer0_outputs(922) <= not(inputs(218));
    layer0_outputs(923) <= (inputs(5)) or (inputs(206));
    layer0_outputs(924) <= '0';
    layer0_outputs(925) <= (inputs(89)) and not (inputs(31));
    layer0_outputs(926) <= not(inputs(131));
    layer0_outputs(927) <= not(inputs(184));
    layer0_outputs(928) <= not((inputs(5)) xor (inputs(169)));
    layer0_outputs(929) <= inputs(197);
    layer0_outputs(930) <= not((inputs(109)) xor (inputs(156)));
    layer0_outputs(931) <= (inputs(163)) xor (inputs(125));
    layer0_outputs(932) <= (inputs(27)) xor (inputs(145));
    layer0_outputs(933) <= not(inputs(166)) or (inputs(225));
    layer0_outputs(934) <= (inputs(7)) or (inputs(22));
    layer0_outputs(935) <= (inputs(120)) and (inputs(113));
    layer0_outputs(936) <= not((inputs(115)) or (inputs(162)));
    layer0_outputs(937) <= not((inputs(76)) and (inputs(107)));
    layer0_outputs(938) <= '0';
    layer0_outputs(939) <= not(inputs(147));
    layer0_outputs(940) <= inputs(145);
    layer0_outputs(941) <= not((inputs(86)) or (inputs(100)));
    layer0_outputs(942) <= '1';
    layer0_outputs(943) <= not((inputs(142)) or (inputs(207)));
    layer0_outputs(944) <= not((inputs(221)) or (inputs(17)));
    layer0_outputs(945) <= not((inputs(64)) or (inputs(66)));
    layer0_outputs(946) <= (inputs(92)) and not (inputs(67));
    layer0_outputs(947) <= (inputs(92)) xor (inputs(1));
    layer0_outputs(948) <= not(inputs(19));
    layer0_outputs(949) <= (inputs(16)) or (inputs(85));
    layer0_outputs(950) <= inputs(133);
    layer0_outputs(951) <= not(inputs(81)) or (inputs(156));
    layer0_outputs(952) <= (inputs(151)) xor (inputs(194));
    layer0_outputs(953) <= (inputs(150)) xor (inputs(103));
    layer0_outputs(954) <= not((inputs(224)) or (inputs(77)));
    layer0_outputs(955) <= not(inputs(232));
    layer0_outputs(956) <= not(inputs(223)) or (inputs(226));
    layer0_outputs(957) <= inputs(111);
    layer0_outputs(958) <= inputs(52);
    layer0_outputs(959) <= not((inputs(143)) or (inputs(67)));
    layer0_outputs(960) <= (inputs(93)) and not (inputs(240));
    layer0_outputs(961) <= (inputs(235)) and not (inputs(132));
    layer0_outputs(962) <= (inputs(131)) and not (inputs(203));
    layer0_outputs(963) <= not((inputs(42)) or (inputs(124)));
    layer0_outputs(964) <= not((inputs(150)) or (inputs(176)));
    layer0_outputs(965) <= (inputs(210)) or (inputs(240));
    layer0_outputs(966) <= inputs(230);
    layer0_outputs(967) <= (inputs(25)) or (inputs(65));
    layer0_outputs(968) <= (inputs(119)) and not (inputs(170));
    layer0_outputs(969) <= (inputs(228)) or (inputs(191));
    layer0_outputs(970) <= (inputs(249)) and not (inputs(239));
    layer0_outputs(971) <= (inputs(135)) or (inputs(65));
    layer0_outputs(972) <= inputs(49);
    layer0_outputs(973) <= not(inputs(21));
    layer0_outputs(974) <= (inputs(43)) xor (inputs(181));
    layer0_outputs(975) <= (inputs(77)) or (inputs(93));
    layer0_outputs(976) <= '1';
    layer0_outputs(977) <= (inputs(97)) and not (inputs(224));
    layer0_outputs(978) <= inputs(162);
    layer0_outputs(979) <= inputs(253);
    layer0_outputs(980) <= (inputs(71)) xor (inputs(83));
    layer0_outputs(981) <= inputs(39);
    layer0_outputs(982) <= not(inputs(169));
    layer0_outputs(983) <= inputs(144);
    layer0_outputs(984) <= inputs(38);
    layer0_outputs(985) <= not(inputs(109)) or (inputs(9));
    layer0_outputs(986) <= inputs(130);
    layer0_outputs(987) <= not(inputs(214));
    layer0_outputs(988) <= '0';
    layer0_outputs(989) <= not(inputs(251));
    layer0_outputs(990) <= inputs(163);
    layer0_outputs(991) <= not(inputs(248));
    layer0_outputs(992) <= (inputs(117)) xor (inputs(234));
    layer0_outputs(993) <= (inputs(18)) xor (inputs(9));
    layer0_outputs(994) <= '0';
    layer0_outputs(995) <= not((inputs(0)) and (inputs(184)));
    layer0_outputs(996) <= inputs(23);
    layer0_outputs(997) <= not(inputs(247)) or (inputs(7));
    layer0_outputs(998) <= not(inputs(212));
    layer0_outputs(999) <= not((inputs(196)) or (inputs(176)));
    layer0_outputs(1000) <= not(inputs(138)) or (inputs(236));
    layer0_outputs(1001) <= not(inputs(107));
    layer0_outputs(1002) <= (inputs(217)) and not (inputs(65));
    layer0_outputs(1003) <= inputs(68);
    layer0_outputs(1004) <= (inputs(217)) and not (inputs(237));
    layer0_outputs(1005) <= inputs(211);
    layer0_outputs(1006) <= inputs(209);
    layer0_outputs(1007) <= not((inputs(250)) or (inputs(109)));
    layer0_outputs(1008) <= not((inputs(105)) or (inputs(106)));
    layer0_outputs(1009) <= not((inputs(33)) and (inputs(227)));
    layer0_outputs(1010) <= (inputs(107)) xor (inputs(197));
    layer0_outputs(1011) <= not(inputs(83));
    layer0_outputs(1012) <= not(inputs(38));
    layer0_outputs(1013) <= inputs(216);
    layer0_outputs(1014) <= (inputs(52)) or (inputs(28));
    layer0_outputs(1015) <= (inputs(193)) and not (inputs(50));
    layer0_outputs(1016) <= (inputs(156)) and (inputs(59));
    layer0_outputs(1017) <= not(inputs(51));
    layer0_outputs(1018) <= (inputs(109)) and not (inputs(207));
    layer0_outputs(1019) <= (inputs(99)) xor (inputs(73));
    layer0_outputs(1020) <= not(inputs(111));
    layer0_outputs(1021) <= not((inputs(77)) or (inputs(35)));
    layer0_outputs(1022) <= inputs(89);
    layer0_outputs(1023) <= inputs(82);
    layer0_outputs(1024) <= not((inputs(238)) or (inputs(50)));
    layer0_outputs(1025) <= '0';
    layer0_outputs(1026) <= inputs(101);
    layer0_outputs(1027) <= not((inputs(204)) or (inputs(240)));
    layer0_outputs(1028) <= '1';
    layer0_outputs(1029) <= (inputs(152)) and not (inputs(28));
    layer0_outputs(1030) <= (inputs(80)) xor (inputs(167));
    layer0_outputs(1031) <= inputs(232);
    layer0_outputs(1032) <= not((inputs(195)) or (inputs(245)));
    layer0_outputs(1033) <= not(inputs(113));
    layer0_outputs(1034) <= not(inputs(126));
    layer0_outputs(1035) <= not((inputs(11)) or (inputs(31)));
    layer0_outputs(1036) <= inputs(90);
    layer0_outputs(1037) <= inputs(147);
    layer0_outputs(1038) <= (inputs(240)) or (inputs(24));
    layer0_outputs(1039) <= (inputs(10)) and not (inputs(88));
    layer0_outputs(1040) <= (inputs(60)) or (inputs(195));
    layer0_outputs(1041) <= (inputs(39)) or (inputs(35));
    layer0_outputs(1042) <= not(inputs(167));
    layer0_outputs(1043) <= '1';
    layer0_outputs(1044) <= not((inputs(174)) or (inputs(176)));
    layer0_outputs(1045) <= not(inputs(75));
    layer0_outputs(1046) <= not(inputs(252));
    layer0_outputs(1047) <= (inputs(129)) or (inputs(59));
    layer0_outputs(1048) <= not(inputs(227));
    layer0_outputs(1049) <= (inputs(61)) and (inputs(11));
    layer0_outputs(1050) <= inputs(163);
    layer0_outputs(1051) <= not((inputs(65)) or (inputs(47)));
    layer0_outputs(1052) <= inputs(66);
    layer0_outputs(1053) <= (inputs(89)) xor (inputs(232));
    layer0_outputs(1054) <= (inputs(13)) and not (inputs(191));
    layer0_outputs(1055) <= not((inputs(225)) xor (inputs(26)));
    layer0_outputs(1056) <= not(inputs(191));
    layer0_outputs(1057) <= not((inputs(89)) xor (inputs(134)));
    layer0_outputs(1058) <= '1';
    layer0_outputs(1059) <= not((inputs(127)) or (inputs(182)));
    layer0_outputs(1060) <= not((inputs(47)) or (inputs(23)));
    layer0_outputs(1061) <= not(inputs(95));
    layer0_outputs(1062) <= not(inputs(214));
    layer0_outputs(1063) <= (inputs(162)) or (inputs(190));
    layer0_outputs(1064) <= inputs(2);
    layer0_outputs(1065) <= (inputs(183)) xor (inputs(109));
    layer0_outputs(1066) <= (inputs(252)) or (inputs(54));
    layer0_outputs(1067) <= inputs(251);
    layer0_outputs(1068) <= not(inputs(121)) or (inputs(129));
    layer0_outputs(1069) <= inputs(190);
    layer0_outputs(1070) <= not((inputs(118)) or (inputs(248)));
    layer0_outputs(1071) <= (inputs(184)) and (inputs(241));
    layer0_outputs(1072) <= inputs(234);
    layer0_outputs(1073) <= not(inputs(37)) or (inputs(234));
    layer0_outputs(1074) <= (inputs(111)) or (inputs(1));
    layer0_outputs(1075) <= (inputs(254)) or (inputs(146));
    layer0_outputs(1076) <= (inputs(179)) or (inputs(49));
    layer0_outputs(1077) <= not(inputs(231));
    layer0_outputs(1078) <= (inputs(86)) or (inputs(109));
    layer0_outputs(1079) <= (inputs(219)) or (inputs(2));
    layer0_outputs(1080) <= not(inputs(44));
    layer0_outputs(1081) <= not(inputs(120));
    layer0_outputs(1082) <= (inputs(179)) and not (inputs(78));
    layer0_outputs(1083) <= not((inputs(35)) or (inputs(247)));
    layer0_outputs(1084) <= inputs(16);
    layer0_outputs(1085) <= not(inputs(206)) or (inputs(48));
    layer0_outputs(1086) <= not(inputs(106)) or (inputs(235));
    layer0_outputs(1087) <= not(inputs(107));
    layer0_outputs(1088) <= not(inputs(50)) or (inputs(61));
    layer0_outputs(1089) <= (inputs(173)) and not (inputs(247));
    layer0_outputs(1090) <= not(inputs(74));
    layer0_outputs(1091) <= (inputs(27)) or (inputs(57));
    layer0_outputs(1092) <= not((inputs(51)) and (inputs(7)));
    layer0_outputs(1093) <= not((inputs(173)) xor (inputs(83)));
    layer0_outputs(1094) <= not(inputs(174));
    layer0_outputs(1095) <= (inputs(53)) or (inputs(9));
    layer0_outputs(1096) <= not((inputs(152)) xor (inputs(165)));
    layer0_outputs(1097) <= not(inputs(167));
    layer0_outputs(1098) <= not(inputs(229));
    layer0_outputs(1099) <= not(inputs(203)) or (inputs(32));
    layer0_outputs(1100) <= inputs(79);
    layer0_outputs(1101) <= inputs(114);
    layer0_outputs(1102) <= (inputs(85)) xor (inputs(113));
    layer0_outputs(1103) <= (inputs(123)) xor (inputs(57));
    layer0_outputs(1104) <= (inputs(56)) and not (inputs(205));
    layer0_outputs(1105) <= (inputs(82)) and not (inputs(152));
    layer0_outputs(1106) <= (inputs(190)) xor (inputs(125));
    layer0_outputs(1107) <= (inputs(146)) xor (inputs(194));
    layer0_outputs(1108) <= not((inputs(79)) or (inputs(164)));
    layer0_outputs(1109) <= (inputs(84)) and not (inputs(160));
    layer0_outputs(1110) <= (inputs(184)) and not (inputs(205));
    layer0_outputs(1111) <= '1';
    layer0_outputs(1112) <= '1';
    layer0_outputs(1113) <= inputs(129);
    layer0_outputs(1114) <= not((inputs(255)) or (inputs(185)));
    layer0_outputs(1115) <= inputs(92);
    layer0_outputs(1116) <= not(inputs(139)) or (inputs(248));
    layer0_outputs(1117) <= not(inputs(120));
    layer0_outputs(1118) <= (inputs(77)) and not (inputs(99));
    layer0_outputs(1119) <= inputs(107);
    layer0_outputs(1120) <= inputs(212);
    layer0_outputs(1121) <= not((inputs(139)) xor (inputs(254)));
    layer0_outputs(1122) <= not(inputs(139));
    layer0_outputs(1123) <= not((inputs(116)) xor (inputs(144)));
    layer0_outputs(1124) <= not(inputs(119)) or (inputs(141));
    layer0_outputs(1125) <= not(inputs(232)) or (inputs(1));
    layer0_outputs(1126) <= not((inputs(201)) xor (inputs(249)));
    layer0_outputs(1127) <= inputs(224);
    layer0_outputs(1128) <= not(inputs(135)) or (inputs(143));
    layer0_outputs(1129) <= (inputs(82)) xor (inputs(36));
    layer0_outputs(1130) <= (inputs(168)) xor (inputs(119));
    layer0_outputs(1131) <= inputs(191);
    layer0_outputs(1132) <= (inputs(63)) or (inputs(119));
    layer0_outputs(1133) <= not((inputs(162)) or (inputs(126)));
    layer0_outputs(1134) <= (inputs(166)) xor (inputs(0));
    layer0_outputs(1135) <= (inputs(245)) xor (inputs(38));
    layer0_outputs(1136) <= (inputs(157)) xor (inputs(21));
    layer0_outputs(1137) <= not(inputs(217));
    layer0_outputs(1138) <= (inputs(42)) and not (inputs(120));
    layer0_outputs(1139) <= inputs(63);
    layer0_outputs(1140) <= (inputs(251)) and not (inputs(160));
    layer0_outputs(1141) <= not((inputs(4)) or (inputs(195)));
    layer0_outputs(1142) <= inputs(19);
    layer0_outputs(1143) <= inputs(238);
    layer0_outputs(1144) <= (inputs(249)) or (inputs(172));
    layer0_outputs(1145) <= not(inputs(194));
    layer0_outputs(1146) <= not((inputs(232)) xor (inputs(22)));
    layer0_outputs(1147) <= not((inputs(230)) or (inputs(206)));
    layer0_outputs(1148) <= not(inputs(220)) or (inputs(240));
    layer0_outputs(1149) <= not(inputs(75)) or (inputs(102));
    layer0_outputs(1150) <= inputs(126);
    layer0_outputs(1151) <= not((inputs(210)) or (inputs(25)));
    layer0_outputs(1152) <= (inputs(116)) xor (inputs(169));
    layer0_outputs(1153) <= inputs(209);
    layer0_outputs(1154) <= not((inputs(144)) or (inputs(32)));
    layer0_outputs(1155) <= inputs(79);
    layer0_outputs(1156) <= not(inputs(158)) or (inputs(87));
    layer0_outputs(1157) <= not((inputs(192)) or (inputs(77)));
    layer0_outputs(1158) <= not(inputs(30)) or (inputs(242));
    layer0_outputs(1159) <= (inputs(136)) and not (inputs(143));
    layer0_outputs(1160) <= not((inputs(14)) xor (inputs(13)));
    layer0_outputs(1161) <= (inputs(186)) and not (inputs(69));
    layer0_outputs(1162) <= inputs(194);
    layer0_outputs(1163) <= (inputs(28)) xor (inputs(37));
    layer0_outputs(1164) <= not((inputs(238)) or (inputs(5)));
    layer0_outputs(1165) <= not((inputs(154)) or (inputs(88)));
    layer0_outputs(1166) <= not(inputs(149));
    layer0_outputs(1167) <= (inputs(167)) and not (inputs(31));
    layer0_outputs(1168) <= not((inputs(161)) xor (inputs(249)));
    layer0_outputs(1169) <= not(inputs(4));
    layer0_outputs(1170) <= not((inputs(209)) or (inputs(114)));
    layer0_outputs(1171) <= (inputs(146)) and not (inputs(149));
    layer0_outputs(1172) <= (inputs(247)) xor (inputs(220));
    layer0_outputs(1173) <= not((inputs(230)) xor (inputs(162)));
    layer0_outputs(1174) <= not((inputs(228)) and (inputs(210)));
    layer0_outputs(1175) <= not(inputs(83)) or (inputs(248));
    layer0_outputs(1176) <= not(inputs(160));
    layer0_outputs(1177) <= not((inputs(112)) xor (inputs(86)));
    layer0_outputs(1178) <= (inputs(53)) or (inputs(6));
    layer0_outputs(1179) <= (inputs(164)) and not (inputs(45));
    layer0_outputs(1180) <= '1';
    layer0_outputs(1181) <= not((inputs(67)) or (inputs(215)));
    layer0_outputs(1182) <= not((inputs(19)) or (inputs(75)));
    layer0_outputs(1183) <= not(inputs(227));
    layer0_outputs(1184) <= not(inputs(217)) or (inputs(1));
    layer0_outputs(1185) <= not((inputs(197)) xor (inputs(162)));
    layer0_outputs(1186) <= not(inputs(97));
    layer0_outputs(1187) <= (inputs(242)) and not (inputs(129));
    layer0_outputs(1188) <= not(inputs(101));
    layer0_outputs(1189) <= (inputs(127)) and not (inputs(169));
    layer0_outputs(1190) <= not(inputs(212));
    layer0_outputs(1191) <= (inputs(24)) and not (inputs(192));
    layer0_outputs(1192) <= not(inputs(56)) or (inputs(201));
    layer0_outputs(1193) <= not((inputs(12)) xor (inputs(36)));
    layer0_outputs(1194) <= inputs(222);
    layer0_outputs(1195) <= inputs(41);
    layer0_outputs(1196) <= inputs(63);
    layer0_outputs(1197) <= (inputs(246)) and not (inputs(0));
    layer0_outputs(1198) <= inputs(115);
    layer0_outputs(1199) <= not((inputs(198)) xor (inputs(244)));
    layer0_outputs(1200) <= not((inputs(225)) or (inputs(5)));
    layer0_outputs(1201) <= not(inputs(108)) or (inputs(240));
    layer0_outputs(1202) <= (inputs(17)) xor (inputs(11));
    layer0_outputs(1203) <= inputs(74);
    layer0_outputs(1204) <= not((inputs(194)) or (inputs(241)));
    layer0_outputs(1205) <= (inputs(177)) xor (inputs(118));
    layer0_outputs(1206) <= not((inputs(220)) xor (inputs(21)));
    layer0_outputs(1207) <= not((inputs(205)) or (inputs(224)));
    layer0_outputs(1208) <= not(inputs(86)) or (inputs(127));
    layer0_outputs(1209) <= (inputs(247)) and (inputs(222));
    layer0_outputs(1210) <= not((inputs(79)) or (inputs(242)));
    layer0_outputs(1211) <= (inputs(178)) or (inputs(146));
    layer0_outputs(1212) <= (inputs(23)) and not (inputs(227));
    layer0_outputs(1213) <= not((inputs(77)) or (inputs(226)));
    layer0_outputs(1214) <= inputs(35);
    layer0_outputs(1215) <= (inputs(26)) and not (inputs(89));
    layer0_outputs(1216) <= not((inputs(55)) xor (inputs(244)));
    layer0_outputs(1217) <= not(inputs(57)) or (inputs(151));
    layer0_outputs(1218) <= not((inputs(117)) xor (inputs(26)));
    layer0_outputs(1219) <= '1';
    layer0_outputs(1220) <= inputs(194);
    layer0_outputs(1221) <= '0';
    layer0_outputs(1222) <= (inputs(231)) and not (inputs(13));
    layer0_outputs(1223) <= not(inputs(113));
    layer0_outputs(1224) <= (inputs(22)) xor (inputs(156));
    layer0_outputs(1225) <= inputs(88);
    layer0_outputs(1226) <= not(inputs(220));
    layer0_outputs(1227) <= not(inputs(117));
    layer0_outputs(1228) <= inputs(246);
    layer0_outputs(1229) <= (inputs(251)) xor (inputs(196));
    layer0_outputs(1230) <= (inputs(110)) xor (inputs(37));
    layer0_outputs(1231) <= not(inputs(90)) or (inputs(164));
    layer0_outputs(1232) <= not(inputs(8));
    layer0_outputs(1233) <= (inputs(59)) or (inputs(238));
    layer0_outputs(1234) <= (inputs(10)) and not (inputs(220));
    layer0_outputs(1235) <= (inputs(193)) xor (inputs(96));
    layer0_outputs(1236) <= (inputs(118)) and not (inputs(33));
    layer0_outputs(1237) <= (inputs(39)) and not (inputs(192));
    layer0_outputs(1238) <= not(inputs(121)) or (inputs(55));
    layer0_outputs(1239) <= (inputs(132)) xor (inputs(71));
    layer0_outputs(1240) <= inputs(147);
    layer0_outputs(1241) <= (inputs(221)) xor (inputs(202));
    layer0_outputs(1242) <= not((inputs(60)) xor (inputs(189)));
    layer0_outputs(1243) <= not((inputs(203)) and (inputs(162)));
    layer0_outputs(1244) <= not((inputs(95)) or (inputs(191)));
    layer0_outputs(1245) <= not((inputs(53)) or (inputs(216)));
    layer0_outputs(1246) <= not(inputs(204));
    layer0_outputs(1247) <= inputs(213);
    layer0_outputs(1248) <= not(inputs(165));
    layer0_outputs(1249) <= not((inputs(186)) xor (inputs(106)));
    layer0_outputs(1250) <= inputs(107);
    layer0_outputs(1251) <= inputs(67);
    layer0_outputs(1252) <= not(inputs(183)) or (inputs(158));
    layer0_outputs(1253) <= (inputs(254)) or (inputs(177));
    layer0_outputs(1254) <= (inputs(175)) xor (inputs(119));
    layer0_outputs(1255) <= not(inputs(101));
    layer0_outputs(1256) <= not(inputs(180)) or (inputs(63));
    layer0_outputs(1257) <= not(inputs(113));
    layer0_outputs(1258) <= (inputs(49)) or (inputs(6));
    layer0_outputs(1259) <= (inputs(170)) or (inputs(146));
    layer0_outputs(1260) <= not(inputs(138));
    layer0_outputs(1261) <= not(inputs(180));
    layer0_outputs(1262) <= (inputs(152)) xor (inputs(255));
    layer0_outputs(1263) <= not((inputs(235)) or (inputs(227)));
    layer0_outputs(1264) <= inputs(147);
    layer0_outputs(1265) <= inputs(72);
    layer0_outputs(1266) <= not(inputs(198));
    layer0_outputs(1267) <= inputs(115);
    layer0_outputs(1268) <= not(inputs(39));
    layer0_outputs(1269) <= not(inputs(46));
    layer0_outputs(1270) <= not(inputs(155));
    layer0_outputs(1271) <= not((inputs(53)) and (inputs(43)));
    layer0_outputs(1272) <= not((inputs(24)) or (inputs(157)));
    layer0_outputs(1273) <= inputs(10);
    layer0_outputs(1274) <= not(inputs(229)) or (inputs(151));
    layer0_outputs(1275) <= not((inputs(92)) xor (inputs(159)));
    layer0_outputs(1276) <= not(inputs(24));
    layer0_outputs(1277) <= (inputs(213)) xor (inputs(128));
    layer0_outputs(1278) <= not(inputs(151));
    layer0_outputs(1279) <= (inputs(76)) and not (inputs(62));
    layer0_outputs(1280) <= not((inputs(66)) and (inputs(4)));
    layer0_outputs(1281) <= not(inputs(25));
    layer0_outputs(1282) <= (inputs(0)) or (inputs(243));
    layer0_outputs(1283) <= not(inputs(115));
    layer0_outputs(1284) <= (inputs(144)) or (inputs(186));
    layer0_outputs(1285) <= inputs(2);
    layer0_outputs(1286) <= not(inputs(81)) or (inputs(177));
    layer0_outputs(1287) <= (inputs(159)) or (inputs(172));
    layer0_outputs(1288) <= inputs(40);
    layer0_outputs(1289) <= (inputs(86)) xor (inputs(105));
    layer0_outputs(1290) <= inputs(52);
    layer0_outputs(1291) <= (inputs(165)) or (inputs(180));
    layer0_outputs(1292) <= (inputs(51)) or (inputs(254));
    layer0_outputs(1293) <= not((inputs(47)) xor (inputs(15)));
    layer0_outputs(1294) <= not((inputs(6)) xor (inputs(157)));
    layer0_outputs(1295) <= not(inputs(122));
    layer0_outputs(1296) <= (inputs(62)) xor (inputs(189));
    layer0_outputs(1297) <= not((inputs(241)) xor (inputs(80)));
    layer0_outputs(1298) <= (inputs(210)) and not (inputs(8));
    layer0_outputs(1299) <= not((inputs(57)) or (inputs(224)));
    layer0_outputs(1300) <= not((inputs(242)) or (inputs(199)));
    layer0_outputs(1301) <= not(inputs(150)) or (inputs(138));
    layer0_outputs(1302) <= not(inputs(214));
    layer0_outputs(1303) <= (inputs(33)) and not (inputs(82));
    layer0_outputs(1304) <= (inputs(62)) or (inputs(185));
    layer0_outputs(1305) <= inputs(206);
    layer0_outputs(1306) <= (inputs(43)) xor (inputs(87));
    layer0_outputs(1307) <= (inputs(73)) and not (inputs(181));
    layer0_outputs(1308) <= not(inputs(136));
    layer0_outputs(1309) <= not((inputs(230)) and (inputs(232)));
    layer0_outputs(1310) <= not(inputs(144)) or (inputs(63));
    layer0_outputs(1311) <= not(inputs(225));
    layer0_outputs(1312) <= not(inputs(235));
    layer0_outputs(1313) <= inputs(66);
    layer0_outputs(1314) <= (inputs(176)) and not (inputs(142));
    layer0_outputs(1315) <= not((inputs(30)) or (inputs(190)));
    layer0_outputs(1316) <= not(inputs(195)) or (inputs(81));
    layer0_outputs(1317) <= (inputs(44)) or (inputs(92));
    layer0_outputs(1318) <= not((inputs(70)) or (inputs(130)));
    layer0_outputs(1319) <= not((inputs(234)) and (inputs(231)));
    layer0_outputs(1320) <= not(inputs(11));
    layer0_outputs(1321) <= not((inputs(212)) xor (inputs(82)));
    layer0_outputs(1322) <= inputs(111);
    layer0_outputs(1323) <= not(inputs(52)) or (inputs(159));
    layer0_outputs(1324) <= not((inputs(66)) xor (inputs(36)));
    layer0_outputs(1325) <= not(inputs(47)) or (inputs(170));
    layer0_outputs(1326) <= not((inputs(249)) and (inputs(248)));
    layer0_outputs(1327) <= inputs(248);
    layer0_outputs(1328) <= not(inputs(98));
    layer0_outputs(1329) <= (inputs(101)) and not (inputs(96));
    layer0_outputs(1330) <= not((inputs(72)) xor (inputs(60)));
    layer0_outputs(1331) <= not((inputs(32)) xor (inputs(70)));
    layer0_outputs(1332) <= not((inputs(3)) or (inputs(41)));
    layer0_outputs(1333) <= not(inputs(241)) or (inputs(183));
    layer0_outputs(1334) <= not(inputs(152));
    layer0_outputs(1335) <= inputs(107);
    layer0_outputs(1336) <= (inputs(13)) or (inputs(111));
    layer0_outputs(1337) <= (inputs(122)) and not (inputs(28));
    layer0_outputs(1338) <= inputs(238);
    layer0_outputs(1339) <= inputs(209);
    layer0_outputs(1340) <= not((inputs(163)) xor (inputs(80)));
    layer0_outputs(1341) <= (inputs(94)) or (inputs(210));
    layer0_outputs(1342) <= inputs(47);
    layer0_outputs(1343) <= (inputs(201)) or (inputs(129));
    layer0_outputs(1344) <= not((inputs(219)) or (inputs(198)));
    layer0_outputs(1345) <= inputs(214);
    layer0_outputs(1346) <= (inputs(227)) and not (inputs(122));
    layer0_outputs(1347) <= (inputs(8)) and not (inputs(5));
    layer0_outputs(1348) <= not(inputs(24)) or (inputs(158));
    layer0_outputs(1349) <= not((inputs(123)) or (inputs(186)));
    layer0_outputs(1350) <= (inputs(107)) xor (inputs(49));
    layer0_outputs(1351) <= not(inputs(242)) or (inputs(150));
    layer0_outputs(1352) <= inputs(199);
    layer0_outputs(1353) <= (inputs(21)) xor (inputs(95));
    layer0_outputs(1354) <= (inputs(220)) and not (inputs(49));
    layer0_outputs(1355) <= not(inputs(98)) or (inputs(225));
    layer0_outputs(1356) <= not((inputs(69)) or (inputs(78)));
    layer0_outputs(1357) <= not((inputs(236)) or (inputs(47)));
    layer0_outputs(1358) <= (inputs(229)) and not (inputs(108));
    layer0_outputs(1359) <= (inputs(49)) or (inputs(104));
    layer0_outputs(1360) <= not(inputs(88));
    layer0_outputs(1361) <= not(inputs(115)) or (inputs(57));
    layer0_outputs(1362) <= not(inputs(136));
    layer0_outputs(1363) <= not(inputs(150));
    layer0_outputs(1364) <= (inputs(149)) or (inputs(181));
    layer0_outputs(1365) <= not(inputs(77));
    layer0_outputs(1366) <= (inputs(140)) xor (inputs(189));
    layer0_outputs(1367) <= (inputs(190)) and not (inputs(58));
    layer0_outputs(1368) <= not(inputs(66)) or (inputs(128));
    layer0_outputs(1369) <= not(inputs(194)) or (inputs(244));
    layer0_outputs(1370) <= not((inputs(198)) or (inputs(168)));
    layer0_outputs(1371) <= not((inputs(112)) or (inputs(139)));
    layer0_outputs(1372) <= (inputs(49)) or (inputs(83));
    layer0_outputs(1373) <= not(inputs(101));
    layer0_outputs(1374) <= (inputs(71)) and not (inputs(175));
    layer0_outputs(1375) <= (inputs(225)) or (inputs(116));
    layer0_outputs(1376) <= '1';
    layer0_outputs(1377) <= not(inputs(229)) or (inputs(94));
    layer0_outputs(1378) <= (inputs(72)) and (inputs(138));
    layer0_outputs(1379) <= inputs(25);
    layer0_outputs(1380) <= inputs(115);
    layer0_outputs(1381) <= not(inputs(154));
    layer0_outputs(1382) <= inputs(44);
    layer0_outputs(1383) <= (inputs(166)) or (inputs(252));
    layer0_outputs(1384) <= not(inputs(255)) or (inputs(48));
    layer0_outputs(1385) <= (inputs(93)) or (inputs(148));
    layer0_outputs(1386) <= (inputs(171)) and not (inputs(77));
    layer0_outputs(1387) <= (inputs(94)) xor (inputs(240));
    layer0_outputs(1388) <= not(inputs(242));
    layer0_outputs(1389) <= not(inputs(52));
    layer0_outputs(1390) <= not((inputs(63)) xor (inputs(156)));
    layer0_outputs(1391) <= (inputs(98)) and not (inputs(170));
    layer0_outputs(1392) <= not(inputs(161));
    layer0_outputs(1393) <= inputs(82);
    layer0_outputs(1394) <= not((inputs(85)) or (inputs(148)));
    layer0_outputs(1395) <= not(inputs(254));
    layer0_outputs(1396) <= inputs(16);
    layer0_outputs(1397) <= not((inputs(131)) or (inputs(83)));
    layer0_outputs(1398) <= inputs(122);
    layer0_outputs(1399) <= (inputs(41)) and not (inputs(226));
    layer0_outputs(1400) <= not(inputs(121)) or (inputs(252));
    layer0_outputs(1401) <= inputs(230);
    layer0_outputs(1402) <= (inputs(135)) or (inputs(199));
    layer0_outputs(1403) <= inputs(197);
    layer0_outputs(1404) <= not((inputs(19)) xor (inputs(85)));
    layer0_outputs(1405) <= not((inputs(217)) or (inputs(244)));
    layer0_outputs(1406) <= not(inputs(122)) or (inputs(206));
    layer0_outputs(1407) <= inputs(76);
    layer0_outputs(1408) <= '0';
    layer0_outputs(1409) <= inputs(44);
    layer0_outputs(1410) <= not((inputs(30)) and (inputs(210)));
    layer0_outputs(1411) <= not((inputs(172)) xor (inputs(17)));
    layer0_outputs(1412) <= (inputs(98)) and not (inputs(140));
    layer0_outputs(1413) <= inputs(208);
    layer0_outputs(1414) <= (inputs(81)) or (inputs(9));
    layer0_outputs(1415) <= (inputs(242)) and (inputs(90));
    layer0_outputs(1416) <= not(inputs(243));
    layer0_outputs(1417) <= (inputs(226)) xor (inputs(158));
    layer0_outputs(1418) <= (inputs(237)) and not (inputs(157));
    layer0_outputs(1419) <= (inputs(40)) or (inputs(32));
    layer0_outputs(1420) <= (inputs(19)) and not (inputs(66));
    layer0_outputs(1421) <= (inputs(50)) and (inputs(234));
    layer0_outputs(1422) <= (inputs(9)) or (inputs(165));
    layer0_outputs(1423) <= (inputs(247)) or (inputs(144));
    layer0_outputs(1424) <= (inputs(142)) xor (inputs(74));
    layer0_outputs(1425) <= (inputs(88)) xor (inputs(152));
    layer0_outputs(1426) <= not(inputs(101));
    layer0_outputs(1427) <= not(inputs(165));
    layer0_outputs(1428) <= not((inputs(153)) or (inputs(198)));
    layer0_outputs(1429) <= (inputs(101)) xor (inputs(206));
    layer0_outputs(1430) <= (inputs(193)) xor (inputs(161));
    layer0_outputs(1431) <= not((inputs(27)) or (inputs(26)));
    layer0_outputs(1432) <= not((inputs(252)) or (inputs(7)));
    layer0_outputs(1433) <= (inputs(225)) or (inputs(227));
    layer0_outputs(1434) <= (inputs(163)) and not (inputs(1));
    layer0_outputs(1435) <= not(inputs(105));
    layer0_outputs(1436) <= not(inputs(246));
    layer0_outputs(1437) <= inputs(209);
    layer0_outputs(1438) <= inputs(240);
    layer0_outputs(1439) <= not(inputs(178)) or (inputs(47));
    layer0_outputs(1440) <= not(inputs(187)) or (inputs(67));
    layer0_outputs(1441) <= not(inputs(130));
    layer0_outputs(1442) <= (inputs(105)) and not (inputs(95));
    layer0_outputs(1443) <= not((inputs(111)) xor (inputs(200)));
    layer0_outputs(1444) <= (inputs(29)) or (inputs(120));
    layer0_outputs(1445) <= inputs(43);
    layer0_outputs(1446) <= inputs(30);
    layer0_outputs(1447) <= (inputs(154)) and not (inputs(65));
    layer0_outputs(1448) <= '1';
    layer0_outputs(1449) <= not((inputs(232)) xor (inputs(22)));
    layer0_outputs(1450) <= (inputs(124)) or (inputs(189));
    layer0_outputs(1451) <= not((inputs(56)) xor (inputs(59)));
    layer0_outputs(1452) <= '0';
    layer0_outputs(1453) <= (inputs(85)) xor (inputs(253));
    layer0_outputs(1454) <= not(inputs(245)) or (inputs(17));
    layer0_outputs(1455) <= not(inputs(214));
    layer0_outputs(1456) <= not(inputs(166));
    layer0_outputs(1457) <= not((inputs(91)) xor (inputs(105)));
    layer0_outputs(1458) <= (inputs(111)) and (inputs(218));
    layer0_outputs(1459) <= not(inputs(117));
    layer0_outputs(1460) <= inputs(7);
    layer0_outputs(1461) <= not(inputs(76)) or (inputs(212));
    layer0_outputs(1462) <= (inputs(12)) or (inputs(50));
    layer0_outputs(1463) <= not((inputs(144)) or (inputs(165)));
    layer0_outputs(1464) <= '1';
    layer0_outputs(1465) <= inputs(118);
    layer0_outputs(1466) <= not(inputs(14)) or (inputs(221));
    layer0_outputs(1467) <= not((inputs(21)) or (inputs(84)));
    layer0_outputs(1468) <= '1';
    layer0_outputs(1469) <= not(inputs(174));
    layer0_outputs(1470) <= not((inputs(211)) xor (inputs(128)));
    layer0_outputs(1471) <= inputs(121);
    layer0_outputs(1472) <= not((inputs(206)) or (inputs(86)));
    layer0_outputs(1473) <= (inputs(168)) xor (inputs(161));
    layer0_outputs(1474) <= (inputs(50)) and (inputs(159));
    layer0_outputs(1475) <= not(inputs(71));
    layer0_outputs(1476) <= not(inputs(232)) or (inputs(125));
    layer0_outputs(1477) <= (inputs(222)) and not (inputs(55));
    layer0_outputs(1478) <= (inputs(188)) and not (inputs(36));
    layer0_outputs(1479) <= (inputs(229)) and not (inputs(131));
    layer0_outputs(1480) <= not(inputs(77));
    layer0_outputs(1481) <= not(inputs(173)) or (inputs(113));
    layer0_outputs(1482) <= (inputs(57)) and not (inputs(20));
    layer0_outputs(1483) <= not((inputs(185)) or (inputs(142)));
    layer0_outputs(1484) <= (inputs(201)) xor (inputs(31));
    layer0_outputs(1485) <= not((inputs(195)) and (inputs(156)));
    layer0_outputs(1486) <= inputs(85);
    layer0_outputs(1487) <= (inputs(170)) xor (inputs(226));
    layer0_outputs(1488) <= not(inputs(75));
    layer0_outputs(1489) <= inputs(224);
    layer0_outputs(1490) <= not(inputs(252));
    layer0_outputs(1491) <= (inputs(27)) and not (inputs(163));
    layer0_outputs(1492) <= (inputs(115)) and not (inputs(226));
    layer0_outputs(1493) <= not(inputs(79));
    layer0_outputs(1494) <= not((inputs(254)) xor (inputs(182)));
    layer0_outputs(1495) <= not((inputs(151)) and (inputs(41)));
    layer0_outputs(1496) <= not(inputs(100));
    layer0_outputs(1497) <= (inputs(148)) or (inputs(117));
    layer0_outputs(1498) <= not(inputs(90));
    layer0_outputs(1499) <= not((inputs(19)) xor (inputs(232)));
    layer0_outputs(1500) <= (inputs(138)) and not (inputs(2));
    layer0_outputs(1501) <= (inputs(13)) and not (inputs(244));
    layer0_outputs(1502) <= not(inputs(115));
    layer0_outputs(1503) <= not((inputs(252)) xor (inputs(182)));
    layer0_outputs(1504) <= not((inputs(192)) or (inputs(12)));
    layer0_outputs(1505) <= (inputs(182)) and not (inputs(108));
    layer0_outputs(1506) <= not((inputs(79)) or (inputs(187)));
    layer0_outputs(1507) <= inputs(226);
    layer0_outputs(1508) <= inputs(201);
    layer0_outputs(1509) <= (inputs(85)) and not (inputs(5));
    layer0_outputs(1510) <= inputs(233);
    layer0_outputs(1511) <= (inputs(48)) xor (inputs(186));
    layer0_outputs(1512) <= '1';
    layer0_outputs(1513) <= (inputs(49)) or (inputs(35));
    layer0_outputs(1514) <= not(inputs(114)) or (inputs(65));
    layer0_outputs(1515) <= inputs(103);
    layer0_outputs(1516) <= not((inputs(126)) or (inputs(18)));
    layer0_outputs(1517) <= (inputs(121)) or (inputs(133));
    layer0_outputs(1518) <= not((inputs(255)) xor (inputs(93)));
    layer0_outputs(1519) <= not(inputs(69)) or (inputs(243));
    layer0_outputs(1520) <= (inputs(192)) xor (inputs(246));
    layer0_outputs(1521) <= not(inputs(80)) or (inputs(73));
    layer0_outputs(1522) <= '1';
    layer0_outputs(1523) <= (inputs(205)) xor (inputs(4));
    layer0_outputs(1524) <= not(inputs(237)) or (inputs(103));
    layer0_outputs(1525) <= (inputs(5)) and not (inputs(250));
    layer0_outputs(1526) <= not((inputs(147)) or (inputs(52)));
    layer0_outputs(1527) <= (inputs(61)) and not (inputs(114));
    layer0_outputs(1528) <= not((inputs(42)) and (inputs(21)));
    layer0_outputs(1529) <= not((inputs(148)) xor (inputs(108)));
    layer0_outputs(1530) <= not((inputs(35)) or (inputs(223)));
    layer0_outputs(1531) <= (inputs(123)) or (inputs(178));
    layer0_outputs(1532) <= (inputs(184)) and (inputs(251));
    layer0_outputs(1533) <= (inputs(81)) or (inputs(91));
    layer0_outputs(1534) <= not(inputs(67));
    layer0_outputs(1535) <= not(inputs(196)) or (inputs(91));
    layer0_outputs(1536) <= not(inputs(79));
    layer0_outputs(1537) <= inputs(152);
    layer0_outputs(1538) <= (inputs(29)) and not (inputs(255));
    layer0_outputs(1539) <= (inputs(86)) and not (inputs(94));
    layer0_outputs(1540) <= (inputs(211)) xor (inputs(119));
    layer0_outputs(1541) <= not((inputs(28)) and (inputs(205)));
    layer0_outputs(1542) <= (inputs(26)) and not (inputs(249));
    layer0_outputs(1543) <= not((inputs(46)) or (inputs(9)));
    layer0_outputs(1544) <= (inputs(218)) and not (inputs(190));
    layer0_outputs(1545) <= inputs(29);
    layer0_outputs(1546) <= not(inputs(89));
    layer0_outputs(1547) <= not(inputs(218));
    layer0_outputs(1548) <= not(inputs(214));
    layer0_outputs(1549) <= (inputs(175)) or (inputs(56));
    layer0_outputs(1550) <= (inputs(176)) or (inputs(177));
    layer0_outputs(1551) <= (inputs(116)) xor (inputs(196));
    layer0_outputs(1552) <= not(inputs(238));
    layer0_outputs(1553) <= not(inputs(51)) or (inputs(2));
    layer0_outputs(1554) <= (inputs(113)) and not (inputs(78));
    layer0_outputs(1555) <= (inputs(214)) xor (inputs(242));
    layer0_outputs(1556) <= not((inputs(161)) xor (inputs(22)));
    layer0_outputs(1557) <= not(inputs(76));
    layer0_outputs(1558) <= (inputs(44)) and not (inputs(25));
    layer0_outputs(1559) <= (inputs(77)) or (inputs(228));
    layer0_outputs(1560) <= (inputs(17)) xor (inputs(97));
    layer0_outputs(1561) <= (inputs(19)) and not (inputs(176));
    layer0_outputs(1562) <= inputs(11);
    layer0_outputs(1563) <= not(inputs(179));
    layer0_outputs(1564) <= (inputs(58)) xor (inputs(233));
    layer0_outputs(1565) <= inputs(176);
    layer0_outputs(1566) <= not(inputs(201));
    layer0_outputs(1567) <= (inputs(64)) and not (inputs(20));
    layer0_outputs(1568) <= not((inputs(248)) or (inputs(81)));
    layer0_outputs(1569) <= inputs(226);
    layer0_outputs(1570) <= not((inputs(76)) or (inputs(81)));
    layer0_outputs(1571) <= (inputs(255)) xor (inputs(225));
    layer0_outputs(1572) <= not(inputs(84));
    layer0_outputs(1573) <= (inputs(196)) and not (inputs(46));
    layer0_outputs(1574) <= not(inputs(56)) or (inputs(70));
    layer0_outputs(1575) <= (inputs(41)) and not (inputs(87));
    layer0_outputs(1576) <= not(inputs(212)) or (inputs(198));
    layer0_outputs(1577) <= not(inputs(7));
    layer0_outputs(1578) <= (inputs(137)) and not (inputs(218));
    layer0_outputs(1579) <= (inputs(182)) and not (inputs(107));
    layer0_outputs(1580) <= not((inputs(51)) or (inputs(93)));
    layer0_outputs(1581) <= (inputs(206)) and not (inputs(239));
    layer0_outputs(1582) <= not(inputs(55));
    layer0_outputs(1583) <= not(inputs(41)) or (inputs(128));
    layer0_outputs(1584) <= not(inputs(11));
    layer0_outputs(1585) <= (inputs(61)) or (inputs(119));
    layer0_outputs(1586) <= (inputs(145)) or (inputs(3));
    layer0_outputs(1587) <= (inputs(74)) and not (inputs(204));
    layer0_outputs(1588) <= inputs(211);
    layer0_outputs(1589) <= not(inputs(150));
    layer0_outputs(1590) <= (inputs(174)) and not (inputs(127));
    layer0_outputs(1591) <= '1';
    layer0_outputs(1592) <= (inputs(148)) xor (inputs(247));
    layer0_outputs(1593) <= inputs(159);
    layer0_outputs(1594) <= not((inputs(153)) or (inputs(13)));
    layer0_outputs(1595) <= not(inputs(188)) or (inputs(232));
    layer0_outputs(1596) <= not((inputs(151)) or (inputs(3)));
    layer0_outputs(1597) <= inputs(130);
    layer0_outputs(1598) <= inputs(146);
    layer0_outputs(1599) <= (inputs(37)) xor (inputs(73));
    layer0_outputs(1600) <= (inputs(135)) or (inputs(146));
    layer0_outputs(1601) <= (inputs(210)) and not (inputs(16));
    layer0_outputs(1602) <= not((inputs(229)) or (inputs(84)));
    layer0_outputs(1603) <= (inputs(127)) or (inputs(190));
    layer0_outputs(1604) <= not(inputs(217)) or (inputs(113));
    layer0_outputs(1605) <= (inputs(185)) xor (inputs(246));
    layer0_outputs(1606) <= (inputs(154)) xor (inputs(19));
    layer0_outputs(1607) <= not((inputs(229)) or (inputs(213)));
    layer0_outputs(1608) <= (inputs(124)) or (inputs(19));
    layer0_outputs(1609) <= not((inputs(52)) or (inputs(2)));
    layer0_outputs(1610) <= not(inputs(205));
    layer0_outputs(1611) <= not(inputs(21)) or (inputs(102));
    layer0_outputs(1612) <= not((inputs(51)) or (inputs(66)));
    layer0_outputs(1613) <= inputs(169);
    layer0_outputs(1614) <= (inputs(198)) and (inputs(60));
    layer0_outputs(1615) <= not(inputs(10));
    layer0_outputs(1616) <= inputs(244);
    layer0_outputs(1617) <= not(inputs(212)) or (inputs(95));
    layer0_outputs(1618) <= not(inputs(89)) or (inputs(34));
    layer0_outputs(1619) <= (inputs(115)) and not (inputs(93));
    layer0_outputs(1620) <= (inputs(58)) or (inputs(20));
    layer0_outputs(1621) <= not((inputs(154)) and (inputs(176)));
    layer0_outputs(1622) <= not(inputs(44));
    layer0_outputs(1623) <= not((inputs(249)) or (inputs(211)));
    layer0_outputs(1624) <= (inputs(47)) or (inputs(138));
    layer0_outputs(1625) <= inputs(97);
    layer0_outputs(1626) <= (inputs(90)) or (inputs(17));
    layer0_outputs(1627) <= inputs(99);
    layer0_outputs(1628) <= not(inputs(140));
    layer0_outputs(1629) <= inputs(182);
    layer0_outputs(1630) <= not(inputs(0));
    layer0_outputs(1631) <= inputs(173);
    layer0_outputs(1632) <= inputs(221);
    layer0_outputs(1633) <= (inputs(64)) or (inputs(233));
    layer0_outputs(1634) <= (inputs(150)) and (inputs(86));
    layer0_outputs(1635) <= not(inputs(188));
    layer0_outputs(1636) <= inputs(193);
    layer0_outputs(1637) <= (inputs(80)) xor (inputs(248));
    layer0_outputs(1638) <= (inputs(194)) and not (inputs(13));
    layer0_outputs(1639) <= (inputs(2)) xor (inputs(192));
    layer0_outputs(1640) <= not((inputs(32)) or (inputs(190)));
    layer0_outputs(1641) <= not(inputs(161));
    layer0_outputs(1642) <= inputs(230);
    layer0_outputs(1643) <= not(inputs(122)) or (inputs(33));
    layer0_outputs(1644) <= not((inputs(245)) or (inputs(218)));
    layer0_outputs(1645) <= (inputs(121)) and not (inputs(84));
    layer0_outputs(1646) <= (inputs(11)) and not (inputs(81));
    layer0_outputs(1647) <= inputs(97);
    layer0_outputs(1648) <= not((inputs(15)) or (inputs(73)));
    layer0_outputs(1649) <= inputs(91);
    layer0_outputs(1650) <= (inputs(151)) or (inputs(135));
    layer0_outputs(1651) <= not((inputs(49)) or (inputs(36)));
    layer0_outputs(1652) <= inputs(74);
    layer0_outputs(1653) <= not((inputs(17)) or (inputs(148)));
    layer0_outputs(1654) <= inputs(136);
    layer0_outputs(1655) <= inputs(151);
    layer0_outputs(1656) <= (inputs(143)) and not (inputs(50));
    layer0_outputs(1657) <= not((inputs(234)) or (inputs(206)));
    layer0_outputs(1658) <= not(inputs(153));
    layer0_outputs(1659) <= not((inputs(252)) xor (inputs(53)));
    layer0_outputs(1660) <= inputs(117);
    layer0_outputs(1661) <= not((inputs(47)) or (inputs(40)));
    layer0_outputs(1662) <= not((inputs(222)) or (inputs(220)));
    layer0_outputs(1663) <= (inputs(28)) and not (inputs(202));
    layer0_outputs(1664) <= inputs(156);
    layer0_outputs(1665) <= not(inputs(228));
    layer0_outputs(1666) <= (inputs(37)) and not (inputs(214));
    layer0_outputs(1667) <= '0';
    layer0_outputs(1668) <= (inputs(181)) or (inputs(48));
    layer0_outputs(1669) <= (inputs(188)) or (inputs(145));
    layer0_outputs(1670) <= (inputs(22)) and not (inputs(159));
    layer0_outputs(1671) <= not(inputs(7)) or (inputs(29));
    layer0_outputs(1672) <= not(inputs(174));
    layer0_outputs(1673) <= inputs(107);
    layer0_outputs(1674) <= (inputs(182)) and not (inputs(192));
    layer0_outputs(1675) <= not((inputs(161)) xor (inputs(163)));
    layer0_outputs(1676) <= not(inputs(148));
    layer0_outputs(1677) <= not(inputs(200)) or (inputs(125));
    layer0_outputs(1678) <= (inputs(238)) xor (inputs(204));
    layer0_outputs(1679) <= (inputs(27)) xor (inputs(109));
    layer0_outputs(1680) <= (inputs(48)) or (inputs(162));
    layer0_outputs(1681) <= (inputs(152)) or (inputs(107));
    layer0_outputs(1682) <= (inputs(138)) xor (inputs(188));
    layer0_outputs(1683) <= '0';
    layer0_outputs(1684) <= (inputs(73)) and not (inputs(14));
    layer0_outputs(1685) <= inputs(221);
    layer0_outputs(1686) <= (inputs(127)) or (inputs(94));
    layer0_outputs(1687) <= not(inputs(182));
    layer0_outputs(1688) <= not(inputs(205));
    layer0_outputs(1689) <= (inputs(161)) xor (inputs(69));
    layer0_outputs(1690) <= not(inputs(62));
    layer0_outputs(1691) <= not(inputs(73)) or (inputs(34));
    layer0_outputs(1692) <= inputs(136);
    layer0_outputs(1693) <= not((inputs(189)) xor (inputs(113)));
    layer0_outputs(1694) <= not(inputs(217));
    layer0_outputs(1695) <= inputs(105);
    layer0_outputs(1696) <= (inputs(183)) and not (inputs(91));
    layer0_outputs(1697) <= (inputs(22)) and not (inputs(79));
    layer0_outputs(1698) <= inputs(140);
    layer0_outputs(1699) <= not(inputs(98));
    layer0_outputs(1700) <= not((inputs(188)) xor (inputs(16)));
    layer0_outputs(1701) <= (inputs(110)) and not (inputs(226));
    layer0_outputs(1702) <= '0';
    layer0_outputs(1703) <= not((inputs(3)) xor (inputs(49)));
    layer0_outputs(1704) <= not((inputs(238)) or (inputs(94)));
    layer0_outputs(1705) <= not((inputs(33)) or (inputs(186)));
    layer0_outputs(1706) <= inputs(14);
    layer0_outputs(1707) <= (inputs(19)) and not (inputs(82));
    layer0_outputs(1708) <= (inputs(20)) and (inputs(223));
    layer0_outputs(1709) <= not(inputs(227)) or (inputs(26));
    layer0_outputs(1710) <= not(inputs(4));
    layer0_outputs(1711) <= (inputs(59)) or (inputs(70));
    layer0_outputs(1712) <= inputs(215);
    layer0_outputs(1713) <= inputs(107);
    layer0_outputs(1714) <= not((inputs(150)) or (inputs(238)));
    layer0_outputs(1715) <= (inputs(68)) and not (inputs(112));
    layer0_outputs(1716) <= not(inputs(14));
    layer0_outputs(1717) <= inputs(14);
    layer0_outputs(1718) <= not(inputs(50));
    layer0_outputs(1719) <= (inputs(89)) and not (inputs(226));
    layer0_outputs(1720) <= '1';
    layer0_outputs(1721) <= not((inputs(220)) or (inputs(178)));
    layer0_outputs(1722) <= (inputs(221)) or (inputs(33));
    layer0_outputs(1723) <= (inputs(179)) and not (inputs(144));
    layer0_outputs(1724) <= (inputs(158)) and not (inputs(185));
    layer0_outputs(1725) <= (inputs(94)) xor (inputs(75));
    layer0_outputs(1726) <= (inputs(156)) and not (inputs(41));
    layer0_outputs(1727) <= (inputs(78)) xor (inputs(108));
    layer0_outputs(1728) <= not(inputs(189)) or (inputs(211));
    layer0_outputs(1729) <= inputs(250);
    layer0_outputs(1730) <= (inputs(161)) or (inputs(221));
    layer0_outputs(1731) <= not(inputs(121)) or (inputs(209));
    layer0_outputs(1732) <= not((inputs(69)) and (inputs(203)));
    layer0_outputs(1733) <= (inputs(127)) or (inputs(122));
    layer0_outputs(1734) <= inputs(92);
    layer0_outputs(1735) <= not(inputs(12)) or (inputs(161));
    layer0_outputs(1736) <= (inputs(196)) xor (inputs(32));
    layer0_outputs(1737) <= (inputs(49)) xor (inputs(53));
    layer0_outputs(1738) <= inputs(176);
    layer0_outputs(1739) <= not((inputs(137)) xor (inputs(190)));
    layer0_outputs(1740) <= inputs(129);
    layer0_outputs(1741) <= (inputs(74)) or (inputs(1));
    layer0_outputs(1742) <= (inputs(200)) and not (inputs(94));
    layer0_outputs(1743) <= not(inputs(212)) or (inputs(75));
    layer0_outputs(1744) <= inputs(25);
    layer0_outputs(1745) <= inputs(92);
    layer0_outputs(1746) <= (inputs(44)) and not (inputs(186));
    layer0_outputs(1747) <= not(inputs(171));
    layer0_outputs(1748) <= not(inputs(228));
    layer0_outputs(1749) <= not(inputs(67));
    layer0_outputs(1750) <= inputs(190);
    layer0_outputs(1751) <= (inputs(12)) and not (inputs(35));
    layer0_outputs(1752) <= (inputs(38)) or (inputs(155));
    layer0_outputs(1753) <= not(inputs(105));
    layer0_outputs(1754) <= not(inputs(183));
    layer0_outputs(1755) <= inputs(57);
    layer0_outputs(1756) <= (inputs(2)) xor (inputs(237));
    layer0_outputs(1757) <= not(inputs(150)) or (inputs(170));
    layer0_outputs(1758) <= '1';
    layer0_outputs(1759) <= not(inputs(129)) or (inputs(72));
    layer0_outputs(1760) <= inputs(21);
    layer0_outputs(1761) <= not((inputs(119)) or (inputs(34)));
    layer0_outputs(1762) <= (inputs(25)) or (inputs(10));
    layer0_outputs(1763) <= (inputs(253)) or (inputs(89));
    layer0_outputs(1764) <= (inputs(10)) and not (inputs(215));
    layer0_outputs(1765) <= (inputs(128)) or (inputs(191));
    layer0_outputs(1766) <= not((inputs(52)) or (inputs(218)));
    layer0_outputs(1767) <= inputs(167);
    layer0_outputs(1768) <= not(inputs(221)) or (inputs(158));
    layer0_outputs(1769) <= not((inputs(42)) xor (inputs(50)));
    layer0_outputs(1770) <= not(inputs(224)) or (inputs(26));
    layer0_outputs(1771) <= inputs(129);
    layer0_outputs(1772) <= not(inputs(151));
    layer0_outputs(1773) <= not(inputs(105)) or (inputs(190));
    layer0_outputs(1774) <= (inputs(44)) or (inputs(204));
    layer0_outputs(1775) <= inputs(145);
    layer0_outputs(1776) <= inputs(210);
    layer0_outputs(1777) <= '1';
    layer0_outputs(1778) <= not(inputs(62));
    layer0_outputs(1779) <= not(inputs(198)) or (inputs(39));
    layer0_outputs(1780) <= not(inputs(58)) or (inputs(239));
    layer0_outputs(1781) <= not((inputs(102)) xor (inputs(23)));
    layer0_outputs(1782) <= not((inputs(141)) xor (inputs(81)));
    layer0_outputs(1783) <= inputs(212);
    layer0_outputs(1784) <= not((inputs(173)) xor (inputs(25)));
    layer0_outputs(1785) <= not((inputs(209)) xor (inputs(239)));
    layer0_outputs(1786) <= not(inputs(11)) or (inputs(218));
    layer0_outputs(1787) <= (inputs(82)) or (inputs(195));
    layer0_outputs(1788) <= not(inputs(178)) or (inputs(17));
    layer0_outputs(1789) <= (inputs(102)) and (inputs(66));
    layer0_outputs(1790) <= (inputs(180)) and not (inputs(114));
    layer0_outputs(1791) <= not(inputs(38));
    layer0_outputs(1792) <= '0';
    layer0_outputs(1793) <= (inputs(117)) xor (inputs(189));
    layer0_outputs(1794) <= inputs(147);
    layer0_outputs(1795) <= not(inputs(130));
    layer0_outputs(1796) <= inputs(147);
    layer0_outputs(1797) <= not((inputs(77)) or (inputs(84)));
    layer0_outputs(1798) <= (inputs(191)) or (inputs(189));
    layer0_outputs(1799) <= not(inputs(179));
    layer0_outputs(1800) <= not(inputs(51));
    layer0_outputs(1801) <= not((inputs(82)) and (inputs(71)));
    layer0_outputs(1802) <= '1';
    layer0_outputs(1803) <= (inputs(224)) or (inputs(174));
    layer0_outputs(1804) <= inputs(29);
    layer0_outputs(1805) <= not((inputs(101)) or (inputs(99)));
    layer0_outputs(1806) <= not(inputs(210)) or (inputs(74));
    layer0_outputs(1807) <= not((inputs(61)) or (inputs(104)));
    layer0_outputs(1808) <= inputs(213);
    layer0_outputs(1809) <= (inputs(20)) xor (inputs(112));
    layer0_outputs(1810) <= inputs(28);
    layer0_outputs(1811) <= not((inputs(51)) xor (inputs(196)));
    layer0_outputs(1812) <= (inputs(137)) xor (inputs(171));
    layer0_outputs(1813) <= not((inputs(167)) or (inputs(2)));
    layer0_outputs(1814) <= (inputs(111)) xor (inputs(84));
    layer0_outputs(1815) <= (inputs(6)) and (inputs(127));
    layer0_outputs(1816) <= (inputs(244)) and not (inputs(4));
    layer0_outputs(1817) <= inputs(101);
    layer0_outputs(1818) <= not((inputs(142)) or (inputs(218)));
    layer0_outputs(1819) <= not(inputs(230));
    layer0_outputs(1820) <= not((inputs(94)) or (inputs(170)));
    layer0_outputs(1821) <= not((inputs(70)) xor (inputs(205)));
    layer0_outputs(1822) <= not((inputs(42)) or (inputs(227)));
    layer0_outputs(1823) <= inputs(202);
    layer0_outputs(1824) <= not((inputs(0)) or (inputs(69)));
    layer0_outputs(1825) <= (inputs(163)) xor (inputs(110));
    layer0_outputs(1826) <= not(inputs(231)) or (inputs(48));
    layer0_outputs(1827) <= not(inputs(138)) or (inputs(205));
    layer0_outputs(1828) <= inputs(119);
    layer0_outputs(1829) <= inputs(221);
    layer0_outputs(1830) <= not((inputs(46)) or (inputs(93)));
    layer0_outputs(1831) <= not((inputs(92)) or (inputs(78)));
    layer0_outputs(1832) <= not(inputs(166));
    layer0_outputs(1833) <= inputs(129);
    layer0_outputs(1834) <= inputs(83);
    layer0_outputs(1835) <= (inputs(191)) or (inputs(216));
    layer0_outputs(1836) <= (inputs(26)) and not (inputs(184));
    layer0_outputs(1837) <= (inputs(96)) or (inputs(237));
    layer0_outputs(1838) <= (inputs(196)) or (inputs(187));
    layer0_outputs(1839) <= not((inputs(246)) xor (inputs(79)));
    layer0_outputs(1840) <= not((inputs(217)) and (inputs(44)));
    layer0_outputs(1841) <= not(inputs(22));
    layer0_outputs(1842) <= not((inputs(212)) or (inputs(41)));
    layer0_outputs(1843) <= not(inputs(90));
    layer0_outputs(1844) <= (inputs(65)) or (inputs(47));
    layer0_outputs(1845) <= not(inputs(127));
    layer0_outputs(1846) <= not(inputs(145)) or (inputs(13));
    layer0_outputs(1847) <= not((inputs(235)) or (inputs(217)));
    layer0_outputs(1848) <= not((inputs(96)) xor (inputs(118)));
    layer0_outputs(1849) <= inputs(118);
    layer0_outputs(1850) <= not((inputs(138)) or (inputs(241)));
    layer0_outputs(1851) <= inputs(165);
    layer0_outputs(1852) <= not(inputs(22));
    layer0_outputs(1853) <= inputs(170);
    layer0_outputs(1854) <= not((inputs(20)) xor (inputs(65)));
    layer0_outputs(1855) <= (inputs(205)) xor (inputs(151));
    layer0_outputs(1856) <= not((inputs(18)) or (inputs(18)));
    layer0_outputs(1857) <= not((inputs(202)) or (inputs(243)));
    layer0_outputs(1858) <= not(inputs(137));
    layer0_outputs(1859) <= (inputs(163)) and (inputs(117));
    layer0_outputs(1860) <= not((inputs(69)) xor (inputs(68)));
    layer0_outputs(1861) <= inputs(197);
    layer0_outputs(1862) <= not(inputs(98));
    layer0_outputs(1863) <= (inputs(182)) or (inputs(0));
    layer0_outputs(1864) <= inputs(79);
    layer0_outputs(1865) <= (inputs(169)) and (inputs(81));
    layer0_outputs(1866) <= inputs(234);
    layer0_outputs(1867) <= not((inputs(42)) and (inputs(39)));
    layer0_outputs(1868) <= not(inputs(58)) or (inputs(71));
    layer0_outputs(1869) <= inputs(133);
    layer0_outputs(1870) <= not(inputs(179)) or (inputs(112));
    layer0_outputs(1871) <= not(inputs(225));
    layer0_outputs(1872) <= not(inputs(9));
    layer0_outputs(1873) <= not(inputs(147));
    layer0_outputs(1874) <= not((inputs(58)) or (inputs(127)));
    layer0_outputs(1875) <= inputs(216);
    layer0_outputs(1876) <= inputs(161);
    layer0_outputs(1877) <= inputs(133);
    layer0_outputs(1878) <= inputs(39);
    layer0_outputs(1879) <= not((inputs(97)) xor (inputs(149)));
    layer0_outputs(1880) <= not((inputs(251)) and (inputs(111)));
    layer0_outputs(1881) <= (inputs(44)) xor (inputs(76));
    layer0_outputs(1882) <= (inputs(59)) and not (inputs(38));
    layer0_outputs(1883) <= (inputs(117)) and (inputs(68));
    layer0_outputs(1884) <= (inputs(118)) xor (inputs(215));
    layer0_outputs(1885) <= not((inputs(92)) xor (inputs(74)));
    layer0_outputs(1886) <= inputs(7);
    layer0_outputs(1887) <= (inputs(20)) and not (inputs(11));
    layer0_outputs(1888) <= (inputs(136)) and not (inputs(91));
    layer0_outputs(1889) <= (inputs(175)) and not (inputs(138));
    layer0_outputs(1890) <= not((inputs(32)) xor (inputs(245)));
    layer0_outputs(1891) <= (inputs(156)) and not (inputs(95));
    layer0_outputs(1892) <= not((inputs(246)) xor (inputs(92)));
    layer0_outputs(1893) <= not(inputs(149)) or (inputs(78));
    layer0_outputs(1894) <= not(inputs(52));
    layer0_outputs(1895) <= not(inputs(74));
    layer0_outputs(1896) <= not((inputs(108)) xor (inputs(144)));
    layer0_outputs(1897) <= (inputs(180)) and not (inputs(142));
    layer0_outputs(1898) <= not((inputs(228)) and (inputs(173)));
    layer0_outputs(1899) <= inputs(146);
    layer0_outputs(1900) <= not((inputs(88)) xor (inputs(167)));
    layer0_outputs(1901) <= not((inputs(11)) or (inputs(79)));
    layer0_outputs(1902) <= (inputs(154)) and not (inputs(236));
    layer0_outputs(1903) <= (inputs(56)) and not (inputs(186));
    layer0_outputs(1904) <= not(inputs(54));
    layer0_outputs(1905) <= (inputs(55)) and not (inputs(171));
    layer0_outputs(1906) <= not(inputs(152)) or (inputs(66));
    layer0_outputs(1907) <= inputs(230);
    layer0_outputs(1908) <= not(inputs(230));
    layer0_outputs(1909) <= not(inputs(13));
    layer0_outputs(1910) <= not(inputs(101));
    layer0_outputs(1911) <= inputs(186);
    layer0_outputs(1912) <= not((inputs(96)) or (inputs(100)));
    layer0_outputs(1913) <= inputs(233);
    layer0_outputs(1914) <= not(inputs(39));
    layer0_outputs(1915) <= not(inputs(77)) or (inputs(158));
    layer0_outputs(1916) <= not(inputs(149)) or (inputs(35));
    layer0_outputs(1917) <= not((inputs(156)) xor (inputs(206)));
    layer0_outputs(1918) <= (inputs(153)) and not (inputs(98));
    layer0_outputs(1919) <= inputs(135);
    layer0_outputs(1920) <= inputs(170);
    layer0_outputs(1921) <= (inputs(222)) xor (inputs(228));
    layer0_outputs(1922) <= inputs(193);
    layer0_outputs(1923) <= inputs(25);
    layer0_outputs(1924) <= (inputs(113)) xor (inputs(99));
    layer0_outputs(1925) <= not((inputs(238)) or (inputs(29)));
    layer0_outputs(1926) <= (inputs(125)) or (inputs(250));
    layer0_outputs(1927) <= inputs(75);
    layer0_outputs(1928) <= inputs(108);
    layer0_outputs(1929) <= (inputs(255)) xor (inputs(10));
    layer0_outputs(1930) <= not((inputs(220)) or (inputs(170)));
    layer0_outputs(1931) <= not((inputs(184)) xor (inputs(233)));
    layer0_outputs(1932) <= (inputs(150)) xor (inputs(47));
    layer0_outputs(1933) <= not((inputs(126)) or (inputs(82)));
    layer0_outputs(1934) <= inputs(102);
    layer0_outputs(1935) <= not(inputs(78));
    layer0_outputs(1936) <= not((inputs(193)) or (inputs(210)));
    layer0_outputs(1937) <= (inputs(89)) xor (inputs(152));
    layer0_outputs(1938) <= not((inputs(108)) or (inputs(84)));
    layer0_outputs(1939) <= (inputs(244)) and not (inputs(96));
    layer0_outputs(1940) <= not((inputs(58)) xor (inputs(179)));
    layer0_outputs(1941) <= inputs(253);
    layer0_outputs(1942) <= not((inputs(244)) and (inputs(31)));
    layer0_outputs(1943) <= (inputs(27)) and not (inputs(17));
    layer0_outputs(1944) <= (inputs(182)) and not (inputs(190));
    layer0_outputs(1945) <= '0';
    layer0_outputs(1946) <= inputs(132);
    layer0_outputs(1947) <= not(inputs(156));
    layer0_outputs(1948) <= not((inputs(97)) and (inputs(154)));
    layer0_outputs(1949) <= not((inputs(53)) xor (inputs(92)));
    layer0_outputs(1950) <= (inputs(194)) xor (inputs(241));
    layer0_outputs(1951) <= inputs(237);
    layer0_outputs(1952) <= (inputs(120)) xor (inputs(25));
    layer0_outputs(1953) <= not((inputs(233)) xor (inputs(185)));
    layer0_outputs(1954) <= not(inputs(112));
    layer0_outputs(1955) <= (inputs(200)) and (inputs(165));
    layer0_outputs(1956) <= (inputs(103)) and not (inputs(77));
    layer0_outputs(1957) <= not(inputs(253)) or (inputs(43));
    layer0_outputs(1958) <= (inputs(36)) xor (inputs(126));
    layer0_outputs(1959) <= not(inputs(233));
    layer0_outputs(1960) <= inputs(44);
    layer0_outputs(1961) <= inputs(113);
    layer0_outputs(1962) <= not(inputs(90));
    layer0_outputs(1963) <= not(inputs(234)) or (inputs(172));
    layer0_outputs(1964) <= (inputs(151)) and not (inputs(3));
    layer0_outputs(1965) <= not(inputs(247));
    layer0_outputs(1966) <= not((inputs(222)) xor (inputs(6)));
    layer0_outputs(1967) <= (inputs(90)) or (inputs(60));
    layer0_outputs(1968) <= not((inputs(6)) or (inputs(166)));
    layer0_outputs(1969) <= (inputs(8)) xor (inputs(112));
    layer0_outputs(1970) <= not((inputs(62)) or (inputs(160)));
    layer0_outputs(1971) <= not(inputs(168));
    layer0_outputs(1972) <= inputs(229);
    layer0_outputs(1973) <= not((inputs(223)) xor (inputs(13)));
    layer0_outputs(1974) <= not(inputs(232));
    layer0_outputs(1975) <= (inputs(73)) and not (inputs(225));
    layer0_outputs(1976) <= (inputs(146)) xor (inputs(242));
    layer0_outputs(1977) <= (inputs(218)) or (inputs(4));
    layer0_outputs(1978) <= inputs(181);
    layer0_outputs(1979) <= not(inputs(176));
    layer0_outputs(1980) <= (inputs(211)) and not (inputs(105));
    layer0_outputs(1981) <= '0';
    layer0_outputs(1982) <= inputs(9);
    layer0_outputs(1983) <= not((inputs(90)) or (inputs(254)));
    layer0_outputs(1984) <= not((inputs(10)) or (inputs(224)));
    layer0_outputs(1985) <= (inputs(159)) and not (inputs(131));
    layer0_outputs(1986) <= (inputs(154)) or (inputs(140));
    layer0_outputs(1987) <= not(inputs(203));
    layer0_outputs(1988) <= (inputs(247)) or (inputs(97));
    layer0_outputs(1989) <= not(inputs(126));
    layer0_outputs(1990) <= (inputs(212)) or (inputs(205));
    layer0_outputs(1991) <= (inputs(159)) or (inputs(212));
    layer0_outputs(1992) <= not(inputs(24));
    layer0_outputs(1993) <= inputs(22);
    layer0_outputs(1994) <= not((inputs(88)) xor (inputs(139)));
    layer0_outputs(1995) <= not((inputs(250)) xor (inputs(156)));
    layer0_outputs(1996) <= not((inputs(246)) or (inputs(173)));
    layer0_outputs(1997) <= inputs(29);
    layer0_outputs(1998) <= (inputs(177)) and not (inputs(141));
    layer0_outputs(1999) <= (inputs(251)) xor (inputs(173));
    layer0_outputs(2000) <= not((inputs(96)) xor (inputs(108)));
    layer0_outputs(2001) <= not(inputs(90)) or (inputs(222));
    layer0_outputs(2002) <= inputs(143);
    layer0_outputs(2003) <= (inputs(126)) and not (inputs(190));
    layer0_outputs(2004) <= (inputs(25)) and not (inputs(162));
    layer0_outputs(2005) <= (inputs(192)) xor (inputs(206));
    layer0_outputs(2006) <= not(inputs(70)) or (inputs(18));
    layer0_outputs(2007) <= inputs(50);
    layer0_outputs(2008) <= not((inputs(137)) xor (inputs(58)));
    layer0_outputs(2009) <= (inputs(160)) xor (inputs(115));
    layer0_outputs(2010) <= not((inputs(7)) xor (inputs(59)));
    layer0_outputs(2011) <= not((inputs(146)) or (inputs(148)));
    layer0_outputs(2012) <= (inputs(49)) xor (inputs(101));
    layer0_outputs(2013) <= inputs(208);
    layer0_outputs(2014) <= (inputs(127)) and not (inputs(95));
    layer0_outputs(2015) <= not(inputs(156));
    layer0_outputs(2016) <= (inputs(225)) and not (inputs(15));
    layer0_outputs(2017) <= (inputs(213)) and not (inputs(174));
    layer0_outputs(2018) <= not(inputs(8)) or (inputs(126));
    layer0_outputs(2019) <= not(inputs(242));
    layer0_outputs(2020) <= not(inputs(218)) or (inputs(75));
    layer0_outputs(2021) <= (inputs(240)) and (inputs(134));
    layer0_outputs(2022) <= (inputs(156)) or (inputs(9));
    layer0_outputs(2023) <= not((inputs(140)) and (inputs(78)));
    layer0_outputs(2024) <= (inputs(16)) or (inputs(2));
    layer0_outputs(2025) <= (inputs(74)) or (inputs(108));
    layer0_outputs(2026) <= (inputs(173)) and not (inputs(95));
    layer0_outputs(2027) <= not(inputs(136)) or (inputs(205));
    layer0_outputs(2028) <= not((inputs(172)) xor (inputs(184)));
    layer0_outputs(2029) <= inputs(235);
    layer0_outputs(2030) <= not(inputs(244));
    layer0_outputs(2031) <= (inputs(243)) or (inputs(225));
    layer0_outputs(2032) <= (inputs(39)) or (inputs(116));
    layer0_outputs(2033) <= (inputs(101)) xor (inputs(69));
    layer0_outputs(2034) <= not(inputs(147));
    layer0_outputs(2035) <= (inputs(189)) and not (inputs(95));
    layer0_outputs(2036) <= inputs(221);
    layer0_outputs(2037) <= (inputs(234)) and not (inputs(91));
    layer0_outputs(2038) <= (inputs(194)) and not (inputs(223));
    layer0_outputs(2039) <= inputs(67);
    layer0_outputs(2040) <= (inputs(183)) and not (inputs(180));
    layer0_outputs(2041) <= not((inputs(161)) or (inputs(75)));
    layer0_outputs(2042) <= (inputs(85)) and not (inputs(223));
    layer0_outputs(2043) <= inputs(62);
    layer0_outputs(2044) <= (inputs(87)) xor (inputs(125));
    layer0_outputs(2045) <= not((inputs(236)) xor (inputs(195)));
    layer0_outputs(2046) <= not(inputs(158));
    layer0_outputs(2047) <= (inputs(43)) or (inputs(97));
    layer0_outputs(2048) <= not(inputs(122));
    layer0_outputs(2049) <= not(inputs(145));
    layer0_outputs(2050) <= not((inputs(130)) or (inputs(244)));
    layer0_outputs(2051) <= not(inputs(87));
    layer0_outputs(2052) <= not((inputs(201)) xor (inputs(221)));
    layer0_outputs(2053) <= (inputs(143)) and not (inputs(96));
    layer0_outputs(2054) <= (inputs(106)) and not (inputs(20));
    layer0_outputs(2055) <= (inputs(7)) and not (inputs(175));
    layer0_outputs(2056) <= inputs(59);
    layer0_outputs(2057) <= (inputs(137)) or (inputs(104));
    layer0_outputs(2058) <= inputs(30);
    layer0_outputs(2059) <= not(inputs(36)) or (inputs(143));
    layer0_outputs(2060) <= (inputs(106)) and not (inputs(204));
    layer0_outputs(2061) <= (inputs(91)) xor (inputs(245));
    layer0_outputs(2062) <= not(inputs(135));
    layer0_outputs(2063) <= inputs(150);
    layer0_outputs(2064) <= not(inputs(23));
    layer0_outputs(2065) <= (inputs(141)) or (inputs(57));
    layer0_outputs(2066) <= inputs(3);
    layer0_outputs(2067) <= not((inputs(168)) xor (inputs(232)));
    layer0_outputs(2068) <= not(inputs(9));
    layer0_outputs(2069) <= inputs(122);
    layer0_outputs(2070) <= not((inputs(58)) or (inputs(176)));
    layer0_outputs(2071) <= inputs(38);
    layer0_outputs(2072) <= inputs(23);
    layer0_outputs(2073) <= not(inputs(147));
    layer0_outputs(2074) <= not(inputs(68));
    layer0_outputs(2075) <= not(inputs(180)) or (inputs(79));
    layer0_outputs(2076) <= inputs(247);
    layer0_outputs(2077) <= inputs(109);
    layer0_outputs(2078) <= not(inputs(233)) or (inputs(86));
    layer0_outputs(2079) <= (inputs(158)) and not (inputs(48));
    layer0_outputs(2080) <= (inputs(222)) or (inputs(31));
    layer0_outputs(2081) <= (inputs(132)) xor (inputs(122));
    layer0_outputs(2082) <= not(inputs(235));
    layer0_outputs(2083) <= (inputs(134)) and not (inputs(17));
    layer0_outputs(2084) <= (inputs(66)) or (inputs(93));
    layer0_outputs(2085) <= inputs(225);
    layer0_outputs(2086) <= not(inputs(176)) or (inputs(95));
    layer0_outputs(2087) <= not(inputs(137));
    layer0_outputs(2088) <= not((inputs(17)) xor (inputs(30)));
    layer0_outputs(2089) <= inputs(20);
    layer0_outputs(2090) <= not(inputs(230));
    layer0_outputs(2091) <= (inputs(124)) or (inputs(68));
    layer0_outputs(2092) <= not((inputs(206)) and (inputs(241)));
    layer0_outputs(2093) <= not((inputs(68)) xor (inputs(195)));
    layer0_outputs(2094) <= not((inputs(14)) or (inputs(115)));
    layer0_outputs(2095) <= not(inputs(6));
    layer0_outputs(2096) <= (inputs(98)) xor (inputs(218));
    layer0_outputs(2097) <= (inputs(101)) and not (inputs(207));
    layer0_outputs(2098) <= (inputs(49)) or (inputs(93));
    layer0_outputs(2099) <= not((inputs(124)) xor (inputs(117)));
    layer0_outputs(2100) <= not(inputs(181)) or (inputs(240));
    layer0_outputs(2101) <= (inputs(147)) xor (inputs(85));
    layer0_outputs(2102) <= inputs(118);
    layer0_outputs(2103) <= not(inputs(107));
    layer0_outputs(2104) <= (inputs(255)) or (inputs(204));
    layer0_outputs(2105) <= not((inputs(155)) or (inputs(162)));
    layer0_outputs(2106) <= (inputs(211)) or (inputs(71));
    layer0_outputs(2107) <= '0';
    layer0_outputs(2108) <= (inputs(15)) and (inputs(153));
    layer0_outputs(2109) <= not((inputs(210)) or (inputs(41)));
    layer0_outputs(2110) <= inputs(150);
    layer0_outputs(2111) <= (inputs(189)) and not (inputs(83));
    layer0_outputs(2112) <= (inputs(84)) and not (inputs(42));
    layer0_outputs(2113) <= not(inputs(7));
    layer0_outputs(2114) <= (inputs(63)) or (inputs(201));
    layer0_outputs(2115) <= not(inputs(166));
    layer0_outputs(2116) <= not((inputs(121)) xor (inputs(162)));
    layer0_outputs(2117) <= (inputs(197)) and not (inputs(124));
    layer0_outputs(2118) <= inputs(147);
    layer0_outputs(2119) <= not(inputs(127)) or (inputs(152));
    layer0_outputs(2120) <= not((inputs(159)) xor (inputs(1)));
    layer0_outputs(2121) <= inputs(101);
    layer0_outputs(2122) <= (inputs(120)) and not (inputs(76));
    layer0_outputs(2123) <= inputs(3);
    layer0_outputs(2124) <= (inputs(165)) and not (inputs(223));
    layer0_outputs(2125) <= not(inputs(194));
    layer0_outputs(2126) <= not(inputs(120));
    layer0_outputs(2127) <= not(inputs(213));
    layer0_outputs(2128) <= not(inputs(98));
    layer0_outputs(2129) <= not(inputs(116));
    layer0_outputs(2130) <= not(inputs(182));
    layer0_outputs(2131) <= not((inputs(198)) or (inputs(3)));
    layer0_outputs(2132) <= inputs(247);
    layer0_outputs(2133) <= inputs(192);
    layer0_outputs(2134) <= not(inputs(114)) or (inputs(172));
    layer0_outputs(2135) <= (inputs(71)) and not (inputs(150));
    layer0_outputs(2136) <= not(inputs(229));
    layer0_outputs(2137) <= (inputs(233)) or (inputs(187));
    layer0_outputs(2138) <= not((inputs(66)) or (inputs(184)));
    layer0_outputs(2139) <= inputs(13);
    layer0_outputs(2140) <= not(inputs(231));
    layer0_outputs(2141) <= (inputs(67)) xor (inputs(24));
    layer0_outputs(2142) <= (inputs(172)) and not (inputs(64));
    layer0_outputs(2143) <= not(inputs(92)) or (inputs(159));
    layer0_outputs(2144) <= inputs(210);
    layer0_outputs(2145) <= not(inputs(135));
    layer0_outputs(2146) <= not((inputs(90)) xor (inputs(206)));
    layer0_outputs(2147) <= not(inputs(105));
    layer0_outputs(2148) <= (inputs(151)) or (inputs(98));
    layer0_outputs(2149) <= not((inputs(89)) or (inputs(148)));
    layer0_outputs(2150) <= inputs(228);
    layer0_outputs(2151) <= (inputs(250)) or (inputs(44));
    layer0_outputs(2152) <= (inputs(23)) and not (inputs(196));
    layer0_outputs(2153) <= (inputs(86)) xor (inputs(154));
    layer0_outputs(2154) <= not(inputs(150)) or (inputs(14));
    layer0_outputs(2155) <= not((inputs(76)) or (inputs(140)));
    layer0_outputs(2156) <= not((inputs(28)) or (inputs(96)));
    layer0_outputs(2157) <= not(inputs(167));
    layer0_outputs(2158) <= not(inputs(119));
    layer0_outputs(2159) <= (inputs(96)) or (inputs(246));
    layer0_outputs(2160) <= inputs(139);
    layer0_outputs(2161) <= inputs(233);
    layer0_outputs(2162) <= not(inputs(214)) or (inputs(162));
    layer0_outputs(2163) <= (inputs(153)) or (inputs(151));
    layer0_outputs(2164) <= (inputs(167)) and not (inputs(255));
    layer0_outputs(2165) <= not(inputs(59));
    layer0_outputs(2166) <= (inputs(123)) or (inputs(140));
    layer0_outputs(2167) <= not(inputs(207));
    layer0_outputs(2168) <= (inputs(233)) and not (inputs(62));
    layer0_outputs(2169) <= (inputs(216)) and not (inputs(104));
    layer0_outputs(2170) <= not((inputs(165)) or (inputs(166)));
    layer0_outputs(2171) <= inputs(239);
    layer0_outputs(2172) <= inputs(39);
    layer0_outputs(2173) <= not((inputs(53)) or (inputs(8)));
    layer0_outputs(2174) <= (inputs(202)) or (inputs(11));
    layer0_outputs(2175) <= (inputs(26)) and not (inputs(213));
    layer0_outputs(2176) <= not(inputs(119));
    layer0_outputs(2177) <= '0';
    layer0_outputs(2178) <= inputs(190);
    layer0_outputs(2179) <= (inputs(104)) and not (inputs(155));
    layer0_outputs(2180) <= not(inputs(101)) or (inputs(160));
    layer0_outputs(2181) <= not(inputs(22));
    layer0_outputs(2182) <= not(inputs(248)) or (inputs(77));
    layer0_outputs(2183) <= not(inputs(44));
    layer0_outputs(2184) <= not(inputs(221));
    layer0_outputs(2185) <= not(inputs(216)) or (inputs(69));
    layer0_outputs(2186) <= inputs(232);
    layer0_outputs(2187) <= not(inputs(4)) or (inputs(218));
    layer0_outputs(2188) <= inputs(134);
    layer0_outputs(2189) <= (inputs(166)) and not (inputs(191));
    layer0_outputs(2190) <= (inputs(132)) xor (inputs(102));
    layer0_outputs(2191) <= not((inputs(215)) xor (inputs(199)));
    layer0_outputs(2192) <= not((inputs(29)) xor (inputs(132)));
    layer0_outputs(2193) <= not(inputs(71)) or (inputs(46));
    layer0_outputs(2194) <= not(inputs(236)) or (inputs(81));
    layer0_outputs(2195) <= not((inputs(39)) and (inputs(112)));
    layer0_outputs(2196) <= (inputs(234)) and not (inputs(123));
    layer0_outputs(2197) <= not((inputs(117)) or (inputs(83)));
    layer0_outputs(2198) <= (inputs(37)) and not (inputs(124));
    layer0_outputs(2199) <= not((inputs(175)) or (inputs(198)));
    layer0_outputs(2200) <= (inputs(147)) or (inputs(163));
    layer0_outputs(2201) <= '1';
    layer0_outputs(2202) <= inputs(62);
    layer0_outputs(2203) <= not(inputs(254));
    layer0_outputs(2204) <= (inputs(30)) or (inputs(26));
    layer0_outputs(2205) <= not(inputs(231)) or (inputs(63));
    layer0_outputs(2206) <= inputs(86);
    layer0_outputs(2207) <= (inputs(119)) and not (inputs(52));
    layer0_outputs(2208) <= inputs(230);
    layer0_outputs(2209) <= not(inputs(229));
    layer0_outputs(2210) <= inputs(144);
    layer0_outputs(2211) <= not((inputs(91)) xor (inputs(108)));
    layer0_outputs(2212) <= (inputs(90)) and not (inputs(116));
    layer0_outputs(2213) <= not(inputs(38));
    layer0_outputs(2214) <= not((inputs(158)) or (inputs(129)));
    layer0_outputs(2215) <= (inputs(40)) or (inputs(32));
    layer0_outputs(2216) <= (inputs(177)) and not (inputs(48));
    layer0_outputs(2217) <= inputs(59);
    layer0_outputs(2218) <= (inputs(180)) or (inputs(236));
    layer0_outputs(2219) <= (inputs(85)) and (inputs(225));
    layer0_outputs(2220) <= (inputs(198)) and not (inputs(123));
    layer0_outputs(2221) <= '1';
    layer0_outputs(2222) <= inputs(25);
    layer0_outputs(2223) <= not((inputs(107)) or (inputs(33)));
    layer0_outputs(2224) <= '1';
    layer0_outputs(2225) <= (inputs(148)) and not (inputs(108));
    layer0_outputs(2226) <= inputs(188);
    layer0_outputs(2227) <= (inputs(209)) and not (inputs(15));
    layer0_outputs(2228) <= (inputs(169)) or (inputs(127));
    layer0_outputs(2229) <= (inputs(184)) or (inputs(82));
    layer0_outputs(2230) <= (inputs(136)) or (inputs(91));
    layer0_outputs(2231) <= not(inputs(166));
    layer0_outputs(2232) <= (inputs(190)) or (inputs(198));
    layer0_outputs(2233) <= (inputs(68)) and not (inputs(175));
    layer0_outputs(2234) <= not(inputs(233));
    layer0_outputs(2235) <= (inputs(254)) or (inputs(151));
    layer0_outputs(2236) <= not(inputs(248)) or (inputs(64));
    layer0_outputs(2237) <= not(inputs(152)) or (inputs(27));
    layer0_outputs(2238) <= not((inputs(139)) xor (inputs(24)));
    layer0_outputs(2239) <= not(inputs(101));
    layer0_outputs(2240) <= not(inputs(124));
    layer0_outputs(2241) <= (inputs(162)) and not (inputs(56));
    layer0_outputs(2242) <= inputs(200);
    layer0_outputs(2243) <= inputs(6);
    layer0_outputs(2244) <= (inputs(219)) and not (inputs(82));
    layer0_outputs(2245) <= (inputs(133)) and (inputs(246));
    layer0_outputs(2246) <= not(inputs(85));
    layer0_outputs(2247) <= not(inputs(162));
    layer0_outputs(2248) <= (inputs(77)) or (inputs(191));
    layer0_outputs(2249) <= inputs(103);
    layer0_outputs(2250) <= not((inputs(147)) xor (inputs(177)));
    layer0_outputs(2251) <= not((inputs(189)) or (inputs(221)));
    layer0_outputs(2252) <= not((inputs(51)) or (inputs(114)));
    layer0_outputs(2253) <= not((inputs(100)) or (inputs(127)));
    layer0_outputs(2254) <= not(inputs(146)) or (inputs(186));
    layer0_outputs(2255) <= inputs(223);
    layer0_outputs(2256) <= inputs(43);
    layer0_outputs(2257) <= not(inputs(233)) or (inputs(10));
    layer0_outputs(2258) <= (inputs(50)) and not (inputs(81));
    layer0_outputs(2259) <= (inputs(48)) xor (inputs(203));
    layer0_outputs(2260) <= (inputs(36)) or (inputs(132));
    layer0_outputs(2261) <= not((inputs(79)) xor (inputs(178)));
    layer0_outputs(2262) <= '0';
    layer0_outputs(2263) <= (inputs(77)) and not (inputs(2));
    layer0_outputs(2264) <= not(inputs(188)) or (inputs(93));
    layer0_outputs(2265) <= (inputs(117)) xor (inputs(69));
    layer0_outputs(2266) <= '1';
    layer0_outputs(2267) <= (inputs(157)) or (inputs(87));
    layer0_outputs(2268) <= (inputs(51)) and not (inputs(132));
    layer0_outputs(2269) <= not((inputs(157)) or (inputs(242)));
    layer0_outputs(2270) <= not(inputs(163));
    layer0_outputs(2271) <= inputs(198);
    layer0_outputs(2272) <= not((inputs(109)) xor (inputs(181)));
    layer0_outputs(2273) <= (inputs(238)) and not (inputs(224));
    layer0_outputs(2274) <= not((inputs(124)) or (inputs(148)));
    layer0_outputs(2275) <= (inputs(87)) and not (inputs(177));
    layer0_outputs(2276) <= not(inputs(174));
    layer0_outputs(2277) <= inputs(238);
    layer0_outputs(2278) <= not((inputs(61)) xor (inputs(23)));
    layer0_outputs(2279) <= (inputs(111)) xor (inputs(230));
    layer0_outputs(2280) <= not(inputs(188)) or (inputs(12));
    layer0_outputs(2281) <= not(inputs(101)) or (inputs(3));
    layer0_outputs(2282) <= not((inputs(78)) or (inputs(191)));
    layer0_outputs(2283) <= '1';
    layer0_outputs(2284) <= (inputs(5)) xor (inputs(159));
    layer0_outputs(2285) <= (inputs(104)) and not (inputs(164));
    layer0_outputs(2286) <= not(inputs(102));
    layer0_outputs(2287) <= not(inputs(218)) or (inputs(12));
    layer0_outputs(2288) <= inputs(77);
    layer0_outputs(2289) <= (inputs(140)) xor (inputs(164));
    layer0_outputs(2290) <= (inputs(88)) and not (inputs(157));
    layer0_outputs(2291) <= (inputs(0)) and (inputs(34));
    layer0_outputs(2292) <= (inputs(157)) and not (inputs(153));
    layer0_outputs(2293) <= not(inputs(226));
    layer0_outputs(2294) <= (inputs(83)) xor (inputs(169));
    layer0_outputs(2295) <= not(inputs(72)) or (inputs(151));
    layer0_outputs(2296) <= '1';
    layer0_outputs(2297) <= not(inputs(169)) or (inputs(12));
    layer0_outputs(2298) <= (inputs(139)) and not (inputs(34));
    layer0_outputs(2299) <= '0';
    layer0_outputs(2300) <= not(inputs(134)) or (inputs(108));
    layer0_outputs(2301) <= inputs(214);
    layer0_outputs(2302) <= inputs(185);
    layer0_outputs(2303) <= (inputs(122)) xor (inputs(158));
    layer0_outputs(2304) <= not((inputs(88)) or (inputs(252)));
    layer0_outputs(2305) <= not(inputs(231));
    layer0_outputs(2306) <= inputs(103);
    layer0_outputs(2307) <= (inputs(246)) xor (inputs(112));
    layer0_outputs(2308) <= not((inputs(2)) or (inputs(32)));
    layer0_outputs(2309) <= not(inputs(0));
    layer0_outputs(2310) <= (inputs(155)) and not (inputs(5));
    layer0_outputs(2311) <= (inputs(109)) and not (inputs(115));
    layer0_outputs(2312) <= inputs(18);
    layer0_outputs(2313) <= not(inputs(48));
    layer0_outputs(2314) <= (inputs(181)) and not (inputs(162));
    layer0_outputs(2315) <= not(inputs(152));
    layer0_outputs(2316) <= (inputs(172)) or (inputs(251));
    layer0_outputs(2317) <= not((inputs(147)) xor (inputs(190)));
    layer0_outputs(2318) <= inputs(232);
    layer0_outputs(2319) <= not((inputs(235)) or (inputs(37)));
    layer0_outputs(2320) <= not((inputs(144)) xor (inputs(211)));
    layer0_outputs(2321) <= not((inputs(241)) or (inputs(249)));
    layer0_outputs(2322) <= (inputs(100)) and not (inputs(224));
    layer0_outputs(2323) <= inputs(217);
    layer0_outputs(2324) <= '1';
    layer0_outputs(2325) <= not((inputs(168)) or (inputs(1)));
    layer0_outputs(2326) <= (inputs(1)) and (inputs(15));
    layer0_outputs(2327) <= not((inputs(29)) or (inputs(15)));
    layer0_outputs(2328) <= not((inputs(99)) or (inputs(165)));
    layer0_outputs(2329) <= inputs(180);
    layer0_outputs(2330) <= not(inputs(103)) or (inputs(179));
    layer0_outputs(2331) <= not(inputs(108));
    layer0_outputs(2332) <= inputs(132);
    layer0_outputs(2333) <= not((inputs(192)) or (inputs(6)));
    layer0_outputs(2334) <= not(inputs(119));
    layer0_outputs(2335) <= (inputs(172)) xor (inputs(221));
    layer0_outputs(2336) <= (inputs(113)) or (inputs(99));
    layer0_outputs(2337) <= not(inputs(211));
    layer0_outputs(2338) <= not(inputs(212));
    layer0_outputs(2339) <= (inputs(104)) and not (inputs(206));
    layer0_outputs(2340) <= not((inputs(235)) and (inputs(218)));
    layer0_outputs(2341) <= not((inputs(209)) or (inputs(5)));
    layer0_outputs(2342) <= (inputs(154)) and not (inputs(250));
    layer0_outputs(2343) <= (inputs(138)) xor (inputs(13));
    layer0_outputs(2344) <= (inputs(196)) or (inputs(252));
    layer0_outputs(2345) <= not(inputs(231));
    layer0_outputs(2346) <= (inputs(206)) and (inputs(183));
    layer0_outputs(2347) <= not((inputs(157)) and (inputs(77)));
    layer0_outputs(2348) <= (inputs(34)) xor (inputs(168));
    layer0_outputs(2349) <= not(inputs(197));
    layer0_outputs(2350) <= not(inputs(184));
    layer0_outputs(2351) <= (inputs(138)) xor (inputs(136));
    layer0_outputs(2352) <= not((inputs(223)) or (inputs(41)));
    layer0_outputs(2353) <= inputs(40);
    layer0_outputs(2354) <= (inputs(135)) or (inputs(134));
    layer0_outputs(2355) <= (inputs(142)) and (inputs(236));
    layer0_outputs(2356) <= not((inputs(70)) xor (inputs(109)));
    layer0_outputs(2357) <= (inputs(149)) and not (inputs(80));
    layer0_outputs(2358) <= inputs(195);
    layer0_outputs(2359) <= not((inputs(161)) or (inputs(212)));
    layer0_outputs(2360) <= (inputs(61)) xor (inputs(23));
    layer0_outputs(2361) <= not((inputs(249)) xor (inputs(102)));
    layer0_outputs(2362) <= not(inputs(108));
    layer0_outputs(2363) <= not(inputs(181)) or (inputs(171));
    layer0_outputs(2364) <= not((inputs(156)) xor (inputs(8)));
    layer0_outputs(2365) <= inputs(57);
    layer0_outputs(2366) <= not((inputs(79)) or (inputs(23)));
    layer0_outputs(2367) <= not((inputs(59)) and (inputs(106)));
    layer0_outputs(2368) <= not(inputs(34)) or (inputs(77));
    layer0_outputs(2369) <= not((inputs(189)) xor (inputs(27)));
    layer0_outputs(2370) <= inputs(34);
    layer0_outputs(2371) <= not((inputs(229)) or (inputs(33)));
    layer0_outputs(2372) <= (inputs(100)) and not (inputs(110));
    layer0_outputs(2373) <= (inputs(220)) or (inputs(212));
    layer0_outputs(2374) <= not(inputs(210));
    layer0_outputs(2375) <= (inputs(29)) and not (inputs(189));
    layer0_outputs(2376) <= inputs(149);
    layer0_outputs(2377) <= inputs(27);
    layer0_outputs(2378) <= not(inputs(41));
    layer0_outputs(2379) <= (inputs(68)) and not (inputs(17));
    layer0_outputs(2380) <= not(inputs(93)) or (inputs(181));
    layer0_outputs(2381) <= not(inputs(75)) or (inputs(255));
    layer0_outputs(2382) <= (inputs(102)) xor (inputs(148));
    layer0_outputs(2383) <= not(inputs(148));
    layer0_outputs(2384) <= not(inputs(241));
    layer0_outputs(2385) <= (inputs(246)) or (inputs(249));
    layer0_outputs(2386) <= not((inputs(63)) xor (inputs(16)));
    layer0_outputs(2387) <= not(inputs(152)) or (inputs(216));
    layer0_outputs(2388) <= (inputs(218)) or (inputs(207));
    layer0_outputs(2389) <= not((inputs(54)) and (inputs(37)));
    layer0_outputs(2390) <= inputs(118);
    layer0_outputs(2391) <= inputs(91);
    layer0_outputs(2392) <= not(inputs(253));
    layer0_outputs(2393) <= not((inputs(32)) xor (inputs(14)));
    layer0_outputs(2394) <= inputs(128);
    layer0_outputs(2395) <= not(inputs(251));
    layer0_outputs(2396) <= not(inputs(24));
    layer0_outputs(2397) <= not(inputs(244)) or (inputs(4));
    layer0_outputs(2398) <= not(inputs(99));
    layer0_outputs(2399) <= (inputs(160)) and not (inputs(254));
    layer0_outputs(2400) <= inputs(219);
    layer0_outputs(2401) <= not((inputs(32)) and (inputs(240)));
    layer0_outputs(2402) <= inputs(131);
    layer0_outputs(2403) <= not((inputs(216)) or (inputs(201)));
    layer0_outputs(2404) <= (inputs(107)) and not (inputs(255));
    layer0_outputs(2405) <= inputs(77);
    layer0_outputs(2406) <= not(inputs(106));
    layer0_outputs(2407) <= (inputs(46)) and (inputs(107));
    layer0_outputs(2408) <= not(inputs(148)) or (inputs(34));
    layer0_outputs(2409) <= not((inputs(82)) xor (inputs(182)));
    layer0_outputs(2410) <= not(inputs(30)) or (inputs(206));
    layer0_outputs(2411) <= (inputs(44)) and (inputs(191));
    layer0_outputs(2412) <= inputs(210);
    layer0_outputs(2413) <= not(inputs(106));
    layer0_outputs(2414) <= not(inputs(88)) or (inputs(143));
    layer0_outputs(2415) <= (inputs(232)) and (inputs(164));
    layer0_outputs(2416) <= not((inputs(25)) or (inputs(189)));
    layer0_outputs(2417) <= inputs(191);
    layer0_outputs(2418) <= inputs(40);
    layer0_outputs(2419) <= inputs(41);
    layer0_outputs(2420) <= not((inputs(232)) xor (inputs(155)));
    layer0_outputs(2421) <= not(inputs(105));
    layer0_outputs(2422) <= not(inputs(216));
    layer0_outputs(2423) <= (inputs(39)) and not (inputs(157));
    layer0_outputs(2424) <= (inputs(85)) and (inputs(88));
    layer0_outputs(2425) <= (inputs(93)) or (inputs(126));
    layer0_outputs(2426) <= (inputs(212)) or (inputs(65));
    layer0_outputs(2427) <= (inputs(41)) xor (inputs(80));
    layer0_outputs(2428) <= (inputs(51)) and not (inputs(54));
    layer0_outputs(2429) <= not((inputs(62)) xor (inputs(228)));
    layer0_outputs(2430) <= (inputs(205)) or (inputs(228));
    layer0_outputs(2431) <= not(inputs(182)) or (inputs(71));
    layer0_outputs(2432) <= '0';
    layer0_outputs(2433) <= (inputs(74)) and (inputs(33));
    layer0_outputs(2434) <= inputs(239);
    layer0_outputs(2435) <= (inputs(115)) xor (inputs(129));
    layer0_outputs(2436) <= (inputs(77)) and not (inputs(132));
    layer0_outputs(2437) <= not(inputs(246));
    layer0_outputs(2438) <= inputs(19);
    layer0_outputs(2439) <= '1';
    layer0_outputs(2440) <= inputs(103);
    layer0_outputs(2441) <= (inputs(116)) and not (inputs(178));
    layer0_outputs(2442) <= inputs(158);
    layer0_outputs(2443) <= not(inputs(115)) or (inputs(180));
    layer0_outputs(2444) <= (inputs(183)) xor (inputs(54));
    layer0_outputs(2445) <= not(inputs(96));
    layer0_outputs(2446) <= not((inputs(175)) xor (inputs(219)));
    layer0_outputs(2447) <= inputs(85);
    layer0_outputs(2448) <= (inputs(12)) or (inputs(34));
    layer0_outputs(2449) <= (inputs(160)) or (inputs(208));
    layer0_outputs(2450) <= (inputs(170)) or (inputs(144));
    layer0_outputs(2451) <= inputs(174);
    layer0_outputs(2452) <= not((inputs(252)) xor (inputs(147)));
    layer0_outputs(2453) <= (inputs(163)) or (inputs(93));
    layer0_outputs(2454) <= (inputs(96)) xor (inputs(30));
    layer0_outputs(2455) <= (inputs(43)) xor (inputs(28));
    layer0_outputs(2456) <= inputs(139);
    layer0_outputs(2457) <= '0';
    layer0_outputs(2458) <= inputs(44);
    layer0_outputs(2459) <= not(inputs(167));
    layer0_outputs(2460) <= (inputs(156)) xor (inputs(123));
    layer0_outputs(2461) <= not(inputs(234));
    layer0_outputs(2462) <= (inputs(114)) xor (inputs(149));
    layer0_outputs(2463) <= not(inputs(104));
    layer0_outputs(2464) <= not((inputs(189)) or (inputs(174)));
    layer0_outputs(2465) <= (inputs(16)) and (inputs(239));
    layer0_outputs(2466) <= (inputs(245)) and not (inputs(49));
    layer0_outputs(2467) <= not(inputs(136));
    layer0_outputs(2468) <= not(inputs(202)) or (inputs(70));
    layer0_outputs(2469) <= not(inputs(153)) or (inputs(65));
    layer0_outputs(2470) <= not(inputs(90)) or (inputs(61));
    layer0_outputs(2471) <= not(inputs(73)) or (inputs(158));
    layer0_outputs(2472) <= not(inputs(215));
    layer0_outputs(2473) <= not(inputs(54));
    layer0_outputs(2474) <= inputs(68);
    layer0_outputs(2475) <= not(inputs(193));
    layer0_outputs(2476) <= (inputs(104)) or (inputs(130));
    layer0_outputs(2477) <= inputs(36);
    layer0_outputs(2478) <= (inputs(123)) and not (inputs(182));
    layer0_outputs(2479) <= not(inputs(186)) or (inputs(33));
    layer0_outputs(2480) <= not(inputs(252)) or (inputs(205));
    layer0_outputs(2481) <= not(inputs(172));
    layer0_outputs(2482) <= inputs(215);
    layer0_outputs(2483) <= (inputs(219)) xor (inputs(155));
    layer0_outputs(2484) <= not((inputs(123)) and (inputs(249)));
    layer0_outputs(2485) <= (inputs(89)) xor (inputs(75));
    layer0_outputs(2486) <= not((inputs(221)) or (inputs(239)));
    layer0_outputs(2487) <= (inputs(181)) and not (inputs(130));
    layer0_outputs(2488) <= (inputs(237)) xor (inputs(116));
    layer0_outputs(2489) <= inputs(90);
    layer0_outputs(2490) <= (inputs(47)) or (inputs(61));
    layer0_outputs(2491) <= not(inputs(40));
    layer0_outputs(2492) <= (inputs(106)) and (inputs(10));
    layer0_outputs(2493) <= not((inputs(99)) or (inputs(95)));
    layer0_outputs(2494) <= (inputs(79)) or (inputs(191));
    layer0_outputs(2495) <= '1';
    layer0_outputs(2496) <= (inputs(61)) xor (inputs(243));
    layer0_outputs(2497) <= inputs(73);
    layer0_outputs(2498) <= (inputs(159)) or (inputs(112));
    layer0_outputs(2499) <= not((inputs(48)) or (inputs(194)));
    layer0_outputs(2500) <= (inputs(177)) or (inputs(204));
    layer0_outputs(2501) <= (inputs(176)) and (inputs(64));
    layer0_outputs(2502) <= not(inputs(116));
    layer0_outputs(2503) <= not((inputs(253)) or (inputs(153)));
    layer0_outputs(2504) <= '1';
    layer0_outputs(2505) <= inputs(230);
    layer0_outputs(2506) <= inputs(239);
    layer0_outputs(2507) <= not((inputs(218)) or (inputs(221)));
    layer0_outputs(2508) <= not(inputs(66)) or (inputs(172));
    layer0_outputs(2509) <= inputs(213);
    layer0_outputs(2510) <= not((inputs(11)) or (inputs(26)));
    layer0_outputs(2511) <= inputs(6);
    layer0_outputs(2512) <= not((inputs(217)) xor (inputs(201)));
    layer0_outputs(2513) <= (inputs(92)) and not (inputs(226));
    layer0_outputs(2514) <= not((inputs(157)) xor (inputs(101)));
    layer0_outputs(2515) <= not((inputs(88)) or (inputs(105)));
    layer0_outputs(2516) <= not((inputs(220)) or (inputs(231)));
    layer0_outputs(2517) <= not(inputs(77)) or (inputs(199));
    layer0_outputs(2518) <= not((inputs(247)) or (inputs(65)));
    layer0_outputs(2519) <= (inputs(171)) or (inputs(223));
    layer0_outputs(2520) <= (inputs(149)) or (inputs(18));
    layer0_outputs(2521) <= not((inputs(111)) xor (inputs(207)));
    layer0_outputs(2522) <= inputs(249);
    layer0_outputs(2523) <= (inputs(43)) or (inputs(164));
    layer0_outputs(2524) <= (inputs(121)) and not (inputs(223));
    layer0_outputs(2525) <= not(inputs(9));
    layer0_outputs(2526) <= not(inputs(188)) or (inputs(107));
    layer0_outputs(2527) <= not((inputs(35)) or (inputs(20)));
    layer0_outputs(2528) <= not(inputs(12));
    layer0_outputs(2529) <= not(inputs(96));
    layer0_outputs(2530) <= '0';
    layer0_outputs(2531) <= not(inputs(214)) or (inputs(21));
    layer0_outputs(2532) <= inputs(170);
    layer0_outputs(2533) <= not(inputs(92)) or (inputs(215));
    layer0_outputs(2534) <= not(inputs(169)) or (inputs(17));
    layer0_outputs(2535) <= (inputs(41)) and (inputs(43));
    layer0_outputs(2536) <= (inputs(216)) and not (inputs(54));
    layer0_outputs(2537) <= '0';
    layer0_outputs(2538) <= not(inputs(35)) or (inputs(112));
    layer0_outputs(2539) <= (inputs(252)) or (inputs(138));
    layer0_outputs(2540) <= inputs(215);
    layer0_outputs(2541) <= not((inputs(31)) or (inputs(154)));
    layer0_outputs(2542) <= not(inputs(63));
    layer0_outputs(2543) <= (inputs(210)) and not (inputs(31));
    layer0_outputs(2544) <= not(inputs(20)) or (inputs(176));
    layer0_outputs(2545) <= (inputs(131)) and (inputs(39));
    layer0_outputs(2546) <= (inputs(108)) or (inputs(100));
    layer0_outputs(2547) <= not(inputs(123));
    layer0_outputs(2548) <= inputs(36);
    layer0_outputs(2549) <= not((inputs(130)) or (inputs(190)));
    layer0_outputs(2550) <= (inputs(97)) xor (inputs(193));
    layer0_outputs(2551) <= (inputs(59)) and not (inputs(59));
    layer0_outputs(2552) <= not((inputs(76)) or (inputs(173)));
    layer0_outputs(2553) <= not(inputs(29));
    layer0_outputs(2554) <= not((inputs(97)) or (inputs(228)));
    layer0_outputs(2555) <= not((inputs(15)) and (inputs(238)));
    layer0_outputs(2556) <= not(inputs(230)) or (inputs(123));
    layer0_outputs(2557) <= inputs(77);
    layer0_outputs(2558) <= '1';
    layer0_outputs(2559) <= (inputs(156)) or (inputs(127));
    layer0_outputs(2560) <= (inputs(205)) or (inputs(95));
    layer0_outputs(2561) <= '1';
    layer0_outputs(2562) <= inputs(7);
    layer0_outputs(2563) <= (inputs(207)) or (inputs(136));
    layer0_outputs(2564) <= not(inputs(61)) or (inputs(0));
    layer0_outputs(2565) <= not((inputs(81)) or (inputs(62)));
    layer0_outputs(2566) <= not((inputs(194)) xor (inputs(24)));
    layer0_outputs(2567) <= (inputs(70)) and not (inputs(205));
    layer0_outputs(2568) <= inputs(38);
    layer0_outputs(2569) <= (inputs(60)) or (inputs(40));
    layer0_outputs(2570) <= (inputs(5)) xor (inputs(64));
    layer0_outputs(2571) <= (inputs(48)) xor (inputs(103));
    layer0_outputs(2572) <= inputs(142);
    layer0_outputs(2573) <= not(inputs(23));
    layer0_outputs(2574) <= not(inputs(109));
    layer0_outputs(2575) <= inputs(18);
    layer0_outputs(2576) <= not(inputs(153));
    layer0_outputs(2577) <= inputs(51);
    layer0_outputs(2578) <= inputs(99);
    layer0_outputs(2579) <= not((inputs(245)) or (inputs(221)));
    layer0_outputs(2580) <= not((inputs(41)) or (inputs(225)));
    layer0_outputs(2581) <= not(inputs(137)) or (inputs(198));
    layer0_outputs(2582) <= not((inputs(142)) xor (inputs(162)));
    layer0_outputs(2583) <= not(inputs(16));
    layer0_outputs(2584) <= (inputs(253)) and not (inputs(31));
    layer0_outputs(2585) <= not(inputs(247));
    layer0_outputs(2586) <= not((inputs(39)) xor (inputs(223)));
    layer0_outputs(2587) <= (inputs(235)) xor (inputs(211));
    layer0_outputs(2588) <= not(inputs(74));
    layer0_outputs(2589) <= (inputs(105)) xor (inputs(163));
    layer0_outputs(2590) <= not(inputs(38)) or (inputs(114));
    layer0_outputs(2591) <= (inputs(78)) xor (inputs(171));
    layer0_outputs(2592) <= inputs(153);
    layer0_outputs(2593) <= (inputs(67)) or (inputs(209));
    layer0_outputs(2594) <= not((inputs(131)) or (inputs(198)));
    layer0_outputs(2595) <= (inputs(218)) xor (inputs(182));
    layer0_outputs(2596) <= (inputs(157)) xor (inputs(124));
    layer0_outputs(2597) <= not(inputs(30)) or (inputs(93));
    layer0_outputs(2598) <= inputs(197);
    layer0_outputs(2599) <= not(inputs(193));
    layer0_outputs(2600) <= not((inputs(3)) or (inputs(125)));
    layer0_outputs(2601) <= not(inputs(109));
    layer0_outputs(2602) <= (inputs(151)) or (inputs(81));
    layer0_outputs(2603) <= not(inputs(146));
    layer0_outputs(2604) <= (inputs(199)) and not (inputs(10));
    layer0_outputs(2605) <= not((inputs(148)) xor (inputs(54)));
    layer0_outputs(2606) <= not((inputs(96)) xor (inputs(54)));
    layer0_outputs(2607) <= not((inputs(200)) or (inputs(3)));
    layer0_outputs(2608) <= inputs(179);
    layer0_outputs(2609) <= not(inputs(73));
    layer0_outputs(2610) <= (inputs(148)) xor (inputs(195));
    layer0_outputs(2611) <= not((inputs(169)) and (inputs(210)));
    layer0_outputs(2612) <= (inputs(158)) xor (inputs(159));
    layer0_outputs(2613) <= not((inputs(195)) or (inputs(76)));
    layer0_outputs(2614) <= not(inputs(87));
    layer0_outputs(2615) <= (inputs(241)) or (inputs(227));
    layer0_outputs(2616) <= (inputs(27)) or (inputs(202));
    layer0_outputs(2617) <= not((inputs(247)) or (inputs(250)));
    layer0_outputs(2618) <= not((inputs(231)) xor (inputs(42)));
    layer0_outputs(2619) <= not(inputs(83)) or (inputs(191));
    layer0_outputs(2620) <= (inputs(160)) xor (inputs(37));
    layer0_outputs(2621) <= (inputs(15)) or (inputs(52));
    layer0_outputs(2622) <= not(inputs(214));
    layer0_outputs(2623) <= inputs(114);
    layer0_outputs(2624) <= not(inputs(9));
    layer0_outputs(2625) <= not(inputs(17)) or (inputs(75));
    layer0_outputs(2626) <= not(inputs(238));
    layer0_outputs(2627) <= not(inputs(210)) or (inputs(133));
    layer0_outputs(2628) <= (inputs(233)) or (inputs(2));
    layer0_outputs(2629) <= not(inputs(141)) or (inputs(110));
    layer0_outputs(2630) <= (inputs(62)) or (inputs(206));
    layer0_outputs(2631) <= (inputs(156)) and not (inputs(225));
    layer0_outputs(2632) <= (inputs(160)) or (inputs(251));
    layer0_outputs(2633) <= not((inputs(181)) or (inputs(14)));
    layer0_outputs(2634) <= (inputs(47)) and not (inputs(235));
    layer0_outputs(2635) <= inputs(182);
    layer0_outputs(2636) <= not(inputs(169));
    layer0_outputs(2637) <= not(inputs(132)) or (inputs(226));
    layer0_outputs(2638) <= not(inputs(195));
    layer0_outputs(2639) <= (inputs(251)) xor (inputs(165));
    layer0_outputs(2640) <= not((inputs(96)) or (inputs(49)));
    layer0_outputs(2641) <= not(inputs(154));
    layer0_outputs(2642) <= (inputs(214)) xor (inputs(172));
    layer0_outputs(2643) <= not((inputs(200)) or (inputs(141)));
    layer0_outputs(2644) <= (inputs(6)) xor (inputs(42));
    layer0_outputs(2645) <= inputs(173);
    layer0_outputs(2646) <= not((inputs(192)) or (inputs(144)));
    layer0_outputs(2647) <= inputs(3);
    layer0_outputs(2648) <= (inputs(188)) xor (inputs(21));
    layer0_outputs(2649) <= not(inputs(12));
    layer0_outputs(2650) <= not((inputs(244)) or (inputs(103)));
    layer0_outputs(2651) <= (inputs(51)) xor (inputs(192));
    layer0_outputs(2652) <= (inputs(200)) or (inputs(151));
    layer0_outputs(2653) <= not(inputs(167));
    layer0_outputs(2654) <= inputs(33);
    layer0_outputs(2655) <= not(inputs(120)) or (inputs(219));
    layer0_outputs(2656) <= not(inputs(109)) or (inputs(115));
    layer0_outputs(2657) <= not((inputs(234)) and (inputs(37)));
    layer0_outputs(2658) <= (inputs(161)) and not (inputs(223));
    layer0_outputs(2659) <= inputs(101);
    layer0_outputs(2660) <= not((inputs(196)) or (inputs(10)));
    layer0_outputs(2661) <= (inputs(173)) and not (inputs(76));
    layer0_outputs(2662) <= (inputs(101)) and not (inputs(124));
    layer0_outputs(2663) <= (inputs(139)) and (inputs(157));
    layer0_outputs(2664) <= (inputs(193)) or (inputs(35));
    layer0_outputs(2665) <= (inputs(35)) and (inputs(217));
    layer0_outputs(2666) <= not((inputs(121)) or (inputs(93)));
    layer0_outputs(2667) <= inputs(59);
    layer0_outputs(2668) <= not(inputs(163)) or (inputs(160));
    layer0_outputs(2669) <= inputs(122);
    layer0_outputs(2670) <= not(inputs(248));
    layer0_outputs(2671) <= not(inputs(197));
    layer0_outputs(2672) <= (inputs(3)) xor (inputs(119));
    layer0_outputs(2673) <= not((inputs(20)) xor (inputs(140)));
    layer0_outputs(2674) <= (inputs(245)) or (inputs(19));
    layer0_outputs(2675) <= not((inputs(175)) or (inputs(201)));
    layer0_outputs(2676) <= not((inputs(145)) xor (inputs(173)));
    layer0_outputs(2677) <= (inputs(123)) xor (inputs(38));
    layer0_outputs(2678) <= not(inputs(85));
    layer0_outputs(2679) <= not((inputs(152)) xor (inputs(164)));
    layer0_outputs(2680) <= not((inputs(251)) or (inputs(106)));
    layer0_outputs(2681) <= not((inputs(211)) or (inputs(212)));
    layer0_outputs(2682) <= inputs(21);
    layer0_outputs(2683) <= not((inputs(156)) or (inputs(126)));
    layer0_outputs(2684) <= not(inputs(59)) or (inputs(159));
    layer0_outputs(2685) <= not(inputs(118));
    layer0_outputs(2686) <= (inputs(70)) xor (inputs(64));
    layer0_outputs(2687) <= (inputs(173)) and not (inputs(45));
    layer0_outputs(2688) <= not(inputs(109));
    layer0_outputs(2689) <= (inputs(166)) xor (inputs(146));
    layer0_outputs(2690) <= (inputs(220)) and not (inputs(100));
    layer0_outputs(2691) <= not(inputs(9)) or (inputs(24));
    layer0_outputs(2692) <= not(inputs(23)) or (inputs(11));
    layer0_outputs(2693) <= not(inputs(18));
    layer0_outputs(2694) <= not((inputs(87)) xor (inputs(69)));
    layer0_outputs(2695) <= (inputs(247)) and not (inputs(47));
    layer0_outputs(2696) <= not((inputs(204)) or (inputs(175)));
    layer0_outputs(2697) <= inputs(154);
    layer0_outputs(2698) <= not(inputs(202)) or (inputs(44));
    layer0_outputs(2699) <= (inputs(62)) and not (inputs(105));
    layer0_outputs(2700) <= inputs(164);
    layer0_outputs(2701) <= inputs(24);
    layer0_outputs(2702) <= not((inputs(196)) or (inputs(235)));
    layer0_outputs(2703) <= not((inputs(38)) or (inputs(169)));
    layer0_outputs(2704) <= not(inputs(184)) or (inputs(250));
    layer0_outputs(2705) <= not(inputs(209)) or (inputs(140));
    layer0_outputs(2706) <= inputs(104);
    layer0_outputs(2707) <= not(inputs(230));
    layer0_outputs(2708) <= not((inputs(161)) xor (inputs(177)));
    layer0_outputs(2709) <= not(inputs(61)) or (inputs(124));
    layer0_outputs(2710) <= (inputs(119)) and not (inputs(142));
    layer0_outputs(2711) <= not(inputs(2)) or (inputs(66));
    layer0_outputs(2712) <= (inputs(102)) or (inputs(202));
    layer0_outputs(2713) <= not(inputs(122)) or (inputs(225));
    layer0_outputs(2714) <= (inputs(205)) and not (inputs(222));
    layer0_outputs(2715) <= (inputs(20)) xor (inputs(48));
    layer0_outputs(2716) <= (inputs(211)) or (inputs(208));
    layer0_outputs(2717) <= (inputs(166)) or (inputs(121));
    layer0_outputs(2718) <= not((inputs(200)) or (inputs(199)));
    layer0_outputs(2719) <= inputs(6);
    layer0_outputs(2720) <= not(inputs(80)) or (inputs(157));
    layer0_outputs(2721) <= not((inputs(169)) or (inputs(216)));
    layer0_outputs(2722) <= inputs(21);
    layer0_outputs(2723) <= inputs(58);
    layer0_outputs(2724) <= inputs(98);
    layer0_outputs(2725) <= not(inputs(121));
    layer0_outputs(2726) <= not((inputs(89)) xor (inputs(18)));
    layer0_outputs(2727) <= '0';
    layer0_outputs(2728) <= inputs(72);
    layer0_outputs(2729) <= (inputs(35)) or (inputs(157));
    layer0_outputs(2730) <= not(inputs(82)) or (inputs(224));
    layer0_outputs(2731) <= not((inputs(85)) or (inputs(66)));
    layer0_outputs(2732) <= (inputs(112)) or (inputs(21));
    layer0_outputs(2733) <= not(inputs(63));
    layer0_outputs(2734) <= inputs(103);
    layer0_outputs(2735) <= (inputs(202)) and not (inputs(91));
    layer0_outputs(2736) <= not((inputs(181)) xor (inputs(211)));
    layer0_outputs(2737) <= not(inputs(158));
    layer0_outputs(2738) <= not(inputs(118)) or (inputs(6));
    layer0_outputs(2739) <= not(inputs(251));
    layer0_outputs(2740) <= (inputs(230)) and not (inputs(165));
    layer0_outputs(2741) <= not(inputs(72));
    layer0_outputs(2742) <= (inputs(250)) or (inputs(6));
    layer0_outputs(2743) <= not((inputs(186)) xor (inputs(101)));
    layer0_outputs(2744) <= not(inputs(23)) or (inputs(129));
    layer0_outputs(2745) <= (inputs(214)) or (inputs(129));
    layer0_outputs(2746) <= (inputs(103)) and not (inputs(108));
    layer0_outputs(2747) <= (inputs(115)) xor (inputs(103));
    layer0_outputs(2748) <= not(inputs(144));
    layer0_outputs(2749) <= not(inputs(132));
    layer0_outputs(2750) <= (inputs(35)) and not (inputs(58));
    layer0_outputs(2751) <= (inputs(183)) and not (inputs(99));
    layer0_outputs(2752) <= (inputs(42)) and not (inputs(16));
    layer0_outputs(2753) <= not(inputs(158)) or (inputs(146));
    layer0_outputs(2754) <= not((inputs(0)) or (inputs(133)));
    layer0_outputs(2755) <= (inputs(46)) xor (inputs(18));
    layer0_outputs(2756) <= not(inputs(187));
    layer0_outputs(2757) <= not((inputs(206)) or (inputs(243)));
    layer0_outputs(2758) <= (inputs(29)) or (inputs(218));
    layer0_outputs(2759) <= not((inputs(148)) xor (inputs(103)));
    layer0_outputs(2760) <= not(inputs(238));
    layer0_outputs(2761) <= inputs(164);
    layer0_outputs(2762) <= inputs(23);
    layer0_outputs(2763) <= not((inputs(253)) or (inputs(147)));
    layer0_outputs(2764) <= not(inputs(106));
    layer0_outputs(2765) <= not(inputs(235)) or (inputs(93));
    layer0_outputs(2766) <= not((inputs(123)) xor (inputs(172)));
    layer0_outputs(2767) <= not((inputs(202)) xor (inputs(65)));
    layer0_outputs(2768) <= (inputs(204)) or (inputs(101));
    layer0_outputs(2769) <= (inputs(189)) or (inputs(2));
    layer0_outputs(2770) <= (inputs(173)) xor (inputs(158));
    layer0_outputs(2771) <= not(inputs(7));
    layer0_outputs(2772) <= (inputs(238)) and not (inputs(207));
    layer0_outputs(2773) <= (inputs(190)) xor (inputs(63));
    layer0_outputs(2774) <= (inputs(187)) or (inputs(18));
    layer0_outputs(2775) <= (inputs(118)) or (inputs(98));
    layer0_outputs(2776) <= not(inputs(53)) or (inputs(102));
    layer0_outputs(2777) <= not(inputs(98));
    layer0_outputs(2778) <= (inputs(100)) xor (inputs(196));
    layer0_outputs(2779) <= not((inputs(209)) xor (inputs(204)));
    layer0_outputs(2780) <= not((inputs(192)) xor (inputs(204)));
    layer0_outputs(2781) <= (inputs(31)) or (inputs(18));
    layer0_outputs(2782) <= not(inputs(80));
    layer0_outputs(2783) <= (inputs(243)) and not (inputs(254));
    layer0_outputs(2784) <= not((inputs(213)) xor (inputs(167)));
    layer0_outputs(2785) <= inputs(169);
    layer0_outputs(2786) <= inputs(139);
    layer0_outputs(2787) <= not(inputs(115));
    layer0_outputs(2788) <= inputs(132);
    layer0_outputs(2789) <= inputs(219);
    layer0_outputs(2790) <= not((inputs(228)) or (inputs(181)));
    layer0_outputs(2791) <= (inputs(144)) or (inputs(247));
    layer0_outputs(2792) <= not((inputs(58)) and (inputs(71)));
    layer0_outputs(2793) <= not((inputs(179)) xor (inputs(177)));
    layer0_outputs(2794) <= (inputs(141)) or (inputs(124));
    layer0_outputs(2795) <= (inputs(249)) xor (inputs(71));
    layer0_outputs(2796) <= not((inputs(229)) xor (inputs(197)));
    layer0_outputs(2797) <= not((inputs(47)) or (inputs(219)));
    layer0_outputs(2798) <= inputs(198);
    layer0_outputs(2799) <= not(inputs(100));
    layer0_outputs(2800) <= not((inputs(224)) and (inputs(42)));
    layer0_outputs(2801) <= not(inputs(23)) or (inputs(91));
    layer0_outputs(2802) <= not((inputs(26)) or (inputs(67)));
    layer0_outputs(2803) <= not(inputs(227)) or (inputs(76));
    layer0_outputs(2804) <= not(inputs(167)) or (inputs(78));
    layer0_outputs(2805) <= (inputs(184)) and not (inputs(103));
    layer0_outputs(2806) <= not(inputs(227));
    layer0_outputs(2807) <= (inputs(95)) or (inputs(11));
    layer0_outputs(2808) <= inputs(190);
    layer0_outputs(2809) <= not(inputs(194)) or (inputs(125));
    layer0_outputs(2810) <= not(inputs(214)) or (inputs(46));
    layer0_outputs(2811) <= (inputs(175)) and not (inputs(1));
    layer0_outputs(2812) <= (inputs(16)) or (inputs(255));
    layer0_outputs(2813) <= (inputs(151)) and not (inputs(125));
    layer0_outputs(2814) <= (inputs(206)) and not (inputs(250));
    layer0_outputs(2815) <= not((inputs(212)) xor (inputs(211)));
    layer0_outputs(2816) <= not(inputs(45));
    layer0_outputs(2817) <= inputs(58);
    layer0_outputs(2818) <= not(inputs(200));
    layer0_outputs(2819) <= not(inputs(51));
    layer0_outputs(2820) <= not(inputs(181));
    layer0_outputs(2821) <= not(inputs(99)) or (inputs(122));
    layer0_outputs(2822) <= inputs(60);
    layer0_outputs(2823) <= not((inputs(185)) or (inputs(251)));
    layer0_outputs(2824) <= '0';
    layer0_outputs(2825) <= (inputs(197)) and not (inputs(208));
    layer0_outputs(2826) <= not(inputs(45));
    layer0_outputs(2827) <= (inputs(198)) xor (inputs(185));
    layer0_outputs(2828) <= not(inputs(74));
    layer0_outputs(2829) <= inputs(37);
    layer0_outputs(2830) <= not(inputs(82));
    layer0_outputs(2831) <= inputs(43);
    layer0_outputs(2832) <= not((inputs(6)) or (inputs(229)));
    layer0_outputs(2833) <= inputs(74);
    layer0_outputs(2834) <= not(inputs(125)) or (inputs(222));
    layer0_outputs(2835) <= inputs(111);
    layer0_outputs(2836) <= not((inputs(159)) or (inputs(12)));
    layer0_outputs(2837) <= not((inputs(5)) xor (inputs(210)));
    layer0_outputs(2838) <= not(inputs(231)) or (inputs(129));
    layer0_outputs(2839) <= (inputs(24)) and not (inputs(237));
    layer0_outputs(2840) <= inputs(23);
    layer0_outputs(2841) <= inputs(57);
    layer0_outputs(2842) <= (inputs(190)) xor (inputs(9));
    layer0_outputs(2843) <= not((inputs(80)) or (inputs(128)));
    layer0_outputs(2844) <= inputs(9);
    layer0_outputs(2845) <= (inputs(144)) and (inputs(82));
    layer0_outputs(2846) <= (inputs(193)) or (inputs(33));
    layer0_outputs(2847) <= (inputs(159)) or (inputs(148));
    layer0_outputs(2848) <= not(inputs(118)) or (inputs(95));
    layer0_outputs(2849) <= inputs(160);
    layer0_outputs(2850) <= (inputs(63)) or (inputs(46));
    layer0_outputs(2851) <= (inputs(30)) and not (inputs(110));
    layer0_outputs(2852) <= inputs(105);
    layer0_outputs(2853) <= not((inputs(129)) or (inputs(219)));
    layer0_outputs(2854) <= inputs(58);
    layer0_outputs(2855) <= not((inputs(100)) xor (inputs(70)));
    layer0_outputs(2856) <= not(inputs(235)) or (inputs(5));
    layer0_outputs(2857) <= not(inputs(180)) or (inputs(112));
    layer0_outputs(2858) <= inputs(67);
    layer0_outputs(2859) <= not((inputs(217)) and (inputs(182)));
    layer0_outputs(2860) <= (inputs(246)) or (inputs(148));
    layer0_outputs(2861) <= not((inputs(201)) or (inputs(251)));
    layer0_outputs(2862) <= (inputs(250)) or (inputs(69));
    layer0_outputs(2863) <= (inputs(188)) and not (inputs(27));
    layer0_outputs(2864) <= not(inputs(151));
    layer0_outputs(2865) <= not(inputs(195));
    layer0_outputs(2866) <= (inputs(196)) xor (inputs(167));
    layer0_outputs(2867) <= not(inputs(65)) or (inputs(252));
    layer0_outputs(2868) <= not(inputs(109));
    layer0_outputs(2869) <= not(inputs(8)) or (inputs(230));
    layer0_outputs(2870) <= not((inputs(151)) or (inputs(1)));
    layer0_outputs(2871) <= (inputs(25)) and not (inputs(14));
    layer0_outputs(2872) <= not((inputs(247)) xor (inputs(175)));
    layer0_outputs(2873) <= (inputs(85)) and not (inputs(248));
    layer0_outputs(2874) <= (inputs(82)) xor (inputs(87));
    layer0_outputs(2875) <= (inputs(3)) or (inputs(178));
    layer0_outputs(2876) <= not(inputs(14));
    layer0_outputs(2877) <= not(inputs(219));
    layer0_outputs(2878) <= (inputs(77)) and not (inputs(30));
    layer0_outputs(2879) <= not(inputs(66));
    layer0_outputs(2880) <= not((inputs(255)) or (inputs(54)));
    layer0_outputs(2881) <= (inputs(196)) and not (inputs(74));
    layer0_outputs(2882) <= not((inputs(42)) or (inputs(169)));
    layer0_outputs(2883) <= not(inputs(95)) or (inputs(43));
    layer0_outputs(2884) <= not((inputs(6)) or (inputs(130)));
    layer0_outputs(2885) <= (inputs(73)) xor (inputs(117));
    layer0_outputs(2886) <= not(inputs(46));
    layer0_outputs(2887) <= (inputs(221)) or (inputs(253));
    layer0_outputs(2888) <= not(inputs(92));
    layer0_outputs(2889) <= inputs(141);
    layer0_outputs(2890) <= (inputs(203)) xor (inputs(84));
    layer0_outputs(2891) <= not(inputs(76));
    layer0_outputs(2892) <= not(inputs(142));
    layer0_outputs(2893) <= (inputs(168)) and (inputs(40));
    layer0_outputs(2894) <= not(inputs(103)) or (inputs(129));
    layer0_outputs(2895) <= inputs(193);
    layer0_outputs(2896) <= not((inputs(146)) or (inputs(35)));
    layer0_outputs(2897) <= not((inputs(241)) xor (inputs(161)));
    layer0_outputs(2898) <= not((inputs(108)) and (inputs(75)));
    layer0_outputs(2899) <= not(inputs(69)) or (inputs(194));
    layer0_outputs(2900) <= (inputs(222)) or (inputs(55));
    layer0_outputs(2901) <= (inputs(18)) or (inputs(166));
    layer0_outputs(2902) <= not((inputs(171)) or (inputs(8)));
    layer0_outputs(2903) <= (inputs(172)) and not (inputs(94));
    layer0_outputs(2904) <= not((inputs(172)) and (inputs(236)));
    layer0_outputs(2905) <= inputs(187);
    layer0_outputs(2906) <= not(inputs(209)) or (inputs(138));
    layer0_outputs(2907) <= not((inputs(202)) and (inputs(7)));
    layer0_outputs(2908) <= (inputs(42)) and not (inputs(219));
    layer0_outputs(2909) <= not(inputs(188)) or (inputs(110));
    layer0_outputs(2910) <= not((inputs(128)) or (inputs(45)));
    layer0_outputs(2911) <= inputs(113);
    layer0_outputs(2912) <= not(inputs(83)) or (inputs(28));
    layer0_outputs(2913) <= not((inputs(137)) xor (inputs(156)));
    layer0_outputs(2914) <= (inputs(231)) and not (inputs(146));
    layer0_outputs(2915) <= not(inputs(26)) or (inputs(226));
    layer0_outputs(2916) <= not(inputs(19));
    layer0_outputs(2917) <= (inputs(192)) xor (inputs(88));
    layer0_outputs(2918) <= inputs(151);
    layer0_outputs(2919) <= not(inputs(30));
    layer0_outputs(2920) <= not((inputs(82)) xor (inputs(177)));
    layer0_outputs(2921) <= not(inputs(231));
    layer0_outputs(2922) <= (inputs(60)) or (inputs(33));
    layer0_outputs(2923) <= not(inputs(82)) or (inputs(251));
    layer0_outputs(2924) <= (inputs(229)) or (inputs(207));
    layer0_outputs(2925) <= inputs(193);
    layer0_outputs(2926) <= not(inputs(200)) or (inputs(79));
    layer0_outputs(2927) <= not((inputs(52)) or (inputs(160)));
    layer0_outputs(2928) <= (inputs(165)) xor (inputs(147));
    layer0_outputs(2929) <= not((inputs(77)) or (inputs(77)));
    layer0_outputs(2930) <= not(inputs(161));
    layer0_outputs(2931) <= (inputs(51)) or (inputs(146));
    layer0_outputs(2932) <= inputs(120);
    layer0_outputs(2933) <= (inputs(30)) or (inputs(140));
    layer0_outputs(2934) <= not(inputs(43)) or (inputs(227));
    layer0_outputs(2935) <= not((inputs(189)) xor (inputs(178)));
    layer0_outputs(2936) <= (inputs(12)) xor (inputs(71));
    layer0_outputs(2937) <= not(inputs(49));
    layer0_outputs(2938) <= not(inputs(18));
    layer0_outputs(2939) <= not((inputs(124)) xor (inputs(113)));
    layer0_outputs(2940) <= not((inputs(200)) or (inputs(109)));
    layer0_outputs(2941) <= inputs(58);
    layer0_outputs(2942) <= (inputs(198)) and (inputs(87));
    layer0_outputs(2943) <= not((inputs(115)) and (inputs(241)));
    layer0_outputs(2944) <= not(inputs(89));
    layer0_outputs(2945) <= inputs(167);
    layer0_outputs(2946) <= not(inputs(123)) or (inputs(205));
    layer0_outputs(2947) <= not(inputs(31)) or (inputs(244));
    layer0_outputs(2948) <= (inputs(197)) and not (inputs(240));
    layer0_outputs(2949) <= (inputs(217)) xor (inputs(93));
    layer0_outputs(2950) <= (inputs(77)) or (inputs(164));
    layer0_outputs(2951) <= not((inputs(142)) or (inputs(203)));
    layer0_outputs(2952) <= (inputs(9)) and not (inputs(145));
    layer0_outputs(2953) <= not(inputs(3)) or (inputs(241));
    layer0_outputs(2954) <= inputs(10);
    layer0_outputs(2955) <= inputs(119);
    layer0_outputs(2956) <= not(inputs(115));
    layer0_outputs(2957) <= not((inputs(162)) xor (inputs(248)));
    layer0_outputs(2958) <= (inputs(228)) or (inputs(148));
    layer0_outputs(2959) <= (inputs(128)) and not (inputs(253));
    layer0_outputs(2960) <= inputs(103);
    layer0_outputs(2961) <= (inputs(184)) xor (inputs(215));
    layer0_outputs(2962) <= not(inputs(131)) or (inputs(13));
    layer0_outputs(2963) <= not(inputs(62)) or (inputs(108));
    layer0_outputs(2964) <= '1';
    layer0_outputs(2965) <= not((inputs(88)) and (inputs(1)));
    layer0_outputs(2966) <= not((inputs(190)) xor (inputs(42)));
    layer0_outputs(2967) <= not(inputs(19)) or (inputs(129));
    layer0_outputs(2968) <= (inputs(22)) xor (inputs(102));
    layer0_outputs(2969) <= (inputs(42)) and not (inputs(146));
    layer0_outputs(2970) <= '1';
    layer0_outputs(2971) <= (inputs(13)) or (inputs(212));
    layer0_outputs(2972) <= not((inputs(70)) or (inputs(73)));
    layer0_outputs(2973) <= (inputs(18)) or (inputs(238));
    layer0_outputs(2974) <= inputs(178);
    layer0_outputs(2975) <= not(inputs(209)) or (inputs(5));
    layer0_outputs(2976) <= not(inputs(196));
    layer0_outputs(2977) <= (inputs(17)) or (inputs(213));
    layer0_outputs(2978) <= (inputs(136)) and not (inputs(208));
    layer0_outputs(2979) <= not((inputs(224)) xor (inputs(206)));
    layer0_outputs(2980) <= (inputs(69)) and not (inputs(77));
    layer0_outputs(2981) <= '0';
    layer0_outputs(2982) <= inputs(202);
    layer0_outputs(2983) <= (inputs(208)) xor (inputs(183));
    layer0_outputs(2984) <= (inputs(252)) or (inputs(81));
    layer0_outputs(2985) <= not((inputs(138)) or (inputs(207)));
    layer0_outputs(2986) <= (inputs(205)) and not (inputs(31));
    layer0_outputs(2987) <= not((inputs(78)) or (inputs(126)));
    layer0_outputs(2988) <= not((inputs(255)) xor (inputs(56)));
    layer0_outputs(2989) <= (inputs(25)) or (inputs(155));
    layer0_outputs(2990) <= (inputs(197)) and not (inputs(112));
    layer0_outputs(2991) <= (inputs(18)) or (inputs(178));
    layer0_outputs(2992) <= (inputs(228)) or (inputs(114));
    layer0_outputs(2993) <= (inputs(222)) xor (inputs(156));
    layer0_outputs(2994) <= inputs(211);
    layer0_outputs(2995) <= (inputs(190)) xor (inputs(238));
    layer0_outputs(2996) <= inputs(162);
    layer0_outputs(2997) <= (inputs(37)) or (inputs(87));
    layer0_outputs(2998) <= '0';
    layer0_outputs(2999) <= not((inputs(191)) or (inputs(235)));
    layer0_outputs(3000) <= (inputs(80)) xor (inputs(60));
    layer0_outputs(3001) <= (inputs(40)) and not (inputs(243));
    layer0_outputs(3002) <= inputs(162);
    layer0_outputs(3003) <= not(inputs(37));
    layer0_outputs(3004) <= not((inputs(0)) or (inputs(12)));
    layer0_outputs(3005) <= (inputs(139)) xor (inputs(189));
    layer0_outputs(3006) <= (inputs(76)) and (inputs(96));
    layer0_outputs(3007) <= inputs(157);
    layer0_outputs(3008) <= not(inputs(220)) or (inputs(244));
    layer0_outputs(3009) <= (inputs(98)) and not (inputs(94));
    layer0_outputs(3010) <= not(inputs(226)) or (inputs(54));
    layer0_outputs(3011) <= not((inputs(70)) xor (inputs(53)));
    layer0_outputs(3012) <= not((inputs(245)) or (inputs(143)));
    layer0_outputs(3013) <= inputs(118);
    layer0_outputs(3014) <= inputs(130);
    layer0_outputs(3015) <= not((inputs(24)) or (inputs(191)));
    layer0_outputs(3016) <= inputs(27);
    layer0_outputs(3017) <= not(inputs(173));
    layer0_outputs(3018) <= (inputs(205)) xor (inputs(95));
    layer0_outputs(3019) <= not(inputs(197));
    layer0_outputs(3020) <= not(inputs(26)) or (inputs(241));
    layer0_outputs(3021) <= (inputs(185)) and (inputs(31));
    layer0_outputs(3022) <= (inputs(85)) and not (inputs(48));
    layer0_outputs(3023) <= not((inputs(102)) or (inputs(69)));
    layer0_outputs(3024) <= (inputs(74)) and not (inputs(197));
    layer0_outputs(3025) <= not((inputs(219)) xor (inputs(37)));
    layer0_outputs(3026) <= inputs(180);
    layer0_outputs(3027) <= not((inputs(181)) xor (inputs(138)));
    layer0_outputs(3028) <= not((inputs(135)) xor (inputs(33)));
    layer0_outputs(3029) <= (inputs(174)) and not (inputs(94));
    layer0_outputs(3030) <= (inputs(150)) and not (inputs(97));
    layer0_outputs(3031) <= inputs(164);
    layer0_outputs(3032) <= inputs(120);
    layer0_outputs(3033) <= not(inputs(84));
    layer0_outputs(3034) <= (inputs(118)) or (inputs(234));
    layer0_outputs(3035) <= (inputs(102)) and not (inputs(234));
    layer0_outputs(3036) <= inputs(90);
    layer0_outputs(3037) <= (inputs(32)) and not (inputs(13));
    layer0_outputs(3038) <= inputs(105);
    layer0_outputs(3039) <= (inputs(137)) and not (inputs(213));
    layer0_outputs(3040) <= inputs(93);
    layer0_outputs(3041) <= not((inputs(137)) xor (inputs(131)));
    layer0_outputs(3042) <= (inputs(170)) xor (inputs(136));
    layer0_outputs(3043) <= (inputs(26)) xor (inputs(36));
    layer0_outputs(3044) <= not(inputs(229));
    layer0_outputs(3045) <= inputs(197);
    layer0_outputs(3046) <= inputs(114);
    layer0_outputs(3047) <= inputs(97);
    layer0_outputs(3048) <= inputs(203);
    layer0_outputs(3049) <= not(inputs(165)) or (inputs(97));
    layer0_outputs(3050) <= not(inputs(41));
    layer0_outputs(3051) <= not((inputs(17)) or (inputs(135)));
    layer0_outputs(3052) <= not(inputs(31));
    layer0_outputs(3053) <= inputs(50);
    layer0_outputs(3054) <= not(inputs(25));
    layer0_outputs(3055) <= inputs(125);
    layer0_outputs(3056) <= not(inputs(27));
    layer0_outputs(3057) <= (inputs(69)) and not (inputs(239));
    layer0_outputs(3058) <= inputs(229);
    layer0_outputs(3059) <= (inputs(27)) and not (inputs(254));
    layer0_outputs(3060) <= not((inputs(70)) or (inputs(159)));
    layer0_outputs(3061) <= not(inputs(160));
    layer0_outputs(3062) <= not(inputs(75)) or (inputs(176));
    layer0_outputs(3063) <= (inputs(168)) or (inputs(49));
    layer0_outputs(3064) <= (inputs(247)) and not (inputs(11));
    layer0_outputs(3065) <= not((inputs(100)) xor (inputs(76)));
    layer0_outputs(3066) <= not(inputs(130));
    layer0_outputs(3067) <= not(inputs(82));
    layer0_outputs(3068) <= not(inputs(208)) or (inputs(174));
    layer0_outputs(3069) <= not((inputs(128)) or (inputs(29)));
    layer0_outputs(3070) <= (inputs(255)) and (inputs(102));
    layer0_outputs(3071) <= not((inputs(84)) or (inputs(46)));
    layer0_outputs(3072) <= (inputs(155)) or (inputs(242));
    layer0_outputs(3073) <= not(inputs(215));
    layer0_outputs(3074) <= inputs(9);
    layer0_outputs(3075) <= (inputs(11)) or (inputs(253));
    layer0_outputs(3076) <= not((inputs(82)) and (inputs(243)));
    layer0_outputs(3077) <= (inputs(3)) or (inputs(219));
    layer0_outputs(3078) <= not(inputs(199)) or (inputs(96));
    layer0_outputs(3079) <= inputs(101);
    layer0_outputs(3080) <= not((inputs(50)) or (inputs(179)));
    layer0_outputs(3081) <= inputs(235);
    layer0_outputs(3082) <= not((inputs(40)) or (inputs(16)));
    layer0_outputs(3083) <= not((inputs(128)) xor (inputs(148)));
    layer0_outputs(3084) <= not(inputs(3));
    layer0_outputs(3085) <= (inputs(7)) and (inputs(25));
    layer0_outputs(3086) <= not((inputs(74)) and (inputs(53)));
    layer0_outputs(3087) <= inputs(178);
    layer0_outputs(3088) <= not((inputs(11)) xor (inputs(46)));
    layer0_outputs(3089) <= not((inputs(207)) or (inputs(126)));
    layer0_outputs(3090) <= not(inputs(95)) or (inputs(205));
    layer0_outputs(3091) <= not(inputs(108));
    layer0_outputs(3092) <= (inputs(60)) and not (inputs(237));
    layer0_outputs(3093) <= (inputs(3)) or (inputs(45));
    layer0_outputs(3094) <= inputs(231);
    layer0_outputs(3095) <= not(inputs(121));
    layer0_outputs(3096) <= (inputs(113)) and not (inputs(16));
    layer0_outputs(3097) <= (inputs(58)) xor (inputs(86));
    layer0_outputs(3098) <= (inputs(246)) xor (inputs(139));
    layer0_outputs(3099) <= not((inputs(166)) or (inputs(145)));
    layer0_outputs(3100) <= inputs(233);
    layer0_outputs(3101) <= not((inputs(58)) xor (inputs(10)));
    layer0_outputs(3102) <= (inputs(241)) and (inputs(79));
    layer0_outputs(3103) <= not((inputs(124)) xor (inputs(205)));
    layer0_outputs(3104) <= not((inputs(243)) or (inputs(217)));
    layer0_outputs(3105) <= inputs(69);
    layer0_outputs(3106) <= (inputs(255)) or (inputs(216));
    layer0_outputs(3107) <= inputs(23);
    layer0_outputs(3108) <= (inputs(97)) or (inputs(112));
    layer0_outputs(3109) <= not((inputs(37)) or (inputs(205)));
    layer0_outputs(3110) <= (inputs(230)) or (inputs(238));
    layer0_outputs(3111) <= not(inputs(83));
    layer0_outputs(3112) <= (inputs(56)) or (inputs(16));
    layer0_outputs(3113) <= inputs(152);
    layer0_outputs(3114) <= not(inputs(29)) or (inputs(176));
    layer0_outputs(3115) <= (inputs(117)) and not (inputs(104));
    layer0_outputs(3116) <= inputs(81);
    layer0_outputs(3117) <= inputs(6);
    layer0_outputs(3118) <= not(inputs(93));
    layer0_outputs(3119) <= not((inputs(211)) xor (inputs(166)));
    layer0_outputs(3120) <= (inputs(195)) and not (inputs(175));
    layer0_outputs(3121) <= not(inputs(114));
    layer0_outputs(3122) <= not(inputs(76)) or (inputs(238));
    layer0_outputs(3123) <= not(inputs(94));
    layer0_outputs(3124) <= (inputs(74)) and not (inputs(147));
    layer0_outputs(3125) <= (inputs(219)) xor (inputs(75));
    layer0_outputs(3126) <= not(inputs(203)) or (inputs(251));
    layer0_outputs(3127) <= (inputs(98)) or (inputs(154));
    layer0_outputs(3128) <= (inputs(142)) xor (inputs(18));
    layer0_outputs(3129) <= inputs(56);
    layer0_outputs(3130) <= (inputs(236)) or (inputs(147));
    layer0_outputs(3131) <= not(inputs(32));
    layer0_outputs(3132) <= (inputs(237)) xor (inputs(19));
    layer0_outputs(3133) <= inputs(208);
    layer0_outputs(3134) <= not((inputs(97)) or (inputs(124)));
    layer0_outputs(3135) <= not(inputs(148));
    layer0_outputs(3136) <= not(inputs(147));
    layer0_outputs(3137) <= not(inputs(165));
    layer0_outputs(3138) <= not((inputs(195)) xor (inputs(89)));
    layer0_outputs(3139) <= (inputs(116)) and not (inputs(194));
    layer0_outputs(3140) <= not(inputs(57));
    layer0_outputs(3141) <= (inputs(151)) and not (inputs(85));
    layer0_outputs(3142) <= not(inputs(72)) or (inputs(15));
    layer0_outputs(3143) <= not(inputs(235));
    layer0_outputs(3144) <= (inputs(234)) or (inputs(158));
    layer0_outputs(3145) <= not(inputs(221));
    layer0_outputs(3146) <= inputs(44);
    layer0_outputs(3147) <= inputs(72);
    layer0_outputs(3148) <= not((inputs(17)) or (inputs(124)));
    layer0_outputs(3149) <= not(inputs(206));
    layer0_outputs(3150) <= inputs(19);
    layer0_outputs(3151) <= not((inputs(202)) xor (inputs(54)));
    layer0_outputs(3152) <= (inputs(200)) and not (inputs(67));
    layer0_outputs(3153) <= (inputs(224)) and not (inputs(122));
    layer0_outputs(3154) <= inputs(31);
    layer0_outputs(3155) <= not((inputs(112)) xor (inputs(26)));
    layer0_outputs(3156) <= not((inputs(194)) xor (inputs(81)));
    layer0_outputs(3157) <= not(inputs(82)) or (inputs(73));
    layer0_outputs(3158) <= (inputs(106)) and not (inputs(18));
    layer0_outputs(3159) <= not((inputs(211)) or (inputs(104)));
    layer0_outputs(3160) <= (inputs(228)) xor (inputs(24));
    layer0_outputs(3161) <= not((inputs(71)) and (inputs(161)));
    layer0_outputs(3162) <= not(inputs(118));
    layer0_outputs(3163) <= not(inputs(23));
    layer0_outputs(3164) <= (inputs(179)) or (inputs(158));
    layer0_outputs(3165) <= (inputs(76)) or (inputs(210));
    layer0_outputs(3166) <= not(inputs(4)) or (inputs(84));
    layer0_outputs(3167) <= not((inputs(48)) or (inputs(151)));
    layer0_outputs(3168) <= inputs(214);
    layer0_outputs(3169) <= not(inputs(240));
    layer0_outputs(3170) <= (inputs(90)) or (inputs(18));
    layer0_outputs(3171) <= not(inputs(107));
    layer0_outputs(3172) <= (inputs(217)) and not (inputs(90));
    layer0_outputs(3173) <= not(inputs(105)) or (inputs(46));
    layer0_outputs(3174) <= (inputs(144)) or (inputs(212));
    layer0_outputs(3175) <= (inputs(205)) and not (inputs(109));
    layer0_outputs(3176) <= (inputs(13)) or (inputs(138));
    layer0_outputs(3177) <= not(inputs(90)) or (inputs(192));
    layer0_outputs(3178) <= inputs(78);
    layer0_outputs(3179) <= not((inputs(51)) or (inputs(129)));
    layer0_outputs(3180) <= (inputs(106)) xor (inputs(136));
    layer0_outputs(3181) <= (inputs(35)) xor (inputs(149));
    layer0_outputs(3182) <= not((inputs(40)) or (inputs(171)));
    layer0_outputs(3183) <= not(inputs(45)) or (inputs(182));
    layer0_outputs(3184) <= not(inputs(27)) or (inputs(3));
    layer0_outputs(3185) <= not(inputs(174));
    layer0_outputs(3186) <= not(inputs(177));
    layer0_outputs(3187) <= (inputs(78)) xor (inputs(63));
    layer0_outputs(3188) <= not(inputs(20)) or (inputs(178));
    layer0_outputs(3189) <= not(inputs(127));
    layer0_outputs(3190) <= not(inputs(138)) or (inputs(49));
    layer0_outputs(3191) <= inputs(20);
    layer0_outputs(3192) <= inputs(78);
    layer0_outputs(3193) <= not(inputs(188));
    layer0_outputs(3194) <= not((inputs(190)) or (inputs(217)));
    layer0_outputs(3195) <= not(inputs(224)) or (inputs(49));
    layer0_outputs(3196) <= (inputs(175)) or (inputs(229));
    layer0_outputs(3197) <= (inputs(200)) and not (inputs(227));
    layer0_outputs(3198) <= (inputs(166)) xor (inputs(196));
    layer0_outputs(3199) <= '1';
    layer0_outputs(3200) <= (inputs(71)) and not (inputs(206));
    layer0_outputs(3201) <= not((inputs(111)) xor (inputs(235)));
    layer0_outputs(3202) <= (inputs(11)) or (inputs(147));
    layer0_outputs(3203) <= not(inputs(151)) or (inputs(157));
    layer0_outputs(3204) <= (inputs(31)) and not (inputs(136));
    layer0_outputs(3205) <= not(inputs(232));
    layer0_outputs(3206) <= (inputs(47)) and not (inputs(209));
    layer0_outputs(3207) <= (inputs(234)) and not (inputs(143));
    layer0_outputs(3208) <= '0';
    layer0_outputs(3209) <= not(inputs(111));
    layer0_outputs(3210) <= not(inputs(184)) or (inputs(192));
    layer0_outputs(3211) <= not((inputs(22)) or (inputs(188)));
    layer0_outputs(3212) <= not(inputs(210)) or (inputs(247));
    layer0_outputs(3213) <= not(inputs(99));
    layer0_outputs(3214) <= not(inputs(63));
    layer0_outputs(3215) <= not(inputs(164));
    layer0_outputs(3216) <= not((inputs(219)) or (inputs(225)));
    layer0_outputs(3217) <= inputs(230);
    layer0_outputs(3218) <= not(inputs(61));
    layer0_outputs(3219) <= (inputs(255)) or (inputs(193));
    layer0_outputs(3220) <= (inputs(63)) xor (inputs(203));
    layer0_outputs(3221) <= not((inputs(214)) or (inputs(97)));
    layer0_outputs(3222) <= not(inputs(58)) or (inputs(186));
    layer0_outputs(3223) <= not((inputs(32)) xor (inputs(132)));
    layer0_outputs(3224) <= not((inputs(3)) or (inputs(4)));
    layer0_outputs(3225) <= not(inputs(248));
    layer0_outputs(3226) <= inputs(37);
    layer0_outputs(3227) <= (inputs(6)) and not (inputs(145));
    layer0_outputs(3228) <= not(inputs(21)) or (inputs(99));
    layer0_outputs(3229) <= '0';
    layer0_outputs(3230) <= (inputs(84)) and (inputs(230));
    layer0_outputs(3231) <= inputs(148);
    layer0_outputs(3232) <= not(inputs(94));
    layer0_outputs(3233) <= inputs(164);
    layer0_outputs(3234) <= not((inputs(169)) xor (inputs(22)));
    layer0_outputs(3235) <= not(inputs(71)) or (inputs(233));
    layer0_outputs(3236) <= not((inputs(149)) xor (inputs(252)));
    layer0_outputs(3237) <= not((inputs(120)) and (inputs(233)));
    layer0_outputs(3238) <= (inputs(71)) or (inputs(128));
    layer0_outputs(3239) <= inputs(208);
    layer0_outputs(3240) <= (inputs(121)) xor (inputs(254));
    layer0_outputs(3241) <= (inputs(84)) and not (inputs(236));
    layer0_outputs(3242) <= inputs(94);
    layer0_outputs(3243) <= inputs(110);
    layer0_outputs(3244) <= (inputs(154)) and not (inputs(242));
    layer0_outputs(3245) <= not(inputs(235));
    layer0_outputs(3246) <= inputs(56);
    layer0_outputs(3247) <= not((inputs(242)) xor (inputs(167)));
    layer0_outputs(3248) <= (inputs(187)) or (inputs(172));
    layer0_outputs(3249) <= (inputs(107)) and not (inputs(141));
    layer0_outputs(3250) <= (inputs(194)) or (inputs(204));
    layer0_outputs(3251) <= not((inputs(233)) or (inputs(5)));
    layer0_outputs(3252) <= inputs(71);
    layer0_outputs(3253) <= not(inputs(30));
    layer0_outputs(3254) <= not((inputs(182)) or (inputs(147)));
    layer0_outputs(3255) <= not((inputs(234)) or (inputs(144)));
    layer0_outputs(3256) <= not((inputs(8)) and (inputs(22)));
    layer0_outputs(3257) <= not(inputs(210));
    layer0_outputs(3258) <= inputs(68);
    layer0_outputs(3259) <= not((inputs(124)) or (inputs(26)));
    layer0_outputs(3260) <= not(inputs(45));
    layer0_outputs(3261) <= not((inputs(196)) or (inputs(230)));
    layer0_outputs(3262) <= not(inputs(88));
    layer0_outputs(3263) <= inputs(246);
    layer0_outputs(3264) <= inputs(118);
    layer0_outputs(3265) <= not(inputs(72));
    layer0_outputs(3266) <= (inputs(153)) or (inputs(127));
    layer0_outputs(3267) <= (inputs(3)) and not (inputs(255));
    layer0_outputs(3268) <= not((inputs(228)) or (inputs(102)));
    layer0_outputs(3269) <= (inputs(63)) xor (inputs(75));
    layer0_outputs(3270) <= (inputs(121)) and not (inputs(164));
    layer0_outputs(3271) <= not((inputs(135)) or (inputs(130)));
    layer0_outputs(3272) <= inputs(108);
    layer0_outputs(3273) <= inputs(8);
    layer0_outputs(3274) <= not(inputs(221));
    layer0_outputs(3275) <= not(inputs(36));
    layer0_outputs(3276) <= not(inputs(251));
    layer0_outputs(3277) <= (inputs(244)) xor (inputs(22));
    layer0_outputs(3278) <= not(inputs(122));
    layer0_outputs(3279) <= not(inputs(19));
    layer0_outputs(3280) <= not(inputs(33));
    layer0_outputs(3281) <= (inputs(10)) and not (inputs(65));
    layer0_outputs(3282) <= not((inputs(138)) or (inputs(30)));
    layer0_outputs(3283) <= not((inputs(177)) or (inputs(67)));
    layer0_outputs(3284) <= not(inputs(154)) or (inputs(116));
    layer0_outputs(3285) <= (inputs(107)) xor (inputs(67));
    layer0_outputs(3286) <= not((inputs(6)) xor (inputs(36)));
    layer0_outputs(3287) <= not((inputs(122)) or (inputs(14)));
    layer0_outputs(3288) <= inputs(157);
    layer0_outputs(3289) <= not(inputs(117));
    layer0_outputs(3290) <= (inputs(146)) and not (inputs(80));
    layer0_outputs(3291) <= inputs(66);
    layer0_outputs(3292) <= '0';
    layer0_outputs(3293) <= inputs(194);
    layer0_outputs(3294) <= not(inputs(212)) or (inputs(90));
    layer0_outputs(3295) <= inputs(185);
    layer0_outputs(3296) <= not((inputs(18)) or (inputs(211)));
    layer0_outputs(3297) <= not((inputs(134)) xor (inputs(101)));
    layer0_outputs(3298) <= (inputs(219)) xor (inputs(52));
    layer0_outputs(3299) <= (inputs(17)) xor (inputs(187));
    layer0_outputs(3300) <= not((inputs(1)) or (inputs(170)));
    layer0_outputs(3301) <= not((inputs(39)) xor (inputs(215)));
    layer0_outputs(3302) <= not(inputs(125));
    layer0_outputs(3303) <= (inputs(158)) or (inputs(100));
    layer0_outputs(3304) <= not((inputs(222)) or (inputs(228)));
    layer0_outputs(3305) <= (inputs(59)) and not (inputs(207));
    layer0_outputs(3306) <= not(inputs(83));
    layer0_outputs(3307) <= not((inputs(18)) or (inputs(31)));
    layer0_outputs(3308) <= not(inputs(84));
    layer0_outputs(3309) <= inputs(145);
    layer0_outputs(3310) <= (inputs(117)) xor (inputs(88));
    layer0_outputs(3311) <= (inputs(255)) or (inputs(198));
    layer0_outputs(3312) <= inputs(115);
    layer0_outputs(3313) <= not(inputs(231));
    layer0_outputs(3314) <= not(inputs(103)) or (inputs(94));
    layer0_outputs(3315) <= (inputs(155)) or (inputs(145));
    layer0_outputs(3316) <= not((inputs(5)) and (inputs(6)));
    layer0_outputs(3317) <= not(inputs(180)) or (inputs(41));
    layer0_outputs(3318) <= (inputs(173)) and not (inputs(169));
    layer0_outputs(3319) <= inputs(21);
    layer0_outputs(3320) <= not(inputs(137));
    layer0_outputs(3321) <= inputs(1);
    layer0_outputs(3322) <= not(inputs(83));
    layer0_outputs(3323) <= not(inputs(88)) or (inputs(79));
    layer0_outputs(3324) <= inputs(127);
    layer0_outputs(3325) <= (inputs(193)) and not (inputs(67));
    layer0_outputs(3326) <= (inputs(10)) and not (inputs(111));
    layer0_outputs(3327) <= not(inputs(58)) or (inputs(183));
    layer0_outputs(3328) <= inputs(166);
    layer0_outputs(3329) <= not(inputs(138));
    layer0_outputs(3330) <= (inputs(179)) or (inputs(109));
    layer0_outputs(3331) <= inputs(225);
    layer0_outputs(3332) <= (inputs(244)) or (inputs(249));
    layer0_outputs(3333) <= (inputs(177)) xor (inputs(216));
    layer0_outputs(3334) <= not(inputs(230));
    layer0_outputs(3335) <= not(inputs(15)) or (inputs(77));
    layer0_outputs(3336) <= not(inputs(233));
    layer0_outputs(3337) <= (inputs(99)) and not (inputs(174));
    layer0_outputs(3338) <= not(inputs(168));
    layer0_outputs(3339) <= not(inputs(163));
    layer0_outputs(3340) <= (inputs(219)) xor (inputs(208));
    layer0_outputs(3341) <= (inputs(129)) or (inputs(174));
    layer0_outputs(3342) <= (inputs(115)) xor (inputs(84));
    layer0_outputs(3343) <= (inputs(195)) or (inputs(196));
    layer0_outputs(3344) <= not(inputs(61));
    layer0_outputs(3345) <= not((inputs(182)) or (inputs(33)));
    layer0_outputs(3346) <= not(inputs(172)) or (inputs(236));
    layer0_outputs(3347) <= not((inputs(93)) xor (inputs(2)));
    layer0_outputs(3348) <= not((inputs(11)) or (inputs(249)));
    layer0_outputs(3349) <= not((inputs(138)) or (inputs(251)));
    layer0_outputs(3350) <= not(inputs(216)) or (inputs(239));
    layer0_outputs(3351) <= not(inputs(228)) or (inputs(42));
    layer0_outputs(3352) <= (inputs(33)) or (inputs(172));
    layer0_outputs(3353) <= (inputs(119)) xor (inputs(159));
    layer0_outputs(3354) <= inputs(101);
    layer0_outputs(3355) <= not(inputs(243));
    layer0_outputs(3356) <= inputs(123);
    layer0_outputs(3357) <= inputs(102);
    layer0_outputs(3358) <= (inputs(204)) and not (inputs(84));
    layer0_outputs(3359) <= not(inputs(15));
    layer0_outputs(3360) <= not(inputs(230));
    layer0_outputs(3361) <= not(inputs(227));
    layer0_outputs(3362) <= (inputs(180)) and not (inputs(165));
    layer0_outputs(3363) <= not((inputs(52)) xor (inputs(95)));
    layer0_outputs(3364) <= not((inputs(219)) xor (inputs(142)));
    layer0_outputs(3365) <= not(inputs(236)) or (inputs(149));
    layer0_outputs(3366) <= inputs(120);
    layer0_outputs(3367) <= not((inputs(214)) xor (inputs(46)));
    layer0_outputs(3368) <= not(inputs(68)) or (inputs(172));
    layer0_outputs(3369) <= inputs(135);
    layer0_outputs(3370) <= not((inputs(3)) or (inputs(21)));
    layer0_outputs(3371) <= not((inputs(120)) xor (inputs(187)));
    layer0_outputs(3372) <= (inputs(39)) and not (inputs(199));
    layer0_outputs(3373) <= not(inputs(3));
    layer0_outputs(3374) <= not(inputs(79)) or (inputs(78));
    layer0_outputs(3375) <= not((inputs(185)) xor (inputs(236)));
    layer0_outputs(3376) <= not(inputs(207)) or (inputs(191));
    layer0_outputs(3377) <= (inputs(226)) and not (inputs(129));
    layer0_outputs(3378) <= not(inputs(162));
    layer0_outputs(3379) <= not(inputs(22)) or (inputs(193));
    layer0_outputs(3380) <= (inputs(132)) and not (inputs(75));
    layer0_outputs(3381) <= (inputs(65)) or (inputs(12));
    layer0_outputs(3382) <= (inputs(248)) and not (inputs(118));
    layer0_outputs(3383) <= not((inputs(224)) or (inputs(232)));
    layer0_outputs(3384) <= (inputs(90)) or (inputs(4));
    layer0_outputs(3385) <= not(inputs(84)) or (inputs(206));
    layer0_outputs(3386) <= not(inputs(244));
    layer0_outputs(3387) <= '1';
    layer0_outputs(3388) <= not((inputs(160)) or (inputs(232)));
    layer0_outputs(3389) <= '1';
    layer0_outputs(3390) <= inputs(35);
    layer0_outputs(3391) <= not((inputs(243)) or (inputs(74)));
    layer0_outputs(3392) <= (inputs(152)) and not (inputs(46));
    layer0_outputs(3393) <= (inputs(83)) or (inputs(45));
    layer0_outputs(3394) <= not(inputs(83)) or (inputs(136));
    layer0_outputs(3395) <= (inputs(123)) and not (inputs(186));
    layer0_outputs(3396) <= not((inputs(42)) xor (inputs(143)));
    layer0_outputs(3397) <= not(inputs(170)) or (inputs(196));
    layer0_outputs(3398) <= not((inputs(201)) xor (inputs(234)));
    layer0_outputs(3399) <= not(inputs(13)) or (inputs(224));
    layer0_outputs(3400) <= not(inputs(195));
    layer0_outputs(3401) <= (inputs(127)) or (inputs(42));
    layer0_outputs(3402) <= inputs(59);
    layer0_outputs(3403) <= not(inputs(180));
    layer0_outputs(3404) <= (inputs(90)) and not (inputs(170));
    layer0_outputs(3405) <= (inputs(223)) and not (inputs(47));
    layer0_outputs(3406) <= not((inputs(53)) or (inputs(246)));
    layer0_outputs(3407) <= not((inputs(236)) xor (inputs(188)));
    layer0_outputs(3408) <= not((inputs(179)) or (inputs(158)));
    layer0_outputs(3409) <= inputs(230);
    layer0_outputs(3410) <= inputs(158);
    layer0_outputs(3411) <= (inputs(101)) and not (inputs(190));
    layer0_outputs(3412) <= not((inputs(232)) or (inputs(176)));
    layer0_outputs(3413) <= (inputs(102)) or (inputs(199));
    layer0_outputs(3414) <= not(inputs(93));
    layer0_outputs(3415) <= not(inputs(248));
    layer0_outputs(3416) <= not(inputs(6));
    layer0_outputs(3417) <= not((inputs(9)) or (inputs(171)));
    layer0_outputs(3418) <= (inputs(149)) and not (inputs(76));
    layer0_outputs(3419) <= (inputs(209)) and not (inputs(141));
    layer0_outputs(3420) <= (inputs(138)) or (inputs(184));
    layer0_outputs(3421) <= not(inputs(195)) or (inputs(112));
    layer0_outputs(3422) <= (inputs(2)) or (inputs(225));
    layer0_outputs(3423) <= not((inputs(161)) and (inputs(51)));
    layer0_outputs(3424) <= (inputs(104)) and not (inputs(170));
    layer0_outputs(3425) <= (inputs(169)) and not (inputs(79));
    layer0_outputs(3426) <= not(inputs(68));
    layer0_outputs(3427) <= (inputs(24)) xor (inputs(159));
    layer0_outputs(3428) <= '0';
    layer0_outputs(3429) <= inputs(106);
    layer0_outputs(3430) <= (inputs(195)) and not (inputs(255));
    layer0_outputs(3431) <= not((inputs(199)) and (inputs(179)));
    layer0_outputs(3432) <= not(inputs(93));
    layer0_outputs(3433) <= not(inputs(107)) or (inputs(37));
    layer0_outputs(3434) <= (inputs(70)) or (inputs(172));
    layer0_outputs(3435) <= inputs(58);
    layer0_outputs(3436) <= not((inputs(224)) and (inputs(86)));
    layer0_outputs(3437) <= not((inputs(68)) or (inputs(102)));
    layer0_outputs(3438) <= (inputs(171)) or (inputs(223));
    layer0_outputs(3439) <= not(inputs(134));
    layer0_outputs(3440) <= not(inputs(34));
    layer0_outputs(3441) <= not(inputs(199)) or (inputs(65));
    layer0_outputs(3442) <= not(inputs(101));
    layer0_outputs(3443) <= not(inputs(103));
    layer0_outputs(3444) <= not((inputs(66)) or (inputs(86)));
    layer0_outputs(3445) <= (inputs(240)) and (inputs(186));
    layer0_outputs(3446) <= (inputs(75)) or (inputs(135));
    layer0_outputs(3447) <= (inputs(205)) and not (inputs(126));
    layer0_outputs(3448) <= (inputs(8)) and not (inputs(208));
    layer0_outputs(3449) <= inputs(142);
    layer0_outputs(3450) <= (inputs(17)) or (inputs(60));
    layer0_outputs(3451) <= not(inputs(208)) or (inputs(12));
    layer0_outputs(3452) <= not(inputs(160)) or (inputs(158));
    layer0_outputs(3453) <= not((inputs(152)) or (inputs(219)));
    layer0_outputs(3454) <= inputs(121);
    layer0_outputs(3455) <= '1';
    layer0_outputs(3456) <= not(inputs(246));
    layer0_outputs(3457) <= (inputs(65)) and not (inputs(209));
    layer0_outputs(3458) <= not((inputs(101)) or (inputs(12)));
    layer0_outputs(3459) <= not(inputs(89)) or (inputs(216));
    layer0_outputs(3460) <= not((inputs(203)) xor (inputs(235)));
    layer0_outputs(3461) <= (inputs(217)) or (inputs(194));
    layer0_outputs(3462) <= not((inputs(247)) or (inputs(174)));
    layer0_outputs(3463) <= (inputs(19)) or (inputs(1));
    layer0_outputs(3464) <= not(inputs(11));
    layer0_outputs(3465) <= (inputs(78)) or (inputs(199));
    layer0_outputs(3466) <= inputs(20);
    layer0_outputs(3467) <= inputs(208);
    layer0_outputs(3468) <= inputs(157);
    layer0_outputs(3469) <= (inputs(169)) and not (inputs(152));
    layer0_outputs(3470) <= inputs(210);
    layer0_outputs(3471) <= (inputs(207)) or (inputs(251));
    layer0_outputs(3472) <= (inputs(224)) xor (inputs(64));
    layer0_outputs(3473) <= (inputs(21)) and not (inputs(162));
    layer0_outputs(3474) <= inputs(87);
    layer0_outputs(3475) <= (inputs(230)) and not (inputs(221));
    layer0_outputs(3476) <= not((inputs(211)) xor (inputs(118)));
    layer0_outputs(3477) <= (inputs(189)) or (inputs(193));
    layer0_outputs(3478) <= inputs(69);
    layer0_outputs(3479) <= (inputs(219)) or (inputs(185));
    layer0_outputs(3480) <= not(inputs(77));
    layer0_outputs(3481) <= not((inputs(70)) xor (inputs(89)));
    layer0_outputs(3482) <= (inputs(180)) xor (inputs(192));
    layer0_outputs(3483) <= not(inputs(169)) or (inputs(131));
    layer0_outputs(3484) <= not(inputs(231));
    layer0_outputs(3485) <= inputs(130);
    layer0_outputs(3486) <= not(inputs(100)) or (inputs(178));
    layer0_outputs(3487) <= not((inputs(219)) xor (inputs(186)));
    layer0_outputs(3488) <= inputs(214);
    layer0_outputs(3489) <= (inputs(87)) and not (inputs(180));
    layer0_outputs(3490) <= not(inputs(186));
    layer0_outputs(3491) <= not(inputs(46));
    layer0_outputs(3492) <= not(inputs(148));
    layer0_outputs(3493) <= not(inputs(237));
    layer0_outputs(3494) <= (inputs(198)) xor (inputs(185));
    layer0_outputs(3495) <= inputs(26);
    layer0_outputs(3496) <= not((inputs(237)) or (inputs(14)));
    layer0_outputs(3497) <= (inputs(212)) or (inputs(232));
    layer0_outputs(3498) <= not((inputs(170)) or (inputs(30)));
    layer0_outputs(3499) <= not(inputs(223));
    layer0_outputs(3500) <= not((inputs(181)) xor (inputs(158)));
    layer0_outputs(3501) <= (inputs(8)) xor (inputs(109));
    layer0_outputs(3502) <= not(inputs(137)) or (inputs(84));
    layer0_outputs(3503) <= (inputs(177)) or (inputs(248));
    layer0_outputs(3504) <= not((inputs(57)) xor (inputs(76)));
    layer0_outputs(3505) <= inputs(31);
    layer0_outputs(3506) <= not((inputs(53)) xor (inputs(88)));
    layer0_outputs(3507) <= not(inputs(144));
    layer0_outputs(3508) <= not((inputs(217)) or (inputs(38)));
    layer0_outputs(3509) <= not(inputs(179)) or (inputs(58));
    layer0_outputs(3510) <= (inputs(0)) or (inputs(255));
    layer0_outputs(3511) <= (inputs(1)) and not (inputs(140));
    layer0_outputs(3512) <= (inputs(119)) and (inputs(25));
    layer0_outputs(3513) <= (inputs(149)) and not (inputs(201));
    layer0_outputs(3514) <= inputs(37);
    layer0_outputs(3515) <= inputs(182);
    layer0_outputs(3516) <= (inputs(30)) xor (inputs(106));
    layer0_outputs(3517) <= (inputs(235)) xor (inputs(16));
    layer0_outputs(3518) <= not((inputs(135)) and (inputs(149)));
    layer0_outputs(3519) <= inputs(171);
    layer0_outputs(3520) <= inputs(116);
    layer0_outputs(3521) <= not((inputs(59)) or (inputs(135)));
    layer0_outputs(3522) <= (inputs(89)) or (inputs(6));
    layer0_outputs(3523) <= inputs(164);
    layer0_outputs(3524) <= inputs(164);
    layer0_outputs(3525) <= (inputs(72)) xor (inputs(117));
    layer0_outputs(3526) <= not((inputs(38)) and (inputs(214)));
    layer0_outputs(3527) <= not(inputs(98));
    layer0_outputs(3528) <= (inputs(0)) xor (inputs(196));
    layer0_outputs(3529) <= not((inputs(29)) or (inputs(71)));
    layer0_outputs(3530) <= inputs(93);
    layer0_outputs(3531) <= (inputs(182)) xor (inputs(212));
    layer0_outputs(3532) <= (inputs(196)) xor (inputs(38));
    layer0_outputs(3533) <= inputs(67);
    layer0_outputs(3534) <= (inputs(159)) xor (inputs(218));
    layer0_outputs(3535) <= inputs(1);
    layer0_outputs(3536) <= (inputs(44)) or (inputs(65));
    layer0_outputs(3537) <= inputs(2);
    layer0_outputs(3538) <= not((inputs(194)) or (inputs(208)));
    layer0_outputs(3539) <= '0';
    layer0_outputs(3540) <= inputs(150);
    layer0_outputs(3541) <= not(inputs(189));
    layer0_outputs(3542) <= not((inputs(18)) or (inputs(182)));
    layer0_outputs(3543) <= not(inputs(75));
    layer0_outputs(3544) <= (inputs(22)) and not (inputs(253));
    layer0_outputs(3545) <= (inputs(89)) and not (inputs(201));
    layer0_outputs(3546) <= not((inputs(168)) or (inputs(242)));
    layer0_outputs(3547) <= not((inputs(171)) or (inputs(149)));
    layer0_outputs(3548) <= not(inputs(250));
    layer0_outputs(3549) <= not((inputs(5)) or (inputs(26)));
    layer0_outputs(3550) <= (inputs(14)) or (inputs(47));
    layer0_outputs(3551) <= (inputs(118)) or (inputs(203));
    layer0_outputs(3552) <= inputs(4);
    layer0_outputs(3553) <= (inputs(57)) and not (inputs(239));
    layer0_outputs(3554) <= (inputs(28)) or (inputs(116));
    layer0_outputs(3555) <= not(inputs(210)) or (inputs(255));
    layer0_outputs(3556) <= not((inputs(113)) or (inputs(192)));
    layer0_outputs(3557) <= not((inputs(31)) or (inputs(27)));
    layer0_outputs(3558) <= (inputs(41)) or (inputs(111));
    layer0_outputs(3559) <= not(inputs(243)) or (inputs(81));
    layer0_outputs(3560) <= (inputs(35)) xor (inputs(24));
    layer0_outputs(3561) <= not(inputs(197));
    layer0_outputs(3562) <= not((inputs(75)) or (inputs(15)));
    layer0_outputs(3563) <= not((inputs(52)) or (inputs(101)));
    layer0_outputs(3564) <= not(inputs(150));
    layer0_outputs(3565) <= (inputs(238)) or (inputs(192));
    layer0_outputs(3566) <= not((inputs(138)) xor (inputs(152)));
    layer0_outputs(3567) <= (inputs(183)) and (inputs(198));
    layer0_outputs(3568) <= (inputs(246)) and not (inputs(126));
    layer0_outputs(3569) <= not(inputs(139)) or (inputs(74));
    layer0_outputs(3570) <= (inputs(209)) and not (inputs(208));
    layer0_outputs(3571) <= '0';
    layer0_outputs(3572) <= (inputs(189)) and not (inputs(221));
    layer0_outputs(3573) <= not(inputs(142)) or (inputs(109));
    layer0_outputs(3574) <= (inputs(62)) and not (inputs(241));
    layer0_outputs(3575) <= not((inputs(235)) and (inputs(107)));
    layer0_outputs(3576) <= not((inputs(64)) xor (inputs(174)));
    layer0_outputs(3577) <= (inputs(186)) xor (inputs(197));
    layer0_outputs(3578) <= (inputs(69)) and not (inputs(202));
    layer0_outputs(3579) <= not((inputs(201)) xor (inputs(89)));
    layer0_outputs(3580) <= '1';
    layer0_outputs(3581) <= not(inputs(6));
    layer0_outputs(3582) <= not((inputs(73)) or (inputs(45)));
    layer0_outputs(3583) <= not((inputs(1)) xor (inputs(105)));
    layer0_outputs(3584) <= not(inputs(77)) or (inputs(201));
    layer0_outputs(3585) <= (inputs(125)) or (inputs(37));
    layer0_outputs(3586) <= (inputs(243)) or (inputs(240));
    layer0_outputs(3587) <= inputs(23);
    layer0_outputs(3588) <= (inputs(111)) or (inputs(182));
    layer0_outputs(3589) <= not(inputs(186)) or (inputs(91));
    layer0_outputs(3590) <= '0';
    layer0_outputs(3591) <= (inputs(197)) and not (inputs(241));
    layer0_outputs(3592) <= not(inputs(175));
    layer0_outputs(3593) <= not((inputs(217)) or (inputs(163)));
    layer0_outputs(3594) <= (inputs(76)) and (inputs(120));
    layer0_outputs(3595) <= inputs(101);
    layer0_outputs(3596) <= (inputs(193)) xor (inputs(181));
    layer0_outputs(3597) <= not(inputs(209));
    layer0_outputs(3598) <= inputs(105);
    layer0_outputs(3599) <= not(inputs(149)) or (inputs(152));
    layer0_outputs(3600) <= (inputs(107)) or (inputs(52));
    layer0_outputs(3601) <= (inputs(254)) or (inputs(131));
    layer0_outputs(3602) <= (inputs(13)) xor (inputs(209));
    layer0_outputs(3603) <= (inputs(168)) and not (inputs(27));
    layer0_outputs(3604) <= not(inputs(110));
    layer0_outputs(3605) <= not(inputs(134)) or (inputs(204));
    layer0_outputs(3606) <= (inputs(232)) and not (inputs(115));
    layer0_outputs(3607) <= not(inputs(41));
    layer0_outputs(3608) <= not(inputs(21));
    layer0_outputs(3609) <= (inputs(234)) or (inputs(16));
    layer0_outputs(3610) <= (inputs(241)) or (inputs(35));
    layer0_outputs(3611) <= not(inputs(70));
    layer0_outputs(3612) <= not(inputs(167)) or (inputs(41));
    layer0_outputs(3613) <= (inputs(58)) and not (inputs(251));
    layer0_outputs(3614) <= inputs(234);
    layer0_outputs(3615) <= inputs(167);
    layer0_outputs(3616) <= '0';
    layer0_outputs(3617) <= (inputs(164)) xor (inputs(111));
    layer0_outputs(3618) <= (inputs(9)) or (inputs(63));
    layer0_outputs(3619) <= '1';
    layer0_outputs(3620) <= inputs(134);
    layer0_outputs(3621) <= (inputs(193)) and not (inputs(26));
    layer0_outputs(3622) <= not(inputs(252)) or (inputs(64));
    layer0_outputs(3623) <= not((inputs(116)) xor (inputs(16)));
    layer0_outputs(3624) <= not(inputs(243));
    layer0_outputs(3625) <= not(inputs(151));
    layer0_outputs(3626) <= inputs(121);
    layer0_outputs(3627) <= not((inputs(115)) xor (inputs(243)));
    layer0_outputs(3628) <= '1';
    layer0_outputs(3629) <= (inputs(189)) or (inputs(213));
    layer0_outputs(3630) <= not(inputs(52)) or (inputs(176));
    layer0_outputs(3631) <= inputs(146);
    layer0_outputs(3632) <= not(inputs(152));
    layer0_outputs(3633) <= not((inputs(174)) and (inputs(189)));
    layer0_outputs(3634) <= inputs(248);
    layer0_outputs(3635) <= inputs(150);
    layer0_outputs(3636) <= (inputs(34)) xor (inputs(143));
    layer0_outputs(3637) <= not((inputs(76)) or (inputs(105)));
    layer0_outputs(3638) <= (inputs(33)) or (inputs(219));
    layer0_outputs(3639) <= not(inputs(25));
    layer0_outputs(3640) <= (inputs(134)) and not (inputs(166));
    layer0_outputs(3641) <= not(inputs(19));
    layer0_outputs(3642) <= not((inputs(219)) or (inputs(173)));
    layer0_outputs(3643) <= not((inputs(147)) or (inputs(8)));
    layer0_outputs(3644) <= '0';
    layer0_outputs(3645) <= (inputs(6)) or (inputs(222));
    layer0_outputs(3646) <= (inputs(33)) and not (inputs(112));
    layer0_outputs(3647) <= not(inputs(17));
    layer0_outputs(3648) <= (inputs(27)) and not (inputs(172));
    layer0_outputs(3649) <= not((inputs(168)) xor (inputs(242)));
    layer0_outputs(3650) <= (inputs(123)) and not (inputs(207));
    layer0_outputs(3651) <= (inputs(48)) or (inputs(235));
    layer0_outputs(3652) <= inputs(30);
    layer0_outputs(3653) <= (inputs(103)) and not (inputs(157));
    layer0_outputs(3654) <= (inputs(85)) and not (inputs(56));
    layer0_outputs(3655) <= not(inputs(253)) or (inputs(78));
    layer0_outputs(3656) <= (inputs(209)) and not (inputs(121));
    layer0_outputs(3657) <= (inputs(212)) or (inputs(132));
    layer0_outputs(3658) <= (inputs(156)) or (inputs(62));
    layer0_outputs(3659) <= not((inputs(181)) xor (inputs(229)));
    layer0_outputs(3660) <= not((inputs(58)) or (inputs(62)));
    layer0_outputs(3661) <= not(inputs(164)) or (inputs(36));
    layer0_outputs(3662) <= not((inputs(48)) or (inputs(1)));
    layer0_outputs(3663) <= '0';
    layer0_outputs(3664) <= (inputs(222)) xor (inputs(2));
    layer0_outputs(3665) <= (inputs(190)) xor (inputs(242));
    layer0_outputs(3666) <= not(inputs(176));
    layer0_outputs(3667) <= (inputs(47)) and not (inputs(236));
    layer0_outputs(3668) <= inputs(182);
    layer0_outputs(3669) <= inputs(84);
    layer0_outputs(3670) <= (inputs(50)) and not (inputs(236));
    layer0_outputs(3671) <= (inputs(203)) and (inputs(152));
    layer0_outputs(3672) <= not((inputs(160)) or (inputs(214)));
    layer0_outputs(3673) <= (inputs(122)) and not (inputs(214));
    layer0_outputs(3674) <= inputs(175);
    layer0_outputs(3675) <= not(inputs(185));
    layer0_outputs(3676) <= (inputs(23)) or (inputs(190));
    layer0_outputs(3677) <= not(inputs(13));
    layer0_outputs(3678) <= not((inputs(176)) or (inputs(164)));
    layer0_outputs(3679) <= not(inputs(105));
    layer0_outputs(3680) <= (inputs(219)) and not (inputs(207));
    layer0_outputs(3681) <= inputs(232);
    layer0_outputs(3682) <= not((inputs(177)) or (inputs(55)));
    layer0_outputs(3683) <= not(inputs(9));
    layer0_outputs(3684) <= not((inputs(210)) xor (inputs(174)));
    layer0_outputs(3685) <= not((inputs(169)) or (inputs(254)));
    layer0_outputs(3686) <= not(inputs(85));
    layer0_outputs(3687) <= (inputs(171)) or (inputs(217));
    layer0_outputs(3688) <= (inputs(186)) or (inputs(203));
    layer0_outputs(3689) <= not(inputs(184));
    layer0_outputs(3690) <= not((inputs(72)) xor (inputs(51)));
    layer0_outputs(3691) <= not((inputs(240)) xor (inputs(127)));
    layer0_outputs(3692) <= not(inputs(153)) or (inputs(225));
    layer0_outputs(3693) <= not((inputs(25)) or (inputs(17)));
    layer0_outputs(3694) <= not((inputs(254)) xor (inputs(21)));
    layer0_outputs(3695) <= not(inputs(193));
    layer0_outputs(3696) <= not(inputs(231)) or (inputs(90));
    layer0_outputs(3697) <= inputs(156);
    layer0_outputs(3698) <= (inputs(197)) and not (inputs(28));
    layer0_outputs(3699) <= (inputs(98)) and not (inputs(191));
    layer0_outputs(3700) <= not(inputs(124));
    layer0_outputs(3701) <= (inputs(219)) or (inputs(6));
    layer0_outputs(3702) <= not(inputs(102));
    layer0_outputs(3703) <= inputs(161);
    layer0_outputs(3704) <= not((inputs(140)) xor (inputs(154)));
    layer0_outputs(3705) <= inputs(154);
    layer0_outputs(3706) <= not((inputs(212)) or (inputs(186)));
    layer0_outputs(3707) <= not(inputs(155)) or (inputs(163));
    layer0_outputs(3708) <= inputs(61);
    layer0_outputs(3709) <= inputs(81);
    layer0_outputs(3710) <= not(inputs(82));
    layer0_outputs(3711) <= (inputs(196)) or (inputs(182));
    layer0_outputs(3712) <= (inputs(139)) or (inputs(158));
    layer0_outputs(3713) <= not(inputs(248));
    layer0_outputs(3714) <= (inputs(229)) and not (inputs(3));
    layer0_outputs(3715) <= (inputs(206)) xor (inputs(127));
    layer0_outputs(3716) <= not(inputs(183)) or (inputs(225));
    layer0_outputs(3717) <= not((inputs(34)) and (inputs(142)));
    layer0_outputs(3718) <= (inputs(85)) and (inputs(85));
    layer0_outputs(3719) <= not(inputs(167));
    layer0_outputs(3720) <= not(inputs(68));
    layer0_outputs(3721) <= not(inputs(125));
    layer0_outputs(3722) <= not(inputs(43)) or (inputs(234));
    layer0_outputs(3723) <= (inputs(168)) and (inputs(247));
    layer0_outputs(3724) <= (inputs(3)) and not (inputs(252));
    layer0_outputs(3725) <= not(inputs(9));
    layer0_outputs(3726) <= (inputs(160)) xor (inputs(81));
    layer0_outputs(3727) <= not(inputs(25));
    layer0_outputs(3728) <= not((inputs(65)) or (inputs(7)));
    layer0_outputs(3729) <= (inputs(20)) xor (inputs(177));
    layer0_outputs(3730) <= (inputs(49)) or (inputs(199));
    layer0_outputs(3731) <= (inputs(196)) and not (inputs(191));
    layer0_outputs(3732) <= (inputs(246)) or (inputs(213));
    layer0_outputs(3733) <= not((inputs(9)) xor (inputs(161)));
    layer0_outputs(3734) <= (inputs(112)) or (inputs(248));
    layer0_outputs(3735) <= (inputs(56)) and (inputs(108));
    layer0_outputs(3736) <= (inputs(185)) or (inputs(123));
    layer0_outputs(3737) <= (inputs(194)) or (inputs(247));
    layer0_outputs(3738) <= (inputs(216)) and not (inputs(246));
    layer0_outputs(3739) <= not(inputs(44)) or (inputs(252));
    layer0_outputs(3740) <= inputs(236);
    layer0_outputs(3741) <= not((inputs(254)) or (inputs(62)));
    layer0_outputs(3742) <= (inputs(138)) xor (inputs(216));
    layer0_outputs(3743) <= not(inputs(60)) or (inputs(81));
    layer0_outputs(3744) <= not(inputs(112));
    layer0_outputs(3745) <= inputs(228);
    layer0_outputs(3746) <= inputs(15);
    layer0_outputs(3747) <= not(inputs(217));
    layer0_outputs(3748) <= (inputs(14)) xor (inputs(126));
    layer0_outputs(3749) <= not(inputs(250));
    layer0_outputs(3750) <= not(inputs(103));
    layer0_outputs(3751) <= inputs(129);
    layer0_outputs(3752) <= (inputs(41)) and not (inputs(66));
    layer0_outputs(3753) <= inputs(2);
    layer0_outputs(3754) <= (inputs(233)) and not (inputs(39));
    layer0_outputs(3755) <= not((inputs(38)) or (inputs(21)));
    layer0_outputs(3756) <= (inputs(149)) and not (inputs(74));
    layer0_outputs(3757) <= not(inputs(115)) or (inputs(206));
    layer0_outputs(3758) <= (inputs(38)) and not (inputs(145));
    layer0_outputs(3759) <= (inputs(28)) and not (inputs(205));
    layer0_outputs(3760) <= not((inputs(62)) xor (inputs(24)));
    layer0_outputs(3761) <= not((inputs(124)) xor (inputs(254)));
    layer0_outputs(3762) <= not((inputs(162)) or (inputs(191)));
    layer0_outputs(3763) <= (inputs(64)) or (inputs(174));
    layer0_outputs(3764) <= (inputs(229)) and not (inputs(15));
    layer0_outputs(3765) <= not((inputs(181)) or (inputs(79)));
    layer0_outputs(3766) <= not(inputs(49));
    layer0_outputs(3767) <= inputs(120);
    layer0_outputs(3768) <= (inputs(195)) and not (inputs(12));
    layer0_outputs(3769) <= not((inputs(211)) xor (inputs(157)));
    layer0_outputs(3770) <= inputs(168);
    layer0_outputs(3771) <= not(inputs(44));
    layer0_outputs(3772) <= not((inputs(255)) or (inputs(49)));
    layer0_outputs(3773) <= not((inputs(66)) xor (inputs(101)));
    layer0_outputs(3774) <= not((inputs(179)) or (inputs(98)));
    layer0_outputs(3775) <= (inputs(175)) or (inputs(79));
    layer0_outputs(3776) <= inputs(88);
    layer0_outputs(3777) <= not(inputs(102));
    layer0_outputs(3778) <= inputs(165);
    layer0_outputs(3779) <= (inputs(58)) and not (inputs(47));
    layer0_outputs(3780) <= not(inputs(101));
    layer0_outputs(3781) <= not((inputs(239)) or (inputs(117)));
    layer0_outputs(3782) <= (inputs(111)) or (inputs(214));
    layer0_outputs(3783) <= not((inputs(198)) or (inputs(243)));
    layer0_outputs(3784) <= '1';
    layer0_outputs(3785) <= (inputs(219)) or (inputs(238));
    layer0_outputs(3786) <= not(inputs(101)) or (inputs(6));
    layer0_outputs(3787) <= (inputs(56)) or (inputs(209));
    layer0_outputs(3788) <= not(inputs(249));
    layer0_outputs(3789) <= inputs(118);
    layer0_outputs(3790) <= (inputs(209)) or (inputs(217));
    layer0_outputs(3791) <= not((inputs(12)) or (inputs(246)));
    layer0_outputs(3792) <= not((inputs(103)) or (inputs(62)));
    layer0_outputs(3793) <= (inputs(182)) and not (inputs(143));
    layer0_outputs(3794) <= not(inputs(166));
    layer0_outputs(3795) <= '0';
    layer0_outputs(3796) <= not((inputs(137)) xor (inputs(151)));
    layer0_outputs(3797) <= inputs(204);
    layer0_outputs(3798) <= inputs(144);
    layer0_outputs(3799) <= inputs(24);
    layer0_outputs(3800) <= (inputs(154)) and (inputs(254));
    layer0_outputs(3801) <= (inputs(106)) and (inputs(26));
    layer0_outputs(3802) <= (inputs(240)) or (inputs(29));
    layer0_outputs(3803) <= inputs(86);
    layer0_outputs(3804) <= (inputs(21)) xor (inputs(80));
    layer0_outputs(3805) <= not(inputs(186)) or (inputs(168));
    layer0_outputs(3806) <= (inputs(58)) or (inputs(194));
    layer0_outputs(3807) <= not(inputs(213));
    layer0_outputs(3808) <= (inputs(167)) and not (inputs(235));
    layer0_outputs(3809) <= inputs(107);
    layer0_outputs(3810) <= not(inputs(3)) or (inputs(81));
    layer0_outputs(3811) <= inputs(142);
    layer0_outputs(3812) <= '1';
    layer0_outputs(3813) <= inputs(134);
    layer0_outputs(3814) <= not(inputs(98)) or (inputs(169));
    layer0_outputs(3815) <= not(inputs(221)) or (inputs(12));
    layer0_outputs(3816) <= inputs(99);
    layer0_outputs(3817) <= not((inputs(101)) xor (inputs(152)));
    layer0_outputs(3818) <= not(inputs(75)) or (inputs(112));
    layer0_outputs(3819) <= not(inputs(235));
    layer0_outputs(3820) <= not((inputs(237)) xor (inputs(64)));
    layer0_outputs(3821) <= not(inputs(95));
    layer0_outputs(3822) <= (inputs(159)) xor (inputs(34));
    layer0_outputs(3823) <= not(inputs(156)) or (inputs(137));
    layer0_outputs(3824) <= not((inputs(210)) and (inputs(171)));
    layer0_outputs(3825) <= not((inputs(107)) and (inputs(73)));
    layer0_outputs(3826) <= not((inputs(234)) or (inputs(143)));
    layer0_outputs(3827) <= (inputs(93)) and not (inputs(229));
    layer0_outputs(3828) <= inputs(25);
    layer0_outputs(3829) <= not(inputs(130));
    layer0_outputs(3830) <= not((inputs(144)) or (inputs(23)));
    layer0_outputs(3831) <= not((inputs(51)) xor (inputs(119)));
    layer0_outputs(3832) <= (inputs(74)) xor (inputs(2));
    layer0_outputs(3833) <= (inputs(208)) and not (inputs(162));
    layer0_outputs(3834) <= inputs(168);
    layer0_outputs(3835) <= (inputs(109)) and not (inputs(137));
    layer0_outputs(3836) <= not(inputs(248)) or (inputs(52));
    layer0_outputs(3837) <= inputs(40);
    layer0_outputs(3838) <= not(inputs(193));
    layer0_outputs(3839) <= (inputs(203)) or (inputs(207));
    layer0_outputs(3840) <= not((inputs(40)) xor (inputs(70)));
    layer0_outputs(3841) <= not((inputs(243)) and (inputs(241)));
    layer0_outputs(3842) <= not(inputs(219)) or (inputs(102));
    layer0_outputs(3843) <= (inputs(21)) and not (inputs(157));
    layer0_outputs(3844) <= (inputs(142)) and not (inputs(171));
    layer0_outputs(3845) <= (inputs(6)) and not (inputs(33));
    layer0_outputs(3846) <= not((inputs(255)) or (inputs(169)));
    layer0_outputs(3847) <= not((inputs(55)) or (inputs(223)));
    layer0_outputs(3848) <= not((inputs(221)) xor (inputs(236)));
    layer0_outputs(3849) <= not((inputs(21)) xor (inputs(150)));
    layer0_outputs(3850) <= (inputs(24)) and not (inputs(225));
    layer0_outputs(3851) <= not((inputs(244)) or (inputs(26)));
    layer0_outputs(3852) <= (inputs(43)) and not (inputs(19));
    layer0_outputs(3853) <= not(inputs(147));
    layer0_outputs(3854) <= not((inputs(15)) or (inputs(169)));
    layer0_outputs(3855) <= not(inputs(87));
    layer0_outputs(3856) <= not(inputs(248)) or (inputs(87));
    layer0_outputs(3857) <= inputs(122);
    layer0_outputs(3858) <= inputs(90);
    layer0_outputs(3859) <= not((inputs(128)) xor (inputs(22)));
    layer0_outputs(3860) <= not(inputs(116)) or (inputs(55));
    layer0_outputs(3861) <= not(inputs(94));
    layer0_outputs(3862) <= (inputs(218)) and not (inputs(32));
    layer0_outputs(3863) <= not(inputs(115));
    layer0_outputs(3864) <= not(inputs(247)) or (inputs(36));
    layer0_outputs(3865) <= inputs(194);
    layer0_outputs(3866) <= not((inputs(51)) xor (inputs(207)));
    layer0_outputs(3867) <= (inputs(150)) xor (inputs(213));
    layer0_outputs(3868) <= (inputs(203)) and not (inputs(7));
    layer0_outputs(3869) <= (inputs(147)) or (inputs(102));
    layer0_outputs(3870) <= inputs(0);
    layer0_outputs(3871) <= not((inputs(234)) xor (inputs(161)));
    layer0_outputs(3872) <= (inputs(92)) and not (inputs(239));
    layer0_outputs(3873) <= (inputs(134)) and (inputs(60));
    layer0_outputs(3874) <= not((inputs(206)) or (inputs(203)));
    layer0_outputs(3875) <= not((inputs(124)) xor (inputs(89)));
    layer0_outputs(3876) <= not((inputs(71)) xor (inputs(254)));
    layer0_outputs(3877) <= not((inputs(67)) and (inputs(8)));
    layer0_outputs(3878) <= inputs(50);
    layer0_outputs(3879) <= '1';
    layer0_outputs(3880) <= (inputs(128)) xor (inputs(172));
    layer0_outputs(3881) <= not((inputs(84)) xor (inputs(9)));
    layer0_outputs(3882) <= not(inputs(137));
    layer0_outputs(3883) <= (inputs(152)) and (inputs(74));
    layer0_outputs(3884) <= not((inputs(110)) xor (inputs(221)));
    layer0_outputs(3885) <= not(inputs(233));
    layer0_outputs(3886) <= (inputs(93)) or (inputs(51));
    layer0_outputs(3887) <= inputs(19);
    layer0_outputs(3888) <= not(inputs(163));
    layer0_outputs(3889) <= inputs(75);
    layer0_outputs(3890) <= not((inputs(131)) or (inputs(203)));
    layer0_outputs(3891) <= (inputs(205)) or (inputs(252));
    layer0_outputs(3892) <= (inputs(67)) or (inputs(185));
    layer0_outputs(3893) <= not(inputs(230)) or (inputs(33));
    layer0_outputs(3894) <= not((inputs(213)) and (inputs(202)));
    layer0_outputs(3895) <= not(inputs(8));
    layer0_outputs(3896) <= inputs(211);
    layer0_outputs(3897) <= not((inputs(52)) or (inputs(37)));
    layer0_outputs(3898) <= (inputs(92)) and not (inputs(238));
    layer0_outputs(3899) <= inputs(110);
    layer0_outputs(3900) <= not(inputs(130));
    layer0_outputs(3901) <= not(inputs(232)) or (inputs(14));
    layer0_outputs(3902) <= not(inputs(68)) or (inputs(16));
    layer0_outputs(3903) <= not((inputs(135)) or (inputs(199)));
    layer0_outputs(3904) <= not(inputs(121));
    layer0_outputs(3905) <= not(inputs(102));
    layer0_outputs(3906) <= not(inputs(128)) or (inputs(238));
    layer0_outputs(3907) <= inputs(221);
    layer0_outputs(3908) <= (inputs(171)) xor (inputs(135));
    layer0_outputs(3909) <= (inputs(141)) xor (inputs(108));
    layer0_outputs(3910) <= (inputs(21)) xor (inputs(175));
    layer0_outputs(3911) <= inputs(55);
    layer0_outputs(3912) <= (inputs(95)) xor (inputs(135));
    layer0_outputs(3913) <= (inputs(130)) or (inputs(34));
    layer0_outputs(3914) <= (inputs(91)) and not (inputs(119));
    layer0_outputs(3915) <= not(inputs(124));
    layer0_outputs(3916) <= inputs(224);
    layer0_outputs(3917) <= (inputs(218)) or (inputs(216));
    layer0_outputs(3918) <= inputs(106);
    layer0_outputs(3919) <= not((inputs(116)) xor (inputs(188)));
    layer0_outputs(3920) <= not(inputs(19));
    layer0_outputs(3921) <= (inputs(194)) and (inputs(138));
    layer0_outputs(3922) <= inputs(249);
    layer0_outputs(3923) <= inputs(166);
    layer0_outputs(3924) <= (inputs(12)) and not (inputs(109));
    layer0_outputs(3925) <= not(inputs(103));
    layer0_outputs(3926) <= inputs(147);
    layer0_outputs(3927) <= not(inputs(69)) or (inputs(116));
    layer0_outputs(3928) <= inputs(19);
    layer0_outputs(3929) <= not((inputs(196)) or (inputs(166)));
    layer0_outputs(3930) <= '1';
    layer0_outputs(3931) <= (inputs(135)) and (inputs(199));
    layer0_outputs(3932) <= inputs(52);
    layer0_outputs(3933) <= not(inputs(28)) or (inputs(207));
    layer0_outputs(3934) <= (inputs(135)) and not (inputs(185));
    layer0_outputs(3935) <= not(inputs(220));
    layer0_outputs(3936) <= (inputs(110)) xor (inputs(32));
    layer0_outputs(3937) <= not((inputs(226)) or (inputs(146)));
    layer0_outputs(3938) <= inputs(56);
    layer0_outputs(3939) <= (inputs(237)) or (inputs(150));
    layer0_outputs(3940) <= not((inputs(122)) or (inputs(163)));
    layer0_outputs(3941) <= (inputs(95)) and (inputs(37));
    layer0_outputs(3942) <= inputs(194);
    layer0_outputs(3943) <= not((inputs(65)) xor (inputs(70)));
    layer0_outputs(3944) <= (inputs(19)) or (inputs(73));
    layer0_outputs(3945) <= (inputs(59)) or (inputs(67));
    layer0_outputs(3946) <= not((inputs(93)) or (inputs(4)));
    layer0_outputs(3947) <= inputs(52);
    layer0_outputs(3948) <= not((inputs(175)) or (inputs(2)));
    layer0_outputs(3949) <= inputs(63);
    layer0_outputs(3950) <= (inputs(0)) or (inputs(71));
    layer0_outputs(3951) <= inputs(182);
    layer0_outputs(3952) <= (inputs(16)) or (inputs(173));
    layer0_outputs(3953) <= inputs(155);
    layer0_outputs(3954) <= not(inputs(61)) or (inputs(149));
    layer0_outputs(3955) <= (inputs(100)) or (inputs(141));
    layer0_outputs(3956) <= (inputs(39)) or (inputs(221));
    layer0_outputs(3957) <= inputs(219);
    layer0_outputs(3958) <= inputs(225);
    layer0_outputs(3959) <= not((inputs(213)) or (inputs(24)));
    layer0_outputs(3960) <= (inputs(9)) and not (inputs(128));
    layer0_outputs(3961) <= not(inputs(149)) or (inputs(143));
    layer0_outputs(3962) <= (inputs(41)) and not (inputs(194));
    layer0_outputs(3963) <= not(inputs(174));
    layer0_outputs(3964) <= '0';
    layer0_outputs(3965) <= not(inputs(168)) or (inputs(241));
    layer0_outputs(3966) <= inputs(85);
    layer0_outputs(3967) <= (inputs(59)) and not (inputs(193));
    layer0_outputs(3968) <= (inputs(22)) or (inputs(55));
    layer0_outputs(3969) <= (inputs(164)) xor (inputs(203));
    layer0_outputs(3970) <= '0';
    layer0_outputs(3971) <= inputs(125);
    layer0_outputs(3972) <= (inputs(161)) or (inputs(146));
    layer0_outputs(3973) <= not(inputs(178));
    layer0_outputs(3974) <= not(inputs(69)) or (inputs(161));
    layer0_outputs(3975) <= (inputs(217)) and not (inputs(34));
    layer0_outputs(3976) <= (inputs(254)) or (inputs(224));
    layer0_outputs(3977) <= not((inputs(24)) or (inputs(33)));
    layer0_outputs(3978) <= inputs(106);
    layer0_outputs(3979) <= not((inputs(238)) or (inputs(109)));
    layer0_outputs(3980) <= not((inputs(67)) or (inputs(174)));
    layer0_outputs(3981) <= not((inputs(26)) xor (inputs(60)));
    layer0_outputs(3982) <= not((inputs(159)) or (inputs(199)));
    layer0_outputs(3983) <= inputs(213);
    layer0_outputs(3984) <= not((inputs(131)) xor (inputs(175)));
    layer0_outputs(3985) <= inputs(173);
    layer0_outputs(3986) <= (inputs(234)) or (inputs(232));
    layer0_outputs(3987) <= not(inputs(24));
    layer0_outputs(3988) <= (inputs(104)) and (inputs(166));
    layer0_outputs(3989) <= inputs(39);
    layer0_outputs(3990) <= not((inputs(37)) xor (inputs(0)));
    layer0_outputs(3991) <= not(inputs(117)) or (inputs(50));
    layer0_outputs(3992) <= (inputs(98)) or (inputs(28));
    layer0_outputs(3993) <= inputs(25);
    layer0_outputs(3994) <= (inputs(6)) and not (inputs(159));
    layer0_outputs(3995) <= (inputs(12)) and (inputs(69));
    layer0_outputs(3996) <= (inputs(55)) and not (inputs(255));
    layer0_outputs(3997) <= not(inputs(74)) or (inputs(169));
    layer0_outputs(3998) <= (inputs(131)) xor (inputs(165));
    layer0_outputs(3999) <= inputs(93);
    layer0_outputs(4000) <= not((inputs(244)) and (inputs(178)));
    layer0_outputs(4001) <= not((inputs(41)) xor (inputs(234)));
    layer0_outputs(4002) <= not((inputs(74)) and (inputs(205)));
    layer0_outputs(4003) <= not(inputs(169));
    layer0_outputs(4004) <= inputs(99);
    layer0_outputs(4005) <= not(inputs(87));
    layer0_outputs(4006) <= not(inputs(115)) or (inputs(46));
    layer0_outputs(4007) <= not((inputs(48)) or (inputs(186)));
    layer0_outputs(4008) <= (inputs(7)) or (inputs(83));
    layer0_outputs(4009) <= (inputs(26)) and not (inputs(147));
    layer0_outputs(4010) <= inputs(211);
    layer0_outputs(4011) <= inputs(91);
    layer0_outputs(4012) <= not(inputs(80));
    layer0_outputs(4013) <= not((inputs(12)) or (inputs(62)));
    layer0_outputs(4014) <= not((inputs(231)) or (inputs(191)));
    layer0_outputs(4015) <= not((inputs(143)) xor (inputs(180)));
    layer0_outputs(4016) <= '1';
    layer0_outputs(4017) <= not((inputs(209)) or (inputs(82)));
    layer0_outputs(4018) <= inputs(223);
    layer0_outputs(4019) <= not(inputs(44));
    layer0_outputs(4020) <= (inputs(186)) or (inputs(19));
    layer0_outputs(4021) <= inputs(46);
    layer0_outputs(4022) <= inputs(100);
    layer0_outputs(4023) <= (inputs(53)) and not (inputs(250));
    layer0_outputs(4024) <= not((inputs(22)) or (inputs(246)));
    layer0_outputs(4025) <= inputs(98);
    layer0_outputs(4026) <= inputs(167);
    layer0_outputs(4027) <= (inputs(159)) or (inputs(235));
    layer0_outputs(4028) <= not(inputs(61));
    layer0_outputs(4029) <= not(inputs(184));
    layer0_outputs(4030) <= inputs(151);
    layer0_outputs(4031) <= inputs(65);
    layer0_outputs(4032) <= '0';
    layer0_outputs(4033) <= not(inputs(241)) or (inputs(78));
    layer0_outputs(4034) <= (inputs(5)) or (inputs(131));
    layer0_outputs(4035) <= inputs(153);
    layer0_outputs(4036) <= not((inputs(165)) xor (inputs(123)));
    layer0_outputs(4037) <= inputs(146);
    layer0_outputs(4038) <= not((inputs(133)) or (inputs(242)));
    layer0_outputs(4039) <= (inputs(223)) and (inputs(100));
    layer0_outputs(4040) <= not((inputs(131)) xor (inputs(20)));
    layer0_outputs(4041) <= (inputs(69)) xor (inputs(82));
    layer0_outputs(4042) <= (inputs(227)) or (inputs(173));
    layer0_outputs(4043) <= inputs(94);
    layer0_outputs(4044) <= not(inputs(172));
    layer0_outputs(4045) <= (inputs(68)) and not (inputs(244));
    layer0_outputs(4046) <= not((inputs(188)) and (inputs(94)));
    layer0_outputs(4047) <= inputs(19);
    layer0_outputs(4048) <= (inputs(167)) or (inputs(5));
    layer0_outputs(4049) <= (inputs(190)) and not (inputs(26));
    layer0_outputs(4050) <= inputs(14);
    layer0_outputs(4051) <= not(inputs(133));
    layer0_outputs(4052) <= inputs(146);
    layer0_outputs(4053) <= not((inputs(11)) or (inputs(50)));
    layer0_outputs(4054) <= not((inputs(72)) and (inputs(226)));
    layer0_outputs(4055) <= inputs(76);
    layer0_outputs(4056) <= (inputs(248)) xor (inputs(105));
    layer0_outputs(4057) <= (inputs(27)) and not (inputs(209));
    layer0_outputs(4058) <= not((inputs(201)) and (inputs(227)));
    layer0_outputs(4059) <= (inputs(249)) or (inputs(150));
    layer0_outputs(4060) <= (inputs(9)) or (inputs(172));
    layer0_outputs(4061) <= (inputs(20)) xor (inputs(156));
    layer0_outputs(4062) <= (inputs(126)) and not (inputs(131));
    layer0_outputs(4063) <= not(inputs(141));
    layer0_outputs(4064) <= not((inputs(225)) or (inputs(247)));
    layer0_outputs(4065) <= not(inputs(105));
    layer0_outputs(4066) <= not((inputs(135)) and (inputs(85)));
    layer0_outputs(4067) <= (inputs(104)) xor (inputs(59));
    layer0_outputs(4068) <= (inputs(154)) and not (inputs(15));
    layer0_outputs(4069) <= not((inputs(140)) and (inputs(12)));
    layer0_outputs(4070) <= (inputs(52)) xor (inputs(48));
    layer0_outputs(4071) <= not(inputs(188));
    layer0_outputs(4072) <= (inputs(158)) and not (inputs(255));
    layer0_outputs(4073) <= (inputs(20)) or (inputs(226));
    layer0_outputs(4074) <= inputs(20);
    layer0_outputs(4075) <= not(inputs(22));
    layer0_outputs(4076) <= not((inputs(151)) and (inputs(136)));
    layer0_outputs(4077) <= not((inputs(40)) xor (inputs(69)));
    layer0_outputs(4078) <= not(inputs(177)) or (inputs(240));
    layer0_outputs(4079) <= not(inputs(218));
    layer0_outputs(4080) <= (inputs(214)) and not (inputs(203));
    layer0_outputs(4081) <= inputs(182);
    layer0_outputs(4082) <= inputs(147);
    layer0_outputs(4083) <= not(inputs(23));
    layer0_outputs(4084) <= (inputs(190)) and not (inputs(65));
    layer0_outputs(4085) <= (inputs(103)) xor (inputs(14));
    layer0_outputs(4086) <= not((inputs(244)) or (inputs(228)));
    layer0_outputs(4087) <= not((inputs(19)) or (inputs(78)));
    layer0_outputs(4088) <= (inputs(38)) and not (inputs(92));
    layer0_outputs(4089) <= not((inputs(111)) or (inputs(53)));
    layer0_outputs(4090) <= not((inputs(72)) xor (inputs(181)));
    layer0_outputs(4091) <= not((inputs(230)) or (inputs(68)));
    layer0_outputs(4092) <= inputs(148);
    layer0_outputs(4093) <= not(inputs(212));
    layer0_outputs(4094) <= not((inputs(47)) or (inputs(73)));
    layer0_outputs(4095) <= (inputs(216)) and not (inputs(128));
    layer0_outputs(4096) <= not(inputs(77));
    layer0_outputs(4097) <= (inputs(56)) and (inputs(207));
    layer0_outputs(4098) <= (inputs(85)) and not (inputs(47));
    layer0_outputs(4099) <= (inputs(186)) and not (inputs(207));
    layer0_outputs(4100) <= (inputs(231)) xor (inputs(105));
    layer0_outputs(4101) <= not((inputs(135)) xor (inputs(122)));
    layer0_outputs(4102) <= not(inputs(74)) or (inputs(196));
    layer0_outputs(4103) <= inputs(57);
    layer0_outputs(4104) <= (inputs(9)) and (inputs(129));
    layer0_outputs(4105) <= not((inputs(117)) xor (inputs(34)));
    layer0_outputs(4106) <= not(inputs(105)) or (inputs(208));
    layer0_outputs(4107) <= not((inputs(11)) and (inputs(134)));
    layer0_outputs(4108) <= not((inputs(193)) or (inputs(9)));
    layer0_outputs(4109) <= (inputs(114)) and not (inputs(252));
    layer0_outputs(4110) <= not(inputs(77));
    layer0_outputs(4111) <= not((inputs(119)) xor (inputs(169)));
    layer0_outputs(4112) <= not(inputs(21));
    layer0_outputs(4113) <= not(inputs(39));
    layer0_outputs(4114) <= not(inputs(144));
    layer0_outputs(4115) <= not(inputs(149));
    layer0_outputs(4116) <= not((inputs(35)) or (inputs(210)));
    layer0_outputs(4117) <= (inputs(51)) or (inputs(37));
    layer0_outputs(4118) <= inputs(249);
    layer0_outputs(4119) <= (inputs(56)) or (inputs(57));
    layer0_outputs(4120) <= not(inputs(220));
    layer0_outputs(4121) <= inputs(117);
    layer0_outputs(4122) <= (inputs(97)) and not (inputs(175));
    layer0_outputs(4123) <= not(inputs(206));
    layer0_outputs(4124) <= not((inputs(42)) xor (inputs(17)));
    layer0_outputs(4125) <= (inputs(217)) and (inputs(0));
    layer0_outputs(4126) <= inputs(163);
    layer0_outputs(4127) <= (inputs(220)) and not (inputs(110));
    layer0_outputs(4128) <= (inputs(183)) or (inputs(32));
    layer0_outputs(4129) <= not(inputs(140)) or (inputs(3));
    layer0_outputs(4130) <= inputs(220);
    layer0_outputs(4131) <= not((inputs(60)) xor (inputs(168)));
    layer0_outputs(4132) <= not(inputs(119));
    layer0_outputs(4133) <= not(inputs(124));
    layer0_outputs(4134) <= not(inputs(163));
    layer0_outputs(4135) <= not(inputs(74)) or (inputs(203));
    layer0_outputs(4136) <= not(inputs(11)) or (inputs(214));
    layer0_outputs(4137) <= (inputs(215)) xor (inputs(94));
    layer0_outputs(4138) <= (inputs(177)) or (inputs(182));
    layer0_outputs(4139) <= (inputs(205)) or (inputs(211));
    layer0_outputs(4140) <= inputs(26);
    layer0_outputs(4141) <= not(inputs(237));
    layer0_outputs(4142) <= not((inputs(155)) xor (inputs(138)));
    layer0_outputs(4143) <= (inputs(105)) or (inputs(84));
    layer0_outputs(4144) <= (inputs(243)) xor (inputs(17));
    layer0_outputs(4145) <= inputs(230);
    layer0_outputs(4146) <= not((inputs(165)) xor (inputs(189)));
    layer0_outputs(4147) <= inputs(252);
    layer0_outputs(4148) <= not((inputs(16)) or (inputs(122)));
    layer0_outputs(4149) <= not(inputs(229));
    layer0_outputs(4150) <= inputs(211);
    layer0_outputs(4151) <= inputs(101);
    layer0_outputs(4152) <= not((inputs(114)) xor (inputs(105)));
    layer0_outputs(4153) <= (inputs(73)) xor (inputs(210));
    layer0_outputs(4154) <= inputs(34);
    layer0_outputs(4155) <= not(inputs(123)) or (inputs(72));
    layer0_outputs(4156) <= not((inputs(90)) or (inputs(47)));
    layer0_outputs(4157) <= not(inputs(58));
    layer0_outputs(4158) <= not(inputs(42)) or (inputs(194));
    layer0_outputs(4159) <= not((inputs(128)) and (inputs(93)));
    layer0_outputs(4160) <= (inputs(121)) or (inputs(20));
    layer0_outputs(4161) <= not((inputs(149)) xor (inputs(97)));
    layer0_outputs(4162) <= not(inputs(195)) or (inputs(30));
    layer0_outputs(4163) <= not(inputs(126)) or (inputs(240));
    layer0_outputs(4164) <= inputs(18);
    layer0_outputs(4165) <= inputs(221);
    layer0_outputs(4166) <= not((inputs(195)) or (inputs(194)));
    layer0_outputs(4167) <= not(inputs(180));
    layer0_outputs(4168) <= not(inputs(183));
    layer0_outputs(4169) <= not(inputs(46)) or (inputs(223));
    layer0_outputs(4170) <= (inputs(77)) xor (inputs(92));
    layer0_outputs(4171) <= not(inputs(99)) or (inputs(68));
    layer0_outputs(4172) <= not((inputs(139)) or (inputs(63)));
    layer0_outputs(4173) <= (inputs(52)) or (inputs(241));
    layer0_outputs(4174) <= not(inputs(200)) or (inputs(94));
    layer0_outputs(4175) <= not((inputs(50)) and (inputs(76)));
    layer0_outputs(4176) <= (inputs(203)) and not (inputs(186));
    layer0_outputs(4177) <= inputs(152);
    layer0_outputs(4178) <= (inputs(142)) xor (inputs(102));
    layer0_outputs(4179) <= (inputs(175)) or (inputs(66));
    layer0_outputs(4180) <= not((inputs(102)) xor (inputs(203)));
    layer0_outputs(4181) <= not(inputs(211));
    layer0_outputs(4182) <= (inputs(78)) or (inputs(42));
    layer0_outputs(4183) <= not(inputs(167)) or (inputs(36));
    layer0_outputs(4184) <= not((inputs(192)) and (inputs(80)));
    layer0_outputs(4185) <= (inputs(32)) xor (inputs(53));
    layer0_outputs(4186) <= not((inputs(252)) or (inputs(115)));
    layer0_outputs(4187) <= inputs(211);
    layer0_outputs(4188) <= (inputs(136)) and not (inputs(1));
    layer0_outputs(4189) <= not((inputs(51)) xor (inputs(90)));
    layer0_outputs(4190) <= not(inputs(71)) or (inputs(188));
    layer0_outputs(4191) <= not((inputs(49)) or (inputs(88)));
    layer0_outputs(4192) <= (inputs(235)) or (inputs(136));
    layer0_outputs(4193) <= not(inputs(76)) or (inputs(195));
    layer0_outputs(4194) <= not(inputs(186));
    layer0_outputs(4195) <= not((inputs(249)) or (inputs(158)));
    layer0_outputs(4196) <= (inputs(81)) xor (inputs(5));
    layer0_outputs(4197) <= inputs(8);
    layer0_outputs(4198) <= not(inputs(203));
    layer0_outputs(4199) <= (inputs(116)) xor (inputs(129));
    layer0_outputs(4200) <= not(inputs(130));
    layer0_outputs(4201) <= not(inputs(221)) or (inputs(120));
    layer0_outputs(4202) <= (inputs(172)) and not (inputs(160));
    layer0_outputs(4203) <= not(inputs(150));
    layer0_outputs(4204) <= not((inputs(82)) or (inputs(8)));
    layer0_outputs(4205) <= not((inputs(64)) or (inputs(213)));
    layer0_outputs(4206) <= not((inputs(74)) xor (inputs(64)));
    layer0_outputs(4207) <= not(inputs(28)) or (inputs(58));
    layer0_outputs(4208) <= inputs(231);
    layer0_outputs(4209) <= not(inputs(173));
    layer0_outputs(4210) <= (inputs(83)) and not (inputs(176));
    layer0_outputs(4211) <= (inputs(99)) or (inputs(12));
    layer0_outputs(4212) <= not(inputs(204)) or (inputs(34));
    layer0_outputs(4213) <= inputs(184);
    layer0_outputs(4214) <= not(inputs(241)) or (inputs(179));
    layer0_outputs(4215) <= not((inputs(212)) or (inputs(168)));
    layer0_outputs(4216) <= not((inputs(108)) xor (inputs(104)));
    layer0_outputs(4217) <= not((inputs(55)) xor (inputs(52)));
    layer0_outputs(4218) <= inputs(95);
    layer0_outputs(4219) <= inputs(145);
    layer0_outputs(4220) <= not((inputs(0)) or (inputs(54)));
    layer0_outputs(4221) <= not((inputs(166)) xor (inputs(205)));
    layer0_outputs(4222) <= '1';
    layer0_outputs(4223) <= not(inputs(2));
    layer0_outputs(4224) <= not((inputs(216)) or (inputs(96)));
    layer0_outputs(4225) <= inputs(165);
    layer0_outputs(4226) <= inputs(127);
    layer0_outputs(4227) <= (inputs(54)) and not (inputs(166));
    layer0_outputs(4228) <= not(inputs(229));
    layer0_outputs(4229) <= not((inputs(10)) or (inputs(50)));
    layer0_outputs(4230) <= (inputs(29)) or (inputs(60));
    layer0_outputs(4231) <= (inputs(86)) xor (inputs(130));
    layer0_outputs(4232) <= (inputs(17)) xor (inputs(186));
    layer0_outputs(4233) <= inputs(35);
    layer0_outputs(4234) <= (inputs(215)) xor (inputs(215));
    layer0_outputs(4235) <= not(inputs(51));
    layer0_outputs(4236) <= (inputs(173)) and (inputs(231));
    layer0_outputs(4237) <= inputs(219);
    layer0_outputs(4238) <= (inputs(151)) and not (inputs(147));
    layer0_outputs(4239) <= (inputs(183)) or (inputs(48));
    layer0_outputs(4240) <= (inputs(185)) xor (inputs(65));
    layer0_outputs(4241) <= inputs(154);
    layer0_outputs(4242) <= '1';
    layer0_outputs(4243) <= not((inputs(194)) or (inputs(83)));
    layer0_outputs(4244) <= (inputs(116)) or (inputs(88));
    layer0_outputs(4245) <= inputs(132);
    layer0_outputs(4246) <= not(inputs(60));
    layer0_outputs(4247) <= (inputs(103)) xor (inputs(229));
    layer0_outputs(4248) <= inputs(214);
    layer0_outputs(4249) <= (inputs(186)) or (inputs(253));
    layer0_outputs(4250) <= not((inputs(178)) or (inputs(78)));
    layer0_outputs(4251) <= (inputs(249)) and not (inputs(169));
    layer0_outputs(4252) <= (inputs(35)) or (inputs(71));
    layer0_outputs(4253) <= (inputs(155)) and not (inputs(7));
    layer0_outputs(4254) <= not(inputs(100));
    layer0_outputs(4255) <= not((inputs(37)) or (inputs(30)));
    layer0_outputs(4256) <= not(inputs(165));
    layer0_outputs(4257) <= not((inputs(15)) xor (inputs(244)));
    layer0_outputs(4258) <= (inputs(218)) xor (inputs(20));
    layer0_outputs(4259) <= (inputs(81)) or (inputs(66));
    layer0_outputs(4260) <= not((inputs(45)) and (inputs(24)));
    layer0_outputs(4261) <= not((inputs(114)) xor (inputs(34)));
    layer0_outputs(4262) <= inputs(119);
    layer0_outputs(4263) <= not((inputs(175)) or (inputs(42)));
    layer0_outputs(4264) <= (inputs(155)) and (inputs(105));
    layer0_outputs(4265) <= not((inputs(106)) or (inputs(23)));
    layer0_outputs(4266) <= (inputs(226)) or (inputs(84));
    layer0_outputs(4267) <= (inputs(7)) and not (inputs(61));
    layer0_outputs(4268) <= (inputs(61)) or (inputs(237));
    layer0_outputs(4269) <= (inputs(10)) xor (inputs(255));
    layer0_outputs(4270) <= (inputs(174)) xor (inputs(239));
    layer0_outputs(4271) <= not((inputs(204)) or (inputs(118)));
    layer0_outputs(4272) <= not(inputs(78));
    layer0_outputs(4273) <= not((inputs(135)) xor (inputs(240)));
    layer0_outputs(4274) <= not((inputs(36)) xor (inputs(0)));
    layer0_outputs(4275) <= inputs(113);
    layer0_outputs(4276) <= not((inputs(137)) or (inputs(10)));
    layer0_outputs(4277) <= not((inputs(239)) or (inputs(248)));
    layer0_outputs(4278) <= not(inputs(141));
    layer0_outputs(4279) <= (inputs(169)) or (inputs(126));
    layer0_outputs(4280) <= not(inputs(233));
    layer0_outputs(4281) <= not(inputs(100));
    layer0_outputs(4282) <= not((inputs(66)) xor (inputs(139)));
    layer0_outputs(4283) <= not((inputs(114)) or (inputs(72)));
    layer0_outputs(4284) <= not((inputs(23)) xor (inputs(55)));
    layer0_outputs(4285) <= inputs(145);
    layer0_outputs(4286) <= (inputs(65)) xor (inputs(198));
    layer0_outputs(4287) <= '0';
    layer0_outputs(4288) <= not(inputs(66)) or (inputs(253));
    layer0_outputs(4289) <= not((inputs(233)) or (inputs(218)));
    layer0_outputs(4290) <= (inputs(98)) xor (inputs(36));
    layer0_outputs(4291) <= not((inputs(128)) xor (inputs(118)));
    layer0_outputs(4292) <= not(inputs(9)) or (inputs(210));
    layer0_outputs(4293) <= not((inputs(196)) or (inputs(97)));
    layer0_outputs(4294) <= (inputs(133)) and not (inputs(21));
    layer0_outputs(4295) <= inputs(30);
    layer0_outputs(4296) <= inputs(243);
    layer0_outputs(4297) <= '1';
    layer0_outputs(4298) <= (inputs(170)) and not (inputs(86));
    layer0_outputs(4299) <= inputs(24);
    layer0_outputs(4300) <= not((inputs(143)) and (inputs(201)));
    layer0_outputs(4301) <= (inputs(170)) xor (inputs(107));
    layer0_outputs(4302) <= not(inputs(5)) or (inputs(190));
    layer0_outputs(4303) <= not(inputs(117));
    layer0_outputs(4304) <= (inputs(208)) or (inputs(211));
    layer0_outputs(4305) <= inputs(51);
    layer0_outputs(4306) <= not(inputs(139)) or (inputs(27));
    layer0_outputs(4307) <= not(inputs(233)) or (inputs(56));
    layer0_outputs(4308) <= not((inputs(28)) or (inputs(5)));
    layer0_outputs(4309) <= (inputs(174)) and not (inputs(101));
    layer0_outputs(4310) <= (inputs(99)) and not (inputs(2));
    layer0_outputs(4311) <= (inputs(17)) or (inputs(147));
    layer0_outputs(4312) <= not((inputs(16)) xor (inputs(36)));
    layer0_outputs(4313) <= inputs(195);
    layer0_outputs(4314) <= not((inputs(222)) xor (inputs(116)));
    layer0_outputs(4315) <= not((inputs(245)) xor (inputs(95)));
    layer0_outputs(4316) <= (inputs(107)) and not (inputs(233));
    layer0_outputs(4317) <= not((inputs(66)) xor (inputs(191)));
    layer0_outputs(4318) <= inputs(167);
    layer0_outputs(4319) <= not((inputs(139)) and (inputs(133)));
    layer0_outputs(4320) <= (inputs(56)) and (inputs(88));
    layer0_outputs(4321) <= (inputs(124)) and not (inputs(22));
    layer0_outputs(4322) <= not((inputs(166)) xor (inputs(184)));
    layer0_outputs(4323) <= not((inputs(168)) xor (inputs(74)));
    layer0_outputs(4324) <= (inputs(233)) and not (inputs(2));
    layer0_outputs(4325) <= inputs(166);
    layer0_outputs(4326) <= (inputs(167)) and not (inputs(68));
    layer0_outputs(4327) <= (inputs(193)) xor (inputs(196));
    layer0_outputs(4328) <= not(inputs(250));
    layer0_outputs(4329) <= (inputs(191)) and (inputs(238));
    layer0_outputs(4330) <= not((inputs(7)) xor (inputs(237)));
    layer0_outputs(4331) <= not((inputs(85)) and (inputs(165)));
    layer0_outputs(4332) <= not(inputs(116));
    layer0_outputs(4333) <= not(inputs(228)) or (inputs(83));
    layer0_outputs(4334) <= not(inputs(118));
    layer0_outputs(4335) <= not(inputs(237));
    layer0_outputs(4336) <= (inputs(141)) and not (inputs(31));
    layer0_outputs(4337) <= not((inputs(224)) xor (inputs(21)));
    layer0_outputs(4338) <= inputs(104);
    layer0_outputs(4339) <= (inputs(194)) or (inputs(222));
    layer0_outputs(4340) <= not((inputs(169)) or (inputs(6)));
    layer0_outputs(4341) <= (inputs(255)) xor (inputs(114));
    layer0_outputs(4342) <= (inputs(107)) xor (inputs(136));
    layer0_outputs(4343) <= not(inputs(40));
    layer0_outputs(4344) <= not((inputs(84)) or (inputs(29)));
    layer0_outputs(4345) <= (inputs(25)) and not (inputs(136));
    layer0_outputs(4346) <= (inputs(214)) or (inputs(96));
    layer0_outputs(4347) <= not(inputs(232));
    layer0_outputs(4348) <= not((inputs(222)) xor (inputs(193)));
    layer0_outputs(4349) <= inputs(5);
    layer0_outputs(4350) <= (inputs(190)) or (inputs(192));
    layer0_outputs(4351) <= (inputs(191)) or (inputs(251));
    layer0_outputs(4352) <= not(inputs(170)) or (inputs(72));
    layer0_outputs(4353) <= inputs(76);
    layer0_outputs(4354) <= not((inputs(122)) and (inputs(91)));
    layer0_outputs(4355) <= not((inputs(183)) xor (inputs(28)));
    layer0_outputs(4356) <= not(inputs(216)) or (inputs(220));
    layer0_outputs(4357) <= not(inputs(111)) or (inputs(1));
    layer0_outputs(4358) <= (inputs(255)) xor (inputs(173));
    layer0_outputs(4359) <= not((inputs(75)) or (inputs(77)));
    layer0_outputs(4360) <= not((inputs(92)) xor (inputs(255)));
    layer0_outputs(4361) <= (inputs(21)) and not (inputs(157));
    layer0_outputs(4362) <= not(inputs(60));
    layer0_outputs(4363) <= (inputs(198)) and not (inputs(183));
    layer0_outputs(4364) <= not((inputs(243)) and (inputs(201)));
    layer0_outputs(4365) <= not((inputs(220)) or (inputs(54)));
    layer0_outputs(4366) <= not((inputs(249)) or (inputs(142)));
    layer0_outputs(4367) <= not(inputs(118));
    layer0_outputs(4368) <= (inputs(100)) and not (inputs(192));
    layer0_outputs(4369) <= '0';
    layer0_outputs(4370) <= inputs(8);
    layer0_outputs(4371) <= (inputs(85)) and not (inputs(125));
    layer0_outputs(4372) <= (inputs(27)) or (inputs(51));
    layer0_outputs(4373) <= not(inputs(113));
    layer0_outputs(4374) <= (inputs(104)) xor (inputs(48));
    layer0_outputs(4375) <= not(inputs(90)) or (inputs(250));
    layer0_outputs(4376) <= not((inputs(45)) xor (inputs(87)));
    layer0_outputs(4377) <= not((inputs(0)) or (inputs(153)));
    layer0_outputs(4378) <= inputs(184);
    layer0_outputs(4379) <= inputs(74);
    layer0_outputs(4380) <= not(inputs(183)) or (inputs(191));
    layer0_outputs(4381) <= inputs(72);
    layer0_outputs(4382) <= not(inputs(59));
    layer0_outputs(4383) <= inputs(73);
    layer0_outputs(4384) <= not(inputs(118));
    layer0_outputs(4385) <= not(inputs(9));
    layer0_outputs(4386) <= not(inputs(104));
    layer0_outputs(4387) <= (inputs(175)) and not (inputs(54));
    layer0_outputs(4388) <= not((inputs(32)) xor (inputs(200)));
    layer0_outputs(4389) <= not((inputs(206)) or (inputs(98)));
    layer0_outputs(4390) <= (inputs(60)) xor (inputs(79));
    layer0_outputs(4391) <= not(inputs(98));
    layer0_outputs(4392) <= inputs(134);
    layer0_outputs(4393) <= not((inputs(172)) or (inputs(130)));
    layer0_outputs(4394) <= (inputs(79)) or (inputs(245));
    layer0_outputs(4395) <= inputs(16);
    layer0_outputs(4396) <= not(inputs(244));
    layer0_outputs(4397) <= not(inputs(176));
    layer0_outputs(4398) <= not((inputs(69)) xor (inputs(83)));
    layer0_outputs(4399) <= inputs(35);
    layer0_outputs(4400) <= (inputs(86)) or (inputs(141));
    layer0_outputs(4401) <= not((inputs(161)) and (inputs(227)));
    layer0_outputs(4402) <= (inputs(34)) xor (inputs(123));
    layer0_outputs(4403) <= inputs(109);
    layer0_outputs(4404) <= not(inputs(98)) or (inputs(94));
    layer0_outputs(4405) <= not((inputs(125)) xor (inputs(88)));
    layer0_outputs(4406) <= not((inputs(230)) xor (inputs(135)));
    layer0_outputs(4407) <= '1';
    layer0_outputs(4408) <= not(inputs(8));
    layer0_outputs(4409) <= not(inputs(99));
    layer0_outputs(4410) <= inputs(104);
    layer0_outputs(4411) <= (inputs(115)) or (inputs(171));
    layer0_outputs(4412) <= not(inputs(93));
    layer0_outputs(4413) <= (inputs(54)) and not (inputs(113));
    layer0_outputs(4414) <= (inputs(32)) xor (inputs(168));
    layer0_outputs(4415) <= not(inputs(178));
    layer0_outputs(4416) <= '0';
    layer0_outputs(4417) <= not((inputs(112)) or (inputs(124)));
    layer0_outputs(4418) <= (inputs(46)) and not (inputs(76));
    layer0_outputs(4419) <= not((inputs(133)) or (inputs(227)));
    layer0_outputs(4420) <= (inputs(237)) or (inputs(87));
    layer0_outputs(4421) <= (inputs(73)) or (inputs(57));
    layer0_outputs(4422) <= not((inputs(114)) or (inputs(145)));
    layer0_outputs(4423) <= (inputs(143)) xor (inputs(212));
    layer0_outputs(4424) <= not(inputs(146));
    layer0_outputs(4425) <= (inputs(137)) xor (inputs(234));
    layer0_outputs(4426) <= not((inputs(87)) xor (inputs(101)));
    layer0_outputs(4427) <= (inputs(238)) xor (inputs(17));
    layer0_outputs(4428) <= (inputs(180)) and not (inputs(128));
    layer0_outputs(4429) <= not((inputs(6)) xor (inputs(52)));
    layer0_outputs(4430) <= inputs(167);
    layer0_outputs(4431) <= (inputs(136)) and not (inputs(61));
    layer0_outputs(4432) <= not((inputs(220)) or (inputs(255)));
    layer0_outputs(4433) <= (inputs(205)) xor (inputs(23));
    layer0_outputs(4434) <= '0';
    layer0_outputs(4435) <= inputs(187);
    layer0_outputs(4436) <= '1';
    layer0_outputs(4437) <= (inputs(111)) or (inputs(220));
    layer0_outputs(4438) <= not((inputs(104)) xor (inputs(59)));
    layer0_outputs(4439) <= (inputs(35)) xor (inputs(11));
    layer0_outputs(4440) <= not(inputs(241));
    layer0_outputs(4441) <= (inputs(101)) or (inputs(145));
    layer0_outputs(4442) <= not((inputs(131)) and (inputs(159)));
    layer0_outputs(4443) <= (inputs(61)) and not (inputs(100));
    layer0_outputs(4444) <= not(inputs(129)) or (inputs(252));
    layer0_outputs(4445) <= not((inputs(45)) xor (inputs(195)));
    layer0_outputs(4446) <= (inputs(187)) xor (inputs(5));
    layer0_outputs(4447) <= not(inputs(70)) or (inputs(194));
    layer0_outputs(4448) <= not(inputs(196)) or (inputs(39));
    layer0_outputs(4449) <= (inputs(49)) xor (inputs(242));
    layer0_outputs(4450) <= (inputs(43)) and not (inputs(221));
    layer0_outputs(4451) <= (inputs(112)) or (inputs(234));
    layer0_outputs(4452) <= inputs(83);
    layer0_outputs(4453) <= (inputs(99)) and not (inputs(79));
    layer0_outputs(4454) <= not(inputs(212));
    layer0_outputs(4455) <= not((inputs(131)) xor (inputs(199)));
    layer0_outputs(4456) <= not(inputs(108));
    layer0_outputs(4457) <= not((inputs(218)) or (inputs(205)));
    layer0_outputs(4458) <= inputs(134);
    layer0_outputs(4459) <= not((inputs(240)) xor (inputs(63)));
    layer0_outputs(4460) <= not((inputs(192)) or (inputs(166)));
    layer0_outputs(4461) <= (inputs(83)) and not (inputs(2));
    layer0_outputs(4462) <= not(inputs(7));
    layer0_outputs(4463) <= inputs(24);
    layer0_outputs(4464) <= (inputs(42)) and not (inputs(211));
    layer0_outputs(4465) <= not(inputs(120)) or (inputs(175));
    layer0_outputs(4466) <= not((inputs(53)) or (inputs(101)));
    layer0_outputs(4467) <= not(inputs(28));
    layer0_outputs(4468) <= inputs(151);
    layer0_outputs(4469) <= (inputs(159)) xor (inputs(224));
    layer0_outputs(4470) <= (inputs(229)) or (inputs(245));
    layer0_outputs(4471) <= not(inputs(194)) or (inputs(253));
    layer0_outputs(4472) <= not(inputs(101));
    layer0_outputs(4473) <= not(inputs(150));
    layer0_outputs(4474) <= (inputs(102)) xor (inputs(38));
    layer0_outputs(4475) <= (inputs(224)) or (inputs(16));
    layer0_outputs(4476) <= inputs(76);
    layer0_outputs(4477) <= (inputs(165)) xor (inputs(240));
    layer0_outputs(4478) <= not(inputs(71));
    layer0_outputs(4479) <= inputs(93);
    layer0_outputs(4480) <= inputs(230);
    layer0_outputs(4481) <= (inputs(194)) or (inputs(171));
    layer0_outputs(4482) <= inputs(85);
    layer0_outputs(4483) <= not(inputs(107));
    layer0_outputs(4484) <= not(inputs(162));
    layer0_outputs(4485) <= inputs(23);
    layer0_outputs(4486) <= not(inputs(121)) or (inputs(57));
    layer0_outputs(4487) <= (inputs(246)) or (inputs(141));
    layer0_outputs(4488) <= not((inputs(41)) or (inputs(57)));
    layer0_outputs(4489) <= not((inputs(82)) xor (inputs(68)));
    layer0_outputs(4490) <= inputs(38);
    layer0_outputs(4491) <= not(inputs(125)) or (inputs(134));
    layer0_outputs(4492) <= inputs(125);
    layer0_outputs(4493) <= (inputs(149)) xor (inputs(148));
    layer0_outputs(4494) <= not((inputs(15)) xor (inputs(69)));
    layer0_outputs(4495) <= (inputs(173)) and (inputs(122));
    layer0_outputs(4496) <= (inputs(56)) and (inputs(119));
    layer0_outputs(4497) <= not(inputs(129));
    layer0_outputs(4498) <= not((inputs(30)) xor (inputs(218)));
    layer0_outputs(4499) <= not(inputs(91)) or (inputs(223));
    layer0_outputs(4500) <= not(inputs(156));
    layer0_outputs(4501) <= not(inputs(60)) or (inputs(104));
    layer0_outputs(4502) <= not((inputs(45)) xor (inputs(18)));
    layer0_outputs(4503) <= not(inputs(105));
    layer0_outputs(4504) <= not((inputs(51)) xor (inputs(239)));
    layer0_outputs(4505) <= inputs(130);
    layer0_outputs(4506) <= not(inputs(9));
    layer0_outputs(4507) <= not((inputs(233)) or (inputs(213)));
    layer0_outputs(4508) <= not(inputs(4)) or (inputs(15));
    layer0_outputs(4509) <= not(inputs(118));
    layer0_outputs(4510) <= inputs(214);
    layer0_outputs(4511) <= not(inputs(232));
    layer0_outputs(4512) <= (inputs(141)) or (inputs(1));
    layer0_outputs(4513) <= (inputs(83)) or (inputs(163));
    layer0_outputs(4514) <= (inputs(115)) and not (inputs(17));
    layer0_outputs(4515) <= (inputs(165)) xor (inputs(23));
    layer0_outputs(4516) <= not(inputs(105)) or (inputs(130));
    layer0_outputs(4517) <= (inputs(216)) and not (inputs(8));
    layer0_outputs(4518) <= not(inputs(217));
    layer0_outputs(4519) <= (inputs(214)) or (inputs(19));
    layer0_outputs(4520) <= (inputs(227)) or (inputs(246));
    layer0_outputs(4521) <= (inputs(89)) and not (inputs(70));
    layer0_outputs(4522) <= (inputs(127)) and not (inputs(88));
    layer0_outputs(4523) <= (inputs(89)) xor (inputs(107));
    layer0_outputs(4524) <= not(inputs(66));
    layer0_outputs(4525) <= not(inputs(163));
    layer0_outputs(4526) <= not(inputs(109)) or (inputs(82));
    layer0_outputs(4527) <= not(inputs(100));
    layer0_outputs(4528) <= not(inputs(200)) or (inputs(63));
    layer0_outputs(4529) <= not(inputs(74));
    layer0_outputs(4530) <= not(inputs(107));
    layer0_outputs(4531) <= not(inputs(3));
    layer0_outputs(4532) <= (inputs(96)) or (inputs(183));
    layer0_outputs(4533) <= not(inputs(182));
    layer0_outputs(4534) <= (inputs(127)) and not (inputs(249));
    layer0_outputs(4535) <= not((inputs(52)) or (inputs(128)));
    layer0_outputs(4536) <= (inputs(52)) or (inputs(94));
    layer0_outputs(4537) <= not(inputs(26)) or (inputs(244));
    layer0_outputs(4538) <= (inputs(180)) or (inputs(32));
    layer0_outputs(4539) <= not((inputs(205)) or (inputs(192)));
    layer0_outputs(4540) <= (inputs(180)) or (inputs(152));
    layer0_outputs(4541) <= (inputs(22)) xor (inputs(147));
    layer0_outputs(4542) <= not((inputs(109)) or (inputs(95)));
    layer0_outputs(4543) <= (inputs(249)) xor (inputs(202));
    layer0_outputs(4544) <= not(inputs(75));
    layer0_outputs(4545) <= (inputs(32)) or (inputs(197));
    layer0_outputs(4546) <= inputs(70);
    layer0_outputs(4547) <= (inputs(254)) and (inputs(234));
    layer0_outputs(4548) <= inputs(224);
    layer0_outputs(4549) <= not(inputs(225)) or (inputs(11));
    layer0_outputs(4550) <= inputs(30);
    layer0_outputs(4551) <= (inputs(247)) and not (inputs(47));
    layer0_outputs(4552) <= inputs(10);
    layer0_outputs(4553) <= not((inputs(18)) xor (inputs(94)));
    layer0_outputs(4554) <= not(inputs(121));
    layer0_outputs(4555) <= inputs(150);
    layer0_outputs(4556) <= not((inputs(76)) xor (inputs(195)));
    layer0_outputs(4557) <= not((inputs(7)) and (inputs(223)));
    layer0_outputs(4558) <= '1';
    layer0_outputs(4559) <= not((inputs(122)) or (inputs(106)));
    layer0_outputs(4560) <= not((inputs(66)) and (inputs(143)));
    layer0_outputs(4561) <= not(inputs(29));
    layer0_outputs(4562) <= not(inputs(109));
    layer0_outputs(4563) <= not((inputs(52)) and (inputs(45)));
    layer0_outputs(4564) <= (inputs(193)) xor (inputs(22));
    layer0_outputs(4565) <= (inputs(54)) and not (inputs(34));
    layer0_outputs(4566) <= (inputs(123)) xor (inputs(157));
    layer0_outputs(4567) <= inputs(248);
    layer0_outputs(4568) <= (inputs(95)) or (inputs(55));
    layer0_outputs(4569) <= not(inputs(97));
    layer0_outputs(4570) <= not(inputs(170)) or (inputs(84));
    layer0_outputs(4571) <= (inputs(181)) or (inputs(212));
    layer0_outputs(4572) <= inputs(192);
    layer0_outputs(4573) <= not(inputs(129));
    layer0_outputs(4574) <= inputs(29);
    layer0_outputs(4575) <= not((inputs(107)) or (inputs(6)));
    layer0_outputs(4576) <= not(inputs(102));
    layer0_outputs(4577) <= inputs(136);
    layer0_outputs(4578) <= not(inputs(108)) or (inputs(31));
    layer0_outputs(4579) <= not(inputs(106));
    layer0_outputs(4580) <= (inputs(105)) and not (inputs(2));
    layer0_outputs(4581) <= (inputs(123)) or (inputs(94));
    layer0_outputs(4582) <= inputs(98);
    layer0_outputs(4583) <= (inputs(28)) or (inputs(0));
    layer0_outputs(4584) <= (inputs(9)) or (inputs(181));
    layer0_outputs(4585) <= not((inputs(58)) xor (inputs(72)));
    layer0_outputs(4586) <= inputs(100);
    layer0_outputs(4587) <= (inputs(218)) xor (inputs(171));
    layer0_outputs(4588) <= inputs(237);
    layer0_outputs(4589) <= not((inputs(102)) xor (inputs(37)));
    layer0_outputs(4590) <= inputs(146);
    layer0_outputs(4591) <= not((inputs(7)) xor (inputs(17)));
    layer0_outputs(4592) <= (inputs(33)) or (inputs(43));
    layer0_outputs(4593) <= (inputs(202)) and not (inputs(143));
    layer0_outputs(4594) <= not((inputs(129)) or (inputs(114)));
    layer0_outputs(4595) <= inputs(232);
    layer0_outputs(4596) <= not((inputs(162)) or (inputs(183)));
    layer0_outputs(4597) <= (inputs(160)) or (inputs(165));
    layer0_outputs(4598) <= not(inputs(213)) or (inputs(166));
    layer0_outputs(4599) <= not(inputs(113));
    layer0_outputs(4600) <= not(inputs(151));
    layer0_outputs(4601) <= (inputs(113)) or (inputs(37));
    layer0_outputs(4602) <= (inputs(47)) or (inputs(226));
    layer0_outputs(4603) <= (inputs(40)) and not (inputs(73));
    layer0_outputs(4604) <= not(inputs(130));
    layer0_outputs(4605) <= inputs(41);
    layer0_outputs(4606) <= inputs(162);
    layer0_outputs(4607) <= not((inputs(212)) or (inputs(144)));
    layer0_outputs(4608) <= inputs(94);
    layer0_outputs(4609) <= (inputs(21)) and not (inputs(84));
    layer0_outputs(4610) <= not((inputs(68)) xor (inputs(160)));
    layer0_outputs(4611) <= not(inputs(110)) or (inputs(251));
    layer0_outputs(4612) <= not(inputs(40)) or (inputs(242));
    layer0_outputs(4613) <= inputs(109);
    layer0_outputs(4614) <= not(inputs(140)) or (inputs(177));
    layer0_outputs(4615) <= not((inputs(157)) or (inputs(85)));
    layer0_outputs(4616) <= (inputs(136)) and not (inputs(115));
    layer0_outputs(4617) <= not(inputs(27));
    layer0_outputs(4618) <= inputs(212);
    layer0_outputs(4619) <= '0';
    layer0_outputs(4620) <= inputs(181);
    layer0_outputs(4621) <= (inputs(91)) and not (inputs(240));
    layer0_outputs(4622) <= (inputs(61)) and (inputs(122));
    layer0_outputs(4623) <= (inputs(155)) and not (inputs(206));
    layer0_outputs(4624) <= (inputs(219)) or (inputs(203));
    layer0_outputs(4625) <= not(inputs(92));
    layer0_outputs(4626) <= not(inputs(220));
    layer0_outputs(4627) <= not(inputs(79));
    layer0_outputs(4628) <= (inputs(237)) xor (inputs(106));
    layer0_outputs(4629) <= not((inputs(79)) or (inputs(117)));
    layer0_outputs(4630) <= not((inputs(215)) or (inputs(231)));
    layer0_outputs(4631) <= not((inputs(69)) or (inputs(63)));
    layer0_outputs(4632) <= not(inputs(116)) or (inputs(126));
    layer0_outputs(4633) <= inputs(246);
    layer0_outputs(4634) <= inputs(145);
    layer0_outputs(4635) <= not((inputs(39)) and (inputs(40)));
    layer0_outputs(4636) <= (inputs(150)) and not (inputs(31));
    layer0_outputs(4637) <= inputs(246);
    layer0_outputs(4638) <= not(inputs(227));
    layer0_outputs(4639) <= not(inputs(92));
    layer0_outputs(4640) <= inputs(246);
    layer0_outputs(4641) <= not((inputs(96)) or (inputs(114)));
    layer0_outputs(4642) <= not(inputs(229)) or (inputs(166));
    layer0_outputs(4643) <= (inputs(69)) and not (inputs(225));
    layer0_outputs(4644) <= not((inputs(199)) or (inputs(153)));
    layer0_outputs(4645) <= inputs(109);
    layer0_outputs(4646) <= (inputs(129)) and (inputs(17));
    layer0_outputs(4647) <= not(inputs(19)) or (inputs(80));
    layer0_outputs(4648) <= not((inputs(143)) xor (inputs(172)));
    layer0_outputs(4649) <= not((inputs(228)) or (inputs(227)));
    layer0_outputs(4650) <= (inputs(153)) and not (inputs(18));
    layer0_outputs(4651) <= (inputs(123)) and (inputs(91));
    layer0_outputs(4652) <= not((inputs(43)) xor (inputs(65)));
    layer0_outputs(4653) <= (inputs(35)) or (inputs(255));
    layer0_outputs(4654) <= (inputs(167)) or (inputs(140));
    layer0_outputs(4655) <= not(inputs(201)) or (inputs(35));
    layer0_outputs(4656) <= not((inputs(178)) or (inputs(127)));
    layer0_outputs(4657) <= inputs(103);
    layer0_outputs(4658) <= not(inputs(117));
    layer0_outputs(4659) <= not((inputs(43)) and (inputs(159)));
    layer0_outputs(4660) <= (inputs(79)) or (inputs(219));
    layer0_outputs(4661) <= not(inputs(99));
    layer0_outputs(4662) <= not((inputs(245)) xor (inputs(103)));
    layer0_outputs(4663) <= not(inputs(85)) or (inputs(250));
    layer0_outputs(4664) <= (inputs(160)) xor (inputs(59));
    layer0_outputs(4665) <= not((inputs(146)) or (inputs(251)));
    layer0_outputs(4666) <= (inputs(146)) and not (inputs(66));
    layer0_outputs(4667) <= (inputs(255)) and not (inputs(96));
    layer0_outputs(4668) <= not(inputs(137)) or (inputs(122));
    layer0_outputs(4669) <= not((inputs(38)) and (inputs(104)));
    layer0_outputs(4670) <= not((inputs(120)) xor (inputs(76)));
    layer0_outputs(4671) <= (inputs(126)) or (inputs(59));
    layer0_outputs(4672) <= (inputs(96)) and not (inputs(250));
    layer0_outputs(4673) <= inputs(90);
    layer0_outputs(4674) <= (inputs(97)) or (inputs(246));
    layer0_outputs(4675) <= not(inputs(164));
    layer0_outputs(4676) <= inputs(67);
    layer0_outputs(4677) <= (inputs(41)) and not (inputs(253));
    layer0_outputs(4678) <= inputs(166);
    layer0_outputs(4679) <= (inputs(137)) xor (inputs(213));
    layer0_outputs(4680) <= not(inputs(195)) or (inputs(120));
    layer0_outputs(4681) <= not(inputs(179)) or (inputs(109));
    layer0_outputs(4682) <= not((inputs(202)) xor (inputs(182)));
    layer0_outputs(4683) <= not(inputs(135));
    layer0_outputs(4684) <= not(inputs(199)) or (inputs(62));
    layer0_outputs(4685) <= (inputs(36)) and (inputs(246));
    layer0_outputs(4686) <= (inputs(178)) or (inputs(185));
    layer0_outputs(4687) <= not(inputs(22));
    layer0_outputs(4688) <= not(inputs(23)) or (inputs(50));
    layer0_outputs(4689) <= (inputs(51)) or (inputs(208));
    layer0_outputs(4690) <= inputs(255);
    layer0_outputs(4691) <= inputs(114);
    layer0_outputs(4692) <= not(inputs(243)) or (inputs(71));
    layer0_outputs(4693) <= (inputs(93)) xor (inputs(234));
    layer0_outputs(4694) <= (inputs(198)) and not (inputs(87));
    layer0_outputs(4695) <= (inputs(130)) or (inputs(78));
    layer0_outputs(4696) <= (inputs(198)) and not (inputs(53));
    layer0_outputs(4697) <= not((inputs(46)) or (inputs(54)));
    layer0_outputs(4698) <= inputs(75);
    layer0_outputs(4699) <= not(inputs(169));
    layer0_outputs(4700) <= not((inputs(234)) or (inputs(25)));
    layer0_outputs(4701) <= (inputs(191)) or (inputs(233));
    layer0_outputs(4702) <= (inputs(181)) or (inputs(96));
    layer0_outputs(4703) <= not(inputs(26));
    layer0_outputs(4704) <= (inputs(114)) and not (inputs(75));
    layer0_outputs(4705) <= not(inputs(136)) or (inputs(238));
    layer0_outputs(4706) <= not(inputs(178)) or (inputs(202));
    layer0_outputs(4707) <= not(inputs(50));
    layer0_outputs(4708) <= not((inputs(163)) or (inputs(220)));
    layer0_outputs(4709) <= (inputs(8)) and (inputs(105));
    layer0_outputs(4710) <= inputs(249);
    layer0_outputs(4711) <= inputs(9);
    layer0_outputs(4712) <= (inputs(126)) xor (inputs(140));
    layer0_outputs(4713) <= not(inputs(177)) or (inputs(249));
    layer0_outputs(4714) <= (inputs(161)) and not (inputs(128));
    layer0_outputs(4715) <= inputs(109);
    layer0_outputs(4716) <= not(inputs(58)) or (inputs(206));
    layer0_outputs(4717) <= (inputs(114)) xor (inputs(117));
    layer0_outputs(4718) <= not(inputs(183)) or (inputs(57));
    layer0_outputs(4719) <= not(inputs(245));
    layer0_outputs(4720) <= inputs(116);
    layer0_outputs(4721) <= (inputs(154)) and (inputs(7));
    layer0_outputs(4722) <= not((inputs(3)) and (inputs(1)));
    layer0_outputs(4723) <= (inputs(37)) or (inputs(18));
    layer0_outputs(4724) <= not((inputs(133)) or (inputs(177)));
    layer0_outputs(4725) <= (inputs(107)) or (inputs(247));
    layer0_outputs(4726) <= not(inputs(85));
    layer0_outputs(4727) <= (inputs(119)) and not (inputs(0));
    layer0_outputs(4728) <= not((inputs(27)) xor (inputs(238)));
    layer0_outputs(4729) <= (inputs(137)) and not (inputs(11));
    layer0_outputs(4730) <= not(inputs(220));
    layer0_outputs(4731) <= not((inputs(96)) and (inputs(58)));
    layer0_outputs(4732) <= not(inputs(151));
    layer0_outputs(4733) <= not(inputs(214)) or (inputs(239));
    layer0_outputs(4734) <= '0';
    layer0_outputs(4735) <= inputs(94);
    layer0_outputs(4736) <= not(inputs(230));
    layer0_outputs(4737) <= not((inputs(204)) xor (inputs(89)));
    layer0_outputs(4738) <= (inputs(190)) and not (inputs(48));
    layer0_outputs(4739) <= not(inputs(25));
    layer0_outputs(4740) <= (inputs(3)) and not (inputs(190));
    layer0_outputs(4741) <= not(inputs(56));
    layer0_outputs(4742) <= (inputs(124)) and not (inputs(236));
    layer0_outputs(4743) <= (inputs(139)) xor (inputs(158));
    layer0_outputs(4744) <= '0';
    layer0_outputs(4745) <= not((inputs(227)) or (inputs(250)));
    layer0_outputs(4746) <= (inputs(146)) or (inputs(145));
    layer0_outputs(4747) <= not(inputs(65)) or (inputs(73));
    layer0_outputs(4748) <= inputs(62);
    layer0_outputs(4749) <= (inputs(236)) xor (inputs(220));
    layer0_outputs(4750) <= inputs(147);
    layer0_outputs(4751) <= (inputs(191)) or (inputs(212));
    layer0_outputs(4752) <= not(inputs(182)) or (inputs(54));
    layer0_outputs(4753) <= (inputs(31)) or (inputs(30));
    layer0_outputs(4754) <= not((inputs(142)) and (inputs(113)));
    layer0_outputs(4755) <= (inputs(101)) and not (inputs(61));
    layer0_outputs(4756) <= (inputs(85)) and not (inputs(124));
    layer0_outputs(4757) <= (inputs(152)) xor (inputs(232));
    layer0_outputs(4758) <= not(inputs(231)) or (inputs(205));
    layer0_outputs(4759) <= (inputs(248)) or (inputs(34));
    layer0_outputs(4760) <= inputs(102);
    layer0_outputs(4761) <= inputs(201);
    layer0_outputs(4762) <= not((inputs(223)) or (inputs(249)));
    layer0_outputs(4763) <= inputs(88);
    layer0_outputs(4764) <= (inputs(196)) and not (inputs(255));
    layer0_outputs(4765) <= inputs(188);
    layer0_outputs(4766) <= (inputs(215)) xor (inputs(122));
    layer0_outputs(4767) <= not(inputs(245)) or (inputs(151));
    layer0_outputs(4768) <= inputs(236);
    layer0_outputs(4769) <= not((inputs(158)) and (inputs(37)));
    layer0_outputs(4770) <= not(inputs(122)) or (inputs(175));
    layer0_outputs(4771) <= not(inputs(32)) or (inputs(222));
    layer0_outputs(4772) <= inputs(210);
    layer0_outputs(4773) <= not((inputs(203)) xor (inputs(169)));
    layer0_outputs(4774) <= (inputs(102)) xor (inputs(131));
    layer0_outputs(4775) <= not((inputs(75)) and (inputs(59)));
    layer0_outputs(4776) <= not((inputs(251)) and (inputs(46)));
    layer0_outputs(4777) <= not(inputs(205));
    layer0_outputs(4778) <= not(inputs(231)) or (inputs(33));
    layer0_outputs(4779) <= not((inputs(57)) and (inputs(6)));
    layer0_outputs(4780) <= (inputs(157)) xor (inputs(5));
    layer0_outputs(4781) <= (inputs(170)) xor (inputs(181));
    layer0_outputs(4782) <= not((inputs(48)) or (inputs(89)));
    layer0_outputs(4783) <= not((inputs(164)) xor (inputs(157)));
    layer0_outputs(4784) <= inputs(218);
    layer0_outputs(4785) <= not(inputs(229));
    layer0_outputs(4786) <= inputs(234);
    layer0_outputs(4787) <= (inputs(98)) or (inputs(156));
    layer0_outputs(4788) <= not(inputs(117));
    layer0_outputs(4789) <= not((inputs(2)) or (inputs(4)));
    layer0_outputs(4790) <= not(inputs(35));
    layer0_outputs(4791) <= (inputs(109)) and not (inputs(223));
    layer0_outputs(4792) <= (inputs(192)) or (inputs(134));
    layer0_outputs(4793) <= not((inputs(177)) or (inputs(100)));
    layer0_outputs(4794) <= (inputs(236)) and not (inputs(94));
    layer0_outputs(4795) <= not((inputs(4)) or (inputs(68)));
    layer0_outputs(4796) <= not((inputs(212)) or (inputs(128)));
    layer0_outputs(4797) <= '1';
    layer0_outputs(4798) <= inputs(63);
    layer0_outputs(4799) <= (inputs(191)) xor (inputs(99));
    layer0_outputs(4800) <= not(inputs(217));
    layer0_outputs(4801) <= inputs(133);
    layer0_outputs(4802) <= not((inputs(64)) xor (inputs(55)));
    layer0_outputs(4803) <= not(inputs(197)) or (inputs(238));
    layer0_outputs(4804) <= inputs(134);
    layer0_outputs(4805) <= (inputs(118)) and (inputs(138));
    layer0_outputs(4806) <= '1';
    layer0_outputs(4807) <= (inputs(227)) or (inputs(97));
    layer0_outputs(4808) <= not((inputs(143)) or (inputs(69)));
    layer0_outputs(4809) <= not((inputs(39)) or (inputs(194)));
    layer0_outputs(4810) <= not((inputs(128)) and (inputs(79)));
    layer0_outputs(4811) <= not((inputs(2)) xor (inputs(132)));
    layer0_outputs(4812) <= not(inputs(54)) or (inputs(12));
    layer0_outputs(4813) <= not(inputs(121)) or (inputs(197));
    layer0_outputs(4814) <= (inputs(174)) and not (inputs(30));
    layer0_outputs(4815) <= not(inputs(211)) or (inputs(57));
    layer0_outputs(4816) <= not(inputs(47)) or (inputs(160));
    layer0_outputs(4817) <= (inputs(123)) xor (inputs(90));
    layer0_outputs(4818) <= (inputs(17)) or (inputs(32));
    layer0_outputs(4819) <= (inputs(25)) or (inputs(110));
    layer0_outputs(4820) <= not((inputs(13)) or (inputs(16)));
    layer0_outputs(4821) <= inputs(59);
    layer0_outputs(4822) <= inputs(109);
    layer0_outputs(4823) <= not(inputs(53));
    layer0_outputs(4824) <= not((inputs(225)) or (inputs(37)));
    layer0_outputs(4825) <= inputs(177);
    layer0_outputs(4826) <= not(inputs(31)) or (inputs(198));
    layer0_outputs(4827) <= not(inputs(202));
    layer0_outputs(4828) <= not(inputs(162));
    layer0_outputs(4829) <= (inputs(56)) and not (inputs(208));
    layer0_outputs(4830) <= not(inputs(196));
    layer0_outputs(4831) <= (inputs(73)) or (inputs(18));
    layer0_outputs(4832) <= '0';
    layer0_outputs(4833) <= not(inputs(150)) or (inputs(183));
    layer0_outputs(4834) <= not(inputs(204));
    layer0_outputs(4835) <= (inputs(122)) or (inputs(150));
    layer0_outputs(4836) <= (inputs(15)) and not (inputs(157));
    layer0_outputs(4837) <= inputs(104);
    layer0_outputs(4838) <= not((inputs(111)) or (inputs(104)));
    layer0_outputs(4839) <= (inputs(85)) xor (inputs(129));
    layer0_outputs(4840) <= inputs(156);
    layer0_outputs(4841) <= not((inputs(79)) or (inputs(20)));
    layer0_outputs(4842) <= (inputs(137)) xor (inputs(164));
    layer0_outputs(4843) <= (inputs(181)) or (inputs(37));
    layer0_outputs(4844) <= (inputs(165)) xor (inputs(29));
    layer0_outputs(4845) <= not(inputs(129));
    layer0_outputs(4846) <= '1';
    layer0_outputs(4847) <= inputs(123);
    layer0_outputs(4848) <= inputs(91);
    layer0_outputs(4849) <= (inputs(71)) or (inputs(139));
    layer0_outputs(4850) <= (inputs(15)) xor (inputs(164));
    layer0_outputs(4851) <= not(inputs(109)) or (inputs(222));
    layer0_outputs(4852) <= not((inputs(181)) or (inputs(45)));
    layer0_outputs(4853) <= inputs(114);
    layer0_outputs(4854) <= not((inputs(184)) or (inputs(143)));
    layer0_outputs(4855) <= (inputs(2)) xor (inputs(190));
    layer0_outputs(4856) <= not((inputs(135)) xor (inputs(143)));
    layer0_outputs(4857) <= not((inputs(201)) or (inputs(176)));
    layer0_outputs(4858) <= (inputs(239)) xor (inputs(84));
    layer0_outputs(4859) <= not(inputs(172));
    layer0_outputs(4860) <= not(inputs(38));
    layer0_outputs(4861) <= (inputs(204)) and not (inputs(110));
    layer0_outputs(4862) <= not(inputs(201)) or (inputs(128));
    layer0_outputs(4863) <= (inputs(57)) and not (inputs(68));
    layer0_outputs(4864) <= (inputs(200)) and not (inputs(10));
    layer0_outputs(4865) <= (inputs(106)) and not (inputs(54));
    layer0_outputs(4866) <= (inputs(113)) and (inputs(178));
    layer0_outputs(4867) <= not(inputs(119));
    layer0_outputs(4868) <= not((inputs(86)) or (inputs(220)));
    layer0_outputs(4869) <= not(inputs(184));
    layer0_outputs(4870) <= inputs(67);
    layer0_outputs(4871) <= not((inputs(222)) or (inputs(165)));
    layer0_outputs(4872) <= not(inputs(209));
    layer0_outputs(4873) <= (inputs(33)) and not (inputs(97));
    layer0_outputs(4874) <= inputs(179);
    layer0_outputs(4875) <= (inputs(218)) and not (inputs(110));
    layer0_outputs(4876) <= (inputs(207)) or (inputs(249));
    layer0_outputs(4877) <= not(inputs(210));
    layer0_outputs(4878) <= (inputs(43)) or (inputs(21));
    layer0_outputs(4879) <= inputs(76);
    layer0_outputs(4880) <= '0';
    layer0_outputs(4881) <= inputs(108);
    layer0_outputs(4882) <= not(inputs(230));
    layer0_outputs(4883) <= not((inputs(232)) xor (inputs(223)));
    layer0_outputs(4884) <= (inputs(34)) and not (inputs(127));
    layer0_outputs(4885) <= not((inputs(38)) xor (inputs(44)));
    layer0_outputs(4886) <= not(inputs(225));
    layer0_outputs(4887) <= (inputs(132)) and not (inputs(205));
    layer0_outputs(4888) <= inputs(120);
    layer0_outputs(4889) <= not(inputs(105));
    layer0_outputs(4890) <= not((inputs(69)) or (inputs(128)));
    layer0_outputs(4891) <= (inputs(74)) or (inputs(66));
    layer0_outputs(4892) <= not(inputs(192)) or (inputs(65));
    layer0_outputs(4893) <= not(inputs(19));
    layer0_outputs(4894) <= not(inputs(26)) or (inputs(50));
    layer0_outputs(4895) <= not(inputs(217)) or (inputs(126));
    layer0_outputs(4896) <= (inputs(38)) xor (inputs(229));
    layer0_outputs(4897) <= (inputs(155)) xor (inputs(141));
    layer0_outputs(4898) <= not((inputs(194)) xor (inputs(9)));
    layer0_outputs(4899) <= (inputs(173)) or (inputs(83));
    layer0_outputs(4900) <= (inputs(16)) or (inputs(185));
    layer0_outputs(4901) <= not(inputs(122)) or (inputs(246));
    layer0_outputs(4902) <= not(inputs(140));
    layer0_outputs(4903) <= not(inputs(220)) or (inputs(114));
    layer0_outputs(4904) <= not((inputs(129)) or (inputs(145)));
    layer0_outputs(4905) <= (inputs(43)) and not (inputs(171));
    layer0_outputs(4906) <= not(inputs(182));
    layer0_outputs(4907) <= (inputs(220)) xor (inputs(237));
    layer0_outputs(4908) <= (inputs(248)) and not (inputs(255));
    layer0_outputs(4909) <= not(inputs(253));
    layer0_outputs(4910) <= not(inputs(185));
    layer0_outputs(4911) <= not(inputs(162)) or (inputs(104));
    layer0_outputs(4912) <= (inputs(6)) xor (inputs(239));
    layer0_outputs(4913) <= (inputs(215)) and not (inputs(140));
    layer0_outputs(4914) <= not(inputs(130));
    layer0_outputs(4915) <= (inputs(217)) xor (inputs(205));
    layer0_outputs(4916) <= inputs(162);
    layer0_outputs(4917) <= not((inputs(1)) or (inputs(55)));
    layer0_outputs(4918) <= inputs(199);
    layer0_outputs(4919) <= (inputs(154)) or (inputs(144));
    layer0_outputs(4920) <= not(inputs(81));
    layer0_outputs(4921) <= not((inputs(249)) xor (inputs(202)));
    layer0_outputs(4922) <= (inputs(134)) or (inputs(80));
    layer0_outputs(4923) <= not((inputs(77)) or (inputs(43)));
    layer0_outputs(4924) <= (inputs(116)) and not (inputs(111));
    layer0_outputs(4925) <= not(inputs(175));
    layer0_outputs(4926) <= not(inputs(215));
    layer0_outputs(4927) <= not(inputs(156)) or (inputs(70));
    layer0_outputs(4928) <= not(inputs(58));
    layer0_outputs(4929) <= not(inputs(100));
    layer0_outputs(4930) <= not(inputs(125));
    layer0_outputs(4931) <= not((inputs(184)) xor (inputs(174)));
    layer0_outputs(4932) <= '0';
    layer0_outputs(4933) <= inputs(150);
    layer0_outputs(4934) <= (inputs(130)) and not (inputs(80));
    layer0_outputs(4935) <= (inputs(221)) and (inputs(42));
    layer0_outputs(4936) <= not(inputs(204)) or (inputs(103));
    layer0_outputs(4937) <= not((inputs(223)) and (inputs(144)));
    layer0_outputs(4938) <= (inputs(121)) and not (inputs(145));
    layer0_outputs(4939) <= not((inputs(195)) or (inputs(175)));
    layer0_outputs(4940) <= (inputs(241)) or (inputs(120));
    layer0_outputs(4941) <= (inputs(86)) xor (inputs(44));
    layer0_outputs(4942) <= (inputs(121)) and not (inputs(191));
    layer0_outputs(4943) <= inputs(209);
    layer0_outputs(4944) <= (inputs(183)) or (inputs(66));
    layer0_outputs(4945) <= inputs(45);
    layer0_outputs(4946) <= (inputs(166)) and not (inputs(3));
    layer0_outputs(4947) <= not((inputs(50)) and (inputs(132)));
    layer0_outputs(4948) <= (inputs(202)) and (inputs(244));
    layer0_outputs(4949) <= not(inputs(129));
    layer0_outputs(4950) <= (inputs(79)) and not (inputs(6));
    layer0_outputs(4951) <= (inputs(169)) and not (inputs(221));
    layer0_outputs(4952) <= not(inputs(91));
    layer0_outputs(4953) <= inputs(25);
    layer0_outputs(4954) <= (inputs(11)) xor (inputs(72));
    layer0_outputs(4955) <= (inputs(244)) and not (inputs(206));
    layer0_outputs(4956) <= not((inputs(180)) or (inputs(38)));
    layer0_outputs(4957) <= not((inputs(38)) or (inputs(158)));
    layer0_outputs(4958) <= not(inputs(249)) or (inputs(62));
    layer0_outputs(4959) <= not(inputs(120)) or (inputs(171));
    layer0_outputs(4960) <= inputs(24);
    layer0_outputs(4961) <= not((inputs(214)) or (inputs(160)));
    layer0_outputs(4962) <= not((inputs(158)) or (inputs(77)));
    layer0_outputs(4963) <= (inputs(104)) and not (inputs(66));
    layer0_outputs(4964) <= (inputs(208)) xor (inputs(179));
    layer0_outputs(4965) <= not(inputs(208));
    layer0_outputs(4966) <= (inputs(90)) or (inputs(51));
    layer0_outputs(4967) <= (inputs(177)) or (inputs(192));
    layer0_outputs(4968) <= not(inputs(230)) or (inputs(75));
    layer0_outputs(4969) <= not((inputs(27)) or (inputs(52)));
    layer0_outputs(4970) <= not(inputs(91));
    layer0_outputs(4971) <= not(inputs(35));
    layer0_outputs(4972) <= not(inputs(75)) or (inputs(18));
    layer0_outputs(4973) <= inputs(20);
    layer0_outputs(4974) <= (inputs(132)) or (inputs(82));
    layer0_outputs(4975) <= (inputs(108)) xor (inputs(66));
    layer0_outputs(4976) <= not(inputs(236));
    layer0_outputs(4977) <= inputs(195);
    layer0_outputs(4978) <= inputs(45);
    layer0_outputs(4979) <= (inputs(82)) or (inputs(155));
    layer0_outputs(4980) <= (inputs(131)) and (inputs(208));
    layer0_outputs(4981) <= not(inputs(28));
    layer0_outputs(4982) <= (inputs(104)) or (inputs(129));
    layer0_outputs(4983) <= not((inputs(251)) or (inputs(118)));
    layer0_outputs(4984) <= (inputs(86)) and not (inputs(254));
    layer0_outputs(4985) <= (inputs(155)) or (inputs(43));
    layer0_outputs(4986) <= inputs(16);
    layer0_outputs(4987) <= not((inputs(249)) or (inputs(126)));
    layer0_outputs(4988) <= not((inputs(109)) xor (inputs(106)));
    layer0_outputs(4989) <= not(inputs(12));
    layer0_outputs(4990) <= (inputs(140)) or (inputs(242));
    layer0_outputs(4991) <= (inputs(85)) xor (inputs(207));
    layer0_outputs(4992) <= not(inputs(53));
    layer0_outputs(4993) <= (inputs(229)) and not (inputs(208));
    layer0_outputs(4994) <= not(inputs(71)) or (inputs(142));
    layer0_outputs(4995) <= inputs(36);
    layer0_outputs(4996) <= (inputs(69)) and not (inputs(230));
    layer0_outputs(4997) <= not(inputs(69)) or (inputs(196));
    layer0_outputs(4998) <= not((inputs(191)) or (inputs(111)));
    layer0_outputs(4999) <= not((inputs(83)) or (inputs(65)));
    layer0_outputs(5000) <= (inputs(138)) xor (inputs(153));
    layer0_outputs(5001) <= not(inputs(220));
    layer0_outputs(5002) <= (inputs(98)) and not (inputs(19));
    layer0_outputs(5003) <= not(inputs(104));
    layer0_outputs(5004) <= (inputs(88)) and not (inputs(63));
    layer0_outputs(5005) <= (inputs(149)) or (inputs(234));
    layer0_outputs(5006) <= (inputs(61)) and not (inputs(16));
    layer0_outputs(5007) <= inputs(209);
    layer0_outputs(5008) <= inputs(149);
    layer0_outputs(5009) <= not(inputs(214));
    layer0_outputs(5010) <= not(inputs(86));
    layer0_outputs(5011) <= '1';
    layer0_outputs(5012) <= (inputs(36)) and not (inputs(127));
    layer0_outputs(5013) <= (inputs(171)) and (inputs(183));
    layer0_outputs(5014) <= not(inputs(179));
    layer0_outputs(5015) <= inputs(164);
    layer0_outputs(5016) <= (inputs(233)) and not (inputs(28));
    layer0_outputs(5017) <= not((inputs(177)) xor (inputs(226)));
    layer0_outputs(5018) <= not(inputs(103));
    layer0_outputs(5019) <= (inputs(82)) and (inputs(114));
    layer0_outputs(5020) <= inputs(3);
    layer0_outputs(5021) <= not((inputs(130)) xor (inputs(107)));
    layer0_outputs(5022) <= (inputs(201)) and (inputs(236));
    layer0_outputs(5023) <= not((inputs(5)) xor (inputs(15)));
    layer0_outputs(5024) <= (inputs(234)) and (inputs(229));
    layer0_outputs(5025) <= (inputs(4)) or (inputs(227));
    layer0_outputs(5026) <= not((inputs(143)) or (inputs(68)));
    layer0_outputs(5027) <= not((inputs(61)) xor (inputs(28)));
    layer0_outputs(5028) <= not(inputs(72)) or (inputs(126));
    layer0_outputs(5029) <= not((inputs(213)) or (inputs(62)));
    layer0_outputs(5030) <= not(inputs(196));
    layer0_outputs(5031) <= (inputs(185)) and (inputs(188));
    layer0_outputs(5032) <= (inputs(242)) xor (inputs(65));
    layer0_outputs(5033) <= not((inputs(25)) xor (inputs(43)));
    layer0_outputs(5034) <= not(inputs(104)) or (inputs(14));
    layer0_outputs(5035) <= not(inputs(247)) or (inputs(110));
    layer0_outputs(5036) <= not((inputs(102)) or (inputs(133)));
    layer0_outputs(5037) <= inputs(106);
    layer0_outputs(5038) <= not(inputs(205));
    layer0_outputs(5039) <= not(inputs(20));
    layer0_outputs(5040) <= inputs(246);
    layer0_outputs(5041) <= (inputs(186)) and not (inputs(108));
    layer0_outputs(5042) <= inputs(208);
    layer0_outputs(5043) <= not(inputs(247));
    layer0_outputs(5044) <= (inputs(201)) xor (inputs(247));
    layer0_outputs(5045) <= not(inputs(243)) or (inputs(105));
    layer0_outputs(5046) <= (inputs(167)) and (inputs(160));
    layer0_outputs(5047) <= not(inputs(195));
    layer0_outputs(5048) <= inputs(27);
    layer0_outputs(5049) <= (inputs(75)) xor (inputs(177));
    layer0_outputs(5050) <= not(inputs(32));
    layer0_outputs(5051) <= not((inputs(234)) xor (inputs(162)));
    layer0_outputs(5052) <= not(inputs(121)) or (inputs(192));
    layer0_outputs(5053) <= inputs(100);
    layer0_outputs(5054) <= (inputs(127)) xor (inputs(152));
    layer0_outputs(5055) <= not((inputs(13)) xor (inputs(176)));
    layer0_outputs(5056) <= not((inputs(25)) or (inputs(112)));
    layer0_outputs(5057) <= inputs(229);
    layer0_outputs(5058) <= not(inputs(74));
    layer0_outputs(5059) <= (inputs(52)) and not (inputs(32));
    layer0_outputs(5060) <= not((inputs(150)) and (inputs(183)));
    layer0_outputs(5061) <= (inputs(70)) and not (inputs(106));
    layer0_outputs(5062) <= (inputs(231)) and (inputs(134));
    layer0_outputs(5063) <= (inputs(151)) and not (inputs(100));
    layer0_outputs(5064) <= (inputs(215)) xor (inputs(153));
    layer0_outputs(5065) <= not(inputs(151)) or (inputs(215));
    layer0_outputs(5066) <= not(inputs(35)) or (inputs(128));
    layer0_outputs(5067) <= (inputs(113)) and not (inputs(27));
    layer0_outputs(5068) <= inputs(92);
    layer0_outputs(5069) <= not(inputs(123)) or (inputs(208));
    layer0_outputs(5070) <= not((inputs(158)) or (inputs(16)));
    layer0_outputs(5071) <= (inputs(201)) or (inputs(157));
    layer0_outputs(5072) <= inputs(210);
    layer0_outputs(5073) <= not((inputs(248)) or (inputs(142)));
    layer0_outputs(5074) <= inputs(55);
    layer0_outputs(5075) <= (inputs(129)) xor (inputs(101));
    layer0_outputs(5076) <= not((inputs(6)) xor (inputs(205)));
    layer0_outputs(5077) <= (inputs(37)) and not (inputs(127));
    layer0_outputs(5078) <= not((inputs(50)) or (inputs(122)));
    layer0_outputs(5079) <= not((inputs(14)) or (inputs(96)));
    layer0_outputs(5080) <= (inputs(105)) xor (inputs(177));
    layer0_outputs(5081) <= not((inputs(186)) or (inputs(115)));
    layer0_outputs(5082) <= (inputs(66)) and not (inputs(143));
    layer0_outputs(5083) <= inputs(89);
    layer0_outputs(5084) <= inputs(142);
    layer0_outputs(5085) <= inputs(169);
    layer0_outputs(5086) <= (inputs(161)) and not (inputs(95));
    layer0_outputs(5087) <= inputs(128);
    layer0_outputs(5088) <= inputs(139);
    layer0_outputs(5089) <= not((inputs(238)) or (inputs(227)));
    layer0_outputs(5090) <= not(inputs(92));
    layer0_outputs(5091) <= (inputs(115)) xor (inputs(64));
    layer0_outputs(5092) <= not(inputs(116)) or (inputs(104));
    layer0_outputs(5093) <= (inputs(217)) and (inputs(0));
    layer0_outputs(5094) <= not(inputs(116)) or (inputs(49));
    layer0_outputs(5095) <= not(inputs(156));
    layer0_outputs(5096) <= inputs(69);
    layer0_outputs(5097) <= inputs(151);
    layer0_outputs(5098) <= (inputs(112)) xor (inputs(156));
    layer0_outputs(5099) <= not(inputs(133)) or (inputs(252));
    layer0_outputs(5100) <= not((inputs(93)) or (inputs(178)));
    layer0_outputs(5101) <= not((inputs(40)) xor (inputs(8)));
    layer0_outputs(5102) <= (inputs(133)) xor (inputs(8));
    layer0_outputs(5103) <= not((inputs(114)) or (inputs(184)));
    layer0_outputs(5104) <= not((inputs(89)) xor (inputs(43)));
    layer0_outputs(5105) <= inputs(113);
    layer0_outputs(5106) <= (inputs(116)) and not (inputs(16));
    layer0_outputs(5107) <= not(inputs(20)) or (inputs(47));
    layer0_outputs(5108) <= (inputs(31)) or (inputs(43));
    layer0_outputs(5109) <= inputs(153);
    layer0_outputs(5110) <= inputs(163);
    layer0_outputs(5111) <= inputs(41);
    layer0_outputs(5112) <= not((inputs(164)) or (inputs(226)));
    layer0_outputs(5113) <= inputs(58);
    layer0_outputs(5114) <= (inputs(54)) xor (inputs(64));
    layer0_outputs(5115) <= not(inputs(129));
    layer0_outputs(5116) <= not((inputs(219)) or (inputs(96)));
    layer0_outputs(5117) <= (inputs(198)) and not (inputs(88));
    layer0_outputs(5118) <= not(inputs(231));
    layer0_outputs(5119) <= not((inputs(134)) xor (inputs(182)));
    layer0_outputs(5120) <= not(inputs(178));
    layer0_outputs(5121) <= (inputs(82)) or (inputs(90));
    layer0_outputs(5122) <= not(inputs(231));
    layer0_outputs(5123) <= (inputs(42)) and not (inputs(0));
    layer0_outputs(5124) <= not(inputs(178));
    layer0_outputs(5125) <= (inputs(23)) xor (inputs(160));
    layer0_outputs(5126) <= not(inputs(152));
    layer0_outputs(5127) <= '1';
    layer0_outputs(5128) <= (inputs(165)) and not (inputs(96));
    layer0_outputs(5129) <= not(inputs(100)) or (inputs(49));
    layer0_outputs(5130) <= inputs(137);
    layer0_outputs(5131) <= (inputs(9)) or (inputs(179));
    layer0_outputs(5132) <= not((inputs(187)) xor (inputs(137)));
    layer0_outputs(5133) <= not((inputs(58)) and (inputs(245)));
    layer0_outputs(5134) <= (inputs(66)) or (inputs(164));
    layer0_outputs(5135) <= inputs(233);
    layer0_outputs(5136) <= (inputs(27)) xor (inputs(131));
    layer0_outputs(5137) <= not(inputs(20));
    layer0_outputs(5138) <= '1';
    layer0_outputs(5139) <= (inputs(98)) xor (inputs(84));
    layer0_outputs(5140) <= not(inputs(208));
    layer0_outputs(5141) <= inputs(153);
    layer0_outputs(5142) <= inputs(130);
    layer0_outputs(5143) <= not(inputs(231)) or (inputs(238));
    layer0_outputs(5144) <= (inputs(148)) xor (inputs(136));
    layer0_outputs(5145) <= not(inputs(103));
    layer0_outputs(5146) <= (inputs(77)) or (inputs(23));
    layer0_outputs(5147) <= (inputs(166)) and (inputs(187));
    layer0_outputs(5148) <= not(inputs(88));
    layer0_outputs(5149) <= (inputs(84)) and not (inputs(204));
    layer0_outputs(5150) <= (inputs(86)) xor (inputs(99));
    layer0_outputs(5151) <= not(inputs(81));
    layer0_outputs(5152) <= not((inputs(91)) xor (inputs(164)));
    layer0_outputs(5153) <= not(inputs(130));
    layer0_outputs(5154) <= inputs(73);
    layer0_outputs(5155) <= inputs(7);
    layer0_outputs(5156) <= (inputs(48)) or (inputs(202));
    layer0_outputs(5157) <= not(inputs(25));
    layer0_outputs(5158) <= not(inputs(181));
    layer0_outputs(5159) <= not((inputs(26)) xor (inputs(41)));
    layer0_outputs(5160) <= (inputs(137)) xor (inputs(167));
    layer0_outputs(5161) <= not(inputs(84)) or (inputs(177));
    layer0_outputs(5162) <= not(inputs(148));
    layer0_outputs(5163) <= (inputs(135)) and (inputs(235));
    layer0_outputs(5164) <= not((inputs(186)) or (inputs(215)));
    layer0_outputs(5165) <= inputs(19);
    layer0_outputs(5166) <= not(inputs(119)) or (inputs(173));
    layer0_outputs(5167) <= not(inputs(186)) or (inputs(47));
    layer0_outputs(5168) <= not((inputs(160)) or (inputs(170)));
    layer0_outputs(5169) <= not(inputs(131)) or (inputs(49));
    layer0_outputs(5170) <= (inputs(166)) or (inputs(154));
    layer0_outputs(5171) <= (inputs(63)) or (inputs(35));
    layer0_outputs(5172) <= not(inputs(198)) or (inputs(11));
    layer0_outputs(5173) <= not((inputs(206)) or (inputs(213)));
    layer0_outputs(5174) <= not(inputs(164));
    layer0_outputs(5175) <= not((inputs(250)) xor (inputs(55)));
    layer0_outputs(5176) <= inputs(101);
    layer0_outputs(5177) <= not(inputs(230));
    layer0_outputs(5178) <= not((inputs(30)) or (inputs(128)));
    layer0_outputs(5179) <= inputs(99);
    layer0_outputs(5180) <= inputs(15);
    layer0_outputs(5181) <= (inputs(131)) or (inputs(54));
    layer0_outputs(5182) <= not((inputs(243)) xor (inputs(22)));
    layer0_outputs(5183) <= inputs(194);
    layer0_outputs(5184) <= not(inputs(53));
    layer0_outputs(5185) <= not((inputs(147)) and (inputs(139)));
    layer0_outputs(5186) <= inputs(196);
    layer0_outputs(5187) <= (inputs(39)) and not (inputs(230));
    layer0_outputs(5188) <= not((inputs(182)) or (inputs(245)));
    layer0_outputs(5189) <= (inputs(104)) xor (inputs(193));
    layer0_outputs(5190) <= '1';
    layer0_outputs(5191) <= inputs(52);
    layer0_outputs(5192) <= (inputs(156)) xor (inputs(4));
    layer0_outputs(5193) <= not(inputs(217));
    layer0_outputs(5194) <= not((inputs(164)) or (inputs(252)));
    layer0_outputs(5195) <= not((inputs(247)) or (inputs(174)));
    layer0_outputs(5196) <= (inputs(189)) and not (inputs(161));
    layer0_outputs(5197) <= not(inputs(192));
    layer0_outputs(5198) <= (inputs(27)) and not (inputs(166));
    layer0_outputs(5199) <= inputs(104);
    layer0_outputs(5200) <= (inputs(210)) and not (inputs(96));
    layer0_outputs(5201) <= not(inputs(26)) or (inputs(112));
    layer0_outputs(5202) <= not(inputs(119));
    layer0_outputs(5203) <= not((inputs(36)) or (inputs(91)));
    layer0_outputs(5204) <= (inputs(59)) xor (inputs(73));
    layer0_outputs(5205) <= (inputs(216)) xor (inputs(195));
    layer0_outputs(5206) <= not(inputs(249)) or (inputs(54));
    layer0_outputs(5207) <= not(inputs(54)) or (inputs(144));
    layer0_outputs(5208) <= inputs(75);
    layer0_outputs(5209) <= not(inputs(53)) or (inputs(205));
    layer0_outputs(5210) <= not(inputs(20));
    layer0_outputs(5211) <= (inputs(65)) or (inputs(138));
    layer0_outputs(5212) <= not(inputs(105));
    layer0_outputs(5213) <= not(inputs(23));
    layer0_outputs(5214) <= not(inputs(114));
    layer0_outputs(5215) <= not(inputs(154)) or (inputs(27));
    layer0_outputs(5216) <= not(inputs(137));
    layer0_outputs(5217) <= not(inputs(3)) or (inputs(128));
    layer0_outputs(5218) <= not(inputs(7));
    layer0_outputs(5219) <= not(inputs(54)) or (inputs(34));
    layer0_outputs(5220) <= not((inputs(226)) or (inputs(21)));
    layer0_outputs(5221) <= inputs(129);
    layer0_outputs(5222) <= not((inputs(255)) xor (inputs(163)));
    layer0_outputs(5223) <= (inputs(209)) or (inputs(118));
    layer0_outputs(5224) <= not(inputs(126));
    layer0_outputs(5225) <= not((inputs(190)) or (inputs(204)));
    layer0_outputs(5226) <= not(inputs(145));
    layer0_outputs(5227) <= not(inputs(42));
    layer0_outputs(5228) <= (inputs(187)) or (inputs(207));
    layer0_outputs(5229) <= not((inputs(227)) or (inputs(219)));
    layer0_outputs(5230) <= (inputs(216)) or (inputs(216));
    layer0_outputs(5231) <= (inputs(169)) and not (inputs(50));
    layer0_outputs(5232) <= (inputs(209)) or (inputs(237));
    layer0_outputs(5233) <= inputs(52);
    layer0_outputs(5234) <= not(inputs(207)) or (inputs(223));
    layer0_outputs(5235) <= inputs(174);
    layer0_outputs(5236) <= not((inputs(204)) xor (inputs(240)));
    layer0_outputs(5237) <= '1';
    layer0_outputs(5238) <= not((inputs(63)) xor (inputs(156)));
    layer0_outputs(5239) <= not(inputs(152));
    layer0_outputs(5240) <= (inputs(231)) and not (inputs(126));
    layer0_outputs(5241) <= not((inputs(196)) xor (inputs(27)));
    layer0_outputs(5242) <= not((inputs(174)) xor (inputs(107)));
    layer0_outputs(5243) <= '1';
    layer0_outputs(5244) <= not((inputs(63)) xor (inputs(199)));
    layer0_outputs(5245) <= not(inputs(230));
    layer0_outputs(5246) <= not((inputs(145)) or (inputs(160)));
    layer0_outputs(5247) <= not((inputs(204)) xor (inputs(225)));
    layer0_outputs(5248) <= not((inputs(65)) or (inputs(179)));
    layer0_outputs(5249) <= (inputs(177)) xor (inputs(144));
    layer0_outputs(5250) <= not(inputs(30));
    layer0_outputs(5251) <= not((inputs(104)) or (inputs(163)));
    layer0_outputs(5252) <= not((inputs(196)) xor (inputs(10)));
    layer0_outputs(5253) <= not(inputs(57)) or (inputs(149));
    layer0_outputs(5254) <= (inputs(68)) xor (inputs(133));
    layer0_outputs(5255) <= not((inputs(21)) or (inputs(43)));
    layer0_outputs(5256) <= (inputs(37)) and not (inputs(223));
    layer0_outputs(5257) <= (inputs(6)) and not (inputs(199));
    layer0_outputs(5258) <= (inputs(247)) or (inputs(88));
    layer0_outputs(5259) <= inputs(113);
    layer0_outputs(5260) <= not((inputs(63)) or (inputs(247)));
    layer0_outputs(5261) <= (inputs(176)) xor (inputs(190));
    layer0_outputs(5262) <= not((inputs(148)) or (inputs(141)));
    layer0_outputs(5263) <= inputs(205);
    layer0_outputs(5264) <= (inputs(52)) and not (inputs(250));
    layer0_outputs(5265) <= not(inputs(194));
    layer0_outputs(5266) <= (inputs(4)) xor (inputs(176));
    layer0_outputs(5267) <= (inputs(0)) and not (inputs(155));
    layer0_outputs(5268) <= (inputs(105)) or (inputs(243));
    layer0_outputs(5269) <= not(inputs(176));
    layer0_outputs(5270) <= (inputs(169)) or (inputs(237));
    layer0_outputs(5271) <= not((inputs(229)) or (inputs(182)));
    layer0_outputs(5272) <= not((inputs(187)) xor (inputs(149)));
    layer0_outputs(5273) <= not(inputs(93));
    layer0_outputs(5274) <= inputs(57);
    layer0_outputs(5275) <= not(inputs(17)) or (inputs(11));
    layer0_outputs(5276) <= (inputs(117)) or (inputs(163));
    layer0_outputs(5277) <= not(inputs(46)) or (inputs(208));
    layer0_outputs(5278) <= inputs(39);
    layer0_outputs(5279) <= not((inputs(53)) xor (inputs(114)));
    layer0_outputs(5280) <= not(inputs(19));
    layer0_outputs(5281) <= inputs(61);
    layer0_outputs(5282) <= inputs(103);
    layer0_outputs(5283) <= (inputs(107)) xor (inputs(90));
    layer0_outputs(5284) <= not((inputs(161)) or (inputs(17)));
    layer0_outputs(5285) <= not(inputs(100)) or (inputs(47));
    layer0_outputs(5286) <= (inputs(254)) or (inputs(252));
    layer0_outputs(5287) <= not((inputs(196)) or (inputs(80)));
    layer0_outputs(5288) <= not((inputs(159)) xor (inputs(31)));
    layer0_outputs(5289) <= not(inputs(138));
    layer0_outputs(5290) <= (inputs(68)) and not (inputs(220));
    layer0_outputs(5291) <= not(inputs(183));
    layer0_outputs(5292) <= not(inputs(181)) or (inputs(237));
    layer0_outputs(5293) <= not(inputs(227));
    layer0_outputs(5294) <= (inputs(245)) or (inputs(175));
    layer0_outputs(5295) <= (inputs(31)) and (inputs(84));
    layer0_outputs(5296) <= not(inputs(34));
    layer0_outputs(5297) <= not(inputs(175));
    layer0_outputs(5298) <= not((inputs(24)) or (inputs(127)));
    layer0_outputs(5299) <= not((inputs(197)) or (inputs(14)));
    layer0_outputs(5300) <= inputs(98);
    layer0_outputs(5301) <= (inputs(35)) or (inputs(140));
    layer0_outputs(5302) <= inputs(57);
    layer0_outputs(5303) <= not(inputs(210));
    layer0_outputs(5304) <= not(inputs(5)) or (inputs(225));
    layer0_outputs(5305) <= not(inputs(139)) or (inputs(248));
    layer0_outputs(5306) <= not(inputs(220));
    layer0_outputs(5307) <= (inputs(103)) and not (inputs(146));
    layer0_outputs(5308) <= not((inputs(177)) and (inputs(210)));
    layer0_outputs(5309) <= inputs(99);
    layer0_outputs(5310) <= (inputs(55)) or (inputs(139));
    layer0_outputs(5311) <= not(inputs(152)) or (inputs(55));
    layer0_outputs(5312) <= (inputs(230)) and (inputs(170));
    layer0_outputs(5313) <= not((inputs(224)) xor (inputs(12)));
    layer0_outputs(5314) <= not((inputs(141)) or (inputs(144)));
    layer0_outputs(5315) <= (inputs(62)) or (inputs(42));
    layer0_outputs(5316) <= not(inputs(184));
    layer0_outputs(5317) <= not(inputs(106));
    layer0_outputs(5318) <= inputs(209);
    layer0_outputs(5319) <= not(inputs(164)) or (inputs(50));
    layer0_outputs(5320) <= (inputs(48)) or (inputs(191));
    layer0_outputs(5321) <= not(inputs(90)) or (inputs(95));
    layer0_outputs(5322) <= not(inputs(253)) or (inputs(81));
    layer0_outputs(5323) <= (inputs(78)) and not (inputs(162));
    layer0_outputs(5324) <= not((inputs(144)) or (inputs(83)));
    layer0_outputs(5325) <= not((inputs(123)) or (inputs(70)));
    layer0_outputs(5326) <= (inputs(249)) or (inputs(1));
    layer0_outputs(5327) <= not(inputs(91));
    layer0_outputs(5328) <= (inputs(27)) and not (inputs(149));
    layer0_outputs(5329) <= (inputs(68)) xor (inputs(105));
    layer0_outputs(5330) <= inputs(40);
    layer0_outputs(5331) <= not(inputs(201)) or (inputs(25));
    layer0_outputs(5332) <= not((inputs(78)) and (inputs(79)));
    layer0_outputs(5333) <= not(inputs(38)) or (inputs(139));
    layer0_outputs(5334) <= not(inputs(95));
    layer0_outputs(5335) <= not((inputs(220)) xor (inputs(161)));
    layer0_outputs(5336) <= (inputs(77)) and not (inputs(49));
    layer0_outputs(5337) <= inputs(118);
    layer0_outputs(5338) <= not(inputs(149));
    layer0_outputs(5339) <= inputs(123);
    layer0_outputs(5340) <= not(inputs(99));
    layer0_outputs(5341) <= inputs(109);
    layer0_outputs(5342) <= (inputs(201)) or (inputs(137));
    layer0_outputs(5343) <= not(inputs(41));
    layer0_outputs(5344) <= not((inputs(125)) xor (inputs(240)));
    layer0_outputs(5345) <= (inputs(42)) or (inputs(2));
    layer0_outputs(5346) <= not((inputs(161)) or (inputs(29)));
    layer0_outputs(5347) <= not(inputs(186)) or (inputs(120));
    layer0_outputs(5348) <= inputs(86);
    layer0_outputs(5349) <= inputs(99);
    layer0_outputs(5350) <= (inputs(88)) or (inputs(194));
    layer0_outputs(5351) <= (inputs(185)) or (inputs(235));
    layer0_outputs(5352) <= (inputs(7)) and not (inputs(86));
    layer0_outputs(5353) <= (inputs(23)) and not (inputs(247));
    layer0_outputs(5354) <= inputs(137);
    layer0_outputs(5355) <= (inputs(61)) or (inputs(5));
    layer0_outputs(5356) <= not(inputs(84)) or (inputs(3));
    layer0_outputs(5357) <= not((inputs(96)) or (inputs(30)));
    layer0_outputs(5358) <= (inputs(139)) and (inputs(139));
    layer0_outputs(5359) <= (inputs(79)) and (inputs(31));
    layer0_outputs(5360) <= not(inputs(77));
    layer0_outputs(5361) <= (inputs(26)) and not (inputs(255));
    layer0_outputs(5362) <= not((inputs(175)) or (inputs(147)));
    layer0_outputs(5363) <= not((inputs(78)) xor (inputs(234)));
    layer0_outputs(5364) <= not(inputs(139)) or (inputs(234));
    layer0_outputs(5365) <= (inputs(136)) or (inputs(148));
    layer0_outputs(5366) <= not(inputs(244));
    layer0_outputs(5367) <= not(inputs(25));
    layer0_outputs(5368) <= (inputs(41)) and not (inputs(48));
    layer0_outputs(5369) <= not(inputs(29));
    layer0_outputs(5370) <= not((inputs(2)) xor (inputs(141)));
    layer0_outputs(5371) <= (inputs(102)) or (inputs(215));
    layer0_outputs(5372) <= (inputs(217)) xor (inputs(166));
    layer0_outputs(5373) <= (inputs(185)) or (inputs(80));
    layer0_outputs(5374) <= (inputs(105)) or (inputs(89));
    layer0_outputs(5375) <= not(inputs(82));
    layer0_outputs(5376) <= inputs(111);
    layer0_outputs(5377) <= inputs(99);
    layer0_outputs(5378) <= inputs(206);
    layer0_outputs(5379) <= (inputs(117)) and not (inputs(205));
    layer0_outputs(5380) <= inputs(174);
    layer0_outputs(5381) <= not(inputs(94));
    layer0_outputs(5382) <= (inputs(56)) and (inputs(244));
    layer0_outputs(5383) <= not(inputs(101)) or (inputs(93));
    layer0_outputs(5384) <= not((inputs(193)) or (inputs(174)));
    layer0_outputs(5385) <= (inputs(105)) and not (inputs(49));
    layer0_outputs(5386) <= (inputs(161)) or (inputs(146));
    layer0_outputs(5387) <= not(inputs(48)) or (inputs(141));
    layer0_outputs(5388) <= not(inputs(148));
    layer0_outputs(5389) <= inputs(178);
    layer0_outputs(5390) <= not(inputs(164));
    layer0_outputs(5391) <= not(inputs(85));
    layer0_outputs(5392) <= (inputs(141)) and not (inputs(92));
    layer0_outputs(5393) <= (inputs(207)) or (inputs(58));
    layer0_outputs(5394) <= inputs(101);
    layer0_outputs(5395) <= inputs(144);
    layer0_outputs(5396) <= (inputs(11)) xor (inputs(51));
    layer0_outputs(5397) <= not(inputs(18));
    layer0_outputs(5398) <= not(inputs(17)) or (inputs(238));
    layer0_outputs(5399) <= not((inputs(229)) or (inputs(191)));
    layer0_outputs(5400) <= not((inputs(66)) or (inputs(112)));
    layer0_outputs(5401) <= not((inputs(28)) or (inputs(34)));
    layer0_outputs(5402) <= (inputs(164)) or (inputs(86));
    layer0_outputs(5403) <= (inputs(211)) or (inputs(189));
    layer0_outputs(5404) <= not((inputs(95)) or (inputs(84)));
    layer0_outputs(5405) <= not(inputs(101));
    layer0_outputs(5406) <= inputs(239);
    layer0_outputs(5407) <= not((inputs(49)) or (inputs(63)));
    layer0_outputs(5408) <= (inputs(224)) and not (inputs(88));
    layer0_outputs(5409) <= not((inputs(83)) xor (inputs(71)));
    layer0_outputs(5410) <= (inputs(0)) or (inputs(128));
    layer0_outputs(5411) <= (inputs(247)) xor (inputs(62));
    layer0_outputs(5412) <= not((inputs(226)) and (inputs(95)));
    layer0_outputs(5413) <= (inputs(163)) and not (inputs(16));
    layer0_outputs(5414) <= not((inputs(253)) or (inputs(189)));
    layer0_outputs(5415) <= not((inputs(64)) or (inputs(255)));
    layer0_outputs(5416) <= inputs(121);
    layer0_outputs(5417) <= not((inputs(53)) xor (inputs(121)));
    layer0_outputs(5418) <= inputs(88);
    layer0_outputs(5419) <= inputs(76);
    layer0_outputs(5420) <= not((inputs(20)) xor (inputs(107)));
    layer0_outputs(5421) <= not(inputs(177)) or (inputs(43));
    layer0_outputs(5422) <= (inputs(85)) and not (inputs(156));
    layer0_outputs(5423) <= not(inputs(182)) or (inputs(45));
    layer0_outputs(5424) <= (inputs(220)) xor (inputs(1));
    layer0_outputs(5425) <= not(inputs(75));
    layer0_outputs(5426) <= not((inputs(201)) or (inputs(218)));
    layer0_outputs(5427) <= inputs(73);
    layer0_outputs(5428) <= (inputs(237)) or (inputs(149));
    layer0_outputs(5429) <= (inputs(141)) and not (inputs(37));
    layer0_outputs(5430) <= (inputs(193)) or (inputs(218));
    layer0_outputs(5431) <= (inputs(37)) and not (inputs(250));
    layer0_outputs(5432) <= inputs(105);
    layer0_outputs(5433) <= inputs(110);
    layer0_outputs(5434) <= (inputs(61)) and not (inputs(113));
    layer0_outputs(5435) <= not(inputs(255)) or (inputs(16));
    layer0_outputs(5436) <= not(inputs(246)) or (inputs(127));
    layer0_outputs(5437) <= '0';
    layer0_outputs(5438) <= inputs(180);
    layer0_outputs(5439) <= not(inputs(197));
    layer0_outputs(5440) <= not((inputs(208)) or (inputs(103)));
    layer0_outputs(5441) <= (inputs(138)) and not (inputs(119));
    layer0_outputs(5442) <= (inputs(22)) xor (inputs(34));
    layer0_outputs(5443) <= (inputs(183)) and not (inputs(238));
    layer0_outputs(5444) <= not(inputs(9)) or (inputs(180));
    layer0_outputs(5445) <= inputs(129);
    layer0_outputs(5446) <= (inputs(231)) xor (inputs(56));
    layer0_outputs(5447) <= not((inputs(51)) or (inputs(107)));
    layer0_outputs(5448) <= '1';
    layer0_outputs(5449) <= not(inputs(179));
    layer0_outputs(5450) <= not(inputs(169));
    layer0_outputs(5451) <= inputs(219);
    layer0_outputs(5452) <= not((inputs(49)) or (inputs(184)));
    layer0_outputs(5453) <= not(inputs(12));
    layer0_outputs(5454) <= (inputs(158)) or (inputs(195));
    layer0_outputs(5455) <= (inputs(67)) and not (inputs(203));
    layer0_outputs(5456) <= (inputs(202)) and not (inputs(113));
    layer0_outputs(5457) <= not(inputs(142)) or (inputs(237));
    layer0_outputs(5458) <= inputs(205);
    layer0_outputs(5459) <= (inputs(0)) xor (inputs(250));
    layer0_outputs(5460) <= (inputs(159)) or (inputs(212));
    layer0_outputs(5461) <= not(inputs(13)) or (inputs(111));
    layer0_outputs(5462) <= not(inputs(86));
    layer0_outputs(5463) <= (inputs(32)) or (inputs(55));
    layer0_outputs(5464) <= not(inputs(210));
    layer0_outputs(5465) <= (inputs(19)) or (inputs(39));
    layer0_outputs(5466) <= not((inputs(68)) and (inputs(133)));
    layer0_outputs(5467) <= (inputs(86)) xor (inputs(20));
    layer0_outputs(5468) <= inputs(85);
    layer0_outputs(5469) <= (inputs(209)) or (inputs(48));
    layer0_outputs(5470) <= not((inputs(24)) and (inputs(194)));
    layer0_outputs(5471) <= not((inputs(59)) xor (inputs(14)));
    layer0_outputs(5472) <= not((inputs(3)) xor (inputs(226)));
    layer0_outputs(5473) <= inputs(132);
    layer0_outputs(5474) <= (inputs(243)) and (inputs(240));
    layer0_outputs(5475) <= (inputs(76)) and not (inputs(108));
    layer0_outputs(5476) <= not(inputs(57));
    layer0_outputs(5477) <= inputs(229);
    layer0_outputs(5478) <= not(inputs(232));
    layer0_outputs(5479) <= not(inputs(219)) or (inputs(109));
    layer0_outputs(5480) <= inputs(143);
    layer0_outputs(5481) <= not(inputs(116));
    layer0_outputs(5482) <= not((inputs(21)) xor (inputs(35)));
    layer0_outputs(5483) <= inputs(86);
    layer0_outputs(5484) <= (inputs(4)) and not (inputs(62));
    layer0_outputs(5485) <= '1';
    layer0_outputs(5486) <= inputs(166);
    layer0_outputs(5487) <= inputs(94);
    layer0_outputs(5488) <= not(inputs(40));
    layer0_outputs(5489) <= not(inputs(216));
    layer0_outputs(5490) <= (inputs(9)) or (inputs(88));
    layer0_outputs(5491) <= (inputs(200)) and not (inputs(84));
    layer0_outputs(5492) <= inputs(225);
    layer0_outputs(5493) <= (inputs(30)) xor (inputs(61));
    layer0_outputs(5494) <= (inputs(214)) or (inputs(56));
    layer0_outputs(5495) <= (inputs(161)) or (inputs(164));
    layer0_outputs(5496) <= inputs(138);
    layer0_outputs(5497) <= not(inputs(119));
    layer0_outputs(5498) <= not((inputs(67)) or (inputs(65)));
    layer0_outputs(5499) <= not((inputs(179)) xor (inputs(121)));
    layer0_outputs(5500) <= not(inputs(132));
    layer0_outputs(5501) <= inputs(104);
    layer0_outputs(5502) <= not(inputs(120));
    layer0_outputs(5503) <= inputs(94);
    layer0_outputs(5504) <= not(inputs(183));
    layer0_outputs(5505) <= (inputs(143)) or (inputs(61));
    layer0_outputs(5506) <= not(inputs(56));
    layer0_outputs(5507) <= not((inputs(93)) or (inputs(121)));
    layer0_outputs(5508) <= not(inputs(105));
    layer0_outputs(5509) <= (inputs(42)) or (inputs(92));
    layer0_outputs(5510) <= not(inputs(85));
    layer0_outputs(5511) <= (inputs(140)) or (inputs(246));
    layer0_outputs(5512) <= not(inputs(180));
    layer0_outputs(5513) <= '0';
    layer0_outputs(5514) <= not(inputs(113));
    layer0_outputs(5515) <= (inputs(35)) or (inputs(2));
    layer0_outputs(5516) <= (inputs(2)) or (inputs(237));
    layer0_outputs(5517) <= not(inputs(45));
    layer0_outputs(5518) <= not(inputs(217)) or (inputs(141));
    layer0_outputs(5519) <= (inputs(237)) or (inputs(146));
    layer0_outputs(5520) <= not(inputs(215)) or (inputs(77));
    layer0_outputs(5521) <= not((inputs(115)) or (inputs(156)));
    layer0_outputs(5522) <= not(inputs(219));
    layer0_outputs(5523) <= inputs(137);
    layer0_outputs(5524) <= (inputs(229)) or (inputs(118));
    layer0_outputs(5525) <= (inputs(242)) and (inputs(228));
    layer0_outputs(5526) <= not((inputs(208)) or (inputs(242)));
    layer0_outputs(5527) <= (inputs(166)) xor (inputs(184));
    layer0_outputs(5528) <= not((inputs(34)) xor (inputs(111)));
    layer0_outputs(5529) <= not(inputs(68)) or (inputs(241));
    layer0_outputs(5530) <= not((inputs(92)) or (inputs(77)));
    layer0_outputs(5531) <= not(inputs(82));
    layer0_outputs(5532) <= not((inputs(68)) or (inputs(223)));
    layer0_outputs(5533) <= '0';
    layer0_outputs(5534) <= (inputs(74)) xor (inputs(77));
    layer0_outputs(5535) <= not(inputs(19));
    layer0_outputs(5536) <= (inputs(209)) or (inputs(216));
    layer0_outputs(5537) <= not((inputs(149)) xor (inputs(184)));
    layer0_outputs(5538) <= inputs(169);
    layer0_outputs(5539) <= not(inputs(105));
    layer0_outputs(5540) <= inputs(25);
    layer0_outputs(5541) <= not(inputs(195));
    layer0_outputs(5542) <= inputs(236);
    layer0_outputs(5543) <= (inputs(116)) and not (inputs(206));
    layer0_outputs(5544) <= not((inputs(236)) xor (inputs(62)));
    layer0_outputs(5545) <= (inputs(115)) or (inputs(115));
    layer0_outputs(5546) <= inputs(120);
    layer0_outputs(5547) <= inputs(252);
    layer0_outputs(5548) <= not(inputs(245));
    layer0_outputs(5549) <= not(inputs(218));
    layer0_outputs(5550) <= not((inputs(200)) xor (inputs(174)));
    layer0_outputs(5551) <= not(inputs(211)) or (inputs(196));
    layer0_outputs(5552) <= inputs(116);
    layer0_outputs(5553) <= not(inputs(103));
    layer0_outputs(5554) <= inputs(40);
    layer0_outputs(5555) <= not(inputs(190)) or (inputs(209));
    layer0_outputs(5556) <= (inputs(182)) xor (inputs(178));
    layer0_outputs(5557) <= not((inputs(28)) or (inputs(14)));
    layer0_outputs(5558) <= (inputs(190)) and not (inputs(29));
    layer0_outputs(5559) <= not((inputs(156)) and (inputs(17)));
    layer0_outputs(5560) <= not((inputs(7)) or (inputs(20)));
    layer0_outputs(5561) <= not(inputs(128));
    layer0_outputs(5562) <= not((inputs(4)) or (inputs(90)));
    layer0_outputs(5563) <= not((inputs(171)) and (inputs(134)));
    layer0_outputs(5564) <= inputs(68);
    layer0_outputs(5565) <= not(inputs(156)) or (inputs(237));
    layer0_outputs(5566) <= not(inputs(124));
    layer0_outputs(5567) <= not(inputs(87)) or (inputs(79));
    layer0_outputs(5568) <= (inputs(1)) or (inputs(220));
    layer0_outputs(5569) <= (inputs(45)) and not (inputs(96));
    layer0_outputs(5570) <= not(inputs(98));
    layer0_outputs(5571) <= (inputs(118)) xor (inputs(157));
    layer0_outputs(5572) <= (inputs(38)) and not (inputs(167));
    layer0_outputs(5573) <= inputs(163);
    layer0_outputs(5574) <= not(inputs(228)) or (inputs(118));
    layer0_outputs(5575) <= (inputs(242)) and not (inputs(202));
    layer0_outputs(5576) <= not((inputs(101)) xor (inputs(99)));
    layer0_outputs(5577) <= inputs(213);
    layer0_outputs(5578) <= not((inputs(221)) or (inputs(181)));
    layer0_outputs(5579) <= not(inputs(127)) or (inputs(221));
    layer0_outputs(5580) <= (inputs(29)) xor (inputs(237));
    layer0_outputs(5581) <= not(inputs(180));
    layer0_outputs(5582) <= inputs(26);
    layer0_outputs(5583) <= (inputs(166)) or (inputs(108));
    layer0_outputs(5584) <= (inputs(73)) xor (inputs(132));
    layer0_outputs(5585) <= (inputs(171)) or (inputs(33));
    layer0_outputs(5586) <= not(inputs(23));
    layer0_outputs(5587) <= not(inputs(184)) or (inputs(1));
    layer0_outputs(5588) <= not(inputs(30));
    layer0_outputs(5589) <= not(inputs(136));
    layer0_outputs(5590) <= not(inputs(234));
    layer0_outputs(5591) <= (inputs(86)) and not (inputs(111));
    layer0_outputs(5592) <= (inputs(122)) xor (inputs(170));
    layer0_outputs(5593) <= not((inputs(154)) and (inputs(122)));
    layer0_outputs(5594) <= (inputs(85)) and not (inputs(224));
    layer0_outputs(5595) <= (inputs(62)) and not (inputs(238));
    layer0_outputs(5596) <= (inputs(117)) or (inputs(239));
    layer0_outputs(5597) <= not(inputs(126));
    layer0_outputs(5598) <= (inputs(0)) and not (inputs(12));
    layer0_outputs(5599) <= not((inputs(33)) or (inputs(48)));
    layer0_outputs(5600) <= not(inputs(102)) or (inputs(242));
    layer0_outputs(5601) <= (inputs(15)) and not (inputs(61));
    layer0_outputs(5602) <= not(inputs(148)) or (inputs(253));
    layer0_outputs(5603) <= (inputs(14)) or (inputs(252));
    layer0_outputs(5604) <= not(inputs(99)) or (inputs(13));
    layer0_outputs(5605) <= not(inputs(142));
    layer0_outputs(5606) <= (inputs(174)) or (inputs(188));
    layer0_outputs(5607) <= not(inputs(204));
    layer0_outputs(5608) <= inputs(247);
    layer0_outputs(5609) <= (inputs(229)) and (inputs(165));
    layer0_outputs(5610) <= not((inputs(162)) or (inputs(145)));
    layer0_outputs(5611) <= not((inputs(77)) or (inputs(199)));
    layer0_outputs(5612) <= (inputs(96)) xor (inputs(104));
    layer0_outputs(5613) <= not(inputs(229));
    layer0_outputs(5614) <= not((inputs(116)) or (inputs(53)));
    layer0_outputs(5615) <= not((inputs(50)) or (inputs(83)));
    layer0_outputs(5616) <= not(inputs(44)) or (inputs(47));
    layer0_outputs(5617) <= not(inputs(209)) or (inputs(191));
    layer0_outputs(5618) <= not((inputs(97)) or (inputs(53)));
    layer0_outputs(5619) <= not((inputs(163)) xor (inputs(190)));
    layer0_outputs(5620) <= (inputs(93)) and (inputs(27));
    layer0_outputs(5621) <= (inputs(132)) and not (inputs(224));
    layer0_outputs(5622) <= (inputs(5)) and (inputs(181));
    layer0_outputs(5623) <= inputs(93);
    layer0_outputs(5624) <= not(inputs(82));
    layer0_outputs(5625) <= not(inputs(97));
    layer0_outputs(5626) <= (inputs(20)) and not (inputs(250));
    layer0_outputs(5627) <= inputs(185);
    layer0_outputs(5628) <= not((inputs(239)) or (inputs(166)));
    layer0_outputs(5629) <= not((inputs(233)) or (inputs(209)));
    layer0_outputs(5630) <= not((inputs(28)) xor (inputs(27)));
    layer0_outputs(5631) <= (inputs(226)) xor (inputs(96));
    layer0_outputs(5632) <= (inputs(9)) and not (inputs(161));
    layer0_outputs(5633) <= inputs(188);
    layer0_outputs(5634) <= (inputs(185)) or (inputs(4));
    layer0_outputs(5635) <= not((inputs(235)) or (inputs(9)));
    layer0_outputs(5636) <= not((inputs(127)) or (inputs(50)));
    layer0_outputs(5637) <= (inputs(73)) and not (inputs(109));
    layer0_outputs(5638) <= not(inputs(164)) or (inputs(63));
    layer0_outputs(5639) <= (inputs(151)) xor (inputs(237));
    layer0_outputs(5640) <= not(inputs(148));
    layer0_outputs(5641) <= not(inputs(217)) or (inputs(94));
    layer0_outputs(5642) <= (inputs(55)) and not (inputs(180));
    layer0_outputs(5643) <= (inputs(129)) xor (inputs(48));
    layer0_outputs(5644) <= not((inputs(102)) or (inputs(203)));
    layer0_outputs(5645) <= not((inputs(200)) or (inputs(200)));
    layer0_outputs(5646) <= not((inputs(254)) or (inputs(199)));
    layer0_outputs(5647) <= (inputs(171)) and not (inputs(50));
    layer0_outputs(5648) <= (inputs(171)) and not (inputs(96));
    layer0_outputs(5649) <= inputs(117);
    layer0_outputs(5650) <= inputs(67);
    layer0_outputs(5651) <= (inputs(254)) xor (inputs(118));
    layer0_outputs(5652) <= inputs(23);
    layer0_outputs(5653) <= not((inputs(115)) and (inputs(196)));
    layer0_outputs(5654) <= (inputs(186)) xor (inputs(138));
    layer0_outputs(5655) <= inputs(250);
    layer0_outputs(5656) <= inputs(195);
    layer0_outputs(5657) <= not((inputs(191)) or (inputs(75)));
    layer0_outputs(5658) <= '1';
    layer0_outputs(5659) <= not(inputs(23)) or (inputs(227));
    layer0_outputs(5660) <= not(inputs(102));
    layer0_outputs(5661) <= (inputs(80)) or (inputs(12));
    layer0_outputs(5662) <= (inputs(71)) or (inputs(48));
    layer0_outputs(5663) <= not(inputs(185)) or (inputs(133));
    layer0_outputs(5664) <= '0';
    layer0_outputs(5665) <= inputs(41);
    layer0_outputs(5666) <= not(inputs(42));
    layer0_outputs(5667) <= not(inputs(21));
    layer0_outputs(5668) <= (inputs(209)) or (inputs(101));
    layer0_outputs(5669) <= not(inputs(151));
    layer0_outputs(5670) <= not(inputs(179)) or (inputs(94));
    layer0_outputs(5671) <= (inputs(134)) or (inputs(222));
    layer0_outputs(5672) <= not((inputs(156)) xor (inputs(213)));
    layer0_outputs(5673) <= (inputs(69)) or (inputs(38));
    layer0_outputs(5674) <= not((inputs(175)) or (inputs(64)));
    layer0_outputs(5675) <= not((inputs(56)) and (inputs(109)));
    layer0_outputs(5676) <= (inputs(14)) or (inputs(239));
    layer0_outputs(5677) <= (inputs(216)) xor (inputs(59));
    layer0_outputs(5678) <= inputs(177);
    layer0_outputs(5679) <= inputs(84);
    layer0_outputs(5680) <= not((inputs(226)) xor (inputs(180)));
    layer0_outputs(5681) <= not(inputs(90));
    layer0_outputs(5682) <= (inputs(207)) xor (inputs(236));
    layer0_outputs(5683) <= not(inputs(88)) or (inputs(129));
    layer0_outputs(5684) <= (inputs(231)) or (inputs(185));
    layer0_outputs(5685) <= not((inputs(119)) xor (inputs(232)));
    layer0_outputs(5686) <= not((inputs(228)) or (inputs(212)));
    layer0_outputs(5687) <= inputs(79);
    layer0_outputs(5688) <= (inputs(138)) and not (inputs(200));
    layer0_outputs(5689) <= (inputs(202)) and not (inputs(120));
    layer0_outputs(5690) <= (inputs(198)) and not (inputs(118));
    layer0_outputs(5691) <= inputs(29);
    layer0_outputs(5692) <= not(inputs(69));
    layer0_outputs(5693) <= inputs(218);
    layer0_outputs(5694) <= inputs(216);
    layer0_outputs(5695) <= '0';
    layer0_outputs(5696) <= '0';
    layer0_outputs(5697) <= not(inputs(233));
    layer0_outputs(5698) <= (inputs(86)) or (inputs(149));
    layer0_outputs(5699) <= inputs(104);
    layer0_outputs(5700) <= (inputs(9)) and (inputs(76));
    layer0_outputs(5701) <= (inputs(10)) or (inputs(61));
    layer0_outputs(5702) <= not((inputs(45)) xor (inputs(75)));
    layer0_outputs(5703) <= inputs(157);
    layer0_outputs(5704) <= (inputs(139)) or (inputs(178));
    layer0_outputs(5705) <= (inputs(110)) or (inputs(3));
    layer0_outputs(5706) <= (inputs(238)) and not (inputs(130));
    layer0_outputs(5707) <= inputs(113);
    layer0_outputs(5708) <= not(inputs(117)) or (inputs(35));
    layer0_outputs(5709) <= (inputs(0)) and not (inputs(241));
    layer0_outputs(5710) <= (inputs(55)) and not (inputs(204));
    layer0_outputs(5711) <= inputs(229);
    layer0_outputs(5712) <= not(inputs(97));
    layer0_outputs(5713) <= (inputs(22)) or (inputs(228));
    layer0_outputs(5714) <= not((inputs(246)) or (inputs(42)));
    layer0_outputs(5715) <= (inputs(226)) and (inputs(236));
    layer0_outputs(5716) <= not(inputs(181));
    layer0_outputs(5717) <= inputs(24);
    layer0_outputs(5718) <= (inputs(167)) xor (inputs(120));
    layer0_outputs(5719) <= (inputs(186)) xor (inputs(185));
    layer0_outputs(5720) <= (inputs(163)) and not (inputs(231));
    layer0_outputs(5721) <= not(inputs(12)) or (inputs(253));
    layer0_outputs(5722) <= (inputs(32)) xor (inputs(6));
    layer0_outputs(5723) <= inputs(136);
    layer0_outputs(5724) <= (inputs(36)) or (inputs(63));
    layer0_outputs(5725) <= not((inputs(106)) xor (inputs(95)));
    layer0_outputs(5726) <= not(inputs(187)) or (inputs(125));
    layer0_outputs(5727) <= (inputs(242)) xor (inputs(53));
    layer0_outputs(5728) <= (inputs(111)) and not (inputs(254));
    layer0_outputs(5729) <= not(inputs(137)) or (inputs(47));
    layer0_outputs(5730) <= not(inputs(35)) or (inputs(129));
    layer0_outputs(5731) <= (inputs(204)) or (inputs(20));
    layer0_outputs(5732) <= (inputs(7)) xor (inputs(210));
    layer0_outputs(5733) <= inputs(60);
    layer0_outputs(5734) <= not(inputs(194));
    layer0_outputs(5735) <= (inputs(155)) xor (inputs(110));
    layer0_outputs(5736) <= (inputs(26)) and not (inputs(222));
    layer0_outputs(5737) <= inputs(165);
    layer0_outputs(5738) <= not((inputs(79)) or (inputs(36)));
    layer0_outputs(5739) <= inputs(224);
    layer0_outputs(5740) <= inputs(168);
    layer0_outputs(5741) <= (inputs(248)) and not (inputs(95));
    layer0_outputs(5742) <= not(inputs(29)) or (inputs(180));
    layer0_outputs(5743) <= not((inputs(130)) or (inputs(144)));
    layer0_outputs(5744) <= '0';
    layer0_outputs(5745) <= not((inputs(233)) xor (inputs(161)));
    layer0_outputs(5746) <= (inputs(107)) or (inputs(175));
    layer0_outputs(5747) <= (inputs(218)) or (inputs(248));
    layer0_outputs(5748) <= not(inputs(87));
    layer0_outputs(5749) <= not(inputs(220));
    layer0_outputs(5750) <= (inputs(37)) and not (inputs(181));
    layer0_outputs(5751) <= inputs(210);
    layer0_outputs(5752) <= not((inputs(150)) or (inputs(18)));
    layer0_outputs(5753) <= not(inputs(82));
    layer0_outputs(5754) <= not(inputs(106));
    layer0_outputs(5755) <= inputs(101);
    layer0_outputs(5756) <= not(inputs(200));
    layer0_outputs(5757) <= (inputs(80)) xor (inputs(163));
    layer0_outputs(5758) <= inputs(164);
    layer0_outputs(5759) <= not((inputs(95)) or (inputs(39)));
    layer0_outputs(5760) <= not(inputs(120));
    layer0_outputs(5761) <= not((inputs(137)) xor (inputs(107)));
    layer0_outputs(5762) <= not((inputs(196)) or (inputs(141)));
    layer0_outputs(5763) <= not((inputs(255)) xor (inputs(31)));
    layer0_outputs(5764) <= inputs(115);
    layer0_outputs(5765) <= '1';
    layer0_outputs(5766) <= not(inputs(125));
    layer0_outputs(5767) <= inputs(94);
    layer0_outputs(5768) <= not((inputs(254)) or (inputs(227)));
    layer0_outputs(5769) <= inputs(195);
    layer0_outputs(5770) <= inputs(243);
    layer0_outputs(5771) <= not(inputs(185));
    layer0_outputs(5772) <= (inputs(117)) or (inputs(114));
    layer0_outputs(5773) <= not((inputs(102)) xor (inputs(49)));
    layer0_outputs(5774) <= not(inputs(99));
    layer0_outputs(5775) <= (inputs(188)) or (inputs(107));
    layer0_outputs(5776) <= '1';
    layer0_outputs(5777) <= not((inputs(239)) xor (inputs(21)));
    layer0_outputs(5778) <= inputs(173);
    layer0_outputs(5779) <= (inputs(65)) or (inputs(134));
    layer0_outputs(5780) <= not(inputs(4)) or (inputs(145));
    layer0_outputs(5781) <= (inputs(142)) and not (inputs(239));
    layer0_outputs(5782) <= not((inputs(146)) xor (inputs(231)));
    layer0_outputs(5783) <= not(inputs(230));
    layer0_outputs(5784) <= (inputs(97)) xor (inputs(255));
    layer0_outputs(5785) <= (inputs(216)) and (inputs(30));
    layer0_outputs(5786) <= not(inputs(124)) or (inputs(111));
    layer0_outputs(5787) <= not(inputs(151));
    layer0_outputs(5788) <= not((inputs(0)) xor (inputs(141)));
    layer0_outputs(5789) <= (inputs(10)) and not (inputs(226));
    layer0_outputs(5790) <= inputs(166);
    layer0_outputs(5791) <= not(inputs(196)) or (inputs(113));
    layer0_outputs(5792) <= not((inputs(62)) xor (inputs(205)));
    layer0_outputs(5793) <= (inputs(43)) and not (inputs(241));
    layer0_outputs(5794) <= inputs(6);
    layer0_outputs(5795) <= not(inputs(108));
    layer0_outputs(5796) <= not((inputs(108)) or (inputs(58)));
    layer0_outputs(5797) <= inputs(135);
    layer0_outputs(5798) <= (inputs(77)) or (inputs(146));
    layer0_outputs(5799) <= inputs(26);
    layer0_outputs(5800) <= inputs(191);
    layer0_outputs(5801) <= not(inputs(107));
    layer0_outputs(5802) <= not(inputs(203)) or (inputs(122));
    layer0_outputs(5803) <= not((inputs(69)) xor (inputs(200)));
    layer0_outputs(5804) <= (inputs(3)) xor (inputs(70));
    layer0_outputs(5805) <= not((inputs(216)) or (inputs(17)));
    layer0_outputs(5806) <= not(inputs(46)) or (inputs(33));
    layer0_outputs(5807) <= (inputs(161)) or (inputs(232));
    layer0_outputs(5808) <= not((inputs(207)) or (inputs(26)));
    layer0_outputs(5809) <= (inputs(245)) and not (inputs(166));
    layer0_outputs(5810) <= (inputs(72)) or (inputs(232));
    layer0_outputs(5811) <= not((inputs(169)) and (inputs(228)));
    layer0_outputs(5812) <= (inputs(73)) and not (inputs(183));
    layer0_outputs(5813) <= (inputs(7)) or (inputs(205));
    layer0_outputs(5814) <= inputs(102);
    layer0_outputs(5815) <= inputs(243);
    layer0_outputs(5816) <= not(inputs(202)) or (inputs(93));
    layer0_outputs(5817) <= not(inputs(126));
    layer0_outputs(5818) <= (inputs(34)) xor (inputs(80));
    layer0_outputs(5819) <= not(inputs(225));
    layer0_outputs(5820) <= not(inputs(158)) or (inputs(15));
    layer0_outputs(5821) <= not(inputs(154)) or (inputs(254));
    layer0_outputs(5822) <= (inputs(23)) xor (inputs(126));
    layer0_outputs(5823) <= inputs(62);
    layer0_outputs(5824) <= not((inputs(199)) or (inputs(244)));
    layer0_outputs(5825) <= not(inputs(228));
    layer0_outputs(5826) <= inputs(114);
    layer0_outputs(5827) <= not((inputs(95)) or (inputs(240)));
    layer0_outputs(5828) <= (inputs(113)) or (inputs(72));
    layer0_outputs(5829) <= not((inputs(250)) xor (inputs(169)));
    layer0_outputs(5830) <= not(inputs(26)) or (inputs(164));
    layer0_outputs(5831) <= not(inputs(167)) or (inputs(39));
    layer0_outputs(5832) <= (inputs(14)) and not (inputs(209));
    layer0_outputs(5833) <= inputs(222);
    layer0_outputs(5834) <= not(inputs(71));
    layer0_outputs(5835) <= inputs(116);
    layer0_outputs(5836) <= (inputs(46)) and not (inputs(89));
    layer0_outputs(5837) <= inputs(153);
    layer0_outputs(5838) <= inputs(17);
    layer0_outputs(5839) <= not((inputs(191)) xor (inputs(148)));
    layer0_outputs(5840) <= inputs(148);
    layer0_outputs(5841) <= (inputs(142)) or (inputs(222));
    layer0_outputs(5842) <= not(inputs(167)) or (inputs(193));
    layer0_outputs(5843) <= not(inputs(247)) or (inputs(182));
    layer0_outputs(5844) <= (inputs(248)) or (inputs(28));
    layer0_outputs(5845) <= inputs(140);
    layer0_outputs(5846) <= (inputs(30)) xor (inputs(53));
    layer0_outputs(5847) <= inputs(55);
    layer0_outputs(5848) <= (inputs(188)) and not (inputs(55));
    layer0_outputs(5849) <= not((inputs(143)) and (inputs(96)));
    layer0_outputs(5850) <= not((inputs(24)) xor (inputs(65)));
    layer0_outputs(5851) <= (inputs(228)) or (inputs(3));
    layer0_outputs(5852) <= (inputs(128)) or (inputs(67));
    layer0_outputs(5853) <= not(inputs(130)) or (inputs(11));
    layer0_outputs(5854) <= not((inputs(57)) or (inputs(42)));
    layer0_outputs(5855) <= not((inputs(99)) or (inputs(113)));
    layer0_outputs(5856) <= not(inputs(149));
    layer0_outputs(5857) <= not(inputs(20));
    layer0_outputs(5858) <= (inputs(206)) xor (inputs(92));
    layer0_outputs(5859) <= (inputs(9)) and not (inputs(210));
    layer0_outputs(5860) <= (inputs(173)) and (inputs(216));
    layer0_outputs(5861) <= not(inputs(91)) or (inputs(80));
    layer0_outputs(5862) <= (inputs(168)) and not (inputs(146));
    layer0_outputs(5863) <= not(inputs(145));
    layer0_outputs(5864) <= not(inputs(46)) or (inputs(109));
    layer0_outputs(5865) <= (inputs(84)) and not (inputs(192));
    layer0_outputs(5866) <= (inputs(7)) or (inputs(40));
    layer0_outputs(5867) <= not((inputs(106)) and (inputs(90)));
    layer0_outputs(5868) <= not(inputs(68)) or (inputs(41));
    layer0_outputs(5869) <= not(inputs(232));
    layer0_outputs(5870) <= (inputs(22)) xor (inputs(69));
    layer0_outputs(5871) <= inputs(148);
    layer0_outputs(5872) <= not(inputs(114));
    layer0_outputs(5873) <= inputs(45);
    layer0_outputs(5874) <= not(inputs(24)) or (inputs(163));
    layer0_outputs(5875) <= inputs(142);
    layer0_outputs(5876) <= not(inputs(251));
    layer0_outputs(5877) <= (inputs(90)) and not (inputs(245));
    layer0_outputs(5878) <= (inputs(245)) and not (inputs(224));
    layer0_outputs(5879) <= not((inputs(254)) xor (inputs(125)));
    layer0_outputs(5880) <= inputs(196);
    layer0_outputs(5881) <= not(inputs(168)) or (inputs(47));
    layer0_outputs(5882) <= not(inputs(104));
    layer0_outputs(5883) <= not((inputs(151)) xor (inputs(253)));
    layer0_outputs(5884) <= (inputs(186)) or (inputs(201));
    layer0_outputs(5885) <= '1';
    layer0_outputs(5886) <= (inputs(25)) xor (inputs(44));
    layer0_outputs(5887) <= not(inputs(98));
    layer0_outputs(5888) <= not(inputs(75));
    layer0_outputs(5889) <= (inputs(207)) xor (inputs(106));
    layer0_outputs(5890) <= inputs(142);
    layer0_outputs(5891) <= not(inputs(202)) or (inputs(43));
    layer0_outputs(5892) <= not(inputs(232));
    layer0_outputs(5893) <= (inputs(19)) or (inputs(2));
    layer0_outputs(5894) <= not((inputs(28)) or (inputs(14)));
    layer0_outputs(5895) <= '0';
    layer0_outputs(5896) <= (inputs(165)) and not (inputs(66));
    layer0_outputs(5897) <= not(inputs(51)) or (inputs(252));
    layer0_outputs(5898) <= not(inputs(24)) or (inputs(192));
    layer0_outputs(5899) <= not(inputs(71)) or (inputs(45));
    layer0_outputs(5900) <= not((inputs(164)) or (inputs(219)));
    layer0_outputs(5901) <= (inputs(27)) xor (inputs(57));
    layer0_outputs(5902) <= '1';
    layer0_outputs(5903) <= inputs(101);
    layer0_outputs(5904) <= inputs(90);
    layer0_outputs(5905) <= (inputs(90)) and not (inputs(187));
    layer0_outputs(5906) <= (inputs(101)) and not (inputs(73));
    layer0_outputs(5907) <= not((inputs(218)) or (inputs(230)));
    layer0_outputs(5908) <= not(inputs(162));
    layer0_outputs(5909) <= not(inputs(213));
    layer0_outputs(5910) <= (inputs(188)) and (inputs(177));
    layer0_outputs(5911) <= (inputs(254)) or (inputs(54));
    layer0_outputs(5912) <= not(inputs(230)) or (inputs(89));
    layer0_outputs(5913) <= (inputs(100)) and not (inputs(80));
    layer0_outputs(5914) <= (inputs(172)) xor (inputs(97));
    layer0_outputs(5915) <= (inputs(57)) and (inputs(221));
    layer0_outputs(5916) <= (inputs(172)) xor (inputs(234));
    layer0_outputs(5917) <= inputs(103);
    layer0_outputs(5918) <= not((inputs(16)) or (inputs(9)));
    layer0_outputs(5919) <= (inputs(197)) and (inputs(156));
    layer0_outputs(5920) <= inputs(94);
    layer0_outputs(5921) <= inputs(195);
    layer0_outputs(5922) <= not(inputs(117));
    layer0_outputs(5923) <= not(inputs(5));
    layer0_outputs(5924) <= (inputs(230)) and not (inputs(107));
    layer0_outputs(5925) <= inputs(55);
    layer0_outputs(5926) <= not(inputs(80));
    layer0_outputs(5927) <= not((inputs(119)) or (inputs(13)));
    layer0_outputs(5928) <= (inputs(52)) and not (inputs(120));
    layer0_outputs(5929) <= (inputs(253)) xor (inputs(75));
    layer0_outputs(5930) <= (inputs(91)) and (inputs(25));
    layer0_outputs(5931) <= not(inputs(142)) or (inputs(220));
    layer0_outputs(5932) <= (inputs(152)) and not (inputs(27));
    layer0_outputs(5933) <= not((inputs(222)) or (inputs(138)));
    layer0_outputs(5934) <= not(inputs(26)) or (inputs(250));
    layer0_outputs(5935) <= not(inputs(68)) or (inputs(222));
    layer0_outputs(5936) <= not(inputs(186));
    layer0_outputs(5937) <= not(inputs(112));
    layer0_outputs(5938) <= (inputs(174)) and (inputs(60));
    layer0_outputs(5939) <= (inputs(158)) or (inputs(244));
    layer0_outputs(5940) <= (inputs(117)) and (inputs(168));
    layer0_outputs(5941) <= inputs(157);
    layer0_outputs(5942) <= not(inputs(121));
    layer0_outputs(5943) <= inputs(223);
    layer0_outputs(5944) <= inputs(153);
    layer0_outputs(5945) <= not((inputs(54)) xor (inputs(52)));
    layer0_outputs(5946) <= not((inputs(189)) or (inputs(32)));
    layer0_outputs(5947) <= not(inputs(110)) or (inputs(123));
    layer0_outputs(5948) <= not(inputs(60)) or (inputs(204));
    layer0_outputs(5949) <= inputs(124);
    layer0_outputs(5950) <= not((inputs(57)) or (inputs(220)));
    layer0_outputs(5951) <= not(inputs(198)) or (inputs(121));
    layer0_outputs(5952) <= (inputs(157)) or (inputs(153));
    layer0_outputs(5953) <= (inputs(172)) and not (inputs(65));
    layer0_outputs(5954) <= not(inputs(240)) or (inputs(27));
    layer0_outputs(5955) <= not((inputs(236)) or (inputs(178)));
    layer0_outputs(5956) <= not(inputs(23));
    layer0_outputs(5957) <= not((inputs(221)) or (inputs(174)));
    layer0_outputs(5958) <= not(inputs(223)) or (inputs(107));
    layer0_outputs(5959) <= not(inputs(78));
    layer0_outputs(5960) <= not(inputs(55));
    layer0_outputs(5961) <= not((inputs(171)) xor (inputs(125)));
    layer0_outputs(5962) <= (inputs(122)) and not (inputs(36));
    layer0_outputs(5963) <= not((inputs(99)) or (inputs(237)));
    layer0_outputs(5964) <= not(inputs(8));
    layer0_outputs(5965) <= not(inputs(248)) or (inputs(26));
    layer0_outputs(5966) <= not(inputs(239));
    layer0_outputs(5967) <= not(inputs(250));
    layer0_outputs(5968) <= (inputs(237)) and (inputs(158));
    layer0_outputs(5969) <= (inputs(130)) and not (inputs(224));
    layer0_outputs(5970) <= (inputs(25)) and (inputs(133));
    layer0_outputs(5971) <= not((inputs(37)) or (inputs(189)));
    layer0_outputs(5972) <= (inputs(7)) and not (inputs(15));
    layer0_outputs(5973) <= inputs(166);
    layer0_outputs(5974) <= not((inputs(59)) or (inputs(111)));
    layer0_outputs(5975) <= inputs(151);
    layer0_outputs(5976) <= not((inputs(64)) or (inputs(133)));
    layer0_outputs(5977) <= (inputs(21)) and not (inputs(251));
    layer0_outputs(5978) <= (inputs(94)) or (inputs(136));
    layer0_outputs(5979) <= inputs(244);
    layer0_outputs(5980) <= inputs(56);
    layer0_outputs(5981) <= (inputs(23)) and not (inputs(19));
    layer0_outputs(5982) <= not(inputs(27));
    layer0_outputs(5983) <= not((inputs(60)) or (inputs(35)));
    layer0_outputs(5984) <= inputs(42);
    layer0_outputs(5985) <= not(inputs(80));
    layer0_outputs(5986) <= (inputs(154)) and not (inputs(33));
    layer0_outputs(5987) <= not((inputs(4)) or (inputs(235)));
    layer0_outputs(5988) <= not(inputs(73));
    layer0_outputs(5989) <= (inputs(216)) or (inputs(36));
    layer0_outputs(5990) <= not(inputs(227));
    layer0_outputs(5991) <= (inputs(169)) and not (inputs(79));
    layer0_outputs(5992) <= inputs(124);
    layer0_outputs(5993) <= not(inputs(129));
    layer0_outputs(5994) <= (inputs(171)) and not (inputs(14));
    layer0_outputs(5995) <= (inputs(184)) xor (inputs(26));
    layer0_outputs(5996) <= (inputs(138)) and not (inputs(198));
    layer0_outputs(5997) <= not((inputs(219)) or (inputs(210)));
    layer0_outputs(5998) <= inputs(92);
    layer0_outputs(5999) <= (inputs(19)) or (inputs(147));
    layer0_outputs(6000) <= not((inputs(123)) and (inputs(203)));
    layer0_outputs(6001) <= not(inputs(124)) or (inputs(78));
    layer0_outputs(6002) <= not((inputs(200)) xor (inputs(100)));
    layer0_outputs(6003) <= (inputs(114)) or (inputs(117));
    layer0_outputs(6004) <= inputs(145);
    layer0_outputs(6005) <= not(inputs(131));
    layer0_outputs(6006) <= not(inputs(245));
    layer0_outputs(6007) <= (inputs(75)) and not (inputs(238));
    layer0_outputs(6008) <= (inputs(189)) or (inputs(126));
    layer0_outputs(6009) <= (inputs(53)) or (inputs(26));
    layer0_outputs(6010) <= not(inputs(25));
    layer0_outputs(6011) <= not(inputs(116)) or (inputs(173));
    layer0_outputs(6012) <= (inputs(131)) and not (inputs(16));
    layer0_outputs(6013) <= not(inputs(57));
    layer0_outputs(6014) <= (inputs(37)) or (inputs(78));
    layer0_outputs(6015) <= not(inputs(99));
    layer0_outputs(6016) <= inputs(238);
    layer0_outputs(6017) <= not((inputs(165)) or (inputs(24)));
    layer0_outputs(6018) <= not(inputs(14));
    layer0_outputs(6019) <= not(inputs(50)) or (inputs(144));
    layer0_outputs(6020) <= not(inputs(172));
    layer0_outputs(6021) <= not(inputs(76)) or (inputs(38));
    layer0_outputs(6022) <= (inputs(247)) or (inputs(201));
    layer0_outputs(6023) <= (inputs(27)) xor (inputs(215));
    layer0_outputs(6024) <= inputs(95);
    layer0_outputs(6025) <= not(inputs(69));
    layer0_outputs(6026) <= '0';
    layer0_outputs(6027) <= (inputs(76)) and (inputs(215));
    layer0_outputs(6028) <= (inputs(120)) and not (inputs(173));
    layer0_outputs(6029) <= not(inputs(88)) or (inputs(192));
    layer0_outputs(6030) <= not(inputs(138)) or (inputs(217));
    layer0_outputs(6031) <= not((inputs(41)) or (inputs(190)));
    layer0_outputs(6032) <= (inputs(239)) or (inputs(122));
    layer0_outputs(6033) <= (inputs(156)) xor (inputs(32));
    layer0_outputs(6034) <= (inputs(125)) and not (inputs(225));
    layer0_outputs(6035) <= not((inputs(217)) or (inputs(209)));
    layer0_outputs(6036) <= (inputs(242)) or (inputs(152));
    layer0_outputs(6037) <= not(inputs(79));
    layer0_outputs(6038) <= not((inputs(149)) xor (inputs(119)));
    layer0_outputs(6039) <= inputs(82);
    layer0_outputs(6040) <= (inputs(39)) or (inputs(223));
    layer0_outputs(6041) <= not(inputs(190));
    layer0_outputs(6042) <= (inputs(115)) xor (inputs(96));
    layer0_outputs(6043) <= not(inputs(6)) or (inputs(81));
    layer0_outputs(6044) <= (inputs(20)) or (inputs(125));
    layer0_outputs(6045) <= (inputs(56)) and not (inputs(227));
    layer0_outputs(6046) <= (inputs(129)) and not (inputs(190));
    layer0_outputs(6047) <= (inputs(67)) or (inputs(116));
    layer0_outputs(6048) <= not((inputs(104)) and (inputs(27)));
    layer0_outputs(6049) <= '0';
    layer0_outputs(6050) <= inputs(34);
    layer0_outputs(6051) <= inputs(87);
    layer0_outputs(6052) <= inputs(223);
    layer0_outputs(6053) <= (inputs(123)) and not (inputs(150));
    layer0_outputs(6054) <= not(inputs(90));
    layer0_outputs(6055) <= inputs(60);
    layer0_outputs(6056) <= (inputs(91)) and not (inputs(160));
    layer0_outputs(6057) <= not((inputs(186)) xor (inputs(145)));
    layer0_outputs(6058) <= not((inputs(47)) or (inputs(13)));
    layer0_outputs(6059) <= '1';
    layer0_outputs(6060) <= not((inputs(237)) or (inputs(127)));
    layer0_outputs(6061) <= not((inputs(51)) or (inputs(184)));
    layer0_outputs(6062) <= (inputs(22)) and not (inputs(147));
    layer0_outputs(6063) <= not((inputs(185)) xor (inputs(218)));
    layer0_outputs(6064) <= not((inputs(61)) or (inputs(211)));
    layer0_outputs(6065) <= not((inputs(78)) xor (inputs(175)));
    layer0_outputs(6066) <= not(inputs(222));
    layer0_outputs(6067) <= not(inputs(245));
    layer0_outputs(6068) <= not(inputs(219));
    layer0_outputs(6069) <= (inputs(125)) xor (inputs(104));
    layer0_outputs(6070) <= inputs(153);
    layer0_outputs(6071) <= (inputs(78)) or (inputs(93));
    layer0_outputs(6072) <= (inputs(139)) and (inputs(125));
    layer0_outputs(6073) <= not((inputs(233)) or (inputs(87)));
    layer0_outputs(6074) <= (inputs(40)) and not (inputs(22));
    layer0_outputs(6075) <= not(inputs(7));
    layer0_outputs(6076) <= (inputs(191)) or (inputs(145));
    layer0_outputs(6077) <= inputs(84);
    layer0_outputs(6078) <= (inputs(234)) and not (inputs(112));
    layer0_outputs(6079) <= not(inputs(108));
    layer0_outputs(6080) <= (inputs(90)) or (inputs(107));
    layer0_outputs(6081) <= (inputs(10)) xor (inputs(19));
    layer0_outputs(6082) <= (inputs(29)) or (inputs(188));
    layer0_outputs(6083) <= not(inputs(120));
    layer0_outputs(6084) <= not(inputs(176));
    layer0_outputs(6085) <= not((inputs(81)) and (inputs(112)));
    layer0_outputs(6086) <= (inputs(230)) xor (inputs(4));
    layer0_outputs(6087) <= (inputs(240)) xor (inputs(240));
    layer0_outputs(6088) <= not(inputs(148));
    layer0_outputs(6089) <= not((inputs(139)) and (inputs(200)));
    layer0_outputs(6090) <= not(inputs(6)) or (inputs(62));
    layer0_outputs(6091) <= not((inputs(222)) or (inputs(153)));
    layer0_outputs(6092) <= not((inputs(101)) or (inputs(222)));
    layer0_outputs(6093) <= not(inputs(183));
    layer0_outputs(6094) <= not(inputs(208)) or (inputs(156));
    layer0_outputs(6095) <= '0';
    layer0_outputs(6096) <= not((inputs(209)) or (inputs(226)));
    layer0_outputs(6097) <= not((inputs(49)) and (inputs(188)));
    layer0_outputs(6098) <= not(inputs(71)) or (inputs(140));
    layer0_outputs(6099) <= inputs(82);
    layer0_outputs(6100) <= not((inputs(48)) xor (inputs(1)));
    layer0_outputs(6101) <= not(inputs(86));
    layer0_outputs(6102) <= not(inputs(139)) or (inputs(6));
    layer0_outputs(6103) <= not(inputs(150)) or (inputs(57));
    layer0_outputs(6104) <= not(inputs(93)) or (inputs(130));
    layer0_outputs(6105) <= not(inputs(226));
    layer0_outputs(6106) <= not((inputs(91)) or (inputs(190)));
    layer0_outputs(6107) <= (inputs(131)) xor (inputs(80));
    layer0_outputs(6108) <= not((inputs(22)) xor (inputs(174)));
    layer0_outputs(6109) <= not(inputs(91));
    layer0_outputs(6110) <= (inputs(142)) and not (inputs(239));
    layer0_outputs(6111) <= (inputs(254)) xor (inputs(10));
    layer0_outputs(6112) <= not(inputs(201));
    layer0_outputs(6113) <= (inputs(121)) or (inputs(97));
    layer0_outputs(6114) <= not((inputs(27)) xor (inputs(22)));
    layer0_outputs(6115) <= inputs(19);
    layer0_outputs(6116) <= (inputs(137)) or (inputs(122));
    layer0_outputs(6117) <= not(inputs(229));
    layer0_outputs(6118) <= inputs(120);
    layer0_outputs(6119) <= not((inputs(103)) or (inputs(181)));
    layer0_outputs(6120) <= not(inputs(103));
    layer0_outputs(6121) <= not(inputs(199));
    layer0_outputs(6122) <= '1';
    layer0_outputs(6123) <= (inputs(240)) or (inputs(1));
    layer0_outputs(6124) <= (inputs(163)) and not (inputs(174));
    layer0_outputs(6125) <= not((inputs(156)) xor (inputs(103)));
    layer0_outputs(6126) <= inputs(189);
    layer0_outputs(6127) <= inputs(90);
    layer0_outputs(6128) <= (inputs(32)) xor (inputs(255));
    layer0_outputs(6129) <= not((inputs(80)) or (inputs(46)));
    layer0_outputs(6130) <= inputs(26);
    layer0_outputs(6131) <= inputs(68);
    layer0_outputs(6132) <= inputs(135);
    layer0_outputs(6133) <= '1';
    layer0_outputs(6134) <= (inputs(52)) or (inputs(98));
    layer0_outputs(6135) <= (inputs(32)) or (inputs(149));
    layer0_outputs(6136) <= not(inputs(87));
    layer0_outputs(6137) <= (inputs(213)) and not (inputs(17));
    layer0_outputs(6138) <= not(inputs(105));
    layer0_outputs(6139) <= inputs(103);
    layer0_outputs(6140) <= not((inputs(141)) or (inputs(169)));
    layer0_outputs(6141) <= not(inputs(21)) or (inputs(5));
    layer0_outputs(6142) <= not((inputs(174)) xor (inputs(85)));
    layer0_outputs(6143) <= inputs(101);
    layer0_outputs(6144) <= not((inputs(43)) xor (inputs(55)));
    layer0_outputs(6145) <= (inputs(4)) or (inputs(13));
    layer0_outputs(6146) <= (inputs(69)) or (inputs(68));
    layer0_outputs(6147) <= (inputs(195)) or (inputs(220));
    layer0_outputs(6148) <= not(inputs(135)) or (inputs(208));
    layer0_outputs(6149) <= not((inputs(203)) xor (inputs(195)));
    layer0_outputs(6150) <= (inputs(13)) or (inputs(224));
    layer0_outputs(6151) <= not((inputs(235)) or (inputs(254)));
    layer0_outputs(6152) <= (inputs(69)) and not (inputs(51));
    layer0_outputs(6153) <= not(inputs(195));
    layer0_outputs(6154) <= not((inputs(230)) xor (inputs(160)));
    layer0_outputs(6155) <= (inputs(200)) and (inputs(172));
    layer0_outputs(6156) <= not(inputs(246));
    layer0_outputs(6157) <= inputs(229);
    layer0_outputs(6158) <= (inputs(134)) or (inputs(239));
    layer0_outputs(6159) <= not(inputs(189));
    layer0_outputs(6160) <= not(inputs(70));
    layer0_outputs(6161) <= not((inputs(185)) xor (inputs(201)));
    layer0_outputs(6162) <= not(inputs(183));
    layer0_outputs(6163) <= inputs(41);
    layer0_outputs(6164) <= (inputs(148)) and not (inputs(221));
    layer0_outputs(6165) <= (inputs(43)) and not (inputs(222));
    layer0_outputs(6166) <= not((inputs(222)) and (inputs(236)));
    layer0_outputs(6167) <= not(inputs(134));
    layer0_outputs(6168) <= (inputs(172)) and not (inputs(110));
    layer0_outputs(6169) <= not(inputs(215)) or (inputs(93));
    layer0_outputs(6170) <= (inputs(82)) xor (inputs(133));
    layer0_outputs(6171) <= not(inputs(197)) or (inputs(215));
    layer0_outputs(6172) <= (inputs(165)) and not (inputs(242));
    layer0_outputs(6173) <= (inputs(228)) and not (inputs(15));
    layer0_outputs(6174) <= (inputs(5)) xor (inputs(53));
    layer0_outputs(6175) <= not((inputs(176)) or (inputs(169)));
    layer0_outputs(6176) <= not(inputs(188)) or (inputs(250));
    layer0_outputs(6177) <= inputs(249);
    layer0_outputs(6178) <= (inputs(132)) or (inputs(248));
    layer0_outputs(6179) <= inputs(69);
    layer0_outputs(6180) <= (inputs(244)) or (inputs(242));
    layer0_outputs(6181) <= (inputs(95)) or (inputs(213));
    layer0_outputs(6182) <= (inputs(16)) or (inputs(154));
    layer0_outputs(6183) <= not(inputs(161)) or (inputs(15));
    layer0_outputs(6184) <= (inputs(100)) or (inputs(10));
    layer0_outputs(6185) <= (inputs(246)) xor (inputs(182));
    layer0_outputs(6186) <= not(inputs(203)) or (inputs(236));
    layer0_outputs(6187) <= inputs(176);
    layer0_outputs(6188) <= not((inputs(127)) or (inputs(170)));
    layer0_outputs(6189) <= (inputs(208)) or (inputs(166));
    layer0_outputs(6190) <= not((inputs(23)) or (inputs(63)));
    layer0_outputs(6191) <= not(inputs(119)) or (inputs(163));
    layer0_outputs(6192) <= not(inputs(239));
    layer0_outputs(6193) <= not(inputs(148));
    layer0_outputs(6194) <= (inputs(154)) xor (inputs(231));
    layer0_outputs(6195) <= (inputs(55)) or (inputs(245));
    layer0_outputs(6196) <= (inputs(106)) and not (inputs(15));
    layer0_outputs(6197) <= not((inputs(138)) xor (inputs(109)));
    layer0_outputs(6198) <= not(inputs(68));
    layer0_outputs(6199) <= not(inputs(126));
    layer0_outputs(6200) <= not(inputs(10));
    layer0_outputs(6201) <= (inputs(75)) and (inputs(36));
    layer0_outputs(6202) <= inputs(178);
    layer0_outputs(6203) <= not((inputs(6)) xor (inputs(225)));
    layer0_outputs(6204) <= (inputs(10)) xor (inputs(138));
    layer0_outputs(6205) <= (inputs(223)) or (inputs(7));
    layer0_outputs(6206) <= (inputs(65)) and (inputs(45));
    layer0_outputs(6207) <= not(inputs(155));
    layer0_outputs(6208) <= not(inputs(225)) or (inputs(237));
    layer0_outputs(6209) <= not(inputs(40)) or (inputs(190));
    layer0_outputs(6210) <= (inputs(30)) and not (inputs(175));
    layer0_outputs(6211) <= inputs(39);
    layer0_outputs(6212) <= not(inputs(174)) or (inputs(13));
    layer0_outputs(6213) <= not(inputs(35));
    layer0_outputs(6214) <= (inputs(158)) or (inputs(32));
    layer0_outputs(6215) <= not((inputs(89)) xor (inputs(168)));
    layer0_outputs(6216) <= (inputs(175)) xor (inputs(46));
    layer0_outputs(6217) <= not((inputs(161)) xor (inputs(164)));
    layer0_outputs(6218) <= (inputs(80)) or (inputs(92));
    layer0_outputs(6219) <= not((inputs(37)) or (inputs(94)));
    layer0_outputs(6220) <= not(inputs(167));
    layer0_outputs(6221) <= not((inputs(194)) and (inputs(18)));
    layer0_outputs(6222) <= '1';
    layer0_outputs(6223) <= (inputs(219)) and not (inputs(130));
    layer0_outputs(6224) <= not((inputs(157)) and (inputs(143)));
    layer0_outputs(6225) <= not((inputs(88)) xor (inputs(146)));
    layer0_outputs(6226) <= not(inputs(230)) or (inputs(77));
    layer0_outputs(6227) <= (inputs(71)) and (inputs(103));
    layer0_outputs(6228) <= not(inputs(131));
    layer0_outputs(6229) <= (inputs(197)) xor (inputs(50));
    layer0_outputs(6230) <= not((inputs(122)) xor (inputs(61)));
    layer0_outputs(6231) <= not(inputs(23)) or (inputs(179));
    layer0_outputs(6232) <= not(inputs(3));
    layer0_outputs(6233) <= (inputs(255)) or (inputs(248));
    layer0_outputs(6234) <= inputs(192);
    layer0_outputs(6235) <= not(inputs(247));
    layer0_outputs(6236) <= not(inputs(119));
    layer0_outputs(6237) <= not((inputs(54)) xor (inputs(38)));
    layer0_outputs(6238) <= not(inputs(166));
    layer0_outputs(6239) <= not((inputs(14)) or (inputs(254)));
    layer0_outputs(6240) <= not(inputs(24));
    layer0_outputs(6241) <= not((inputs(222)) or (inputs(72)));
    layer0_outputs(6242) <= not((inputs(207)) or (inputs(161)));
    layer0_outputs(6243) <= not((inputs(28)) or (inputs(123)));
    layer0_outputs(6244) <= (inputs(249)) xor (inputs(86));
    layer0_outputs(6245) <= (inputs(68)) or (inputs(32));
    layer0_outputs(6246) <= not(inputs(92));
    layer0_outputs(6247) <= inputs(254);
    layer0_outputs(6248) <= not(inputs(125)) or (inputs(222));
    layer0_outputs(6249) <= not(inputs(111));
    layer0_outputs(6250) <= (inputs(229)) and not (inputs(42));
    layer0_outputs(6251) <= not(inputs(9)) or (inputs(129));
    layer0_outputs(6252) <= inputs(39);
    layer0_outputs(6253) <= not((inputs(198)) or (inputs(64)));
    layer0_outputs(6254) <= inputs(113);
    layer0_outputs(6255) <= (inputs(119)) and not (inputs(126));
    layer0_outputs(6256) <= not(inputs(3));
    layer0_outputs(6257) <= not(inputs(61)) or (inputs(129));
    layer0_outputs(6258) <= not(inputs(227));
    layer0_outputs(6259) <= not(inputs(0)) or (inputs(4));
    layer0_outputs(6260) <= (inputs(61)) or (inputs(239));
    layer0_outputs(6261) <= (inputs(193)) or (inputs(246));
    layer0_outputs(6262) <= not(inputs(172));
    layer0_outputs(6263) <= (inputs(203)) and not (inputs(1));
    layer0_outputs(6264) <= inputs(104);
    layer0_outputs(6265) <= not((inputs(67)) or (inputs(5)));
    layer0_outputs(6266) <= (inputs(143)) or (inputs(77));
    layer0_outputs(6267) <= inputs(121);
    layer0_outputs(6268) <= '0';
    layer0_outputs(6269) <= inputs(183);
    layer0_outputs(6270) <= not(inputs(9));
    layer0_outputs(6271) <= not((inputs(44)) xor (inputs(209)));
    layer0_outputs(6272) <= (inputs(92)) xor (inputs(19));
    layer0_outputs(6273) <= inputs(55);
    layer0_outputs(6274) <= not(inputs(155));
    layer0_outputs(6275) <= inputs(141);
    layer0_outputs(6276) <= not(inputs(250));
    layer0_outputs(6277) <= not((inputs(221)) or (inputs(20)));
    layer0_outputs(6278) <= not(inputs(150)) or (inputs(208));
    layer0_outputs(6279) <= inputs(100);
    layer0_outputs(6280) <= not(inputs(184)) or (inputs(245));
    layer0_outputs(6281) <= (inputs(17)) and (inputs(126));
    layer0_outputs(6282) <= not(inputs(226));
    layer0_outputs(6283) <= (inputs(9)) or (inputs(160));
    layer0_outputs(6284) <= not(inputs(77)) or (inputs(80));
    layer0_outputs(6285) <= not(inputs(153)) or (inputs(174));
    layer0_outputs(6286) <= not(inputs(184)) or (inputs(131));
    layer0_outputs(6287) <= (inputs(184)) xor (inputs(176));
    layer0_outputs(6288) <= not((inputs(70)) and (inputs(73)));
    layer0_outputs(6289) <= inputs(230);
    layer0_outputs(6290) <= not(inputs(153));
    layer0_outputs(6291) <= not(inputs(40));
    layer0_outputs(6292) <= not(inputs(216));
    layer0_outputs(6293) <= inputs(1);
    layer0_outputs(6294) <= (inputs(188)) or (inputs(216));
    layer0_outputs(6295) <= (inputs(129)) and not (inputs(10));
    layer0_outputs(6296) <= not((inputs(72)) or (inputs(93)));
    layer0_outputs(6297) <= inputs(2);
    layer0_outputs(6298) <= not((inputs(79)) xor (inputs(37)));
    layer0_outputs(6299) <= (inputs(212)) and (inputs(200));
    layer0_outputs(6300) <= not((inputs(49)) xor (inputs(228)));
    layer0_outputs(6301) <= (inputs(253)) and not (inputs(95));
    layer0_outputs(6302) <= not((inputs(206)) xor (inputs(87)));
    layer0_outputs(6303) <= '0';
    layer0_outputs(6304) <= not(inputs(39));
    layer0_outputs(6305) <= (inputs(149)) and not (inputs(33));
    layer0_outputs(6306) <= not(inputs(41));
    layer0_outputs(6307) <= inputs(109);
    layer0_outputs(6308) <= inputs(202);
    layer0_outputs(6309) <= not((inputs(21)) or (inputs(87)));
    layer0_outputs(6310) <= not((inputs(171)) xor (inputs(205)));
    layer0_outputs(6311) <= not((inputs(148)) and (inputs(26)));
    layer0_outputs(6312) <= (inputs(136)) xor (inputs(21));
    layer0_outputs(6313) <= (inputs(63)) or (inputs(55));
    layer0_outputs(6314) <= not((inputs(101)) or (inputs(180)));
    layer0_outputs(6315) <= not(inputs(18)) or (inputs(63));
    layer0_outputs(6316) <= (inputs(160)) or (inputs(66));
    layer0_outputs(6317) <= not((inputs(173)) xor (inputs(69)));
    layer0_outputs(6318) <= inputs(25);
    layer0_outputs(6319) <= not((inputs(92)) or (inputs(93)));
    layer0_outputs(6320) <= (inputs(169)) or (inputs(64));
    layer0_outputs(6321) <= not((inputs(163)) or (inputs(148)));
    layer0_outputs(6322) <= not((inputs(4)) xor (inputs(148)));
    layer0_outputs(6323) <= not(inputs(92)) or (inputs(241));
    layer0_outputs(6324) <= inputs(89);
    layer0_outputs(6325) <= (inputs(51)) xor (inputs(52));
    layer0_outputs(6326) <= not((inputs(171)) and (inputs(198)));
    layer0_outputs(6327) <= '1';
    layer0_outputs(6328) <= inputs(157);
    layer0_outputs(6329) <= (inputs(207)) and not (inputs(128));
    layer0_outputs(6330) <= not(inputs(100));
    layer0_outputs(6331) <= (inputs(52)) and not (inputs(175));
    layer0_outputs(6332) <= not(inputs(177)) or (inputs(14));
    layer0_outputs(6333) <= not((inputs(103)) xor (inputs(97)));
    layer0_outputs(6334) <= not((inputs(17)) or (inputs(90)));
    layer0_outputs(6335) <= not(inputs(24)) or (inputs(241));
    layer0_outputs(6336) <= not(inputs(152));
    layer0_outputs(6337) <= (inputs(85)) and not (inputs(27));
    layer0_outputs(6338) <= (inputs(58)) or (inputs(183));
    layer0_outputs(6339) <= not((inputs(10)) or (inputs(127)));
    layer0_outputs(6340) <= not((inputs(35)) or (inputs(13)));
    layer0_outputs(6341) <= not(inputs(85)) or (inputs(160));
    layer0_outputs(6342) <= (inputs(32)) and not (inputs(25));
    layer0_outputs(6343) <= (inputs(28)) xor (inputs(138));
    layer0_outputs(6344) <= (inputs(137)) and not (inputs(96));
    layer0_outputs(6345) <= (inputs(81)) or (inputs(89));
    layer0_outputs(6346) <= inputs(123);
    layer0_outputs(6347) <= not(inputs(190));
    layer0_outputs(6348) <= not((inputs(88)) xor (inputs(56)));
    layer0_outputs(6349) <= not(inputs(182));
    layer0_outputs(6350) <= (inputs(184)) and (inputs(232));
    layer0_outputs(6351) <= not(inputs(170));
    layer0_outputs(6352) <= not(inputs(42));
    layer0_outputs(6353) <= not((inputs(80)) or (inputs(104)));
    layer0_outputs(6354) <= not(inputs(235)) or (inputs(15));
    layer0_outputs(6355) <= inputs(76);
    layer0_outputs(6356) <= (inputs(226)) xor (inputs(65));
    layer0_outputs(6357) <= (inputs(38)) xor (inputs(207));
    layer0_outputs(6358) <= not(inputs(108)) or (inputs(66));
    layer0_outputs(6359) <= not((inputs(127)) or (inputs(131)));
    layer0_outputs(6360) <= inputs(248);
    layer0_outputs(6361) <= not((inputs(179)) or (inputs(208)));
    layer0_outputs(6362) <= not(inputs(126)) or (inputs(130));
    layer0_outputs(6363) <= (inputs(172)) and not (inputs(113));
    layer0_outputs(6364) <= inputs(121);
    layer0_outputs(6365) <= not(inputs(212)) or (inputs(238));
    layer0_outputs(6366) <= not(inputs(114));
    layer0_outputs(6367) <= not((inputs(76)) or (inputs(44)));
    layer0_outputs(6368) <= not(inputs(82));
    layer0_outputs(6369) <= inputs(193);
    layer0_outputs(6370) <= inputs(107);
    layer0_outputs(6371) <= not(inputs(251));
    layer0_outputs(6372) <= (inputs(172)) and not (inputs(6));
    layer0_outputs(6373) <= inputs(124);
    layer0_outputs(6374) <= not(inputs(249));
    layer0_outputs(6375) <= inputs(164);
    layer0_outputs(6376) <= not((inputs(187)) xor (inputs(105)));
    layer0_outputs(6377) <= not((inputs(179)) xor (inputs(177)));
    layer0_outputs(6378) <= not((inputs(216)) xor (inputs(248)));
    layer0_outputs(6379) <= (inputs(121)) and not (inputs(97));
    layer0_outputs(6380) <= (inputs(133)) and not (inputs(218));
    layer0_outputs(6381) <= not((inputs(16)) or (inputs(29)));
    layer0_outputs(6382) <= not((inputs(61)) xor (inputs(37)));
    layer0_outputs(6383) <= not(inputs(19)) or (inputs(208));
    layer0_outputs(6384) <= (inputs(155)) and not (inputs(253));
    layer0_outputs(6385) <= not(inputs(166));
    layer0_outputs(6386) <= not(inputs(100)) or (inputs(253));
    layer0_outputs(6387) <= (inputs(89)) or (inputs(220));
    layer0_outputs(6388) <= (inputs(173)) and not (inputs(100));
    layer0_outputs(6389) <= not((inputs(158)) xor (inputs(117)));
    layer0_outputs(6390) <= not((inputs(203)) xor (inputs(65)));
    layer0_outputs(6391) <= (inputs(231)) xor (inputs(27));
    layer0_outputs(6392) <= (inputs(207)) xor (inputs(149));
    layer0_outputs(6393) <= not((inputs(246)) and (inputs(195)));
    layer0_outputs(6394) <= not(inputs(231)) or (inputs(106));
    layer0_outputs(6395) <= not(inputs(75));
    layer0_outputs(6396) <= not(inputs(53)) or (inputs(243));
    layer0_outputs(6397) <= (inputs(48)) or (inputs(149));
    layer0_outputs(6398) <= not(inputs(56));
    layer0_outputs(6399) <= not(inputs(94));
    layer0_outputs(6400) <= not(inputs(110)) or (inputs(182));
    layer0_outputs(6401) <= not(inputs(40));
    layer0_outputs(6402) <= (inputs(77)) or (inputs(92));
    layer0_outputs(6403) <= not((inputs(55)) and (inputs(154)));
    layer0_outputs(6404) <= not(inputs(72));
    layer0_outputs(6405) <= (inputs(36)) xor (inputs(200));
    layer0_outputs(6406) <= (inputs(31)) or (inputs(45));
    layer0_outputs(6407) <= not(inputs(239));
    layer0_outputs(6408) <= inputs(72);
    layer0_outputs(6409) <= not((inputs(196)) and (inputs(201)));
    layer0_outputs(6410) <= inputs(100);
    layer0_outputs(6411) <= (inputs(179)) xor (inputs(222));
    layer0_outputs(6412) <= (inputs(130)) or (inputs(153));
    layer0_outputs(6413) <= not(inputs(39)) or (inputs(178));
    layer0_outputs(6414) <= not((inputs(133)) xor (inputs(131)));
    layer0_outputs(6415) <= not(inputs(59)) or (inputs(239));
    layer0_outputs(6416) <= (inputs(155)) xor (inputs(41));
    layer0_outputs(6417) <= (inputs(178)) and not (inputs(124));
    layer0_outputs(6418) <= not((inputs(5)) or (inputs(43)));
    layer0_outputs(6419) <= (inputs(171)) and not (inputs(132));
    layer0_outputs(6420) <= not(inputs(148)) or (inputs(178));
    layer0_outputs(6421) <= not((inputs(250)) or (inputs(229)));
    layer0_outputs(6422) <= inputs(8);
    layer0_outputs(6423) <= not((inputs(5)) xor (inputs(45)));
    layer0_outputs(6424) <= not(inputs(145));
    layer0_outputs(6425) <= inputs(76);
    layer0_outputs(6426) <= not(inputs(153)) or (inputs(62));
    layer0_outputs(6427) <= not(inputs(23)) or (inputs(190));
    layer0_outputs(6428) <= not(inputs(36)) or (inputs(187));
    layer0_outputs(6429) <= not((inputs(163)) xor (inputs(198)));
    layer0_outputs(6430) <= (inputs(36)) and not (inputs(234));
    layer0_outputs(6431) <= not((inputs(194)) or (inputs(11)));
    layer0_outputs(6432) <= not(inputs(222)) or (inputs(31));
    layer0_outputs(6433) <= (inputs(61)) xor (inputs(28));
    layer0_outputs(6434) <= not(inputs(137)) or (inputs(155));
    layer0_outputs(6435) <= (inputs(121)) or (inputs(35));
    layer0_outputs(6436) <= not(inputs(62));
    layer0_outputs(6437) <= (inputs(203)) and not (inputs(28));
    layer0_outputs(6438) <= not(inputs(180));
    layer0_outputs(6439) <= (inputs(109)) and not (inputs(12));
    layer0_outputs(6440) <= not(inputs(219));
    layer0_outputs(6441) <= (inputs(90)) and not (inputs(71));
    layer0_outputs(6442) <= not(inputs(246)) or (inputs(14));
    layer0_outputs(6443) <= inputs(250);
    layer0_outputs(6444) <= not(inputs(171)) or (inputs(223));
    layer0_outputs(6445) <= (inputs(64)) and not (inputs(131));
    layer0_outputs(6446) <= (inputs(42)) and (inputs(85));
    layer0_outputs(6447) <= not(inputs(139));
    layer0_outputs(6448) <= inputs(113);
    layer0_outputs(6449) <= not(inputs(140));
    layer0_outputs(6450) <= not((inputs(132)) xor (inputs(137)));
    layer0_outputs(6451) <= (inputs(178)) or (inputs(81));
    layer0_outputs(6452) <= not(inputs(182));
    layer0_outputs(6453) <= inputs(95);
    layer0_outputs(6454) <= not(inputs(118)) or (inputs(4));
    layer0_outputs(6455) <= not(inputs(31)) or (inputs(52));
    layer0_outputs(6456) <= inputs(59);
    layer0_outputs(6457) <= not(inputs(1));
    layer0_outputs(6458) <= (inputs(18)) or (inputs(56));
    layer0_outputs(6459) <= (inputs(254)) xor (inputs(207));
    layer0_outputs(6460) <= (inputs(182)) or (inputs(44));
    layer0_outputs(6461) <= (inputs(84)) xor (inputs(224));
    layer0_outputs(6462) <= (inputs(126)) or (inputs(18));
    layer0_outputs(6463) <= (inputs(223)) or (inputs(84));
    layer0_outputs(6464) <= (inputs(23)) or (inputs(36));
    layer0_outputs(6465) <= (inputs(214)) and (inputs(132));
    layer0_outputs(6466) <= (inputs(95)) xor (inputs(57));
    layer0_outputs(6467) <= (inputs(199)) and not (inputs(86));
    layer0_outputs(6468) <= (inputs(175)) and not (inputs(26));
    layer0_outputs(6469) <= (inputs(191)) or (inputs(8));
    layer0_outputs(6470) <= not((inputs(249)) xor (inputs(231)));
    layer0_outputs(6471) <= inputs(60);
    layer0_outputs(6472) <= (inputs(2)) xor (inputs(15));
    layer0_outputs(6473) <= (inputs(223)) or (inputs(62));
    layer0_outputs(6474) <= (inputs(230)) or (inputs(229));
    layer0_outputs(6475) <= inputs(41);
    layer0_outputs(6476) <= inputs(62);
    layer0_outputs(6477) <= (inputs(211)) or (inputs(143));
    layer0_outputs(6478) <= not((inputs(143)) xor (inputs(139)));
    layer0_outputs(6479) <= (inputs(152)) or (inputs(237));
    layer0_outputs(6480) <= not(inputs(166));
    layer0_outputs(6481) <= not((inputs(12)) or (inputs(94)));
    layer0_outputs(6482) <= inputs(44);
    layer0_outputs(6483) <= not((inputs(175)) xor (inputs(253)));
    layer0_outputs(6484) <= '0';
    layer0_outputs(6485) <= not(inputs(200)) or (inputs(239));
    layer0_outputs(6486) <= (inputs(78)) xor (inputs(179));
    layer0_outputs(6487) <= '1';
    layer0_outputs(6488) <= (inputs(71)) and not (inputs(138));
    layer0_outputs(6489) <= not(inputs(117));
    layer0_outputs(6490) <= inputs(114);
    layer0_outputs(6491) <= inputs(229);
    layer0_outputs(6492) <= not((inputs(238)) xor (inputs(47)));
    layer0_outputs(6493) <= not(inputs(162));
    layer0_outputs(6494) <= not(inputs(182));
    layer0_outputs(6495) <= not(inputs(5));
    layer0_outputs(6496) <= not(inputs(205));
    layer0_outputs(6497) <= not(inputs(65));
    layer0_outputs(6498) <= (inputs(53)) or (inputs(25));
    layer0_outputs(6499) <= not(inputs(97));
    layer0_outputs(6500) <= (inputs(165)) and not (inputs(240));
    layer0_outputs(6501) <= not((inputs(30)) or (inputs(190)));
    layer0_outputs(6502) <= (inputs(109)) or (inputs(131));
    layer0_outputs(6503) <= not(inputs(162));
    layer0_outputs(6504) <= '0';
    layer0_outputs(6505) <= not((inputs(189)) and (inputs(5)));
    layer0_outputs(6506) <= inputs(123);
    layer0_outputs(6507) <= (inputs(21)) or (inputs(33));
    layer0_outputs(6508) <= not(inputs(119));
    layer0_outputs(6509) <= inputs(36);
    layer0_outputs(6510) <= not(inputs(68));
    layer0_outputs(6511) <= (inputs(209)) and not (inputs(71));
    layer0_outputs(6512) <= not(inputs(130));
    layer0_outputs(6513) <= not(inputs(248));
    layer0_outputs(6514) <= not(inputs(143)) or (inputs(32));
    layer0_outputs(6515) <= (inputs(243)) and (inputs(219));
    layer0_outputs(6516) <= not(inputs(231));
    layer0_outputs(6517) <= inputs(197);
    layer0_outputs(6518) <= not(inputs(222)) or (inputs(15));
    layer0_outputs(6519) <= not(inputs(200));
    layer0_outputs(6520) <= not(inputs(149)) or (inputs(106));
    layer0_outputs(6521) <= (inputs(154)) or (inputs(81));
    layer0_outputs(6522) <= (inputs(170)) or (inputs(128));
    layer0_outputs(6523) <= not((inputs(72)) xor (inputs(15)));
    layer0_outputs(6524) <= (inputs(142)) or (inputs(11));
    layer0_outputs(6525) <= not(inputs(181));
    layer0_outputs(6526) <= not((inputs(204)) or (inputs(217)));
    layer0_outputs(6527) <= not((inputs(126)) xor (inputs(155)));
    layer0_outputs(6528) <= (inputs(212)) and (inputs(76));
    layer0_outputs(6529) <= not((inputs(191)) xor (inputs(110)));
    layer0_outputs(6530) <= (inputs(36)) and not (inputs(165));
    layer0_outputs(6531) <= not(inputs(56)) or (inputs(4));
    layer0_outputs(6532) <= inputs(123);
    layer0_outputs(6533) <= (inputs(179)) and (inputs(244));
    layer0_outputs(6534) <= (inputs(170)) or (inputs(175));
    layer0_outputs(6535) <= inputs(91);
    layer0_outputs(6536) <= (inputs(248)) or (inputs(125));
    layer0_outputs(6537) <= not((inputs(81)) and (inputs(134)));
    layer0_outputs(6538) <= inputs(157);
    layer0_outputs(6539) <= not(inputs(139)) or (inputs(42));
    layer0_outputs(6540) <= not(inputs(70));
    layer0_outputs(6541) <= not(inputs(209));
    layer0_outputs(6542) <= not(inputs(138)) or (inputs(214));
    layer0_outputs(6543) <= not(inputs(69));
    layer0_outputs(6544) <= '1';
    layer0_outputs(6545) <= not((inputs(85)) or (inputs(115)));
    layer0_outputs(6546) <= (inputs(133)) xor (inputs(98));
    layer0_outputs(6547) <= not(inputs(184));
    layer0_outputs(6548) <= not(inputs(89));
    layer0_outputs(6549) <= inputs(113);
    layer0_outputs(6550) <= not(inputs(211)) or (inputs(58));
    layer0_outputs(6551) <= not(inputs(242));
    layer0_outputs(6552) <= (inputs(40)) or (inputs(62));
    layer0_outputs(6553) <= (inputs(87)) xor (inputs(100));
    layer0_outputs(6554) <= (inputs(199)) or (inputs(134));
    layer0_outputs(6555) <= inputs(115);
    layer0_outputs(6556) <= (inputs(141)) or (inputs(188));
    layer0_outputs(6557) <= inputs(126);
    layer0_outputs(6558) <= not((inputs(2)) or (inputs(1)));
    layer0_outputs(6559) <= (inputs(211)) or (inputs(160));
    layer0_outputs(6560) <= not(inputs(178));
    layer0_outputs(6561) <= inputs(41);
    layer0_outputs(6562) <= (inputs(195)) and not (inputs(62));
    layer0_outputs(6563) <= not((inputs(244)) or (inputs(228)));
    layer0_outputs(6564) <= (inputs(87)) and not (inputs(185));
    layer0_outputs(6565) <= inputs(193);
    layer0_outputs(6566) <= (inputs(26)) and not (inputs(133));
    layer0_outputs(6567) <= not((inputs(91)) xor (inputs(142)));
    layer0_outputs(6568) <= (inputs(7)) and not (inputs(174));
    layer0_outputs(6569) <= inputs(173);
    layer0_outputs(6570) <= (inputs(171)) and not (inputs(53));
    layer0_outputs(6571) <= (inputs(22)) or (inputs(33));
    layer0_outputs(6572) <= inputs(134);
    layer0_outputs(6573) <= not((inputs(80)) or (inputs(99)));
    layer0_outputs(6574) <= not((inputs(195)) or (inputs(50)));
    layer0_outputs(6575) <= (inputs(105)) and not (inputs(192));
    layer0_outputs(6576) <= not(inputs(136));
    layer0_outputs(6577) <= (inputs(2)) or (inputs(231));
    layer0_outputs(6578) <= not(inputs(108));
    layer0_outputs(6579) <= (inputs(175)) or (inputs(212));
    layer0_outputs(6580) <= (inputs(121)) or (inputs(255));
    layer0_outputs(6581) <= not((inputs(210)) or (inputs(213)));
    layer0_outputs(6582) <= not(inputs(98));
    layer0_outputs(6583) <= not((inputs(19)) or (inputs(150)));
    layer0_outputs(6584) <= (inputs(75)) and (inputs(25));
    layer0_outputs(6585) <= not((inputs(119)) or (inputs(15)));
    layer0_outputs(6586) <= '0';
    layer0_outputs(6587) <= (inputs(166)) or (inputs(80));
    layer0_outputs(6588) <= (inputs(120)) or (inputs(14));
    layer0_outputs(6589) <= not(inputs(135));
    layer0_outputs(6590) <= not((inputs(156)) or (inputs(216)));
    layer0_outputs(6591) <= not(inputs(127)) or (inputs(190));
    layer0_outputs(6592) <= not((inputs(213)) or (inputs(223)));
    layer0_outputs(6593) <= (inputs(158)) xor (inputs(118));
    layer0_outputs(6594) <= (inputs(62)) xor (inputs(36));
    layer0_outputs(6595) <= inputs(29);
    layer0_outputs(6596) <= not((inputs(144)) xor (inputs(46)));
    layer0_outputs(6597) <= not(inputs(77));
    layer0_outputs(6598) <= inputs(191);
    layer0_outputs(6599) <= (inputs(177)) or (inputs(17));
    layer0_outputs(6600) <= inputs(91);
    layer0_outputs(6601) <= not((inputs(233)) or (inputs(44)));
    layer0_outputs(6602) <= not(inputs(245));
    layer0_outputs(6603) <= (inputs(221)) and not (inputs(128));
    layer0_outputs(6604) <= not(inputs(133));
    layer0_outputs(6605) <= not(inputs(158)) or (inputs(254));
    layer0_outputs(6606) <= inputs(113);
    layer0_outputs(6607) <= not(inputs(8)) or (inputs(212));
    layer0_outputs(6608) <= not(inputs(52));
    layer0_outputs(6609) <= (inputs(157)) or (inputs(28));
    layer0_outputs(6610) <= (inputs(24)) and not (inputs(146));
    layer0_outputs(6611) <= inputs(69);
    layer0_outputs(6612) <= inputs(197);
    layer0_outputs(6613) <= (inputs(205)) xor (inputs(187));
    layer0_outputs(6614) <= not((inputs(102)) and (inputs(104)));
    layer0_outputs(6615) <= not(inputs(245)) or (inputs(3));
    layer0_outputs(6616) <= inputs(176);
    layer0_outputs(6617) <= (inputs(164)) and (inputs(195));
    layer0_outputs(6618) <= not((inputs(89)) xor (inputs(148)));
    layer0_outputs(6619) <= (inputs(125)) xor (inputs(16));
    layer0_outputs(6620) <= not(inputs(161));
    layer0_outputs(6621) <= not((inputs(237)) or (inputs(243)));
    layer0_outputs(6622) <= not((inputs(97)) xor (inputs(47)));
    layer0_outputs(6623) <= (inputs(141)) or (inputs(198));
    layer0_outputs(6624) <= inputs(194);
    layer0_outputs(6625) <= (inputs(239)) xor (inputs(224));
    layer0_outputs(6626) <= '1';
    layer0_outputs(6627) <= (inputs(77)) and not (inputs(18));
    layer0_outputs(6628) <= (inputs(20)) xor (inputs(193));
    layer0_outputs(6629) <= not(inputs(85));
    layer0_outputs(6630) <= inputs(176);
    layer0_outputs(6631) <= not(inputs(202));
    layer0_outputs(6632) <= not(inputs(232));
    layer0_outputs(6633) <= not((inputs(143)) or (inputs(197)));
    layer0_outputs(6634) <= not(inputs(7));
    layer0_outputs(6635) <= not(inputs(14));
    layer0_outputs(6636) <= not((inputs(214)) or (inputs(247)));
    layer0_outputs(6637) <= inputs(139);
    layer0_outputs(6638) <= not((inputs(127)) or (inputs(176)));
    layer0_outputs(6639) <= not(inputs(102));
    layer0_outputs(6640) <= (inputs(214)) xor (inputs(246));
    layer0_outputs(6641) <= (inputs(66)) or (inputs(232));
    layer0_outputs(6642) <= inputs(139);
    layer0_outputs(6643) <= not(inputs(180));
    layer0_outputs(6644) <= not(inputs(244)) or (inputs(29));
    layer0_outputs(6645) <= not((inputs(75)) or (inputs(6)));
    layer0_outputs(6646) <= (inputs(231)) and not (inputs(30));
    layer0_outputs(6647) <= not(inputs(28));
    layer0_outputs(6648) <= inputs(176);
    layer0_outputs(6649) <= (inputs(174)) and (inputs(250));
    layer0_outputs(6650) <= not((inputs(106)) or (inputs(14)));
    layer0_outputs(6651) <= not((inputs(88)) xor (inputs(124)));
    layer0_outputs(6652) <= not(inputs(68));
    layer0_outputs(6653) <= not(inputs(198));
    layer0_outputs(6654) <= not((inputs(19)) or (inputs(127)));
    layer0_outputs(6655) <= (inputs(141)) and (inputs(105));
    layer0_outputs(6656) <= not((inputs(125)) or (inputs(17)));
    layer0_outputs(6657) <= inputs(32);
    layer0_outputs(6658) <= (inputs(24)) and not (inputs(130));
    layer0_outputs(6659) <= (inputs(85)) and not (inputs(32));
    layer0_outputs(6660) <= not(inputs(85));
    layer0_outputs(6661) <= not((inputs(210)) xor (inputs(179)));
    layer0_outputs(6662) <= (inputs(220)) and (inputs(251));
    layer0_outputs(6663) <= not((inputs(126)) or (inputs(197)));
    layer0_outputs(6664) <= not((inputs(228)) xor (inputs(136)));
    layer0_outputs(6665) <= not((inputs(245)) or (inputs(239)));
    layer0_outputs(6666) <= not(inputs(41)) or (inputs(11));
    layer0_outputs(6667) <= inputs(85);
    layer0_outputs(6668) <= not((inputs(164)) or (inputs(198)));
    layer0_outputs(6669) <= not((inputs(95)) or (inputs(247)));
    layer0_outputs(6670) <= inputs(196);
    layer0_outputs(6671) <= not(inputs(213)) or (inputs(89));
    layer0_outputs(6672) <= not(inputs(142));
    layer0_outputs(6673) <= inputs(212);
    layer0_outputs(6674) <= not(inputs(164));
    layer0_outputs(6675) <= not((inputs(201)) or (inputs(196)));
    layer0_outputs(6676) <= (inputs(160)) or (inputs(206));
    layer0_outputs(6677) <= (inputs(211)) xor (inputs(177));
    layer0_outputs(6678) <= (inputs(106)) and not (inputs(31));
    layer0_outputs(6679) <= not(inputs(23));
    layer0_outputs(6680) <= not((inputs(15)) xor (inputs(168)));
    layer0_outputs(6681) <= inputs(115);
    layer0_outputs(6682) <= (inputs(46)) or (inputs(10));
    layer0_outputs(6683) <= (inputs(59)) or (inputs(109));
    layer0_outputs(6684) <= not(inputs(124)) or (inputs(243));
    layer0_outputs(6685) <= not((inputs(22)) and (inputs(226)));
    layer0_outputs(6686) <= (inputs(8)) xor (inputs(85));
    layer0_outputs(6687) <= not((inputs(232)) and (inputs(91)));
    layer0_outputs(6688) <= not(inputs(157)) or (inputs(14));
    layer0_outputs(6689) <= (inputs(103)) xor (inputs(208));
    layer0_outputs(6690) <= (inputs(222)) or (inputs(250));
    layer0_outputs(6691) <= (inputs(147)) xor (inputs(234));
    layer0_outputs(6692) <= (inputs(1)) xor (inputs(108));
    layer0_outputs(6693) <= inputs(48);
    layer0_outputs(6694) <= not((inputs(196)) xor (inputs(7)));
    layer0_outputs(6695) <= not(inputs(199));
    layer0_outputs(6696) <= not(inputs(86));
    layer0_outputs(6697) <= (inputs(10)) and not (inputs(210));
    layer0_outputs(6698) <= not(inputs(253));
    layer0_outputs(6699) <= not((inputs(175)) xor (inputs(160)));
    layer0_outputs(6700) <= inputs(125);
    layer0_outputs(6701) <= not((inputs(120)) xor (inputs(69)));
    layer0_outputs(6702) <= not(inputs(121));
    layer0_outputs(6703) <= inputs(84);
    layer0_outputs(6704) <= inputs(131);
    layer0_outputs(6705) <= not((inputs(9)) xor (inputs(208)));
    layer0_outputs(6706) <= not((inputs(242)) xor (inputs(170)));
    layer0_outputs(6707) <= not(inputs(86)) or (inputs(237));
    layer0_outputs(6708) <= inputs(54);
    layer0_outputs(6709) <= (inputs(14)) and not (inputs(177));
    layer0_outputs(6710) <= inputs(181);
    layer0_outputs(6711) <= (inputs(199)) and not (inputs(76));
    layer0_outputs(6712) <= not((inputs(224)) or (inputs(184)));
    layer0_outputs(6713) <= not(inputs(22));
    layer0_outputs(6714) <= (inputs(4)) or (inputs(94));
    layer0_outputs(6715) <= (inputs(135)) and not (inputs(70));
    layer0_outputs(6716) <= not(inputs(136)) or (inputs(100));
    layer0_outputs(6717) <= not(inputs(58));
    layer0_outputs(6718) <= (inputs(20)) and not (inputs(85));
    layer0_outputs(6719) <= (inputs(126)) or (inputs(142));
    layer0_outputs(6720) <= not((inputs(190)) or (inputs(80)));
    layer0_outputs(6721) <= (inputs(85)) and not (inputs(78));
    layer0_outputs(6722) <= not((inputs(17)) xor (inputs(81)));
    layer0_outputs(6723) <= (inputs(43)) and (inputs(104));
    layer0_outputs(6724) <= inputs(69);
    layer0_outputs(6725) <= not((inputs(8)) xor (inputs(159)));
    layer0_outputs(6726) <= not(inputs(6));
    layer0_outputs(6727) <= not((inputs(181)) or (inputs(49)));
    layer0_outputs(6728) <= inputs(212);
    layer0_outputs(6729) <= inputs(201);
    layer0_outputs(6730) <= not(inputs(36));
    layer0_outputs(6731) <= not((inputs(42)) xor (inputs(31)));
    layer0_outputs(6732) <= not((inputs(26)) xor (inputs(102)));
    layer0_outputs(6733) <= inputs(233);
    layer0_outputs(6734) <= inputs(149);
    layer0_outputs(6735) <= inputs(189);
    layer0_outputs(6736) <= not(inputs(58)) or (inputs(233));
    layer0_outputs(6737) <= not(inputs(167));
    layer0_outputs(6738) <= not(inputs(232));
    layer0_outputs(6739) <= not(inputs(44)) or (inputs(135));
    layer0_outputs(6740) <= (inputs(34)) xor (inputs(151));
    layer0_outputs(6741) <= (inputs(7)) and not (inputs(197));
    layer0_outputs(6742) <= inputs(207);
    layer0_outputs(6743) <= inputs(87);
    layer0_outputs(6744) <= inputs(135);
    layer0_outputs(6745) <= not(inputs(243));
    layer0_outputs(6746) <= not(inputs(23)) or (inputs(146));
    layer0_outputs(6747) <= (inputs(154)) and not (inputs(141));
    layer0_outputs(6748) <= (inputs(22)) or (inputs(236));
    layer0_outputs(6749) <= not(inputs(99));
    layer0_outputs(6750) <= not(inputs(106));
    layer0_outputs(6751) <= not((inputs(130)) or (inputs(214)));
    layer0_outputs(6752) <= (inputs(55)) xor (inputs(71));
    layer0_outputs(6753) <= not(inputs(179));
    layer0_outputs(6754) <= (inputs(62)) or (inputs(80));
    layer0_outputs(6755) <= not((inputs(160)) or (inputs(142)));
    layer0_outputs(6756) <= not((inputs(0)) xor (inputs(7)));
    layer0_outputs(6757) <= not((inputs(123)) xor (inputs(89)));
    layer0_outputs(6758) <= not(inputs(36)) or (inputs(223));
    layer0_outputs(6759) <= not(inputs(248));
    layer0_outputs(6760) <= not((inputs(97)) and (inputs(30)));
    layer0_outputs(6761) <= not(inputs(53));
    layer0_outputs(6762) <= not((inputs(108)) or (inputs(18)));
    layer0_outputs(6763) <= inputs(69);
    layer0_outputs(6764) <= not(inputs(208));
    layer0_outputs(6765) <= not((inputs(88)) and (inputs(172)));
    layer0_outputs(6766) <= (inputs(245)) or (inputs(249));
    layer0_outputs(6767) <= not((inputs(109)) xor (inputs(167)));
    layer0_outputs(6768) <= inputs(254);
    layer0_outputs(6769) <= (inputs(222)) xor (inputs(121));
    layer0_outputs(6770) <= (inputs(16)) xor (inputs(52));
    layer0_outputs(6771) <= not(inputs(87));
    layer0_outputs(6772) <= not((inputs(43)) xor (inputs(70)));
    layer0_outputs(6773) <= inputs(181);
    layer0_outputs(6774) <= not(inputs(229));
    layer0_outputs(6775) <= (inputs(51)) or (inputs(31));
    layer0_outputs(6776) <= (inputs(36)) xor (inputs(82));
    layer0_outputs(6777) <= inputs(173);
    layer0_outputs(6778) <= (inputs(205)) and not (inputs(239));
    layer0_outputs(6779) <= (inputs(218)) and not (inputs(136));
    layer0_outputs(6780) <= not(inputs(187));
    layer0_outputs(6781) <= (inputs(88)) and not (inputs(210));
    layer0_outputs(6782) <= (inputs(139)) and not (inputs(174));
    layer0_outputs(6783) <= (inputs(138)) and not (inputs(75));
    layer0_outputs(6784) <= not((inputs(35)) or (inputs(80)));
    layer0_outputs(6785) <= not((inputs(160)) or (inputs(141)));
    layer0_outputs(6786) <= not((inputs(132)) or (inputs(62)));
    layer0_outputs(6787) <= not(inputs(23));
    layer0_outputs(6788) <= not((inputs(197)) xor (inputs(96)));
    layer0_outputs(6789) <= not((inputs(205)) or (inputs(215)));
    layer0_outputs(6790) <= inputs(232);
    layer0_outputs(6791) <= inputs(17);
    layer0_outputs(6792) <= inputs(215);
    layer0_outputs(6793) <= (inputs(187)) or (inputs(169));
    layer0_outputs(6794) <= not(inputs(113));
    layer0_outputs(6795) <= inputs(89);
    layer0_outputs(6796) <= (inputs(137)) xor (inputs(148));
    layer0_outputs(6797) <= (inputs(20)) and not (inputs(159));
    layer0_outputs(6798) <= not((inputs(201)) or (inputs(232)));
    layer0_outputs(6799) <= not(inputs(187)) or (inputs(110));
    layer0_outputs(6800) <= inputs(34);
    layer0_outputs(6801) <= not(inputs(94)) or (inputs(82));
    layer0_outputs(6802) <= not((inputs(119)) or (inputs(219)));
    layer0_outputs(6803) <= not(inputs(110));
    layer0_outputs(6804) <= not((inputs(145)) and (inputs(211)));
    layer0_outputs(6805) <= inputs(69);
    layer0_outputs(6806) <= (inputs(215)) or (inputs(115));
    layer0_outputs(6807) <= (inputs(114)) and not (inputs(66));
    layer0_outputs(6808) <= not(inputs(109));
    layer0_outputs(6809) <= inputs(82);
    layer0_outputs(6810) <= not(inputs(66)) or (inputs(250));
    layer0_outputs(6811) <= inputs(98);
    layer0_outputs(6812) <= (inputs(32)) and not (inputs(225));
    layer0_outputs(6813) <= not((inputs(77)) and (inputs(106)));
    layer0_outputs(6814) <= (inputs(238)) or (inputs(5));
    layer0_outputs(6815) <= (inputs(215)) and not (inputs(33));
    layer0_outputs(6816) <= not(inputs(67));
    layer0_outputs(6817) <= not(inputs(180)) or (inputs(15));
    layer0_outputs(6818) <= not(inputs(231)) or (inputs(208));
    layer0_outputs(6819) <= not(inputs(60)) or (inputs(194));
    layer0_outputs(6820) <= inputs(128);
    layer0_outputs(6821) <= '0';
    layer0_outputs(6822) <= (inputs(131)) and not (inputs(164));
    layer0_outputs(6823) <= not((inputs(54)) and (inputs(175)));
    layer0_outputs(6824) <= (inputs(49)) and not (inputs(121));
    layer0_outputs(6825) <= not(inputs(182));
    layer0_outputs(6826) <= not(inputs(204)) or (inputs(168));
    layer0_outputs(6827) <= inputs(179);
    layer0_outputs(6828) <= (inputs(159)) or (inputs(170));
    layer0_outputs(6829) <= inputs(48);
    layer0_outputs(6830) <= (inputs(210)) or (inputs(192));
    layer0_outputs(6831) <= not((inputs(134)) or (inputs(234)));
    layer0_outputs(6832) <= not(inputs(255));
    layer0_outputs(6833) <= not(inputs(106));
    layer0_outputs(6834) <= not(inputs(232)) or (inputs(86));
    layer0_outputs(6835) <= (inputs(179)) or (inputs(168));
    layer0_outputs(6836) <= (inputs(5)) or (inputs(207));
    layer0_outputs(6837) <= not(inputs(216));
    layer0_outputs(6838) <= not(inputs(146));
    layer0_outputs(6839) <= not((inputs(244)) or (inputs(19)));
    layer0_outputs(6840) <= not(inputs(154)) or (inputs(147));
    layer0_outputs(6841) <= inputs(13);
    layer0_outputs(6842) <= (inputs(105)) and (inputs(84));
    layer0_outputs(6843) <= (inputs(207)) or (inputs(150));
    layer0_outputs(6844) <= (inputs(8)) xor (inputs(130));
    layer0_outputs(6845) <= not((inputs(152)) or (inputs(253)));
    layer0_outputs(6846) <= not((inputs(60)) xor (inputs(49)));
    layer0_outputs(6847) <= inputs(73);
    layer0_outputs(6848) <= '0';
    layer0_outputs(6849) <= inputs(92);
    layer0_outputs(6850) <= (inputs(144)) or (inputs(155));
    layer0_outputs(6851) <= '0';
    layer0_outputs(6852) <= not(inputs(19)) or (inputs(175));
    layer0_outputs(6853) <= not((inputs(54)) xor (inputs(51)));
    layer0_outputs(6854) <= (inputs(15)) or (inputs(13));
    layer0_outputs(6855) <= not(inputs(201));
    layer0_outputs(6856) <= not((inputs(62)) or (inputs(41)));
    layer0_outputs(6857) <= (inputs(80)) and (inputs(97));
    layer0_outputs(6858) <= inputs(164);
    layer0_outputs(6859) <= (inputs(81)) or (inputs(173));
    layer0_outputs(6860) <= not(inputs(102));
    layer0_outputs(6861) <= inputs(163);
    layer0_outputs(6862) <= (inputs(99)) xor (inputs(101));
    layer0_outputs(6863) <= not((inputs(195)) or (inputs(192)));
    layer0_outputs(6864) <= inputs(225);
    layer0_outputs(6865) <= (inputs(206)) xor (inputs(18));
    layer0_outputs(6866) <= (inputs(56)) or (inputs(23));
    layer0_outputs(6867) <= not((inputs(134)) or (inputs(251)));
    layer0_outputs(6868) <= not(inputs(70));
    layer0_outputs(6869) <= not((inputs(172)) xor (inputs(146)));
    layer0_outputs(6870) <= inputs(113);
    layer0_outputs(6871) <= (inputs(137)) or (inputs(228));
    layer0_outputs(6872) <= inputs(218);
    layer0_outputs(6873) <= inputs(124);
    layer0_outputs(6874) <= not(inputs(79));
    layer0_outputs(6875) <= (inputs(40)) and not (inputs(98));
    layer0_outputs(6876) <= (inputs(247)) xor (inputs(184));
    layer0_outputs(6877) <= not(inputs(71));
    layer0_outputs(6878) <= (inputs(126)) or (inputs(55));
    layer0_outputs(6879) <= not((inputs(197)) or (inputs(5)));
    layer0_outputs(6880) <= not((inputs(219)) or (inputs(223)));
    layer0_outputs(6881) <= inputs(219);
    layer0_outputs(6882) <= (inputs(43)) and not (inputs(5));
    layer0_outputs(6883) <= not(inputs(147));
    layer0_outputs(6884) <= (inputs(74)) or (inputs(98));
    layer0_outputs(6885) <= inputs(144);
    layer0_outputs(6886) <= (inputs(251)) or (inputs(74));
    layer0_outputs(6887) <= (inputs(56)) or (inputs(84));
    layer0_outputs(6888) <= (inputs(149)) or (inputs(193));
    layer0_outputs(6889) <= not(inputs(28));
    layer0_outputs(6890) <= not((inputs(122)) or (inputs(20)));
    layer0_outputs(6891) <= inputs(186);
    layer0_outputs(6892) <= not((inputs(106)) or (inputs(154)));
    layer0_outputs(6893) <= (inputs(212)) or (inputs(49));
    layer0_outputs(6894) <= (inputs(211)) or (inputs(176));
    layer0_outputs(6895) <= (inputs(76)) xor (inputs(90));
    layer0_outputs(6896) <= inputs(35);
    layer0_outputs(6897) <= not((inputs(228)) xor (inputs(10)));
    layer0_outputs(6898) <= (inputs(214)) or (inputs(6));
    layer0_outputs(6899) <= not(inputs(82));
    layer0_outputs(6900) <= not((inputs(87)) or (inputs(187)));
    layer0_outputs(6901) <= not(inputs(211));
    layer0_outputs(6902) <= not(inputs(85));
    layer0_outputs(6903) <= (inputs(222)) or (inputs(142));
    layer0_outputs(6904) <= not((inputs(92)) or (inputs(209)));
    layer0_outputs(6905) <= inputs(166);
    layer0_outputs(6906) <= '1';
    layer0_outputs(6907) <= (inputs(175)) xor (inputs(9));
    layer0_outputs(6908) <= not(inputs(187)) or (inputs(31));
    layer0_outputs(6909) <= (inputs(15)) xor (inputs(217));
    layer0_outputs(6910) <= not(inputs(154));
    layer0_outputs(6911) <= (inputs(7)) or (inputs(111));
    layer0_outputs(6912) <= not(inputs(131));
    layer0_outputs(6913) <= not((inputs(103)) or (inputs(87)));
    layer0_outputs(6914) <= not(inputs(88));
    layer0_outputs(6915) <= (inputs(50)) xor (inputs(238));
    layer0_outputs(6916) <= not(inputs(243));
    layer0_outputs(6917) <= not(inputs(46));
    layer0_outputs(6918) <= not((inputs(197)) or (inputs(82)));
    layer0_outputs(6919) <= not((inputs(114)) xor (inputs(107)));
    layer0_outputs(6920) <= not((inputs(223)) and (inputs(224)));
    layer0_outputs(6921) <= not(inputs(165)) or (inputs(222));
    layer0_outputs(6922) <= not((inputs(83)) xor (inputs(16)));
    layer0_outputs(6923) <= (inputs(94)) xor (inputs(201));
    layer0_outputs(6924) <= not(inputs(165));
    layer0_outputs(6925) <= not(inputs(71));
    layer0_outputs(6926) <= not((inputs(83)) and (inputs(105)));
    layer0_outputs(6927) <= '0';
    layer0_outputs(6928) <= not(inputs(230));
    layer0_outputs(6929) <= not(inputs(101)) or (inputs(21));
    layer0_outputs(6930) <= not(inputs(113));
    layer0_outputs(6931) <= (inputs(25)) xor (inputs(98));
    layer0_outputs(6932) <= (inputs(185)) and not (inputs(61));
    layer0_outputs(6933) <= not(inputs(86));
    layer0_outputs(6934) <= not(inputs(151));
    layer0_outputs(6935) <= '1';
    layer0_outputs(6936) <= not((inputs(36)) or (inputs(21)));
    layer0_outputs(6937) <= not(inputs(64));
    layer0_outputs(6938) <= (inputs(97)) xor (inputs(76));
    layer0_outputs(6939) <= not(inputs(119));
    layer0_outputs(6940) <= not(inputs(60));
    layer0_outputs(6941) <= not(inputs(36));
    layer0_outputs(6942) <= (inputs(210)) and not (inputs(152));
    layer0_outputs(6943) <= not((inputs(162)) or (inputs(29)));
    layer0_outputs(6944) <= inputs(99);
    layer0_outputs(6945) <= not((inputs(115)) and (inputs(122)));
    layer0_outputs(6946) <= not(inputs(87)) or (inputs(239));
    layer0_outputs(6947) <= not(inputs(20));
    layer0_outputs(6948) <= not((inputs(253)) or (inputs(133)));
    layer0_outputs(6949) <= (inputs(136)) or (inputs(233));
    layer0_outputs(6950) <= not(inputs(167)) or (inputs(16));
    layer0_outputs(6951) <= (inputs(157)) and not (inputs(10));
    layer0_outputs(6952) <= (inputs(95)) xor (inputs(54));
    layer0_outputs(6953) <= '1';
    layer0_outputs(6954) <= (inputs(88)) and not (inputs(2));
    layer0_outputs(6955) <= (inputs(188)) xor (inputs(185));
    layer0_outputs(6956) <= (inputs(48)) or (inputs(28));
    layer0_outputs(6957) <= (inputs(99)) xor (inputs(214));
    layer0_outputs(6958) <= not(inputs(141));
    layer0_outputs(6959) <= not(inputs(35));
    layer0_outputs(6960) <= inputs(167);
    layer0_outputs(6961) <= (inputs(151)) xor (inputs(197));
    layer0_outputs(6962) <= not(inputs(176));
    layer0_outputs(6963) <= not(inputs(37));
    layer0_outputs(6964) <= not(inputs(81));
    layer0_outputs(6965) <= not(inputs(22)) or (inputs(160));
    layer0_outputs(6966) <= not(inputs(143));
    layer0_outputs(6967) <= inputs(147);
    layer0_outputs(6968) <= not((inputs(150)) xor (inputs(103)));
    layer0_outputs(6969) <= inputs(121);
    layer0_outputs(6970) <= not(inputs(117));
    layer0_outputs(6971) <= inputs(116);
    layer0_outputs(6972) <= not(inputs(98));
    layer0_outputs(6973) <= (inputs(202)) and not (inputs(78));
    layer0_outputs(6974) <= (inputs(168)) and not (inputs(79));
    layer0_outputs(6975) <= not(inputs(165)) or (inputs(90));
    layer0_outputs(6976) <= (inputs(79)) or (inputs(106));
    layer0_outputs(6977) <= inputs(52);
    layer0_outputs(6978) <= not((inputs(59)) or (inputs(111)));
    layer0_outputs(6979) <= not(inputs(215)) or (inputs(67));
    layer0_outputs(6980) <= inputs(188);
    layer0_outputs(6981) <= inputs(106);
    layer0_outputs(6982) <= not(inputs(99));
    layer0_outputs(6983) <= (inputs(242)) and not (inputs(13));
    layer0_outputs(6984) <= (inputs(213)) and (inputs(113));
    layer0_outputs(6985) <= (inputs(129)) or (inputs(203));
    layer0_outputs(6986) <= inputs(66);
    layer0_outputs(6987) <= not(inputs(6)) or (inputs(128));
    layer0_outputs(6988) <= (inputs(155)) and (inputs(108));
    layer0_outputs(6989) <= (inputs(114)) or (inputs(70));
    layer0_outputs(6990) <= not(inputs(229));
    layer0_outputs(6991) <= not((inputs(239)) and (inputs(13)));
    layer0_outputs(6992) <= (inputs(86)) and not (inputs(78));
    layer0_outputs(6993) <= inputs(253);
    layer0_outputs(6994) <= not(inputs(196)) or (inputs(124));
    layer0_outputs(6995) <= (inputs(90)) and not (inputs(65));
    layer0_outputs(6996) <= inputs(237);
    layer0_outputs(6997) <= (inputs(32)) or (inputs(210));
    layer0_outputs(6998) <= (inputs(176)) or (inputs(94));
    layer0_outputs(6999) <= (inputs(114)) or (inputs(225));
    layer0_outputs(7000) <= inputs(67);
    layer0_outputs(7001) <= not(inputs(109));
    layer0_outputs(7002) <= not((inputs(172)) or (inputs(213)));
    layer0_outputs(7003) <= not(inputs(103)) or (inputs(114));
    layer0_outputs(7004) <= (inputs(188)) or (inputs(2));
    layer0_outputs(7005) <= not(inputs(19)) or (inputs(144));
    layer0_outputs(7006) <= inputs(112);
    layer0_outputs(7007) <= (inputs(83)) and not (inputs(220));
    layer0_outputs(7008) <= inputs(253);
    layer0_outputs(7009) <= (inputs(38)) and not (inputs(206));
    layer0_outputs(7010) <= inputs(24);
    layer0_outputs(7011) <= inputs(253);
    layer0_outputs(7012) <= inputs(146);
    layer0_outputs(7013) <= not(inputs(28));
    layer0_outputs(7014) <= not(inputs(171));
    layer0_outputs(7015) <= not((inputs(84)) or (inputs(102)));
    layer0_outputs(7016) <= (inputs(129)) and not (inputs(122));
    layer0_outputs(7017) <= '1';
    layer0_outputs(7018) <= not((inputs(180)) xor (inputs(178)));
    layer0_outputs(7019) <= (inputs(95)) and not (inputs(4));
    layer0_outputs(7020) <= inputs(59);
    layer0_outputs(7021) <= not(inputs(121));
    layer0_outputs(7022) <= not(inputs(21)) or (inputs(46));
    layer0_outputs(7023) <= not((inputs(205)) or (inputs(43)));
    layer0_outputs(7024) <= not(inputs(3)) or (inputs(249));
    layer0_outputs(7025) <= (inputs(63)) or (inputs(124));
    layer0_outputs(7026) <= not((inputs(200)) xor (inputs(133)));
    layer0_outputs(7027) <= not((inputs(108)) or (inputs(0)));
    layer0_outputs(7028) <= not(inputs(40));
    layer0_outputs(7029) <= (inputs(29)) xor (inputs(11));
    layer0_outputs(7030) <= not((inputs(32)) or (inputs(214)));
    layer0_outputs(7031) <= inputs(37);
    layer0_outputs(7032) <= (inputs(34)) or (inputs(75));
    layer0_outputs(7033) <= (inputs(72)) xor (inputs(26));
    layer0_outputs(7034) <= (inputs(189)) or (inputs(201));
    layer0_outputs(7035) <= not((inputs(240)) or (inputs(223)));
    layer0_outputs(7036) <= not(inputs(99));
    layer0_outputs(7037) <= (inputs(80)) or (inputs(65));
    layer0_outputs(7038) <= not(inputs(183));
    layer0_outputs(7039) <= (inputs(186)) or (inputs(112));
    layer0_outputs(7040) <= (inputs(127)) and not (inputs(64));
    layer0_outputs(7041) <= not(inputs(245));
    layer0_outputs(7042) <= inputs(113);
    layer0_outputs(7043) <= (inputs(91)) or (inputs(113));
    layer0_outputs(7044) <= '0';
    layer0_outputs(7045) <= not(inputs(229));
    layer0_outputs(7046) <= inputs(124);
    layer0_outputs(7047) <= (inputs(24)) xor (inputs(134));
    layer0_outputs(7048) <= not((inputs(213)) or (inputs(213)));
    layer0_outputs(7049) <= (inputs(217)) xor (inputs(91));
    layer0_outputs(7050) <= not((inputs(120)) xor (inputs(88)));
    layer0_outputs(7051) <= not(inputs(89)) or (inputs(81));
    layer0_outputs(7052) <= (inputs(247)) or (inputs(229));
    layer0_outputs(7053) <= inputs(249);
    layer0_outputs(7054) <= not((inputs(34)) or (inputs(23)));
    layer0_outputs(7055) <= not(inputs(157));
    layer0_outputs(7056) <= inputs(34);
    layer0_outputs(7057) <= (inputs(216)) xor (inputs(48));
    layer0_outputs(7058) <= not(inputs(22)) or (inputs(249));
    layer0_outputs(7059) <= (inputs(38)) xor (inputs(7));
    layer0_outputs(7060) <= not((inputs(110)) or (inputs(13)));
    layer0_outputs(7061) <= (inputs(113)) and not (inputs(115));
    layer0_outputs(7062) <= (inputs(14)) xor (inputs(49));
    layer0_outputs(7063) <= (inputs(163)) xor (inputs(116));
    layer0_outputs(7064) <= not(inputs(89));
    layer0_outputs(7065) <= (inputs(199)) and not (inputs(184));
    layer0_outputs(7066) <= '1';
    layer0_outputs(7067) <= not(inputs(162));
    layer0_outputs(7068) <= not((inputs(13)) and (inputs(243)));
    layer0_outputs(7069) <= not((inputs(35)) or (inputs(95)));
    layer0_outputs(7070) <= inputs(106);
    layer0_outputs(7071) <= inputs(61);
    layer0_outputs(7072) <= not((inputs(149)) xor (inputs(209)));
    layer0_outputs(7073) <= not((inputs(119)) or (inputs(87)));
    layer0_outputs(7074) <= (inputs(23)) and not (inputs(164));
    layer0_outputs(7075) <= inputs(202);
    layer0_outputs(7076) <= (inputs(70)) and not (inputs(200));
    layer0_outputs(7077) <= not(inputs(3)) or (inputs(190));
    layer0_outputs(7078) <= not(inputs(8));
    layer0_outputs(7079) <= (inputs(155)) or (inputs(116));
    layer0_outputs(7080) <= not(inputs(170)) or (inputs(98));
    layer0_outputs(7081) <= not((inputs(214)) or (inputs(184)));
    layer0_outputs(7082) <= not(inputs(171)) or (inputs(13));
    layer0_outputs(7083) <= inputs(145);
    layer0_outputs(7084) <= (inputs(56)) xor (inputs(231));
    layer0_outputs(7085) <= (inputs(191)) or (inputs(158));
    layer0_outputs(7086) <= not((inputs(220)) xor (inputs(87)));
    layer0_outputs(7087) <= (inputs(81)) or (inputs(133));
    layer0_outputs(7088) <= not((inputs(26)) and (inputs(164)));
    layer0_outputs(7089) <= not(inputs(26)) or (inputs(229));
    layer0_outputs(7090) <= not(inputs(246)) or (inputs(61));
    layer0_outputs(7091) <= (inputs(179)) and not (inputs(107));
    layer0_outputs(7092) <= (inputs(86)) or (inputs(235));
    layer0_outputs(7093) <= (inputs(138)) or (inputs(237));
    layer0_outputs(7094) <= not(inputs(61)) or (inputs(144));
    layer0_outputs(7095) <= not(inputs(45));
    layer0_outputs(7096) <= not((inputs(157)) or (inputs(96)));
    layer0_outputs(7097) <= (inputs(114)) xor (inputs(186));
    layer0_outputs(7098) <= (inputs(202)) xor (inputs(61));
    layer0_outputs(7099) <= not((inputs(198)) or (inputs(32)));
    layer0_outputs(7100) <= inputs(254);
    layer0_outputs(7101) <= not(inputs(228));
    layer0_outputs(7102) <= inputs(203);
    layer0_outputs(7103) <= not(inputs(168));
    layer0_outputs(7104) <= not(inputs(245));
    layer0_outputs(7105) <= not(inputs(29));
    layer0_outputs(7106) <= (inputs(155)) xor (inputs(202));
    layer0_outputs(7107) <= not(inputs(101)) or (inputs(19));
    layer0_outputs(7108) <= not(inputs(213));
    layer0_outputs(7109) <= (inputs(167)) and not (inputs(113));
    layer0_outputs(7110) <= (inputs(233)) and not (inputs(142));
    layer0_outputs(7111) <= (inputs(200)) or (inputs(84));
    layer0_outputs(7112) <= not(inputs(251));
    layer0_outputs(7113) <= (inputs(116)) or (inputs(102));
    layer0_outputs(7114) <= (inputs(149)) and not (inputs(190));
    layer0_outputs(7115) <= not((inputs(140)) xor (inputs(15)));
    layer0_outputs(7116) <= not((inputs(119)) xor (inputs(86)));
    layer0_outputs(7117) <= (inputs(108)) and not (inputs(31));
    layer0_outputs(7118) <= not(inputs(150));
    layer0_outputs(7119) <= (inputs(93)) and (inputs(194));
    layer0_outputs(7120) <= inputs(26);
    layer0_outputs(7121) <= not(inputs(161));
    layer0_outputs(7122) <= (inputs(243)) or (inputs(109));
    layer0_outputs(7123) <= (inputs(168)) and not (inputs(129));
    layer0_outputs(7124) <= inputs(151);
    layer0_outputs(7125) <= (inputs(153)) or (inputs(245));
    layer0_outputs(7126) <= (inputs(212)) and not (inputs(149));
    layer0_outputs(7127) <= (inputs(80)) xor (inputs(48));
    layer0_outputs(7128) <= not((inputs(160)) xor (inputs(97)));
    layer0_outputs(7129) <= (inputs(187)) and not (inputs(1));
    layer0_outputs(7130) <= not(inputs(90)) or (inputs(201));
    layer0_outputs(7131) <= not(inputs(220)) or (inputs(94));
    layer0_outputs(7132) <= not((inputs(79)) xor (inputs(92)));
    layer0_outputs(7133) <= inputs(147);
    layer0_outputs(7134) <= not(inputs(127));
    layer0_outputs(7135) <= inputs(196);
    layer0_outputs(7136) <= (inputs(14)) and not (inputs(134));
    layer0_outputs(7137) <= (inputs(202)) and not (inputs(23));
    layer0_outputs(7138) <= inputs(177);
    layer0_outputs(7139) <= inputs(131);
    layer0_outputs(7140) <= (inputs(75)) or (inputs(54));
    layer0_outputs(7141) <= (inputs(111)) or (inputs(131));
    layer0_outputs(7142) <= not(inputs(13));
    layer0_outputs(7143) <= not(inputs(142));
    layer0_outputs(7144) <= (inputs(130)) and (inputs(11));
    layer0_outputs(7145) <= (inputs(38)) xor (inputs(143));
    layer0_outputs(7146) <= inputs(195);
    layer0_outputs(7147) <= not(inputs(230));
    layer0_outputs(7148) <= not((inputs(146)) or (inputs(204)));
    layer0_outputs(7149) <= '1';
    layer0_outputs(7150) <= not(inputs(130));
    layer0_outputs(7151) <= (inputs(157)) and not (inputs(29));
    layer0_outputs(7152) <= (inputs(99)) and not (inputs(47));
    layer0_outputs(7153) <= (inputs(177)) or (inputs(160));
    layer0_outputs(7154) <= not((inputs(111)) or (inputs(150)));
    layer0_outputs(7155) <= not(inputs(13)) or (inputs(145));
    layer0_outputs(7156) <= (inputs(71)) and (inputs(67));
    layer0_outputs(7157) <= not(inputs(117));
    layer0_outputs(7158) <= (inputs(198)) xor (inputs(230));
    layer0_outputs(7159) <= not((inputs(158)) or (inputs(159)));
    layer0_outputs(7160) <= (inputs(9)) xor (inputs(127));
    layer0_outputs(7161) <= inputs(167);
    layer0_outputs(7162) <= (inputs(152)) xor (inputs(90));
    layer0_outputs(7163) <= '0';
    layer0_outputs(7164) <= (inputs(141)) or (inputs(50));
    layer0_outputs(7165) <= inputs(131);
    layer0_outputs(7166) <= inputs(180);
    layer0_outputs(7167) <= not((inputs(140)) xor (inputs(202)));
    layer0_outputs(7168) <= not(inputs(106));
    layer0_outputs(7169) <= inputs(186);
    layer0_outputs(7170) <= not(inputs(160)) or (inputs(72));
    layer0_outputs(7171) <= inputs(42);
    layer0_outputs(7172) <= (inputs(195)) xor (inputs(224));
    layer0_outputs(7173) <= not(inputs(70)) or (inputs(33));
    layer0_outputs(7174) <= (inputs(218)) xor (inputs(65));
    layer0_outputs(7175) <= inputs(22);
    layer0_outputs(7176) <= inputs(241);
    layer0_outputs(7177) <= (inputs(73)) and not (inputs(224));
    layer0_outputs(7178) <= (inputs(164)) and not (inputs(12));
    layer0_outputs(7179) <= not(inputs(228));
    layer0_outputs(7180) <= not(inputs(175)) or (inputs(128));
    layer0_outputs(7181) <= not(inputs(177));
    layer0_outputs(7182) <= (inputs(20)) and not (inputs(146));
    layer0_outputs(7183) <= (inputs(245)) and (inputs(199));
    layer0_outputs(7184) <= (inputs(55)) or (inputs(176));
    layer0_outputs(7185) <= (inputs(112)) or (inputs(29));
    layer0_outputs(7186) <= '1';
    layer0_outputs(7187) <= (inputs(227)) or (inputs(232));
    layer0_outputs(7188) <= not(inputs(71));
    layer0_outputs(7189) <= (inputs(138)) or (inputs(239));
    layer0_outputs(7190) <= not(inputs(174));
    layer0_outputs(7191) <= (inputs(103)) or (inputs(220));
    layer0_outputs(7192) <= (inputs(210)) or (inputs(8));
    layer0_outputs(7193) <= not((inputs(231)) xor (inputs(184)));
    layer0_outputs(7194) <= not(inputs(91));
    layer0_outputs(7195) <= (inputs(90)) or (inputs(110));
    layer0_outputs(7196) <= not((inputs(29)) xor (inputs(12)));
    layer0_outputs(7197) <= (inputs(40)) and not (inputs(160));
    layer0_outputs(7198) <= not(inputs(133));
    layer0_outputs(7199) <= (inputs(182)) or (inputs(131));
    layer0_outputs(7200) <= inputs(116);
    layer0_outputs(7201) <= (inputs(106)) and not (inputs(94));
    layer0_outputs(7202) <= (inputs(164)) or (inputs(238));
    layer0_outputs(7203) <= not(inputs(228)) or (inputs(125));
    layer0_outputs(7204) <= (inputs(249)) and not (inputs(170));
    layer0_outputs(7205) <= (inputs(154)) xor (inputs(123));
    layer0_outputs(7206) <= (inputs(234)) xor (inputs(96));
    layer0_outputs(7207) <= (inputs(243)) and not (inputs(144));
    layer0_outputs(7208) <= not(inputs(246)) or (inputs(76));
    layer0_outputs(7209) <= inputs(23);
    layer0_outputs(7210) <= not((inputs(31)) or (inputs(170)));
    layer0_outputs(7211) <= not(inputs(28)) or (inputs(252));
    layer0_outputs(7212) <= not(inputs(25));
    layer0_outputs(7213) <= not((inputs(48)) or (inputs(77)));
    layer0_outputs(7214) <= inputs(122);
    layer0_outputs(7215) <= (inputs(1)) xor (inputs(140));
    layer0_outputs(7216) <= (inputs(93)) and not (inputs(81));
    layer0_outputs(7217) <= not(inputs(5)) or (inputs(30));
    layer0_outputs(7218) <= (inputs(118)) xor (inputs(87));
    layer0_outputs(7219) <= not((inputs(221)) or (inputs(216)));
    layer0_outputs(7220) <= inputs(143);
    layer0_outputs(7221) <= not(inputs(74));
    layer0_outputs(7222) <= (inputs(135)) and not (inputs(229));
    layer0_outputs(7223) <= not((inputs(121)) xor (inputs(169)));
    layer0_outputs(7224) <= not((inputs(133)) and (inputs(153)));
    layer0_outputs(7225) <= not(inputs(145));
    layer0_outputs(7226) <= not(inputs(146));
    layer0_outputs(7227) <= not((inputs(97)) xor (inputs(85)));
    layer0_outputs(7228) <= not((inputs(206)) and (inputs(2)));
    layer0_outputs(7229) <= not((inputs(171)) or (inputs(219)));
    layer0_outputs(7230) <= not((inputs(83)) or (inputs(37)));
    layer0_outputs(7231) <= not(inputs(230));
    layer0_outputs(7232) <= '0';
    layer0_outputs(7233) <= inputs(178);
    layer0_outputs(7234) <= not(inputs(209)) or (inputs(67));
    layer0_outputs(7235) <= inputs(47);
    layer0_outputs(7236) <= not(inputs(206)) or (inputs(45));
    layer0_outputs(7237) <= inputs(91);
    layer0_outputs(7238) <= not((inputs(165)) xor (inputs(192)));
    layer0_outputs(7239) <= (inputs(131)) xor (inputs(134));
    layer0_outputs(7240) <= (inputs(55)) and not (inputs(31));
    layer0_outputs(7241) <= inputs(95);
    layer0_outputs(7242) <= not((inputs(37)) xor (inputs(21)));
    layer0_outputs(7243) <= not(inputs(66)) or (inputs(33));
    layer0_outputs(7244) <= not(inputs(47)) or (inputs(147));
    layer0_outputs(7245) <= not((inputs(133)) or (inputs(132)));
    layer0_outputs(7246) <= not((inputs(125)) or (inputs(253)));
    layer0_outputs(7247) <= not(inputs(95)) or (inputs(237));
    layer0_outputs(7248) <= not(inputs(123));
    layer0_outputs(7249) <= not(inputs(68)) or (inputs(63));
    layer0_outputs(7250) <= not((inputs(73)) xor (inputs(91)));
    layer0_outputs(7251) <= '1';
    layer0_outputs(7252) <= inputs(128);
    layer0_outputs(7253) <= (inputs(34)) xor (inputs(56));
    layer0_outputs(7254) <= (inputs(63)) and not (inputs(14));
    layer0_outputs(7255) <= not(inputs(41)) or (inputs(85));
    layer0_outputs(7256) <= (inputs(167)) and (inputs(151));
    layer0_outputs(7257) <= (inputs(164)) and (inputs(64));
    layer0_outputs(7258) <= not(inputs(198));
    layer0_outputs(7259) <= not(inputs(74));
    layer0_outputs(7260) <= (inputs(180)) xor (inputs(193));
    layer0_outputs(7261) <= not(inputs(134)) or (inputs(72));
    layer0_outputs(7262) <= (inputs(3)) or (inputs(46));
    layer0_outputs(7263) <= not(inputs(130));
    layer0_outputs(7264) <= inputs(251);
    layer0_outputs(7265) <= (inputs(204)) and not (inputs(16));
    layer0_outputs(7266) <= (inputs(217)) xor (inputs(150));
    layer0_outputs(7267) <= inputs(166);
    layer0_outputs(7268) <= not((inputs(162)) or (inputs(96)));
    layer0_outputs(7269) <= (inputs(196)) or (inputs(85));
    layer0_outputs(7270) <= not((inputs(172)) or (inputs(157)));
    layer0_outputs(7271) <= (inputs(8)) and not (inputs(220));
    layer0_outputs(7272) <= not(inputs(207));
    layer0_outputs(7273) <= (inputs(42)) xor (inputs(205));
    layer0_outputs(7274) <= not(inputs(142));
    layer0_outputs(7275) <= not((inputs(115)) xor (inputs(44)));
    layer0_outputs(7276) <= not((inputs(141)) or (inputs(132)));
    layer0_outputs(7277) <= not(inputs(109));
    layer0_outputs(7278) <= inputs(52);
    layer0_outputs(7279) <= (inputs(100)) and not (inputs(41));
    layer0_outputs(7280) <= (inputs(75)) or (inputs(136));
    layer0_outputs(7281) <= (inputs(80)) or (inputs(148));
    layer0_outputs(7282) <= (inputs(250)) or (inputs(153));
    layer0_outputs(7283) <= not((inputs(163)) and (inputs(126)));
    layer0_outputs(7284) <= '0';
    layer0_outputs(7285) <= not((inputs(97)) xor (inputs(81)));
    layer0_outputs(7286) <= inputs(64);
    layer0_outputs(7287) <= not((inputs(37)) or (inputs(95)));
    layer0_outputs(7288) <= not((inputs(143)) xor (inputs(248)));
    layer0_outputs(7289) <= not(inputs(181)) or (inputs(188));
    layer0_outputs(7290) <= not(inputs(89)) or (inputs(68));
    layer0_outputs(7291) <= not(inputs(151));
    layer0_outputs(7292) <= '0';
    layer0_outputs(7293) <= not((inputs(197)) or (inputs(123)));
    layer0_outputs(7294) <= not((inputs(209)) or (inputs(182)));
    layer0_outputs(7295) <= (inputs(171)) xor (inputs(37));
    layer0_outputs(7296) <= (inputs(49)) xor (inputs(220));
    layer0_outputs(7297) <= (inputs(155)) and not (inputs(197));
    layer0_outputs(7298) <= not(inputs(192));
    layer0_outputs(7299) <= not(inputs(247)) or (inputs(95));
    layer0_outputs(7300) <= inputs(65);
    layer0_outputs(7301) <= not((inputs(188)) xor (inputs(246)));
    layer0_outputs(7302) <= not((inputs(181)) or (inputs(251)));
    layer0_outputs(7303) <= not(inputs(37)) or (inputs(176));
    layer0_outputs(7304) <= not(inputs(130)) or (inputs(71));
    layer0_outputs(7305) <= '0';
    layer0_outputs(7306) <= inputs(54);
    layer0_outputs(7307) <= not(inputs(57));
    layer0_outputs(7308) <= not(inputs(69));
    layer0_outputs(7309) <= not((inputs(25)) or (inputs(18)));
    layer0_outputs(7310) <= inputs(229);
    layer0_outputs(7311) <= (inputs(95)) or (inputs(33));
    layer0_outputs(7312) <= not((inputs(242)) or (inputs(138)));
    layer0_outputs(7313) <= not((inputs(215)) xor (inputs(207)));
    layer0_outputs(7314) <= not(inputs(148));
    layer0_outputs(7315) <= (inputs(39)) and not (inputs(217));
    layer0_outputs(7316) <= inputs(190);
    layer0_outputs(7317) <= '0';
    layer0_outputs(7318) <= (inputs(148)) and not (inputs(206));
    layer0_outputs(7319) <= (inputs(165)) or (inputs(188));
    layer0_outputs(7320) <= not((inputs(202)) xor (inputs(144)));
    layer0_outputs(7321) <= not(inputs(195));
    layer0_outputs(7322) <= not(inputs(210));
    layer0_outputs(7323) <= inputs(53);
    layer0_outputs(7324) <= inputs(74);
    layer0_outputs(7325) <= inputs(13);
    layer0_outputs(7326) <= inputs(99);
    layer0_outputs(7327) <= not(inputs(137)) or (inputs(111));
    layer0_outputs(7328) <= '0';
    layer0_outputs(7329) <= inputs(130);
    layer0_outputs(7330) <= not(inputs(45)) or (inputs(18));
    layer0_outputs(7331) <= not(inputs(229));
    layer0_outputs(7332) <= (inputs(53)) and not (inputs(126));
    layer0_outputs(7333) <= (inputs(196)) xor (inputs(243));
    layer0_outputs(7334) <= not((inputs(135)) or (inputs(183)));
    layer0_outputs(7335) <= not((inputs(8)) xor (inputs(39)));
    layer0_outputs(7336) <= not(inputs(177));
    layer0_outputs(7337) <= (inputs(157)) or (inputs(10));
    layer0_outputs(7338) <= (inputs(140)) and (inputs(114));
    layer0_outputs(7339) <= not((inputs(74)) or (inputs(73)));
    layer0_outputs(7340) <= not(inputs(98));
    layer0_outputs(7341) <= (inputs(187)) xor (inputs(195));
    layer0_outputs(7342) <= (inputs(89)) xor (inputs(97));
    layer0_outputs(7343) <= (inputs(24)) and not (inputs(250));
    layer0_outputs(7344) <= not(inputs(24)) or (inputs(242));
    layer0_outputs(7345) <= not(inputs(46)) or (inputs(187));
    layer0_outputs(7346) <= (inputs(53)) xor (inputs(185));
    layer0_outputs(7347) <= (inputs(232)) xor (inputs(160));
    layer0_outputs(7348) <= (inputs(95)) or (inputs(170));
    layer0_outputs(7349) <= (inputs(9)) xor (inputs(217));
    layer0_outputs(7350) <= not(inputs(119));
    layer0_outputs(7351) <= (inputs(140)) and (inputs(136));
    layer0_outputs(7352) <= (inputs(49)) xor (inputs(233));
    layer0_outputs(7353) <= '0';
    layer0_outputs(7354) <= (inputs(34)) xor (inputs(173));
    layer0_outputs(7355) <= not((inputs(65)) or (inputs(165)));
    layer0_outputs(7356) <= inputs(167);
    layer0_outputs(7357) <= not((inputs(104)) or (inputs(238)));
    layer0_outputs(7358) <= not((inputs(193)) or (inputs(211)));
    layer0_outputs(7359) <= inputs(62);
    layer0_outputs(7360) <= (inputs(182)) or (inputs(231));
    layer0_outputs(7361) <= inputs(73);
    layer0_outputs(7362) <= not(inputs(131));
    layer0_outputs(7363) <= (inputs(105)) and not (inputs(143));
    layer0_outputs(7364) <= not(inputs(95));
    layer0_outputs(7365) <= not((inputs(135)) or (inputs(75)));
    layer0_outputs(7366) <= inputs(214);
    layer0_outputs(7367) <= (inputs(126)) or (inputs(201));
    layer0_outputs(7368) <= not(inputs(0)) or (inputs(179));
    layer0_outputs(7369) <= (inputs(119)) and not (inputs(159));
    layer0_outputs(7370) <= not(inputs(3)) or (inputs(33));
    layer0_outputs(7371) <= inputs(53);
    layer0_outputs(7372) <= not((inputs(204)) xor (inputs(197)));
    layer0_outputs(7373) <= not(inputs(17)) or (inputs(128));
    layer0_outputs(7374) <= not(inputs(59)) or (inputs(178));
    layer0_outputs(7375) <= (inputs(118)) and not (inputs(149));
    layer0_outputs(7376) <= not(inputs(199)) or (inputs(53));
    layer0_outputs(7377) <= not(inputs(84));
    layer0_outputs(7378) <= (inputs(19)) or (inputs(188));
    layer0_outputs(7379) <= not((inputs(141)) and (inputs(158)));
    layer0_outputs(7380) <= not(inputs(179)) or (inputs(35));
    layer0_outputs(7381) <= (inputs(112)) or (inputs(34));
    layer0_outputs(7382) <= (inputs(213)) or (inputs(249));
    layer0_outputs(7383) <= (inputs(114)) and not (inputs(221));
    layer0_outputs(7384) <= not((inputs(234)) and (inputs(140)));
    layer0_outputs(7385) <= (inputs(158)) and not (inputs(112));
    layer0_outputs(7386) <= not(inputs(68));
    layer0_outputs(7387) <= not((inputs(125)) or (inputs(47)));
    layer0_outputs(7388) <= not((inputs(62)) or (inputs(195)));
    layer0_outputs(7389) <= (inputs(69)) and (inputs(186));
    layer0_outputs(7390) <= inputs(167);
    layer0_outputs(7391) <= inputs(98);
    layer0_outputs(7392) <= not((inputs(234)) xor (inputs(107)));
    layer0_outputs(7393) <= inputs(100);
    layer0_outputs(7394) <= inputs(183);
    layer0_outputs(7395) <= '1';
    layer0_outputs(7396) <= (inputs(69)) and not (inputs(224));
    layer0_outputs(7397) <= inputs(168);
    layer0_outputs(7398) <= not((inputs(14)) xor (inputs(56)));
    layer0_outputs(7399) <= (inputs(157)) or (inputs(9));
    layer0_outputs(7400) <= not(inputs(162)) or (inputs(64));
    layer0_outputs(7401) <= not((inputs(245)) or (inputs(98)));
    layer0_outputs(7402) <= not(inputs(75));
    layer0_outputs(7403) <= (inputs(185)) xor (inputs(218));
    layer0_outputs(7404) <= inputs(167);
    layer0_outputs(7405) <= not((inputs(96)) or (inputs(165)));
    layer0_outputs(7406) <= (inputs(202)) or (inputs(18));
    layer0_outputs(7407) <= (inputs(63)) or (inputs(233));
    layer0_outputs(7408) <= not((inputs(222)) xor (inputs(180)));
    layer0_outputs(7409) <= (inputs(77)) or (inputs(3));
    layer0_outputs(7410) <= not((inputs(188)) xor (inputs(221)));
    layer0_outputs(7411) <= not((inputs(188)) xor (inputs(129)));
    layer0_outputs(7412) <= not(inputs(54));
    layer0_outputs(7413) <= (inputs(252)) and (inputs(252));
    layer0_outputs(7414) <= '1';
    layer0_outputs(7415) <= (inputs(246)) or (inputs(229));
    layer0_outputs(7416) <= not(inputs(219));
    layer0_outputs(7417) <= inputs(105);
    layer0_outputs(7418) <= not((inputs(182)) or (inputs(226)));
    layer0_outputs(7419) <= (inputs(96)) or (inputs(238));
    layer0_outputs(7420) <= (inputs(224)) and not (inputs(30));
    layer0_outputs(7421) <= not(inputs(163));
    layer0_outputs(7422) <= not(inputs(22));
    layer0_outputs(7423) <= not(inputs(94)) or (inputs(153));
    layer0_outputs(7424) <= not((inputs(178)) or (inputs(24)));
    layer0_outputs(7425) <= not((inputs(38)) and (inputs(102)));
    layer0_outputs(7426) <= (inputs(231)) or (inputs(246));
    layer0_outputs(7427) <= not(inputs(100));
    layer0_outputs(7428) <= not((inputs(5)) xor (inputs(70)));
    layer0_outputs(7429) <= (inputs(11)) and (inputs(131));
    layer0_outputs(7430) <= (inputs(12)) and not (inputs(79));
    layer0_outputs(7431) <= (inputs(7)) or (inputs(204));
    layer0_outputs(7432) <= inputs(183);
    layer0_outputs(7433) <= not((inputs(216)) or (inputs(226)));
    layer0_outputs(7434) <= inputs(226);
    layer0_outputs(7435) <= inputs(121);
    layer0_outputs(7436) <= (inputs(74)) and not (inputs(201));
    layer0_outputs(7437) <= (inputs(163)) and not (inputs(222));
    layer0_outputs(7438) <= inputs(151);
    layer0_outputs(7439) <= '0';
    layer0_outputs(7440) <= not(inputs(120));
    layer0_outputs(7441) <= not((inputs(102)) xor (inputs(169)));
    layer0_outputs(7442) <= inputs(169);
    layer0_outputs(7443) <= not(inputs(210)) or (inputs(139));
    layer0_outputs(7444) <= not(inputs(130));
    layer0_outputs(7445) <= '1';
    layer0_outputs(7446) <= not((inputs(45)) or (inputs(108)));
    layer0_outputs(7447) <= inputs(179);
    layer0_outputs(7448) <= not(inputs(247));
    layer0_outputs(7449) <= inputs(140);
    layer0_outputs(7450) <= not(inputs(49));
    layer0_outputs(7451) <= (inputs(228)) and not (inputs(86));
    layer0_outputs(7452) <= not((inputs(84)) xor (inputs(38)));
    layer0_outputs(7453) <= not((inputs(223)) or (inputs(206)));
    layer0_outputs(7454) <= inputs(10);
    layer0_outputs(7455) <= not(inputs(91)) or (inputs(159));
    layer0_outputs(7456) <= not(inputs(130)) or (inputs(237));
    layer0_outputs(7457) <= inputs(134);
    layer0_outputs(7458) <= not(inputs(194)) or (inputs(122));
    layer0_outputs(7459) <= inputs(73);
    layer0_outputs(7460) <= (inputs(113)) xor (inputs(36));
    layer0_outputs(7461) <= (inputs(219)) or (inputs(162));
    layer0_outputs(7462) <= not((inputs(78)) and (inputs(43)));
    layer0_outputs(7463) <= '0';
    layer0_outputs(7464) <= not(inputs(38));
    layer0_outputs(7465) <= not(inputs(53)) or (inputs(13));
    layer0_outputs(7466) <= inputs(175);
    layer0_outputs(7467) <= not((inputs(71)) xor (inputs(45)));
    layer0_outputs(7468) <= (inputs(92)) or (inputs(246));
    layer0_outputs(7469) <= not(inputs(59)) or (inputs(253));
    layer0_outputs(7470) <= inputs(112);
    layer0_outputs(7471) <= (inputs(207)) or (inputs(62));
    layer0_outputs(7472) <= (inputs(17)) and (inputs(144));
    layer0_outputs(7473) <= not((inputs(254)) and (inputs(168)));
    layer0_outputs(7474) <= not(inputs(222));
    layer0_outputs(7475) <= not((inputs(216)) or (inputs(228)));
    layer0_outputs(7476) <= inputs(19);
    layer0_outputs(7477) <= not(inputs(117));
    layer0_outputs(7478) <= not(inputs(92));
    layer0_outputs(7479) <= not(inputs(53));
    layer0_outputs(7480) <= not(inputs(214)) or (inputs(52));
    layer0_outputs(7481) <= (inputs(141)) or (inputs(219));
    layer0_outputs(7482) <= inputs(26);
    layer0_outputs(7483) <= not((inputs(211)) xor (inputs(110)));
    layer0_outputs(7484) <= (inputs(222)) xor (inputs(251));
    layer0_outputs(7485) <= (inputs(45)) and not (inputs(240));
    layer0_outputs(7486) <= not((inputs(243)) xor (inputs(197)));
    layer0_outputs(7487) <= (inputs(97)) or (inputs(109));
    layer0_outputs(7488) <= (inputs(212)) xor (inputs(180));
    layer0_outputs(7489) <= not((inputs(240)) or (inputs(30)));
    layer0_outputs(7490) <= inputs(134);
    layer0_outputs(7491) <= not((inputs(89)) or (inputs(120)));
    layer0_outputs(7492) <= not((inputs(136)) xor (inputs(26)));
    layer0_outputs(7493) <= not(inputs(158));
    layer0_outputs(7494) <= (inputs(27)) and not (inputs(209));
    layer0_outputs(7495) <= inputs(92);
    layer0_outputs(7496) <= (inputs(213)) or (inputs(211));
    layer0_outputs(7497) <= not(inputs(175));
    layer0_outputs(7498) <= (inputs(114)) or (inputs(99));
    layer0_outputs(7499) <= not(inputs(159));
    layer0_outputs(7500) <= inputs(80);
    layer0_outputs(7501) <= (inputs(154)) and not (inputs(78));
    layer0_outputs(7502) <= not((inputs(243)) or (inputs(150)));
    layer0_outputs(7503) <= not(inputs(232));
    layer0_outputs(7504) <= '0';
    layer0_outputs(7505) <= not((inputs(105)) xor (inputs(203)));
    layer0_outputs(7506) <= (inputs(128)) or (inputs(76));
    layer0_outputs(7507) <= not((inputs(189)) or (inputs(29)));
    layer0_outputs(7508) <= inputs(77);
    layer0_outputs(7509) <= '0';
    layer0_outputs(7510) <= (inputs(80)) or (inputs(82));
    layer0_outputs(7511) <= (inputs(116)) or (inputs(149));
    layer0_outputs(7512) <= (inputs(9)) and not (inputs(226));
    layer0_outputs(7513) <= not((inputs(252)) or (inputs(56)));
    layer0_outputs(7514) <= not(inputs(120));
    layer0_outputs(7515) <= (inputs(132)) and not (inputs(32));
    layer0_outputs(7516) <= not(inputs(40)) or (inputs(153));
    layer0_outputs(7517) <= (inputs(191)) or (inputs(140));
    layer0_outputs(7518) <= not(inputs(9));
    layer0_outputs(7519) <= (inputs(228)) and (inputs(116));
    layer0_outputs(7520) <= (inputs(180)) or (inputs(66));
    layer0_outputs(7521) <= not((inputs(86)) or (inputs(154)));
    layer0_outputs(7522) <= (inputs(87)) and not (inputs(188));
    layer0_outputs(7523) <= not(inputs(45)) or (inputs(191));
    layer0_outputs(7524) <= not((inputs(93)) xor (inputs(35)));
    layer0_outputs(7525) <= not(inputs(161));
    layer0_outputs(7526) <= (inputs(211)) and (inputs(45));
    layer0_outputs(7527) <= inputs(122);
    layer0_outputs(7528) <= not((inputs(97)) or (inputs(92)));
    layer0_outputs(7529) <= inputs(120);
    layer0_outputs(7530) <= inputs(162);
    layer0_outputs(7531) <= not((inputs(250)) or (inputs(134)));
    layer0_outputs(7532) <= not(inputs(104));
    layer0_outputs(7533) <= not((inputs(130)) xor (inputs(255)));
    layer0_outputs(7534) <= (inputs(246)) and (inputs(107));
    layer0_outputs(7535) <= (inputs(236)) and not (inputs(50));
    layer0_outputs(7536) <= not(inputs(204));
    layer0_outputs(7537) <= not(inputs(121)) or (inputs(244));
    layer0_outputs(7538) <= inputs(130);
    layer0_outputs(7539) <= (inputs(177)) and not (inputs(139));
    layer0_outputs(7540) <= not((inputs(172)) and (inputs(196)));
    layer0_outputs(7541) <= inputs(66);
    layer0_outputs(7542) <= not(inputs(167));
    layer0_outputs(7543) <= not(inputs(225));
    layer0_outputs(7544) <= inputs(89);
    layer0_outputs(7545) <= not(inputs(51)) or (inputs(143));
    layer0_outputs(7546) <= not(inputs(89));
    layer0_outputs(7547) <= inputs(211);
    layer0_outputs(7548) <= not(inputs(70));
    layer0_outputs(7549) <= not(inputs(125));
    layer0_outputs(7550) <= not(inputs(94));
    layer0_outputs(7551) <= inputs(57);
    layer0_outputs(7552) <= (inputs(219)) and not (inputs(151));
    layer0_outputs(7553) <= inputs(161);
    layer0_outputs(7554) <= (inputs(21)) xor (inputs(231));
    layer0_outputs(7555) <= not(inputs(185)) or (inputs(31));
    layer0_outputs(7556) <= not((inputs(217)) or (inputs(184)));
    layer0_outputs(7557) <= (inputs(72)) and not (inputs(50));
    layer0_outputs(7558) <= not(inputs(210));
    layer0_outputs(7559) <= not((inputs(143)) or (inputs(224)));
    layer0_outputs(7560) <= (inputs(126)) or (inputs(131));
    layer0_outputs(7561) <= not(inputs(110));
    layer0_outputs(7562) <= not((inputs(209)) xor (inputs(96)));
    layer0_outputs(7563) <= not((inputs(71)) or (inputs(93)));
    layer0_outputs(7564) <= '0';
    layer0_outputs(7565) <= inputs(69);
    layer0_outputs(7566) <= (inputs(75)) and not (inputs(158));
    layer0_outputs(7567) <= inputs(24);
    layer0_outputs(7568) <= (inputs(117)) and not (inputs(57));
    layer0_outputs(7569) <= inputs(8);
    layer0_outputs(7570) <= not((inputs(44)) xor (inputs(90)));
    layer0_outputs(7571) <= not((inputs(47)) or (inputs(106)));
    layer0_outputs(7572) <= not(inputs(100));
    layer0_outputs(7573) <= (inputs(227)) xor (inputs(108));
    layer0_outputs(7574) <= not((inputs(221)) or (inputs(182)));
    layer0_outputs(7575) <= (inputs(1)) xor (inputs(183));
    layer0_outputs(7576) <= not(inputs(203));
    layer0_outputs(7577) <= inputs(225);
    layer0_outputs(7578) <= (inputs(227)) or (inputs(71));
    layer0_outputs(7579) <= not((inputs(138)) xor (inputs(77)));
    layer0_outputs(7580) <= inputs(210);
    layer0_outputs(7581) <= (inputs(172)) and (inputs(228));
    layer0_outputs(7582) <= '0';
    layer0_outputs(7583) <= not((inputs(180)) or (inputs(68)));
    layer0_outputs(7584) <= (inputs(153)) and not (inputs(77));
    layer0_outputs(7585) <= inputs(231);
    layer0_outputs(7586) <= inputs(62);
    layer0_outputs(7587) <= (inputs(61)) or (inputs(20));
    layer0_outputs(7588) <= (inputs(111)) xor (inputs(123));
    layer0_outputs(7589) <= not((inputs(216)) and (inputs(72)));
    layer0_outputs(7590) <= not(inputs(231)) or (inputs(237));
    layer0_outputs(7591) <= not(inputs(171)) or (inputs(2));
    layer0_outputs(7592) <= (inputs(221)) xor (inputs(128));
    layer0_outputs(7593) <= (inputs(194)) or (inputs(85));
    layer0_outputs(7594) <= (inputs(0)) and not (inputs(55));
    layer0_outputs(7595) <= not((inputs(90)) xor (inputs(249)));
    layer0_outputs(7596) <= (inputs(82)) or (inputs(115));
    layer0_outputs(7597) <= (inputs(187)) and not (inputs(149));
    layer0_outputs(7598) <= not(inputs(41));
    layer0_outputs(7599) <= (inputs(15)) or (inputs(12));
    layer0_outputs(7600) <= (inputs(150)) or (inputs(41));
    layer0_outputs(7601) <= (inputs(95)) or (inputs(76));
    layer0_outputs(7602) <= not(inputs(13));
    layer0_outputs(7603) <= (inputs(247)) and not (inputs(69));
    layer0_outputs(7604) <= inputs(162);
    layer0_outputs(7605) <= not(inputs(29)) or (inputs(43));
    layer0_outputs(7606) <= inputs(77);
    layer0_outputs(7607) <= (inputs(37)) and not (inputs(83));
    layer0_outputs(7608) <= inputs(62);
    layer0_outputs(7609) <= not(inputs(136)) or (inputs(238));
    layer0_outputs(7610) <= not(inputs(156));
    layer0_outputs(7611) <= inputs(165);
    layer0_outputs(7612) <= not(inputs(102));
    layer0_outputs(7613) <= not((inputs(216)) xor (inputs(232)));
    layer0_outputs(7614) <= not((inputs(202)) and (inputs(77)));
    layer0_outputs(7615) <= (inputs(136)) and not (inputs(250));
    layer0_outputs(7616) <= not((inputs(123)) or (inputs(51)));
    layer0_outputs(7617) <= not(inputs(176));
    layer0_outputs(7618) <= inputs(120);
    layer0_outputs(7619) <= not((inputs(199)) or (inputs(179)));
    layer0_outputs(7620) <= inputs(180);
    layer0_outputs(7621) <= not(inputs(137)) or (inputs(189));
    layer0_outputs(7622) <= not((inputs(20)) or (inputs(68)));
    layer0_outputs(7623) <= not((inputs(45)) xor (inputs(11)));
    layer0_outputs(7624) <= not((inputs(163)) xor (inputs(137)));
    layer0_outputs(7625) <= not((inputs(182)) and (inputs(198)));
    layer0_outputs(7626) <= not((inputs(8)) or (inputs(47)));
    layer0_outputs(7627) <= (inputs(242)) xor (inputs(215));
    layer0_outputs(7628) <= (inputs(4)) xor (inputs(114));
    layer0_outputs(7629) <= not((inputs(11)) or (inputs(83)));
    layer0_outputs(7630) <= '1';
    layer0_outputs(7631) <= (inputs(185)) xor (inputs(234));
    layer0_outputs(7632) <= (inputs(156)) and not (inputs(255));
    layer0_outputs(7633) <= not(inputs(113)) or (inputs(223));
    layer0_outputs(7634) <= not(inputs(168)) or (inputs(158));
    layer0_outputs(7635) <= not((inputs(45)) or (inputs(7)));
    layer0_outputs(7636) <= inputs(113);
    layer0_outputs(7637) <= (inputs(43)) xor (inputs(46));
    layer0_outputs(7638) <= inputs(229);
    layer0_outputs(7639) <= inputs(33);
    layer0_outputs(7640) <= inputs(216);
    layer0_outputs(7641) <= (inputs(45)) xor (inputs(125));
    layer0_outputs(7642) <= (inputs(154)) xor (inputs(158));
    layer0_outputs(7643) <= not((inputs(154)) xor (inputs(72)));
    layer0_outputs(7644) <= (inputs(32)) or (inputs(164));
    layer0_outputs(7645) <= inputs(14);
    layer0_outputs(7646) <= (inputs(220)) or (inputs(197));
    layer0_outputs(7647) <= (inputs(189)) or (inputs(2));
    layer0_outputs(7648) <= not(inputs(34));
    layer0_outputs(7649) <= not((inputs(82)) or (inputs(147)));
    layer0_outputs(7650) <= (inputs(35)) and (inputs(142));
    layer0_outputs(7651) <= not((inputs(208)) or (inputs(223)));
    layer0_outputs(7652) <= (inputs(21)) or (inputs(219));
    layer0_outputs(7653) <= inputs(168);
    layer0_outputs(7654) <= (inputs(69)) and not (inputs(243));
    layer0_outputs(7655) <= inputs(147);
    layer0_outputs(7656) <= inputs(162);
    layer0_outputs(7657) <= not((inputs(181)) or (inputs(141)));
    layer0_outputs(7658) <= (inputs(75)) or (inputs(222));
    layer0_outputs(7659) <= not((inputs(23)) and (inputs(134)));
    layer0_outputs(7660) <= inputs(211);
    layer0_outputs(7661) <= not(inputs(25));
    layer0_outputs(7662) <= not((inputs(91)) xor (inputs(19)));
    layer0_outputs(7663) <= not((inputs(220)) xor (inputs(253)));
    layer0_outputs(7664) <= not(inputs(126));
    layer0_outputs(7665) <= not((inputs(160)) xor (inputs(86)));
    layer0_outputs(7666) <= inputs(212);
    layer0_outputs(7667) <= not(inputs(151));
    layer0_outputs(7668) <= inputs(48);
    layer0_outputs(7669) <= inputs(165);
    layer0_outputs(7670) <= not(inputs(186)) or (inputs(246));
    layer0_outputs(7671) <= (inputs(42)) and not (inputs(224));
    layer0_outputs(7672) <= (inputs(132)) or (inputs(114));
    layer0_outputs(7673) <= (inputs(77)) or (inputs(108));
    layer0_outputs(7674) <= (inputs(24)) and not (inputs(5));
    layer0_outputs(7675) <= inputs(202);
    layer0_outputs(7676) <= (inputs(60)) and not (inputs(112));
    layer0_outputs(7677) <= '1';
    layer0_outputs(7678) <= not((inputs(193)) xor (inputs(238)));
    layer0_outputs(7679) <= (inputs(202)) or (inputs(159));
    layer0_outputs(7680) <= (inputs(82)) or (inputs(240));
    layer0_outputs(7681) <= not((inputs(241)) or (inputs(247)));
    layer0_outputs(7682) <= inputs(24);
    layer0_outputs(7683) <= not(inputs(186)) or (inputs(16));
    layer0_outputs(7684) <= inputs(7);
    layer0_outputs(7685) <= (inputs(180)) or (inputs(168));
    layer0_outputs(7686) <= (inputs(225)) or (inputs(145));
    layer0_outputs(7687) <= not((inputs(206)) or (inputs(50)));
    layer0_outputs(7688) <= (inputs(42)) xor (inputs(10));
    layer0_outputs(7689) <= (inputs(172)) or (inputs(187));
    layer0_outputs(7690) <= inputs(225);
    layer0_outputs(7691) <= not(inputs(211)) or (inputs(16));
    layer0_outputs(7692) <= not((inputs(24)) or (inputs(247)));
    layer0_outputs(7693) <= inputs(119);
    layer0_outputs(7694) <= not(inputs(27));
    layer0_outputs(7695) <= not(inputs(189)) or (inputs(33));
    layer0_outputs(7696) <= inputs(160);
    layer0_outputs(7697) <= not(inputs(85)) or (inputs(226));
    layer0_outputs(7698) <= not((inputs(224)) or (inputs(135)));
    layer0_outputs(7699) <= (inputs(91)) and not (inputs(160));
    layer0_outputs(7700) <= not((inputs(101)) xor (inputs(99)));
    layer0_outputs(7701) <= not(inputs(241)) or (inputs(66));
    layer0_outputs(7702) <= (inputs(21)) and not (inputs(44));
    layer0_outputs(7703) <= not(inputs(252));
    layer0_outputs(7704) <= (inputs(196)) or (inputs(37));
    layer0_outputs(7705) <= not(inputs(183));
    layer0_outputs(7706) <= inputs(234);
    layer0_outputs(7707) <= not(inputs(229));
    layer0_outputs(7708) <= (inputs(70)) or (inputs(183));
    layer0_outputs(7709) <= not(inputs(106)) or (inputs(128));
    layer0_outputs(7710) <= (inputs(126)) and not (inputs(106));
    layer0_outputs(7711) <= inputs(245);
    layer0_outputs(7712) <= not(inputs(34));
    layer0_outputs(7713) <= not((inputs(94)) or (inputs(8)));
    layer0_outputs(7714) <= '1';
    layer0_outputs(7715) <= not(inputs(219));
    layer0_outputs(7716) <= (inputs(101)) or (inputs(228));
    layer0_outputs(7717) <= inputs(7);
    layer0_outputs(7718) <= (inputs(57)) and not (inputs(252));
    layer0_outputs(7719) <= not((inputs(237)) and (inputs(156)));
    layer0_outputs(7720) <= not(inputs(241));
    layer0_outputs(7721) <= (inputs(177)) xor (inputs(246));
    layer0_outputs(7722) <= inputs(86);
    layer0_outputs(7723) <= not(inputs(216));
    layer0_outputs(7724) <= (inputs(39)) or (inputs(223));
    layer0_outputs(7725) <= not(inputs(2));
    layer0_outputs(7726) <= (inputs(171)) xor (inputs(202));
    layer0_outputs(7727) <= (inputs(124)) xor (inputs(63));
    layer0_outputs(7728) <= inputs(235);
    layer0_outputs(7729) <= not(inputs(86)) or (inputs(93));
    layer0_outputs(7730) <= inputs(55);
    layer0_outputs(7731) <= (inputs(224)) or (inputs(236));
    layer0_outputs(7732) <= (inputs(191)) or (inputs(104));
    layer0_outputs(7733) <= not(inputs(147)) or (inputs(50));
    layer0_outputs(7734) <= not((inputs(19)) or (inputs(123)));
    layer0_outputs(7735) <= not((inputs(40)) xor (inputs(111)));
    layer0_outputs(7736) <= (inputs(190)) or (inputs(176));
    layer0_outputs(7737) <= not((inputs(125)) or (inputs(137)));
    layer0_outputs(7738) <= not(inputs(101)) or (inputs(185));
    layer0_outputs(7739) <= not((inputs(71)) or (inputs(159)));
    layer0_outputs(7740) <= (inputs(135)) and not (inputs(26));
    layer0_outputs(7741) <= not(inputs(111)) or (inputs(2));
    layer0_outputs(7742) <= (inputs(161)) and (inputs(233));
    layer0_outputs(7743) <= (inputs(83)) or (inputs(121));
    layer0_outputs(7744) <= not(inputs(53)) or (inputs(27));
    layer0_outputs(7745) <= not(inputs(100));
    layer0_outputs(7746) <= (inputs(84)) and not (inputs(205));
    layer0_outputs(7747) <= not(inputs(64)) or (inputs(249));
    layer0_outputs(7748) <= inputs(205);
    layer0_outputs(7749) <= not((inputs(146)) and (inputs(130)));
    layer0_outputs(7750) <= not((inputs(124)) xor (inputs(36)));
    layer0_outputs(7751) <= (inputs(178)) xor (inputs(116));
    layer0_outputs(7752) <= (inputs(16)) and not (inputs(16));
    layer0_outputs(7753) <= inputs(161);
    layer0_outputs(7754) <= (inputs(13)) or (inputs(236));
    layer0_outputs(7755) <= not(inputs(68));
    layer0_outputs(7756) <= (inputs(108)) xor (inputs(50));
    layer0_outputs(7757) <= (inputs(184)) and not (inputs(116));
    layer0_outputs(7758) <= not(inputs(123)) or (inputs(195));
    layer0_outputs(7759) <= (inputs(196)) and not (inputs(123));
    layer0_outputs(7760) <= not(inputs(65)) or (inputs(141));
    layer0_outputs(7761) <= (inputs(172)) and not (inputs(94));
    layer0_outputs(7762) <= (inputs(74)) and not (inputs(158));
    layer0_outputs(7763) <= inputs(73);
    layer0_outputs(7764) <= not(inputs(42));
    layer0_outputs(7765) <= inputs(78);
    layer0_outputs(7766) <= inputs(25);
    layer0_outputs(7767) <= (inputs(170)) xor (inputs(106));
    layer0_outputs(7768) <= (inputs(78)) and not (inputs(166));
    layer0_outputs(7769) <= not(inputs(228));
    layer0_outputs(7770) <= (inputs(234)) xor (inputs(61));
    layer0_outputs(7771) <= not(inputs(229)) or (inputs(66));
    layer0_outputs(7772) <= not((inputs(54)) or (inputs(193)));
    layer0_outputs(7773) <= inputs(83);
    layer0_outputs(7774) <= inputs(102);
    layer0_outputs(7775) <= (inputs(134)) or (inputs(89));
    layer0_outputs(7776) <= not(inputs(91));
    layer0_outputs(7777) <= not(inputs(246));
    layer0_outputs(7778) <= (inputs(43)) and not (inputs(204));
    layer0_outputs(7779) <= (inputs(9)) and not (inputs(144));
    layer0_outputs(7780) <= inputs(161);
    layer0_outputs(7781) <= inputs(132);
    layer0_outputs(7782) <= (inputs(174)) or (inputs(204));
    layer0_outputs(7783) <= not(inputs(92)) or (inputs(209));
    layer0_outputs(7784) <= (inputs(143)) xor (inputs(10));
    layer0_outputs(7785) <= not(inputs(146));
    layer0_outputs(7786) <= (inputs(71)) xor (inputs(21));
    layer0_outputs(7787) <= (inputs(253)) xor (inputs(18));
    layer0_outputs(7788) <= not(inputs(76));
    layer0_outputs(7789) <= not((inputs(148)) or (inputs(93)));
    layer0_outputs(7790) <= (inputs(27)) and not (inputs(166));
    layer0_outputs(7791) <= not(inputs(24));
    layer0_outputs(7792) <= inputs(197);
    layer0_outputs(7793) <= (inputs(2)) or (inputs(223));
    layer0_outputs(7794) <= not((inputs(142)) or (inputs(84)));
    layer0_outputs(7795) <= inputs(30);
    layer0_outputs(7796) <= (inputs(64)) and (inputs(49));
    layer0_outputs(7797) <= '0';
    layer0_outputs(7798) <= (inputs(204)) and not (inputs(40));
    layer0_outputs(7799) <= (inputs(235)) xor (inputs(150));
    layer0_outputs(7800) <= inputs(29);
    layer0_outputs(7801) <= inputs(57);
    layer0_outputs(7802) <= not(inputs(120));
    layer0_outputs(7803) <= inputs(123);
    layer0_outputs(7804) <= not(inputs(38));
    layer0_outputs(7805) <= not((inputs(212)) or (inputs(238)));
    layer0_outputs(7806) <= not(inputs(193));
    layer0_outputs(7807) <= (inputs(44)) and not (inputs(176));
    layer0_outputs(7808) <= not(inputs(60)) or (inputs(118));
    layer0_outputs(7809) <= inputs(119);
    layer0_outputs(7810) <= not((inputs(67)) or (inputs(218)));
    layer0_outputs(7811) <= inputs(70);
    layer0_outputs(7812) <= inputs(29);
    layer0_outputs(7813) <= not((inputs(179)) or (inputs(170)));
    layer0_outputs(7814) <= (inputs(162)) or (inputs(24));
    layer0_outputs(7815) <= not(inputs(210));
    layer0_outputs(7816) <= inputs(91);
    layer0_outputs(7817) <= (inputs(71)) xor (inputs(218));
    layer0_outputs(7818) <= not(inputs(133));
    layer0_outputs(7819) <= (inputs(54)) xor (inputs(252));
    layer0_outputs(7820) <= (inputs(68)) xor (inputs(51));
    layer0_outputs(7821) <= not((inputs(217)) or (inputs(208)));
    layer0_outputs(7822) <= inputs(194);
    layer0_outputs(7823) <= (inputs(188)) or (inputs(86));
    layer0_outputs(7824) <= (inputs(182)) or (inputs(83));
    layer0_outputs(7825) <= (inputs(54)) and not (inputs(29));
    layer0_outputs(7826) <= not((inputs(35)) xor (inputs(192)));
    layer0_outputs(7827) <= not(inputs(160));
    layer0_outputs(7828) <= not(inputs(249));
    layer0_outputs(7829) <= (inputs(61)) and not (inputs(132));
    layer0_outputs(7830) <= not(inputs(241));
    layer0_outputs(7831) <= not(inputs(100));
    layer0_outputs(7832) <= not((inputs(171)) and (inputs(178)));
    layer0_outputs(7833) <= inputs(250);
    layer0_outputs(7834) <= (inputs(239)) or (inputs(176));
    layer0_outputs(7835) <= not((inputs(231)) or (inputs(94)));
    layer0_outputs(7836) <= not(inputs(114));
    layer0_outputs(7837) <= not(inputs(179));
    layer0_outputs(7838) <= '0';
    layer0_outputs(7839) <= not(inputs(56));
    layer0_outputs(7840) <= not(inputs(227));
    layer0_outputs(7841) <= inputs(7);
    layer0_outputs(7842) <= not((inputs(26)) xor (inputs(207)));
    layer0_outputs(7843) <= (inputs(96)) and (inputs(224));
    layer0_outputs(7844) <= (inputs(42)) or (inputs(214));
    layer0_outputs(7845) <= (inputs(36)) or (inputs(126));
    layer0_outputs(7846) <= not((inputs(169)) xor (inputs(149)));
    layer0_outputs(7847) <= not((inputs(222)) xor (inputs(62)));
    layer0_outputs(7848) <= not((inputs(23)) or (inputs(6)));
    layer0_outputs(7849) <= not(inputs(28)) or (inputs(192));
    layer0_outputs(7850) <= (inputs(141)) and not (inputs(222));
    layer0_outputs(7851) <= (inputs(127)) xor (inputs(27));
    layer0_outputs(7852) <= (inputs(143)) or (inputs(3));
    layer0_outputs(7853) <= (inputs(202)) xor (inputs(213));
    layer0_outputs(7854) <= not((inputs(96)) xor (inputs(130)));
    layer0_outputs(7855) <= not(inputs(119));
    layer0_outputs(7856) <= (inputs(65)) or (inputs(68));
    layer0_outputs(7857) <= (inputs(68)) or (inputs(125));
    layer0_outputs(7858) <= not((inputs(65)) or (inputs(238)));
    layer0_outputs(7859) <= not((inputs(23)) or (inputs(225)));
    layer0_outputs(7860) <= (inputs(155)) or (inputs(18));
    layer0_outputs(7861) <= (inputs(204)) or (inputs(174));
    layer0_outputs(7862) <= '0';
    layer0_outputs(7863) <= not(inputs(80));
    layer0_outputs(7864) <= (inputs(101)) and (inputs(198));
    layer0_outputs(7865) <= (inputs(121)) and (inputs(212));
    layer0_outputs(7866) <= (inputs(4)) and not (inputs(176));
    layer0_outputs(7867) <= not(inputs(140));
    layer0_outputs(7868) <= not((inputs(110)) or (inputs(3)));
    layer0_outputs(7869) <= not(inputs(9));
    layer0_outputs(7870) <= '1';
    layer0_outputs(7871) <= not(inputs(136)) or (inputs(241));
    layer0_outputs(7872) <= inputs(74);
    layer0_outputs(7873) <= (inputs(244)) and not (inputs(35));
    layer0_outputs(7874) <= not(inputs(149));
    layer0_outputs(7875) <= not(inputs(8)) or (inputs(83));
    layer0_outputs(7876) <= inputs(105);
    layer0_outputs(7877) <= '0';
    layer0_outputs(7878) <= not(inputs(41));
    layer0_outputs(7879) <= (inputs(117)) or (inputs(87));
    layer0_outputs(7880) <= '0';
    layer0_outputs(7881) <= inputs(0);
    layer0_outputs(7882) <= (inputs(204)) and not (inputs(127));
    layer0_outputs(7883) <= not(inputs(68)) or (inputs(18));
    layer0_outputs(7884) <= not((inputs(103)) xor (inputs(255)));
    layer0_outputs(7885) <= not(inputs(166));
    layer0_outputs(7886) <= not((inputs(196)) or (inputs(53)));
    layer0_outputs(7887) <= (inputs(248)) or (inputs(192));
    layer0_outputs(7888) <= inputs(76);
    layer0_outputs(7889) <= (inputs(45)) or (inputs(88));
    layer0_outputs(7890) <= '1';
    layer0_outputs(7891) <= (inputs(42)) and not (inputs(162));
    layer0_outputs(7892) <= not(inputs(22)) or (inputs(81));
    layer0_outputs(7893) <= (inputs(180)) or (inputs(23));
    layer0_outputs(7894) <= not((inputs(232)) or (inputs(211)));
    layer0_outputs(7895) <= (inputs(59)) or (inputs(109));
    layer0_outputs(7896) <= not(inputs(113));
    layer0_outputs(7897) <= not((inputs(190)) xor (inputs(211)));
    layer0_outputs(7898) <= not((inputs(63)) xor (inputs(18)));
    layer0_outputs(7899) <= (inputs(249)) or (inputs(100));
    layer0_outputs(7900) <= inputs(167);
    layer0_outputs(7901) <= not((inputs(1)) or (inputs(55)));
    layer0_outputs(7902) <= not(inputs(113));
    layer0_outputs(7903) <= not((inputs(129)) or (inputs(203)));
    layer0_outputs(7904) <= not(inputs(199)) or (inputs(13));
    layer0_outputs(7905) <= inputs(248);
    layer0_outputs(7906) <= (inputs(187)) or (inputs(154));
    layer0_outputs(7907) <= not((inputs(54)) and (inputs(112)));
    layer0_outputs(7908) <= inputs(37);
    layer0_outputs(7909) <= not((inputs(41)) or (inputs(35)));
    layer0_outputs(7910) <= not((inputs(102)) or (inputs(97)));
    layer0_outputs(7911) <= not(inputs(134));
    layer0_outputs(7912) <= not((inputs(14)) or (inputs(151)));
    layer0_outputs(7913) <= not((inputs(177)) or (inputs(245)));
    layer0_outputs(7914) <= not((inputs(11)) xor (inputs(98)));
    layer0_outputs(7915) <= not(inputs(34)) or (inputs(239));
    layer0_outputs(7916) <= inputs(30);
    layer0_outputs(7917) <= not(inputs(224)) or (inputs(125));
    layer0_outputs(7918) <= not((inputs(71)) xor (inputs(101)));
    layer0_outputs(7919) <= inputs(86);
    layer0_outputs(7920) <= (inputs(181)) and not (inputs(108));
    layer0_outputs(7921) <= not(inputs(164));
    layer0_outputs(7922) <= (inputs(26)) and not (inputs(163));
    layer0_outputs(7923) <= (inputs(185)) and not (inputs(52));
    layer0_outputs(7924) <= not(inputs(23));
    layer0_outputs(7925) <= not(inputs(9));
    layer0_outputs(7926) <= not(inputs(146)) or (inputs(138));
    layer0_outputs(7927) <= (inputs(64)) and (inputs(208));
    layer0_outputs(7928) <= not((inputs(115)) and (inputs(213)));
    layer0_outputs(7929) <= inputs(203);
    layer0_outputs(7930) <= not(inputs(142));
    layer0_outputs(7931) <= not((inputs(158)) or (inputs(63)));
    layer0_outputs(7932) <= not((inputs(38)) xor (inputs(72)));
    layer0_outputs(7933) <= inputs(10);
    layer0_outputs(7934) <= not((inputs(240)) and (inputs(236)));
    layer0_outputs(7935) <= (inputs(88)) and not (inputs(49));
    layer0_outputs(7936) <= (inputs(79)) or (inputs(218));
    layer0_outputs(7937) <= inputs(123);
    layer0_outputs(7938) <= not(inputs(223));
    layer0_outputs(7939) <= (inputs(197)) or (inputs(144));
    layer0_outputs(7940) <= not(inputs(25));
    layer0_outputs(7941) <= not((inputs(151)) or (inputs(1)));
    layer0_outputs(7942) <= not(inputs(178));
    layer0_outputs(7943) <= (inputs(159)) or (inputs(161));
    layer0_outputs(7944) <= (inputs(224)) or (inputs(250));
    layer0_outputs(7945) <= not(inputs(91));
    layer0_outputs(7946) <= (inputs(231)) and not (inputs(220));
    layer0_outputs(7947) <= not(inputs(167));
    layer0_outputs(7948) <= not(inputs(48));
    layer0_outputs(7949) <= (inputs(229)) and not (inputs(136));
    layer0_outputs(7950) <= (inputs(205)) xor (inputs(10));
    layer0_outputs(7951) <= not((inputs(144)) or (inputs(49)));
    layer0_outputs(7952) <= (inputs(74)) or (inputs(110));
    layer0_outputs(7953) <= inputs(56);
    layer0_outputs(7954) <= inputs(114);
    layer0_outputs(7955) <= not(inputs(164));
    layer0_outputs(7956) <= inputs(211);
    layer0_outputs(7957) <= not(inputs(183)) or (inputs(15));
    layer0_outputs(7958) <= not((inputs(228)) or (inputs(148)));
    layer0_outputs(7959) <= not((inputs(251)) or (inputs(85)));
    layer0_outputs(7960) <= (inputs(170)) and not (inputs(32));
    layer0_outputs(7961) <= (inputs(148)) and not (inputs(178));
    layer0_outputs(7962) <= inputs(173);
    layer0_outputs(7963) <= (inputs(36)) and not (inputs(148));
    layer0_outputs(7964) <= not(inputs(217));
    layer0_outputs(7965) <= inputs(39);
    layer0_outputs(7966) <= (inputs(1)) xor (inputs(222));
    layer0_outputs(7967) <= inputs(209);
    layer0_outputs(7968) <= not(inputs(83));
    layer0_outputs(7969) <= not((inputs(50)) and (inputs(64)));
    layer0_outputs(7970) <= not((inputs(198)) xor (inputs(249)));
    layer0_outputs(7971) <= not(inputs(222));
    layer0_outputs(7972) <= not((inputs(171)) xor (inputs(1)));
    layer0_outputs(7973) <= (inputs(193)) and not (inputs(81));
    layer0_outputs(7974) <= not(inputs(22));
    layer0_outputs(7975) <= (inputs(248)) and not (inputs(251));
    layer0_outputs(7976) <= not(inputs(218));
    layer0_outputs(7977) <= not(inputs(139));
    layer0_outputs(7978) <= inputs(79);
    layer0_outputs(7979) <= (inputs(20)) xor (inputs(176));
    layer0_outputs(7980) <= not(inputs(179));
    layer0_outputs(7981) <= (inputs(161)) or (inputs(215));
    layer0_outputs(7982) <= (inputs(100)) or (inputs(174));
    layer0_outputs(7983) <= inputs(229);
    layer0_outputs(7984) <= inputs(181);
    layer0_outputs(7985) <= not(inputs(150));
    layer0_outputs(7986) <= (inputs(193)) and not (inputs(245));
    layer0_outputs(7987) <= (inputs(172)) or (inputs(33));
    layer0_outputs(7988) <= (inputs(144)) and not (inputs(62));
    layer0_outputs(7989) <= '1';
    layer0_outputs(7990) <= (inputs(16)) xor (inputs(248));
    layer0_outputs(7991) <= not((inputs(10)) or (inputs(141)));
    layer0_outputs(7992) <= not((inputs(157)) or (inputs(101)));
    layer0_outputs(7993) <= (inputs(236)) and not (inputs(249));
    layer0_outputs(7994) <= (inputs(171)) or (inputs(98));
    layer0_outputs(7995) <= inputs(91);
    layer0_outputs(7996) <= (inputs(115)) and not (inputs(202));
    layer0_outputs(7997) <= not(inputs(195));
    layer0_outputs(7998) <= not((inputs(17)) or (inputs(45)));
    layer0_outputs(7999) <= not((inputs(126)) xor (inputs(48)));
    layer0_outputs(8000) <= inputs(30);
    layer0_outputs(8001) <= not(inputs(169)) or (inputs(15));
    layer0_outputs(8002) <= not(inputs(49)) or (inputs(1));
    layer0_outputs(8003) <= not(inputs(186)) or (inputs(192));
    layer0_outputs(8004) <= (inputs(62)) or (inputs(33));
    layer0_outputs(8005) <= not(inputs(59));
    layer0_outputs(8006) <= not(inputs(16));
    layer0_outputs(8007) <= (inputs(88)) and not (inputs(147));
    layer0_outputs(8008) <= not(inputs(41));
    layer0_outputs(8009) <= (inputs(255)) or (inputs(147));
    layer0_outputs(8010) <= (inputs(184)) and not (inputs(78));
    layer0_outputs(8011) <= (inputs(245)) or (inputs(81));
    layer0_outputs(8012) <= not((inputs(125)) xor (inputs(86)));
    layer0_outputs(8013) <= not(inputs(68)) or (inputs(166));
    layer0_outputs(8014) <= (inputs(173)) and not (inputs(16));
    layer0_outputs(8015) <= (inputs(220)) and not (inputs(91));
    layer0_outputs(8016) <= not((inputs(194)) xor (inputs(123)));
    layer0_outputs(8017) <= not((inputs(61)) or (inputs(95)));
    layer0_outputs(8018) <= (inputs(75)) and (inputs(79));
    layer0_outputs(8019) <= (inputs(248)) or (inputs(208));
    layer0_outputs(8020) <= not((inputs(80)) xor (inputs(6)));
    layer0_outputs(8021) <= not((inputs(102)) xor (inputs(148)));
    layer0_outputs(8022) <= inputs(188);
    layer0_outputs(8023) <= not(inputs(87)) or (inputs(64));
    layer0_outputs(8024) <= (inputs(208)) and not (inputs(0));
    layer0_outputs(8025) <= not((inputs(190)) or (inputs(95)));
    layer0_outputs(8026) <= not(inputs(98));
    layer0_outputs(8027) <= not(inputs(107)) or (inputs(114));
    layer0_outputs(8028) <= not((inputs(206)) xor (inputs(175)));
    layer0_outputs(8029) <= not((inputs(196)) or (inputs(33)));
    layer0_outputs(8030) <= not(inputs(24));
    layer0_outputs(8031) <= (inputs(179)) and not (inputs(17));
    layer0_outputs(8032) <= not((inputs(227)) xor (inputs(1)));
    layer0_outputs(8033) <= not((inputs(18)) xor (inputs(195)));
    layer0_outputs(8034) <= (inputs(199)) xor (inputs(181));
    layer0_outputs(8035) <= not((inputs(114)) or (inputs(91)));
    layer0_outputs(8036) <= inputs(127);
    layer0_outputs(8037) <= not((inputs(159)) xor (inputs(101)));
    layer0_outputs(8038) <= (inputs(0)) and not (inputs(255));
    layer0_outputs(8039) <= (inputs(36)) xor (inputs(128));
    layer0_outputs(8040) <= inputs(246);
    layer0_outputs(8041) <= not((inputs(126)) or (inputs(236)));
    layer0_outputs(8042) <= not((inputs(207)) or (inputs(227)));
    layer0_outputs(8043) <= inputs(25);
    layer0_outputs(8044) <= not(inputs(79));
    layer0_outputs(8045) <= not(inputs(45)) or (inputs(55));
    layer0_outputs(8046) <= not((inputs(157)) xor (inputs(115)));
    layer0_outputs(8047) <= '0';
    layer0_outputs(8048) <= not((inputs(251)) or (inputs(245)));
    layer0_outputs(8049) <= (inputs(234)) and not (inputs(165));
    layer0_outputs(8050) <= (inputs(23)) xor (inputs(66));
    layer0_outputs(8051) <= not(inputs(173)) or (inputs(178));
    layer0_outputs(8052) <= not(inputs(221));
    layer0_outputs(8053) <= inputs(121);
    layer0_outputs(8054) <= not(inputs(59));
    layer0_outputs(8055) <= not(inputs(82));
    layer0_outputs(8056) <= (inputs(157)) xor (inputs(36));
    layer0_outputs(8057) <= inputs(180);
    layer0_outputs(8058) <= (inputs(204)) xor (inputs(225));
    layer0_outputs(8059) <= '0';
    layer0_outputs(8060) <= not(inputs(130)) or (inputs(222));
    layer0_outputs(8061) <= not(inputs(142));
    layer0_outputs(8062) <= not(inputs(69));
    layer0_outputs(8063) <= inputs(164);
    layer0_outputs(8064) <= (inputs(194)) xor (inputs(235));
    layer0_outputs(8065) <= not(inputs(90));
    layer0_outputs(8066) <= (inputs(149)) xor (inputs(189));
    layer0_outputs(8067) <= inputs(82);
    layer0_outputs(8068) <= (inputs(28)) and (inputs(69));
    layer0_outputs(8069) <= not(inputs(41));
    layer0_outputs(8070) <= not(inputs(222));
    layer0_outputs(8071) <= not(inputs(201));
    layer0_outputs(8072) <= (inputs(251)) and not (inputs(241));
    layer0_outputs(8073) <= (inputs(65)) or (inputs(83));
    layer0_outputs(8074) <= not((inputs(143)) and (inputs(60)));
    layer0_outputs(8075) <= (inputs(55)) and not (inputs(34));
    layer0_outputs(8076) <= (inputs(196)) or (inputs(248));
    layer0_outputs(8077) <= not(inputs(220)) or (inputs(87));
    layer0_outputs(8078) <= inputs(10);
    layer0_outputs(8079) <= not((inputs(13)) or (inputs(144)));
    layer0_outputs(8080) <= inputs(67);
    layer0_outputs(8081) <= not(inputs(67)) or (inputs(73));
    layer0_outputs(8082) <= not((inputs(197)) or (inputs(7)));
    layer0_outputs(8083) <= not(inputs(206)) or (inputs(112));
    layer0_outputs(8084) <= not((inputs(255)) or (inputs(143)));
    layer0_outputs(8085) <= (inputs(123)) and not (inputs(178));
    layer0_outputs(8086) <= not((inputs(246)) xor (inputs(169)));
    layer0_outputs(8087) <= not(inputs(129)) or (inputs(102));
    layer0_outputs(8088) <= not(inputs(90));
    layer0_outputs(8089) <= not(inputs(214)) or (inputs(123));
    layer0_outputs(8090) <= (inputs(123)) or (inputs(20));
    layer0_outputs(8091) <= not(inputs(57)) or (inputs(188));
    layer0_outputs(8092) <= inputs(142);
    layer0_outputs(8093) <= inputs(232);
    layer0_outputs(8094) <= (inputs(176)) xor (inputs(171));
    layer0_outputs(8095) <= (inputs(63)) or (inputs(48));
    layer0_outputs(8096) <= not(inputs(166));
    layer0_outputs(8097) <= not((inputs(52)) or (inputs(206)));
    layer0_outputs(8098) <= (inputs(190)) and (inputs(45));
    layer0_outputs(8099) <= (inputs(103)) xor (inputs(73));
    layer0_outputs(8100) <= not((inputs(181)) or (inputs(65)));
    layer0_outputs(8101) <= (inputs(229)) and not (inputs(95));
    layer0_outputs(8102) <= inputs(40);
    layer0_outputs(8103) <= not(inputs(35)) or (inputs(83));
    layer0_outputs(8104) <= not((inputs(193)) or (inputs(2)));
    layer0_outputs(8105) <= not(inputs(74));
    layer0_outputs(8106) <= not(inputs(158));
    layer0_outputs(8107) <= not((inputs(104)) or (inputs(174)));
    layer0_outputs(8108) <= not(inputs(162));
    layer0_outputs(8109) <= not(inputs(24)) or (inputs(228));
    layer0_outputs(8110) <= not((inputs(125)) xor (inputs(240)));
    layer0_outputs(8111) <= not(inputs(133)) or (inputs(31));
    layer0_outputs(8112) <= not(inputs(223)) or (inputs(200));
    layer0_outputs(8113) <= not(inputs(104)) or (inputs(167));
    layer0_outputs(8114) <= (inputs(122)) xor (inputs(239));
    layer0_outputs(8115) <= not((inputs(137)) and (inputs(209)));
    layer0_outputs(8116) <= (inputs(117)) and not (inputs(147));
    layer0_outputs(8117) <= (inputs(40)) or (inputs(23));
    layer0_outputs(8118) <= not(inputs(156));
    layer0_outputs(8119) <= not(inputs(163)) or (inputs(83));
    layer0_outputs(8120) <= (inputs(169)) xor (inputs(50));
    layer0_outputs(8121) <= (inputs(215)) or (inputs(237));
    layer0_outputs(8122) <= not(inputs(87)) or (inputs(34));
    layer0_outputs(8123) <= not(inputs(1));
    layer0_outputs(8124) <= not((inputs(163)) xor (inputs(170)));
    layer0_outputs(8125) <= not((inputs(121)) xor (inputs(101)));
    layer0_outputs(8126) <= inputs(112);
    layer0_outputs(8127) <= not((inputs(104)) xor (inputs(148)));
    layer0_outputs(8128) <= inputs(177);
    layer0_outputs(8129) <= inputs(78);
    layer0_outputs(8130) <= (inputs(69)) or (inputs(208));
    layer0_outputs(8131) <= not(inputs(176)) or (inputs(35));
    layer0_outputs(8132) <= inputs(136);
    layer0_outputs(8133) <= not((inputs(138)) or (inputs(165)));
    layer0_outputs(8134) <= (inputs(155)) xor (inputs(238));
    layer0_outputs(8135) <= not(inputs(206));
    layer0_outputs(8136) <= (inputs(240)) xor (inputs(21));
    layer0_outputs(8137) <= not(inputs(123));
    layer0_outputs(8138) <= '1';
    layer0_outputs(8139) <= not((inputs(71)) xor (inputs(227)));
    layer0_outputs(8140) <= (inputs(231)) and not (inputs(140));
    layer0_outputs(8141) <= inputs(22);
    layer0_outputs(8142) <= not(inputs(151));
    layer0_outputs(8143) <= (inputs(0)) xor (inputs(246));
    layer0_outputs(8144) <= not((inputs(19)) xor (inputs(72)));
    layer0_outputs(8145) <= inputs(212);
    layer0_outputs(8146) <= (inputs(124)) and not (inputs(12));
    layer0_outputs(8147) <= (inputs(224)) or (inputs(137));
    layer0_outputs(8148) <= not(inputs(68)) or (inputs(106));
    layer0_outputs(8149) <= (inputs(95)) or (inputs(61));
    layer0_outputs(8150) <= (inputs(2)) or (inputs(35));
    layer0_outputs(8151) <= (inputs(29)) or (inputs(188));
    layer0_outputs(8152) <= not(inputs(111));
    layer0_outputs(8153) <= inputs(250);
    layer0_outputs(8154) <= (inputs(85)) or (inputs(194));
    layer0_outputs(8155) <= not((inputs(51)) or (inputs(112)));
    layer0_outputs(8156) <= not(inputs(90)) or (inputs(239));
    layer0_outputs(8157) <= not((inputs(64)) or (inputs(214)));
    layer0_outputs(8158) <= (inputs(192)) and not (inputs(251));
    layer0_outputs(8159) <= inputs(110);
    layer0_outputs(8160) <= (inputs(203)) xor (inputs(171));
    layer0_outputs(8161) <= (inputs(178)) and not (inputs(60));
    layer0_outputs(8162) <= not((inputs(156)) xor (inputs(157)));
    layer0_outputs(8163) <= not((inputs(67)) xor (inputs(69)));
    layer0_outputs(8164) <= inputs(206);
    layer0_outputs(8165) <= (inputs(189)) and not (inputs(254));
    layer0_outputs(8166) <= not(inputs(142));
    layer0_outputs(8167) <= (inputs(7)) and not (inputs(225));
    layer0_outputs(8168) <= not((inputs(52)) xor (inputs(33)));
    layer0_outputs(8169) <= inputs(110);
    layer0_outputs(8170) <= not((inputs(140)) and (inputs(131)));
    layer0_outputs(8171) <= not(inputs(119));
    layer0_outputs(8172) <= (inputs(218)) and not (inputs(25));
    layer0_outputs(8173) <= not(inputs(22));
    layer0_outputs(8174) <= not((inputs(152)) or (inputs(177)));
    layer0_outputs(8175) <= not(inputs(44));
    layer0_outputs(8176) <= not(inputs(14));
    layer0_outputs(8177) <= not(inputs(234)) or (inputs(78));
    layer0_outputs(8178) <= not((inputs(234)) xor (inputs(62)));
    layer0_outputs(8179) <= (inputs(197)) and not (inputs(116));
    layer0_outputs(8180) <= not(inputs(230)) or (inputs(156));
    layer0_outputs(8181) <= (inputs(29)) and not (inputs(32));
    layer0_outputs(8182) <= inputs(62);
    layer0_outputs(8183) <= not(inputs(129)) or (inputs(223));
    layer0_outputs(8184) <= not(inputs(243)) or (inputs(14));
    layer0_outputs(8185) <= (inputs(126)) or (inputs(242));
    layer0_outputs(8186) <= not(inputs(41)) or (inputs(127));
    layer0_outputs(8187) <= (inputs(63)) xor (inputs(248));
    layer0_outputs(8188) <= not((inputs(195)) or (inputs(239)));
    layer0_outputs(8189) <= not((inputs(7)) xor (inputs(74)));
    layer0_outputs(8190) <= not(inputs(137)) or (inputs(28));
    layer0_outputs(8191) <= (inputs(96)) xor (inputs(23));
    layer0_outputs(8192) <= (inputs(234)) or (inputs(194));
    layer0_outputs(8193) <= (inputs(248)) or (inputs(65));
    layer0_outputs(8194) <= not((inputs(58)) or (inputs(59)));
    layer0_outputs(8195) <= (inputs(86)) and (inputs(176));
    layer0_outputs(8196) <= not((inputs(179)) or (inputs(176)));
    layer0_outputs(8197) <= inputs(0);
    layer0_outputs(8198) <= (inputs(202)) or (inputs(241));
    layer0_outputs(8199) <= (inputs(247)) and not (inputs(22));
    layer0_outputs(8200) <= (inputs(99)) and (inputs(83));
    layer0_outputs(8201) <= not(inputs(204)) or (inputs(225));
    layer0_outputs(8202) <= inputs(118);
    layer0_outputs(8203) <= not(inputs(165)) or (inputs(255));
    layer0_outputs(8204) <= (inputs(200)) and (inputs(197));
    layer0_outputs(8205) <= not(inputs(213)) or (inputs(206));
    layer0_outputs(8206) <= (inputs(159)) xor (inputs(214));
    layer0_outputs(8207) <= (inputs(182)) and not (inputs(8));
    layer0_outputs(8208) <= '1';
    layer0_outputs(8209) <= (inputs(131)) or (inputs(12));
    layer0_outputs(8210) <= not(inputs(119)) or (inputs(0));
    layer0_outputs(8211) <= not(inputs(210)) or (inputs(254));
    layer0_outputs(8212) <= not(inputs(54));
    layer0_outputs(8213) <= not(inputs(97)) or (inputs(62));
    layer0_outputs(8214) <= (inputs(170)) or (inputs(165));
    layer0_outputs(8215) <= inputs(196);
    layer0_outputs(8216) <= (inputs(88)) or (inputs(223));
    layer0_outputs(8217) <= inputs(83);
    layer0_outputs(8218) <= (inputs(178)) or (inputs(92));
    layer0_outputs(8219) <= not(inputs(76));
    layer0_outputs(8220) <= not(inputs(181));
    layer0_outputs(8221) <= (inputs(225)) and not (inputs(63));
    layer0_outputs(8222) <= not(inputs(149)) or (inputs(207));
    layer0_outputs(8223) <= not(inputs(154));
    layer0_outputs(8224) <= not(inputs(66));
    layer0_outputs(8225) <= inputs(198);
    layer0_outputs(8226) <= not((inputs(13)) xor (inputs(57)));
    layer0_outputs(8227) <= not(inputs(194));
    layer0_outputs(8228) <= (inputs(20)) and (inputs(242));
    layer0_outputs(8229) <= not((inputs(111)) or (inputs(13)));
    layer0_outputs(8230) <= (inputs(39)) and not (inputs(226));
    layer0_outputs(8231) <= (inputs(20)) xor (inputs(65));
    layer0_outputs(8232) <= (inputs(159)) or (inputs(26));
    layer0_outputs(8233) <= (inputs(160)) and not (inputs(137));
    layer0_outputs(8234) <= not(inputs(56));
    layer0_outputs(8235) <= not(inputs(46));
    layer0_outputs(8236) <= inputs(119);
    layer0_outputs(8237) <= (inputs(74)) and not (inputs(47));
    layer0_outputs(8238) <= not((inputs(149)) xor (inputs(138)));
    layer0_outputs(8239) <= inputs(50);
    layer0_outputs(8240) <= not(inputs(47)) or (inputs(221));
    layer0_outputs(8241) <= not(inputs(113));
    layer0_outputs(8242) <= (inputs(89)) and not (inputs(209));
    layer0_outputs(8243) <= not((inputs(6)) xor (inputs(133)));
    layer0_outputs(8244) <= (inputs(245)) xor (inputs(213));
    layer0_outputs(8245) <= (inputs(195)) xor (inputs(211));
    layer0_outputs(8246) <= (inputs(102)) and not (inputs(73));
    layer0_outputs(8247) <= not(inputs(44));
    layer0_outputs(8248) <= inputs(22);
    layer0_outputs(8249) <= (inputs(216)) and not (inputs(44));
    layer0_outputs(8250) <= not(inputs(176));
    layer0_outputs(8251) <= not(inputs(217));
    layer0_outputs(8252) <= not((inputs(22)) or (inputs(36)));
    layer0_outputs(8253) <= (inputs(162)) and not (inputs(64));
    layer0_outputs(8254) <= not(inputs(221)) or (inputs(152));
    layer0_outputs(8255) <= inputs(91);
    layer0_outputs(8256) <= not((inputs(230)) xor (inputs(195)));
    layer0_outputs(8257) <= (inputs(50)) or (inputs(115));
    layer0_outputs(8258) <= inputs(152);
    layer0_outputs(8259) <= not(inputs(93)) or (inputs(79));
    layer0_outputs(8260) <= (inputs(10)) xor (inputs(254));
    layer0_outputs(8261) <= (inputs(88)) and (inputs(44));
    layer0_outputs(8262) <= (inputs(172)) xor (inputs(115));
    layer0_outputs(8263) <= not(inputs(116));
    layer0_outputs(8264) <= '1';
    layer0_outputs(8265) <= not((inputs(135)) and (inputs(5)));
    layer0_outputs(8266) <= (inputs(118)) or (inputs(234));
    layer0_outputs(8267) <= not((inputs(252)) or (inputs(39)));
    layer0_outputs(8268) <= inputs(160);
    layer0_outputs(8269) <= not(inputs(246));
    layer0_outputs(8270) <= not(inputs(77));
    layer0_outputs(8271) <= not(inputs(45)) or (inputs(138));
    layer0_outputs(8272) <= not((inputs(57)) or (inputs(240)));
    layer0_outputs(8273) <= (inputs(130)) and (inputs(211));
    layer0_outputs(8274) <= not((inputs(94)) xor (inputs(219)));
    layer0_outputs(8275) <= '1';
    layer0_outputs(8276) <= not((inputs(197)) xor (inputs(1)));
    layer0_outputs(8277) <= (inputs(73)) and not (inputs(15));
    layer0_outputs(8278) <= (inputs(107)) or (inputs(37));
    layer0_outputs(8279) <= not(inputs(55)) or (inputs(132));
    layer0_outputs(8280) <= not(inputs(20)) or (inputs(188));
    layer0_outputs(8281) <= inputs(150);
    layer0_outputs(8282) <= (inputs(27)) xor (inputs(166));
    layer0_outputs(8283) <= not(inputs(252));
    layer0_outputs(8284) <= not((inputs(193)) or (inputs(161)));
    layer0_outputs(8285) <= (inputs(89)) xor (inputs(118));
    layer0_outputs(8286) <= inputs(118);
    layer0_outputs(8287) <= (inputs(122)) and not (inputs(112));
    layer0_outputs(8288) <= not(inputs(174));
    layer0_outputs(8289) <= (inputs(234)) xor (inputs(221));
    layer0_outputs(8290) <= not(inputs(247));
    layer0_outputs(8291) <= inputs(22);
    layer0_outputs(8292) <= not(inputs(110)) or (inputs(243));
    layer0_outputs(8293) <= inputs(85);
    layer0_outputs(8294) <= not(inputs(70));
    layer0_outputs(8295) <= (inputs(144)) or (inputs(100));
    layer0_outputs(8296) <= (inputs(64)) or (inputs(82));
    layer0_outputs(8297) <= not((inputs(18)) xor (inputs(4)));
    layer0_outputs(8298) <= not((inputs(79)) or (inputs(221)));
    layer0_outputs(8299) <= not(inputs(137)) or (inputs(88));
    layer0_outputs(8300) <= (inputs(130)) and (inputs(178));
    layer0_outputs(8301) <= not((inputs(117)) or (inputs(48)));
    layer0_outputs(8302) <= not((inputs(62)) and (inputs(86)));
    layer0_outputs(8303) <= (inputs(248)) and not (inputs(199));
    layer0_outputs(8304) <= not((inputs(129)) or (inputs(83)));
    layer0_outputs(8305) <= not((inputs(25)) and (inputs(244)));
    layer0_outputs(8306) <= (inputs(131)) and not (inputs(229));
    layer0_outputs(8307) <= (inputs(79)) xor (inputs(125));
    layer0_outputs(8308) <= not(inputs(104));
    layer0_outputs(8309) <= (inputs(134)) and not (inputs(93));
    layer0_outputs(8310) <= not(inputs(51));
    layer0_outputs(8311) <= inputs(252);
    layer0_outputs(8312) <= inputs(181);
    layer0_outputs(8313) <= inputs(93);
    layer0_outputs(8314) <= not((inputs(153)) and (inputs(243)));
    layer0_outputs(8315) <= (inputs(37)) and not (inputs(209));
    layer0_outputs(8316) <= not((inputs(213)) or (inputs(19)));
    layer0_outputs(8317) <= not(inputs(203)) or (inputs(87));
    layer0_outputs(8318) <= (inputs(195)) or (inputs(70));
    layer0_outputs(8319) <= (inputs(10)) or (inputs(227));
    layer0_outputs(8320) <= inputs(255);
    layer0_outputs(8321) <= not(inputs(217)) or (inputs(86));
    layer0_outputs(8322) <= (inputs(164)) and not (inputs(88));
    layer0_outputs(8323) <= (inputs(170)) or (inputs(145));
    layer0_outputs(8324) <= inputs(91);
    layer0_outputs(8325) <= not(inputs(73)) or (inputs(4));
    layer0_outputs(8326) <= (inputs(219)) or (inputs(150));
    layer0_outputs(8327) <= not(inputs(97));
    layer0_outputs(8328) <= not((inputs(92)) or (inputs(2)));
    layer0_outputs(8329) <= not(inputs(246));
    layer0_outputs(8330) <= inputs(233);
    layer0_outputs(8331) <= not((inputs(248)) or (inputs(192)));
    layer0_outputs(8332) <= not(inputs(62));
    layer0_outputs(8333) <= (inputs(27)) xor (inputs(160));
    layer0_outputs(8334) <= not(inputs(31));
    layer0_outputs(8335) <= not(inputs(115));
    layer0_outputs(8336) <= not(inputs(232)) or (inputs(101));
    layer0_outputs(8337) <= not(inputs(179));
    layer0_outputs(8338) <= (inputs(20)) xor (inputs(80));
    layer0_outputs(8339) <= not((inputs(34)) and (inputs(156)));
    layer0_outputs(8340) <= inputs(157);
    layer0_outputs(8341) <= not(inputs(83));
    layer0_outputs(8342) <= (inputs(185)) xor (inputs(196));
    layer0_outputs(8343) <= not(inputs(121)) or (inputs(174));
    layer0_outputs(8344) <= (inputs(14)) or (inputs(83));
    layer0_outputs(8345) <= (inputs(77)) and not (inputs(198));
    layer0_outputs(8346) <= (inputs(215)) and (inputs(214));
    layer0_outputs(8347) <= inputs(189);
    layer0_outputs(8348) <= (inputs(214)) or (inputs(232));
    layer0_outputs(8349) <= not((inputs(206)) xor (inputs(165)));
    layer0_outputs(8350) <= not(inputs(78));
    layer0_outputs(8351) <= (inputs(253)) or (inputs(75));
    layer0_outputs(8352) <= not((inputs(199)) xor (inputs(241)));
    layer0_outputs(8353) <= not(inputs(166));
    layer0_outputs(8354) <= (inputs(121)) or (inputs(82));
    layer0_outputs(8355) <= not(inputs(137)) or (inputs(242));
    layer0_outputs(8356) <= inputs(140);
    layer0_outputs(8357) <= '1';
    layer0_outputs(8358) <= inputs(197);
    layer0_outputs(8359) <= not((inputs(197)) xor (inputs(58)));
    layer0_outputs(8360) <= (inputs(219)) and not (inputs(122));
    layer0_outputs(8361) <= inputs(142);
    layer0_outputs(8362) <= inputs(39);
    layer0_outputs(8363) <= inputs(25);
    layer0_outputs(8364) <= inputs(114);
    layer0_outputs(8365) <= (inputs(73)) xor (inputs(170));
    layer0_outputs(8366) <= not((inputs(13)) or (inputs(216)));
    layer0_outputs(8367) <= (inputs(133)) and not (inputs(253));
    layer0_outputs(8368) <= inputs(196);
    layer0_outputs(8369) <= inputs(184);
    layer0_outputs(8370) <= not((inputs(140)) or (inputs(58)));
    layer0_outputs(8371) <= inputs(139);
    layer0_outputs(8372) <= inputs(107);
    layer0_outputs(8373) <= not(inputs(204)) or (inputs(252));
    layer0_outputs(8374) <= not(inputs(172)) or (inputs(57));
    layer0_outputs(8375) <= (inputs(30)) and (inputs(143));
    layer0_outputs(8376) <= not((inputs(247)) or (inputs(124)));
    layer0_outputs(8377) <= not(inputs(109));
    layer0_outputs(8378) <= not((inputs(84)) or (inputs(85)));
    layer0_outputs(8379) <= not(inputs(70)) or (inputs(127));
    layer0_outputs(8380) <= not((inputs(193)) xor (inputs(227)));
    layer0_outputs(8381) <= (inputs(213)) or (inputs(205));
    layer0_outputs(8382) <= not((inputs(192)) or (inputs(177)));
    layer0_outputs(8383) <= not(inputs(115)) or (inputs(57));
    layer0_outputs(8384) <= not(inputs(211)) or (inputs(92));
    layer0_outputs(8385) <= not(inputs(82));
    layer0_outputs(8386) <= not(inputs(172)) or (inputs(239));
    layer0_outputs(8387) <= inputs(237);
    layer0_outputs(8388) <= inputs(155);
    layer0_outputs(8389) <= inputs(76);
    layer0_outputs(8390) <= inputs(78);
    layer0_outputs(8391) <= not(inputs(35));
    layer0_outputs(8392) <= (inputs(7)) or (inputs(177));
    layer0_outputs(8393) <= not(inputs(194));
    layer0_outputs(8394) <= (inputs(127)) or (inputs(163));
    layer0_outputs(8395) <= (inputs(132)) xor (inputs(168));
    layer0_outputs(8396) <= not(inputs(231));
    layer0_outputs(8397) <= not(inputs(54));
    layer0_outputs(8398) <= not((inputs(74)) or (inputs(4)));
    layer0_outputs(8399) <= (inputs(109)) and (inputs(56));
    layer0_outputs(8400) <= inputs(230);
    layer0_outputs(8401) <= inputs(40);
    layer0_outputs(8402) <= (inputs(118)) or (inputs(244));
    layer0_outputs(8403) <= not(inputs(228));
    layer0_outputs(8404) <= inputs(74);
    layer0_outputs(8405) <= not((inputs(33)) xor (inputs(121)));
    layer0_outputs(8406) <= (inputs(218)) or (inputs(236));
    layer0_outputs(8407) <= (inputs(132)) or (inputs(163));
    layer0_outputs(8408) <= not(inputs(90));
    layer0_outputs(8409) <= (inputs(239)) or (inputs(213));
    layer0_outputs(8410) <= (inputs(95)) or (inputs(102));
    layer0_outputs(8411) <= not(inputs(174)) or (inputs(189));
    layer0_outputs(8412) <= not((inputs(232)) or (inputs(87)));
    layer0_outputs(8413) <= not(inputs(84)) or (inputs(242));
    layer0_outputs(8414) <= (inputs(112)) and not (inputs(249));
    layer0_outputs(8415) <= (inputs(78)) xor (inputs(149));
    layer0_outputs(8416) <= not(inputs(182));
    layer0_outputs(8417) <= (inputs(159)) and not (inputs(67));
    layer0_outputs(8418) <= not(inputs(13));
    layer0_outputs(8419) <= '0';
    layer0_outputs(8420) <= not(inputs(214)) or (inputs(33));
    layer0_outputs(8421) <= (inputs(20)) and not (inputs(88));
    layer0_outputs(8422) <= inputs(192);
    layer0_outputs(8423) <= (inputs(116)) xor (inputs(200));
    layer0_outputs(8424) <= not(inputs(53)) or (inputs(240));
    layer0_outputs(8425) <= not(inputs(13));
    layer0_outputs(8426) <= not(inputs(148));
    layer0_outputs(8427) <= (inputs(61)) and not (inputs(190));
    layer0_outputs(8428) <= (inputs(26)) and not (inputs(250));
    layer0_outputs(8429) <= not((inputs(38)) xor (inputs(250)));
    layer0_outputs(8430) <= (inputs(135)) and not (inputs(18));
    layer0_outputs(8431) <= not(inputs(154)) or (inputs(192));
    layer0_outputs(8432) <= not((inputs(59)) xor (inputs(168)));
    layer0_outputs(8433) <= not((inputs(47)) or (inputs(193)));
    layer0_outputs(8434) <= not(inputs(228)) or (inputs(109));
    layer0_outputs(8435) <= (inputs(151)) and (inputs(250));
    layer0_outputs(8436) <= not(inputs(58)) or (inputs(184));
    layer0_outputs(8437) <= '0';
    layer0_outputs(8438) <= not((inputs(157)) xor (inputs(15)));
    layer0_outputs(8439) <= not(inputs(161)) or (inputs(94));
    layer0_outputs(8440) <= not((inputs(249)) xor (inputs(126)));
    layer0_outputs(8441) <= not(inputs(221));
    layer0_outputs(8442) <= (inputs(84)) xor (inputs(112));
    layer0_outputs(8443) <= (inputs(24)) and not (inputs(255));
    layer0_outputs(8444) <= not((inputs(4)) or (inputs(147)));
    layer0_outputs(8445) <= (inputs(31)) or (inputs(52));
    layer0_outputs(8446) <= not((inputs(141)) or (inputs(179)));
    layer0_outputs(8447) <= inputs(38);
    layer0_outputs(8448) <= not(inputs(237));
    layer0_outputs(8449) <= inputs(153);
    layer0_outputs(8450) <= not((inputs(234)) or (inputs(201)));
    layer0_outputs(8451) <= not(inputs(121));
    layer0_outputs(8452) <= '1';
    layer0_outputs(8453) <= (inputs(131)) xor (inputs(102));
    layer0_outputs(8454) <= inputs(132);
    layer0_outputs(8455) <= (inputs(239)) or (inputs(181));
    layer0_outputs(8456) <= inputs(230);
    layer0_outputs(8457) <= not(inputs(59));
    layer0_outputs(8458) <= not((inputs(209)) and (inputs(193)));
    layer0_outputs(8459) <= (inputs(110)) xor (inputs(61));
    layer0_outputs(8460) <= inputs(230);
    layer0_outputs(8461) <= (inputs(11)) or (inputs(196));
    layer0_outputs(8462) <= not(inputs(29));
    layer0_outputs(8463) <= not(inputs(189)) or (inputs(184));
    layer0_outputs(8464) <= not(inputs(7));
    layer0_outputs(8465) <= not(inputs(116));
    layer0_outputs(8466) <= not(inputs(113));
    layer0_outputs(8467) <= (inputs(173)) and not (inputs(83));
    layer0_outputs(8468) <= inputs(136);
    layer0_outputs(8469) <= (inputs(204)) and not (inputs(65));
    layer0_outputs(8470) <= (inputs(149)) xor (inputs(241));
    layer0_outputs(8471) <= inputs(55);
    layer0_outputs(8472) <= (inputs(179)) or (inputs(237));
    layer0_outputs(8473) <= (inputs(215)) and not (inputs(132));
    layer0_outputs(8474) <= inputs(203);
    layer0_outputs(8475) <= not(inputs(147)) or (inputs(142));
    layer0_outputs(8476) <= not(inputs(166)) or (inputs(209));
    layer0_outputs(8477) <= not(inputs(140)) or (inputs(178));
    layer0_outputs(8478) <= not((inputs(60)) or (inputs(37)));
    layer0_outputs(8479) <= not(inputs(81)) or (inputs(169));
    layer0_outputs(8480) <= (inputs(235)) and not (inputs(100));
    layer0_outputs(8481) <= not(inputs(141));
    layer0_outputs(8482) <= inputs(146);
    layer0_outputs(8483) <= (inputs(199)) and not (inputs(40));
    layer0_outputs(8484) <= (inputs(128)) xor (inputs(246));
    layer0_outputs(8485) <= inputs(222);
    layer0_outputs(8486) <= (inputs(75)) and not (inputs(209));
    layer0_outputs(8487) <= '0';
    layer0_outputs(8488) <= not(inputs(183)) or (inputs(208));
    layer0_outputs(8489) <= (inputs(239)) or (inputs(228));
    layer0_outputs(8490) <= '1';
    layer0_outputs(8491) <= not(inputs(40));
    layer0_outputs(8492) <= not((inputs(208)) or (inputs(244)));
    layer0_outputs(8493) <= not(inputs(10));
    layer0_outputs(8494) <= (inputs(207)) or (inputs(167));
    layer0_outputs(8495) <= not(inputs(223));
    layer0_outputs(8496) <= not((inputs(204)) xor (inputs(147)));
    layer0_outputs(8497) <= not((inputs(204)) and (inputs(39)));
    layer0_outputs(8498) <= not(inputs(148));
    layer0_outputs(8499) <= (inputs(174)) and not (inputs(237));
    layer0_outputs(8500) <= (inputs(117)) and not (inputs(251));
    layer0_outputs(8501) <= not(inputs(126));
    layer0_outputs(8502) <= not(inputs(227));
    layer0_outputs(8503) <= (inputs(11)) or (inputs(82));
    layer0_outputs(8504) <= not(inputs(100)) or (inputs(223));
    layer0_outputs(8505) <= not((inputs(253)) or (inputs(182)));
    layer0_outputs(8506) <= not(inputs(22));
    layer0_outputs(8507) <= (inputs(240)) or (inputs(188));
    layer0_outputs(8508) <= not((inputs(61)) xor (inputs(63)));
    layer0_outputs(8509) <= (inputs(47)) xor (inputs(3));
    layer0_outputs(8510) <= inputs(110);
    layer0_outputs(8511) <= not((inputs(253)) xor (inputs(52)));
    layer0_outputs(8512) <= not((inputs(38)) or (inputs(62)));
    layer0_outputs(8513) <= (inputs(143)) and not (inputs(194));
    layer0_outputs(8514) <= (inputs(12)) and not (inputs(221));
    layer0_outputs(8515) <= inputs(230);
    layer0_outputs(8516) <= (inputs(97)) or (inputs(254));
    layer0_outputs(8517) <= not((inputs(170)) or (inputs(230)));
    layer0_outputs(8518) <= inputs(111);
    layer0_outputs(8519) <= (inputs(147)) xor (inputs(184));
    layer0_outputs(8520) <= (inputs(46)) or (inputs(232));
    layer0_outputs(8521) <= (inputs(151)) or (inputs(77));
    layer0_outputs(8522) <= (inputs(72)) and not (inputs(62));
    layer0_outputs(8523) <= inputs(115);
    layer0_outputs(8524) <= not((inputs(5)) and (inputs(178)));
    layer0_outputs(8525) <= not(inputs(51)) or (inputs(145));
    layer0_outputs(8526) <= (inputs(18)) or (inputs(185));
    layer0_outputs(8527) <= not(inputs(100));
    layer0_outputs(8528) <= not(inputs(221)) or (inputs(94));
    layer0_outputs(8529) <= not((inputs(72)) or (inputs(249)));
    layer0_outputs(8530) <= (inputs(39)) and not (inputs(173));
    layer0_outputs(8531) <= (inputs(100)) or (inputs(249));
    layer0_outputs(8532) <= '1';
    layer0_outputs(8533) <= (inputs(121)) xor (inputs(251));
    layer0_outputs(8534) <= not(inputs(30));
    layer0_outputs(8535) <= not((inputs(56)) or (inputs(210)));
    layer0_outputs(8536) <= (inputs(13)) and not (inputs(239));
    layer0_outputs(8537) <= (inputs(8)) xor (inputs(189));
    layer0_outputs(8538) <= (inputs(118)) xor (inputs(149));
    layer0_outputs(8539) <= (inputs(143)) and not (inputs(239));
    layer0_outputs(8540) <= not((inputs(100)) or (inputs(113)));
    layer0_outputs(8541) <= not(inputs(78));
    layer0_outputs(8542) <= inputs(193);
    layer0_outputs(8543) <= not((inputs(194)) or (inputs(198)));
    layer0_outputs(8544) <= (inputs(188)) xor (inputs(136));
    layer0_outputs(8545) <= (inputs(100)) xor (inputs(126));
    layer0_outputs(8546) <= (inputs(161)) xor (inputs(152));
    layer0_outputs(8547) <= inputs(26);
    layer0_outputs(8548) <= (inputs(55)) and not (inputs(35));
    layer0_outputs(8549) <= (inputs(31)) xor (inputs(67));
    layer0_outputs(8550) <= not((inputs(94)) and (inputs(130)));
    layer0_outputs(8551) <= (inputs(198)) and not (inputs(42));
    layer0_outputs(8552) <= (inputs(36)) or (inputs(50));
    layer0_outputs(8553) <= inputs(130);
    layer0_outputs(8554) <= (inputs(100)) xor (inputs(72));
    layer0_outputs(8555) <= (inputs(60)) xor (inputs(143));
    layer0_outputs(8556) <= inputs(215);
    layer0_outputs(8557) <= not(inputs(254));
    layer0_outputs(8558) <= inputs(121);
    layer0_outputs(8559) <= not(inputs(95)) or (inputs(129));
    layer0_outputs(8560) <= not(inputs(213));
    layer0_outputs(8561) <= (inputs(250)) or (inputs(210));
    layer0_outputs(8562) <= not(inputs(80));
    layer0_outputs(8563) <= inputs(17);
    layer0_outputs(8564) <= (inputs(157)) and not (inputs(61));
    layer0_outputs(8565) <= inputs(215);
    layer0_outputs(8566) <= '0';
    layer0_outputs(8567) <= inputs(53);
    layer0_outputs(8568) <= not((inputs(202)) or (inputs(218)));
    layer0_outputs(8569) <= (inputs(48)) and not (inputs(12));
    layer0_outputs(8570) <= '0';
    layer0_outputs(8571) <= inputs(24);
    layer0_outputs(8572) <= not(inputs(168)) or (inputs(34));
    layer0_outputs(8573) <= not((inputs(78)) xor (inputs(248)));
    layer0_outputs(8574) <= (inputs(18)) and not (inputs(199));
    layer0_outputs(8575) <= inputs(235);
    layer0_outputs(8576) <= inputs(211);
    layer0_outputs(8577) <= not(inputs(142)) or (inputs(220));
    layer0_outputs(8578) <= (inputs(153)) and not (inputs(38));
    layer0_outputs(8579) <= not((inputs(237)) and (inputs(218)));
    layer0_outputs(8580) <= not((inputs(252)) or (inputs(177)));
    layer0_outputs(8581) <= not((inputs(119)) or (inputs(121)));
    layer0_outputs(8582) <= (inputs(211)) or (inputs(84));
    layer0_outputs(8583) <= not((inputs(218)) xor (inputs(115)));
    layer0_outputs(8584) <= not((inputs(27)) xor (inputs(233)));
    layer0_outputs(8585) <= (inputs(56)) and not (inputs(18));
    layer0_outputs(8586) <= not((inputs(230)) or (inputs(223)));
    layer0_outputs(8587) <= not(inputs(99));
    layer0_outputs(8588) <= inputs(196);
    layer0_outputs(8589) <= not((inputs(103)) and (inputs(89)));
    layer0_outputs(8590) <= inputs(81);
    layer0_outputs(8591) <= not((inputs(76)) xor (inputs(109)));
    layer0_outputs(8592) <= not(inputs(120));
    layer0_outputs(8593) <= not((inputs(152)) and (inputs(86)));
    layer0_outputs(8594) <= not(inputs(212)) or (inputs(76));
    layer0_outputs(8595) <= (inputs(176)) xor (inputs(138));
    layer0_outputs(8596) <= (inputs(133)) and not (inputs(13));
    layer0_outputs(8597) <= not((inputs(192)) or (inputs(216)));
    layer0_outputs(8598) <= not(inputs(132));
    layer0_outputs(8599) <= (inputs(2)) or (inputs(156));
    layer0_outputs(8600) <= (inputs(186)) or (inputs(163));
    layer0_outputs(8601) <= not(inputs(61));
    layer0_outputs(8602) <= (inputs(250)) and not (inputs(75));
    layer0_outputs(8603) <= not((inputs(214)) or (inputs(188)));
    layer0_outputs(8604) <= inputs(209);
    layer0_outputs(8605) <= not((inputs(59)) xor (inputs(131)));
    layer0_outputs(8606) <= (inputs(108)) or (inputs(253));
    layer0_outputs(8607) <= not(inputs(137)) or (inputs(102));
    layer0_outputs(8608) <= not((inputs(222)) or (inputs(5)));
    layer0_outputs(8609) <= not(inputs(187)) or (inputs(223));
    layer0_outputs(8610) <= (inputs(178)) xor (inputs(249));
    layer0_outputs(8611) <= not((inputs(146)) xor (inputs(70)));
    layer0_outputs(8612) <= not((inputs(68)) or (inputs(114)));
    layer0_outputs(8613) <= (inputs(186)) and (inputs(48));
    layer0_outputs(8614) <= (inputs(191)) and not (inputs(14));
    layer0_outputs(8615) <= (inputs(25)) and not (inputs(159));
    layer0_outputs(8616) <= (inputs(213)) xor (inputs(122));
    layer0_outputs(8617) <= not(inputs(151));
    layer0_outputs(8618) <= (inputs(131)) and not (inputs(35));
    layer0_outputs(8619) <= (inputs(7)) xor (inputs(69));
    layer0_outputs(8620) <= not((inputs(212)) and (inputs(215)));
    layer0_outputs(8621) <= not((inputs(3)) xor (inputs(139)));
    layer0_outputs(8622) <= (inputs(229)) and not (inputs(143));
    layer0_outputs(8623) <= not((inputs(71)) or (inputs(227)));
    layer0_outputs(8624) <= not((inputs(177)) or (inputs(11)));
    layer0_outputs(8625) <= inputs(184);
    layer0_outputs(8626) <= not(inputs(153));
    layer0_outputs(8627) <= (inputs(134)) xor (inputs(87));
    layer0_outputs(8628) <= (inputs(98)) and (inputs(134));
    layer0_outputs(8629) <= not(inputs(64));
    layer0_outputs(8630) <= inputs(130);
    layer0_outputs(8631) <= not(inputs(198));
    layer0_outputs(8632) <= not((inputs(188)) or (inputs(75)));
    layer0_outputs(8633) <= not(inputs(182)) or (inputs(97));
    layer0_outputs(8634) <= not(inputs(148));
    layer0_outputs(8635) <= inputs(164);
    layer0_outputs(8636) <= (inputs(237)) or (inputs(145));
    layer0_outputs(8637) <= not((inputs(199)) or (inputs(8)));
    layer0_outputs(8638) <= inputs(46);
    layer0_outputs(8639) <= inputs(193);
    layer0_outputs(8640) <= (inputs(191)) or (inputs(189));
    layer0_outputs(8641) <= (inputs(103)) and not (inputs(163));
    layer0_outputs(8642) <= (inputs(64)) and not (inputs(112));
    layer0_outputs(8643) <= not((inputs(17)) or (inputs(182)));
    layer0_outputs(8644) <= '0';
    layer0_outputs(8645) <= (inputs(119)) xor (inputs(106));
    layer0_outputs(8646) <= not(inputs(128));
    layer0_outputs(8647) <= not((inputs(194)) xor (inputs(247)));
    layer0_outputs(8648) <= (inputs(179)) or (inputs(87));
    layer0_outputs(8649) <= inputs(22);
    layer0_outputs(8650) <= not((inputs(26)) xor (inputs(64)));
    layer0_outputs(8651) <= not((inputs(227)) or (inputs(132)));
    layer0_outputs(8652) <= inputs(18);
    layer0_outputs(8653) <= inputs(45);
    layer0_outputs(8654) <= (inputs(55)) and (inputs(49));
    layer0_outputs(8655) <= not((inputs(202)) or (inputs(233)));
    layer0_outputs(8656) <= inputs(207);
    layer0_outputs(8657) <= (inputs(230)) and not (inputs(56));
    layer0_outputs(8658) <= not(inputs(139)) or (inputs(163));
    layer0_outputs(8659) <= (inputs(184)) and not (inputs(163));
    layer0_outputs(8660) <= not((inputs(207)) xor (inputs(19)));
    layer0_outputs(8661) <= inputs(168);
    layer0_outputs(8662) <= inputs(197);
    layer0_outputs(8663) <= not((inputs(240)) xor (inputs(213)));
    layer0_outputs(8664) <= (inputs(233)) and not (inputs(96));
    layer0_outputs(8665) <= not(inputs(118));
    layer0_outputs(8666) <= inputs(187);
    layer0_outputs(8667) <= not(inputs(253));
    layer0_outputs(8668) <= not(inputs(85));
    layer0_outputs(8669) <= (inputs(247)) and not (inputs(177));
    layer0_outputs(8670) <= (inputs(72)) xor (inputs(46));
    layer0_outputs(8671) <= not(inputs(8)) or (inputs(249));
    layer0_outputs(8672) <= (inputs(186)) and not (inputs(110));
    layer0_outputs(8673) <= inputs(211);
    layer0_outputs(8674) <= (inputs(110)) or (inputs(253));
    layer0_outputs(8675) <= inputs(205);
    layer0_outputs(8676) <= not(inputs(105)) or (inputs(209));
    layer0_outputs(8677) <= (inputs(226)) xor (inputs(181));
    layer0_outputs(8678) <= (inputs(36)) or (inputs(255));
    layer0_outputs(8679) <= not((inputs(75)) or (inputs(154)));
    layer0_outputs(8680) <= not(inputs(51));
    layer0_outputs(8681) <= not(inputs(22));
    layer0_outputs(8682) <= '1';
    layer0_outputs(8683) <= inputs(203);
    layer0_outputs(8684) <= (inputs(174)) or (inputs(245));
    layer0_outputs(8685) <= not(inputs(230));
    layer0_outputs(8686) <= not(inputs(207));
    layer0_outputs(8687) <= (inputs(42)) or (inputs(155));
    layer0_outputs(8688) <= inputs(85);
    layer0_outputs(8689) <= not(inputs(150));
    layer0_outputs(8690) <= '1';
    layer0_outputs(8691) <= not((inputs(187)) xor (inputs(183)));
    layer0_outputs(8692) <= not((inputs(80)) or (inputs(64)));
    layer0_outputs(8693) <= not((inputs(187)) or (inputs(98)));
    layer0_outputs(8694) <= (inputs(145)) and not (inputs(79));
    layer0_outputs(8695) <= not(inputs(247));
    layer0_outputs(8696) <= inputs(71);
    layer0_outputs(8697) <= not((inputs(139)) or (inputs(45)));
    layer0_outputs(8698) <= inputs(167);
    layer0_outputs(8699) <= (inputs(96)) or (inputs(150));
    layer0_outputs(8700) <= not(inputs(87)) or (inputs(49));
    layer0_outputs(8701) <= (inputs(178)) or (inputs(252));
    layer0_outputs(8702) <= not((inputs(66)) xor (inputs(25)));
    layer0_outputs(8703) <= not((inputs(96)) or (inputs(129)));
    layer0_outputs(8704) <= not(inputs(99));
    layer0_outputs(8705) <= inputs(162);
    layer0_outputs(8706) <= inputs(177);
    layer0_outputs(8707) <= not(inputs(200));
    layer0_outputs(8708) <= (inputs(93)) and not (inputs(17));
    layer0_outputs(8709) <= (inputs(118)) and not (inputs(133));
    layer0_outputs(8710) <= (inputs(71)) and not (inputs(246));
    layer0_outputs(8711) <= not(inputs(4));
    layer0_outputs(8712) <= not((inputs(124)) and (inputs(44)));
    layer0_outputs(8713) <= not((inputs(33)) or (inputs(192)));
    layer0_outputs(8714) <= (inputs(228)) or (inputs(10));
    layer0_outputs(8715) <= not(inputs(114));
    layer0_outputs(8716) <= not((inputs(157)) xor (inputs(4)));
    layer0_outputs(8717) <= not((inputs(1)) or (inputs(180)));
    layer0_outputs(8718) <= not(inputs(40));
    layer0_outputs(8719) <= inputs(67);
    layer0_outputs(8720) <= not(inputs(20));
    layer0_outputs(8721) <= (inputs(228)) or (inputs(230));
    layer0_outputs(8722) <= not(inputs(179));
    layer0_outputs(8723) <= not(inputs(145));
    layer0_outputs(8724) <= (inputs(146)) or (inputs(105));
    layer0_outputs(8725) <= not(inputs(18)) or (inputs(14));
    layer0_outputs(8726) <= inputs(103);
    layer0_outputs(8727) <= (inputs(220)) or (inputs(197));
    layer0_outputs(8728) <= not((inputs(189)) and (inputs(122)));
    layer0_outputs(8729) <= not((inputs(104)) or (inputs(192)));
    layer0_outputs(8730) <= (inputs(198)) xor (inputs(175));
    layer0_outputs(8731) <= inputs(43);
    layer0_outputs(8732) <= not(inputs(11));
    layer0_outputs(8733) <= not(inputs(156));
    layer0_outputs(8734) <= inputs(204);
    layer0_outputs(8735) <= inputs(188);
    layer0_outputs(8736) <= (inputs(36)) or (inputs(32));
    layer0_outputs(8737) <= not((inputs(96)) xor (inputs(83)));
    layer0_outputs(8738) <= not(inputs(132));
    layer0_outputs(8739) <= (inputs(251)) or (inputs(88));
    layer0_outputs(8740) <= inputs(111);
    layer0_outputs(8741) <= (inputs(28)) and not (inputs(160));
    layer0_outputs(8742) <= inputs(83);
    layer0_outputs(8743) <= not(inputs(91)) or (inputs(23));
    layer0_outputs(8744) <= (inputs(96)) xor (inputs(209));
    layer0_outputs(8745) <= not(inputs(202)) or (inputs(59));
    layer0_outputs(8746) <= not((inputs(114)) or (inputs(58)));
    layer0_outputs(8747) <= (inputs(146)) xor (inputs(104));
    layer0_outputs(8748) <= not(inputs(230));
    layer0_outputs(8749) <= (inputs(203)) and not (inputs(47));
    layer0_outputs(8750) <= (inputs(162)) or (inputs(94));
    layer0_outputs(8751) <= not(inputs(105));
    layer0_outputs(8752) <= not(inputs(152));
    layer0_outputs(8753) <= not(inputs(206));
    layer0_outputs(8754) <= not((inputs(64)) or (inputs(182)));
    layer0_outputs(8755) <= not(inputs(173)) or (inputs(158));
    layer0_outputs(8756) <= (inputs(0)) or (inputs(247));
    layer0_outputs(8757) <= not((inputs(163)) or (inputs(247)));
    layer0_outputs(8758) <= (inputs(176)) xor (inputs(45));
    layer0_outputs(8759) <= not(inputs(25));
    layer0_outputs(8760) <= (inputs(185)) xor (inputs(138));
    layer0_outputs(8761) <= (inputs(162)) or (inputs(91));
    layer0_outputs(8762) <= not(inputs(176));
    layer0_outputs(8763) <= not(inputs(246)) or (inputs(126));
    layer0_outputs(8764) <= inputs(78);
    layer0_outputs(8765) <= '1';
    layer0_outputs(8766) <= inputs(176);
    layer0_outputs(8767) <= (inputs(224)) and not (inputs(214));
    layer0_outputs(8768) <= not(inputs(117));
    layer0_outputs(8769) <= not((inputs(91)) or (inputs(240)));
    layer0_outputs(8770) <= not(inputs(94)) or (inputs(35));
    layer0_outputs(8771) <= not(inputs(86));
    layer0_outputs(8772) <= (inputs(207)) xor (inputs(142));
    layer0_outputs(8773) <= (inputs(233)) and not (inputs(46));
    layer0_outputs(8774) <= not((inputs(217)) and (inputs(204)));
    layer0_outputs(8775) <= not(inputs(59));
    layer0_outputs(8776) <= not(inputs(48));
    layer0_outputs(8777) <= not(inputs(197)) or (inputs(78));
    layer0_outputs(8778) <= '0';
    layer0_outputs(8779) <= (inputs(155)) and not (inputs(42));
    layer0_outputs(8780) <= (inputs(165)) or (inputs(248));
    layer0_outputs(8781) <= (inputs(165)) and not (inputs(59));
    layer0_outputs(8782) <= not(inputs(167)) or (inputs(47));
    layer0_outputs(8783) <= (inputs(254)) or (inputs(255));
    layer0_outputs(8784) <= (inputs(48)) or (inputs(234));
    layer0_outputs(8785) <= (inputs(35)) and not (inputs(173));
    layer0_outputs(8786) <= not((inputs(163)) or (inputs(134)));
    layer0_outputs(8787) <= (inputs(92)) xor (inputs(19));
    layer0_outputs(8788) <= not(inputs(44));
    layer0_outputs(8789) <= '0';
    layer0_outputs(8790) <= (inputs(38)) xor (inputs(193));
    layer0_outputs(8791) <= not(inputs(32));
    layer0_outputs(8792) <= not((inputs(201)) or (inputs(249)));
    layer0_outputs(8793) <= inputs(30);
    layer0_outputs(8794) <= inputs(231);
    layer0_outputs(8795) <= not(inputs(133));
    layer0_outputs(8796) <= (inputs(148)) and not (inputs(130));
    layer0_outputs(8797) <= (inputs(124)) or (inputs(111));
    layer0_outputs(8798) <= (inputs(236)) and (inputs(17));
    layer0_outputs(8799) <= (inputs(149)) and not (inputs(2));
    layer0_outputs(8800) <= not(inputs(232));
    layer0_outputs(8801) <= not((inputs(53)) xor (inputs(59)));
    layer0_outputs(8802) <= (inputs(210)) or (inputs(145));
    layer0_outputs(8803) <= not(inputs(88));
    layer0_outputs(8804) <= (inputs(198)) or (inputs(149));
    layer0_outputs(8805) <= '1';
    layer0_outputs(8806) <= (inputs(14)) and not (inputs(5));
    layer0_outputs(8807) <= not(inputs(132)) or (inputs(201));
    layer0_outputs(8808) <= (inputs(167)) and not (inputs(143));
    layer0_outputs(8809) <= (inputs(176)) or (inputs(247));
    layer0_outputs(8810) <= '1';
    layer0_outputs(8811) <= not(inputs(136));
    layer0_outputs(8812) <= not((inputs(73)) xor (inputs(96)));
    layer0_outputs(8813) <= (inputs(211)) and not (inputs(68));
    layer0_outputs(8814) <= (inputs(52)) or (inputs(95));
    layer0_outputs(8815) <= not((inputs(145)) or (inputs(171)));
    layer0_outputs(8816) <= not(inputs(173)) or (inputs(111));
    layer0_outputs(8817) <= '0';
    layer0_outputs(8818) <= not((inputs(73)) and (inputs(184)));
    layer0_outputs(8819) <= not(inputs(207));
    layer0_outputs(8820) <= not(inputs(165)) or (inputs(192));
    layer0_outputs(8821) <= inputs(108);
    layer0_outputs(8822) <= (inputs(91)) or (inputs(108));
    layer0_outputs(8823) <= not(inputs(74)) or (inputs(145));
    layer0_outputs(8824) <= not(inputs(213));
    layer0_outputs(8825) <= (inputs(204)) xor (inputs(67));
    layer0_outputs(8826) <= not(inputs(245));
    layer0_outputs(8827) <= (inputs(86)) or (inputs(91));
    layer0_outputs(8828) <= not((inputs(64)) xor (inputs(240)));
    layer0_outputs(8829) <= not(inputs(14));
    layer0_outputs(8830) <= (inputs(248)) or (inputs(157));
    layer0_outputs(8831) <= not(inputs(86));
    layer0_outputs(8832) <= not(inputs(20));
    layer0_outputs(8833) <= inputs(240);
    layer0_outputs(8834) <= not(inputs(116)) or (inputs(208));
    layer0_outputs(8835) <= (inputs(118)) xor (inputs(51));
    layer0_outputs(8836) <= not((inputs(40)) or (inputs(14)));
    layer0_outputs(8837) <= not((inputs(232)) xor (inputs(70)));
    layer0_outputs(8838) <= (inputs(135)) and not (inputs(160));
    layer0_outputs(8839) <= (inputs(210)) and not (inputs(130));
    layer0_outputs(8840) <= (inputs(125)) and not (inputs(254));
    layer0_outputs(8841) <= not(inputs(110));
    layer0_outputs(8842) <= not(inputs(232));
    layer0_outputs(8843) <= not((inputs(145)) or (inputs(42)));
    layer0_outputs(8844) <= not((inputs(110)) xor (inputs(32)));
    layer0_outputs(8845) <= not((inputs(90)) xor (inputs(34)));
    layer0_outputs(8846) <= not(inputs(212));
    layer0_outputs(8847) <= not(inputs(6));
    layer0_outputs(8848) <= inputs(56);
    layer0_outputs(8849) <= not(inputs(141)) or (inputs(157));
    layer0_outputs(8850) <= not(inputs(177)) or (inputs(32));
    layer0_outputs(8851) <= (inputs(248)) and not (inputs(168));
    layer0_outputs(8852) <= (inputs(3)) xor (inputs(33));
    layer0_outputs(8853) <= not((inputs(197)) xor (inputs(242)));
    layer0_outputs(8854) <= not((inputs(97)) or (inputs(192)));
    layer0_outputs(8855) <= not(inputs(87)) or (inputs(244));
    layer0_outputs(8856) <= not(inputs(4));
    layer0_outputs(8857) <= (inputs(135)) or (inputs(236));
    layer0_outputs(8858) <= not(inputs(217));
    layer0_outputs(8859) <= not(inputs(116));
    layer0_outputs(8860) <= not(inputs(60));
    layer0_outputs(8861) <= inputs(193);
    layer0_outputs(8862) <= inputs(114);
    layer0_outputs(8863) <= inputs(67);
    layer0_outputs(8864) <= inputs(108);
    layer0_outputs(8865) <= (inputs(187)) and not (inputs(28));
    layer0_outputs(8866) <= not(inputs(253));
    layer0_outputs(8867) <= not(inputs(169)) or (inputs(226));
    layer0_outputs(8868) <= not(inputs(161)) or (inputs(2));
    layer0_outputs(8869) <= not((inputs(188)) or (inputs(189)));
    layer0_outputs(8870) <= '1';
    layer0_outputs(8871) <= inputs(117);
    layer0_outputs(8872) <= inputs(163);
    layer0_outputs(8873) <= not(inputs(21)) or (inputs(114));
    layer0_outputs(8874) <= not(inputs(230));
    layer0_outputs(8875) <= not((inputs(187)) or (inputs(111)));
    layer0_outputs(8876) <= not(inputs(125));
    layer0_outputs(8877) <= not(inputs(152)) or (inputs(64));
    layer0_outputs(8878) <= not(inputs(102));
    layer0_outputs(8879) <= inputs(212);
    layer0_outputs(8880) <= (inputs(99)) and not (inputs(250));
    layer0_outputs(8881) <= inputs(93);
    layer0_outputs(8882) <= not((inputs(115)) xor (inputs(203)));
    layer0_outputs(8883) <= not(inputs(94));
    layer0_outputs(8884) <= not((inputs(106)) xor (inputs(97)));
    layer0_outputs(8885) <= not(inputs(93));
    layer0_outputs(8886) <= not(inputs(34)) or (inputs(145));
    layer0_outputs(8887) <= not((inputs(171)) xor (inputs(159)));
    layer0_outputs(8888) <= not((inputs(119)) and (inputs(178)));
    layer0_outputs(8889) <= not((inputs(250)) or (inputs(204)));
    layer0_outputs(8890) <= not((inputs(249)) or (inputs(206)));
    layer0_outputs(8891) <= (inputs(207)) and not (inputs(97));
    layer0_outputs(8892) <= (inputs(145)) or (inputs(229));
    layer0_outputs(8893) <= not(inputs(210));
    layer0_outputs(8894) <= not((inputs(147)) or (inputs(226)));
    layer0_outputs(8895) <= not(inputs(81));
    layer0_outputs(8896) <= not(inputs(184));
    layer0_outputs(8897) <= not(inputs(88)) or (inputs(110));
    layer0_outputs(8898) <= inputs(57);
    layer0_outputs(8899) <= inputs(43);
    layer0_outputs(8900) <= (inputs(64)) or (inputs(222));
    layer0_outputs(8901) <= not((inputs(176)) or (inputs(41)));
    layer0_outputs(8902) <= not(inputs(228)) or (inputs(8));
    layer0_outputs(8903) <= (inputs(9)) xor (inputs(63));
    layer0_outputs(8904) <= not((inputs(169)) and (inputs(136)));
    layer0_outputs(8905) <= not(inputs(244)) or (inputs(103));
    layer0_outputs(8906) <= inputs(110);
    layer0_outputs(8907) <= (inputs(122)) xor (inputs(156));
    layer0_outputs(8908) <= not(inputs(218)) or (inputs(90));
    layer0_outputs(8909) <= inputs(133);
    layer0_outputs(8910) <= not(inputs(93));
    layer0_outputs(8911) <= inputs(114);
    layer0_outputs(8912) <= (inputs(50)) or (inputs(127));
    layer0_outputs(8913) <= (inputs(145)) xor (inputs(116));
    layer0_outputs(8914) <= not((inputs(240)) and (inputs(191)));
    layer0_outputs(8915) <= not((inputs(190)) xor (inputs(10)));
    layer0_outputs(8916) <= (inputs(200)) xor (inputs(16));
    layer0_outputs(8917) <= not((inputs(75)) or (inputs(159)));
    layer0_outputs(8918) <= inputs(147);
    layer0_outputs(8919) <= not(inputs(217)) or (inputs(74));
    layer0_outputs(8920) <= (inputs(0)) xor (inputs(193));
    layer0_outputs(8921) <= not(inputs(152));
    layer0_outputs(8922) <= (inputs(169)) or (inputs(168));
    layer0_outputs(8923) <= not((inputs(128)) or (inputs(122)));
    layer0_outputs(8924) <= not((inputs(40)) xor (inputs(130)));
    layer0_outputs(8925) <= inputs(191);
    layer0_outputs(8926) <= not(inputs(250));
    layer0_outputs(8927) <= (inputs(197)) and not (inputs(202));
    layer0_outputs(8928) <= not(inputs(95));
    layer0_outputs(8929) <= (inputs(221)) and not (inputs(110));
    layer0_outputs(8930) <= inputs(230);
    layer0_outputs(8931) <= (inputs(229)) and not (inputs(135));
    layer0_outputs(8932) <= not(inputs(23));
    layer0_outputs(8933) <= inputs(84);
    layer0_outputs(8934) <= inputs(248);
    layer0_outputs(8935) <= (inputs(215)) and (inputs(115));
    layer0_outputs(8936) <= (inputs(84)) and not (inputs(111));
    layer0_outputs(8937) <= not((inputs(22)) or (inputs(10)));
    layer0_outputs(8938) <= '0';
    layer0_outputs(8939) <= not(inputs(180)) or (inputs(103));
    layer0_outputs(8940) <= inputs(131);
    layer0_outputs(8941) <= not(inputs(84));
    layer0_outputs(8942) <= not((inputs(162)) xor (inputs(189)));
    layer0_outputs(8943) <= inputs(180);
    layer0_outputs(8944) <= not(inputs(199)) or (inputs(98));
    layer0_outputs(8945) <= not(inputs(187)) or (inputs(147));
    layer0_outputs(8946) <= not(inputs(0)) or (inputs(156));
    layer0_outputs(8947) <= inputs(214);
    layer0_outputs(8948) <= inputs(114);
    layer0_outputs(8949) <= not(inputs(246));
    layer0_outputs(8950) <= (inputs(106)) and not (inputs(195));
    layer0_outputs(8951) <= inputs(87);
    layer0_outputs(8952) <= not((inputs(11)) and (inputs(93)));
    layer0_outputs(8953) <= inputs(98);
    layer0_outputs(8954) <= not((inputs(30)) and (inputs(56)));
    layer0_outputs(8955) <= inputs(23);
    layer0_outputs(8956) <= (inputs(180)) xor (inputs(183));
    layer0_outputs(8957) <= inputs(125);
    layer0_outputs(8958) <= (inputs(56)) and not (inputs(6));
    layer0_outputs(8959) <= (inputs(83)) xor (inputs(76));
    layer0_outputs(8960) <= (inputs(170)) or (inputs(129));
    layer0_outputs(8961) <= not(inputs(249));
    layer0_outputs(8962) <= inputs(97);
    layer0_outputs(8963) <= not(inputs(54)) or (inputs(233));
    layer0_outputs(8964) <= inputs(234);
    layer0_outputs(8965) <= (inputs(72)) and not (inputs(34));
    layer0_outputs(8966) <= not(inputs(146));
    layer0_outputs(8967) <= not(inputs(158));
    layer0_outputs(8968) <= not(inputs(231));
    layer0_outputs(8969) <= (inputs(155)) or (inputs(249));
    layer0_outputs(8970) <= (inputs(90)) or (inputs(76));
    layer0_outputs(8971) <= (inputs(157)) or (inputs(122));
    layer0_outputs(8972) <= not(inputs(139)) or (inputs(145));
    layer0_outputs(8973) <= inputs(222);
    layer0_outputs(8974) <= (inputs(57)) xor (inputs(110));
    layer0_outputs(8975) <= (inputs(63)) or (inputs(58));
    layer0_outputs(8976) <= (inputs(123)) and not (inputs(212));
    layer0_outputs(8977) <= not(inputs(171));
    layer0_outputs(8978) <= (inputs(179)) and not (inputs(96));
    layer0_outputs(8979) <= not((inputs(190)) or (inputs(60)));
    layer0_outputs(8980) <= (inputs(251)) or (inputs(63));
    layer0_outputs(8981) <= not(inputs(90));
    layer0_outputs(8982) <= (inputs(72)) xor (inputs(44));
    layer0_outputs(8983) <= '1';
    layer0_outputs(8984) <= not(inputs(0));
    layer0_outputs(8985) <= (inputs(212)) or (inputs(81));
    layer0_outputs(8986) <= not((inputs(84)) or (inputs(50)));
    layer0_outputs(8987) <= (inputs(224)) and not (inputs(241));
    layer0_outputs(8988) <= not(inputs(103));
    layer0_outputs(8989) <= inputs(99);
    layer0_outputs(8990) <= (inputs(117)) and not (inputs(2));
    layer0_outputs(8991) <= (inputs(43)) and not (inputs(161));
    layer0_outputs(8992) <= not(inputs(66));
    layer0_outputs(8993) <= not((inputs(32)) or (inputs(63)));
    layer0_outputs(8994) <= not(inputs(43)) or (inputs(220));
    layer0_outputs(8995) <= (inputs(246)) and not (inputs(120));
    layer0_outputs(8996) <= (inputs(24)) and (inputs(106));
    layer0_outputs(8997) <= (inputs(221)) or (inputs(236));
    layer0_outputs(8998) <= (inputs(146)) or (inputs(176));
    layer0_outputs(8999) <= not((inputs(118)) or (inputs(199)));
    layer0_outputs(9000) <= not(inputs(39)) or (inputs(246));
    layer0_outputs(9001) <= inputs(104);
    layer0_outputs(9002) <= (inputs(67)) or (inputs(113));
    layer0_outputs(9003) <= not((inputs(12)) xor (inputs(100)));
    layer0_outputs(9004) <= (inputs(94)) xor (inputs(126));
    layer0_outputs(9005) <= not(inputs(190)) or (inputs(223));
    layer0_outputs(9006) <= (inputs(175)) or (inputs(141));
    layer0_outputs(9007) <= (inputs(144)) xor (inputs(178));
    layer0_outputs(9008) <= '0';
    layer0_outputs(9009) <= not((inputs(222)) or (inputs(187)));
    layer0_outputs(9010) <= not((inputs(64)) xor (inputs(24)));
    layer0_outputs(9011) <= not(inputs(83));
    layer0_outputs(9012) <= inputs(96);
    layer0_outputs(9013) <= not((inputs(80)) xor (inputs(77)));
    layer0_outputs(9014) <= not((inputs(59)) or (inputs(2)));
    layer0_outputs(9015) <= not(inputs(156)) or (inputs(254));
    layer0_outputs(9016) <= (inputs(125)) or (inputs(123));
    layer0_outputs(9017) <= (inputs(227)) or (inputs(208));
    layer0_outputs(9018) <= (inputs(42)) and not (inputs(133));
    layer0_outputs(9019) <= inputs(146);
    layer0_outputs(9020) <= inputs(232);
    layer0_outputs(9021) <= inputs(47);
    layer0_outputs(9022) <= not(inputs(83)) or (inputs(199));
    layer0_outputs(9023) <= not(inputs(130));
    layer0_outputs(9024) <= (inputs(157)) xor (inputs(78));
    layer0_outputs(9025) <= inputs(8);
    layer0_outputs(9026) <= not(inputs(66));
    layer0_outputs(9027) <= (inputs(23)) and not (inputs(174));
    layer0_outputs(9028) <= (inputs(143)) xor (inputs(204));
    layer0_outputs(9029) <= not(inputs(81)) or (inputs(178));
    layer0_outputs(9030) <= not((inputs(172)) or (inputs(128)));
    layer0_outputs(9031) <= not(inputs(84));
    layer0_outputs(9032) <= not((inputs(132)) or (inputs(146)));
    layer0_outputs(9033) <= not((inputs(1)) xor (inputs(43)));
    layer0_outputs(9034) <= not((inputs(82)) xor (inputs(203)));
    layer0_outputs(9035) <= not(inputs(51)) or (inputs(223));
    layer0_outputs(9036) <= not(inputs(66)) or (inputs(156));
    layer0_outputs(9037) <= (inputs(87)) xor (inputs(132));
    layer0_outputs(9038) <= (inputs(218)) and not (inputs(94));
    layer0_outputs(9039) <= not(inputs(75)) or (inputs(150));
    layer0_outputs(9040) <= (inputs(169)) or (inputs(70));
    layer0_outputs(9041) <= not((inputs(103)) or (inputs(159)));
    layer0_outputs(9042) <= (inputs(83)) or (inputs(168));
    layer0_outputs(9043) <= inputs(193);
    layer0_outputs(9044) <= inputs(189);
    layer0_outputs(9045) <= (inputs(1)) or (inputs(34));
    layer0_outputs(9046) <= not((inputs(219)) or (inputs(192)));
    layer0_outputs(9047) <= not(inputs(54)) or (inputs(158));
    layer0_outputs(9048) <= not(inputs(98));
    layer0_outputs(9049) <= not((inputs(134)) or (inputs(171)));
    layer0_outputs(9050) <= inputs(216);
    layer0_outputs(9051) <= (inputs(125)) and not (inputs(186));
    layer0_outputs(9052) <= (inputs(132)) and not (inputs(136));
    layer0_outputs(9053) <= inputs(158);
    layer0_outputs(9054) <= inputs(25);
    layer0_outputs(9055) <= not((inputs(219)) or (inputs(192)));
    layer0_outputs(9056) <= not((inputs(0)) xor (inputs(209)));
    layer0_outputs(9057) <= not(inputs(178));
    layer0_outputs(9058) <= not(inputs(11)) or (inputs(32));
    layer0_outputs(9059) <= not(inputs(84));
    layer0_outputs(9060) <= (inputs(58)) and not (inputs(37));
    layer0_outputs(9061) <= not(inputs(193));
    layer0_outputs(9062) <= (inputs(187)) and not (inputs(54));
    layer0_outputs(9063) <= not((inputs(212)) or (inputs(208)));
    layer0_outputs(9064) <= (inputs(98)) or (inputs(160));
    layer0_outputs(9065) <= '1';
    layer0_outputs(9066) <= (inputs(48)) xor (inputs(254));
    layer0_outputs(9067) <= (inputs(168)) or (inputs(233));
    layer0_outputs(9068) <= inputs(135);
    layer0_outputs(9069) <= not(inputs(80)) or (inputs(159));
    layer0_outputs(9070) <= not((inputs(14)) xor (inputs(45)));
    layer0_outputs(9071) <= not((inputs(205)) or (inputs(44)));
    layer0_outputs(9072) <= not(inputs(248));
    layer0_outputs(9073) <= not(inputs(181));
    layer0_outputs(9074) <= inputs(118);
    layer0_outputs(9075) <= (inputs(195)) and (inputs(59));
    layer0_outputs(9076) <= (inputs(215)) and not (inputs(253));
    layer0_outputs(9077) <= (inputs(100)) and not (inputs(202));
    layer0_outputs(9078) <= '0';
    layer0_outputs(9079) <= not(inputs(43)) or (inputs(179));
    layer0_outputs(9080) <= not((inputs(1)) or (inputs(162)));
    layer0_outputs(9081) <= (inputs(57)) or (inputs(202));
    layer0_outputs(9082) <= (inputs(83)) and not (inputs(249));
    layer0_outputs(9083) <= not(inputs(229));
    layer0_outputs(9084) <= (inputs(246)) xor (inputs(40));
    layer0_outputs(9085) <= (inputs(30)) or (inputs(67));
    layer0_outputs(9086) <= (inputs(39)) and (inputs(154));
    layer0_outputs(9087) <= not(inputs(201));
    layer0_outputs(9088) <= (inputs(116)) xor (inputs(129));
    layer0_outputs(9089) <= not((inputs(92)) or (inputs(239)));
    layer0_outputs(9090) <= not(inputs(217));
    layer0_outputs(9091) <= (inputs(161)) or (inputs(80));
    layer0_outputs(9092) <= not(inputs(241));
    layer0_outputs(9093) <= not(inputs(57));
    layer0_outputs(9094) <= not((inputs(37)) or (inputs(50)));
    layer0_outputs(9095) <= (inputs(46)) xor (inputs(18));
    layer0_outputs(9096) <= inputs(119);
    layer0_outputs(9097) <= not(inputs(92)) or (inputs(4));
    layer0_outputs(9098) <= not(inputs(107));
    layer0_outputs(9099) <= not((inputs(95)) and (inputs(145)));
    layer0_outputs(9100) <= not(inputs(170));
    layer0_outputs(9101) <= inputs(89);
    layer0_outputs(9102) <= not((inputs(249)) and (inputs(135)));
    layer0_outputs(9103) <= not(inputs(254));
    layer0_outputs(9104) <= inputs(124);
    layer0_outputs(9105) <= (inputs(242)) or (inputs(221));
    layer0_outputs(9106) <= not((inputs(56)) or (inputs(86)));
    layer0_outputs(9107) <= not(inputs(205)) or (inputs(87));
    layer0_outputs(9108) <= not(inputs(67)) or (inputs(235));
    layer0_outputs(9109) <= not((inputs(209)) or (inputs(252)));
    layer0_outputs(9110) <= inputs(56);
    layer0_outputs(9111) <= inputs(203);
    layer0_outputs(9112) <= not((inputs(25)) xor (inputs(47)));
    layer0_outputs(9113) <= not(inputs(146)) or (inputs(47));
    layer0_outputs(9114) <= not(inputs(89));
    layer0_outputs(9115) <= not((inputs(242)) xor (inputs(194)));
    layer0_outputs(9116) <= (inputs(74)) or (inputs(77));
    layer0_outputs(9117) <= not((inputs(177)) or (inputs(85)));
    layer0_outputs(9118) <= (inputs(32)) and not (inputs(223));
    layer0_outputs(9119) <= not((inputs(3)) or (inputs(137)));
    layer0_outputs(9120) <= inputs(103);
    layer0_outputs(9121) <= not(inputs(221));
    layer0_outputs(9122) <= inputs(178);
    layer0_outputs(9123) <= inputs(203);
    layer0_outputs(9124) <= (inputs(142)) xor (inputs(20));
    layer0_outputs(9125) <= not(inputs(129));
    layer0_outputs(9126) <= not((inputs(135)) or (inputs(78)));
    layer0_outputs(9127) <= not(inputs(215)) or (inputs(41));
    layer0_outputs(9128) <= inputs(23);
    layer0_outputs(9129) <= not(inputs(125)) or (inputs(241));
    layer0_outputs(9130) <= (inputs(124)) and (inputs(236));
    layer0_outputs(9131) <= (inputs(13)) xor (inputs(243));
    layer0_outputs(9132) <= not(inputs(105)) or (inputs(149));
    layer0_outputs(9133) <= not(inputs(231)) or (inputs(252));
    layer0_outputs(9134) <= (inputs(52)) and not (inputs(56));
    layer0_outputs(9135) <= not(inputs(54));
    layer0_outputs(9136) <= not(inputs(181)) or (inputs(63));
    layer0_outputs(9137) <= inputs(134);
    layer0_outputs(9138) <= inputs(205);
    layer0_outputs(9139) <= (inputs(213)) and not (inputs(165));
    layer0_outputs(9140) <= (inputs(14)) or (inputs(97));
    layer0_outputs(9141) <= (inputs(204)) xor (inputs(26));
    layer0_outputs(9142) <= not((inputs(48)) or (inputs(122)));
    layer0_outputs(9143) <= (inputs(73)) or (inputs(198));
    layer0_outputs(9144) <= (inputs(144)) xor (inputs(53));
    layer0_outputs(9145) <= not(inputs(67)) or (inputs(54));
    layer0_outputs(9146) <= (inputs(57)) and not (inputs(33));
    layer0_outputs(9147) <= not(inputs(91));
    layer0_outputs(9148) <= (inputs(0)) and not (inputs(138));
    layer0_outputs(9149) <= not(inputs(113));
    layer0_outputs(9150) <= (inputs(146)) xor (inputs(183));
    layer0_outputs(9151) <= not((inputs(87)) or (inputs(86)));
    layer0_outputs(9152) <= inputs(145);
    layer0_outputs(9153) <= inputs(103);
    layer0_outputs(9154) <= not(inputs(39));
    layer0_outputs(9155) <= (inputs(244)) and (inputs(215));
    layer0_outputs(9156) <= not((inputs(74)) xor (inputs(88)));
    layer0_outputs(9157) <= not((inputs(168)) xor (inputs(199)));
    layer0_outputs(9158) <= (inputs(245)) and not (inputs(189));
    layer0_outputs(9159) <= not((inputs(27)) xor (inputs(245)));
    layer0_outputs(9160) <= (inputs(13)) and not (inputs(160));
    layer0_outputs(9161) <= inputs(36);
    layer0_outputs(9162) <= not((inputs(165)) xor (inputs(61)));
    layer0_outputs(9163) <= (inputs(149)) and (inputs(244));
    layer0_outputs(9164) <= not((inputs(132)) xor (inputs(237)));
    layer0_outputs(9165) <= not((inputs(123)) or (inputs(29)));
    layer0_outputs(9166) <= not(inputs(163));
    layer0_outputs(9167) <= (inputs(177)) and not (inputs(177));
    layer0_outputs(9168) <= not(inputs(56)) or (inputs(140));
    layer0_outputs(9169) <= not(inputs(206)) or (inputs(82));
    layer0_outputs(9170) <= not((inputs(139)) or (inputs(153)));
    layer0_outputs(9171) <= not((inputs(160)) and (inputs(193)));
    layer0_outputs(9172) <= not((inputs(251)) xor (inputs(17)));
    layer0_outputs(9173) <= not(inputs(230)) or (inputs(147));
    layer0_outputs(9174) <= not((inputs(180)) or (inputs(191)));
    layer0_outputs(9175) <= (inputs(223)) or (inputs(72));
    layer0_outputs(9176) <= (inputs(155)) or (inputs(225));
    layer0_outputs(9177) <= inputs(60);
    layer0_outputs(9178) <= not(inputs(52)) or (inputs(135));
    layer0_outputs(9179) <= (inputs(152)) or (inputs(62));
    layer0_outputs(9180) <= (inputs(29)) or (inputs(146));
    layer0_outputs(9181) <= not((inputs(76)) xor (inputs(57)));
    layer0_outputs(9182) <= (inputs(167)) and not (inputs(52));
    layer0_outputs(9183) <= not(inputs(134)) or (inputs(200));
    layer0_outputs(9184) <= (inputs(105)) or (inputs(96));
    layer0_outputs(9185) <= (inputs(30)) xor (inputs(188));
    layer0_outputs(9186) <= not(inputs(192)) or (inputs(11));
    layer0_outputs(9187) <= not(inputs(4));
    layer0_outputs(9188) <= not(inputs(142)) or (inputs(6));
    layer0_outputs(9189) <= (inputs(5)) and not (inputs(255));
    layer0_outputs(9190) <= not(inputs(20));
    layer0_outputs(9191) <= inputs(77);
    layer0_outputs(9192) <= not(inputs(233)) or (inputs(110));
    layer0_outputs(9193) <= not((inputs(245)) and (inputs(21)));
    layer0_outputs(9194) <= not((inputs(223)) xor (inputs(143)));
    layer0_outputs(9195) <= not(inputs(248));
    layer0_outputs(9196) <= not(inputs(39));
    layer0_outputs(9197) <= not((inputs(110)) or (inputs(197)));
    layer0_outputs(9198) <= '0';
    layer0_outputs(9199) <= (inputs(63)) or (inputs(216));
    layer0_outputs(9200) <= inputs(133);
    layer0_outputs(9201) <= not((inputs(186)) or (inputs(132)));
    layer0_outputs(9202) <= (inputs(136)) xor (inputs(156));
    layer0_outputs(9203) <= (inputs(177)) xor (inputs(75));
    layer0_outputs(9204) <= not(inputs(218)) or (inputs(107));
    layer0_outputs(9205) <= '0';
    layer0_outputs(9206) <= (inputs(167)) or (inputs(157));
    layer0_outputs(9207) <= (inputs(129)) and (inputs(158));
    layer0_outputs(9208) <= inputs(135);
    layer0_outputs(9209) <= (inputs(172)) or (inputs(203));
    layer0_outputs(9210) <= not(inputs(145));
    layer0_outputs(9211) <= (inputs(233)) xor (inputs(58));
    layer0_outputs(9212) <= not(inputs(117));
    layer0_outputs(9213) <= (inputs(193)) or (inputs(195));
    layer0_outputs(9214) <= not(inputs(151)) or (inputs(109));
    layer0_outputs(9215) <= (inputs(119)) xor (inputs(186));
    layer0_outputs(9216) <= (inputs(218)) xor (inputs(114));
    layer0_outputs(9217) <= not(inputs(228)) or (inputs(49));
    layer0_outputs(9218) <= (inputs(249)) and not (inputs(146));
    layer0_outputs(9219) <= (inputs(94)) and not (inputs(12));
    layer0_outputs(9220) <= (inputs(179)) or (inputs(196));
    layer0_outputs(9221) <= not(inputs(166)) or (inputs(4));
    layer0_outputs(9222) <= not(inputs(183)) or (inputs(54));
    layer0_outputs(9223) <= (inputs(118)) xor (inputs(87));
    layer0_outputs(9224) <= (inputs(82)) and not (inputs(242));
    layer0_outputs(9225) <= (inputs(130)) xor (inputs(167));
    layer0_outputs(9226) <= not((inputs(55)) xor (inputs(11)));
    layer0_outputs(9227) <= inputs(110);
    layer0_outputs(9228) <= not((inputs(116)) or (inputs(157)));
    layer0_outputs(9229) <= (inputs(176)) xor (inputs(18));
    layer0_outputs(9230) <= (inputs(198)) or (inputs(148));
    layer0_outputs(9231) <= not((inputs(110)) xor (inputs(16)));
    layer0_outputs(9232) <= (inputs(48)) and not (inputs(193));
    layer0_outputs(9233) <= (inputs(24)) and (inputs(25));
    layer0_outputs(9234) <= not((inputs(248)) and (inputs(169)));
    layer0_outputs(9235) <= (inputs(130)) xor (inputs(22));
    layer0_outputs(9236) <= not(inputs(105)) or (inputs(17));
    layer0_outputs(9237) <= not(inputs(10));
    layer0_outputs(9238) <= not(inputs(129));
    layer0_outputs(9239) <= not(inputs(181)) or (inputs(144));
    layer0_outputs(9240) <= inputs(89);
    layer0_outputs(9241) <= not((inputs(81)) or (inputs(12)));
    layer0_outputs(9242) <= (inputs(153)) xor (inputs(140));
    layer0_outputs(9243) <= not((inputs(12)) or (inputs(134)));
    layer0_outputs(9244) <= not((inputs(23)) xor (inputs(187)));
    layer0_outputs(9245) <= not(inputs(157)) or (inputs(17));
    layer0_outputs(9246) <= not(inputs(122)) or (inputs(179));
    layer0_outputs(9247) <= (inputs(226)) or (inputs(178));
    layer0_outputs(9248) <= not((inputs(167)) or (inputs(152)));
    layer0_outputs(9249) <= not((inputs(74)) or (inputs(128)));
    layer0_outputs(9250) <= not((inputs(181)) xor (inputs(133)));
    layer0_outputs(9251) <= not((inputs(64)) xor (inputs(90)));
    layer0_outputs(9252) <= (inputs(93)) or (inputs(8));
    layer0_outputs(9253) <= not(inputs(78));
    layer0_outputs(9254) <= not((inputs(211)) xor (inputs(38)));
    layer0_outputs(9255) <= (inputs(63)) or (inputs(86));
    layer0_outputs(9256) <= inputs(107);
    layer0_outputs(9257) <= (inputs(45)) or (inputs(185));
    layer0_outputs(9258) <= (inputs(95)) and (inputs(189));
    layer0_outputs(9259) <= not((inputs(24)) or (inputs(94)));
    layer0_outputs(9260) <= (inputs(168)) or (inputs(250));
    layer0_outputs(9261) <= (inputs(84)) and not (inputs(8));
    layer0_outputs(9262) <= not((inputs(51)) or (inputs(31)));
    layer0_outputs(9263) <= not(inputs(147)) or (inputs(228));
    layer0_outputs(9264) <= (inputs(34)) xor (inputs(7));
    layer0_outputs(9265) <= inputs(155);
    layer0_outputs(9266) <= not(inputs(113));
    layer0_outputs(9267) <= (inputs(154)) and not (inputs(76));
    layer0_outputs(9268) <= (inputs(176)) and (inputs(219));
    layer0_outputs(9269) <= inputs(106);
    layer0_outputs(9270) <= not(inputs(128)) or (inputs(238));
    layer0_outputs(9271) <= not(inputs(231));
    layer0_outputs(9272) <= not(inputs(52));
    layer0_outputs(9273) <= (inputs(151)) and (inputs(85));
    layer0_outputs(9274) <= not(inputs(149));
    layer0_outputs(9275) <= inputs(8);
    layer0_outputs(9276) <= not((inputs(223)) or (inputs(229)));
    layer0_outputs(9277) <= (inputs(67)) or (inputs(185));
    layer0_outputs(9278) <= not(inputs(187));
    layer0_outputs(9279) <= (inputs(41)) or (inputs(80));
    layer0_outputs(9280) <= not(inputs(124));
    layer0_outputs(9281) <= (inputs(191)) or (inputs(88));
    layer0_outputs(9282) <= not(inputs(96));
    layer0_outputs(9283) <= (inputs(242)) and (inputs(70));
    layer0_outputs(9284) <= not((inputs(141)) or (inputs(189)));
    layer0_outputs(9285) <= inputs(162);
    layer0_outputs(9286) <= not(inputs(196));
    layer0_outputs(9287) <= (inputs(217)) and not (inputs(108));
    layer0_outputs(9288) <= inputs(131);
    layer0_outputs(9289) <= not(inputs(67));
    layer0_outputs(9290) <= (inputs(40)) or (inputs(47));
    layer0_outputs(9291) <= inputs(247);
    layer0_outputs(9292) <= inputs(25);
    layer0_outputs(9293) <= (inputs(217)) and not (inputs(96));
    layer0_outputs(9294) <= (inputs(16)) or (inputs(90));
    layer0_outputs(9295) <= inputs(28);
    layer0_outputs(9296) <= (inputs(73)) xor (inputs(71));
    layer0_outputs(9297) <= inputs(12);
    layer0_outputs(9298) <= (inputs(5)) xor (inputs(79));
    layer0_outputs(9299) <= not(inputs(134)) or (inputs(158));
    layer0_outputs(9300) <= (inputs(178)) and not (inputs(47));
    layer0_outputs(9301) <= inputs(135);
    layer0_outputs(9302) <= not(inputs(140));
    layer0_outputs(9303) <= not(inputs(209));
    layer0_outputs(9304) <= inputs(249);
    layer0_outputs(9305) <= not(inputs(173));
    layer0_outputs(9306) <= not((inputs(121)) xor (inputs(180)));
    layer0_outputs(9307) <= inputs(36);
    layer0_outputs(9308) <= not(inputs(249));
    layer0_outputs(9309) <= not(inputs(162));
    layer0_outputs(9310) <= not(inputs(44));
    layer0_outputs(9311) <= not(inputs(165));
    layer0_outputs(9312) <= (inputs(173)) xor (inputs(131));
    layer0_outputs(9313) <= not(inputs(130));
    layer0_outputs(9314) <= (inputs(8)) and not (inputs(74));
    layer0_outputs(9315) <= inputs(22);
    layer0_outputs(9316) <= inputs(109);
    layer0_outputs(9317) <= (inputs(11)) xor (inputs(9));
    layer0_outputs(9318) <= not(inputs(69)) or (inputs(48));
    layer0_outputs(9319) <= not(inputs(70)) or (inputs(62));
    layer0_outputs(9320) <= (inputs(243)) and (inputs(169));
    layer0_outputs(9321) <= (inputs(208)) or (inputs(111));
    layer0_outputs(9322) <= not((inputs(90)) xor (inputs(29)));
    layer0_outputs(9323) <= inputs(17);
    layer0_outputs(9324) <= (inputs(40)) and not (inputs(81));
    layer0_outputs(9325) <= inputs(34);
    layer0_outputs(9326) <= (inputs(54)) or (inputs(180));
    layer0_outputs(9327) <= inputs(126);
    layer0_outputs(9328) <= (inputs(49)) xor (inputs(234));
    layer0_outputs(9329) <= not(inputs(76));
    layer0_outputs(9330) <= not((inputs(70)) or (inputs(112)));
    layer0_outputs(9331) <= '1';
    layer0_outputs(9332) <= not((inputs(196)) and (inputs(100)));
    layer0_outputs(9333) <= (inputs(39)) and not (inputs(88));
    layer0_outputs(9334) <= not((inputs(74)) xor (inputs(215)));
    layer0_outputs(9335) <= not(inputs(200)) or (inputs(201));
    layer0_outputs(9336) <= (inputs(199)) xor (inputs(185));
    layer0_outputs(9337) <= (inputs(42)) or (inputs(14));
    layer0_outputs(9338) <= not((inputs(54)) or (inputs(65)));
    layer0_outputs(9339) <= (inputs(6)) or (inputs(145));
    layer0_outputs(9340) <= (inputs(187)) and not (inputs(10));
    layer0_outputs(9341) <= (inputs(246)) or (inputs(189));
    layer0_outputs(9342) <= (inputs(188)) or (inputs(211));
    layer0_outputs(9343) <= not((inputs(37)) or (inputs(192)));
    layer0_outputs(9344) <= (inputs(219)) xor (inputs(103));
    layer0_outputs(9345) <= (inputs(91)) xor (inputs(218));
    layer0_outputs(9346) <= not(inputs(51)) or (inputs(225));
    layer0_outputs(9347) <= (inputs(225)) xor (inputs(175));
    layer0_outputs(9348) <= not(inputs(138));
    layer0_outputs(9349) <= inputs(39);
    layer0_outputs(9350) <= not(inputs(113));
    layer0_outputs(9351) <= inputs(146);
    layer0_outputs(9352) <= '1';
    layer0_outputs(9353) <= (inputs(121)) and not (inputs(244));
    layer0_outputs(9354) <= (inputs(46)) xor (inputs(73));
    layer0_outputs(9355) <= not(inputs(40)) or (inputs(193));
    layer0_outputs(9356) <= not(inputs(207)) or (inputs(177));
    layer0_outputs(9357) <= inputs(210);
    layer0_outputs(9358) <= (inputs(225)) or (inputs(162));
    layer0_outputs(9359) <= inputs(122);
    layer0_outputs(9360) <= (inputs(89)) and not (inputs(160));
    layer0_outputs(9361) <= not((inputs(245)) or (inputs(235)));
    layer0_outputs(9362) <= not((inputs(174)) or (inputs(199)));
    layer0_outputs(9363) <= (inputs(34)) xor (inputs(235));
    layer0_outputs(9364) <= not(inputs(206));
    layer0_outputs(9365) <= inputs(45);
    layer0_outputs(9366) <= (inputs(51)) or (inputs(207));
    layer0_outputs(9367) <= not((inputs(7)) xor (inputs(79)));
    layer0_outputs(9368) <= not(inputs(160));
    layer0_outputs(9369) <= not(inputs(78));
    layer0_outputs(9370) <= inputs(62);
    layer0_outputs(9371) <= not((inputs(164)) and (inputs(186)));
    layer0_outputs(9372) <= not((inputs(53)) xor (inputs(51)));
    layer0_outputs(9373) <= inputs(148);
    layer0_outputs(9374) <= not((inputs(126)) or (inputs(1)));
    layer0_outputs(9375) <= (inputs(132)) and (inputs(72));
    layer0_outputs(9376) <= not(inputs(186)) or (inputs(48));
    layer0_outputs(9377) <= not((inputs(33)) xor (inputs(49)));
    layer0_outputs(9378) <= inputs(197);
    layer0_outputs(9379) <= inputs(230);
    layer0_outputs(9380) <= not((inputs(241)) xor (inputs(46)));
    layer0_outputs(9381) <= (inputs(142)) or (inputs(112));
    layer0_outputs(9382) <= not(inputs(68)) or (inputs(173));
    layer0_outputs(9383) <= not(inputs(212));
    layer0_outputs(9384) <= (inputs(47)) or (inputs(60));
    layer0_outputs(9385) <= not((inputs(13)) and (inputs(12)));
    layer0_outputs(9386) <= (inputs(18)) and not (inputs(175));
    layer0_outputs(9387) <= (inputs(78)) xor (inputs(127));
    layer0_outputs(9388) <= (inputs(106)) and not (inputs(232));
    layer0_outputs(9389) <= not((inputs(183)) or (inputs(64)));
    layer0_outputs(9390) <= inputs(179);
    layer0_outputs(9391) <= inputs(198);
    layer0_outputs(9392) <= inputs(14);
    layer0_outputs(9393) <= (inputs(168)) xor (inputs(179));
    layer0_outputs(9394) <= not((inputs(11)) or (inputs(104)));
    layer0_outputs(9395) <= not((inputs(181)) or (inputs(239)));
    layer0_outputs(9396) <= (inputs(9)) and not (inputs(15));
    layer0_outputs(9397) <= (inputs(48)) or (inputs(172));
    layer0_outputs(9398) <= '1';
    layer0_outputs(9399) <= '1';
    layer0_outputs(9400) <= inputs(209);
    layer0_outputs(9401) <= not(inputs(245)) or (inputs(20));
    layer0_outputs(9402) <= not((inputs(4)) xor (inputs(118)));
    layer0_outputs(9403) <= (inputs(12)) or (inputs(195));
    layer0_outputs(9404) <= (inputs(135)) and not (inputs(110));
    layer0_outputs(9405) <= (inputs(46)) or (inputs(190));
    layer0_outputs(9406) <= not((inputs(144)) xor (inputs(164)));
    layer0_outputs(9407) <= (inputs(183)) and not (inputs(117));
    layer0_outputs(9408) <= (inputs(131)) and not (inputs(250));
    layer0_outputs(9409) <= not(inputs(105));
    layer0_outputs(9410) <= not((inputs(6)) xor (inputs(69)));
    layer0_outputs(9411) <= inputs(93);
    layer0_outputs(9412) <= not((inputs(191)) xor (inputs(180)));
    layer0_outputs(9413) <= not(inputs(145));
    layer0_outputs(9414) <= not(inputs(36));
    layer0_outputs(9415) <= not(inputs(97));
    layer0_outputs(9416) <= not(inputs(183)) or (inputs(140));
    layer0_outputs(9417) <= (inputs(242)) xor (inputs(124));
    layer0_outputs(9418) <= (inputs(86)) and not (inputs(94));
    layer0_outputs(9419) <= not((inputs(6)) or (inputs(17)));
    layer0_outputs(9420) <= inputs(78);
    layer0_outputs(9421) <= (inputs(190)) and not (inputs(191));
    layer0_outputs(9422) <= not(inputs(8));
    layer0_outputs(9423) <= not((inputs(44)) xor (inputs(59)));
    layer0_outputs(9424) <= inputs(88);
    layer0_outputs(9425) <= (inputs(49)) and not (inputs(138));
    layer0_outputs(9426) <= not(inputs(85));
    layer0_outputs(9427) <= not((inputs(251)) or (inputs(228)));
    layer0_outputs(9428) <= not(inputs(110)) or (inputs(32));
    layer0_outputs(9429) <= inputs(232);
    layer0_outputs(9430) <= not((inputs(98)) xor (inputs(194)));
    layer0_outputs(9431) <= not(inputs(37)) or (inputs(180));
    layer0_outputs(9432) <= not(inputs(123)) or (inputs(151));
    layer0_outputs(9433) <= not((inputs(46)) or (inputs(248)));
    layer0_outputs(9434) <= not(inputs(236));
    layer0_outputs(9435) <= not(inputs(110));
    layer0_outputs(9436) <= (inputs(207)) or (inputs(79));
    layer0_outputs(9437) <= not((inputs(224)) or (inputs(247)));
    layer0_outputs(9438) <= (inputs(201)) or (inputs(17));
    layer0_outputs(9439) <= (inputs(60)) xor (inputs(91));
    layer0_outputs(9440) <= inputs(34);
    layer0_outputs(9441) <= (inputs(238)) xor (inputs(131));
    layer0_outputs(9442) <= (inputs(99)) xor (inputs(227));
    layer0_outputs(9443) <= not((inputs(120)) or (inputs(135)));
    layer0_outputs(9444) <= not((inputs(57)) xor (inputs(173)));
    layer0_outputs(9445) <= (inputs(36)) and not (inputs(156));
    layer0_outputs(9446) <= not(inputs(2)) or (inputs(86));
    layer0_outputs(9447) <= (inputs(180)) or (inputs(245));
    layer0_outputs(9448) <= not((inputs(113)) xor (inputs(84)));
    layer0_outputs(9449) <= not((inputs(108)) or (inputs(16)));
    layer0_outputs(9450) <= (inputs(250)) and not (inputs(11));
    layer0_outputs(9451) <= not(inputs(114)) or (inputs(80));
    layer0_outputs(9452) <= not((inputs(193)) or (inputs(244)));
    layer0_outputs(9453) <= (inputs(154)) and not (inputs(5));
    layer0_outputs(9454) <= not(inputs(15));
    layer0_outputs(9455) <= not(inputs(25));
    layer0_outputs(9456) <= inputs(88);
    layer0_outputs(9457) <= not(inputs(59));
    layer0_outputs(9458) <= not((inputs(171)) or (inputs(27)));
    layer0_outputs(9459) <= not((inputs(32)) or (inputs(17)));
    layer0_outputs(9460) <= inputs(118);
    layer0_outputs(9461) <= inputs(25);
    layer0_outputs(9462) <= (inputs(22)) xor (inputs(9));
    layer0_outputs(9463) <= not(inputs(231));
    layer0_outputs(9464) <= (inputs(243)) or (inputs(9));
    layer0_outputs(9465) <= inputs(25);
    layer0_outputs(9466) <= inputs(102);
    layer0_outputs(9467) <= '1';
    layer0_outputs(9468) <= inputs(81);
    layer0_outputs(9469) <= (inputs(156)) and not (inputs(127));
    layer0_outputs(9470) <= not((inputs(10)) or (inputs(125)));
    layer0_outputs(9471) <= inputs(53);
    layer0_outputs(9472) <= not(inputs(189));
    layer0_outputs(9473) <= (inputs(211)) xor (inputs(198));
    layer0_outputs(9474) <= (inputs(235)) and (inputs(5));
    layer0_outputs(9475) <= inputs(232);
    layer0_outputs(9476) <= inputs(84);
    layer0_outputs(9477) <= not(inputs(112));
    layer0_outputs(9478) <= (inputs(47)) or (inputs(31));
    layer0_outputs(9479) <= not(inputs(89)) or (inputs(115));
    layer0_outputs(9480) <= not(inputs(164));
    layer0_outputs(9481) <= not(inputs(248));
    layer0_outputs(9482) <= not(inputs(128));
    layer0_outputs(9483) <= inputs(217);
    layer0_outputs(9484) <= not((inputs(113)) xor (inputs(244)));
    layer0_outputs(9485) <= not(inputs(44)) or (inputs(95));
    layer0_outputs(9486) <= not((inputs(44)) and (inputs(159)));
    layer0_outputs(9487) <= '0';
    layer0_outputs(9488) <= not(inputs(250));
    layer0_outputs(9489) <= inputs(87);
    layer0_outputs(9490) <= not(inputs(124));
    layer0_outputs(9491) <= inputs(71);
    layer0_outputs(9492) <= (inputs(88)) and not (inputs(36));
    layer0_outputs(9493) <= not((inputs(78)) xor (inputs(76)));
    layer0_outputs(9494) <= (inputs(131)) and not (inputs(192));
    layer0_outputs(9495) <= not(inputs(187));
    layer0_outputs(9496) <= not(inputs(42)) or (inputs(80));
    layer0_outputs(9497) <= not(inputs(122));
    layer0_outputs(9498) <= not((inputs(222)) or (inputs(221)));
    layer0_outputs(9499) <= not((inputs(20)) and (inputs(187)));
    layer0_outputs(9500) <= (inputs(177)) or (inputs(213));
    layer0_outputs(9501) <= (inputs(4)) or (inputs(168));
    layer0_outputs(9502) <= (inputs(236)) and not (inputs(32));
    layer0_outputs(9503) <= not(inputs(107));
    layer0_outputs(9504) <= (inputs(218)) and not (inputs(133));
    layer0_outputs(9505) <= not(inputs(120));
    layer0_outputs(9506) <= not((inputs(226)) or (inputs(212)));
    layer0_outputs(9507) <= (inputs(169)) and not (inputs(117));
    layer0_outputs(9508) <= not((inputs(72)) or (inputs(170)));
    layer0_outputs(9509) <= (inputs(93)) xor (inputs(106));
    layer0_outputs(9510) <= inputs(124);
    layer0_outputs(9511) <= (inputs(27)) xor (inputs(91));
    layer0_outputs(9512) <= (inputs(167)) or (inputs(210));
    layer0_outputs(9513) <= not(inputs(60)) or (inputs(205));
    layer0_outputs(9514) <= not((inputs(233)) or (inputs(88)));
    layer0_outputs(9515) <= inputs(16);
    layer0_outputs(9516) <= (inputs(75)) and not (inputs(159));
    layer0_outputs(9517) <= not((inputs(71)) or (inputs(64)));
    layer0_outputs(9518) <= not(inputs(25));
    layer0_outputs(9519) <= not((inputs(104)) or (inputs(218)));
    layer0_outputs(9520) <= (inputs(139)) and not (inputs(0));
    layer0_outputs(9521) <= '1';
    layer0_outputs(9522) <= not((inputs(167)) or (inputs(243)));
    layer0_outputs(9523) <= '1';
    layer0_outputs(9524) <= not((inputs(150)) or (inputs(189)));
    layer0_outputs(9525) <= not((inputs(60)) xor (inputs(145)));
    layer0_outputs(9526) <= not(inputs(61));
    layer0_outputs(9527) <= not(inputs(60)) or (inputs(80));
    layer0_outputs(9528) <= not((inputs(228)) and (inputs(226)));
    layer0_outputs(9529) <= not(inputs(65)) or (inputs(111));
    layer0_outputs(9530) <= not((inputs(99)) or (inputs(46)));
    layer0_outputs(9531) <= not((inputs(23)) xor (inputs(243)));
    layer0_outputs(9532) <= not(inputs(60)) or (inputs(2));
    layer0_outputs(9533) <= not(inputs(159)) or (inputs(12));
    layer0_outputs(9534) <= (inputs(208)) or (inputs(248));
    layer0_outputs(9535) <= not(inputs(85));
    layer0_outputs(9536) <= (inputs(240)) and not (inputs(90));
    layer0_outputs(9537) <= '1';
    layer0_outputs(9538) <= (inputs(214)) or (inputs(176));
    layer0_outputs(9539) <= (inputs(18)) and not (inputs(79));
    layer0_outputs(9540) <= not(inputs(99));
    layer0_outputs(9541) <= (inputs(76)) and (inputs(10));
    layer0_outputs(9542) <= not(inputs(213));
    layer0_outputs(9543) <= not((inputs(183)) xor (inputs(69)));
    layer0_outputs(9544) <= (inputs(177)) xor (inputs(3));
    layer0_outputs(9545) <= not((inputs(168)) or (inputs(113)));
    layer0_outputs(9546) <= not(inputs(4));
    layer0_outputs(9547) <= not(inputs(212)) or (inputs(38));
    layer0_outputs(9548) <= not((inputs(113)) or (inputs(27)));
    layer0_outputs(9549) <= (inputs(226)) xor (inputs(243));
    layer0_outputs(9550) <= not(inputs(93));
    layer0_outputs(9551) <= not(inputs(107));
    layer0_outputs(9552) <= (inputs(61)) or (inputs(236));
    layer0_outputs(9553) <= not(inputs(13));
    layer0_outputs(9554) <= not(inputs(172));
    layer0_outputs(9555) <= inputs(130);
    layer0_outputs(9556) <= (inputs(102)) and not (inputs(226));
    layer0_outputs(9557) <= inputs(92);
    layer0_outputs(9558) <= not(inputs(104)) or (inputs(68));
    layer0_outputs(9559) <= not(inputs(152));
    layer0_outputs(9560) <= not(inputs(235));
    layer0_outputs(9561) <= not(inputs(216));
    layer0_outputs(9562) <= not(inputs(65));
    layer0_outputs(9563) <= (inputs(108)) and not (inputs(225));
    layer0_outputs(9564) <= not(inputs(191)) or (inputs(27));
    layer0_outputs(9565) <= not(inputs(242));
    layer0_outputs(9566) <= (inputs(24)) xor (inputs(55));
    layer0_outputs(9567) <= (inputs(116)) or (inputs(119));
    layer0_outputs(9568) <= not((inputs(192)) xor (inputs(151)));
    layer0_outputs(9569) <= (inputs(162)) or (inputs(216));
    layer0_outputs(9570) <= inputs(102);
    layer0_outputs(9571) <= not((inputs(167)) or (inputs(238)));
    layer0_outputs(9572) <= not((inputs(158)) xor (inputs(117)));
    layer0_outputs(9573) <= '1';
    layer0_outputs(9574) <= not((inputs(93)) or (inputs(183)));
    layer0_outputs(9575) <= not(inputs(118));
    layer0_outputs(9576) <= not((inputs(190)) or (inputs(63)));
    layer0_outputs(9577) <= not((inputs(224)) or (inputs(213)));
    layer0_outputs(9578) <= not((inputs(97)) xor (inputs(147)));
    layer0_outputs(9579) <= (inputs(121)) or (inputs(239));
    layer0_outputs(9580) <= not((inputs(164)) xor (inputs(195)));
    layer0_outputs(9581) <= (inputs(192)) xor (inputs(174));
    layer0_outputs(9582) <= not((inputs(222)) or (inputs(25)));
    layer0_outputs(9583) <= not((inputs(99)) xor (inputs(121)));
    layer0_outputs(9584) <= '0';
    layer0_outputs(9585) <= not(inputs(7)) or (inputs(71));
    layer0_outputs(9586) <= (inputs(73)) and not (inputs(255));
    layer0_outputs(9587) <= not((inputs(6)) xor (inputs(133)));
    layer0_outputs(9588) <= not((inputs(67)) or (inputs(77)));
    layer0_outputs(9589) <= not(inputs(104)) or (inputs(251));
    layer0_outputs(9590) <= not(inputs(210)) or (inputs(163));
    layer0_outputs(9591) <= inputs(214);
    layer0_outputs(9592) <= not(inputs(146));
    layer0_outputs(9593) <= not(inputs(117)) or (inputs(139));
    layer0_outputs(9594) <= not((inputs(23)) xor (inputs(231)));
    layer0_outputs(9595) <= inputs(113);
    layer0_outputs(9596) <= not(inputs(22));
    layer0_outputs(9597) <= (inputs(195)) xor (inputs(199));
    layer0_outputs(9598) <= '0';
    layer0_outputs(9599) <= (inputs(121)) xor (inputs(231));
    layer0_outputs(9600) <= not(inputs(39));
    layer0_outputs(9601) <= (inputs(40)) and not (inputs(222));
    layer0_outputs(9602) <= (inputs(138)) and not (inputs(179));
    layer0_outputs(9603) <= (inputs(94)) and not (inputs(255));
    layer0_outputs(9604) <= not(inputs(86));
    layer0_outputs(9605) <= inputs(19);
    layer0_outputs(9606) <= not((inputs(105)) or (inputs(62)));
    layer0_outputs(9607) <= not((inputs(56)) xor (inputs(168)));
    layer0_outputs(9608) <= (inputs(11)) or (inputs(108));
    layer0_outputs(9609) <= (inputs(20)) xor (inputs(78));
    layer0_outputs(9610) <= not(inputs(74));
    layer0_outputs(9611) <= not((inputs(108)) xor (inputs(6)));
    layer0_outputs(9612) <= not(inputs(39));
    layer0_outputs(9613) <= inputs(74);
    layer0_outputs(9614) <= not(inputs(237)) or (inputs(251));
    layer0_outputs(9615) <= (inputs(51)) xor (inputs(98));
    layer0_outputs(9616) <= (inputs(85)) or (inputs(82));
    layer0_outputs(9617) <= (inputs(255)) or (inputs(122));
    layer0_outputs(9618) <= not(inputs(163));
    layer0_outputs(9619) <= inputs(92);
    layer0_outputs(9620) <= (inputs(64)) and (inputs(211));
    layer0_outputs(9621) <= not((inputs(92)) xor (inputs(32)));
    layer0_outputs(9622) <= inputs(157);
    layer0_outputs(9623) <= (inputs(162)) and not (inputs(34));
    layer0_outputs(9624) <= not((inputs(254)) or (inputs(201)));
    layer0_outputs(9625) <= (inputs(29)) and not (inputs(117));
    layer0_outputs(9626) <= (inputs(183)) and (inputs(185));
    layer0_outputs(9627) <= not((inputs(169)) xor (inputs(150)));
    layer0_outputs(9628) <= not((inputs(80)) xor (inputs(19)));
    layer0_outputs(9629) <= not(inputs(229));
    layer0_outputs(9630) <= (inputs(27)) and not (inputs(200));
    layer0_outputs(9631) <= not(inputs(161));
    layer0_outputs(9632) <= not(inputs(21)) or (inputs(160));
    layer0_outputs(9633) <= inputs(57);
    layer0_outputs(9634) <= not(inputs(144));
    layer0_outputs(9635) <= not((inputs(87)) or (inputs(105)));
    layer0_outputs(9636) <= inputs(147);
    layer0_outputs(9637) <= not((inputs(147)) or (inputs(208)));
    layer0_outputs(9638) <= not(inputs(135));
    layer0_outputs(9639) <= (inputs(215)) and not (inputs(76));
    layer0_outputs(9640) <= (inputs(50)) xor (inputs(238));
    layer0_outputs(9641) <= (inputs(16)) or (inputs(59));
    layer0_outputs(9642) <= inputs(217);
    layer0_outputs(9643) <= inputs(68);
    layer0_outputs(9644) <= not((inputs(7)) xor (inputs(88)));
    layer0_outputs(9645) <= not((inputs(180)) xor (inputs(135)));
    layer0_outputs(9646) <= (inputs(220)) or (inputs(186));
    layer0_outputs(9647) <= (inputs(8)) or (inputs(48));
    layer0_outputs(9648) <= not(inputs(161)) or (inputs(47));
    layer0_outputs(9649) <= inputs(73);
    layer0_outputs(9650) <= not(inputs(119));
    layer0_outputs(9651) <= not((inputs(255)) or (inputs(31)));
    layer0_outputs(9652) <= not((inputs(28)) xor (inputs(251)));
    layer0_outputs(9653) <= not(inputs(220));
    layer0_outputs(9654) <= inputs(101);
    layer0_outputs(9655) <= (inputs(112)) or (inputs(183));
    layer0_outputs(9656) <= (inputs(3)) and not (inputs(53));
    layer0_outputs(9657) <= not(inputs(104)) or (inputs(212));
    layer0_outputs(9658) <= (inputs(253)) or (inputs(232));
    layer0_outputs(9659) <= (inputs(64)) or (inputs(152));
    layer0_outputs(9660) <= inputs(44);
    layer0_outputs(9661) <= not((inputs(185)) or (inputs(187)));
    layer0_outputs(9662) <= (inputs(97)) xor (inputs(74));
    layer0_outputs(9663) <= inputs(26);
    layer0_outputs(9664) <= not(inputs(117));
    layer0_outputs(9665) <= not((inputs(58)) or (inputs(24)));
    layer0_outputs(9666) <= (inputs(37)) and not (inputs(237));
    layer0_outputs(9667) <= not((inputs(251)) or (inputs(252)));
    layer0_outputs(9668) <= (inputs(159)) and not (inputs(111));
    layer0_outputs(9669) <= not(inputs(82)) or (inputs(16));
    layer0_outputs(9670) <= inputs(37);
    layer0_outputs(9671) <= (inputs(243)) or (inputs(98));
    layer0_outputs(9672) <= not((inputs(35)) and (inputs(36)));
    layer0_outputs(9673) <= (inputs(237)) and not (inputs(143));
    layer0_outputs(9674) <= (inputs(231)) and not (inputs(41));
    layer0_outputs(9675) <= inputs(185);
    layer0_outputs(9676) <= not((inputs(246)) and (inputs(75)));
    layer0_outputs(9677) <= not((inputs(8)) or (inputs(174)));
    layer0_outputs(9678) <= not((inputs(207)) or (inputs(200)));
    layer0_outputs(9679) <= (inputs(249)) or (inputs(114));
    layer0_outputs(9680) <= not((inputs(36)) xor (inputs(92)));
    layer0_outputs(9681) <= inputs(23);
    layer0_outputs(9682) <= (inputs(252)) or (inputs(164));
    layer0_outputs(9683) <= not(inputs(168)) or (inputs(24));
    layer0_outputs(9684) <= inputs(124);
    layer0_outputs(9685) <= (inputs(253)) or (inputs(133));
    layer0_outputs(9686) <= not((inputs(10)) or (inputs(5)));
    layer0_outputs(9687) <= not(inputs(162)) or (inputs(96));
    layer0_outputs(9688) <= not(inputs(167));
    layer0_outputs(9689) <= inputs(180);
    layer0_outputs(9690) <= not(inputs(203));
    layer0_outputs(9691) <= not((inputs(21)) and (inputs(113)));
    layer0_outputs(9692) <= inputs(107);
    layer0_outputs(9693) <= inputs(230);
    layer0_outputs(9694) <= (inputs(5)) and not (inputs(0));
    layer0_outputs(9695) <= (inputs(7)) and not (inputs(147));
    layer0_outputs(9696) <= not((inputs(137)) xor (inputs(119)));
    layer0_outputs(9697) <= inputs(35);
    layer0_outputs(9698) <= not(inputs(180)) or (inputs(33));
    layer0_outputs(9699) <= not((inputs(24)) and (inputs(90)));
    layer0_outputs(9700) <= (inputs(162)) xor (inputs(147));
    layer0_outputs(9701) <= inputs(59);
    layer0_outputs(9702) <= inputs(44);
    layer0_outputs(9703) <= not(inputs(226));
    layer0_outputs(9704) <= not(inputs(183)) or (inputs(133));
    layer0_outputs(9705) <= not((inputs(62)) or (inputs(214)));
    layer0_outputs(9706) <= (inputs(4)) xor (inputs(101));
    layer0_outputs(9707) <= inputs(166);
    layer0_outputs(9708) <= not(inputs(188)) or (inputs(47));
    layer0_outputs(9709) <= inputs(9);
    layer0_outputs(9710) <= (inputs(1)) xor (inputs(136));
    layer0_outputs(9711) <= not(inputs(17));
    layer0_outputs(9712) <= not(inputs(198)) or (inputs(191));
    layer0_outputs(9713) <= not(inputs(162));
    layer0_outputs(9714) <= '1';
    layer0_outputs(9715) <= (inputs(215)) and not (inputs(254));
    layer0_outputs(9716) <= not(inputs(79));
    layer0_outputs(9717) <= not(inputs(18));
    layer0_outputs(9718) <= not(inputs(27));
    layer0_outputs(9719) <= inputs(117);
    layer0_outputs(9720) <= inputs(104);
    layer0_outputs(9721) <= not(inputs(221));
    layer0_outputs(9722) <= not((inputs(40)) or (inputs(174)));
    layer0_outputs(9723) <= not((inputs(2)) and (inputs(109)));
    layer0_outputs(9724) <= inputs(126);
    layer0_outputs(9725) <= not(inputs(141));
    layer0_outputs(9726) <= (inputs(38)) or (inputs(212));
    layer0_outputs(9727) <= (inputs(49)) or (inputs(231));
    layer0_outputs(9728) <= (inputs(92)) and not (inputs(179));
    layer0_outputs(9729) <= not((inputs(50)) xor (inputs(47)));
    layer0_outputs(9730) <= not(inputs(41)) or (inputs(164));
    layer0_outputs(9731) <= (inputs(166)) or (inputs(149));
    layer0_outputs(9732) <= not(inputs(236));
    layer0_outputs(9733) <= (inputs(22)) and (inputs(228));
    layer0_outputs(9734) <= not(inputs(182));
    layer0_outputs(9735) <= (inputs(89)) xor (inputs(107));
    layer0_outputs(9736) <= (inputs(242)) or (inputs(176));
    layer0_outputs(9737) <= (inputs(8)) and not (inputs(128));
    layer0_outputs(9738) <= (inputs(180)) and not (inputs(159));
    layer0_outputs(9739) <= not(inputs(236)) or (inputs(139));
    layer0_outputs(9740) <= not((inputs(199)) or (inputs(252)));
    layer0_outputs(9741) <= not(inputs(200));
    layer0_outputs(9742) <= inputs(130);
    layer0_outputs(9743) <= inputs(158);
    layer0_outputs(9744) <= not(inputs(178));
    layer0_outputs(9745) <= not((inputs(118)) or (inputs(225)));
    layer0_outputs(9746) <= '1';
    layer0_outputs(9747) <= (inputs(140)) and not (inputs(237));
    layer0_outputs(9748) <= not(inputs(98)) or (inputs(123));
    layer0_outputs(9749) <= (inputs(232)) and not (inputs(64));
    layer0_outputs(9750) <= not((inputs(185)) xor (inputs(134)));
    layer0_outputs(9751) <= (inputs(171)) and not (inputs(45));
    layer0_outputs(9752) <= not((inputs(173)) xor (inputs(187)));
    layer0_outputs(9753) <= (inputs(150)) or (inputs(83));
    layer0_outputs(9754) <= (inputs(225)) or (inputs(148));
    layer0_outputs(9755) <= inputs(198);
    layer0_outputs(9756) <= (inputs(7)) or (inputs(204));
    layer0_outputs(9757) <= not((inputs(156)) or (inputs(145)));
    layer0_outputs(9758) <= not((inputs(75)) or (inputs(21)));
    layer0_outputs(9759) <= inputs(163);
    layer0_outputs(9760) <= inputs(231);
    layer0_outputs(9761) <= not((inputs(221)) xor (inputs(249)));
    layer0_outputs(9762) <= not((inputs(62)) or (inputs(48)));
    layer0_outputs(9763) <= not(inputs(163)) or (inputs(74));
    layer0_outputs(9764) <= not(inputs(36)) or (inputs(216));
    layer0_outputs(9765) <= (inputs(190)) xor (inputs(32));
    layer0_outputs(9766) <= (inputs(235)) or (inputs(251));
    layer0_outputs(9767) <= not((inputs(127)) or (inputs(219)));
    layer0_outputs(9768) <= inputs(81);
    layer0_outputs(9769) <= inputs(132);
    layer0_outputs(9770) <= (inputs(146)) xor (inputs(238));
    layer0_outputs(9771) <= (inputs(18)) or (inputs(181));
    layer0_outputs(9772) <= not((inputs(11)) xor (inputs(31)));
    layer0_outputs(9773) <= (inputs(46)) or (inputs(177));
    layer0_outputs(9774) <= inputs(59);
    layer0_outputs(9775) <= inputs(27);
    layer0_outputs(9776) <= not(inputs(237)) or (inputs(241));
    layer0_outputs(9777) <= not(inputs(27)) or (inputs(163));
    layer0_outputs(9778) <= not(inputs(226)) or (inputs(120));
    layer0_outputs(9779) <= inputs(81);
    layer0_outputs(9780) <= inputs(88);
    layer0_outputs(9781) <= (inputs(103)) and not (inputs(206));
    layer0_outputs(9782) <= (inputs(66)) or (inputs(163));
    layer0_outputs(9783) <= (inputs(89)) xor (inputs(222));
    layer0_outputs(9784) <= not(inputs(229));
    layer0_outputs(9785) <= (inputs(158)) and (inputs(189));
    layer0_outputs(9786) <= (inputs(246)) or (inputs(128));
    layer0_outputs(9787) <= (inputs(12)) and not (inputs(157));
    layer0_outputs(9788) <= (inputs(126)) and not (inputs(219));
    layer0_outputs(9789) <= not((inputs(82)) xor (inputs(85)));
    layer0_outputs(9790) <= not(inputs(105)) or (inputs(22));
    layer0_outputs(9791) <= not(inputs(186)) or (inputs(43));
    layer0_outputs(9792) <= inputs(25);
    layer0_outputs(9793) <= (inputs(132)) or (inputs(246));
    layer0_outputs(9794) <= not(inputs(172));
    layer0_outputs(9795) <= not(inputs(241));
    layer0_outputs(9796) <= not(inputs(173));
    layer0_outputs(9797) <= not(inputs(153));
    layer0_outputs(9798) <= (inputs(152)) or (inputs(144));
    layer0_outputs(9799) <= not((inputs(128)) and (inputs(143)));
    layer0_outputs(9800) <= not(inputs(248));
    layer0_outputs(9801) <= inputs(186);
    layer0_outputs(9802) <= not(inputs(63));
    layer0_outputs(9803) <= not(inputs(229)) or (inputs(175));
    layer0_outputs(9804) <= not(inputs(210)) or (inputs(239));
    layer0_outputs(9805) <= not((inputs(121)) or (inputs(106)));
    layer0_outputs(9806) <= inputs(163);
    layer0_outputs(9807) <= inputs(231);
    layer0_outputs(9808) <= not(inputs(111));
    layer0_outputs(9809) <= not(inputs(74)) or (inputs(164));
    layer0_outputs(9810) <= inputs(75);
    layer0_outputs(9811) <= (inputs(87)) or (inputs(242));
    layer0_outputs(9812) <= (inputs(160)) or (inputs(38));
    layer0_outputs(9813) <= not((inputs(216)) xor (inputs(111)));
    layer0_outputs(9814) <= not((inputs(155)) xor (inputs(198)));
    layer0_outputs(9815) <= inputs(181);
    layer0_outputs(9816) <= not(inputs(165));
    layer0_outputs(9817) <= not(inputs(142));
    layer0_outputs(9818) <= not((inputs(117)) and (inputs(201)));
    layer0_outputs(9819) <= not(inputs(227));
    layer0_outputs(9820) <= not((inputs(24)) xor (inputs(21)));
    layer0_outputs(9821) <= (inputs(207)) xor (inputs(77));
    layer0_outputs(9822) <= not((inputs(194)) or (inputs(175)));
    layer0_outputs(9823) <= not(inputs(46));
    layer0_outputs(9824) <= not(inputs(39)) or (inputs(26));
    layer0_outputs(9825) <= (inputs(141)) and (inputs(235));
    layer0_outputs(9826) <= not((inputs(4)) xor (inputs(254)));
    layer0_outputs(9827) <= not((inputs(102)) xor (inputs(175)));
    layer0_outputs(9828) <= (inputs(37)) and not (inputs(220));
    layer0_outputs(9829) <= (inputs(88)) xor (inputs(23));
    layer0_outputs(9830) <= (inputs(110)) and not (inputs(136));
    layer0_outputs(9831) <= not(inputs(202));
    layer0_outputs(9832) <= not(inputs(86));
    layer0_outputs(9833) <= (inputs(164)) or (inputs(80));
    layer0_outputs(9834) <= (inputs(177)) or (inputs(81));
    layer0_outputs(9835) <= inputs(57);
    layer0_outputs(9836) <= not((inputs(70)) and (inputs(214)));
    layer0_outputs(9837) <= (inputs(63)) or (inputs(226));
    layer0_outputs(9838) <= (inputs(141)) and not (inputs(155));
    layer0_outputs(9839) <= not((inputs(195)) or (inputs(68)));
    layer0_outputs(9840) <= not(inputs(75)) or (inputs(34));
    layer0_outputs(9841) <= not(inputs(78));
    layer0_outputs(9842) <= inputs(214);
    layer0_outputs(9843) <= (inputs(228)) xor (inputs(143));
    layer0_outputs(9844) <= inputs(76);
    layer0_outputs(9845) <= (inputs(228)) and not (inputs(5));
    layer0_outputs(9846) <= inputs(26);
    layer0_outputs(9847) <= (inputs(108)) or (inputs(9));
    layer0_outputs(9848) <= inputs(121);
    layer0_outputs(9849) <= (inputs(61)) or (inputs(197));
    layer0_outputs(9850) <= (inputs(112)) or (inputs(172));
    layer0_outputs(9851) <= not((inputs(195)) and (inputs(10)));
    layer0_outputs(9852) <= (inputs(176)) and not (inputs(64));
    layer0_outputs(9853) <= not(inputs(158));
    layer0_outputs(9854) <= (inputs(187)) or (inputs(88));
    layer0_outputs(9855) <= inputs(22);
    layer0_outputs(9856) <= not(inputs(108));
    layer0_outputs(9857) <= not((inputs(150)) or (inputs(10)));
    layer0_outputs(9858) <= not((inputs(162)) or (inputs(146)));
    layer0_outputs(9859) <= inputs(37);
    layer0_outputs(9860) <= '1';
    layer0_outputs(9861) <= (inputs(87)) and (inputs(170));
    layer0_outputs(9862) <= (inputs(106)) and not (inputs(158));
    layer0_outputs(9863) <= not(inputs(82)) or (inputs(75));
    layer0_outputs(9864) <= not(inputs(221));
    layer0_outputs(9865) <= (inputs(24)) and not (inputs(236));
    layer0_outputs(9866) <= (inputs(242)) xor (inputs(180));
    layer0_outputs(9867) <= not(inputs(103));
    layer0_outputs(9868) <= not((inputs(221)) or (inputs(192)));
    layer0_outputs(9869) <= inputs(233);
    layer0_outputs(9870) <= not((inputs(129)) xor (inputs(102)));
    layer0_outputs(9871) <= not(inputs(100));
    layer0_outputs(9872) <= not(inputs(218));
    layer0_outputs(9873) <= inputs(117);
    layer0_outputs(9874) <= (inputs(178)) or (inputs(159));
    layer0_outputs(9875) <= (inputs(247)) and not (inputs(106));
    layer0_outputs(9876) <= not(inputs(186));
    layer0_outputs(9877) <= not(inputs(85));
    layer0_outputs(9878) <= (inputs(166)) and not (inputs(176));
    layer0_outputs(9879) <= (inputs(86)) xor (inputs(36));
    layer0_outputs(9880) <= not((inputs(65)) and (inputs(32)));
    layer0_outputs(9881) <= (inputs(64)) xor (inputs(161));
    layer0_outputs(9882) <= not(inputs(35)) or (inputs(100));
    layer0_outputs(9883) <= (inputs(112)) or (inputs(97));
    layer0_outputs(9884) <= not((inputs(171)) or (inputs(85)));
    layer0_outputs(9885) <= not((inputs(187)) xor (inputs(101)));
    layer0_outputs(9886) <= not(inputs(142));
    layer0_outputs(9887) <= not(inputs(119));
    layer0_outputs(9888) <= not(inputs(150));
    layer0_outputs(9889) <= '0';
    layer0_outputs(9890) <= inputs(133);
    layer0_outputs(9891) <= (inputs(193)) and not (inputs(2));
    layer0_outputs(9892) <= not(inputs(85));
    layer0_outputs(9893) <= not(inputs(113)) or (inputs(4));
    layer0_outputs(9894) <= not((inputs(191)) or (inputs(182)));
    layer0_outputs(9895) <= not((inputs(38)) and (inputs(99)));
    layer0_outputs(9896) <= not(inputs(93)) or (inputs(224));
    layer0_outputs(9897) <= not((inputs(112)) and (inputs(128)));
    layer0_outputs(9898) <= inputs(16);
    layer0_outputs(9899) <= inputs(8);
    layer0_outputs(9900) <= (inputs(136)) and not (inputs(96));
    layer0_outputs(9901) <= not((inputs(237)) or (inputs(23)));
    layer0_outputs(9902) <= inputs(124);
    layer0_outputs(9903) <= not((inputs(92)) xor (inputs(79)));
    layer0_outputs(9904) <= (inputs(122)) and not (inputs(35));
    layer0_outputs(9905) <= (inputs(130)) xor (inputs(103));
    layer0_outputs(9906) <= (inputs(63)) or (inputs(250));
    layer0_outputs(9907) <= inputs(177);
    layer0_outputs(9908) <= inputs(59);
    layer0_outputs(9909) <= (inputs(228)) or (inputs(51));
    layer0_outputs(9910) <= (inputs(27)) and not (inputs(181));
    layer0_outputs(9911) <= not(inputs(84));
    layer0_outputs(9912) <= (inputs(174)) xor (inputs(133));
    layer0_outputs(9913) <= inputs(14);
    layer0_outputs(9914) <= not(inputs(213));
    layer0_outputs(9915) <= inputs(211);
    layer0_outputs(9916) <= not((inputs(96)) xor (inputs(42)));
    layer0_outputs(9917) <= not((inputs(242)) or (inputs(248)));
    layer0_outputs(9918) <= inputs(162);
    layer0_outputs(9919) <= inputs(196);
    layer0_outputs(9920) <= not(inputs(238)) or (inputs(209));
    layer0_outputs(9921) <= inputs(248);
    layer0_outputs(9922) <= not((inputs(174)) or (inputs(61)));
    layer0_outputs(9923) <= (inputs(144)) xor (inputs(1));
    layer0_outputs(9924) <= not(inputs(152));
    layer0_outputs(9925) <= not(inputs(231));
    layer0_outputs(9926) <= not(inputs(246));
    layer0_outputs(9927) <= (inputs(230)) and not (inputs(146));
    layer0_outputs(9928) <= not(inputs(231));
    layer0_outputs(9929) <= (inputs(57)) or (inputs(193));
    layer0_outputs(9930) <= inputs(143);
    layer0_outputs(9931) <= (inputs(14)) xor (inputs(183));
    layer0_outputs(9932) <= (inputs(142)) and (inputs(82));
    layer0_outputs(9933) <= (inputs(89)) xor (inputs(209));
    layer0_outputs(9934) <= not(inputs(20));
    layer0_outputs(9935) <= not((inputs(25)) xor (inputs(80)));
    layer0_outputs(9936) <= (inputs(95)) and not (inputs(135));
    layer0_outputs(9937) <= not(inputs(179)) or (inputs(212));
    layer0_outputs(9938) <= '0';
    layer0_outputs(9939) <= not(inputs(230));
    layer0_outputs(9940) <= (inputs(99)) or (inputs(14));
    layer0_outputs(9941) <= (inputs(178)) xor (inputs(188));
    layer0_outputs(9942) <= (inputs(91)) and (inputs(30));
    layer0_outputs(9943) <= not((inputs(171)) and (inputs(228)));
    layer0_outputs(9944) <= (inputs(89)) and not (inputs(202));
    layer0_outputs(9945) <= inputs(174);
    layer0_outputs(9946) <= not(inputs(202));
    layer0_outputs(9947) <= not(inputs(153));
    layer0_outputs(9948) <= not(inputs(120)) or (inputs(32));
    layer0_outputs(9949) <= (inputs(158)) or (inputs(19));
    layer0_outputs(9950) <= (inputs(138)) or (inputs(15));
    layer0_outputs(9951) <= not(inputs(199)) or (inputs(76));
    layer0_outputs(9952) <= (inputs(63)) or (inputs(142));
    layer0_outputs(9953) <= (inputs(7)) or (inputs(60));
    layer0_outputs(9954) <= inputs(10);
    layer0_outputs(9955) <= inputs(122);
    layer0_outputs(9956) <= (inputs(196)) and not (inputs(61));
    layer0_outputs(9957) <= (inputs(46)) and not (inputs(188));
    layer0_outputs(9958) <= (inputs(239)) or (inputs(200));
    layer0_outputs(9959) <= not(inputs(43));
    layer0_outputs(9960) <= not(inputs(201)) or (inputs(27));
    layer0_outputs(9961) <= (inputs(232)) and not (inputs(255));
    layer0_outputs(9962) <= not(inputs(30)) or (inputs(254));
    layer0_outputs(9963) <= inputs(87);
    layer0_outputs(9964) <= not((inputs(93)) xor (inputs(2)));
    layer0_outputs(9965) <= inputs(23);
    layer0_outputs(9966) <= (inputs(34)) or (inputs(255));
    layer0_outputs(9967) <= (inputs(216)) xor (inputs(189));
    layer0_outputs(9968) <= (inputs(89)) and not (inputs(192));
    layer0_outputs(9969) <= not((inputs(160)) xor (inputs(131)));
    layer0_outputs(9970) <= not((inputs(102)) or (inputs(101)));
    layer0_outputs(9971) <= not(inputs(2));
    layer0_outputs(9972) <= (inputs(111)) xor (inputs(76));
    layer0_outputs(9973) <= not(inputs(150)) or (inputs(73));
    layer0_outputs(9974) <= not(inputs(33));
    layer0_outputs(9975) <= inputs(34);
    layer0_outputs(9976) <= (inputs(93)) xor (inputs(233));
    layer0_outputs(9977) <= (inputs(180)) xor (inputs(88));
    layer0_outputs(9978) <= inputs(243);
    layer0_outputs(9979) <= not(inputs(203));
    layer0_outputs(9980) <= not(inputs(232));
    layer0_outputs(9981) <= not(inputs(68));
    layer0_outputs(9982) <= not((inputs(16)) or (inputs(160)));
    layer0_outputs(9983) <= not(inputs(134)) or (inputs(14));
    layer0_outputs(9984) <= (inputs(90)) and not (inputs(118));
    layer0_outputs(9985) <= (inputs(32)) xor (inputs(60));
    layer0_outputs(9986) <= inputs(41);
    layer0_outputs(9987) <= not(inputs(50)) or (inputs(167));
    layer0_outputs(9988) <= not((inputs(184)) or (inputs(184)));
    layer0_outputs(9989) <= (inputs(218)) and not (inputs(63));
    layer0_outputs(9990) <= not((inputs(65)) or (inputs(29)));
    layer0_outputs(9991) <= not(inputs(179)) or (inputs(55));
    layer0_outputs(9992) <= not(inputs(104));
    layer0_outputs(9993) <= (inputs(147)) xor (inputs(153));
    layer0_outputs(9994) <= not(inputs(52)) or (inputs(72));
    layer0_outputs(9995) <= not(inputs(89));
    layer0_outputs(9996) <= not(inputs(26)) or (inputs(219));
    layer0_outputs(9997) <= not((inputs(113)) or (inputs(163)));
    layer0_outputs(9998) <= not(inputs(6));
    layer0_outputs(9999) <= (inputs(239)) and not (inputs(46));
    layer0_outputs(10000) <= not(inputs(139)) or (inputs(73));
    layer0_outputs(10001) <= not(inputs(71));
    layer0_outputs(10002) <= not(inputs(157)) or (inputs(182));
    layer0_outputs(10003) <= not(inputs(121)) or (inputs(156));
    layer0_outputs(10004) <= inputs(18);
    layer0_outputs(10005) <= not(inputs(212));
    layer0_outputs(10006) <= (inputs(177)) xor (inputs(92));
    layer0_outputs(10007) <= not(inputs(164));
    layer0_outputs(10008) <= (inputs(175)) and not (inputs(72));
    layer0_outputs(10009) <= not((inputs(21)) xor (inputs(204)));
    layer0_outputs(10010) <= not(inputs(183));
    layer0_outputs(10011) <= not(inputs(36));
    layer0_outputs(10012) <= (inputs(10)) or (inputs(1));
    layer0_outputs(10013) <= inputs(163);
    layer0_outputs(10014) <= inputs(44);
    layer0_outputs(10015) <= inputs(70);
    layer0_outputs(10016) <= not(inputs(175));
    layer0_outputs(10017) <= (inputs(155)) and not (inputs(26));
    layer0_outputs(10018) <= (inputs(162)) and (inputs(249));
    layer0_outputs(10019) <= inputs(100);
    layer0_outputs(10020) <= inputs(115);
    layer0_outputs(10021) <= (inputs(94)) and (inputs(92));
    layer0_outputs(10022) <= (inputs(150)) or (inputs(204));
    layer0_outputs(10023) <= not(inputs(142));
    layer0_outputs(10024) <= not((inputs(47)) or (inputs(46)));
    layer0_outputs(10025) <= (inputs(171)) or (inputs(208));
    layer0_outputs(10026) <= inputs(194);
    layer0_outputs(10027) <= not(inputs(154));
    layer0_outputs(10028) <= inputs(165);
    layer0_outputs(10029) <= inputs(122);
    layer0_outputs(10030) <= inputs(215);
    layer0_outputs(10031) <= not(inputs(114));
    layer0_outputs(10032) <= (inputs(187)) and not (inputs(143));
    layer0_outputs(10033) <= not((inputs(172)) or (inputs(79)));
    layer0_outputs(10034) <= not((inputs(109)) or (inputs(93)));
    layer0_outputs(10035) <= (inputs(116)) and not (inputs(4));
    layer0_outputs(10036) <= (inputs(172)) and not (inputs(54));
    layer0_outputs(10037) <= (inputs(236)) or (inputs(173));
    layer0_outputs(10038) <= not((inputs(22)) xor (inputs(50)));
    layer0_outputs(10039) <= (inputs(141)) and not (inputs(5));
    layer0_outputs(10040) <= (inputs(165)) xor (inputs(76));
    layer0_outputs(10041) <= (inputs(70)) xor (inputs(34));
    layer0_outputs(10042) <= (inputs(0)) and not (inputs(216));
    layer0_outputs(10043) <= not((inputs(56)) xor (inputs(30)));
    layer0_outputs(10044) <= (inputs(171)) xor (inputs(88));
    layer0_outputs(10045) <= not(inputs(114));
    layer0_outputs(10046) <= not(inputs(87));
    layer0_outputs(10047) <= not(inputs(99)) or (inputs(15));
    layer0_outputs(10048) <= inputs(191);
    layer0_outputs(10049) <= not((inputs(74)) xor (inputs(72)));
    layer0_outputs(10050) <= (inputs(42)) xor (inputs(118));
    layer0_outputs(10051) <= inputs(56);
    layer0_outputs(10052) <= (inputs(239)) and not (inputs(175));
    layer0_outputs(10053) <= inputs(99);
    layer0_outputs(10054) <= (inputs(142)) or (inputs(217));
    layer0_outputs(10055) <= inputs(232);
    layer0_outputs(10056) <= (inputs(108)) or (inputs(81));
    layer0_outputs(10057) <= inputs(5);
    layer0_outputs(10058) <= (inputs(252)) xor (inputs(127));
    layer0_outputs(10059) <= not((inputs(127)) or (inputs(201)));
    layer0_outputs(10060) <= inputs(133);
    layer0_outputs(10061) <= (inputs(236)) or (inputs(196));
    layer0_outputs(10062) <= not((inputs(4)) or (inputs(51)));
    layer0_outputs(10063) <= not(inputs(229));
    layer0_outputs(10064) <= (inputs(58)) or (inputs(97));
    layer0_outputs(10065) <= not(inputs(87)) or (inputs(19));
    layer0_outputs(10066) <= '1';
    layer0_outputs(10067) <= not((inputs(206)) xor (inputs(7)));
    layer0_outputs(10068) <= (inputs(210)) or (inputs(220));
    layer0_outputs(10069) <= '0';
    layer0_outputs(10070) <= inputs(216);
    layer0_outputs(10071) <= (inputs(66)) and not (inputs(107));
    layer0_outputs(10072) <= (inputs(195)) xor (inputs(189));
    layer0_outputs(10073) <= inputs(98);
    layer0_outputs(10074) <= not(inputs(88));
    layer0_outputs(10075) <= inputs(103);
    layer0_outputs(10076) <= inputs(151);
    layer0_outputs(10077) <= (inputs(88)) and (inputs(8));
    layer0_outputs(10078) <= inputs(52);
    layer0_outputs(10079) <= (inputs(66)) or (inputs(38));
    layer0_outputs(10080) <= not((inputs(64)) xor (inputs(112)));
    layer0_outputs(10081) <= not((inputs(192)) xor (inputs(90)));
    layer0_outputs(10082) <= inputs(66);
    layer0_outputs(10083) <= (inputs(234)) and (inputs(41));
    layer0_outputs(10084) <= (inputs(74)) xor (inputs(253));
    layer0_outputs(10085) <= (inputs(109)) or (inputs(78));
    layer0_outputs(10086) <= not((inputs(179)) xor (inputs(128)));
    layer0_outputs(10087) <= (inputs(176)) or (inputs(141));
    layer0_outputs(10088) <= (inputs(42)) and not (inputs(69));
    layer0_outputs(10089) <= not((inputs(35)) or (inputs(243)));
    layer0_outputs(10090) <= not(inputs(12)) or (inputs(154));
    layer0_outputs(10091) <= not((inputs(179)) or (inputs(188)));
    layer0_outputs(10092) <= (inputs(69)) xor (inputs(112));
    layer0_outputs(10093) <= not((inputs(118)) or (inputs(205)));
    layer0_outputs(10094) <= inputs(14);
    layer0_outputs(10095) <= not((inputs(86)) or (inputs(78)));
    layer0_outputs(10096) <= inputs(41);
    layer0_outputs(10097) <= (inputs(30)) or (inputs(182));
    layer0_outputs(10098) <= (inputs(72)) and (inputs(9));
    layer0_outputs(10099) <= inputs(102);
    layer0_outputs(10100) <= not(inputs(100));
    layer0_outputs(10101) <= (inputs(234)) or (inputs(217));
    layer0_outputs(10102) <= inputs(77);
    layer0_outputs(10103) <= not(inputs(120));
    layer0_outputs(10104) <= not(inputs(162));
    layer0_outputs(10105) <= not(inputs(54));
    layer0_outputs(10106) <= not((inputs(150)) and (inputs(181)));
    layer0_outputs(10107) <= not((inputs(173)) xor (inputs(194)));
    layer0_outputs(10108) <= not((inputs(43)) xor (inputs(11)));
    layer0_outputs(10109) <= not((inputs(187)) xor (inputs(116)));
    layer0_outputs(10110) <= not((inputs(197)) or (inputs(158)));
    layer0_outputs(10111) <= inputs(197);
    layer0_outputs(10112) <= not(inputs(235));
    layer0_outputs(10113) <= not(inputs(44));
    layer0_outputs(10114) <= not((inputs(145)) or (inputs(116)));
    layer0_outputs(10115) <= not((inputs(196)) xor (inputs(44)));
    layer0_outputs(10116) <= not((inputs(143)) xor (inputs(139)));
    layer0_outputs(10117) <= (inputs(204)) and (inputs(233));
    layer0_outputs(10118) <= inputs(5);
    layer0_outputs(10119) <= not((inputs(252)) xor (inputs(83)));
    layer0_outputs(10120) <= not((inputs(51)) or (inputs(52)));
    layer0_outputs(10121) <= not(inputs(131));
    layer0_outputs(10122) <= not((inputs(196)) or (inputs(220)));
    layer0_outputs(10123) <= inputs(125);
    layer0_outputs(10124) <= inputs(217);
    layer0_outputs(10125) <= not((inputs(81)) or (inputs(225)));
    layer0_outputs(10126) <= (inputs(72)) xor (inputs(67));
    layer0_outputs(10127) <= (inputs(35)) and (inputs(4));
    layer0_outputs(10128) <= not(inputs(227));
    layer0_outputs(10129) <= not(inputs(25));
    layer0_outputs(10130) <= inputs(104);
    layer0_outputs(10131) <= not(inputs(28)) or (inputs(193));
    layer0_outputs(10132) <= (inputs(57)) or (inputs(37));
    layer0_outputs(10133) <= inputs(23);
    layer0_outputs(10134) <= (inputs(202)) and not (inputs(37));
    layer0_outputs(10135) <= not((inputs(193)) xor (inputs(247)));
    layer0_outputs(10136) <= inputs(144);
    layer0_outputs(10137) <= (inputs(219)) and (inputs(131));
    layer0_outputs(10138) <= (inputs(95)) and not (inputs(241));
    layer0_outputs(10139) <= not(inputs(29)) or (inputs(144));
    layer0_outputs(10140) <= inputs(163);
    layer0_outputs(10141) <= '0';
    layer0_outputs(10142) <= not((inputs(131)) xor (inputs(161)));
    layer0_outputs(10143) <= not(inputs(36));
    layer0_outputs(10144) <= (inputs(212)) and (inputs(162));
    layer0_outputs(10145) <= not(inputs(153));
    layer0_outputs(10146) <= inputs(198);
    layer0_outputs(10147) <= inputs(193);
    layer0_outputs(10148) <= not((inputs(193)) xor (inputs(240)));
    layer0_outputs(10149) <= not(inputs(147)) or (inputs(208));
    layer0_outputs(10150) <= (inputs(204)) and not (inputs(254));
    layer0_outputs(10151) <= (inputs(180)) and not (inputs(1));
    layer0_outputs(10152) <= (inputs(5)) or (inputs(28));
    layer0_outputs(10153) <= (inputs(137)) and not (inputs(18));
    layer0_outputs(10154) <= (inputs(132)) xor (inputs(51));
    layer0_outputs(10155) <= inputs(120);
    layer0_outputs(10156) <= not((inputs(194)) xor (inputs(65)));
    layer0_outputs(10157) <= not(inputs(26));
    layer0_outputs(10158) <= (inputs(131)) or (inputs(78));
    layer0_outputs(10159) <= (inputs(171)) xor (inputs(19));
    layer0_outputs(10160) <= not((inputs(207)) xor (inputs(23)));
    layer0_outputs(10161) <= not((inputs(187)) and (inputs(202)));
    layer0_outputs(10162) <= inputs(54);
    layer0_outputs(10163) <= inputs(247);
    layer0_outputs(10164) <= not(inputs(7)) or (inputs(86));
    layer0_outputs(10165) <= not((inputs(206)) or (inputs(190)));
    layer0_outputs(10166) <= inputs(74);
    layer0_outputs(10167) <= (inputs(248)) and not (inputs(63));
    layer0_outputs(10168) <= (inputs(120)) and not (inputs(165));
    layer0_outputs(10169) <= '1';
    layer0_outputs(10170) <= inputs(167);
    layer0_outputs(10171) <= (inputs(46)) xor (inputs(5));
    layer0_outputs(10172) <= not(inputs(114)) or (inputs(191));
    layer0_outputs(10173) <= not((inputs(38)) or (inputs(239)));
    layer0_outputs(10174) <= inputs(13);
    layer0_outputs(10175) <= not((inputs(29)) or (inputs(225)));
    layer0_outputs(10176) <= (inputs(42)) and (inputs(133));
    layer0_outputs(10177) <= (inputs(152)) or (inputs(124));
    layer0_outputs(10178) <= not(inputs(115));
    layer0_outputs(10179) <= inputs(37);
    layer0_outputs(10180) <= not(inputs(22));
    layer0_outputs(10181) <= not((inputs(248)) or (inputs(163)));
    layer0_outputs(10182) <= not(inputs(240)) or (inputs(78));
    layer0_outputs(10183) <= not(inputs(1));
    layer0_outputs(10184) <= not((inputs(126)) or (inputs(48)));
    layer0_outputs(10185) <= inputs(25);
    layer0_outputs(10186) <= inputs(54);
    layer0_outputs(10187) <= inputs(249);
    layer0_outputs(10188) <= (inputs(183)) or (inputs(237));
    layer0_outputs(10189) <= not((inputs(140)) xor (inputs(196)));
    layer0_outputs(10190) <= (inputs(53)) xor (inputs(34));
    layer0_outputs(10191) <= (inputs(243)) or (inputs(204));
    layer0_outputs(10192) <= not((inputs(169)) xor (inputs(129)));
    layer0_outputs(10193) <= inputs(89);
    layer0_outputs(10194) <= (inputs(172)) and not (inputs(17));
    layer0_outputs(10195) <= inputs(8);
    layer0_outputs(10196) <= not((inputs(72)) or (inputs(64)));
    layer0_outputs(10197) <= (inputs(128)) or (inputs(66));
    layer0_outputs(10198) <= not((inputs(80)) or (inputs(118)));
    layer0_outputs(10199) <= not((inputs(236)) and (inputs(35)));
    layer0_outputs(10200) <= inputs(87);
    layer0_outputs(10201) <= (inputs(29)) and not (inputs(226));
    layer0_outputs(10202) <= (inputs(186)) or (inputs(17));
    layer0_outputs(10203) <= inputs(69);
    layer0_outputs(10204) <= not(inputs(9)) or (inputs(143));
    layer0_outputs(10205) <= not(inputs(254));
    layer0_outputs(10206) <= '0';
    layer0_outputs(10207) <= not((inputs(67)) xor (inputs(82)));
    layer0_outputs(10208) <= not(inputs(67));
    layer0_outputs(10209) <= (inputs(184)) or (inputs(165));
    layer0_outputs(10210) <= not((inputs(206)) or (inputs(205)));
    layer0_outputs(10211) <= (inputs(89)) and not (inputs(250));
    layer0_outputs(10212) <= (inputs(222)) xor (inputs(78));
    layer0_outputs(10213) <= not(inputs(231)) or (inputs(30));
    layer0_outputs(10214) <= not((inputs(28)) or (inputs(100)));
    layer0_outputs(10215) <= not(inputs(131));
    layer0_outputs(10216) <= not(inputs(50));
    layer0_outputs(10217) <= inputs(104);
    layer0_outputs(10218) <= not((inputs(55)) xor (inputs(114)));
    layer0_outputs(10219) <= not((inputs(4)) or (inputs(34)));
    layer0_outputs(10220) <= not(inputs(172));
    layer0_outputs(10221) <= not((inputs(0)) xor (inputs(50)));
    layer0_outputs(10222) <= not((inputs(158)) xor (inputs(106)));
    layer0_outputs(10223) <= (inputs(120)) and not (inputs(9));
    layer0_outputs(10224) <= (inputs(105)) and not (inputs(236));
    layer0_outputs(10225) <= (inputs(28)) and not (inputs(254));
    layer0_outputs(10226) <= (inputs(191)) and not (inputs(166));
    layer0_outputs(10227) <= not(inputs(54));
    layer0_outputs(10228) <= not(inputs(141));
    layer0_outputs(10229) <= (inputs(76)) or (inputs(135));
    layer0_outputs(10230) <= (inputs(127)) and not (inputs(252));
    layer0_outputs(10231) <= not((inputs(91)) or (inputs(108)));
    layer0_outputs(10232) <= (inputs(103)) or (inputs(226));
    layer0_outputs(10233) <= not((inputs(181)) or (inputs(1)));
    layer0_outputs(10234) <= inputs(30);
    layer0_outputs(10235) <= inputs(33);
    layer0_outputs(10236) <= not(inputs(216));
    layer0_outputs(10237) <= not(inputs(100));
    layer0_outputs(10238) <= not(inputs(79)) or (inputs(190));
    layer0_outputs(10239) <= (inputs(113)) and not (inputs(111));
    outputs(0) <= (layer0_outputs(333)) or (layer0_outputs(2974));
    outputs(1) <= not((layer0_outputs(2196)) xor (layer0_outputs(3350)));
    outputs(2) <= (layer0_outputs(7747)) and not (layer0_outputs(509));
    outputs(3) <= (layer0_outputs(8588)) xor (layer0_outputs(7564));
    outputs(4) <= (layer0_outputs(3872)) or (layer0_outputs(4473));
    outputs(5) <= not(layer0_outputs(9435));
    outputs(6) <= not(layer0_outputs(9013));
    outputs(7) <= not((layer0_outputs(3640)) xor (layer0_outputs(2189)));
    outputs(8) <= not(layer0_outputs(6306));
    outputs(9) <= (layer0_outputs(1357)) and not (layer0_outputs(4129));
    outputs(10) <= not(layer0_outputs(8901));
    outputs(11) <= not((layer0_outputs(8460)) xor (layer0_outputs(4558)));
    outputs(12) <= not(layer0_outputs(8481));
    outputs(13) <= not((layer0_outputs(7550)) and (layer0_outputs(6540)));
    outputs(14) <= not((layer0_outputs(9425)) or (layer0_outputs(3900)));
    outputs(15) <= layer0_outputs(782);
    outputs(16) <= (layer0_outputs(7857)) and (layer0_outputs(295));
    outputs(17) <= not(layer0_outputs(4773));
    outputs(18) <= layer0_outputs(1423);
    outputs(19) <= '0';
    outputs(20) <= layer0_outputs(8422);
    outputs(21) <= not((layer0_outputs(2786)) or (layer0_outputs(2517)));
    outputs(22) <= not(layer0_outputs(2001)) or (layer0_outputs(8036));
    outputs(23) <= (layer0_outputs(231)) xor (layer0_outputs(7443));
    outputs(24) <= not(layer0_outputs(2970)) or (layer0_outputs(1334));
    outputs(25) <= not(layer0_outputs(2939));
    outputs(26) <= (layer0_outputs(2005)) xor (layer0_outputs(522));
    outputs(27) <= layer0_outputs(94);
    outputs(28) <= not(layer0_outputs(3334));
    outputs(29) <= not((layer0_outputs(3425)) and (layer0_outputs(9840)));
    outputs(30) <= layer0_outputs(7195);
    outputs(31) <= not(layer0_outputs(1665)) or (layer0_outputs(8291));
    outputs(32) <= not((layer0_outputs(8754)) xor (layer0_outputs(8451)));
    outputs(33) <= not(layer0_outputs(4773));
    outputs(34) <= layer0_outputs(4903);
    outputs(35) <= layer0_outputs(4516);
    outputs(36) <= not(layer0_outputs(3773));
    outputs(37) <= not(layer0_outputs(509));
    outputs(38) <= (layer0_outputs(4053)) xor (layer0_outputs(1413));
    outputs(39) <= not(layer0_outputs(9208));
    outputs(40) <= (layer0_outputs(9364)) and not (layer0_outputs(4620));
    outputs(41) <= not((layer0_outputs(1707)) xor (layer0_outputs(6345)));
    outputs(42) <= not((layer0_outputs(3209)) xor (layer0_outputs(1279)));
    outputs(43) <= layer0_outputs(4505);
    outputs(44) <= not(layer0_outputs(6587));
    outputs(45) <= layer0_outputs(2515);
    outputs(46) <= not(layer0_outputs(5944));
    outputs(47) <= not(layer0_outputs(1537));
    outputs(48) <= not(layer0_outputs(9371)) or (layer0_outputs(9227));
    outputs(49) <= layer0_outputs(2131);
    outputs(50) <= not((layer0_outputs(1445)) xor (layer0_outputs(4328)));
    outputs(51) <= (layer0_outputs(8993)) and not (layer0_outputs(4272));
    outputs(52) <= (layer0_outputs(9971)) xor (layer0_outputs(1956));
    outputs(53) <= not(layer0_outputs(9032));
    outputs(54) <= (layer0_outputs(1198)) or (layer0_outputs(7892));
    outputs(55) <= not(layer0_outputs(6150));
    outputs(56) <= layer0_outputs(3528);
    outputs(57) <= layer0_outputs(426);
    outputs(58) <= not((layer0_outputs(1425)) or (layer0_outputs(3626)));
    outputs(59) <= not((layer0_outputs(5377)) xor (layer0_outputs(837)));
    outputs(60) <= (layer0_outputs(3616)) or (layer0_outputs(9559));
    outputs(61) <= not(layer0_outputs(6219));
    outputs(62) <= not(layer0_outputs(7298)) or (layer0_outputs(9331));
    outputs(63) <= (layer0_outputs(7768)) or (layer0_outputs(3435));
    outputs(64) <= not(layer0_outputs(8659));
    outputs(65) <= layer0_outputs(1988);
    outputs(66) <= (layer0_outputs(7912)) xor (layer0_outputs(1022));
    outputs(67) <= (layer0_outputs(9408)) or (layer0_outputs(7864));
    outputs(68) <= (layer0_outputs(6324)) xor (layer0_outputs(4377));
    outputs(69) <= (layer0_outputs(3335)) and not (layer0_outputs(6783));
    outputs(70) <= layer0_outputs(1768);
    outputs(71) <= not((layer0_outputs(6070)) and (layer0_outputs(7861)));
    outputs(72) <= layer0_outputs(6214);
    outputs(73) <= layer0_outputs(10159);
    outputs(74) <= (layer0_outputs(5520)) or (layer0_outputs(1967));
    outputs(75) <= (layer0_outputs(5067)) or (layer0_outputs(2147));
    outputs(76) <= layer0_outputs(7441);
    outputs(77) <= not(layer0_outputs(2347));
    outputs(78) <= not(layer0_outputs(6868));
    outputs(79) <= (layer0_outputs(8328)) xor (layer0_outputs(1933));
    outputs(80) <= not(layer0_outputs(4373));
    outputs(81) <= not(layer0_outputs(6199));
    outputs(82) <= '1';
    outputs(83) <= not(layer0_outputs(7540));
    outputs(84) <= (layer0_outputs(969)) and not (layer0_outputs(368));
    outputs(85) <= (layer0_outputs(8749)) xor (layer0_outputs(672));
    outputs(86) <= layer0_outputs(3174);
    outputs(87) <= not((layer0_outputs(3744)) xor (layer0_outputs(8174)));
    outputs(88) <= layer0_outputs(9443);
    outputs(89) <= not(layer0_outputs(3378));
    outputs(90) <= layer0_outputs(7644);
    outputs(91) <= not(layer0_outputs(9323)) or (layer0_outputs(4880));
    outputs(92) <= (layer0_outputs(553)) or (layer0_outputs(7642));
    outputs(93) <= layer0_outputs(8070);
    outputs(94) <= not(layer0_outputs(2247));
    outputs(95) <= layer0_outputs(6178);
    outputs(96) <= not((layer0_outputs(3941)) xor (layer0_outputs(6161)));
    outputs(97) <= not(layer0_outputs(7121)) or (layer0_outputs(3926));
    outputs(98) <= layer0_outputs(6850);
    outputs(99) <= (layer0_outputs(3299)) xor (layer0_outputs(7886));
    outputs(100) <= layer0_outputs(10096);
    outputs(101) <= not(layer0_outputs(7444));
    outputs(102) <= not((layer0_outputs(2991)) xor (layer0_outputs(7837)));
    outputs(103) <= layer0_outputs(1241);
    outputs(104) <= layer0_outputs(7261);
    outputs(105) <= not(layer0_outputs(396));
    outputs(106) <= not(layer0_outputs(5837));
    outputs(107) <= layer0_outputs(6110);
    outputs(108) <= not((layer0_outputs(2948)) xor (layer0_outputs(8532)));
    outputs(109) <= layer0_outputs(4975);
    outputs(110) <= not(layer0_outputs(6395));
    outputs(111) <= layer0_outputs(542);
    outputs(112) <= (layer0_outputs(6720)) and (layer0_outputs(4718));
    outputs(113) <= layer0_outputs(8761);
    outputs(114) <= (layer0_outputs(10165)) and not (layer0_outputs(5990));
    outputs(115) <= not(layer0_outputs(8164));
    outputs(116) <= not(layer0_outputs(2671));
    outputs(117) <= not(layer0_outputs(2165));
    outputs(118) <= not(layer0_outputs(3978));
    outputs(119) <= layer0_outputs(6508);
    outputs(120) <= not(layer0_outputs(4030));
    outputs(121) <= not((layer0_outputs(9682)) xor (layer0_outputs(4113)));
    outputs(122) <= layer0_outputs(9770);
    outputs(123) <= not(layer0_outputs(3615));
    outputs(124) <= not(layer0_outputs(9997));
    outputs(125) <= layer0_outputs(1686);
    outputs(126) <= not(layer0_outputs(5947));
    outputs(127) <= not((layer0_outputs(4754)) and (layer0_outputs(4318)));
    outputs(128) <= layer0_outputs(9688);
    outputs(129) <= not(layer0_outputs(9548));
    outputs(130) <= layer0_outputs(6673);
    outputs(131) <= not(layer0_outputs(1874));
    outputs(132) <= (layer0_outputs(916)) and (layer0_outputs(7753));
    outputs(133) <= (layer0_outputs(9505)) and not (layer0_outputs(8018));
    outputs(134) <= (layer0_outputs(9723)) and not (layer0_outputs(9702));
    outputs(135) <= not((layer0_outputs(4501)) and (layer0_outputs(5565)));
    outputs(136) <= layer0_outputs(4092);
    outputs(137) <= not(layer0_outputs(4817));
    outputs(138) <= layer0_outputs(5938);
    outputs(139) <= not((layer0_outputs(9129)) and (layer0_outputs(6509)));
    outputs(140) <= layer0_outputs(3999);
    outputs(141) <= (layer0_outputs(7406)) xor (layer0_outputs(2104));
    outputs(142) <= (layer0_outputs(9611)) xor (layer0_outputs(8909));
    outputs(143) <= (layer0_outputs(9849)) or (layer0_outputs(7046));
    outputs(144) <= not((layer0_outputs(880)) and (layer0_outputs(8685)));
    outputs(145) <= (layer0_outputs(7504)) or (layer0_outputs(7315));
    outputs(146) <= (layer0_outputs(2841)) and (layer0_outputs(2581));
    outputs(147) <= layer0_outputs(690);
    outputs(148) <= (layer0_outputs(3991)) xor (layer0_outputs(8479));
    outputs(149) <= not(layer0_outputs(5516));
    outputs(150) <= (layer0_outputs(7778)) or (layer0_outputs(9485));
    outputs(151) <= (layer0_outputs(1368)) and not (layer0_outputs(10097));
    outputs(152) <= (layer0_outputs(8508)) xor (layer0_outputs(79));
    outputs(153) <= (layer0_outputs(5707)) or (layer0_outputs(4887));
    outputs(154) <= (layer0_outputs(2653)) and (layer0_outputs(431));
    outputs(155) <= layer0_outputs(7083);
    outputs(156) <= (layer0_outputs(9804)) xor (layer0_outputs(157));
    outputs(157) <= not(layer0_outputs(1020)) or (layer0_outputs(7294));
    outputs(158) <= not((layer0_outputs(641)) or (layer0_outputs(3743)));
    outputs(159) <= not(layer0_outputs(4507));
    outputs(160) <= not((layer0_outputs(9656)) or (layer0_outputs(6267)));
    outputs(161) <= not((layer0_outputs(3978)) or (layer0_outputs(10005)));
    outputs(162) <= not(layer0_outputs(5912));
    outputs(163) <= (layer0_outputs(9851)) or (layer0_outputs(1593));
    outputs(164) <= (layer0_outputs(410)) and not (layer0_outputs(1853));
    outputs(165) <= not(layer0_outputs(3690));
    outputs(166) <= not((layer0_outputs(3642)) xor (layer0_outputs(334)));
    outputs(167) <= layer0_outputs(9341);
    outputs(168) <= not(layer0_outputs(9223));
    outputs(169) <= (layer0_outputs(1640)) xor (layer0_outputs(1625));
    outputs(170) <= (layer0_outputs(8525)) and not (layer0_outputs(2851));
    outputs(171) <= not((layer0_outputs(596)) or (layer0_outputs(5130)));
    outputs(172) <= layer0_outputs(8931);
    outputs(173) <= not(layer0_outputs(10121));
    outputs(174) <= not(layer0_outputs(1134));
    outputs(175) <= layer0_outputs(358);
    outputs(176) <= not(layer0_outputs(8258));
    outputs(177) <= not(layer0_outputs(29));
    outputs(178) <= layer0_outputs(4276);
    outputs(179) <= layer0_outputs(5395);
    outputs(180) <= not((layer0_outputs(5616)) and (layer0_outputs(5636)));
    outputs(181) <= layer0_outputs(6849);
    outputs(182) <= not(layer0_outputs(2063));
    outputs(183) <= not(layer0_outputs(8147));
    outputs(184) <= not(layer0_outputs(7590));
    outputs(185) <= layer0_outputs(2950);
    outputs(186) <= (layer0_outputs(6179)) or (layer0_outputs(7703));
    outputs(187) <= layer0_outputs(624);
    outputs(188) <= layer0_outputs(3546);
    outputs(189) <= (layer0_outputs(3293)) and not (layer0_outputs(8541));
    outputs(190) <= (layer0_outputs(2965)) and not (layer0_outputs(7568));
    outputs(191) <= not(layer0_outputs(3814));
    outputs(192) <= layer0_outputs(6820);
    outputs(193) <= not(layer0_outputs(8162));
    outputs(194) <= not(layer0_outputs(8329));
    outputs(195) <= (layer0_outputs(8448)) and (layer0_outputs(1594));
    outputs(196) <= (layer0_outputs(5884)) xor (layer0_outputs(1384));
    outputs(197) <= not((layer0_outputs(4443)) xor (layer0_outputs(5102)));
    outputs(198) <= not(layer0_outputs(3044));
    outputs(199) <= not(layer0_outputs(2898));
    outputs(200) <= not(layer0_outputs(4147));
    outputs(201) <= not(layer0_outputs(3122));
    outputs(202) <= not((layer0_outputs(336)) xor (layer0_outputs(6472)));
    outputs(203) <= layer0_outputs(8833);
    outputs(204) <= not(layer0_outputs(3791));
    outputs(205) <= not((layer0_outputs(7163)) and (layer0_outputs(6768)));
    outputs(206) <= (layer0_outputs(1464)) xor (layer0_outputs(2378));
    outputs(207) <= layer0_outputs(6290);
    outputs(208) <= layer0_outputs(4568);
    outputs(209) <= not(layer0_outputs(9328));
    outputs(210) <= (layer0_outputs(3440)) and (layer0_outputs(47));
    outputs(211) <= layer0_outputs(3453);
    outputs(212) <= layer0_outputs(9638);
    outputs(213) <= layer0_outputs(2121);
    outputs(214) <= not(layer0_outputs(2978));
    outputs(215) <= not((layer0_outputs(1045)) and (layer0_outputs(5743)));
    outputs(216) <= not((layer0_outputs(3284)) xor (layer0_outputs(134)));
    outputs(217) <= not(layer0_outputs(6217));
    outputs(218) <= not(layer0_outputs(8060)) or (layer0_outputs(6522));
    outputs(219) <= (layer0_outputs(5878)) and not (layer0_outputs(4963));
    outputs(220) <= layer0_outputs(9589);
    outputs(221) <= (layer0_outputs(3739)) xor (layer0_outputs(2590));
    outputs(222) <= layer0_outputs(6706);
    outputs(223) <= (layer0_outputs(3761)) xor (layer0_outputs(9110));
    outputs(224) <= not((layer0_outputs(4659)) xor (layer0_outputs(6536)));
    outputs(225) <= not((layer0_outputs(2694)) or (layer0_outputs(6409)));
    outputs(226) <= not(layer0_outputs(6834));
    outputs(227) <= layer0_outputs(2267);
    outputs(228) <= not(layer0_outputs(3805));
    outputs(229) <= not(layer0_outputs(4885)) or (layer0_outputs(2613));
    outputs(230) <= layer0_outputs(4764);
    outputs(231) <= (layer0_outputs(5621)) and not (layer0_outputs(791));
    outputs(232) <= (layer0_outputs(7828)) xor (layer0_outputs(9217));
    outputs(233) <= not((layer0_outputs(6237)) xor (layer0_outputs(5876)));
    outputs(234) <= (layer0_outputs(4480)) and not (layer0_outputs(1613));
    outputs(235) <= not((layer0_outputs(5653)) and (layer0_outputs(2709)));
    outputs(236) <= not(layer0_outputs(2155));
    outputs(237) <= not((layer0_outputs(4738)) xor (layer0_outputs(1670)));
    outputs(238) <= layer0_outputs(4799);
    outputs(239) <= (layer0_outputs(5254)) and not (layer0_outputs(6443));
    outputs(240) <= not((layer0_outputs(9172)) xor (layer0_outputs(5151)));
    outputs(241) <= not(layer0_outputs(5932));
    outputs(242) <= (layer0_outputs(7514)) and (layer0_outputs(3998));
    outputs(243) <= not(layer0_outputs(7739));
    outputs(244) <= (layer0_outputs(3684)) xor (layer0_outputs(6117));
    outputs(245) <= layer0_outputs(1363);
    outputs(246) <= not(layer0_outputs(10168));
    outputs(247) <= not(layer0_outputs(2258));
    outputs(248) <= (layer0_outputs(7844)) and not (layer0_outputs(4709));
    outputs(249) <= layer0_outputs(3028);
    outputs(250) <= (layer0_outputs(10146)) xor (layer0_outputs(6614));
    outputs(251) <= layer0_outputs(6261);
    outputs(252) <= not((layer0_outputs(10094)) xor (layer0_outputs(2563)));
    outputs(253) <= (layer0_outputs(392)) and not (layer0_outputs(2382));
    outputs(254) <= (layer0_outputs(7223)) and not (layer0_outputs(8628));
    outputs(255) <= (layer0_outputs(9246)) and (layer0_outputs(6086));
    outputs(256) <= layer0_outputs(5336);
    outputs(257) <= not(layer0_outputs(9325)) or (layer0_outputs(5410));
    outputs(258) <= layer0_outputs(3806);
    outputs(259) <= (layer0_outputs(3955)) or (layer0_outputs(1683));
    outputs(260) <= not(layer0_outputs(9244)) or (layer0_outputs(665));
    outputs(261) <= not(layer0_outputs(3550));
    outputs(262) <= layer0_outputs(804);
    outputs(263) <= not(layer0_outputs(8061));
    outputs(264) <= not(layer0_outputs(694));
    outputs(265) <= not((layer0_outputs(6021)) and (layer0_outputs(9270)));
    outputs(266) <= not(layer0_outputs(5199)) or (layer0_outputs(2761));
    outputs(267) <= (layer0_outputs(7758)) and not (layer0_outputs(3319));
    outputs(268) <= not(layer0_outputs(8468));
    outputs(269) <= not((layer0_outputs(9174)) or (layer0_outputs(1895)));
    outputs(270) <= not(layer0_outputs(5182));
    outputs(271) <= layer0_outputs(2459);
    outputs(272) <= (layer0_outputs(8799)) xor (layer0_outputs(3751));
    outputs(273) <= not(layer0_outputs(10124)) or (layer0_outputs(7269));
    outputs(274) <= not(layer0_outputs(519));
    outputs(275) <= (layer0_outputs(6464)) xor (layer0_outputs(5209));
    outputs(276) <= layer0_outputs(6047);
    outputs(277) <= not((layer0_outputs(9410)) or (layer0_outputs(4427)));
    outputs(278) <= not(layer0_outputs(9428));
    outputs(279) <= not((layer0_outputs(7225)) and (layer0_outputs(7423)));
    outputs(280) <= not(layer0_outputs(5199));
    outputs(281) <= not(layer0_outputs(6602));
    outputs(282) <= layer0_outputs(10167);
    outputs(283) <= not((layer0_outputs(770)) or (layer0_outputs(4414)));
    outputs(284) <= not(layer0_outputs(5605));
    outputs(285) <= (layer0_outputs(3542)) and not (layer0_outputs(113));
    outputs(286) <= (layer0_outputs(7364)) xor (layer0_outputs(4438));
    outputs(287) <= (layer0_outputs(77)) or (layer0_outputs(3685));
    outputs(288) <= not(layer0_outputs(6687));
    outputs(289) <= (layer0_outputs(7350)) and not (layer0_outputs(4164));
    outputs(290) <= not(layer0_outputs(8801));
    outputs(291) <= layer0_outputs(4608);
    outputs(292) <= not(layer0_outputs(9523)) or (layer0_outputs(3806));
    outputs(293) <= (layer0_outputs(3798)) and not (layer0_outputs(3970));
    outputs(294) <= layer0_outputs(624);
    outputs(295) <= layer0_outputs(7291);
    outputs(296) <= layer0_outputs(5389);
    outputs(297) <= not(layer0_outputs(8876));
    outputs(298) <= not(layer0_outputs(4711));
    outputs(299) <= layer0_outputs(517);
    outputs(300) <= not(layer0_outputs(8430));
    outputs(301) <= not(layer0_outputs(6503));
    outputs(302) <= not(layer0_outputs(9363));
    outputs(303) <= not(layer0_outputs(2524));
    outputs(304) <= not(layer0_outputs(3456));
    outputs(305) <= layer0_outputs(8355);
    outputs(306) <= (layer0_outputs(370)) xor (layer0_outputs(7302));
    outputs(307) <= not((layer0_outputs(9468)) and (layer0_outputs(2953)));
    outputs(308) <= not(layer0_outputs(8132));
    outputs(309) <= layer0_outputs(9907);
    outputs(310) <= layer0_outputs(438);
    outputs(311) <= layer0_outputs(5728);
    outputs(312) <= not(layer0_outputs(8900));
    outputs(313) <= not((layer0_outputs(3862)) xor (layer0_outputs(10236)));
    outputs(314) <= (layer0_outputs(3338)) and (layer0_outputs(6860));
    outputs(315) <= not(layer0_outputs(3506));
    outputs(316) <= layer0_outputs(5433);
    outputs(317) <= not(layer0_outputs(531)) or (layer0_outputs(8154));
    outputs(318) <= layer0_outputs(9619);
    outputs(319) <= not(layer0_outputs(337)) or (layer0_outputs(2686));
    outputs(320) <= (layer0_outputs(6296)) xor (layer0_outputs(4921));
    outputs(321) <= (layer0_outputs(3085)) or (layer0_outputs(7166));
    outputs(322) <= not(layer0_outputs(4678));
    outputs(323) <= (layer0_outputs(2680)) and (layer0_outputs(3345));
    outputs(324) <= layer0_outputs(8308);
    outputs(325) <= not((layer0_outputs(1732)) and (layer0_outputs(9208)));
    outputs(326) <= not(layer0_outputs(9401));
    outputs(327) <= (layer0_outputs(3435)) and not (layer0_outputs(4945));
    outputs(328) <= not((layer0_outputs(8436)) xor (layer0_outputs(6627)));
    outputs(329) <= not((layer0_outputs(498)) or (layer0_outputs(4892)));
    outputs(330) <= layer0_outputs(1366);
    outputs(331) <= not((layer0_outputs(4914)) and (layer0_outputs(3374)));
    outputs(332) <= (layer0_outputs(2084)) and not (layer0_outputs(9839));
    outputs(333) <= (layer0_outputs(837)) or (layer0_outputs(8511));
    outputs(334) <= not(layer0_outputs(5664)) or (layer0_outputs(9795));
    outputs(335) <= not((layer0_outputs(4652)) and (layer0_outputs(3123)));
    outputs(336) <= (layer0_outputs(7302)) or (layer0_outputs(467));
    outputs(337) <= not(layer0_outputs(2620));
    outputs(338) <= not(layer0_outputs(4631)) or (layer0_outputs(6494));
    outputs(339) <= not(layer0_outputs(5196));
    outputs(340) <= not((layer0_outputs(1895)) and (layer0_outputs(4382)));
    outputs(341) <= not(layer0_outputs(1502)) or (layer0_outputs(2847));
    outputs(342) <= not(layer0_outputs(6883));
    outputs(343) <= not((layer0_outputs(9187)) and (layer0_outputs(9438)));
    outputs(344) <= not(layer0_outputs(58));
    outputs(345) <= layer0_outputs(7588);
    outputs(346) <= layer0_outputs(639);
    outputs(347) <= layer0_outputs(7441);
    outputs(348) <= not((layer0_outputs(3414)) and (layer0_outputs(4970)));
    outputs(349) <= not((layer0_outputs(2783)) and (layer0_outputs(8885)));
    outputs(350) <= (layer0_outputs(8940)) and not (layer0_outputs(2058));
    outputs(351) <= not((layer0_outputs(1641)) xor (layer0_outputs(7114)));
    outputs(352) <= not(layer0_outputs(177));
    outputs(353) <= (layer0_outputs(3459)) and not (layer0_outputs(7767));
    outputs(354) <= not(layer0_outputs(2100));
    outputs(355) <= not((layer0_outputs(2451)) xor (layer0_outputs(1351)));
    outputs(356) <= not(layer0_outputs(3473));
    outputs(357) <= (layer0_outputs(8443)) and not (layer0_outputs(6821));
    outputs(358) <= layer0_outputs(3904);
    outputs(359) <= not(layer0_outputs(4972));
    outputs(360) <= not(layer0_outputs(6032));
    outputs(361) <= (layer0_outputs(409)) xor (layer0_outputs(1151));
    outputs(362) <= layer0_outputs(8626);
    outputs(363) <= (layer0_outputs(3357)) xor (layer0_outputs(9311));
    outputs(364) <= layer0_outputs(8907);
    outputs(365) <= not((layer0_outputs(2495)) xor (layer0_outputs(8688)));
    outputs(366) <= layer0_outputs(9248);
    outputs(367) <= layer0_outputs(606);
    outputs(368) <= not(layer0_outputs(8326));
    outputs(369) <= layer0_outputs(5942);
    outputs(370) <= layer0_outputs(7857);
    outputs(371) <= not((layer0_outputs(10170)) or (layer0_outputs(3789)));
    outputs(372) <= not((layer0_outputs(7397)) or (layer0_outputs(1696)));
    outputs(373) <= layer0_outputs(3094);
    outputs(374) <= not(layer0_outputs(8086));
    outputs(375) <= (layer0_outputs(6215)) and (layer0_outputs(1466));
    outputs(376) <= (layer0_outputs(1312)) and (layer0_outputs(627));
    outputs(377) <= not((layer0_outputs(6206)) or (layer0_outputs(4972)));
    outputs(378) <= not(layer0_outputs(4949));
    outputs(379) <= not(layer0_outputs(5530)) or (layer0_outputs(1876));
    outputs(380) <= layer0_outputs(2567);
    outputs(381) <= not((layer0_outputs(3991)) xor (layer0_outputs(7012)));
    outputs(382) <= not((layer0_outputs(1476)) and (layer0_outputs(9307)));
    outputs(383) <= not((layer0_outputs(5671)) and (layer0_outputs(3019)));
    outputs(384) <= layer0_outputs(7918);
    outputs(385) <= layer0_outputs(4955);
    outputs(386) <= (layer0_outputs(8671)) and not (layer0_outputs(3570));
    outputs(387) <= layer0_outputs(6955);
    outputs(388) <= layer0_outputs(3904);
    outputs(389) <= not(layer0_outputs(9309)) or (layer0_outputs(7736));
    outputs(390) <= not(layer0_outputs(5790));
    outputs(391) <= not((layer0_outputs(169)) xor (layer0_outputs(3546)));
    outputs(392) <= (layer0_outputs(385)) xor (layer0_outputs(8878));
    outputs(393) <= (layer0_outputs(8786)) xor (layer0_outputs(8821));
    outputs(394) <= not(layer0_outputs(6838));
    outputs(395) <= (layer0_outputs(8851)) xor (layer0_outputs(8197));
    outputs(396) <= layer0_outputs(6702);
    outputs(397) <= layer0_outputs(296);
    outputs(398) <= layer0_outputs(9603);
    outputs(399) <= not(layer0_outputs(6620)) or (layer0_outputs(3698));
    outputs(400) <= (layer0_outputs(7696)) or (layer0_outputs(2460));
    outputs(401) <= not(layer0_outputs(580));
    outputs(402) <= not(layer0_outputs(9808)) or (layer0_outputs(643));
    outputs(403) <= not((layer0_outputs(6079)) or (layer0_outputs(7249)));
    outputs(404) <= not((layer0_outputs(3513)) or (layer0_outputs(999)));
    outputs(405) <= (layer0_outputs(6655)) xor (layer0_outputs(1175));
    outputs(406) <= layer0_outputs(10000);
    outputs(407) <= layer0_outputs(3496);
    outputs(408) <= layer0_outputs(8947);
    outputs(409) <= not(layer0_outputs(1143));
    outputs(410) <= (layer0_outputs(3850)) xor (layer0_outputs(2560));
    outputs(411) <= not(layer0_outputs(5550));
    outputs(412) <= (layer0_outputs(6836)) xor (layer0_outputs(4229));
    outputs(413) <= not(layer0_outputs(7029));
    outputs(414) <= not(layer0_outputs(6228));
    outputs(415) <= layer0_outputs(3679);
    outputs(416) <= not(layer0_outputs(5431));
    outputs(417) <= (layer0_outputs(8745)) and not (layer0_outputs(2603));
    outputs(418) <= not(layer0_outputs(7561));
    outputs(419) <= (layer0_outputs(1362)) and (layer0_outputs(7468));
    outputs(420) <= layer0_outputs(5807);
    outputs(421) <= not(layer0_outputs(2000));
    outputs(422) <= layer0_outputs(6557);
    outputs(423) <= layer0_outputs(4735);
    outputs(424) <= (layer0_outputs(628)) xor (layer0_outputs(3925));
    outputs(425) <= layer0_outputs(845);
    outputs(426) <= not(layer0_outputs(9579));
    outputs(427) <= not(layer0_outputs(8033)) or (layer0_outputs(9874));
    outputs(428) <= layer0_outputs(5746);
    outputs(429) <= layer0_outputs(6938);
    outputs(430) <= not((layer0_outputs(475)) and (layer0_outputs(3567)));
    outputs(431) <= not(layer0_outputs(4357));
    outputs(432) <= not(layer0_outputs(9406));
    outputs(433) <= not((layer0_outputs(8641)) xor (layer0_outputs(8661)));
    outputs(434) <= not((layer0_outputs(2643)) and (layer0_outputs(9422)));
    outputs(435) <= not((layer0_outputs(2815)) and (layer0_outputs(6364)));
    outputs(436) <= (layer0_outputs(967)) xor (layer0_outputs(10202));
    outputs(437) <= layer0_outputs(6465);
    outputs(438) <= not((layer0_outputs(4533)) xor (layer0_outputs(4327)));
    outputs(439) <= not((layer0_outputs(3842)) and (layer0_outputs(2364)));
    outputs(440) <= layer0_outputs(61);
    outputs(441) <= not(layer0_outputs(1795)) or (layer0_outputs(6889));
    outputs(442) <= layer0_outputs(3882);
    outputs(443) <= layer0_outputs(9555);
    outputs(444) <= (layer0_outputs(6975)) xor (layer0_outputs(6350));
    outputs(445) <= (layer0_outputs(4492)) and not (layer0_outputs(8846));
    outputs(446) <= not(layer0_outputs(5130));
    outputs(447) <= not(layer0_outputs(6264));
    outputs(448) <= (layer0_outputs(4474)) and not (layer0_outputs(7254));
    outputs(449) <= not(layer0_outputs(9318)) or (layer0_outputs(4003));
    outputs(450) <= layer0_outputs(1322);
    outputs(451) <= not(layer0_outputs(357));
    outputs(452) <= layer0_outputs(2958);
    outputs(453) <= (layer0_outputs(6613)) and (layer0_outputs(8713));
    outputs(454) <= not(layer0_outputs(2317));
    outputs(455) <= (layer0_outputs(3318)) and not (layer0_outputs(8625));
    outputs(456) <= not((layer0_outputs(9094)) xor (layer0_outputs(6682)));
    outputs(457) <= (layer0_outputs(1907)) and not (layer0_outputs(3921));
    outputs(458) <= not((layer0_outputs(1391)) xor (layer0_outputs(4051)));
    outputs(459) <= not(layer0_outputs(8793));
    outputs(460) <= layer0_outputs(2210);
    outputs(461) <= layer0_outputs(344);
    outputs(462) <= not(layer0_outputs(7824)) or (layer0_outputs(3892));
    outputs(463) <= layer0_outputs(266);
    outputs(464) <= not(layer0_outputs(9531)) or (layer0_outputs(688));
    outputs(465) <= layer0_outputs(2157);
    outputs(466) <= not(layer0_outputs(5783));
    outputs(467) <= layer0_outputs(6533);
    outputs(468) <= not((layer0_outputs(877)) and (layer0_outputs(121)));
    outputs(469) <= layer0_outputs(2062);
    outputs(470) <= (layer0_outputs(5681)) xor (layer0_outputs(9596));
    outputs(471) <= not((layer0_outputs(6328)) xor (layer0_outputs(6102)));
    outputs(472) <= not(layer0_outputs(5561));
    outputs(473) <= layer0_outputs(4509);
    outputs(474) <= (layer0_outputs(5587)) or (layer0_outputs(2631));
    outputs(475) <= (layer0_outputs(3178)) xor (layer0_outputs(1928));
    outputs(476) <= (layer0_outputs(8456)) and not (layer0_outputs(3404));
    outputs(477) <= not(layer0_outputs(2808)) or (layer0_outputs(1488));
    outputs(478) <= layer0_outputs(1163);
    outputs(479) <= (layer0_outputs(2297)) xor (layer0_outputs(8951));
    outputs(480) <= not((layer0_outputs(2376)) xor (layer0_outputs(1004)));
    outputs(481) <= not(layer0_outputs(3730));
    outputs(482) <= not(layer0_outputs(1176)) or (layer0_outputs(6177));
    outputs(483) <= not(layer0_outputs(593));
    outputs(484) <= not((layer0_outputs(2994)) xor (layer0_outputs(7571)));
    outputs(485) <= (layer0_outputs(10013)) and (layer0_outputs(2904));
    outputs(486) <= not(layer0_outputs(6399));
    outputs(487) <= not(layer0_outputs(2595)) or (layer0_outputs(8732));
    outputs(488) <= not(layer0_outputs(6228));
    outputs(489) <= not(layer0_outputs(9916));
    outputs(490) <= (layer0_outputs(3382)) and not (layer0_outputs(2734));
    outputs(491) <= not(layer0_outputs(8550));
    outputs(492) <= not(layer0_outputs(3232));
    outputs(493) <= (layer0_outputs(3913)) xor (layer0_outputs(9288));
    outputs(494) <= layer0_outputs(7721);
    outputs(495) <= not(layer0_outputs(7660)) or (layer0_outputs(7506));
    outputs(496) <= not(layer0_outputs(7584));
    outputs(497) <= layer0_outputs(10103);
    outputs(498) <= not((layer0_outputs(6320)) xor (layer0_outputs(7430)));
    outputs(499) <= not((layer0_outputs(6400)) and (layer0_outputs(9896)));
    outputs(500) <= not((layer0_outputs(6192)) xor (layer0_outputs(2503)));
    outputs(501) <= layer0_outputs(8714);
    outputs(502) <= (layer0_outputs(4506)) and not (layer0_outputs(37));
    outputs(503) <= not(layer0_outputs(387));
    outputs(504) <= not((layer0_outputs(9640)) or (layer0_outputs(7777)));
    outputs(505) <= (layer0_outputs(4517)) xor (layer0_outputs(5562));
    outputs(506) <= layer0_outputs(5066);
    outputs(507) <= (layer0_outputs(438)) and (layer0_outputs(7026));
    outputs(508) <= (layer0_outputs(6926)) and not (layer0_outputs(1436));
    outputs(509) <= layer0_outputs(977);
    outputs(510) <= not(layer0_outputs(2369)) or (layer0_outputs(974));
    outputs(511) <= not(layer0_outputs(3471)) or (layer0_outputs(5784));
    outputs(512) <= layer0_outputs(1053);
    outputs(513) <= not(layer0_outputs(9096));
    outputs(514) <= (layer0_outputs(1448)) and not (layer0_outputs(1067));
    outputs(515) <= layer0_outputs(10145);
    outputs(516) <= layer0_outputs(8218);
    outputs(517) <= layer0_outputs(7672);
    outputs(518) <= (layer0_outputs(2527)) and not (layer0_outputs(2034));
    outputs(519) <= not((layer0_outputs(1544)) xor (layer0_outputs(6164)));
    outputs(520) <= layer0_outputs(9285);
    outputs(521) <= not((layer0_outputs(3030)) xor (layer0_outputs(705)));
    outputs(522) <= not((layer0_outputs(3184)) or (layer0_outputs(2502)));
    outputs(523) <= layer0_outputs(3634);
    outputs(524) <= not(layer0_outputs(418)) or (layer0_outputs(4790));
    outputs(525) <= not((layer0_outputs(619)) and (layer0_outputs(7826)));
    outputs(526) <= (layer0_outputs(1046)) and not (layer0_outputs(5862));
    outputs(527) <= not(layer0_outputs(4059)) or (layer0_outputs(4683));
    outputs(528) <= layer0_outputs(9473);
    outputs(529) <= layer0_outputs(1146);
    outputs(530) <= (layer0_outputs(6410)) and (layer0_outputs(1288));
    outputs(531) <= layer0_outputs(5809);
    outputs(532) <= not(layer0_outputs(9245)) or (layer0_outputs(9633));
    outputs(533) <= not(layer0_outputs(2579));
    outputs(534) <= not(layer0_outputs(5541));
    outputs(535) <= (layer0_outputs(3903)) xor (layer0_outputs(4763));
    outputs(536) <= layer0_outputs(960);
    outputs(537) <= layer0_outputs(4321);
    outputs(538) <= not(layer0_outputs(9368));
    outputs(539) <= layer0_outputs(796);
    outputs(540) <= (layer0_outputs(7011)) xor (layer0_outputs(6750));
    outputs(541) <= layer0_outputs(8293);
    outputs(542) <= not(layer0_outputs(1767));
    outputs(543) <= not(layer0_outputs(9893)) or (layer0_outputs(2419));
    outputs(544) <= (layer0_outputs(3945)) or (layer0_outputs(219));
    outputs(545) <= not(layer0_outputs(579));
    outputs(546) <= layer0_outputs(5044);
    outputs(547) <= not(layer0_outputs(1655));
    outputs(548) <= not((layer0_outputs(1864)) or (layer0_outputs(9068)));
    outputs(549) <= not((layer0_outputs(10219)) xor (layer0_outputs(2486)));
    outputs(550) <= layer0_outputs(182);
    outputs(551) <= not(layer0_outputs(8746));
    outputs(552) <= (layer0_outputs(9408)) and not (layer0_outputs(205));
    outputs(553) <= not(layer0_outputs(8733));
    outputs(554) <= (layer0_outputs(3384)) xor (layer0_outputs(47));
    outputs(555) <= (layer0_outputs(9776)) and not (layer0_outputs(1820));
    outputs(556) <= layer0_outputs(3320);
    outputs(557) <= layer0_outputs(481);
    outputs(558) <= layer0_outputs(7327);
    outputs(559) <= '1';
    outputs(560) <= layer0_outputs(1772);
    outputs(561) <= not(layer0_outputs(9484)) or (layer0_outputs(8865));
    outputs(562) <= (layer0_outputs(5985)) and (layer0_outputs(5039));
    outputs(563) <= (layer0_outputs(10030)) or (layer0_outputs(2543));
    outputs(564) <= not(layer0_outputs(6512));
    outputs(565) <= layer0_outputs(7141);
    outputs(566) <= not(layer0_outputs(4804));
    outputs(567) <= layer0_outputs(4285);
    outputs(568) <= not(layer0_outputs(3934));
    outputs(569) <= not(layer0_outputs(3537));
    outputs(570) <= not((layer0_outputs(7580)) xor (layer0_outputs(9169)));
    outputs(571) <= not(layer0_outputs(8521));
    outputs(572) <= (layer0_outputs(3086)) xor (layer0_outputs(7211));
    outputs(573) <= (layer0_outputs(7712)) and (layer0_outputs(7605));
    outputs(574) <= not(layer0_outputs(3360));
    outputs(575) <= (layer0_outputs(5068)) or (layer0_outputs(1727));
    outputs(576) <= layer0_outputs(4320);
    outputs(577) <= not((layer0_outputs(5385)) or (layer0_outputs(203)));
    outputs(578) <= not(layer0_outputs(9131)) or (layer0_outputs(1738));
    outputs(579) <= layer0_outputs(9627);
    outputs(580) <= not(layer0_outputs(6776));
    outputs(581) <= not(layer0_outputs(7733));
    outputs(582) <= layer0_outputs(1106);
    outputs(583) <= not(layer0_outputs(2439)) or (layer0_outputs(4867));
    outputs(584) <= not(layer0_outputs(8722)) or (layer0_outputs(263));
    outputs(585) <= not(layer0_outputs(1425));
    outputs(586) <= (layer0_outputs(5313)) and not (layer0_outputs(6919));
    outputs(587) <= layer0_outputs(2300);
    outputs(588) <= not((layer0_outputs(318)) xor (layer0_outputs(9405)));
    outputs(589) <= not(layer0_outputs(4026));
    outputs(590) <= not(layer0_outputs(96));
    outputs(591) <= (layer0_outputs(9785)) or (layer0_outputs(3372));
    outputs(592) <= (layer0_outputs(7705)) and (layer0_outputs(1658));
    outputs(593) <= not(layer0_outputs(7664));
    outputs(594) <= (layer0_outputs(1595)) and not (layer0_outputs(5718));
    outputs(595) <= not((layer0_outputs(8007)) xor (layer0_outputs(7325)));
    outputs(596) <= (layer0_outputs(4205)) xor (layer0_outputs(3705));
    outputs(597) <= layer0_outputs(6434);
    outputs(598) <= layer0_outputs(7520);
    outputs(599) <= layer0_outputs(143);
    outputs(600) <= layer0_outputs(4683);
    outputs(601) <= (layer0_outputs(1917)) xor (layer0_outputs(7719));
    outputs(602) <= not(layer0_outputs(8494));
    outputs(603) <= not((layer0_outputs(4919)) xor (layer0_outputs(10002)));
    outputs(604) <= not(layer0_outputs(8838));
    outputs(605) <= (layer0_outputs(5811)) xor (layer0_outputs(5479));
    outputs(606) <= not(layer0_outputs(7854)) or (layer0_outputs(1477));
    outputs(607) <= (layer0_outputs(10179)) xor (layer0_outputs(9498));
    outputs(608) <= layer0_outputs(7083);
    outputs(609) <= not((layer0_outputs(1061)) xor (layer0_outputs(3040)));
    outputs(610) <= not((layer0_outputs(4196)) and (layer0_outputs(5219)));
    outputs(611) <= not(layer0_outputs(1696));
    outputs(612) <= not((layer0_outputs(7800)) xor (layer0_outputs(2571)));
    outputs(613) <= not((layer0_outputs(1329)) xor (layer0_outputs(6826)));
    outputs(614) <= not(layer0_outputs(2987));
    outputs(615) <= layer0_outputs(7334);
    outputs(616) <= layer0_outputs(419);
    outputs(617) <= layer0_outputs(8921);
    outputs(618) <= not(layer0_outputs(5734));
    outputs(619) <= not((layer0_outputs(5840)) xor (layer0_outputs(9035)));
    outputs(620) <= (layer0_outputs(4820)) and not (layer0_outputs(9501));
    outputs(621) <= (layer0_outputs(7483)) xor (layer0_outputs(3508));
    outputs(622) <= layer0_outputs(5317);
    outputs(623) <= not(layer0_outputs(6398)) or (layer0_outputs(6165));
    outputs(624) <= (layer0_outputs(1857)) or (layer0_outputs(2402));
    outputs(625) <= (layer0_outputs(4065)) or (layer0_outputs(2510));
    outputs(626) <= not(layer0_outputs(9037));
    outputs(627) <= not(layer0_outputs(10076));
    outputs(628) <= not(layer0_outputs(4580));
    outputs(629) <= layer0_outputs(4148);
    outputs(630) <= not(layer0_outputs(614));
    outputs(631) <= layer0_outputs(1353);
    outputs(632) <= not((layer0_outputs(9937)) xor (layer0_outputs(8926)));
    outputs(633) <= not(layer0_outputs(7143)) or (layer0_outputs(6882));
    outputs(634) <= not(layer0_outputs(1033));
    outputs(635) <= layer0_outputs(7016);
    outputs(636) <= not(layer0_outputs(1576));
    outputs(637) <= not(layer0_outputs(881));
    outputs(638) <= not(layer0_outputs(1190));
    outputs(639) <= not(layer0_outputs(1392));
    outputs(640) <= not((layer0_outputs(1631)) xor (layer0_outputs(4436)));
    outputs(641) <= layer0_outputs(9122);
    outputs(642) <= not(layer0_outputs(6310));
    outputs(643) <= layer0_outputs(4717);
    outputs(644) <= layer0_outputs(2515);
    outputs(645) <= not(layer0_outputs(7704)) or (layer0_outputs(9852));
    outputs(646) <= layer0_outputs(3025);
    outputs(647) <= not((layer0_outputs(9493)) or (layer0_outputs(3808)));
    outputs(648) <= not((layer0_outputs(1352)) xor (layer0_outputs(2042)));
    outputs(649) <= layer0_outputs(6892);
    outputs(650) <= (layer0_outputs(7236)) and not (layer0_outputs(4117));
    outputs(651) <= layer0_outputs(781);
    outputs(652) <= not((layer0_outputs(1799)) and (layer0_outputs(9744)));
    outputs(653) <= layer0_outputs(9700);
    outputs(654) <= layer0_outputs(3238);
    outputs(655) <= (layer0_outputs(5472)) xor (layer0_outputs(2448));
    outputs(656) <= not((layer0_outputs(7740)) or (layer0_outputs(6118)));
    outputs(657) <= (layer0_outputs(1574)) xor (layer0_outputs(7901));
    outputs(658) <= not(layer0_outputs(4));
    outputs(659) <= layer0_outputs(6648);
    outputs(660) <= not(layer0_outputs(750));
    outputs(661) <= layer0_outputs(8787);
    outputs(662) <= layer0_outputs(6486);
    outputs(663) <= not((layer0_outputs(4947)) xor (layer0_outputs(7918)));
    outputs(664) <= layer0_outputs(6125);
    outputs(665) <= not((layer0_outputs(5455)) xor (layer0_outputs(8406)));
    outputs(666) <= not(layer0_outputs(4333)) or (layer0_outputs(6007));
    outputs(667) <= not((layer0_outputs(7358)) or (layer0_outputs(6572)));
    outputs(668) <= not(layer0_outputs(6377));
    outputs(669) <= not(layer0_outputs(4325));
    outputs(670) <= not(layer0_outputs(8016));
    outputs(671) <= (layer0_outputs(3165)) and not (layer0_outputs(6116));
    outputs(672) <= not((layer0_outputs(7190)) xor (layer0_outputs(7581)));
    outputs(673) <= not((layer0_outputs(8449)) or (layer0_outputs(348)));
    outputs(674) <= layer0_outputs(3287);
    outputs(675) <= not((layer0_outputs(7400)) and (layer0_outputs(7048)));
    outputs(676) <= not(layer0_outputs(129));
    outputs(677) <= not((layer0_outputs(2872)) or (layer0_outputs(8194)));
    outputs(678) <= layer0_outputs(6480);
    outputs(679) <= (layer0_outputs(6027)) and (layer0_outputs(4337));
    outputs(680) <= not(layer0_outputs(9432)) or (layer0_outputs(9985));
    outputs(681) <= layer0_outputs(1206);
    outputs(682) <= not((layer0_outputs(3107)) xor (layer0_outputs(213)));
    outputs(683) <= not((layer0_outputs(9691)) and (layer0_outputs(4713)));
    outputs(684) <= not(layer0_outputs(9836));
    outputs(685) <= not(layer0_outputs(2834));
    outputs(686) <= not((layer0_outputs(4164)) or (layer0_outputs(10225)));
    outputs(687) <= (layer0_outputs(1384)) xor (layer0_outputs(7388));
    outputs(688) <= not(layer0_outputs(9451));
    outputs(689) <= (layer0_outputs(9544)) or (layer0_outputs(8031));
    outputs(690) <= (layer0_outputs(8387)) xor (layer0_outputs(4687));
    outputs(691) <= layer0_outputs(5075);
    outputs(692) <= (layer0_outputs(3104)) and not (layer0_outputs(5308));
    outputs(693) <= (layer0_outputs(8575)) xor (layer0_outputs(6066));
    outputs(694) <= not((layer0_outputs(3505)) or (layer0_outputs(3366)));
    outputs(695) <= (layer0_outputs(10117)) xor (layer0_outputs(6165));
    outputs(696) <= not(layer0_outputs(1884));
    outputs(697) <= not((layer0_outputs(7744)) and (layer0_outputs(7421)));
    outputs(698) <= layer0_outputs(403);
    outputs(699) <= layer0_outputs(5554);
    outputs(700) <= layer0_outputs(3779);
    outputs(701) <= not(layer0_outputs(7529));
    outputs(702) <= (layer0_outputs(3485)) xor (layer0_outputs(846));
    outputs(703) <= not(layer0_outputs(7836)) or (layer0_outputs(2959));
    outputs(704) <= not((layer0_outputs(458)) xor (layer0_outputs(1864)));
    outputs(705) <= (layer0_outputs(9151)) xor (layer0_outputs(1226));
    outputs(706) <= not(layer0_outputs(9392));
    outputs(707) <= not(layer0_outputs(7577));
    outputs(708) <= (layer0_outputs(2598)) or (layer0_outputs(3450));
    outputs(709) <= layer0_outputs(599);
    outputs(710) <= not(layer0_outputs(3207));
    outputs(711) <= layer0_outputs(1495);
    outputs(712) <= not((layer0_outputs(545)) xor (layer0_outputs(2137)));
    outputs(713) <= not(layer0_outputs(9171));
    outputs(714) <= (layer0_outputs(3364)) xor (layer0_outputs(1267));
    outputs(715) <= layer0_outputs(2415);
    outputs(716) <= not((layer0_outputs(2618)) xor (layer0_outputs(3401)));
    outputs(717) <= not((layer0_outputs(6635)) xor (layer0_outputs(1840)));
    outputs(718) <= not(layer0_outputs(4966)) or (layer0_outputs(1793));
    outputs(719) <= not(layer0_outputs(6144));
    outputs(720) <= not(layer0_outputs(3342));
    outputs(721) <= layer0_outputs(7802);
    outputs(722) <= not(layer0_outputs(5319));
    outputs(723) <= not(layer0_outputs(7072));
    outputs(724) <= not(layer0_outputs(8651));
    outputs(725) <= not((layer0_outputs(9073)) xor (layer0_outputs(8998)));
    outputs(726) <= not(layer0_outputs(2812)) or (layer0_outputs(4197));
    outputs(727) <= not((layer0_outputs(8044)) xor (layer0_outputs(3711)));
    outputs(728) <= not(layer0_outputs(9728));
    outputs(729) <= (layer0_outputs(9416)) xor (layer0_outputs(1707));
    outputs(730) <= not(layer0_outputs(4283));
    outputs(731) <= not(layer0_outputs(5618));
    outputs(732) <= not((layer0_outputs(1054)) or (layer0_outputs(473)));
    outputs(733) <= not(layer0_outputs(711));
    outputs(734) <= not(layer0_outputs(7499));
    outputs(735) <= not(layer0_outputs(5723));
    outputs(736) <= layer0_outputs(6107);
    outputs(737) <= not(layer0_outputs(82));
    outputs(738) <= not(layer0_outputs(7456));
    outputs(739) <= layer0_outputs(3564);
    outputs(740) <= not(layer0_outputs(3660));
    outputs(741) <= layer0_outputs(1195);
    outputs(742) <= not((layer0_outputs(5794)) xor (layer0_outputs(3824)));
    outputs(743) <= layer0_outputs(8298);
    outputs(744) <= not(layer0_outputs(4391));
    outputs(745) <= not(layer0_outputs(4444));
    outputs(746) <= layer0_outputs(484);
    outputs(747) <= not(layer0_outputs(3661)) or (layer0_outputs(7073));
    outputs(748) <= layer0_outputs(3143);
    outputs(749) <= not((layer0_outputs(840)) xor (layer0_outputs(1471)));
    outputs(750) <= not(layer0_outputs(8373)) or (layer0_outputs(4022));
    outputs(751) <= layer0_outputs(7098);
    outputs(752) <= layer0_outputs(2928);
    outputs(753) <= not(layer0_outputs(2036));
    outputs(754) <= (layer0_outputs(7119)) or (layer0_outputs(1150));
    outputs(755) <= not(layer0_outputs(8396));
    outputs(756) <= not(layer0_outputs(6212));
    outputs(757) <= layer0_outputs(4199);
    outputs(758) <= not(layer0_outputs(6669)) or (layer0_outputs(402));
    outputs(759) <= (layer0_outputs(7365)) and not (layer0_outputs(7336));
    outputs(760) <= '1';
    outputs(761) <= not((layer0_outputs(5654)) xor (layer0_outputs(5001)));
    outputs(762) <= not(layer0_outputs(5653));
    outputs(763) <= layer0_outputs(9553);
    outputs(764) <= not((layer0_outputs(6420)) xor (layer0_outputs(2911)));
    outputs(765) <= not(layer0_outputs(4162));
    outputs(766) <= not(layer0_outputs(7999));
    outputs(767) <= (layer0_outputs(2713)) and not (layer0_outputs(2060));
    outputs(768) <= not(layer0_outputs(1217)) or (layer0_outputs(10064));
    outputs(769) <= layer0_outputs(120);
    outputs(770) <= not((layer0_outputs(9308)) xor (layer0_outputs(7722)));
    outputs(771) <= not(layer0_outputs(7749));
    outputs(772) <= not((layer0_outputs(3534)) xor (layer0_outputs(6721)));
    outputs(773) <= not(layer0_outputs(9781));
    outputs(774) <= layer0_outputs(3397);
    outputs(775) <= (layer0_outputs(2172)) and (layer0_outputs(5732));
    outputs(776) <= (layer0_outputs(10132)) and (layer0_outputs(2216));
    outputs(777) <= layer0_outputs(4036);
    outputs(778) <= not((layer0_outputs(4968)) xor (layer0_outputs(1835)));
    outputs(779) <= layer0_outputs(4226);
    outputs(780) <= (layer0_outputs(6380)) xor (layer0_outputs(9851));
    outputs(781) <= not(layer0_outputs(6958));
    outputs(782) <= not(layer0_outputs(3298)) or (layer0_outputs(5727));
    outputs(783) <= layer0_outputs(4712);
    outputs(784) <= (layer0_outputs(6286)) and not (layer0_outputs(5523));
    outputs(785) <= layer0_outputs(6589);
    outputs(786) <= not(layer0_outputs(7926));
    outputs(787) <= not(layer0_outputs(3476));
    outputs(788) <= not(layer0_outputs(5353));
    outputs(789) <= not(layer0_outputs(1896));
    outputs(790) <= not(layer0_outputs(9259));
    outputs(791) <= (layer0_outputs(726)) and not (layer0_outputs(2338));
    outputs(792) <= not((layer0_outputs(1688)) xor (layer0_outputs(3749)));
    outputs(793) <= (layer0_outputs(1738)) or (layer0_outputs(8882));
    outputs(794) <= not((layer0_outputs(8032)) xor (layer0_outputs(799)));
    outputs(795) <= layer0_outputs(6164);
    outputs(796) <= (layer0_outputs(3707)) and not (layer0_outputs(9182));
    outputs(797) <= '1';
    outputs(798) <= (layer0_outputs(5842)) and not (layer0_outputs(2592));
    outputs(799) <= not(layer0_outputs(2381));
    outputs(800) <= not(layer0_outputs(6242));
    outputs(801) <= layer0_outputs(2817);
    outputs(802) <= (layer0_outputs(7814)) and not (layer0_outputs(1828));
    outputs(803) <= not((layer0_outputs(7859)) xor (layer0_outputs(5001)));
    outputs(804) <= not(layer0_outputs(356));
    outputs(805) <= not(layer0_outputs(6479));
    outputs(806) <= layer0_outputs(388);
    outputs(807) <= layer0_outputs(2847);
    outputs(808) <= not((layer0_outputs(5315)) xor (layer0_outputs(9355)));
    outputs(809) <= not(layer0_outputs(8812));
    outputs(810) <= not((layer0_outputs(7490)) xor (layer0_outputs(6543)));
    outputs(811) <= (layer0_outputs(4465)) and not (layer0_outputs(7484));
    outputs(812) <= layer0_outputs(5467);
    outputs(813) <= (layer0_outputs(3899)) or (layer0_outputs(7220));
    outputs(814) <= not(layer0_outputs(5899));
    outputs(815) <= layer0_outputs(4273);
    outputs(816) <= (layer0_outputs(6197)) xor (layer0_outputs(1121));
    outputs(817) <= not(layer0_outputs(6435));
    outputs(818) <= layer0_outputs(1833);
    outputs(819) <= not(layer0_outputs(10201));
    outputs(820) <= not((layer0_outputs(2992)) xor (layer0_outputs(6480)));
    outputs(821) <= not(layer0_outputs(8466));
    outputs(822) <= not(layer0_outputs(4627)) or (layer0_outputs(277));
    outputs(823) <= not((layer0_outputs(1898)) and (layer0_outputs(4548)));
    outputs(824) <= (layer0_outputs(5400)) and (layer0_outputs(4915));
    outputs(825) <= not(layer0_outputs(3067)) or (layer0_outputs(5749));
    outputs(826) <= (layer0_outputs(2977)) or (layer0_outputs(3055));
    outputs(827) <= layer0_outputs(9894);
    outputs(828) <= not((layer0_outputs(5675)) and (layer0_outputs(4675)));
    outputs(829) <= not((layer0_outputs(910)) or (layer0_outputs(5346)));
    outputs(830) <= (layer0_outputs(9420)) xor (layer0_outputs(4981));
    outputs(831) <= layer0_outputs(3196);
    outputs(832) <= not(layer0_outputs(8634)) or (layer0_outputs(2146));
    outputs(833) <= not((layer0_outputs(9228)) or (layer0_outputs(5118)));
    outputs(834) <= layer0_outputs(5274);
    outputs(835) <= (layer0_outputs(1357)) and not (layer0_outputs(6078));
    outputs(836) <= not(layer0_outputs(8857));
    outputs(837) <= not((layer0_outputs(5488)) and (layer0_outputs(4007)));
    outputs(838) <= not(layer0_outputs(2122));
    outputs(839) <= not(layer0_outputs(7741));
    outputs(840) <= not(layer0_outputs(8723));
    outputs(841) <= not(layer0_outputs(3255)) or (layer0_outputs(1816));
    outputs(842) <= layer0_outputs(2699);
    outputs(843) <= not((layer0_outputs(3358)) or (layer0_outputs(3353)));
    outputs(844) <= not(layer0_outputs(9413));
    outputs(845) <= (layer0_outputs(6119)) and not (layer0_outputs(5604));
    outputs(846) <= not(layer0_outputs(1154)) or (layer0_outputs(9389));
    outputs(847) <= not(layer0_outputs(1650));
    outputs(848) <= layer0_outputs(7239);
    outputs(849) <= (layer0_outputs(1266)) and (layer0_outputs(9052));
    outputs(850) <= layer0_outputs(3523);
    outputs(851) <= layer0_outputs(359);
    outputs(852) <= layer0_outputs(8774);
    outputs(853) <= not((layer0_outputs(699)) xor (layer0_outputs(1196)));
    outputs(854) <= not(layer0_outputs(5047));
    outputs(855) <= not(layer0_outputs(1997));
    outputs(856) <= not(layer0_outputs(4392));
    outputs(857) <= not((layer0_outputs(5406)) and (layer0_outputs(4612)));
    outputs(858) <= not(layer0_outputs(4406));
    outputs(859) <= not(layer0_outputs(6916));
    outputs(860) <= not((layer0_outputs(7397)) or (layer0_outputs(4154)));
    outputs(861) <= layer0_outputs(5508);
    outputs(862) <= not(layer0_outputs(9648));
    outputs(863) <= not(layer0_outputs(6804));
    outputs(864) <= layer0_outputs(6840);
    outputs(865) <= not((layer0_outputs(10071)) xor (layer0_outputs(9445)));
    outputs(866) <= layer0_outputs(9830);
    outputs(867) <= layer0_outputs(4980);
    outputs(868) <= layer0_outputs(259);
    outputs(869) <= layer0_outputs(9575);
    outputs(870) <= not(layer0_outputs(4593));
    outputs(871) <= (layer0_outputs(4685)) and (layer0_outputs(5902));
    outputs(872) <= not((layer0_outputs(1305)) or (layer0_outputs(6658)));
    outputs(873) <= layer0_outputs(4556);
    outputs(874) <= layer0_outputs(6528);
    outputs(875) <= not((layer0_outputs(622)) xor (layer0_outputs(5089)));
    outputs(876) <= (layer0_outputs(7576)) and not (layer0_outputs(7544));
    outputs(877) <= not((layer0_outputs(3586)) xor (layer0_outputs(6643)));
    outputs(878) <= (layer0_outputs(1688)) and not (layer0_outputs(152));
    outputs(879) <= not(layer0_outputs(1672)) or (layer0_outputs(616));
    outputs(880) <= (layer0_outputs(6932)) or (layer0_outputs(5631));
    outputs(881) <= not(layer0_outputs(139)) or (layer0_outputs(6884));
    outputs(882) <= not(layer0_outputs(1402));
    outputs(883) <= layer0_outputs(2908);
    outputs(884) <= layer0_outputs(8728);
    outputs(885) <= not(layer0_outputs(5561)) or (layer0_outputs(6611));
    outputs(886) <= not(layer0_outputs(160));
    outputs(887) <= layer0_outputs(3337);
    outputs(888) <= not(layer0_outputs(9383));
    outputs(889) <= (layer0_outputs(7242)) and (layer0_outputs(9389));
    outputs(890) <= not(layer0_outputs(8887));
    outputs(891) <= not(layer0_outputs(5381));
    outputs(892) <= not((layer0_outputs(4364)) xor (layer0_outputs(3799)));
    outputs(893) <= layer0_outputs(4522);
    outputs(894) <= layer0_outputs(155);
    outputs(895) <= not((layer0_outputs(3215)) and (layer0_outputs(1763)));
    outputs(896) <= layer0_outputs(5882);
    outputs(897) <= layer0_outputs(9569);
    outputs(898) <= layer0_outputs(7178);
    outputs(899) <= not(layer0_outputs(2209));
    outputs(900) <= (layer0_outputs(3841)) xor (layer0_outputs(340));
    outputs(901) <= not((layer0_outputs(7897)) or (layer0_outputs(478)));
    outputs(902) <= not(layer0_outputs(6248));
    outputs(903) <= not((layer0_outputs(10189)) xor (layer0_outputs(180)));
    outputs(904) <= (layer0_outputs(6744)) xor (layer0_outputs(2368));
    outputs(905) <= (layer0_outputs(2857)) xor (layer0_outputs(4000));
    outputs(906) <= not((layer0_outputs(9712)) xor (layer0_outputs(5389)));
    outputs(907) <= layer0_outputs(4321);
    outputs(908) <= (layer0_outputs(2222)) xor (layer0_outputs(6387));
    outputs(909) <= not((layer0_outputs(3073)) and (layer0_outputs(6470)));
    outputs(910) <= layer0_outputs(9019);
    outputs(911) <= not(layer0_outputs(7410));
    outputs(912) <= (layer0_outputs(4636)) xor (layer0_outputs(3583));
    outputs(913) <= not(layer0_outputs(3825)) or (layer0_outputs(7006));
    outputs(914) <= layer0_outputs(8811);
    outputs(915) <= (layer0_outputs(5078)) and not (layer0_outputs(7862));
    outputs(916) <= (layer0_outputs(7275)) and (layer0_outputs(2693));
    outputs(917) <= layer0_outputs(4284);
    outputs(918) <= not(layer0_outputs(2420)) or (layer0_outputs(2457));
    outputs(919) <= (layer0_outputs(3572)) xor (layer0_outputs(6506));
    outputs(920) <= layer0_outputs(1113);
    outputs(921) <= not(layer0_outputs(7225));
    outputs(922) <= layer0_outputs(331);
    outputs(923) <= not(layer0_outputs(4578));
    outputs(924) <= not(layer0_outputs(7568));
    outputs(925) <= layer0_outputs(317);
    outputs(926) <= (layer0_outputs(2870)) and not (layer0_outputs(8114));
    outputs(927) <= '1';
    outputs(928) <= layer0_outputs(2017);
    outputs(929) <= not((layer0_outputs(6514)) and (layer0_outputs(1722)));
    outputs(930) <= not(layer0_outputs(8365));
    outputs(931) <= not(layer0_outputs(3864));
    outputs(932) <= not(layer0_outputs(8642));
    outputs(933) <= not(layer0_outputs(3221));
    outputs(934) <= (layer0_outputs(3877)) xor (layer0_outputs(6590));
    outputs(935) <= not((layer0_outputs(5363)) and (layer0_outputs(941)));
    outputs(936) <= not((layer0_outputs(9301)) or (layer0_outputs(3958)));
    outputs(937) <= not(layer0_outputs(336));
    outputs(938) <= (layer0_outputs(4388)) and not (layer0_outputs(1487));
    outputs(939) <= not(layer0_outputs(3089));
    outputs(940) <= not((layer0_outputs(7966)) or (layer0_outputs(6879)));
    outputs(941) <= (layer0_outputs(7137)) or (layer0_outputs(9152));
    outputs(942) <= not((layer0_outputs(4228)) or (layer0_outputs(1695)));
    outputs(943) <= (layer0_outputs(2075)) xor (layer0_outputs(5088));
    outputs(944) <= (layer0_outputs(1210)) xor (layer0_outputs(6727));
    outputs(945) <= not(layer0_outputs(2694));
    outputs(946) <= (layer0_outputs(8617)) and not (layer0_outputs(3208));
    outputs(947) <= (layer0_outputs(9616)) and (layer0_outputs(6283));
    outputs(948) <= (layer0_outputs(3075)) xor (layer0_outputs(1664));
    outputs(949) <= layer0_outputs(6562);
    outputs(950) <= not(layer0_outputs(2531)) or (layer0_outputs(721));
    outputs(951) <= not(layer0_outputs(6935)) or (layer0_outputs(140));
    outputs(952) <= (layer0_outputs(604)) xor (layer0_outputs(9361));
    outputs(953) <= layer0_outputs(1434);
    outputs(954) <= layer0_outputs(3243);
    outputs(955) <= not(layer0_outputs(395));
    outputs(956) <= layer0_outputs(3320);
    outputs(957) <= not((layer0_outputs(3322)) xor (layer0_outputs(3035)));
    outputs(958) <= not(layer0_outputs(6057));
    outputs(959) <= (layer0_outputs(806)) and not (layer0_outputs(2671));
    outputs(960) <= layer0_outputs(4170);
    outputs(961) <= layer0_outputs(3488);
    outputs(962) <= (layer0_outputs(2824)) or (layer0_outputs(6027));
    outputs(963) <= layer0_outputs(9524);
    outputs(964) <= not(layer0_outputs(6203)) or (layer0_outputs(3332));
    outputs(965) <= not((layer0_outputs(725)) xor (layer0_outputs(4529)));
    outputs(966) <= layer0_outputs(328);
    outputs(967) <= (layer0_outputs(3997)) and not (layer0_outputs(3206));
    outputs(968) <= not((layer0_outputs(5538)) or (layer0_outputs(2179)));
    outputs(969) <= not(layer0_outputs(5109));
    outputs(970) <= not((layer0_outputs(6422)) xor (layer0_outputs(8188)));
    outputs(971) <= not(layer0_outputs(971));
    outputs(972) <= (layer0_outputs(7787)) xor (layer0_outputs(9429));
    outputs(973) <= not((layer0_outputs(7449)) xor (layer0_outputs(8020)));
    outputs(974) <= layer0_outputs(9764);
    outputs(975) <= (layer0_outputs(3210)) and not (layer0_outputs(1516));
    outputs(976) <= not((layer0_outputs(1538)) or (layer0_outputs(6319)));
    outputs(977) <= not(layer0_outputs(4835)) or (layer0_outputs(1869));
    outputs(978) <= not((layer0_outputs(2779)) xor (layer0_outputs(9027)));
    outputs(979) <= layer0_outputs(4698);
    outputs(980) <= layer0_outputs(5152);
    outputs(981) <= (layer0_outputs(8448)) and (layer0_outputs(1687));
    outputs(982) <= (layer0_outputs(1882)) or (layer0_outputs(5828));
    outputs(983) <= not(layer0_outputs(1995)) or (layer0_outputs(7849));
    outputs(984) <= not(layer0_outputs(874));
    outputs(985) <= not(layer0_outputs(9426)) or (layer0_outputs(6304));
    outputs(986) <= (layer0_outputs(8595)) xor (layer0_outputs(9821));
    outputs(987) <= layer0_outputs(3449);
    outputs(988) <= not(layer0_outputs(7465));
    outputs(989) <= not(layer0_outputs(8698));
    outputs(990) <= not((layer0_outputs(445)) or (layer0_outputs(4338)));
    outputs(991) <= (layer0_outputs(4707)) and not (layer0_outputs(1181));
    outputs(992) <= not(layer0_outputs(5222));
    outputs(993) <= not((layer0_outputs(1410)) xor (layer0_outputs(810)));
    outputs(994) <= not(layer0_outputs(4096));
    outputs(995) <= layer0_outputs(5382);
    outputs(996) <= layer0_outputs(5902);
    outputs(997) <= (layer0_outputs(3196)) and (layer0_outputs(7437));
    outputs(998) <= not(layer0_outputs(4598));
    outputs(999) <= not((layer0_outputs(1186)) or (layer0_outputs(2734)));
    outputs(1000) <= (layer0_outputs(1731)) and not (layer0_outputs(6978));
    outputs(1001) <= (layer0_outputs(5678)) xor (layer0_outputs(9390));
    outputs(1002) <= layer0_outputs(311);
    outputs(1003) <= layer0_outputs(7975);
    outputs(1004) <= not(layer0_outputs(5174));
    outputs(1005) <= not(layer0_outputs(7263));
    outputs(1006) <= layer0_outputs(1042);
    outputs(1007) <= layer0_outputs(408);
    outputs(1008) <= not(layer0_outputs(429)) or (layer0_outputs(7846));
    outputs(1009) <= (layer0_outputs(4400)) or (layer0_outputs(8129));
    outputs(1010) <= not((layer0_outputs(6745)) and (layer0_outputs(4936)));
    outputs(1011) <= not(layer0_outputs(4599)) or (layer0_outputs(570));
    outputs(1012) <= not((layer0_outputs(4628)) or (layer0_outputs(7419)));
    outputs(1013) <= (layer0_outputs(1099)) xor (layer0_outputs(4770));
    outputs(1014) <= not((layer0_outputs(7678)) and (layer0_outputs(6800)));
    outputs(1015) <= layer0_outputs(9761);
    outputs(1016) <= not(layer0_outputs(5425));
    outputs(1017) <= (layer0_outputs(2505)) and not (layer0_outputs(10155));
    outputs(1018) <= not(layer0_outputs(3494));
    outputs(1019) <= not(layer0_outputs(7161));
    outputs(1020) <= layer0_outputs(471);
    outputs(1021) <= layer0_outputs(10191);
    outputs(1022) <= layer0_outputs(1741);
    outputs(1023) <= not(layer0_outputs(6929));
    outputs(1024) <= layer0_outputs(7757);
    outputs(1025) <= (layer0_outputs(7207)) and not (layer0_outputs(1618));
    outputs(1026) <= (layer0_outputs(9268)) and not (layer0_outputs(1400));
    outputs(1027) <= (layer0_outputs(3370)) and (layer0_outputs(4192));
    outputs(1028) <= not(layer0_outputs(9277));
    outputs(1029) <= (layer0_outputs(4271)) and (layer0_outputs(5262));
    outputs(1030) <= not((layer0_outputs(1491)) or (layer0_outputs(5373)));
    outputs(1031) <= (layer0_outputs(10115)) and not (layer0_outputs(4060));
    outputs(1032) <= (layer0_outputs(6852)) and not (layer0_outputs(9793));
    outputs(1033) <= not((layer0_outputs(7354)) or (layer0_outputs(5110)));
    outputs(1034) <= (layer0_outputs(3920)) and not (layer0_outputs(310));
    outputs(1035) <= not((layer0_outputs(3688)) or (layer0_outputs(4536)));
    outputs(1036) <= (layer0_outputs(5936)) and (layer0_outputs(10120));
    outputs(1037) <= not((layer0_outputs(59)) xor (layer0_outputs(7110)));
    outputs(1038) <= (layer0_outputs(10224)) and not (layer0_outputs(6034));
    outputs(1039) <= (layer0_outputs(5968)) and not (layer0_outputs(5757));
    outputs(1040) <= not((layer0_outputs(9706)) or (layer0_outputs(6530)));
    outputs(1041) <= (layer0_outputs(7853)) and not (layer0_outputs(3142));
    outputs(1042) <= (layer0_outputs(7635)) and (layer0_outputs(7267));
    outputs(1043) <= (layer0_outputs(5360)) and (layer0_outputs(1193));
    outputs(1044) <= layer0_outputs(4320);
    outputs(1045) <= (layer0_outputs(9475)) and (layer0_outputs(6094));
    outputs(1046) <= layer0_outputs(4546);
    outputs(1047) <= (layer0_outputs(6344)) and not (layer0_outputs(6518));
    outputs(1048) <= layer0_outputs(843);
    outputs(1049) <= (layer0_outputs(2173)) and not (layer0_outputs(8418));
    outputs(1050) <= not((layer0_outputs(3226)) xor (layer0_outputs(5223)));
    outputs(1051) <= (layer0_outputs(6537)) and not (layer0_outputs(9953));
    outputs(1052) <= (layer0_outputs(4261)) xor (layer0_outputs(3340));
    outputs(1053) <= (layer0_outputs(6470)) xor (layer0_outputs(6867));
    outputs(1054) <= (layer0_outputs(3000)) xor (layer0_outputs(8965));
    outputs(1055) <= (layer0_outputs(1747)) and (layer0_outputs(9112));
    outputs(1056) <= not(layer0_outputs(6184));
    outputs(1057) <= not((layer0_outputs(762)) or (layer0_outputs(3145)));
    outputs(1058) <= not((layer0_outputs(2548)) or (layer0_outputs(879)));
    outputs(1059) <= '0';
    outputs(1060) <= not((layer0_outputs(4796)) xor (layer0_outputs(7293)));
    outputs(1061) <= layer0_outputs(9431);
    outputs(1062) <= (layer0_outputs(10213)) and not (layer0_outputs(6903));
    outputs(1063) <= not((layer0_outputs(6371)) and (layer0_outputs(3479)));
    outputs(1064) <= '0';
    outputs(1065) <= (layer0_outputs(2122)) or (layer0_outputs(2355));
    outputs(1066) <= not((layer0_outputs(3323)) or (layer0_outputs(5379)));
    outputs(1067) <= (layer0_outputs(10067)) and (layer0_outputs(1246));
    outputs(1068) <= (layer0_outputs(6004)) xor (layer0_outputs(6660));
    outputs(1069) <= (layer0_outputs(936)) and not (layer0_outputs(2732));
    outputs(1070) <= (layer0_outputs(9165)) xor (layer0_outputs(8902));
    outputs(1071) <= '0';
    outputs(1072) <= (layer0_outputs(4053)) and (layer0_outputs(6358));
    outputs(1073) <= (layer0_outputs(939)) and (layer0_outputs(9725));
    outputs(1074) <= (layer0_outputs(3234)) and not (layer0_outputs(7962));
    outputs(1075) <= (layer0_outputs(5976)) and (layer0_outputs(3662));
    outputs(1076) <= layer0_outputs(2731);
    outputs(1077) <= layer0_outputs(9162);
    outputs(1078) <= (layer0_outputs(9147)) xor (layer0_outputs(2193));
    outputs(1079) <= not(layer0_outputs(7346));
    outputs(1080) <= (layer0_outputs(2551)) xor (layer0_outputs(1176));
    outputs(1081) <= (layer0_outputs(3131)) and not (layer0_outputs(5253));
    outputs(1082) <= not((layer0_outputs(9605)) or (layer0_outputs(568)));
    outputs(1083) <= not((layer0_outputs(4819)) or (layer0_outputs(5941)));
    outputs(1084) <= (layer0_outputs(5307)) and not (layer0_outputs(102));
    outputs(1085) <= (layer0_outputs(2672)) and (layer0_outputs(6442));
    outputs(1086) <= not((layer0_outputs(888)) or (layer0_outputs(2860)));
    outputs(1087) <= (layer0_outputs(8659)) and (layer0_outputs(1030));
    outputs(1088) <= (layer0_outputs(8087)) and (layer0_outputs(789));
    outputs(1089) <= layer0_outputs(8201);
    outputs(1090) <= (layer0_outputs(2164)) and (layer0_outputs(1749));
    outputs(1091) <= (layer0_outputs(6025)) and (layer0_outputs(9870));
    outputs(1092) <= layer0_outputs(4524);
    outputs(1093) <= not((layer0_outputs(4732)) xor (layer0_outputs(9453)));
    outputs(1094) <= not(layer0_outputs(7704));
    outputs(1095) <= not((layer0_outputs(5103)) or (layer0_outputs(3393)));
    outputs(1096) <= (layer0_outputs(1932)) and (layer0_outputs(5140));
    outputs(1097) <= layer0_outputs(1394);
    outputs(1098) <= (layer0_outputs(4088)) and not (layer0_outputs(1723));
    outputs(1099) <= not((layer0_outputs(1261)) or (layer0_outputs(7802)));
    outputs(1100) <= layer0_outputs(4087);
    outputs(1101) <= (layer0_outputs(8016)) and (layer0_outputs(1822));
    outputs(1102) <= not(layer0_outputs(2293));
    outputs(1103) <= (layer0_outputs(9976)) xor (layer0_outputs(4993));
    outputs(1104) <= not((layer0_outputs(176)) or (layer0_outputs(4437)));
    outputs(1105) <= layer0_outputs(5372);
    outputs(1106) <= not(layer0_outputs(4737));
    outputs(1107) <= (layer0_outputs(8612)) and not (layer0_outputs(4889));
    outputs(1108) <= not((layer0_outputs(4522)) or (layer0_outputs(3995)));
    outputs(1109) <= layer0_outputs(6227);
    outputs(1110) <= (layer0_outputs(1294)) and not (layer0_outputs(3699));
    outputs(1111) <= layer0_outputs(8767);
    outputs(1112) <= not(layer0_outputs(1969));
    outputs(1113) <= (layer0_outputs(8029)) and not (layer0_outputs(6121));
    outputs(1114) <= not(layer0_outputs(6343));
    outputs(1115) <= (layer0_outputs(2351)) and not (layer0_outputs(3258));
    outputs(1116) <= not((layer0_outputs(6174)) or (layer0_outputs(1815)));
    outputs(1117) <= not((layer0_outputs(2103)) xor (layer0_outputs(4377)));
    outputs(1118) <= not((layer0_outputs(2520)) xor (layer0_outputs(1184)));
    outputs(1119) <= layer0_outputs(5340);
    outputs(1120) <= (layer0_outputs(9146)) and not (layer0_outputs(6071));
    outputs(1121) <= (layer0_outputs(9237)) and not (layer0_outputs(4538));
    outputs(1122) <= layer0_outputs(8097);
    outputs(1123) <= (layer0_outputs(7571)) and (layer0_outputs(8792));
    outputs(1124) <= (layer0_outputs(210)) and not (layer0_outputs(1906));
    outputs(1125) <= not((layer0_outputs(6412)) xor (layer0_outputs(6585)));
    outputs(1126) <= not((layer0_outputs(611)) or (layer0_outputs(10037)));
    outputs(1127) <= (layer0_outputs(2814)) xor (layer0_outputs(670));
    outputs(1128) <= not(layer0_outputs(2033));
    outputs(1129) <= (layer0_outputs(4739)) xor (layer0_outputs(2065));
    outputs(1130) <= (layer0_outputs(3317)) and not (layer0_outputs(3712));
    outputs(1131) <= (layer0_outputs(730)) and not (layer0_outputs(1531));
    outputs(1132) <= (layer0_outputs(9980)) xor (layer0_outputs(3603));
    outputs(1133) <= (layer0_outputs(1121)) and not (layer0_outputs(1453));
    outputs(1134) <= not((layer0_outputs(4844)) or (layer0_outputs(724)));
    outputs(1135) <= not(layer0_outputs(7631));
    outputs(1136) <= (layer0_outputs(3915)) and not (layer0_outputs(5468));
    outputs(1137) <= not((layer0_outputs(8165)) or (layer0_outputs(8897)));
    outputs(1138) <= (layer0_outputs(5028)) and not (layer0_outputs(6519));
    outputs(1139) <= layer0_outputs(3182);
    outputs(1140) <= not(layer0_outputs(7164));
    outputs(1141) <= (layer0_outputs(3738)) or (layer0_outputs(7428));
    outputs(1142) <= not(layer0_outputs(4008));
    outputs(1143) <= (layer0_outputs(4542)) and (layer0_outputs(7629));
    outputs(1144) <= not((layer0_outputs(3867)) or (layer0_outputs(7658)));
    outputs(1145) <= not((layer0_outputs(7442)) xor (layer0_outputs(350)));
    outputs(1146) <= (layer0_outputs(8541)) and (layer0_outputs(7439));
    outputs(1147) <= not(layer0_outputs(239)) or (layer0_outputs(1532));
    outputs(1148) <= not((layer0_outputs(1792)) xor (layer0_outputs(2581)));
    outputs(1149) <= (layer0_outputs(6798)) and (layer0_outputs(5438));
    outputs(1150) <= (layer0_outputs(6588)) and not (layer0_outputs(3816));
    outputs(1151) <= (layer0_outputs(9533)) and not (layer0_outputs(3910));
    outputs(1152) <= (layer0_outputs(2345)) and not (layer0_outputs(5301));
    outputs(1153) <= not(layer0_outputs(3504));
    outputs(1154) <= not(layer0_outputs(7498));
    outputs(1155) <= not((layer0_outputs(8375)) or (layer0_outputs(1716)));
    outputs(1156) <= (layer0_outputs(5334)) and not (layer0_outputs(1492));
    outputs(1157) <= not(layer0_outputs(2233));
    outputs(1158) <= (layer0_outputs(7430)) xor (layer0_outputs(5465));
    outputs(1159) <= (layer0_outputs(3052)) and not (layer0_outputs(3926));
    outputs(1160) <= layer0_outputs(6372);
    outputs(1161) <= not((layer0_outputs(3473)) or (layer0_outputs(6894)));
    outputs(1162) <= (layer0_outputs(5971)) and (layer0_outputs(3406));
    outputs(1163) <= (layer0_outputs(9529)) and (layer0_outputs(4611));
    outputs(1164) <= (layer0_outputs(5409)) and not (layer0_outputs(717));
    outputs(1165) <= not((layer0_outputs(1010)) or (layer0_outputs(306)));
    outputs(1166) <= not(layer0_outputs(2664));
    outputs(1167) <= (layer0_outputs(3984)) and (layer0_outputs(10051));
    outputs(1168) <= (layer0_outputs(3750)) and not (layer0_outputs(4775));
    outputs(1169) <= not(layer0_outputs(8615));
    outputs(1170) <= (layer0_outputs(6441)) and (layer0_outputs(8103));
    outputs(1171) <= (layer0_outputs(2516)) and not (layer0_outputs(6812));
    outputs(1172) <= not(layer0_outputs(10001));
    outputs(1173) <= not((layer0_outputs(7351)) or (layer0_outputs(9275)));
    outputs(1174) <= not(layer0_outputs(7727));
    outputs(1175) <= (layer0_outputs(8837)) and not (layer0_outputs(2072));
    outputs(1176) <= layer0_outputs(9354);
    outputs(1177) <= not(layer0_outputs(6880));
    outputs(1178) <= (layer0_outputs(6259)) xor (layer0_outputs(2164));
    outputs(1179) <= (layer0_outputs(2493)) and not (layer0_outputs(9552));
    outputs(1180) <= not((layer0_outputs(3442)) xor (layer0_outputs(3830)));
    outputs(1181) <= (layer0_outputs(4929)) and not (layer0_outputs(7218));
    outputs(1182) <= layer0_outputs(9858);
    outputs(1183) <= not(layer0_outputs(449));
    outputs(1184) <= not((layer0_outputs(8189)) or (layer0_outputs(9793)));
    outputs(1185) <= not(layer0_outputs(2768));
    outputs(1186) <= not((layer0_outputs(1684)) xor (layer0_outputs(188)));
    outputs(1187) <= (layer0_outputs(6252)) xor (layer0_outputs(1733));
    outputs(1188) <= layer0_outputs(1067);
    outputs(1189) <= not((layer0_outputs(601)) xor (layer0_outputs(3361)));
    outputs(1190) <= layer0_outputs(2604);
    outputs(1191) <= not(layer0_outputs(7343));
    outputs(1192) <= (layer0_outputs(8648)) and not (layer0_outputs(3636));
    outputs(1193) <= layer0_outputs(10215);
    outputs(1194) <= (layer0_outputs(1514)) and (layer0_outputs(7835));
    outputs(1195) <= (layer0_outputs(1103)) and not (layer0_outputs(510));
    outputs(1196) <= (layer0_outputs(6949)) and not (layer0_outputs(2370));
    outputs(1197) <= (layer0_outputs(1170)) and (layer0_outputs(5299));
    outputs(1198) <= not((layer0_outputs(1921)) or (layer0_outputs(6147)));
    outputs(1199) <= (layer0_outputs(5773)) and not (layer0_outputs(7064));
    outputs(1200) <= (layer0_outputs(2061)) and not (layer0_outputs(3873));
    outputs(1201) <= (layer0_outputs(1108)) and (layer0_outputs(4904));
    outputs(1202) <= not((layer0_outputs(8936)) or (layer0_outputs(1560)));
    outputs(1203) <= (layer0_outputs(4081)) xor (layer0_outputs(9502));
    outputs(1204) <= layer0_outputs(9026);
    outputs(1205) <= (layer0_outputs(5054)) or (layer0_outputs(7590));
    outputs(1206) <= (layer0_outputs(8723)) and (layer0_outputs(5213));
    outputs(1207) <= '0';
    outputs(1208) <= (layer0_outputs(4850)) and not (layer0_outputs(4434));
    outputs(1209) <= (layer0_outputs(6647)) xor (layer0_outputs(3384));
    outputs(1210) <= (layer0_outputs(918)) xor (layer0_outputs(8122));
    outputs(1211) <= not(layer0_outputs(5537));
    outputs(1212) <= (layer0_outputs(7579)) and not (layer0_outputs(2144));
    outputs(1213) <= layer0_outputs(5159);
    outputs(1214) <= (layer0_outputs(1284)) xor (layer0_outputs(4365));
    outputs(1215) <= not((layer0_outputs(2757)) xor (layer0_outputs(1712)));
    outputs(1216) <= (layer0_outputs(575)) and not (layer0_outputs(1962));
    outputs(1217) <= (layer0_outputs(3017)) and not (layer0_outputs(9918));
    outputs(1218) <= layer0_outputs(10167);
    outputs(1219) <= (layer0_outputs(10108)) and not (layer0_outputs(5729));
    outputs(1220) <= (layer0_outputs(3451)) and not (layer0_outputs(2096));
    outputs(1221) <= not(layer0_outputs(1589));
    outputs(1222) <= not(layer0_outputs(8453));
    outputs(1223) <= (layer0_outputs(878)) and not (layer0_outputs(70));
    outputs(1224) <= layer0_outputs(4876);
    outputs(1225) <= not((layer0_outputs(3160)) xor (layer0_outputs(6440)));
    outputs(1226) <= (layer0_outputs(7886)) and (layer0_outputs(2128));
    outputs(1227) <= (layer0_outputs(6324)) and not (layer0_outputs(6290));
    outputs(1228) <= not((layer0_outputs(2134)) xor (layer0_outputs(4669)));
    outputs(1229) <= not(layer0_outputs(8902)) or (layer0_outputs(9201));
    outputs(1230) <= not(layer0_outputs(2991));
    outputs(1231) <= (layer0_outputs(504)) and not (layer0_outputs(9517));
    outputs(1232) <= not((layer0_outputs(6354)) xor (layer0_outputs(1629)));
    outputs(1233) <= (layer0_outputs(3367)) xor (layer0_outputs(4238));
    outputs(1234) <= not((layer0_outputs(9583)) xor (layer0_outputs(7002)));
    outputs(1235) <= not((layer0_outputs(6730)) xor (layer0_outputs(8254)));
    outputs(1236) <= not((layer0_outputs(2288)) xor (layer0_outputs(4295)));
    outputs(1237) <= layer0_outputs(9063);
    outputs(1238) <= (layer0_outputs(3173)) xor (layer0_outputs(8898));
    outputs(1239) <= (layer0_outputs(6970)) and not (layer0_outputs(3952));
    outputs(1240) <= not(layer0_outputs(9514));
    outputs(1241) <= (layer0_outputs(5904)) and not (layer0_outputs(4541));
    outputs(1242) <= not(layer0_outputs(2716));
    outputs(1243) <= not((layer0_outputs(10)) or (layer0_outputs(9312)));
    outputs(1244) <= not((layer0_outputs(6686)) or (layer0_outputs(618)));
    outputs(1245) <= not((layer0_outputs(3724)) or (layer0_outputs(1107)));
    outputs(1246) <= (layer0_outputs(1186)) xor (layer0_outputs(9062));
    outputs(1247) <= (layer0_outputs(3148)) and (layer0_outputs(7924));
    outputs(1248) <= not((layer0_outputs(2033)) or (layer0_outputs(1285)));
    outputs(1249) <= not(layer0_outputs(6244));
    outputs(1250) <= (layer0_outputs(5027)) and not (layer0_outputs(8501));
    outputs(1251) <= (layer0_outputs(1104)) and not (layer0_outputs(586));
    outputs(1252) <= (layer0_outputs(1972)) xor (layer0_outputs(9284));
    outputs(1253) <= not((layer0_outputs(5941)) or (layer0_outputs(4145)));
    outputs(1254) <= not(layer0_outputs(1096));
    outputs(1255) <= (layer0_outputs(5644)) and (layer0_outputs(5692));
    outputs(1256) <= (layer0_outputs(7529)) and (layer0_outputs(7243));
    outputs(1257) <= (layer0_outputs(493)) and not (layer0_outputs(7117));
    outputs(1258) <= not(layer0_outputs(3502));
    outputs(1259) <= (layer0_outputs(5407)) and not (layer0_outputs(6482));
    outputs(1260) <= (layer0_outputs(2795)) xor (layer0_outputs(8243));
    outputs(1261) <= not((layer0_outputs(8398)) xor (layer0_outputs(1782)));
    outputs(1262) <= not(layer0_outputs(228));
    outputs(1263) <= (layer0_outputs(6145)) xor (layer0_outputs(9344));
    outputs(1264) <= (layer0_outputs(4859)) and not (layer0_outputs(275));
    outputs(1265) <= not(layer0_outputs(4211));
    outputs(1266) <= not(layer0_outputs(6446));
    outputs(1267) <= layer0_outputs(1558);
    outputs(1268) <= (layer0_outputs(6699)) and not (layer0_outputs(7679));
    outputs(1269) <= (layer0_outputs(8248)) xor (layer0_outputs(1356));
    outputs(1270) <= layer0_outputs(9594);
    outputs(1271) <= not(layer0_outputs(5731));
    outputs(1272) <= (layer0_outputs(7450)) and not (layer0_outputs(8352));
    outputs(1273) <= not((layer0_outputs(2219)) or (layer0_outputs(4885)));
    outputs(1274) <= (layer0_outputs(6675)) and not (layer0_outputs(9065));
    outputs(1275) <= (layer0_outputs(4726)) and not (layer0_outputs(5883));
    outputs(1276) <= not(layer0_outputs(7814));
    outputs(1277) <= (layer0_outputs(2923)) and not (layer0_outputs(9397));
    outputs(1278) <= (layer0_outputs(6727)) and (layer0_outputs(9993));
    outputs(1279) <= (layer0_outputs(3541)) and (layer0_outputs(7266));
    outputs(1280) <= (layer0_outputs(5269)) and not (layer0_outputs(777));
    outputs(1281) <= (layer0_outputs(6756)) and not (layer0_outputs(3035));
    outputs(1282) <= (layer0_outputs(4429)) and (layer0_outputs(7082));
    outputs(1283) <= (layer0_outputs(5329)) and not (layer0_outputs(1513));
    outputs(1284) <= not(layer0_outputs(8154));
    outputs(1285) <= (layer0_outputs(4016)) and not (layer0_outputs(6985));
    outputs(1286) <= not(layer0_outputs(932));
    outputs(1287) <= not((layer0_outputs(4613)) or (layer0_outputs(3299)));
    outputs(1288) <= (layer0_outputs(4188)) and not (layer0_outputs(10016));
    outputs(1289) <= (layer0_outputs(1671)) and not (layer0_outputs(7139));
    outputs(1290) <= (layer0_outputs(8070)) and (layer0_outputs(4494));
    outputs(1291) <= not(layer0_outputs(10043));
    outputs(1292) <= not((layer0_outputs(9514)) or (layer0_outputs(8957)));
    outputs(1293) <= (layer0_outputs(2759)) and not (layer0_outputs(8581));
    outputs(1294) <= (layer0_outputs(2927)) and (layer0_outputs(7066));
    outputs(1295) <= not((layer0_outputs(9486)) or (layer0_outputs(4911)));
    outputs(1296) <= layer0_outputs(9618);
    outputs(1297) <= not(layer0_outputs(6410));
    outputs(1298) <= (layer0_outputs(5662)) and not (layer0_outputs(7492));
    outputs(1299) <= layer0_outputs(9628);
    outputs(1300) <= layer0_outputs(4040);
    outputs(1301) <= (layer0_outputs(662)) xor (layer0_outputs(4206));
    outputs(1302) <= not((layer0_outputs(8027)) or (layer0_outputs(3756)));
    outputs(1303) <= (layer0_outputs(4675)) and not (layer0_outputs(1385));
    outputs(1304) <= not((layer0_outputs(4012)) xor (layer0_outputs(2749)));
    outputs(1305) <= (layer0_outputs(9117)) and not (layer0_outputs(8654));
    outputs(1306) <= not((layer0_outputs(9721)) and (layer0_outputs(4026)));
    outputs(1307) <= not((layer0_outputs(9456)) xor (layer0_outputs(2544)));
    outputs(1308) <= (layer0_outputs(1617)) and not (layer0_outputs(1314));
    outputs(1309) <= (layer0_outputs(9637)) and not (layer0_outputs(3516));
    outputs(1310) <= not(layer0_outputs(10040));
    outputs(1311) <= (layer0_outputs(856)) and not (layer0_outputs(3697));
    outputs(1312) <= layer0_outputs(3301);
    outputs(1313) <= (layer0_outputs(6853)) and (layer0_outputs(8578));
    outputs(1314) <= '0';
    outputs(1315) <= (layer0_outputs(9885)) and (layer0_outputs(5560));
    outputs(1316) <= (layer0_outputs(9398)) and (layer0_outputs(6713));
    outputs(1317) <= (layer0_outputs(9344)) and not (layer0_outputs(9124));
    outputs(1318) <= not((layer0_outputs(6187)) or (layer0_outputs(207)));
    outputs(1319) <= not((layer0_outputs(1544)) xor (layer0_outputs(32)));
    outputs(1320) <= (layer0_outputs(9092)) xor (layer0_outputs(205));
    outputs(1321) <= (layer0_outputs(9459)) and not (layer0_outputs(2022));
    outputs(1322) <= (layer0_outputs(184)) and not (layer0_outputs(3245));
    outputs(1323) <= (layer0_outputs(5743)) and not (layer0_outputs(1937));
    outputs(1324) <= (layer0_outputs(10095)) xor (layer0_outputs(7652));
    outputs(1325) <= (layer0_outputs(8030)) xor (layer0_outputs(8974));
    outputs(1326) <= (layer0_outputs(6645)) and not (layer0_outputs(42));
    outputs(1327) <= (layer0_outputs(2481)) and not (layer0_outputs(9118));
    outputs(1328) <= not((layer0_outputs(4463)) or (layer0_outputs(175)));
    outputs(1329) <= not((layer0_outputs(8234)) xor (layer0_outputs(7070)));
    outputs(1330) <= (layer0_outputs(9497)) and not (layer0_outputs(2807));
    outputs(1331) <= layer0_outputs(2398);
    outputs(1332) <= (layer0_outputs(250)) and (layer0_outputs(1490));
    outputs(1333) <= not((layer0_outputs(9336)) xor (layer0_outputs(9299)));
    outputs(1334) <= (layer0_outputs(4228)) and not (layer0_outputs(2428));
    outputs(1335) <= (layer0_outputs(8224)) and (layer0_outputs(6736));
    outputs(1336) <= (layer0_outputs(8725)) and (layer0_outputs(6550));
    outputs(1337) <= (layer0_outputs(8377)) and not (layer0_outputs(4662));
    outputs(1338) <= not(layer0_outputs(6498));
    outputs(1339) <= (layer0_outputs(659)) and (layer0_outputs(2212));
    outputs(1340) <= (layer0_outputs(1482)) xor (layer0_outputs(3602));
    outputs(1341) <= (layer0_outputs(6066)) and not (layer0_outputs(2485));
    outputs(1342) <= (layer0_outputs(6073)) xor (layer0_outputs(5911));
    outputs(1343) <= (layer0_outputs(4864)) and not (layer0_outputs(3887));
    outputs(1344) <= not((layer0_outputs(2804)) xor (layer0_outputs(9801)));
    outputs(1345) <= (layer0_outputs(7557)) and not (layer0_outputs(8039));
    outputs(1346) <= not(layer0_outputs(2077));
    outputs(1347) <= not((layer0_outputs(8436)) or (layer0_outputs(7067)));
    outputs(1348) <= (layer0_outputs(1938)) and (layer0_outputs(342));
    outputs(1349) <= (layer0_outputs(8810)) and not (layer0_outputs(2427));
    outputs(1350) <= (layer0_outputs(4648)) and (layer0_outputs(4646));
    outputs(1351) <= (layer0_outputs(8041)) xor (layer0_outputs(3612));
    outputs(1352) <= not((layer0_outputs(6392)) or (layer0_outputs(2456)));
    outputs(1353) <= (layer0_outputs(3497)) and not (layer0_outputs(398));
    outputs(1354) <= not((layer0_outputs(5261)) or (layer0_outputs(5291)));
    outputs(1355) <= (layer0_outputs(4642)) and not (layer0_outputs(3420));
    outputs(1356) <= (layer0_outputs(2765)) xor (layer0_outputs(2097));
    outputs(1357) <= layer0_outputs(5907);
    outputs(1358) <= layer0_outputs(8522);
    outputs(1359) <= not(layer0_outputs(8139));
    outputs(1360) <= (layer0_outputs(8008)) and not (layer0_outputs(4356));
    outputs(1361) <= not(layer0_outputs(5736));
    outputs(1362) <= (layer0_outputs(362)) and not (layer0_outputs(7510));
    outputs(1363) <= (layer0_outputs(7942)) and (layer0_outputs(1926));
    outputs(1364) <= (layer0_outputs(6478)) and (layer0_outputs(7222));
    outputs(1365) <= not(layer0_outputs(6548));
    outputs(1366) <= (layer0_outputs(7384)) and not (layer0_outputs(10025));
    outputs(1367) <= (layer0_outputs(3118)) and not (layer0_outputs(2456));
    outputs(1368) <= (layer0_outputs(5093)) and not (layer0_outputs(7517));
    outputs(1369) <= (layer0_outputs(901)) and not (layer0_outputs(8484));
    outputs(1370) <= (layer0_outputs(6383)) and not (layer0_outputs(2450));
    outputs(1371) <= (layer0_outputs(7646)) and not (layer0_outputs(9213));
    outputs(1372) <= (layer0_outputs(1426)) and not (layer0_outputs(8805));
    outputs(1373) <= (layer0_outputs(8234)) xor (layer0_outputs(3587));
    outputs(1374) <= not((layer0_outputs(2899)) xor (layer0_outputs(3900)));
    outputs(1375) <= (layer0_outputs(5100)) and not (layer0_outputs(3305));
    outputs(1376) <= not((layer0_outputs(9966)) or (layer0_outputs(5760)));
    outputs(1377) <= (layer0_outputs(6140)) and not (layer0_outputs(8257));
    outputs(1378) <= not((layer0_outputs(7233)) or (layer0_outputs(5493)));
    outputs(1379) <= not((layer0_outputs(8014)) or (layer0_outputs(6204)));
    outputs(1380) <= (layer0_outputs(1695)) and not (layer0_outputs(1429));
    outputs(1381) <= (layer0_outputs(4445)) and not (layer0_outputs(655));
    outputs(1382) <= not(layer0_outputs(6384));
    outputs(1383) <= (layer0_outputs(9391)) and (layer0_outputs(8901));
    outputs(1384) <= not((layer0_outputs(1076)) xor (layer0_outputs(7166)));
    outputs(1385) <= (layer0_outputs(2689)) and (layer0_outputs(8716));
    outputs(1386) <= layer0_outputs(3589);
    outputs(1387) <= (layer0_outputs(5302)) xor (layer0_outputs(9016));
    outputs(1388) <= not((layer0_outputs(8714)) or (layer0_outputs(638)));
    outputs(1389) <= (layer0_outputs(3183)) xor (layer0_outputs(2794));
    outputs(1390) <= (layer0_outputs(5119)) and not (layer0_outputs(10035));
    outputs(1391) <= not((layer0_outputs(9922)) xor (layer0_outputs(5638)));
    outputs(1392) <= not((layer0_outputs(9950)) xor (layer0_outputs(6191)));
    outputs(1393) <= (layer0_outputs(1201)) xor (layer0_outputs(3241));
    outputs(1394) <= (layer0_outputs(6823)) and not (layer0_outputs(975));
    outputs(1395) <= (layer0_outputs(2939)) and (layer0_outputs(6274));
    outputs(1396) <= (layer0_outputs(4326)) and (layer0_outputs(4663));
    outputs(1397) <= (layer0_outputs(8730)) and not (layer0_outputs(7292));
    outputs(1398) <= (layer0_outputs(6854)) and not (layer0_outputs(913));
    outputs(1399) <= (layer0_outputs(7222)) or (layer0_outputs(1981));
    outputs(1400) <= (layer0_outputs(4589)) and (layer0_outputs(3604));
    outputs(1401) <= not((layer0_outputs(1936)) xor (layer0_outputs(1297)));
    outputs(1402) <= not(layer0_outputs(8226));
    outputs(1403) <= not(layer0_outputs(8529));
    outputs(1404) <= not(layer0_outputs(9640));
    outputs(1405) <= (layer0_outputs(6495)) and not (layer0_outputs(3352));
    outputs(1406) <= (layer0_outputs(6023)) and (layer0_outputs(7251));
    outputs(1407) <= (layer0_outputs(6158)) and not (layer0_outputs(5778));
    outputs(1408) <= not(layer0_outputs(9703));
    outputs(1409) <= not(layer0_outputs(5967));
    outputs(1410) <= not((layer0_outputs(5222)) xor (layer0_outputs(3033)));
    outputs(1411) <= (layer0_outputs(719)) and not (layer0_outputs(10085));
    outputs(1412) <= not(layer0_outputs(5923)) or (layer0_outputs(3912));
    outputs(1413) <= (layer0_outputs(6396)) and not (layer0_outputs(4430));
    outputs(1414) <= not((layer0_outputs(7929)) or (layer0_outputs(2620)));
    outputs(1415) <= (layer0_outputs(6918)) and (layer0_outputs(3122));
    outputs(1416) <= (layer0_outputs(4059)) and (layer0_outputs(904));
    outputs(1417) <= not((layer0_outputs(1347)) or (layer0_outputs(2989)));
    outputs(1418) <= (layer0_outputs(8438)) and not (layer0_outputs(8890));
    outputs(1419) <= not((layer0_outputs(3816)) or (layer0_outputs(8920)));
    outputs(1420) <= not((layer0_outputs(8687)) or (layer0_outputs(4735)));
    outputs(1421) <= not((layer0_outputs(8352)) or (layer0_outputs(1040)));
    outputs(1422) <= (layer0_outputs(45)) and not (layer0_outputs(4101));
    outputs(1423) <= (layer0_outputs(2865)) and (layer0_outputs(4114));
    outputs(1424) <= not((layer0_outputs(5509)) xor (layer0_outputs(71)));
    outputs(1425) <= (layer0_outputs(4971)) and (layer0_outputs(7931));
    outputs(1426) <= not((layer0_outputs(9334)) xor (layer0_outputs(312)));
    outputs(1427) <= not(layer0_outputs(8892));
    outputs(1428) <= not((layer0_outputs(3771)) xor (layer0_outputs(6943)));
    outputs(1429) <= not((layer0_outputs(9951)) or (layer0_outputs(5937)));
    outputs(1430) <= (layer0_outputs(8318)) xor (layer0_outputs(5482));
    outputs(1431) <= not(layer0_outputs(8552));
    outputs(1432) <= (layer0_outputs(8747)) and (layer0_outputs(8945));
    outputs(1433) <= layer0_outputs(6803);
    outputs(1434) <= not((layer0_outputs(403)) or (layer0_outputs(2227)));
    outputs(1435) <= (layer0_outputs(5517)) xor (layer0_outputs(5237));
    outputs(1436) <= (layer0_outputs(3809)) xor (layer0_outputs(6382));
    outputs(1437) <= (layer0_outputs(2612)) and not (layer0_outputs(6260));
    outputs(1438) <= (layer0_outputs(1133)) and not (layer0_outputs(7087));
    outputs(1439) <= not((layer0_outputs(4960)) or (layer0_outputs(2260)));
    outputs(1440) <= (layer0_outputs(4180)) and not (layer0_outputs(2559));
    outputs(1441) <= (layer0_outputs(7025)) xor (layer0_outputs(4560));
    outputs(1442) <= (layer0_outputs(3458)) and (layer0_outputs(4963));
    outputs(1443) <= layer0_outputs(3103);
    outputs(1444) <= not((layer0_outputs(2985)) xor (layer0_outputs(8601)));
    outputs(1445) <= (layer0_outputs(4330)) and not (layer0_outputs(6993));
    outputs(1446) <= (layer0_outputs(3575)) and (layer0_outputs(4707));
    outputs(1447) <= layer0_outputs(4078);
    outputs(1448) <= (layer0_outputs(2766)) and not (layer0_outputs(2265));
    outputs(1449) <= (layer0_outputs(9585)) and not (layer0_outputs(5585));
    outputs(1450) <= not((layer0_outputs(7917)) xor (layer0_outputs(95)));
    outputs(1451) <= layer0_outputs(8221);
    outputs(1452) <= layer0_outputs(8832);
    outputs(1453) <= layer0_outputs(4243);
    outputs(1454) <= not(layer0_outputs(7494));
    outputs(1455) <= (layer0_outputs(1098)) and (layer0_outputs(174));
    outputs(1456) <= '0';
    outputs(1457) <= (layer0_outputs(1083)) and not (layer0_outputs(794));
    outputs(1458) <= not(layer0_outputs(10012));
    outputs(1459) <= (layer0_outputs(8029)) and not (layer0_outputs(4673));
    outputs(1460) <= (layer0_outputs(1011)) and (layer0_outputs(2380));
    outputs(1461) <= '0';
    outputs(1462) <= (layer0_outputs(7932)) and not (layer0_outputs(9002));
    outputs(1463) <= not(layer0_outputs(5096));
    outputs(1464) <= not((layer0_outputs(7679)) or (layer0_outputs(9650)));
    outputs(1465) <= (layer0_outputs(9031)) and not (layer0_outputs(1478));
    outputs(1466) <= (layer0_outputs(9343)) and not (layer0_outputs(7689));
    outputs(1467) <= not((layer0_outputs(9450)) xor (layer0_outputs(5634)));
    outputs(1468) <= (layer0_outputs(3567)) and not (layer0_outputs(3971));
    outputs(1469) <= not((layer0_outputs(3954)) xor (layer0_outputs(3346)));
    outputs(1470) <= (layer0_outputs(1611)) and (layer0_outputs(354));
    outputs(1471) <= (layer0_outputs(7558)) and (layer0_outputs(4046));
    outputs(1472) <= layer0_outputs(3988);
    outputs(1473) <= not((layer0_outputs(848)) or (layer0_outputs(9134)));
    outputs(1474) <= (layer0_outputs(1903)) xor (layer0_outputs(3650));
    outputs(1475) <= (layer0_outputs(5273)) and (layer0_outputs(5517));
    outputs(1476) <= not((layer0_outputs(7667)) xor (layer0_outputs(8407)));
    outputs(1477) <= (layer0_outputs(1800)) and not (layer0_outputs(3315));
    outputs(1478) <= not(layer0_outputs(9387));
    outputs(1479) <= not((layer0_outputs(2616)) or (layer0_outputs(3670)));
    outputs(1480) <= (layer0_outputs(1651)) and not (layer0_outputs(5621));
    outputs(1481) <= layer0_outputs(7578);
    outputs(1482) <= not((layer0_outputs(10139)) or (layer0_outputs(579)));
    outputs(1483) <= layer0_outputs(6262);
    outputs(1484) <= layer0_outputs(4969);
    outputs(1485) <= not(layer0_outputs(1582));
    outputs(1486) <= not((layer0_outputs(5234)) or (layer0_outputs(6807)));
    outputs(1487) <= (layer0_outputs(456)) and (layer0_outputs(3101));
    outputs(1488) <= (layer0_outputs(6922)) and not (layer0_outputs(4380));
    outputs(1489) <= (layer0_outputs(1818)) and not (layer0_outputs(9544));
    outputs(1490) <= layer0_outputs(7992);
    outputs(1491) <= (layer0_outputs(1178)) xor (layer0_outputs(9337));
    outputs(1492) <= not((layer0_outputs(6778)) xor (layer0_outputs(3960)));
    outputs(1493) <= (layer0_outputs(5029)) and not (layer0_outputs(721));
    outputs(1494) <= (layer0_outputs(6005)) and not (layer0_outputs(2968));
    outputs(1495) <= not((layer0_outputs(10010)) or (layer0_outputs(7476)));
    outputs(1496) <= not(layer0_outputs(559));
    outputs(1497) <= not((layer0_outputs(5882)) or (layer0_outputs(6353)));
    outputs(1498) <= layer0_outputs(4317);
    outputs(1499) <= layer0_outputs(7078);
    outputs(1500) <= (layer0_outputs(1151)) and (layer0_outputs(3931));
    outputs(1501) <= layer0_outputs(2008);
    outputs(1502) <= not((layer0_outputs(10233)) xor (layer0_outputs(2161)));
    outputs(1503) <= layer0_outputs(9878);
    outputs(1504) <= (layer0_outputs(6367)) and (layer0_outputs(7559));
    outputs(1505) <= (layer0_outputs(2644)) and not (layer0_outputs(6845));
    outputs(1506) <= (layer0_outputs(8612)) and not (layer0_outputs(7716));
    outputs(1507) <= (layer0_outputs(7900)) and not (layer0_outputs(2344));
    outputs(1508) <= (layer0_outputs(2276)) and not (layer0_outputs(2829));
    outputs(1509) <= not((layer0_outputs(8657)) or (layer0_outputs(7075)));
    outputs(1510) <= (layer0_outputs(4115)) and (layer0_outputs(2748));
    outputs(1511) <= not((layer0_outputs(4721)) xor (layer0_outputs(4051)));
    outputs(1512) <= not(layer0_outputs(5417));
    outputs(1513) <= (layer0_outputs(5140)) and (layer0_outputs(2912));
    outputs(1514) <= (layer0_outputs(3858)) or (layer0_outputs(5004));
    outputs(1515) <= not((layer0_outputs(5919)) or (layer0_outputs(43)));
    outputs(1516) <= (layer0_outputs(1808)) xor (layer0_outputs(2681));
    outputs(1517) <= (layer0_outputs(309)) xor (layer0_outputs(10231));
    outputs(1518) <= not(layer0_outputs(9461));
    outputs(1519) <= (layer0_outputs(8315)) xor (layer0_outputs(3398));
    outputs(1520) <= (layer0_outputs(5947)) and not (layer0_outputs(1095));
    outputs(1521) <= layer0_outputs(6361);
    outputs(1522) <= not((layer0_outputs(3810)) xor (layer0_outputs(9981)));
    outputs(1523) <= (layer0_outputs(5863)) and not (layer0_outputs(1993));
    outputs(1524) <= not((layer0_outputs(8353)) xor (layer0_outputs(3605)));
    outputs(1525) <= (layer0_outputs(1879)) and not (layer0_outputs(8095));
    outputs(1526) <= (layer0_outputs(5383)) and (layer0_outputs(4390));
    outputs(1527) <= not((layer0_outputs(4919)) xor (layer0_outputs(8988)));
    outputs(1528) <= not(layer0_outputs(8139));
    outputs(1529) <= not(layer0_outputs(5885));
    outputs(1530) <= not(layer0_outputs(8890));
    outputs(1531) <= layer0_outputs(5104);
    outputs(1532) <= not((layer0_outputs(1870)) xor (layer0_outputs(4033)));
    outputs(1533) <= (layer0_outputs(8527)) and not (layer0_outputs(3262));
    outputs(1534) <= not((layer0_outputs(8779)) or (layer0_outputs(9307)));
    outputs(1535) <= not((layer0_outputs(4380)) xor (layer0_outputs(965)));
    outputs(1536) <= (layer0_outputs(6060)) and (layer0_outputs(3614));
    outputs(1537) <= not(layer0_outputs(7295));
    outputs(1538) <= not((layer0_outputs(4206)) or (layer0_outputs(5476)));
    outputs(1539) <= (layer0_outputs(1674)) and not (layer0_outputs(4294));
    outputs(1540) <= (layer0_outputs(5365)) xor (layer0_outputs(2677));
    outputs(1541) <= (layer0_outputs(8142)) xor (layer0_outputs(9150));
    outputs(1542) <= (layer0_outputs(5588)) and not (layer0_outputs(8157));
    outputs(1543) <= (layer0_outputs(5710)) and not (layer0_outputs(6777));
    outputs(1544) <= not((layer0_outputs(2801)) xor (layer0_outputs(7952)));
    outputs(1545) <= (layer0_outputs(1944)) and (layer0_outputs(4250));
    outputs(1546) <= (layer0_outputs(6940)) xor (layer0_outputs(3265));
    outputs(1547) <= layer0_outputs(8522);
    outputs(1548) <= not((layer0_outputs(724)) xor (layer0_outputs(688)));
    outputs(1549) <= not((layer0_outputs(10195)) or (layer0_outputs(5836)));
    outputs(1550) <= (layer0_outputs(241)) and (layer0_outputs(468));
    outputs(1551) <= not(layer0_outputs(3520));
    outputs(1552) <= (layer0_outputs(7122)) and not (layer0_outputs(2895));
    outputs(1553) <= not(layer0_outputs(707));
    outputs(1554) <= (layer0_outputs(6199)) xor (layer0_outputs(676));
    outputs(1555) <= layer0_outputs(4914);
    outputs(1556) <= layer0_outputs(3151);
    outputs(1557) <= (layer0_outputs(7902)) and not (layer0_outputs(4731));
    outputs(1558) <= (layer0_outputs(9661)) and not (layer0_outputs(9765));
    outputs(1559) <= (layer0_outputs(264)) and not (layer0_outputs(2989));
    outputs(1560) <= not((layer0_outputs(3519)) or (layer0_outputs(9788)));
    outputs(1561) <= (layer0_outputs(1022)) and not (layer0_outputs(2409));
    outputs(1562) <= not(layer0_outputs(9325));
    outputs(1563) <= (layer0_outputs(4629)) and not (layer0_outputs(7076));
    outputs(1564) <= (layer0_outputs(7097)) xor (layer0_outputs(5692));
    outputs(1565) <= layer0_outputs(7799);
    outputs(1566) <= not((layer0_outputs(6731)) xor (layer0_outputs(4178)));
    outputs(1567) <= (layer0_outputs(8784)) and not (layer0_outputs(4931));
    outputs(1568) <= not((layer0_outputs(9975)) or (layer0_outputs(1407)));
    outputs(1569) <= (layer0_outputs(4056)) and not (layer0_outputs(3341));
    outputs(1570) <= (layer0_outputs(7935)) xor (layer0_outputs(170));
    outputs(1571) <= (layer0_outputs(7187)) and not (layer0_outputs(3266));
    outputs(1572) <= (layer0_outputs(6089)) and (layer0_outputs(4243));
    outputs(1573) <= (layer0_outputs(6743)) or (layer0_outputs(9182));
    outputs(1574) <= not((layer0_outputs(5799)) or (layer0_outputs(4805)));
    outputs(1575) <= (layer0_outputs(945)) and not (layer0_outputs(4679));
    outputs(1576) <= (layer0_outputs(8223)) and not (layer0_outputs(2570));
    outputs(1577) <= (layer0_outputs(8822)) xor (layer0_outputs(3771));
    outputs(1578) <= (layer0_outputs(105)) and (layer0_outputs(9482));
    outputs(1579) <= not(layer0_outputs(9566));
    outputs(1580) <= layer0_outputs(1797);
    outputs(1581) <= (layer0_outputs(5786)) and (layer0_outputs(1529));
    outputs(1582) <= layer0_outputs(9942);
    outputs(1583) <= (layer0_outputs(7818)) and (layer0_outputs(10221));
    outputs(1584) <= not(layer0_outputs(5460));
    outputs(1585) <= not((layer0_outputs(4060)) xor (layer0_outputs(7383)));
    outputs(1586) <= (layer0_outputs(7651)) and not (layer0_outputs(8790));
    outputs(1587) <= (layer0_outputs(5614)) and (layer0_outputs(1659));
    outputs(1588) <= (layer0_outputs(4288)) and not (layer0_outputs(9077));
    outputs(1589) <= (layer0_outputs(959)) and (layer0_outputs(7997));
    outputs(1590) <= not(layer0_outputs(1224));
    outputs(1591) <= layer0_outputs(6690);
    outputs(1592) <= (layer0_outputs(3728)) and not (layer0_outputs(7632));
    outputs(1593) <= (layer0_outputs(6092)) and not (layer0_outputs(9082));
    outputs(1594) <= (layer0_outputs(8155)) and not (layer0_outputs(1064));
    outputs(1595) <= (layer0_outputs(5223)) xor (layer0_outputs(7093));
    outputs(1596) <= '0';
    outputs(1597) <= (layer0_outputs(3660)) and not (layer0_outputs(5387));
    outputs(1598) <= (layer0_outputs(1692)) and (layer0_outputs(9921));
    outputs(1599) <= not((layer0_outputs(8454)) or (layer0_outputs(7097)));
    outputs(1600) <= (layer0_outputs(8021)) and not (layer0_outputs(7986));
    outputs(1601) <= layer0_outputs(4728);
    outputs(1602) <= not((layer0_outputs(3355)) or (layer0_outputs(8729)));
    outputs(1603) <= (layer0_outputs(8949)) and (layer0_outputs(2639));
    outputs(1604) <= not((layer0_outputs(8640)) or (layer0_outputs(1429)));
    outputs(1605) <= (layer0_outputs(8965)) and (layer0_outputs(8501));
    outputs(1606) <= not((layer0_outputs(6181)) or (layer0_outputs(9168)));
    outputs(1607) <= (layer0_outputs(9573)) and not (layer0_outputs(5798));
    outputs(1608) <= '0';
    outputs(1609) <= not((layer0_outputs(4660)) or (layer0_outputs(3503)));
    outputs(1610) <= (layer0_outputs(1917)) and not (layer0_outputs(73));
    outputs(1611) <= layer0_outputs(8148);
    outputs(1612) <= (layer0_outputs(1276)) and not (layer0_outputs(9999));
    outputs(1613) <= (layer0_outputs(3893)) and not (layer0_outputs(9091));
    outputs(1614) <= not((layer0_outputs(10087)) or (layer0_outputs(4995)));
    outputs(1615) <= not((layer0_outputs(7709)) xor (layer0_outputs(6227)));
    outputs(1616) <= layer0_outputs(7974);
    outputs(1617) <= (layer0_outputs(6163)) xor (layer0_outputs(4678));
    outputs(1618) <= (layer0_outputs(8638)) and not (layer0_outputs(8752));
    outputs(1619) <= (layer0_outputs(6375)) xor (layer0_outputs(35));
    outputs(1620) <= (layer0_outputs(6574)) and not (layer0_outputs(3501));
    outputs(1621) <= (layer0_outputs(2705)) and not (layer0_outputs(1240));
    outputs(1622) <= (layer0_outputs(8875)) xor (layer0_outputs(172));
    outputs(1623) <= (layer0_outputs(165)) xor (layer0_outputs(10042));
    outputs(1624) <= not(layer0_outputs(4912));
    outputs(1625) <= not(layer0_outputs(1694));
    outputs(1626) <= (layer0_outputs(1010)) and (layer0_outputs(8580));
    outputs(1627) <= not((layer0_outputs(1691)) xor (layer0_outputs(9695)));
    outputs(1628) <= (layer0_outputs(8042)) xor (layer0_outputs(4194));
    outputs(1629) <= (layer0_outputs(10156)) and not (layer0_outputs(2781));
    outputs(1630) <= layer0_outputs(8378);
    outputs(1631) <= (layer0_outputs(3490)) and (layer0_outputs(1795));
    outputs(1632) <= (layer0_outputs(4254)) and (layer0_outputs(3589));
    outputs(1633) <= not(layer0_outputs(6701));
    outputs(1634) <= '0';
    outputs(1635) <= (layer0_outputs(9963)) and not (layer0_outputs(9604));
    outputs(1636) <= (layer0_outputs(3695)) and (layer0_outputs(10189));
    outputs(1637) <= (layer0_outputs(10062)) and not (layer0_outputs(3715));
    outputs(1638) <= (layer0_outputs(3653)) and not (layer0_outputs(6130));
    outputs(1639) <= (layer0_outputs(8021)) and (layer0_outputs(1555));
    outputs(1640) <= layer0_outputs(3259);
    outputs(1641) <= (layer0_outputs(9909)) xor (layer0_outputs(5366));
    outputs(1642) <= (layer0_outputs(1981)) and not (layer0_outputs(8754));
    outputs(1643) <= not((layer0_outputs(7471)) or (layer0_outputs(8822)));
    outputs(1644) <= (layer0_outputs(9713)) and (layer0_outputs(3424));
    outputs(1645) <= layer0_outputs(9509);
    outputs(1646) <= layer0_outputs(6759);
    outputs(1647) <= (layer0_outputs(9074)) xor (layer0_outputs(6322));
    outputs(1648) <= not(layer0_outputs(69));
    outputs(1649) <= (layer0_outputs(3598)) and (layer0_outputs(8301));
    outputs(1650) <= (layer0_outputs(1385)) xor (layer0_outputs(5472));
    outputs(1651) <= (layer0_outputs(8047)) and not (layer0_outputs(4993));
    outputs(1652) <= (layer0_outputs(4902)) and not (layer0_outputs(5986));
    outputs(1653) <= (layer0_outputs(6981)) xor (layer0_outputs(9249));
    outputs(1654) <= not(layer0_outputs(4801));
    outputs(1655) <= not((layer0_outputs(992)) and (layer0_outputs(2088)));
    outputs(1656) <= (layer0_outputs(3710)) and not (layer0_outputs(8256));
    outputs(1657) <= (layer0_outputs(2041)) and (layer0_outputs(5857));
    outputs(1658) <= layer0_outputs(9266);
    outputs(1659) <= not((layer0_outputs(781)) xor (layer0_outputs(1343)));
    outputs(1660) <= not((layer0_outputs(4549)) or (layer0_outputs(2832)));
    outputs(1661) <= not((layer0_outputs(1101)) or (layer0_outputs(2038)));
    outputs(1662) <= not((layer0_outputs(5895)) xor (layer0_outputs(8771)));
    outputs(1663) <= not((layer0_outputs(10089)) xor (layer0_outputs(30)));
    outputs(1664) <= (layer0_outputs(10219)) and (layer0_outputs(2308));
    outputs(1665) <= not(layer0_outputs(4474));
    outputs(1666) <= layer0_outputs(2326);
    outputs(1667) <= (layer0_outputs(7521)) xor (layer0_outputs(863));
    outputs(1668) <= (layer0_outputs(198)) and not (layer0_outputs(2248));
    outputs(1669) <= (layer0_outputs(1952)) and not (layer0_outputs(1486));
    outputs(1670) <= not(layer0_outputs(8212)) or (layer0_outputs(3931));
    outputs(1671) <= (layer0_outputs(6688)) and (layer0_outputs(10038));
    outputs(1672) <= (layer0_outputs(2857)) and not (layer0_outputs(8855));
    outputs(1673) <= layer0_outputs(2527);
    outputs(1674) <= not((layer0_outputs(7317)) or (layer0_outputs(9114)));
    outputs(1675) <= layer0_outputs(2230);
    outputs(1676) <= not(layer0_outputs(6148)) or (layer0_outputs(6052));
    outputs(1677) <= not(layer0_outputs(5553)) or (layer0_outputs(1209));
    outputs(1678) <= not((layer0_outputs(6893)) or (layer0_outputs(8567)));
    outputs(1679) <= layer0_outputs(9322);
    outputs(1680) <= (layer0_outputs(5217)) and not (layer0_outputs(9235));
    outputs(1681) <= layer0_outputs(8759);
    outputs(1682) <= layer0_outputs(7640);
    outputs(1683) <= (layer0_outputs(5427)) xor (layer0_outputs(9038));
    outputs(1684) <= (layer0_outputs(10002)) and not (layer0_outputs(6822));
    outputs(1685) <= (layer0_outputs(2106)) and (layer0_outputs(1580));
    outputs(1686) <= not(layer0_outputs(4221));
    outputs(1687) <= (layer0_outputs(9417)) and not (layer0_outputs(7155));
    outputs(1688) <= not(layer0_outputs(4023));
    outputs(1689) <= layer0_outputs(6762);
    outputs(1690) <= layer0_outputs(4489);
    outputs(1691) <= not((layer0_outputs(4111)) or (layer0_outputs(1025)));
    outputs(1692) <= layer0_outputs(2902);
    outputs(1693) <= not(layer0_outputs(9643));
    outputs(1694) <= (layer0_outputs(1397)) and (layer0_outputs(1556));
    outputs(1695) <= not(layer0_outputs(8547));
    outputs(1696) <= (layer0_outputs(6230)) and not (layer0_outputs(249));
    outputs(1697) <= (layer0_outputs(4896)) and (layer0_outputs(9423));
    outputs(1698) <= (layer0_outputs(10034)) and (layer0_outputs(2823));
    outputs(1699) <= (layer0_outputs(2002)) and not (layer0_outputs(3330));
    outputs(1700) <= (layer0_outputs(2361)) and not (layer0_outputs(8925));
    outputs(1701) <= not((layer0_outputs(8980)) or (layer0_outputs(8962)));
    outputs(1702) <= '0';
    outputs(1703) <= (layer0_outputs(2880)) and not (layer0_outputs(5685));
    outputs(1704) <= (layer0_outputs(8966)) and not (layer0_outputs(8134));
    outputs(1705) <= (layer0_outputs(1828)) and not (layer0_outputs(5852));
    outputs(1706) <= not((layer0_outputs(8784)) xor (layer0_outputs(9505)));
    outputs(1707) <= not(layer0_outputs(814));
    outputs(1708) <= not((layer0_outputs(8607)) or (layer0_outputs(8785)));
    outputs(1709) <= not((layer0_outputs(484)) xor (layer0_outputs(6292)));
    outputs(1710) <= (layer0_outputs(4466)) and (layer0_outputs(2676));
    outputs(1711) <= (layer0_outputs(7964)) xor (layer0_outputs(1041));
    outputs(1712) <= (layer0_outputs(9458)) and not (layer0_outputs(2786));
    outputs(1713) <= not((layer0_outputs(6323)) xor (layer0_outputs(928)));
    outputs(1714) <= (layer0_outputs(375)) and not (layer0_outputs(9357));
    outputs(1715) <= (layer0_outputs(3163)) and not (layer0_outputs(6851));
    outputs(1716) <= (layer0_outputs(3080)) and not (layer0_outputs(246));
    outputs(1717) <= (layer0_outputs(7089)) and not (layer0_outputs(2322));
    outputs(1718) <= (layer0_outputs(973)) and (layer0_outputs(3541));
    outputs(1719) <= (layer0_outputs(4014)) and not (layer0_outputs(380));
    outputs(1720) <= not((layer0_outputs(9233)) or (layer0_outputs(3891)));
    outputs(1721) <= (layer0_outputs(2235)) and not (layer0_outputs(7628));
    outputs(1722) <= (layer0_outputs(8702)) and not (layer0_outputs(5378));
    outputs(1723) <= not(layer0_outputs(4241));
    outputs(1724) <= layer0_outputs(4941);
    outputs(1725) <= (layer0_outputs(4743)) and (layer0_outputs(5603));
    outputs(1726) <= (layer0_outputs(3623)) and (layer0_outputs(8));
    outputs(1727) <= layer0_outputs(2105);
    outputs(1728) <= (layer0_outputs(7386)) and (layer0_outputs(1044));
    outputs(1729) <= (layer0_outputs(963)) and not (layer0_outputs(6797));
    outputs(1730) <= not(layer0_outputs(1372));
    outputs(1731) <= not(layer0_outputs(2203));
    outputs(1732) <= not((layer0_outputs(2940)) xor (layer0_outputs(9437)));
    outputs(1733) <= not((layer0_outputs(9085)) xor (layer0_outputs(7348)));
    outputs(1734) <= (layer0_outputs(3930)) and not (layer0_outputs(4259));
    outputs(1735) <= not(layer0_outputs(6181));
    outputs(1736) <= not((layer0_outputs(4298)) xor (layer0_outputs(1713)));
    outputs(1737) <= '0';
    outputs(1738) <= not(layer0_outputs(6916));
    outputs(1739) <= layer0_outputs(7927);
    outputs(1740) <= layer0_outputs(8483);
    outputs(1741) <= not((layer0_outputs(8164)) or (layer0_outputs(7514)));
    outputs(1742) <= (layer0_outputs(8133)) and not (layer0_outputs(9929));
    outputs(1743) <= (layer0_outputs(7369)) and not (layer0_outputs(3408));
    outputs(1744) <= not((layer0_outputs(2535)) or (layer0_outputs(1765)));
    outputs(1745) <= (layer0_outputs(139)) and (layer0_outputs(5922));
    outputs(1746) <= not((layer0_outputs(6782)) or (layer0_outputs(1450)));
    outputs(1747) <= (layer0_outputs(8378)) and (layer0_outputs(9629));
    outputs(1748) <= (layer0_outputs(2990)) and (layer0_outputs(8414));
    outputs(1749) <= (layer0_outputs(4255)) and not (layer0_outputs(1908));
    outputs(1750) <= not((layer0_outputs(8159)) or (layer0_outputs(4358)));
    outputs(1751) <= not(layer0_outputs(4310));
    outputs(1752) <= not(layer0_outputs(4090));
    outputs(1753) <= (layer0_outputs(3884)) and not (layer0_outputs(1503));
    outputs(1754) <= not(layer0_outputs(5606));
    outputs(1755) <= (layer0_outputs(3609)) xor (layer0_outputs(7317));
    outputs(1756) <= not(layer0_outputs(1216));
    outputs(1757) <= (layer0_outputs(1092)) and not (layer0_outputs(7667));
    outputs(1758) <= (layer0_outputs(5849)) and not (layer0_outputs(5819));
    outputs(1759) <= (layer0_outputs(8777)) and not (layer0_outputs(8959));
    outputs(1760) <= layer0_outputs(8680);
    outputs(1761) <= (layer0_outputs(2549)) and (layer0_outputs(1262));
    outputs(1762) <= '0';
    outputs(1763) <= layer0_outputs(9884);
    outputs(1764) <= not((layer0_outputs(4923)) xor (layer0_outputs(1868)));
    outputs(1765) <= (layer0_outputs(8243)) and not (layer0_outputs(9792));
    outputs(1766) <= not((layer0_outputs(9577)) or (layer0_outputs(6279)));
    outputs(1767) <= (layer0_outputs(3186)) and not (layer0_outputs(7357));
    outputs(1768) <= (layer0_outputs(5872)) and (layer0_outputs(3439));
    outputs(1769) <= (layer0_outputs(81)) and not (layer0_outputs(3000));
    outputs(1770) <= (layer0_outputs(9435)) and not (layer0_outputs(7798));
    outputs(1771) <= (layer0_outputs(4957)) and not (layer0_outputs(9684));
    outputs(1772) <= layer0_outputs(8645);
    outputs(1773) <= (layer0_outputs(8675)) xor (layer0_outputs(7436));
    outputs(1774) <= (layer0_outputs(2179)) and (layer0_outputs(8807));
    outputs(1775) <= (layer0_outputs(2901)) xor (layer0_outputs(5099));
    outputs(1776) <= (layer0_outputs(9463)) and (layer0_outputs(10080));
    outputs(1777) <= not((layer0_outputs(2846)) or (layer0_outputs(7501)));
    outputs(1778) <= (layer0_outputs(8018)) xor (layer0_outputs(2156));
    outputs(1779) <= (layer0_outputs(4828)) and (layer0_outputs(3256));
    outputs(1780) <= layer0_outputs(1699);
    outputs(1781) <= (layer0_outputs(5570)) and (layer0_outputs(9587));
    outputs(1782) <= (layer0_outputs(7712)) and not (layer0_outputs(3248));
    outputs(1783) <= (layer0_outputs(5076)) and not (layer0_outputs(7759));
    outputs(1784) <= not((layer0_outputs(4459)) xor (layer0_outputs(8048)));
    outputs(1785) <= (layer0_outputs(9686)) and not (layer0_outputs(2718));
    outputs(1786) <= not((layer0_outputs(4067)) or (layer0_outputs(5091)));
    outputs(1787) <= not((layer0_outputs(5833)) or (layer0_outputs(3178)));
    outputs(1788) <= (layer0_outputs(233)) and not (layer0_outputs(6450));
    outputs(1789) <= (layer0_outputs(6945)) and not (layer0_outputs(1809));
    outputs(1790) <= not((layer0_outputs(6430)) or (layer0_outputs(699)));
    outputs(1791) <= (layer0_outputs(7707)) and (layer0_outputs(6314));
    outputs(1792) <= (layer0_outputs(4063)) and (layer0_outputs(9103));
    outputs(1793) <= (layer0_outputs(6936)) and (layer0_outputs(9250));
    outputs(1794) <= (layer0_outputs(3499)) and not (layer0_outputs(6316));
    outputs(1795) <= (layer0_outputs(10217)) and not (layer0_outputs(976));
    outputs(1796) <= (layer0_outputs(7075)) xor (layer0_outputs(2220));
    outputs(1797) <= (layer0_outputs(5909)) and not (layer0_outputs(4355));
    outputs(1798) <= layer0_outputs(9935);
    outputs(1799) <= (layer0_outputs(74)) and not (layer0_outputs(4279));
    outputs(1800) <= not((layer0_outputs(8599)) or (layer0_outputs(7007)));
    outputs(1801) <= not((layer0_outputs(465)) or (layer0_outputs(6640)));
    outputs(1802) <= not((layer0_outputs(8613)) or (layer0_outputs(4297)));
    outputs(1803) <= not((layer0_outputs(8690)) or (layer0_outputs(3254)));
    outputs(1804) <= not((layer0_outputs(5036)) xor (layer0_outputs(3109)));
    outputs(1805) <= (layer0_outputs(9003)) and not (layer0_outputs(2788));
    outputs(1806) <= (layer0_outputs(1345)) xor (layer0_outputs(1908));
    outputs(1807) <= (layer0_outputs(2552)) and not (layer0_outputs(215));
    outputs(1808) <= not(layer0_outputs(1380));
    outputs(1809) <= not((layer0_outputs(3315)) or (layer0_outputs(2808)));
    outputs(1810) <= layer0_outputs(6210);
    outputs(1811) <= (layer0_outputs(387)) and not (layer0_outputs(8700));
    outputs(1812) <= not((layer0_outputs(7383)) or (layer0_outputs(8441)));
    outputs(1813) <= (layer0_outputs(5428)) and not (layer0_outputs(8256));
    outputs(1814) <= (layer0_outputs(7217)) and not (layer0_outputs(5859));
    outputs(1815) <= (layer0_outputs(741)) and not (layer0_outputs(8231));
    outputs(1816) <= not((layer0_outputs(1018)) or (layer0_outputs(3028)));
    outputs(1817) <= (layer0_outputs(9783)) and not (layer0_outputs(4257));
    outputs(1818) <= not(layer0_outputs(7112));
    outputs(1819) <= (layer0_outputs(3373)) and not (layer0_outputs(6474));
    outputs(1820) <= not((layer0_outputs(7808)) or (layer0_outputs(6044)));
    outputs(1821) <= not(layer0_outputs(3));
    outputs(1822) <= not(layer0_outputs(791));
    outputs(1823) <= layer0_outputs(9424);
    outputs(1824) <= not((layer0_outputs(3645)) or (layer0_outputs(5977)));
    outputs(1825) <= (layer0_outputs(417)) and not (layer0_outputs(7970));
    outputs(1826) <= not((layer0_outputs(1403)) xor (layer0_outputs(908)));
    outputs(1827) <= not(layer0_outputs(8635)) or (layer0_outputs(7737));
    outputs(1828) <= not((layer0_outputs(9995)) or (layer0_outputs(1794)));
    outputs(1829) <= layer0_outputs(9083);
    outputs(1830) <= not((layer0_outputs(7104)) or (layer0_outputs(7811)));
    outputs(1831) <= (layer0_outputs(3728)) and (layer0_outputs(2059));
    outputs(1832) <= not(layer0_outputs(7652));
    outputs(1833) <= '0';
    outputs(1834) <= layer0_outputs(587);
    outputs(1835) <= (layer0_outputs(6278)) xor (layer0_outputs(7211));
    outputs(1836) <= (layer0_outputs(5197)) and (layer0_outputs(6065));
    outputs(1837) <= not((layer0_outputs(1198)) or (layer0_outputs(2411)));
    outputs(1838) <= layer0_outputs(4710);
    outputs(1839) <= layer0_outputs(630);
    outputs(1840) <= not((layer0_outputs(6119)) xor (layer0_outputs(5230)));
    outputs(1841) <= (layer0_outputs(8710)) and not (layer0_outputs(2294));
    outputs(1842) <= (layer0_outputs(3637)) xor (layer0_outputs(10173));
    outputs(1843) <= (layer0_outputs(2859)) and not (layer0_outputs(3016));
    outputs(1844) <= not((layer0_outputs(803)) or (layer0_outputs(3648)));
    outputs(1845) <= not(layer0_outputs(9084));
    outputs(1846) <= (layer0_outputs(8278)) and not (layer0_outputs(7585));
    outputs(1847) <= (layer0_outputs(307)) and (layer0_outputs(6138));
    outputs(1848) <= (layer0_outputs(5225)) and not (layer0_outputs(5623));
    outputs(1849) <= (layer0_outputs(3375)) and not (layer0_outputs(5240));
    outputs(1850) <= (layer0_outputs(7747)) and not (layer0_outputs(5807));
    outputs(1851) <= (layer0_outputs(5796)) and not (layer0_outputs(5736));
    outputs(1852) <= not((layer0_outputs(2755)) or (layer0_outputs(2070)));
    outputs(1853) <= not((layer0_outputs(5669)) and (layer0_outputs(7981)));
    outputs(1854) <= (layer0_outputs(3206)) and (layer0_outputs(1132));
    outputs(1855) <= not((layer0_outputs(9213)) or (layer0_outputs(3822)));
    outputs(1856) <= '0';
    outputs(1857) <= not((layer0_outputs(6182)) or (layer0_outputs(6754)));
    outputs(1858) <= (layer0_outputs(86)) and not (layer0_outputs(8958));
    outputs(1859) <= (layer0_outputs(8002)) and not (layer0_outputs(1511));
    outputs(1860) <= (layer0_outputs(3008)) and not (layer0_outputs(1760));
    outputs(1861) <= (layer0_outputs(6271)) xor (layer0_outputs(5123));
    outputs(1862) <= not((layer0_outputs(3612)) or (layer0_outputs(9923)));
    outputs(1863) <= (layer0_outputs(9934)) and (layer0_outputs(8939));
    outputs(1864) <= (layer0_outputs(974)) xor (layer0_outputs(6197));
    outputs(1865) <= layer0_outputs(5039);
    outputs(1866) <= not((layer0_outputs(657)) xor (layer0_outputs(4909)));
    outputs(1867) <= not((layer0_outputs(9478)) or (layer0_outputs(4780)));
    outputs(1868) <= (layer0_outputs(7789)) and not (layer0_outputs(9255));
    outputs(1869) <= (layer0_outputs(3702)) xor (layer0_outputs(6239));
    outputs(1870) <= (layer0_outputs(400)) and (layer0_outputs(5314));
    outputs(1871) <= (layer0_outputs(4172)) and not (layer0_outputs(696));
    outputs(1872) <= layer0_outputs(5157);
    outputs(1873) <= not((layer0_outputs(6082)) xor (layer0_outputs(3314)));
    outputs(1874) <= not(layer0_outputs(806));
    outputs(1875) <= not((layer0_outputs(8499)) or (layer0_outputs(4695)));
    outputs(1876) <= (layer0_outputs(8732)) and not (layer0_outputs(1307));
    outputs(1877) <= not(layer0_outputs(3524)) or (layer0_outputs(4708));
    outputs(1878) <= (layer0_outputs(328)) xor (layer0_outputs(8410));
    outputs(1879) <= not((layer0_outputs(6388)) or (layer0_outputs(3782)));
    outputs(1880) <= (layer0_outputs(4329)) and (layer0_outputs(23));
    outputs(1881) <= (layer0_outputs(864)) and not (layer0_outputs(871));
    outputs(1882) <= not((layer0_outputs(3671)) or (layer0_outputs(642)));
    outputs(1883) <= (layer0_outputs(712)) and not (layer0_outputs(3226));
    outputs(1884) <= (layer0_outputs(4359)) and (layer0_outputs(4971));
    outputs(1885) <= (layer0_outputs(9599)) and not (layer0_outputs(9835));
    outputs(1886) <= (layer0_outputs(8299)) xor (layer0_outputs(7658));
    outputs(1887) <= not((layer0_outputs(6262)) xor (layer0_outputs(3091)));
    outputs(1888) <= (layer0_outputs(1185)) and (layer0_outputs(4852));
    outputs(1889) <= not((layer0_outputs(1252)) or (layer0_outputs(2523)));
    outputs(1890) <= not(layer0_outputs(6793));
    outputs(1891) <= not((layer0_outputs(9366)) or (layer0_outputs(6599)));
    outputs(1892) <= not((layer0_outputs(1774)) or (layer0_outputs(8539)));
    outputs(1893) <= (layer0_outputs(7826)) and (layer0_outputs(5918));
    outputs(1894) <= layer0_outputs(7335);
    outputs(1895) <= not((layer0_outputs(9725)) xor (layer0_outputs(700)));
    outputs(1896) <= (layer0_outputs(7245)) and not (layer0_outputs(2257));
    outputs(1897) <= (layer0_outputs(18)) and not (layer0_outputs(4953));
    outputs(1898) <= not(layer0_outputs(2174));
    outputs(1899) <= not(layer0_outputs(5960));
    outputs(1900) <= (layer0_outputs(5079)) and (layer0_outputs(7944));
    outputs(1901) <= not((layer0_outputs(6369)) or (layer0_outputs(6490)));
    outputs(1902) <= not(layer0_outputs(3885));
    outputs(1903) <= (layer0_outputs(7758)) and not (layer0_outputs(7416));
    outputs(1904) <= not(layer0_outputs(569)) or (layer0_outputs(7109));
    outputs(1905) <= (layer0_outputs(4498)) and not (layer0_outputs(9139));
    outputs(1906) <= not((layer0_outputs(1393)) or (layer0_outputs(7589)));
    outputs(1907) <= not((layer0_outputs(8392)) or (layer0_outputs(1109)));
    outputs(1908) <= not(layer0_outputs(6891));
    outputs(1909) <= not((layer0_outputs(1779)) or (layer0_outputs(9736)));
    outputs(1910) <= (layer0_outputs(441)) and not (layer0_outputs(486));
    outputs(1911) <= not((layer0_outputs(562)) or (layer0_outputs(2575)));
    outputs(1912) <= not((layer0_outputs(5948)) xor (layer0_outputs(206)));
    outputs(1913) <= (layer0_outputs(6408)) and (layer0_outputs(5022));
    outputs(1914) <= (layer0_outputs(3084)) and not (layer0_outputs(6297));
    outputs(1915) <= not(layer0_outputs(2723));
    outputs(1916) <= not((layer0_outputs(21)) or (layer0_outputs(8823)));
    outputs(1917) <= (layer0_outputs(7413)) and not (layer0_outputs(8957));
    outputs(1918) <= not((layer0_outputs(1079)) or (layer0_outputs(7289)));
    outputs(1919) <= (layer0_outputs(4722)) and (layer0_outputs(9160));
    outputs(1920) <= (layer0_outputs(9803)) and not (layer0_outputs(4031));
    outputs(1921) <= (layer0_outputs(2655)) and not (layer0_outputs(4125));
    outputs(1922) <= layer0_outputs(5056);
    outputs(1923) <= (layer0_outputs(6740)) and not (layer0_outputs(9134));
    outputs(1924) <= (layer0_outputs(5637)) and (layer0_outputs(5144));
    outputs(1925) <= layer0_outputs(6510);
    outputs(1926) <= not((layer0_outputs(9279)) and (layer0_outputs(470)));
    outputs(1927) <= (layer0_outputs(4782)) xor (layer0_outputs(9447));
    outputs(1928) <= not((layer0_outputs(3255)) xor (layer0_outputs(4138)));
    outputs(1929) <= (layer0_outputs(4235)) and (layer0_outputs(6063));
    outputs(1930) <= not((layer0_outputs(951)) xor (layer0_outputs(1901)));
    outputs(1931) <= not((layer0_outputs(426)) or (layer0_outputs(1258)));
    outputs(1932) <= (layer0_outputs(8155)) and not (layer0_outputs(3191));
    outputs(1933) <= layer0_outputs(6348);
    outputs(1934) <= not(layer0_outputs(5858));
    outputs(1935) <= (layer0_outputs(7298)) and (layer0_outputs(2416));
    outputs(1936) <= (layer0_outputs(6638)) and (layer0_outputs(1609));
    outputs(1937) <= (layer0_outputs(8302)) and not (layer0_outputs(4752));
    outputs(1938) <= not((layer0_outputs(5410)) or (layer0_outputs(8447)));
    outputs(1939) <= (layer0_outputs(5777)) and (layer0_outputs(299));
    outputs(1940) <= (layer0_outputs(1850)) xor (layer0_outputs(9177));
    outputs(1941) <= layer0_outputs(6636);
    outputs(1942) <= (layer0_outputs(2998)) and not (layer0_outputs(940));
    outputs(1943) <= (layer0_outputs(2852)) and (layer0_outputs(5677));
    outputs(1944) <= not((layer0_outputs(1170)) xor (layer0_outputs(2)));
    outputs(1945) <= (layer0_outputs(760)) and not (layer0_outputs(655));
    outputs(1946) <= (layer0_outputs(9625)) and (layer0_outputs(6588));
    outputs(1947) <= (layer0_outputs(1570)) and (layer0_outputs(1044));
    outputs(1948) <= not(layer0_outputs(50));
    outputs(1949) <= (layer0_outputs(1424)) and not (layer0_outputs(7870));
    outputs(1950) <= not(layer0_outputs(8760));
    outputs(1951) <= (layer0_outputs(8181)) and (layer0_outputs(2314));
    outputs(1952) <= (layer0_outputs(4431)) and not (layer0_outputs(4329));
    outputs(1953) <= (layer0_outputs(7401)) and not (layer0_outputs(4298));
    outputs(1954) <= (layer0_outputs(8951)) and not (layer0_outputs(191));
    outputs(1955) <= not((layer0_outputs(2422)) xor (layer0_outputs(10105)));
    outputs(1956) <= (layer0_outputs(5982)) and (layer0_outputs(5527));
    outputs(1957) <= (layer0_outputs(3221)) and (layer0_outputs(2594));
    outputs(1958) <= (layer0_outputs(1633)) and (layer0_outputs(6582));
    outputs(1959) <= (layer0_outputs(1973)) and not (layer0_outputs(9140));
    outputs(1960) <= (layer0_outputs(445)) and not (layer0_outputs(6331));
    outputs(1961) <= (layer0_outputs(853)) xor (layer0_outputs(7982));
    outputs(1962) <= not((layer0_outputs(7022)) xor (layer0_outputs(2057)));
    outputs(1963) <= not(layer0_outputs(3788));
    outputs(1964) <= layer0_outputs(2068);
    outputs(1965) <= layer0_outputs(7486);
    outputs(1966) <= (layer0_outputs(6167)) xor (layer0_outputs(9843));
    outputs(1967) <= (layer0_outputs(6960)) and (layer0_outputs(136));
    outputs(1968) <= (layer0_outputs(4864)) and not (layer0_outputs(3817));
    outputs(1969) <= not((layer0_outputs(6107)) or (layer0_outputs(2430)));
    outputs(1970) <= (layer0_outputs(9729)) and not (layer0_outputs(8830));
    outputs(1971) <= (layer0_outputs(7240)) and (layer0_outputs(8049));
    outputs(1972) <= layer0_outputs(3650);
    outputs(1973) <= (layer0_outputs(6057)) and not (layer0_outputs(4609));
    outputs(1974) <= not((layer0_outputs(1698)) or (layer0_outputs(8160)));
    outputs(1975) <= (layer0_outputs(9356)) and not (layer0_outputs(598));
    outputs(1976) <= (layer0_outputs(9211)) and not (layer0_outputs(9062));
    outputs(1977) <= (layer0_outputs(1785)) and (layer0_outputs(3604));
    outputs(1978) <= not((layer0_outputs(4791)) xor (layer0_outputs(4433)));
    outputs(1979) <= not((layer0_outputs(1530)) xor (layer0_outputs(4663)));
    outputs(1980) <= (layer0_outputs(6622)) and not (layer0_outputs(639));
    outputs(1981) <= not((layer0_outputs(9033)) xor (layer0_outputs(892)));
    outputs(1982) <= (layer0_outputs(2885)) and not (layer0_outputs(8589));
    outputs(1983) <= not((layer0_outputs(3676)) or (layer0_outputs(9425)));
    outputs(1984) <= not(layer0_outputs(10182));
    outputs(1985) <= (layer0_outputs(755)) and not (layer0_outputs(5495));
    outputs(1986) <= not((layer0_outputs(294)) xor (layer0_outputs(8309)));
    outputs(1987) <= not((layer0_outputs(5266)) or (layer0_outputs(179)));
    outputs(1988) <= '0';
    outputs(1989) <= not(layer0_outputs(3048));
    outputs(1990) <= not((layer0_outputs(4870)) or (layer0_outputs(2091)));
    outputs(1991) <= (layer0_outputs(4246)) and not (layer0_outputs(4979));
    outputs(1992) <= layer0_outputs(6198);
    outputs(1993) <= '0';
    outputs(1994) <= not((layer0_outputs(9773)) or (layer0_outputs(8531)));
    outputs(1995) <= (layer0_outputs(6069)) and not (layer0_outputs(4441));
    outputs(1996) <= (layer0_outputs(2627)) and (layer0_outputs(99));
    outputs(1997) <= not(layer0_outputs(1669));
    outputs(1998) <= not((layer0_outputs(3619)) or (layer0_outputs(4907)));
    outputs(1999) <= not(layer0_outputs(8476));
    outputs(2000) <= layer0_outputs(1781);
    outputs(2001) <= (layer0_outputs(7575)) and not (layer0_outputs(2995));
    outputs(2002) <= not((layer0_outputs(10029)) xor (layer0_outputs(521)));
    outputs(2003) <= (layer0_outputs(2127)) and (layer0_outputs(3154));
    outputs(2004) <= layer0_outputs(211);
    outputs(2005) <= (layer0_outputs(5471)) and not (layer0_outputs(10004));
    outputs(2006) <= (layer0_outputs(9708)) and not (layer0_outputs(1430));
    outputs(2007) <= not(layer0_outputs(808));
    outputs(2008) <= layer0_outputs(1528);
    outputs(2009) <= not((layer0_outputs(6531)) or (layer0_outputs(6818)));
    outputs(2010) <= '0';
    outputs(2011) <= (layer0_outputs(1481)) and not (layer0_outputs(6980));
    outputs(2012) <= '0';
    outputs(2013) <= (layer0_outputs(4851)) and not (layer0_outputs(5007));
    outputs(2014) <= (layer0_outputs(4703)) and not (layer0_outputs(1771));
    outputs(2015) <= (layer0_outputs(4826)) and not (layer0_outputs(2550));
    outputs(2016) <= not((layer0_outputs(2426)) or (layer0_outputs(8073)));
    outputs(2017) <= (layer0_outputs(9106)) and not (layer0_outputs(8050));
    outputs(2018) <= (layer0_outputs(9495)) and not (layer0_outputs(6719));
    outputs(2019) <= not((layer0_outputs(4844)) or (layer0_outputs(8863)));
    outputs(2020) <= layer0_outputs(1126);
    outputs(2021) <= (layer0_outputs(5287)) and not (layer0_outputs(8987));
    outputs(2022) <= layer0_outputs(5586);
    outputs(2023) <= (layer0_outputs(104)) and not (layer0_outputs(330));
    outputs(2024) <= not(layer0_outputs(2022));
    outputs(2025) <= (layer0_outputs(5026)) and not (layer0_outputs(7409));
    outputs(2026) <= not(layer0_outputs(6770)) or (layer0_outputs(2291));
    outputs(2027) <= (layer0_outputs(5521)) and not (layer0_outputs(5136));
    outputs(2028) <= (layer0_outputs(1299)) xor (layer0_outputs(6121));
    outputs(2029) <= not(layer0_outputs(1451));
    outputs(2030) <= layer0_outputs(998);
    outputs(2031) <= (layer0_outputs(7874)) and (layer0_outputs(897));
    outputs(2032) <= layer0_outputs(333);
    outputs(2033) <= (layer0_outputs(7812)) and not (layer0_outputs(6103));
    outputs(2034) <= (layer0_outputs(6312)) and not (layer0_outputs(4109));
    outputs(2035) <= layer0_outputs(8162);
    outputs(2036) <= (layer0_outputs(7914)) and not (layer0_outputs(5098));
    outputs(2037) <= (layer0_outputs(8370)) and not (layer0_outputs(4179));
    outputs(2038) <= not(layer0_outputs(4959)) or (layer0_outputs(4646));
    outputs(2039) <= (layer0_outputs(9015)) and (layer0_outputs(1157));
    outputs(2040) <= (layer0_outputs(3347)) and (layer0_outputs(6124));
    outputs(2041) <= (layer0_outputs(5933)) xor (layer0_outputs(8970));
    outputs(2042) <= not((layer0_outputs(5518)) or (layer0_outputs(6648)));
    outputs(2043) <= not((layer0_outputs(9436)) or (layer0_outputs(6952)));
    outputs(2044) <= (layer0_outputs(6633)) and (layer0_outputs(1411));
    outputs(2045) <= (layer0_outputs(3194)) and not (layer0_outputs(5651));
    outputs(2046) <= not(layer0_outputs(6704));
    outputs(2047) <= (layer0_outputs(8757)) xor (layer0_outputs(4073));
    outputs(2048) <= not(layer0_outputs(8502));
    outputs(2049) <= not(layer0_outputs(9561)) or (layer0_outputs(2242));
    outputs(2050) <= not(layer0_outputs(8939));
    outputs(2051) <= (layer0_outputs(5758)) or (layer0_outputs(3720));
    outputs(2052) <= not(layer0_outputs(3594));
    outputs(2053) <= not(layer0_outputs(2870)) or (layer0_outputs(6320));
    outputs(2054) <= not(layer0_outputs(9109));
    outputs(2055) <= not(layer0_outputs(6811));
    outputs(2056) <= layer0_outputs(7107);
    outputs(2057) <= (layer0_outputs(1816)) xor (layer0_outputs(9656));
    outputs(2058) <= not(layer0_outputs(1185));
    outputs(2059) <= not((layer0_outputs(1750)) xor (layer0_outputs(3885)));
    outputs(2060) <= not(layer0_outputs(1589));
    outputs(2061) <= layer0_outputs(7125);
    outputs(2062) <= layer0_outputs(638);
    outputs(2063) <= layer0_outputs(7427);
    outputs(2064) <= not(layer0_outputs(6651)) or (layer0_outputs(1129));
    outputs(2065) <= not(layer0_outputs(316)) or (layer0_outputs(4617));
    outputs(2066) <= layer0_outputs(4889);
    outputs(2067) <= not(layer0_outputs(8200));
    outputs(2068) <= (layer0_outputs(2636)) xor (layer0_outputs(9546));
    outputs(2069) <= not(layer0_outputs(8071));
    outputs(2070) <= not((layer0_outputs(4202)) or (layer0_outputs(3760)));
    outputs(2071) <= layer0_outputs(54);
    outputs(2072) <= (layer0_outputs(6595)) xor (layer0_outputs(10023));
    outputs(2073) <= (layer0_outputs(9697)) xor (layer0_outputs(6138));
    outputs(2074) <= not(layer0_outputs(6019)) or (layer0_outputs(903));
    outputs(2075) <= not((layer0_outputs(4962)) xor (layer0_outputs(8462)));
    outputs(2076) <= not(layer0_outputs(7418));
    outputs(2077) <= (layer0_outputs(6462)) xor (layer0_outputs(2557));
    outputs(2078) <= not(layer0_outputs(2125));
    outputs(2079) <= (layer0_outputs(8253)) and not (layer0_outputs(3326));
    outputs(2080) <= not((layer0_outputs(9185)) xor (layer0_outputs(5380)));
    outputs(2081) <= not((layer0_outputs(4432)) and (layer0_outputs(5674)));
    outputs(2082) <= layer0_outputs(8704);
    outputs(2083) <= not((layer0_outputs(4558)) xor (layer0_outputs(9125)));
    outputs(2084) <= not(layer0_outputs(5574));
    outputs(2085) <= not(layer0_outputs(7485));
    outputs(2086) <= (layer0_outputs(1592)) and not (layer0_outputs(7650));
    outputs(2087) <= not(layer0_outputs(21));
    outputs(2088) <= (layer0_outputs(6397)) xor (layer0_outputs(2545));
    outputs(2089) <= not((layer0_outputs(5652)) xor (layer0_outputs(2473)));
    outputs(2090) <= (layer0_outputs(4068)) or (layer0_outputs(9165));
    outputs(2091) <= not(layer0_outputs(3145));
    outputs(2092) <= (layer0_outputs(1381)) xor (layer0_outputs(9257));
    outputs(2093) <= not(layer0_outputs(1141));
    outputs(2094) <= not(layer0_outputs(2054));
    outputs(2095) <= layer0_outputs(5129);
    outputs(2096) <= not(layer0_outputs(9740));
    outputs(2097) <= not(layer0_outputs(5608)) or (layer0_outputs(4218));
    outputs(2098) <= not(layer0_outputs(1936));
    outputs(2099) <= not((layer0_outputs(4868)) or (layer0_outputs(1740)));
    outputs(2100) <= (layer0_outputs(5667)) xor (layer0_outputs(5766));
    outputs(2101) <= not(layer0_outputs(5000));
    outputs(2102) <= layer0_outputs(9150);
    outputs(2103) <= (layer0_outputs(3031)) or (layer0_outputs(7756));
    outputs(2104) <= not((layer0_outputs(2905)) xor (layer0_outputs(991)));
    outputs(2105) <= not(layer0_outputs(816));
    outputs(2106) <= layer0_outputs(9512);
    outputs(2107) <= not(layer0_outputs(8933));
    outputs(2108) <= (layer0_outputs(3041)) and (layer0_outputs(9897));
    outputs(2109) <= not(layer0_outputs(5452));
    outputs(2110) <= layer0_outputs(3045);
    outputs(2111) <= (layer0_outputs(2300)) and not (layer0_outputs(8344));
    outputs(2112) <= not((layer0_outputs(6116)) and (layer0_outputs(6361)));
    outputs(2113) <= (layer0_outputs(4535)) and not (layer0_outputs(5045));
    outputs(2114) <= not((layer0_outputs(9758)) xor (layer0_outputs(5825)));
    outputs(2115) <= not(layer0_outputs(7683));
    outputs(2116) <= layer0_outputs(5277);
    outputs(2117) <= layer0_outputs(1449);
    outputs(2118) <= not((layer0_outputs(9876)) and (layer0_outputs(1868)));
    outputs(2119) <= not(layer0_outputs(4988));
    outputs(2120) <= not(layer0_outputs(9901));
    outputs(2121) <= (layer0_outputs(276)) xor (layer0_outputs(3113));
    outputs(2122) <= not((layer0_outputs(9057)) and (layer0_outputs(8002)));
    outputs(2123) <= layer0_outputs(615);
    outputs(2124) <= not((layer0_outputs(3590)) xor (layer0_outputs(324)));
    outputs(2125) <= layer0_outputs(9407);
    outputs(2126) <= layer0_outputs(6011);
    outputs(2127) <= layer0_outputs(1066);
    outputs(2128) <= layer0_outputs(2642);
    outputs(2129) <= not((layer0_outputs(8116)) or (layer0_outputs(584)));
    outputs(2130) <= not((layer0_outputs(5194)) and (layer0_outputs(1703)));
    outputs(2131) <= not(layer0_outputs(226)) or (layer0_outputs(4900));
    outputs(2132) <= (layer0_outputs(5046)) xor (layer0_outputs(9989));
    outputs(2133) <= not(layer0_outputs(1596));
    outputs(2134) <= not((layer0_outputs(4021)) xor (layer0_outputs(3775)));
    outputs(2135) <= not(layer0_outputs(3820));
    outputs(2136) <= layer0_outputs(10028);
    outputs(2137) <= not((layer0_outputs(272)) xor (layer0_outputs(4563)));
    outputs(2138) <= not((layer0_outputs(1311)) and (layer0_outputs(7806)));
    outputs(2139) <= not(layer0_outputs(3455)) or (layer0_outputs(3839));
    outputs(2140) <= not(layer0_outputs(7525)) or (layer0_outputs(6342));
    outputs(2141) <= (layer0_outputs(2554)) xor (layer0_outputs(9116));
    outputs(2142) <= layer0_outputs(9289);
    outputs(2143) <= layer0_outputs(194);
    outputs(2144) <= layer0_outputs(7984);
    outputs(2145) <= layer0_outputs(7106);
    outputs(2146) <= (layer0_outputs(2738)) and (layer0_outputs(8339));
    outputs(2147) <= not((layer0_outputs(2040)) xor (layer0_outputs(3421)));
    outputs(2148) <= layer0_outputs(4845);
    outputs(2149) <= not((layer0_outputs(8316)) xor (layer0_outputs(57)));
    outputs(2150) <= (layer0_outputs(5605)) and not (layer0_outputs(7743));
    outputs(2151) <= layer0_outputs(2887);
    outputs(2152) <= not((layer0_outputs(7778)) xor (layer0_outputs(2695)));
    outputs(2153) <= not((layer0_outputs(4693)) xor (layer0_outputs(4324)));
    outputs(2154) <= layer0_outputs(7015);
    outputs(2155) <= not(layer0_outputs(258)) or (layer0_outputs(3430));
    outputs(2156) <= not(layer0_outputs(3492));
    outputs(2157) <= layer0_outputs(6202);
    outputs(2158) <= (layer0_outputs(1211)) xor (layer0_outputs(939));
    outputs(2159) <= not(layer0_outputs(8835));
    outputs(2160) <= layer0_outputs(7469);
    outputs(2161) <= not((layer0_outputs(5354)) xor (layer0_outputs(9939)));
    outputs(2162) <= layer0_outputs(1081);
    outputs(2163) <= not(layer0_outputs(3695));
    outputs(2164) <= not(layer0_outputs(6723));
    outputs(2165) <= not(layer0_outputs(5850));
    outputs(2166) <= not(layer0_outputs(4526)) or (layer0_outputs(2449));
    outputs(2167) <= not((layer0_outputs(4839)) xor (layer0_outputs(9492)));
    outputs(2168) <= layer0_outputs(5033);
    outputs(2169) <= not(layer0_outputs(6965)) or (layer0_outputs(2171));
    outputs(2170) <= not(layer0_outputs(4982));
    outputs(2171) <= not(layer0_outputs(4897));
    outputs(2172) <= not((layer0_outputs(6127)) and (layer0_outputs(8681)));
    outputs(2173) <= not((layer0_outputs(3189)) xor (layer0_outputs(6917)));
    outputs(2174) <= not(layer0_outputs(5826));
    outputs(2175) <= not(layer0_outputs(2019)) or (layer0_outputs(5722));
    outputs(2176) <= layer0_outputs(668);
    outputs(2177) <= layer0_outputs(1680);
    outputs(2178) <= not(layer0_outputs(9732));
    outputs(2179) <= not((layer0_outputs(1928)) or (layer0_outputs(2784)));
    outputs(2180) <= layer0_outputs(2614);
    outputs(2181) <= not(layer0_outputs(2185)) or (layer0_outputs(2346));
    outputs(2182) <= not((layer0_outputs(3794)) xor (layer0_outputs(7318)));
    outputs(2183) <= layer0_outputs(5462);
    outputs(2184) <= not((layer0_outputs(4367)) xor (layer0_outputs(10031)));
    outputs(2185) <= not(layer0_outputs(6551));
    outputs(2186) <= layer0_outputs(8408);
    outputs(2187) <= (layer0_outputs(9438)) and not (layer0_outputs(9240));
    outputs(2188) <= not(layer0_outputs(2319));
    outputs(2189) <= layer0_outputs(2670);
    outputs(2190) <= (layer0_outputs(1939)) or (layer0_outputs(6676));
    outputs(2191) <= (layer0_outputs(4423)) and not (layer0_outputs(10053));
    outputs(2192) <= not(layer0_outputs(816));
    outputs(2193) <= not((layer0_outputs(1804)) xor (layer0_outputs(10134)));
    outputs(2194) <= '1';
    outputs(2195) <= (layer0_outputs(2757)) xor (layer0_outputs(8667));
    outputs(2196) <= not(layer0_outputs(3421));
    outputs(2197) <= not(layer0_outputs(5174));
    outputs(2198) <= (layer0_outputs(954)) xor (layer0_outputs(9680));
    outputs(2199) <= not(layer0_outputs(9244));
    outputs(2200) <= layer0_outputs(503);
    outputs(2201) <= not(layer0_outputs(6080));
    outputs(2202) <= not(layer0_outputs(2957));
    outputs(2203) <= not(layer0_outputs(7774));
    outputs(2204) <= not(layer0_outputs(6440));
    outputs(2205) <= not(layer0_outputs(1653)) or (layer0_outputs(7575));
    outputs(2206) <= layer0_outputs(5453);
    outputs(2207) <= not((layer0_outputs(1439)) and (layer0_outputs(7827)));
    outputs(2208) <= layer0_outputs(2855);
    outputs(2209) <= not(layer0_outputs(833));
    outputs(2210) <= (layer0_outputs(2410)) xor (layer0_outputs(2465));
    outputs(2211) <= not(layer0_outputs(1248));
    outputs(2212) <= (layer0_outputs(3136)) xor (layer0_outputs(9803));
    outputs(2213) <= (layer0_outputs(9823)) and not (layer0_outputs(9074));
    outputs(2214) <= layer0_outputs(2398);
    outputs(2215) <= (layer0_outputs(2103)) xor (layer0_outputs(10089));
    outputs(2216) <= not(layer0_outputs(10098));
    outputs(2217) <= not(layer0_outputs(1552));
    outputs(2218) <= not(layer0_outputs(3079));
    outputs(2219) <= (layer0_outputs(5405)) and not (layer0_outputs(7599));
    outputs(2220) <= layer0_outputs(8576);
    outputs(2221) <= not(layer0_outputs(4720));
    outputs(2222) <= (layer0_outputs(2324)) or (layer0_outputs(7017));
    outputs(2223) <= not(layer0_outputs(2659));
    outputs(2224) <= layer0_outputs(1123);
    outputs(2225) <= not(layer0_outputs(4256));
    outputs(2226) <= not(layer0_outputs(1027)) or (layer0_outputs(5856));
    outputs(2227) <= not((layer0_outputs(6904)) and (layer0_outputs(7382)));
    outputs(2228) <= not(layer0_outputs(6345));
    outputs(2229) <= not(layer0_outputs(4695));
    outputs(2230) <= (layer0_outputs(2684)) xor (layer0_outputs(4386));
    outputs(2231) <= (layer0_outputs(9125)) and not (layer0_outputs(3014));
    outputs(2232) <= not(layer0_outputs(9734));
    outputs(2233) <= (layer0_outputs(8527)) and not (layer0_outputs(906));
    outputs(2234) <= not(layer0_outputs(2442));
    outputs(2235) <= not(layer0_outputs(9838));
    outputs(2236) <= (layer0_outputs(685)) and (layer0_outputs(6129));
    outputs(2237) <= not((layer0_outputs(6288)) xor (layer0_outputs(9236)));
    outputs(2238) <= layer0_outputs(2196);
    outputs(2239) <= (layer0_outputs(4503)) or (layer0_outputs(1138));
    outputs(2240) <= not(layer0_outputs(4052)) or (layer0_outputs(1436));
    outputs(2241) <= layer0_outputs(5921);
    outputs(2242) <= (layer0_outputs(1422)) xor (layer0_outputs(312));
    outputs(2243) <= (layer0_outputs(6386)) and (layer0_outputs(7602));
    outputs(2244) <= (layer0_outputs(3625)) xor (layer0_outputs(7786));
    outputs(2245) <= (layer0_outputs(34)) xor (layer0_outputs(847));
    outputs(2246) <= layer0_outputs(9948);
    outputs(2247) <= layer0_outputs(8163);
    outputs(2248) <= layer0_outputs(8584);
    outputs(2249) <= not(layer0_outputs(7885));
    outputs(2250) <= not(layer0_outputs(5300));
    outputs(2251) <= layer0_outputs(9431);
    outputs(2252) <= not((layer0_outputs(8937)) xor (layer0_outputs(9819)));
    outputs(2253) <= not((layer0_outputs(3182)) xor (layer0_outputs(7708)));
    outputs(2254) <= not(layer0_outputs(3838));
    outputs(2255) <= layer0_outputs(5438);
    outputs(2256) <= not(layer0_outputs(9187)) or (layer0_outputs(520));
    outputs(2257) <= not(layer0_outputs(397)) or (layer0_outputs(260));
    outputs(2258) <= not(layer0_outputs(4727));
    outputs(2259) <= layer0_outputs(7206);
    outputs(2260) <= not(layer0_outputs(6432));
    outputs(2261) <= layer0_outputs(4061);
    outputs(2262) <= not((layer0_outputs(2020)) and (layer0_outputs(5782)));
    outputs(2263) <= not(layer0_outputs(2403));
    outputs(2264) <= (layer0_outputs(3271)) and (layer0_outputs(6327));
    outputs(2265) <= not((layer0_outputs(6152)) xor (layer0_outputs(9468)));
    outputs(2266) <= layer0_outputs(6489);
    outputs(2267) <= not(layer0_outputs(6012));
    outputs(2268) <= not((layer0_outputs(9622)) or (layer0_outputs(6954)));
    outputs(2269) <= not(layer0_outputs(8894));
    outputs(2270) <= layer0_outputs(8768);
    outputs(2271) <= (layer0_outputs(1039)) or (layer0_outputs(9759));
    outputs(2272) <= not(layer0_outputs(2339));
    outputs(2273) <= not((layer0_outputs(6624)) xor (layer0_outputs(731)));
    outputs(2274) <= not(layer0_outputs(8660)) or (layer0_outputs(7757));
    outputs(2275) <= not(layer0_outputs(1363));
    outputs(2276) <= layer0_outputs(8843);
    outputs(2277) <= (layer0_outputs(10164)) xor (layer0_outputs(472));
    outputs(2278) <= (layer0_outputs(4082)) or (layer0_outputs(7270));
    outputs(2279) <= not(layer0_outputs(7899));
    outputs(2280) <= not(layer0_outputs(564));
    outputs(2281) <= (layer0_outputs(7773)) xor (layer0_outputs(1371));
    outputs(2282) <= not(layer0_outputs(1344));
    outputs(2283) <= not(layer0_outputs(75)) or (layer0_outputs(6748));
    outputs(2284) <= not((layer0_outputs(8602)) xor (layer0_outputs(5612)));
    outputs(2285) <= (layer0_outputs(4107)) xor (layer0_outputs(4493));
    outputs(2286) <= layer0_outputs(3688);
    outputs(2287) <= not((layer0_outputs(8579)) and (layer0_outputs(1916)));
    outputs(2288) <= not(layer0_outputs(6560));
    outputs(2289) <= (layer0_outputs(7745)) and (layer0_outputs(1861));
    outputs(2290) <= layer0_outputs(3175);
    outputs(2291) <= not(layer0_outputs(6452)) or (layer0_outputs(1976));
    outputs(2292) <= layer0_outputs(5128);
    outputs(2293) <= (layer0_outputs(6040)) xor (layer0_outputs(1069));
    outputs(2294) <= layer0_outputs(3207);
    outputs(2295) <= not(layer0_outputs(3286));
    outputs(2296) <= not(layer0_outputs(7342)) or (layer0_outputs(6848));
    outputs(2297) <= (layer0_outputs(6414)) and not (layer0_outputs(2703));
    outputs(2298) <= layer0_outputs(8145);
    outputs(2299) <= not((layer0_outputs(9381)) or (layer0_outputs(10224)));
    outputs(2300) <= layer0_outputs(2787);
    outputs(2301) <= layer0_outputs(2956);
    outputs(2302) <= layer0_outputs(9415);
    outputs(2303) <= not((layer0_outputs(217)) and (layer0_outputs(8321)));
    outputs(2304) <= (layer0_outputs(1905)) xor (layer0_outputs(3443));
    outputs(2305) <= not(layer0_outputs(4004));
    outputs(2306) <= not(layer0_outputs(3955));
    outputs(2307) <= layer0_outputs(4714);
    outputs(2308) <= (layer0_outputs(8272)) xor (layer0_outputs(2089));
    outputs(2309) <= not((layer0_outputs(5281)) xor (layer0_outputs(10187)));
    outputs(2310) <= layer0_outputs(8189);
    outputs(2311) <= (layer0_outputs(1848)) and not (layer0_outputs(8364));
    outputs(2312) <= not(layer0_outputs(3622)) or (layer0_outputs(2690));
    outputs(2313) <= (layer0_outputs(379)) and (layer0_outputs(3717));
    outputs(2314) <= not(layer0_outputs(8502));
    outputs(2315) <= layer0_outputs(8808);
    outputs(2316) <= (layer0_outputs(3335)) and (layer0_outputs(9324));
    outputs(2317) <= layer0_outputs(7488);
    outputs(2318) <= layer0_outputs(8474);
    outputs(2319) <= layer0_outputs(4254);
    outputs(2320) <= not((layer0_outputs(9216)) xor (layer0_outputs(4463)));
    outputs(2321) <= (layer0_outputs(1244)) xor (layer0_outputs(9653));
    outputs(2322) <= not(layer0_outputs(7975));
    outputs(2323) <= not(layer0_outputs(9864)) or (layer0_outputs(3645));
    outputs(2324) <= not(layer0_outputs(658));
    outputs(2325) <= not(layer0_outputs(1266));
    outputs(2326) <= (layer0_outputs(6544)) xor (layer0_outputs(8903));
    outputs(2327) <= not(layer0_outputs(3803));
    outputs(2328) <= not(layer0_outputs(8497));
    outputs(2329) <= layer0_outputs(6696);
    outputs(2330) <= layer0_outputs(376);
    outputs(2331) <= layer0_outputs(1419);
    outputs(2332) <= not((layer0_outputs(1489)) xor (layer0_outputs(5387)));
    outputs(2333) <= not((layer0_outputs(5886)) xor (layer0_outputs(6568)));
    outputs(2334) <= not(layer0_outputs(3212)) or (layer0_outputs(4880));
    outputs(2335) <= (layer0_outputs(7264)) xor (layer0_outputs(8338));
    outputs(2336) <= layer0_outputs(1106);
    outputs(2337) <= layer0_outputs(2918);
    outputs(2338) <= (layer0_outputs(8025)) xor (layer0_outputs(3641));
    outputs(2339) <= not((layer0_outputs(7879)) or (layer0_outputs(8514)));
    outputs(2340) <= layer0_outputs(9530);
    outputs(2341) <= not(layer0_outputs(5574));
    outputs(2342) <= (layer0_outputs(3883)) xor (layer0_outputs(9096));
    outputs(2343) <= layer0_outputs(3213);
    outputs(2344) <= layer0_outputs(5753);
    outputs(2345) <= not((layer0_outputs(2796)) or (layer0_outputs(9768)));
    outputs(2346) <= layer0_outputs(7442);
    outputs(2347) <= layer0_outputs(3563);
    outputs(2348) <= not((layer0_outputs(6925)) xor (layer0_outputs(6340)));
    outputs(2349) <= layer0_outputs(5790);
    outputs(2350) <= not(layer0_outputs(3762));
    outputs(2351) <= not((layer0_outputs(15)) or (layer0_outputs(5971)));
    outputs(2352) <= not(layer0_outputs(1726));
    outputs(2353) <= layer0_outputs(7304);
    outputs(2354) <= not((layer0_outputs(6535)) and (layer0_outputs(1583)));
    outputs(2355) <= not(layer0_outputs(2285));
    outputs(2356) <= layer0_outputs(1505);
    outputs(2357) <= (layer0_outputs(5625)) and (layer0_outputs(8138));
    outputs(2358) <= not(layer0_outputs(7014));
    outputs(2359) <= (layer0_outputs(349)) xor (layer0_outputs(7055));
    outputs(2360) <= not(layer0_outputs(9879));
    outputs(2361) <= layer0_outputs(4126);
    outputs(2362) <= not(layer0_outputs(7905));
    outputs(2363) <= layer0_outputs(10237);
    outputs(2364) <= layer0_outputs(2232);
    outputs(2365) <= (layer0_outputs(8734)) and not (layer0_outputs(5808));
    outputs(2366) <= not((layer0_outputs(2212)) xor (layer0_outputs(2656)));
    outputs(2367) <= not(layer0_outputs(6407)) or (layer0_outputs(1958));
    outputs(2368) <= layer0_outputs(9754);
    outputs(2369) <= layer0_outputs(3577);
    outputs(2370) <= not(layer0_outputs(8553));
    outputs(2371) <= not(layer0_outputs(6699)) or (layer0_outputs(76));
    outputs(2372) <= layer0_outputs(4204);
    outputs(2373) <= layer0_outputs(2200);
    outputs(2374) <= layer0_outputs(2761);
    outputs(2375) <= not(layer0_outputs(1610)) or (layer0_outputs(3565));
    outputs(2376) <= not((layer0_outputs(2868)) or (layer0_outputs(7574)));
    outputs(2377) <= not((layer0_outputs(5167)) and (layer0_outputs(835)));
    outputs(2378) <= not((layer0_outputs(8948)) or (layer0_outputs(9624)));
    outputs(2379) <= not((layer0_outputs(569)) xor (layer0_outputs(8563)));
    outputs(2380) <= not(layer0_outputs(5432));
    outputs(2381) <= not(layer0_outputs(543));
    outputs(2382) <= not(layer0_outputs(4364)) or (layer0_outputs(2117));
    outputs(2383) <= not(layer0_outputs(7946)) or (layer0_outputs(994));
    outputs(2384) <= layer0_outputs(5813);
    outputs(2385) <= layer0_outputs(2543);
    outputs(2386) <= layer0_outputs(6565);
    outputs(2387) <= not((layer0_outputs(2395)) xor (layer0_outputs(2035)));
    outputs(2388) <= (layer0_outputs(5240)) or (layer0_outputs(8024));
    outputs(2389) <= layer0_outputs(1179);
    outputs(2390) <= not(layer0_outputs(2325)) or (layer0_outputs(5627));
    outputs(2391) <= layer0_outputs(3506);
    outputs(2392) <= not(layer0_outputs(6782));
    outputs(2393) <= not((layer0_outputs(8992)) xor (layer0_outputs(6937)));
    outputs(2394) <= not(layer0_outputs(9955)) or (layer0_outputs(5441));
    outputs(2395) <= not(layer0_outputs(116));
    outputs(2396) <= not(layer0_outputs(2476));
    outputs(2397) <= not(layer0_outputs(257));
    outputs(2398) <= not(layer0_outputs(8948));
    outputs(2399) <= not((layer0_outputs(6652)) xor (layer0_outputs(4080)));
    outputs(2400) <= layer0_outputs(2915);
    outputs(2401) <= (layer0_outputs(526)) xor (layer0_outputs(612));
    outputs(2402) <= layer0_outputs(6794);
    outputs(2403) <= not((layer0_outputs(4208)) xor (layer0_outputs(7706)));
    outputs(2404) <= (layer0_outputs(8493)) xor (layer0_outputs(6476));
    outputs(2405) <= not(layer0_outputs(5608));
    outputs(2406) <= not(layer0_outputs(9120));
    outputs(2407) <= not(layer0_outputs(3820));
    outputs(2408) <= layer0_outputs(7580);
    outputs(2409) <= (layer0_outputs(7551)) xor (layer0_outputs(3326));
    outputs(2410) <= not(layer0_outputs(4455));
    outputs(2411) <= not(layer0_outputs(10014));
    outputs(2412) <= not(layer0_outputs(5829));
    outputs(2413) <= (layer0_outputs(5145)) or (layer0_outputs(5134));
    outputs(2414) <= not(layer0_outputs(7586));
    outputs(2415) <= layer0_outputs(9482);
    outputs(2416) <= not(layer0_outputs(335));
    outputs(2417) <= not(layer0_outputs(93));
    outputs(2418) <= not(layer0_outputs(415));
    outputs(2419) <= (layer0_outputs(6349)) xor (layer0_outputs(6604));
    outputs(2420) <= (layer0_outputs(10176)) xor (layer0_outputs(6259));
    outputs(2421) <= layer0_outputs(6356);
    outputs(2422) <= not(layer0_outputs(1813));
    outputs(2423) <= (layer0_outputs(2484)) and not (layer0_outputs(7812));
    outputs(2424) <= layer0_outputs(3855);
    outputs(2425) <= not(layer0_outputs(8962));
    outputs(2426) <= layer0_outputs(930);
    outputs(2427) <= not(layer0_outputs(1877));
    outputs(2428) <= not(layer0_outputs(5549));
    outputs(2429) <= layer0_outputs(9970);
    outputs(2430) <= layer0_outputs(6389);
    outputs(2431) <= not((layer0_outputs(2672)) or (layer0_outputs(8934)));
    outputs(2432) <= layer0_outputs(6892);
    outputs(2433) <= not((layer0_outputs(367)) xor (layer0_outputs(2854)));
    outputs(2434) <= (layer0_outputs(5573)) or (layer0_outputs(4784));
    outputs(2435) <= (layer0_outputs(3385)) and not (layer0_outputs(7522));
    outputs(2436) <= layer0_outputs(5186);
    outputs(2437) <= layer0_outputs(1638);
    outputs(2438) <= not(layer0_outputs(6664));
    outputs(2439) <= not((layer0_outputs(5494)) xor (layer0_outputs(4090)));
    outputs(2440) <= not((layer0_outputs(8267)) xor (layer0_outputs(1182)));
    outputs(2441) <= layer0_outputs(2335);
    outputs(2442) <= not(layer0_outputs(8242));
    outputs(2443) <= not(layer0_outputs(4681));
    outputs(2444) <= (layer0_outputs(6281)) xor (layer0_outputs(6874));
    outputs(2445) <= not((layer0_outputs(16)) xor (layer0_outputs(5043)));
    outputs(2446) <= (layer0_outputs(2748)) and (layer0_outputs(2106));
    outputs(2447) <= not(layer0_outputs(6108));
    outputs(2448) <= layer0_outputs(2323);
    outputs(2449) <= layer0_outputs(4943);
    outputs(2450) <= layer0_outputs(7973);
    outputs(2451) <= (layer0_outputs(8839)) and not (layer0_outputs(6277));
    outputs(2452) <= (layer0_outputs(3081)) or (layer0_outputs(2812));
    outputs(2453) <= layer0_outputs(9509);
    outputs(2454) <= not(layer0_outputs(227)) or (layer0_outputs(159));
    outputs(2455) <= not((layer0_outputs(3211)) xor (layer0_outputs(4787)));
    outputs(2456) <= layer0_outputs(5351);
    outputs(2457) <= not(layer0_outputs(4877));
    outputs(2458) <= layer0_outputs(1863);
    outputs(2459) <= layer0_outputs(499);
    outputs(2460) <= not(layer0_outputs(1700)) or (layer0_outputs(3586));
    outputs(2461) <= layer0_outputs(961);
    outputs(2462) <= layer0_outputs(3260);
    outputs(2463) <= not(layer0_outputs(3803)) or (layer0_outputs(9132));
    outputs(2464) <= not((layer0_outputs(4)) xor (layer0_outputs(4676)));
    outputs(2465) <= (layer0_outputs(383)) xor (layer0_outputs(9310));
    outputs(2466) <= not((layer0_outputs(9961)) and (layer0_outputs(2498)));
    outputs(2467) <= layer0_outputs(566);
    outputs(2468) <= layer0_outputs(9731);
    outputs(2469) <= (layer0_outputs(2785)) and not (layer0_outputs(5144));
    outputs(2470) <= not(layer0_outputs(5307));
    outputs(2471) <= layer0_outputs(8376);
    outputs(2472) <= not(layer0_outputs(7985));
    outputs(2473) <= not(layer0_outputs(9781)) or (layer0_outputs(8636));
    outputs(2474) <= layer0_outputs(7135);
    outputs(2475) <= (layer0_outputs(4604)) and not (layer0_outputs(3230));
    outputs(2476) <= (layer0_outputs(3205)) xor (layer0_outputs(4539));
    outputs(2477) <= not(layer0_outputs(7971)) or (layer0_outputs(3656));
    outputs(2478) <= layer0_outputs(6876);
    outputs(2479) <= not(layer0_outputs(1251)) or (layer0_outputs(5373));
    outputs(2480) <= not((layer0_outputs(6090)) and (layer0_outputs(8028)));
    outputs(2481) <= not(layer0_outputs(147));
    outputs(2482) <= (layer0_outputs(301)) or (layer0_outputs(6677));
    outputs(2483) <= not(layer0_outputs(4903));
    outputs(2484) <= layer0_outputs(4417);
    outputs(2485) <= not(layer0_outputs(4141));
    outputs(2486) <= (layer0_outputs(3214)) xor (layer0_outputs(9136));
    outputs(2487) <= layer0_outputs(1371);
    outputs(2488) <= (layer0_outputs(3114)) xor (layer0_outputs(890));
    outputs(2489) <= layer0_outputs(7230);
    outputs(2490) <= not(layer0_outputs(6438));
    outputs(2491) <= not(layer0_outputs(1114));
    outputs(2492) <= not(layer0_outputs(5512));
    outputs(2493) <= not((layer0_outputs(6685)) and (layer0_outputs(2599)));
    outputs(2494) <= not(layer0_outputs(4181));
    outputs(2495) <= layer0_outputs(128);
    outputs(2496) <= (layer0_outputs(9253)) and not (layer0_outputs(5109));
    outputs(2497) <= not((layer0_outputs(2073)) xor (layer0_outputs(284)));
    outputs(2498) <= (layer0_outputs(5231)) or (layer0_outputs(4428));
    outputs(2499) <= (layer0_outputs(818)) xor (layer0_outputs(2567));
    outputs(2500) <= layer0_outputs(5720);
    outputs(2501) <= (layer0_outputs(8941)) and not (layer0_outputs(4457));
    outputs(2502) <= not(layer0_outputs(3201));
    outputs(2503) <= not(layer0_outputs(7329));
    outputs(2504) <= not(layer0_outputs(1871));
    outputs(2505) <= not(layer0_outputs(6798));
    outputs(2506) <= (layer0_outputs(9772)) or (layer0_outputs(4953));
    outputs(2507) <= not(layer0_outputs(5108)) or (layer0_outputs(6180));
    outputs(2508) <= not((layer0_outputs(7495)) xor (layer0_outputs(5088)));
    outputs(2509) <= (layer0_outputs(2049)) xor (layer0_outputs(2978));
    outputs(2510) <= layer0_outputs(441);
    outputs(2511) <= (layer0_outputs(9380)) and (layer0_outputs(9372));
    outputs(2512) <= layer0_outputs(5624);
    outputs(2513) <= not(layer0_outputs(4871));
    outputs(2514) <= not(layer0_outputs(2476));
    outputs(2515) <= not((layer0_outputs(6067)) xor (layer0_outputs(8627)));
    outputs(2516) <= not(layer0_outputs(2148)) or (layer0_outputs(6773));
    outputs(2517) <= layer0_outputs(6048);
    outputs(2518) <= layer0_outputs(5870);
    outputs(2519) <= layer0_outputs(10028);
    outputs(2520) <= (layer0_outputs(7010)) xor (layer0_outputs(6632));
    outputs(2521) <= (layer0_outputs(2025)) xor (layer0_outputs(6746));
    outputs(2522) <= layer0_outputs(2789);
    outputs(2523) <= layer0_outputs(1418);
    outputs(2524) <= not(layer0_outputs(4022));
    outputs(2525) <= not(layer0_outputs(366));
    outputs(2526) <= not((layer0_outputs(6755)) xor (layer0_outputs(1258)));
    outputs(2527) <= not(layer0_outputs(4077)) or (layer0_outputs(6996));
    outputs(2528) <= not(layer0_outputs(250));
    outputs(2529) <= not(layer0_outputs(7636));
    outputs(2530) <= layer0_outputs(5993);
    outputs(2531) <= (layer0_outputs(152)) xor (layer0_outputs(1335));
    outputs(2532) <= not(layer0_outputs(5445));
    outputs(2533) <= (layer0_outputs(7217)) and not (layer0_outputs(6772));
    outputs(2534) <= layer0_outputs(2010);
    outputs(2535) <= not((layer0_outputs(4024)) xor (layer0_outputs(6839)));
    outputs(2536) <= layer0_outputs(4291);
    outputs(2537) <= not(layer0_outputs(5791));
    outputs(2538) <= (layer0_outputs(1434)) xor (layer0_outputs(3631));
    outputs(2539) <= not((layer0_outputs(1547)) and (layer0_outputs(7543)));
    outputs(2540) <= not(layer0_outputs(4077));
    outputs(2541) <= not(layer0_outputs(3789));
    outputs(2542) <= (layer0_outputs(9350)) and (layer0_outputs(7612));
    outputs(2543) <= (layer0_outputs(66)) or (layer0_outputs(3939));
    outputs(2544) <= (layer0_outputs(628)) or (layer0_outputs(9069));
    outputs(2545) <= (layer0_outputs(4996)) xor (layer0_outputs(369));
    outputs(2546) <= not((layer0_outputs(46)) and (layer0_outputs(6426)));
    outputs(2547) <= not((layer0_outputs(5859)) or (layer0_outputs(7976)));
    outputs(2548) <= not((layer0_outputs(5755)) or (layer0_outputs(9741)));
    outputs(2549) <= not(layer0_outputs(2775));
    outputs(2550) <= layer0_outputs(4339);
    outputs(2551) <= layer0_outputs(8878);
    outputs(2552) <= (layer0_outputs(9532)) xor (layer0_outputs(3356));
    outputs(2553) <= (layer0_outputs(5238)) and not (layer0_outputs(2194));
    outputs(2554) <= layer0_outputs(1838);
    outputs(2555) <= (layer0_outputs(2181)) xor (layer0_outputs(9201));
    outputs(2556) <= not(layer0_outputs(4862));
    outputs(2557) <= not(layer0_outputs(4978));
    outputs(2558) <= not(layer0_outputs(6448));
    outputs(2559) <= (layer0_outputs(5023)) or (layer0_outputs(4480));
    outputs(2560) <= not(layer0_outputs(8143));
    outputs(2561) <= not((layer0_outputs(2920)) or (layer0_outputs(5598)));
    outputs(2562) <= layer0_outputs(5064);
    outputs(2563) <= not(layer0_outputs(5306));
    outputs(2564) <= not(layer0_outputs(6764));
    outputs(2565) <= not(layer0_outputs(6099));
    outputs(2566) <= not(layer0_outputs(1200));
    outputs(2567) <= not(layer0_outputs(8741)) or (layer0_outputs(1606));
    outputs(2568) <= (layer0_outputs(9481)) and (layer0_outputs(6607));
    outputs(2569) <= (layer0_outputs(2749)) and not (layer0_outputs(8146));
    outputs(2570) <= not(layer0_outputs(8104));
    outputs(2571) <= not((layer0_outputs(339)) xor (layer0_outputs(9368)));
    outputs(2572) <= layer0_outputs(9569);
    outputs(2573) <= layer0_outputs(212);
    outputs(2574) <= layer0_outputs(7296);
    outputs(2575) <= layer0_outputs(501);
    outputs(2576) <= layer0_outputs(8037);
    outputs(2577) <= not(layer0_outputs(9197));
    outputs(2578) <= not(layer0_outputs(4210));
    outputs(2579) <= (layer0_outputs(3069)) and (layer0_outputs(4627));
    outputs(2580) <= not(layer0_outputs(2446));
    outputs(2581) <= layer0_outputs(5510);
    outputs(2582) <= layer0_outputs(1790);
    outputs(2583) <= not((layer0_outputs(512)) and (layer0_outputs(560)));
    outputs(2584) <= not(layer0_outputs(6544)) or (layer0_outputs(4477));
    outputs(2585) <= not((layer0_outputs(6661)) and (layer0_outputs(4634)));
    outputs(2586) <= not(layer0_outputs(6971));
    outputs(2587) <= (layer0_outputs(7793)) or (layer0_outputs(2982));
    outputs(2588) <= not(layer0_outputs(7868));
    outputs(2589) <= layer0_outputs(9433);
    outputs(2590) <= layer0_outputs(9215);
    outputs(2591) <= not(layer0_outputs(5089));
    outputs(2592) <= not((layer0_outputs(2291)) xor (layer0_outputs(1714)));
    outputs(2593) <= layer0_outputs(8335);
    outputs(2594) <= (layer0_outputs(3348)) xor (layer0_outputs(4479));
    outputs(2595) <= not(layer0_outputs(9722)) or (layer0_outputs(3405));
    outputs(2596) <= not((layer0_outputs(2601)) xor (layer0_outputs(5264)));
    outputs(2597) <= not((layer0_outputs(8089)) or (layer0_outputs(1023)));
    outputs(2598) <= (layer0_outputs(5332)) and not (layer0_outputs(7954));
    outputs(2599) <= not(layer0_outputs(5734));
    outputs(2600) <= (layer0_outputs(2239)) and (layer0_outputs(7096));
    outputs(2601) <= not(layer0_outputs(3526));
    outputs(2602) <= (layer0_outputs(5588)) or (layer0_outputs(3087));
    outputs(2603) <= not(layer0_outputs(10038));
    outputs(2604) <= not(layer0_outputs(9571));
    outputs(2605) <= layer0_outputs(1364);
    outputs(2606) <= layer0_outputs(5708);
    outputs(2607) <= (layer0_outputs(3763)) or (layer0_outputs(3976));
    outputs(2608) <= layer0_outputs(9966);
    outputs(2609) <= (layer0_outputs(2519)) and not (layer0_outputs(4744));
    outputs(2610) <= not(layer0_outputs(5322)) or (layer0_outputs(8698));
    outputs(2611) <= not(layer0_outputs(3748));
    outputs(2612) <= not((layer0_outputs(4118)) xor (layer0_outputs(3897)));
    outputs(2613) <= (layer0_outputs(156)) and (layer0_outputs(9048));
    outputs(2614) <= layer0_outputs(1938);
    outputs(2615) <= not(layer0_outputs(1591)) or (layer0_outputs(6997));
    outputs(2616) <= not(layer0_outputs(1053));
    outputs(2617) <= not((layer0_outputs(9581)) xor (layer0_outputs(3050)));
    outputs(2618) <= not(layer0_outputs(277)) or (layer0_outputs(5577));
    outputs(2619) <= layer0_outputs(8179);
    outputs(2620) <= not(layer0_outputs(103));
    outputs(2621) <= not(layer0_outputs(1870));
    outputs(2622) <= layer0_outputs(236);
    outputs(2623) <= not(layer0_outputs(3202)) or (layer0_outputs(616));
    outputs(2624) <= layer0_outputs(6136);
    outputs(2625) <= (layer0_outputs(4812)) xor (layer0_outputs(6270));
    outputs(2626) <= not(layer0_outputs(2638));
    outputs(2627) <= not(layer0_outputs(5571));
    outputs(2628) <= layer0_outputs(2528);
    outputs(2629) <= not(layer0_outputs(9630)) or (layer0_outputs(8311));
    outputs(2630) <= (layer0_outputs(5690)) or (layer0_outputs(4950));
    outputs(2631) <= layer0_outputs(9328);
    outputs(2632) <= not(layer0_outputs(9912));
    outputs(2633) <= not((layer0_outputs(3582)) xor (layer0_outputs(6808)));
    outputs(2634) <= not((layer0_outputs(1095)) xor (layer0_outputs(1187)));
    outputs(2635) <= not((layer0_outputs(8755)) and (layer0_outputs(8866)));
    outputs(2636) <= (layer0_outputs(6363)) xor (layer0_outputs(2017));
    outputs(2637) <= not((layer0_outputs(6761)) xor (layer0_outputs(8050)));
    outputs(2638) <= layer0_outputs(7377);
    outputs(2639) <= not((layer0_outputs(829)) xor (layer0_outputs(9466)));
    outputs(2640) <= not((layer0_outputs(2009)) or (layer0_outputs(2663)));
    outputs(2641) <= layer0_outputs(7347);
    outputs(2642) <= (layer0_outputs(2539)) xor (layer0_outputs(286));
    outputs(2643) <= (layer0_outputs(3511)) or (layer0_outputs(5125));
    outputs(2644) <= not((layer0_outputs(3060)) xor (layer0_outputs(5930)));
    outputs(2645) <= not((layer0_outputs(9506)) and (layer0_outputs(5526)));
    outputs(2646) <= not((layer0_outputs(2090)) xor (layer0_outputs(9747)));
    outputs(2647) <= (layer0_outputs(3698)) or (layer0_outputs(5320));
    outputs(2648) <= layer0_outputs(5887);
    outputs(2649) <= not(layer0_outputs(189));
    outputs(2650) <= not((layer0_outputs(6158)) xor (layer0_outputs(1365)));
    outputs(2651) <= not((layer0_outputs(3082)) xor (layer0_outputs(8205)));
    outputs(2652) <= (layer0_outputs(478)) xor (layer0_outputs(442));
    outputs(2653) <= not(layer0_outputs(8544));
    outputs(2654) <= layer0_outputs(3686);
    outputs(2655) <= not(layer0_outputs(8976));
    outputs(2656) <= layer0_outputs(6814);
    outputs(2657) <= not(layer0_outputs(6354)) or (layer0_outputs(1976));
    outputs(2658) <= not((layer0_outputs(6322)) xor (layer0_outputs(8510)));
    outputs(2659) <= not((layer0_outputs(4601)) and (layer0_outputs(1983)));
    outputs(2660) <= not(layer0_outputs(1881));
    outputs(2661) <= not(layer0_outputs(3395));
    outputs(2662) <= not(layer0_outputs(1679));
    outputs(2663) <= not(layer0_outputs(6254));
    outputs(2664) <= not(layer0_outputs(3644));
    outputs(2665) <= not(layer0_outputs(8523));
    outputs(2666) <= layer0_outputs(8263);
    outputs(2667) <= not(layer0_outputs(9510));
    outputs(2668) <= not((layer0_outputs(4760)) or (layer0_outputs(5826)));
    outputs(2669) <= (layer0_outputs(583)) and not (layer0_outputs(7555));
    outputs(2670) <= layer0_outputs(6317);
    outputs(2671) <= (layer0_outputs(2994)) and not (layer0_outputs(6809));
    outputs(2672) <= (layer0_outputs(736)) xor (layer0_outputs(4075));
    outputs(2673) <= not(layer0_outputs(549));
    outputs(2674) <= not(layer0_outputs(7904));
    outputs(2675) <= layer0_outputs(8587);
    outputs(2676) <= layer0_outputs(3615);
    outputs(2677) <= (layer0_outputs(8697)) and not (layer0_outputs(2394));
    outputs(2678) <= layer0_outputs(5862);
    outputs(2679) <= not(layer0_outputs(800)) or (layer0_outputs(9067));
    outputs(2680) <= not(layer0_outputs(2442));
    outputs(2681) <= not(layer0_outputs(4869));
    outputs(2682) <= not(layer0_outputs(6220)) or (layer0_outputs(2700));
    outputs(2683) <= not(layer0_outputs(5179));
    outputs(2684) <= layer0_outputs(5945);
    outputs(2685) <= (layer0_outputs(5890)) xor (layer0_outputs(6148));
    outputs(2686) <= layer0_outputs(1632);
    outputs(2687) <= layer0_outputs(2197);
    outputs(2688) <= not(layer0_outputs(1832)) or (layer0_outputs(1507));
    outputs(2689) <= not(layer0_outputs(9767));
    outputs(2690) <= not(layer0_outputs(6547));
    outputs(2691) <= not((layer0_outputs(1622)) xor (layer0_outputs(1055)));
    outputs(2692) <= not(layer0_outputs(2524));
    outputs(2693) <= layer0_outputs(1130);
    outputs(2694) <= layer0_outputs(757);
    outputs(2695) <= layer0_outputs(4599);
    outputs(2696) <= layer0_outputs(65);
    outputs(2697) <= layer0_outputs(8290);
    outputs(2698) <= layer0_outputs(2899);
    outputs(2699) <= not(layer0_outputs(4340)) or (layer0_outputs(5682));
    outputs(2700) <= not(layer0_outputs(5236));
    outputs(2701) <= layer0_outputs(6630);
    outputs(2702) <= layer0_outputs(780);
    outputs(2703) <= not(layer0_outputs(1924));
    outputs(2704) <= not((layer0_outputs(8909)) and (layer0_outputs(2125)));
    outputs(2705) <= (layer0_outputs(3327)) and not (layer0_outputs(4924));
    outputs(2706) <= not((layer0_outputs(389)) and (layer0_outputs(8586)));
    outputs(2707) <= not(layer0_outputs(9905));
    outputs(2708) <= (layer0_outputs(4952)) or (layer0_outputs(1221));
    outputs(2709) <= (layer0_outputs(7728)) and (layer0_outputs(7664));
    outputs(2710) <= layer0_outputs(72);
    outputs(2711) <= (layer0_outputs(6151)) xor (layer0_outputs(7426));
    outputs(2712) <= layer0_outputs(3011);
    outputs(2713) <= not((layer0_outputs(48)) and (layer0_outputs(3937)));
    outputs(2714) <= layer0_outputs(5858);
    outputs(2715) <= not(layer0_outputs(4514));
    outputs(2716) <= (layer0_outputs(2739)) xor (layer0_outputs(5851));
    outputs(2717) <= not((layer0_outputs(1612)) xor (layer0_outputs(1670)));
    outputs(2718) <= (layer0_outputs(3860)) and not (layer0_outputs(801));
    outputs(2719) <= layer0_outputs(0);
    outputs(2720) <= not((layer0_outputs(3046)) and (layer0_outputs(6991)));
    outputs(2721) <= (layer0_outputs(10016)) xor (layer0_outputs(9046));
    outputs(2722) <= (layer0_outputs(8228)) or (layer0_outputs(8198));
    outputs(2723) <= not((layer0_outputs(8153)) or (layer0_outputs(1036)));
    outputs(2724) <= (layer0_outputs(4716)) or (layer0_outputs(1305));
    outputs(2725) <= (layer0_outputs(1680)) and not (layer0_outputs(970));
    outputs(2726) <= not((layer0_outputs(2306)) and (layer0_outputs(2392)));
    outputs(2727) <= layer0_outputs(273);
    outputs(2728) <= not(layer0_outputs(677));
    outputs(2729) <= not(layer0_outputs(1252)) or (layer0_outputs(3293));
    outputs(2730) <= (layer0_outputs(5026)) xor (layer0_outputs(8670));
    outputs(2731) <= layer0_outputs(2990);
    outputs(2732) <= (layer0_outputs(798)) and not (layer0_outputs(5797));
    outputs(2733) <= layer0_outputs(8412);
    outputs(2734) <= not(layer0_outputs(7815));
    outputs(2735) <= layer0_outputs(2905);
    outputs(2736) <= not(layer0_outputs(9883));
    outputs(2737) <= not((layer0_outputs(2007)) xor (layer0_outputs(4458)));
    outputs(2738) <= not((layer0_outputs(242)) xor (layer0_outputs(922)));
    outputs(2739) <= layer0_outputs(1220);
    outputs(2740) <= not((layer0_outputs(1538)) or (layer0_outputs(8536)));
    outputs(2741) <= not((layer0_outputs(9876)) and (layer0_outputs(9850)));
    outputs(2742) <= (layer0_outputs(828)) xor (layer0_outputs(992));
    outputs(2743) <= not(layer0_outputs(2960));
    outputs(2744) <= layer0_outputs(1897);
    outputs(2745) <= not(layer0_outputs(1427)) or (layer0_outputs(3377));
    outputs(2746) <= not((layer0_outputs(10116)) xor (layer0_outputs(5557)));
    outputs(2747) <= layer0_outputs(5456);
    outputs(2748) <= layer0_outputs(756);
    outputs(2749) <= not(layer0_outputs(5505));
    outputs(2750) <= (layer0_outputs(8537)) xor (layer0_outputs(2053));
    outputs(2751) <= not((layer0_outputs(7598)) xor (layer0_outputs(7121)));
    outputs(2752) <= layer0_outputs(4334);
    outputs(2753) <= not((layer0_outputs(2450)) xor (layer0_outputs(6502)));
    outputs(2754) <= layer0_outputs(6356);
    outputs(2755) <= (layer0_outputs(4560)) and not (layer0_outputs(3124));
    outputs(2756) <= layer0_outputs(7920);
    outputs(2757) <= (layer0_outputs(1007)) xor (layer0_outputs(9653));
    outputs(2758) <= layer0_outputs(31);
    outputs(2759) <= not(layer0_outputs(8307));
    outputs(2760) <= not(layer0_outputs(1324)) or (layer0_outputs(641));
    outputs(2761) <= layer0_outputs(3588);
    outputs(2762) <= not((layer0_outputs(9496)) xor (layer0_outputs(2692)));
    outputs(2763) <= not((layer0_outputs(6975)) and (layer0_outputs(8184)));
    outputs(2764) <= layer0_outputs(6079);
    outputs(2765) <= not(layer0_outputs(9395));
    outputs(2766) <= (layer0_outputs(10045)) and (layer0_outputs(4061));
    outputs(2767) <= not(layer0_outputs(5956));
    outputs(2768) <= layer0_outputs(581);
    outputs(2769) <= not(layer0_outputs(2270)) or (layer0_outputs(8179));
    outputs(2770) <= not(layer0_outputs(7671)) or (layer0_outputs(7440));
    outputs(2771) <= layer0_outputs(3088);
    outputs(2772) <= layer0_outputs(10214);
    outputs(2773) <= (layer0_outputs(5012)) xor (layer0_outputs(825));
    outputs(2774) <= not((layer0_outputs(10021)) or (layer0_outputs(3590)));
    outputs(2775) <= not(layer0_outputs(2906));
    outputs(2776) <= not(layer0_outputs(9190));
    outputs(2777) <= not(layer0_outputs(3852));
    outputs(2778) <= layer0_outputs(4249);
    outputs(2779) <= layer0_outputs(9131);
    outputs(2780) <= layer0_outputs(8895);
    outputs(2781) <= layer0_outputs(7447);
    outputs(2782) <= not((layer0_outputs(10073)) or (layer0_outputs(9574)));
    outputs(2783) <= layer0_outputs(9022);
    outputs(2784) <= layer0_outputs(10006);
    outputs(2785) <= (layer0_outputs(5917)) xor (layer0_outputs(4447));
    outputs(2786) <= not(layer0_outputs(1096)) or (layer0_outputs(9298));
    outputs(2787) <= layer0_outputs(7736);
    outputs(2788) <= not(layer0_outputs(8543));
    outputs(2789) <= layer0_outputs(2329);
    outputs(2790) <= not(layer0_outputs(3125));
    outputs(2791) <= not(layer0_outputs(3303));
    outputs(2792) <= layer0_outputs(2370);
    outputs(2793) <= layer0_outputs(6922);
    outputs(2794) <= not(layer0_outputs(8089)) or (layer0_outputs(10188));
    outputs(2795) <= not(layer0_outputs(294));
    outputs(2796) <= not(layer0_outputs(794));
    outputs(2797) <= layer0_outputs(29);
    outputs(2798) <= not((layer0_outputs(4421)) xor (layer0_outputs(2977)));
    outputs(2799) <= not(layer0_outputs(4440)) or (layer0_outputs(8507));
    outputs(2800) <= layer0_outputs(1825);
    outputs(2801) <= (layer0_outputs(9877)) and not (layer0_outputs(4945));
    outputs(2802) <= not((layer0_outputs(2340)) and (layer0_outputs(8261)));
    outputs(2803) <= (layer0_outputs(8489)) and not (layer0_outputs(4050));
    outputs(2804) <= not(layer0_outputs(4205)) or (layer0_outputs(10021));
    outputs(2805) <= (layer0_outputs(6982)) and not (layer0_outputs(8630));
    outputs(2806) <= layer0_outputs(7825);
    outputs(2807) <= (layer0_outputs(4644)) xor (layer0_outputs(8265));
    outputs(2808) <= not(layer0_outputs(6659));
    outputs(2809) <= not(layer0_outputs(7522));
    outputs(2810) <= layer0_outputs(1328);
    outputs(2811) <= (layer0_outputs(6639)) and not (layer0_outputs(5594));
    outputs(2812) <= not(layer0_outputs(3595));
    outputs(2813) <= layer0_outputs(6414);
    outputs(2814) <= layer0_outputs(3289);
    outputs(2815) <= layer0_outputs(8455);
    outputs(2816) <= (layer0_outputs(5885)) and not (layer0_outputs(2245));
    outputs(2817) <= (layer0_outputs(3467)) or (layer0_outputs(5117));
    outputs(2818) <= not(layer0_outputs(2270)) or (layer0_outputs(2242));
    outputs(2819) <= not(layer0_outputs(6112));
    outputs(2820) <= (layer0_outputs(4114)) xor (layer0_outputs(10174));
    outputs(2821) <= not(layer0_outputs(7957));
    outputs(2822) <= not(layer0_outputs(4275));
    outputs(2823) <= layer0_outputs(9970);
    outputs(2824) <= layer0_outputs(1569);
    outputs(2825) <= not(layer0_outputs(10200));
    outputs(2826) <= (layer0_outputs(1177)) or (layer0_outputs(2111));
    outputs(2827) <= not(layer0_outputs(7641));
    outputs(2828) <= not(layer0_outputs(944));
    outputs(2829) <= not((layer0_outputs(4485)) xor (layer0_outputs(8930)));
    outputs(2830) <= layer0_outputs(1502);
    outputs(2831) <= layer0_outputs(49);
    outputs(2832) <= not(layer0_outputs(3848));
    outputs(2833) <= not((layer0_outputs(1137)) xor (layer0_outputs(3726)));
    outputs(2834) <= (layer0_outputs(2434)) or (layer0_outputs(210));
    outputs(2835) <= not(layer0_outputs(6407)) or (layer0_outputs(10151));
    outputs(2836) <= not(layer0_outputs(3131)) or (layer0_outputs(7353));
    outputs(2837) <= not((layer0_outputs(8190)) and (layer0_outputs(5489)));
    outputs(2838) <= not(layer0_outputs(4607)) or (layer0_outputs(5363));
    outputs(2839) <= (layer0_outputs(8282)) or (layer0_outputs(811));
    outputs(2840) <= not(layer0_outputs(6541)) or (layer0_outputs(9334));
    outputs(2841) <= not((layer0_outputs(3136)) xor (layer0_outputs(230)));
    outputs(2842) <= not(layer0_outputs(3821)) or (layer0_outputs(6933));
    outputs(2843) <= layer0_outputs(5357);
    outputs(2844) <= not((layer0_outputs(5522)) xor (layer0_outputs(1500)));
    outputs(2845) <= layer0_outputs(2560);
    outputs(2846) <= not(layer0_outputs(5629)) or (layer0_outputs(1682));
    outputs(2847) <= not(layer0_outputs(3884));
    outputs(2848) <= layer0_outputs(4332);
    outputs(2849) <= layer0_outputs(8715);
    outputs(2850) <= layer0_outputs(9597);
    outputs(2851) <= not(layer0_outputs(7744)) or (layer0_outputs(8592));
    outputs(2852) <= not((layer0_outputs(9604)) xor (layer0_outputs(3399)));
    outputs(2853) <= layer0_outputs(0);
    outputs(2854) <= not(layer0_outputs(7723)) or (layer0_outputs(4232));
    outputs(2855) <= not(layer0_outputs(6649)) or (layer0_outputs(2547));
    outputs(2856) <= not(layer0_outputs(3296));
    outputs(2857) <= not(layer0_outputs(541));
    outputs(2858) <= not(layer0_outputs(9184));
    outputs(2859) <= not(layer0_outputs(6863));
    outputs(2860) <= layer0_outputs(8504);
    outputs(2861) <= not((layer0_outputs(1675)) and (layer0_outputs(6563)));
    outputs(2862) <= not(layer0_outputs(5752));
    outputs(2863) <= not(layer0_outputs(1535));
    outputs(2864) <= (layer0_outputs(5362)) xor (layer0_outputs(8801));
    outputs(2865) <= (layer0_outputs(3529)) and not (layer0_outputs(3078));
    outputs(2866) <= (layer0_outputs(3552)) xor (layer0_outputs(1292));
    outputs(2867) <= not(layer0_outputs(5107)) or (layer0_outputs(7102));
    outputs(2868) <= layer0_outputs(8600);
    outputs(2869) <= not(layer0_outputs(8838));
    outputs(2870) <= layer0_outputs(8973);
    outputs(2871) <= (layer0_outputs(6749)) and (layer0_outputs(1999));
    outputs(2872) <= not(layer0_outputs(2267));
    outputs(2873) <= not(layer0_outputs(3490)) or (layer0_outputs(7644));
    outputs(2874) <= not((layer0_outputs(9952)) or (layer0_outputs(4236)));
    outputs(2875) <= layer0_outputs(5660);
    outputs(2876) <= not(layer0_outputs(185));
    outputs(2877) <= not(layer0_outputs(9740)) or (layer0_outputs(4065));
    outputs(2878) <= not(layer0_outputs(5271));
    outputs(2879) <= (layer0_outputs(3722)) and not (layer0_outputs(7391));
    outputs(2880) <= not((layer0_outputs(2461)) xor (layer0_outputs(6126)));
    outputs(2881) <= not(layer0_outputs(9511));
    outputs(2882) <= not((layer0_outputs(8497)) and (layer0_outputs(1164)));
    outputs(2883) <= not(layer0_outputs(9239));
    outputs(2884) <= not(layer0_outputs(8403));
    outputs(2885) <= not(layer0_outputs(4626)) or (layer0_outputs(772));
    outputs(2886) <= (layer0_outputs(7392)) xor (layer0_outputs(2723));
    outputs(2887) <= (layer0_outputs(735)) and not (layer0_outputs(8078));
    outputs(2888) <= not(layer0_outputs(8707));
    outputs(2889) <= layer0_outputs(4005);
    outputs(2890) <= layer0_outputs(4304);
    outputs(2891) <= (layer0_outputs(4278)) or (layer0_outputs(2204));
    outputs(2892) <= (layer0_outputs(6272)) and (layer0_outputs(5927));
    outputs(2893) <= layer0_outputs(930);
    outputs(2894) <= (layer0_outputs(2842)) xor (layer0_outputs(3055));
    outputs(2895) <= layer0_outputs(4291);
    outputs(2896) <= not((layer0_outputs(8339)) xor (layer0_outputs(5324)));
    outputs(2897) <= layer0_outputs(3077);
    outputs(2898) <= not((layer0_outputs(1169)) xor (layer0_outputs(8232)));
    outputs(2899) <= not((layer0_outputs(7022)) xor (layer0_outputs(7278)));
    outputs(2900) <= (layer0_outputs(4107)) and (layer0_outputs(6813));
    outputs(2901) <= not((layer0_outputs(2418)) xor (layer0_outputs(3388)));
    outputs(2902) <= (layer0_outputs(5340)) and not (layer0_outputs(6074));
    outputs(2903) <= (layer0_outputs(4466)) xor (layer0_outputs(4449));
    outputs(2904) <= not(layer0_outputs(1085)) or (layer0_outputs(1839));
    outputs(2905) <= not((layer0_outputs(8611)) xor (layer0_outputs(9812)));
    outputs(2906) <= (layer0_outputs(4587)) and (layer0_outputs(3730));
    outputs(2907) <= (layer0_outputs(7724)) or (layer0_outputs(2843));
    outputs(2908) <= not(layer0_outputs(198));
    outputs(2909) <= not(layer0_outputs(7435));
    outputs(2910) <= layer0_outputs(460);
    outputs(2911) <= layer0_outputs(2608);
    outputs(2912) <= not((layer0_outputs(8917)) xor (layer0_outputs(5239)));
    outputs(2913) <= not(layer0_outputs(462));
    outputs(2914) <= not(layer0_outputs(1199));
    outputs(2915) <= not(layer0_outputs(4056));
    outputs(2916) <= (layer0_outputs(1918)) and not (layer0_outputs(2157));
    outputs(2917) <= not(layer0_outputs(761));
    outputs(2918) <= not(layer0_outputs(6072));
    outputs(2919) <= (layer0_outputs(8802)) and (layer0_outputs(2830));
    outputs(2920) <= not((layer0_outputs(3697)) xor (layer0_outputs(3281)));
    outputs(2921) <= (layer0_outputs(7103)) xor (layer0_outputs(4736));
    outputs(2922) <= (layer0_outputs(5473)) xor (layer0_outputs(9576));
    outputs(2923) <= not(layer0_outputs(7200));
    outputs(2924) <= (layer0_outputs(1315)) xor (layer0_outputs(2728));
    outputs(2925) <= not(layer0_outputs(548));
    outputs(2926) <= (layer0_outputs(6226)) xor (layer0_outputs(6205));
    outputs(2927) <= (layer0_outputs(1910)) or (layer0_outputs(5156));
    outputs(2928) <= layer0_outputs(4426);
    outputs(2929) <= (layer0_outputs(275)) xor (layer0_outputs(8223));
    outputs(2930) <= not(layer0_outputs(9261));
    outputs(2931) <= layer0_outputs(4350);
    outputs(2932) <= not(layer0_outputs(3364)) or (layer0_outputs(8392));
    outputs(2933) <= (layer0_outputs(1954)) and not (layer0_outputs(4215));
    outputs(2934) <= (layer0_outputs(2051)) or (layer0_outputs(10235));
    outputs(2935) <= not(layer0_outputs(7617)) or (layer0_outputs(2616));
    outputs(2936) <= not(layer0_outputs(9024)) or (layer0_outputs(4623));
    outputs(2937) <= (layer0_outputs(156)) and (layer0_outputs(3491));
    outputs(2938) <= (layer0_outputs(7692)) xor (layer0_outputs(9749));
    outputs(2939) <= layer0_outputs(9504);
    outputs(2940) <= not((layer0_outputs(6626)) xor (layer0_outputs(9348)));
    outputs(2941) <= not(layer0_outputs(4586));
    outputs(2942) <= layer0_outputs(871);
    outputs(2943) <= (layer0_outputs(7010)) and (layer0_outputs(14));
    outputs(2944) <= (layer0_outputs(9226)) and (layer0_outputs(3963));
    outputs(2945) <= layer0_outputs(3358);
    outputs(2946) <= not(layer0_outputs(2076));
    outputs(2947) <= layer0_outputs(9771);
    outputs(2948) <= layer0_outputs(3843);
    outputs(2949) <= (layer0_outputs(9606)) and not (layer0_outputs(9700));
    outputs(2950) <= layer0_outputs(4001);
    outputs(2951) <= layer0_outputs(2281);
    outputs(2952) <= layer0_outputs(6750);
    outputs(2953) <= not((layer0_outputs(6169)) or (layer0_outputs(7375)));
    outputs(2954) <= layer0_outputs(3831);
    outputs(2955) <= not(layer0_outputs(341));
    outputs(2956) <= not((layer0_outputs(7673)) and (layer0_outputs(3559)));
    outputs(2957) <= not(layer0_outputs(3494));
    outputs(2958) <= not(layer0_outputs(8580));
    outputs(2959) <= not(layer0_outputs(3247));
    outputs(2960) <= not((layer0_outputs(6483)) and (layer0_outputs(3927)));
    outputs(2961) <= (layer0_outputs(3362)) xor (layer0_outputs(3447));
    outputs(2962) <= layer0_outputs(9958);
    outputs(2963) <= not(layer0_outputs(9286));
    outputs(2964) <= layer0_outputs(2848);
    outputs(2965) <= (layer0_outputs(5288)) and not (layer0_outputs(8620));
    outputs(2966) <= not(layer0_outputs(4976));
    outputs(2967) <= layer0_outputs(4132);
    outputs(2968) <= not(layer0_outputs(8643));
    outputs(2969) <= not(layer0_outputs(9163)) or (layer0_outputs(7339));
    outputs(2970) <= not(layer0_outputs(3580)) or (layer0_outputs(228));
    outputs(2971) <= layer0_outputs(5049);
    outputs(2972) <= not(layer0_outputs(7772)) or (layer0_outputs(5230));
    outputs(2973) <= (layer0_outputs(199)) xor (layer0_outputs(1985));
    outputs(2974) <= not(layer0_outputs(5160));
    outputs(2975) <= not(layer0_outputs(5803)) or (layer0_outputs(5320));
    outputs(2976) <= (layer0_outputs(5446)) and not (layer0_outputs(3844));
    outputs(2977) <= layer0_outputs(8836);
    outputs(2978) <= not((layer0_outputs(4732)) and (layer0_outputs(1454)));
    outputs(2979) <= not((layer0_outputs(9665)) xor (layer0_outputs(7775)));
    outputs(2980) <= layer0_outputs(2141);
    outputs(2981) <= (layer0_outputs(6572)) or (layer0_outputs(8369));
    outputs(2982) <= (layer0_outputs(5951)) xor (layer0_outputs(7947));
    outputs(2983) <= (layer0_outputs(1521)) and (layer0_outputs(8192));
    outputs(2984) <= layer0_outputs(5033);
    outputs(2985) <= not(layer0_outputs(1713));
    outputs(2986) <= layer0_outputs(3981);
    outputs(2987) <= not(layer0_outputs(7519));
    outputs(2988) <= layer0_outputs(9895);
    outputs(2989) <= (layer0_outputs(4010)) and (layer0_outputs(2348));
    outputs(2990) <= (layer0_outputs(5615)) xor (layer0_outputs(1133));
    outputs(2991) <= not((layer0_outputs(5258)) xor (layer0_outputs(5352)));
    outputs(2992) <= layer0_outputs(1588);
    outputs(2993) <= not(layer0_outputs(9560)) or (layer0_outputs(4019));
    outputs(2994) <= layer0_outputs(3087);
    outputs(2995) <= not(layer0_outputs(1312));
    outputs(2996) <= not(layer0_outputs(820));
    outputs(2997) <= not(layer0_outputs(6908));
    outputs(2998) <= not(layer0_outputs(7670));
    outputs(2999) <= not((layer0_outputs(9434)) xor (layer0_outputs(10071)));
    outputs(3000) <= not(layer0_outputs(5835));
    outputs(3001) <= not((layer0_outputs(3847)) and (layer0_outputs(2693)));
    outputs(3002) <= layer0_outputs(4576);
    outputs(3003) <= layer0_outputs(3750);
    outputs(3004) <= not((layer0_outputs(5702)) and (layer0_outputs(3257)));
    outputs(3005) <= not((layer0_outputs(2203)) and (layer0_outputs(4333)));
    outputs(3006) <= not((layer0_outputs(41)) xor (layer0_outputs(9564)));
    outputs(3007) <= not(layer0_outputs(4942));
    outputs(3008) <= (layer0_outputs(10197)) xor (layer0_outputs(3481));
    outputs(3009) <= layer0_outputs(3610);
    outputs(3010) <= not((layer0_outputs(9180)) or (layer0_outputs(8618)));
    outputs(3011) <= not(layer0_outputs(3796)) or (layer0_outputs(10083));
    outputs(3012) <= (layer0_outputs(5774)) and (layer0_outputs(4920));
    outputs(3013) <= not((layer0_outputs(9913)) or (layer0_outputs(162)));
    outputs(3014) <= not(layer0_outputs(6550));
    outputs(3015) <= not(layer0_outputs(7393));
    outputs(3016) <= not(layer0_outputs(5699));
    outputs(3017) <= not((layer0_outputs(1899)) xor (layer0_outputs(7132)));
    outputs(3018) <= not((layer0_outputs(6323)) xor (layer0_outputs(2412)));
    outputs(3019) <= not(layer0_outputs(5810)) or (layer0_outputs(2277));
    outputs(3020) <= (layer0_outputs(5436)) and not (layer0_outputs(2394));
    outputs(3021) <= layer0_outputs(2295);
    outputs(3022) <= not(layer0_outputs(3992));
    outputs(3023) <= not((layer0_outputs(7153)) xor (layer0_outputs(852)));
    outputs(3024) <= not(layer0_outputs(2526)) or (layer0_outputs(7684));
    outputs(3025) <= layer0_outputs(5553);
    outputs(3026) <= not((layer0_outputs(9085)) xor (layer0_outputs(381)));
    outputs(3027) <= not((layer0_outputs(9020)) xor (layer0_outputs(6447)));
    outputs(3028) <= not((layer0_outputs(8629)) and (layer0_outputs(7605)));
    outputs(3029) <= (layer0_outputs(8017)) or (layer0_outputs(2666));
    outputs(3030) <= layer0_outputs(961);
    outputs(3031) <= layer0_outputs(8831);
    outputs(3032) <= not(layer0_outputs(9051));
    outputs(3033) <= layer0_outputs(2329);
    outputs(3034) <= not((layer0_outputs(1190)) or (layer0_outputs(267)));
    outputs(3035) <= (layer0_outputs(7655)) xor (layer0_outputs(5099));
    outputs(3036) <= not(layer0_outputs(656));
    outputs(3037) <= not((layer0_outputs(6712)) or (layer0_outputs(5087)));
    outputs(3038) <= (layer0_outputs(6330)) and not (layer0_outputs(6951));
    outputs(3039) <= layer0_outputs(1217);
    outputs(3040) <= (layer0_outputs(10124)) or (layer0_outputs(9393));
    outputs(3041) <= not(layer0_outputs(5105));
    outputs(3042) <= (layer0_outputs(4303)) xor (layer0_outputs(1421));
    outputs(3043) <= (layer0_outputs(386)) and (layer0_outputs(5508));
    outputs(3044) <= not(layer0_outputs(10092)) or (layer0_outputs(5031));
    outputs(3045) <= not((layer0_outputs(404)) xor (layer0_outputs(8972)));
    outputs(3046) <= not(layer0_outputs(7181));
    outputs(3047) <= not(layer0_outputs(1205));
    outputs(3048) <= layer0_outputs(7731);
    outputs(3049) <= layer0_outputs(1622);
    outputs(3050) <= (layer0_outputs(9925)) xor (layer0_outputs(8012));
    outputs(3051) <= not(layer0_outputs(609));
    outputs(3052) <= not(layer0_outputs(4151));
    outputs(3053) <= layer0_outputs(5063);
    outputs(3054) <= not(layer0_outputs(6664));
    outputs(3055) <= not(layer0_outputs(3139));
    outputs(3056) <= not(layer0_outputs(7942)) or (layer0_outputs(6173));
    outputs(3057) <= not(layer0_outputs(1528)) or (layer0_outputs(4311));
    outputs(3058) <= layer0_outputs(2169);
    outputs(3059) <= not(layer0_outputs(6720)) or (layer0_outputs(7793));
    outputs(3060) <= not(layer0_outputs(2763)) or (layer0_outputs(4948));
    outputs(3061) <= layer0_outputs(3923);
    outputs(3062) <= layer0_outputs(7595);
    outputs(3063) <= not(layer0_outputs(8345));
    outputs(3064) <= not(layer0_outputs(1278));
    outputs(3065) <= not(layer0_outputs(3353));
    outputs(3066) <= layer0_outputs(9501);
    outputs(3067) <= (layer0_outputs(6624)) and (layer0_outputs(2568));
    outputs(3068) <= not(layer0_outputs(9088));
    outputs(3069) <= layer0_outputs(1390);
    outputs(3070) <= not((layer0_outputs(1479)) xor (layer0_outputs(9713)));
    outputs(3071) <= not(layer0_outputs(5211));
    outputs(3072) <= not(layer0_outputs(9804)) or (layer0_outputs(2728));
    outputs(3073) <= not(layer0_outputs(6236));
    outputs(3074) <= layer0_outputs(5652);
    outputs(3075) <= not(layer0_outputs(2485));
    outputs(3076) <= not((layer0_outputs(4741)) xor (layer0_outputs(5368)));
    outputs(3077) <= not(layer0_outputs(7536));
    outputs(3078) <= layer0_outputs(9026);
    outputs(3079) <= layer0_outputs(7597);
    outputs(3080) <= not(layer0_outputs(7759));
    outputs(3081) <= not((layer0_outputs(3517)) xor (layer0_outputs(6952)));
    outputs(3082) <= not(layer0_outputs(3411));
    outputs(3083) <= (layer0_outputs(5157)) xor (layer0_outputs(243));
    outputs(3084) <= not(layer0_outputs(8860)) or (layer0_outputs(4202));
    outputs(3085) <= (layer0_outputs(9423)) and (layer0_outputs(7537));
    outputs(3086) <= not(layer0_outputs(5497));
    outputs(3087) <= not(layer0_outputs(5015));
    outputs(3088) <= layer0_outputs(8675);
    outputs(3089) <= layer0_outputs(2961);
    outputs(3090) <= not(layer0_outputs(2276)) or (layer0_outputs(9601));
    outputs(3091) <= not((layer0_outputs(2468)) and (layer0_outputs(6347)));
    outputs(3092) <= layer0_outputs(2138);
    outputs(3093) <= not(layer0_outputs(1325)) or (layer0_outputs(9025));
    outputs(3094) <= not(layer0_outputs(5689));
    outputs(3095) <= (layer0_outputs(1863)) xor (layer0_outputs(3186));
    outputs(3096) <= layer0_outputs(7405);
    outputs(3097) <= layer0_outputs(2111);
    outputs(3098) <= not((layer0_outputs(2393)) xor (layer0_outputs(111)));
    outputs(3099) <= (layer0_outputs(3480)) xor (layer0_outputs(10196));
    outputs(3100) <= not(layer0_outputs(4902));
    outputs(3101) <= not(layer0_outputs(4376));
    outputs(3102) <= (layer0_outputs(1605)) and not (layer0_outputs(3043));
    outputs(3103) <= layer0_outputs(595);
    outputs(3104) <= not(layer0_outputs(8589));
    outputs(3105) <= not(layer0_outputs(7524)) or (layer0_outputs(9938));
    outputs(3106) <= layer0_outputs(5953);
    outputs(3107) <= (layer0_outputs(8129)) or (layer0_outputs(7434));
    outputs(3108) <= (layer0_outputs(68)) and not (layer0_outputs(3268));
    outputs(3109) <= not(layer0_outputs(7847));
    outputs(3110) <= layer0_outputs(6689);
    outputs(3111) <= not(layer0_outputs(5270));
    outputs(3112) <= (layer0_outputs(245)) and not (layer0_outputs(468));
    outputs(3113) <= not((layer0_outputs(6605)) and (layer0_outputs(4428)));
    outputs(3114) <= not((layer0_outputs(471)) xor (layer0_outputs(7751)));
    outputs(3115) <= not((layer0_outputs(3474)) xor (layer0_outputs(7788)));
    outputs(3116) <= layer0_outputs(8389);
    outputs(3117) <= layer0_outputs(8245);
    outputs(3118) <= layer0_outputs(9191);
    outputs(3119) <= not((layer0_outputs(4399)) xor (layer0_outputs(6075)));
    outputs(3120) <= not((layer0_outputs(3947)) xor (layer0_outputs(549)));
    outputs(3121) <= not(layer0_outputs(8554));
    outputs(3122) <= layer0_outputs(644);
    outputs(3123) <= not(layer0_outputs(2656)) or (layer0_outputs(9994));
    outputs(3124) <= not((layer0_outputs(10018)) xor (layer0_outputs(263)));
    outputs(3125) <= layer0_outputs(168);
    outputs(3126) <= not(layer0_outputs(10190));
    outputs(3127) <= not(layer0_outputs(9995));
    outputs(3128) <= (layer0_outputs(2920)) and not (layer0_outputs(576));
    outputs(3129) <= not((layer0_outputs(2685)) xor (layer0_outputs(6599)));
    outputs(3130) <= not(layer0_outputs(693));
    outputs(3131) <= not(layer0_outputs(5502));
    outputs(3132) <= (layer0_outputs(600)) xor (layer0_outputs(4039));
    outputs(3133) <= not(layer0_outputs(6257));
    outputs(3134) <= not(layer0_outputs(7530));
    outputs(3135) <= (layer0_outputs(9059)) and not (layer0_outputs(5539));
    outputs(3136) <= (layer0_outputs(4236)) or (layer0_outputs(10153));
    outputs(3137) <= (layer0_outputs(1901)) xor (layer0_outputs(6277));
    outputs(3138) <= not(layer0_outputs(2444));
    outputs(3139) <= (layer0_outputs(9149)) and not (layer0_outputs(6967));
    outputs(3140) <= (layer0_outputs(1563)) xor (layer0_outputs(7897));
    outputs(3141) <= not(layer0_outputs(3654));
    outputs(3142) <= not(layer0_outputs(5737));
    outputs(3143) <= (layer0_outputs(9990)) xor (layer0_outputs(3296));
    outputs(3144) <= not((layer0_outputs(8156)) or (layer0_outputs(3057)));
    outputs(3145) <= (layer0_outputs(4009)) and not (layer0_outputs(2982));
    outputs(3146) <= layer0_outputs(2231);
    outputs(3147) <= (layer0_outputs(2316)) and (layer0_outputs(9011));
    outputs(3148) <= not(layer0_outputs(9555));
    outputs(3149) <= not(layer0_outputs(5818));
    outputs(3150) <= not((layer0_outputs(2716)) xor (layer0_outputs(9983)));
    outputs(3151) <= (layer0_outputs(7215)) and not (layer0_outputs(7440));
    outputs(3152) <= (layer0_outputs(3837)) and (layer0_outputs(3611));
    outputs(3153) <= not(layer0_outputs(8621));
    outputs(3154) <= (layer0_outputs(3500)) and not (layer0_outputs(986));
    outputs(3155) <= layer0_outputs(1821);
    outputs(3156) <= not((layer0_outputs(6067)) and (layer0_outputs(9962)));
    outputs(3157) <= layer0_outputs(8222);
    outputs(3158) <= not(layer0_outputs(4375));
    outputs(3159) <= (layer0_outputs(1191)) and not (layer0_outputs(8113));
    outputs(3160) <= layer0_outputs(5703);
    outputs(3161) <= not(layer0_outputs(5264));
    outputs(3162) <= (layer0_outputs(2439)) and not (layer0_outputs(3392));
    outputs(3163) <= not((layer0_outputs(2627)) xor (layer0_outputs(8467)));
    outputs(3164) <= (layer0_outputs(3849)) xor (layer0_outputs(2919));
    outputs(3165) <= (layer0_outputs(7947)) xor (layer0_outputs(1006));
    outputs(3166) <= (layer0_outputs(8304)) and (layer0_outputs(4684));
    outputs(3167) <= layer0_outputs(2917);
    outputs(3168) <= not((layer0_outputs(1758)) and (layer0_outputs(1267)));
    outputs(3169) <= layer0_outputs(6491);
    outputs(3170) <= not(layer0_outputs(6587));
    outputs(3171) <= not(layer0_outputs(2101));
    outputs(3172) <= layer0_outputs(9241);
    outputs(3173) <= not(layer0_outputs(6703));
    outputs(3174) <= not(layer0_outputs(3528));
    outputs(3175) <= layer0_outputs(4394);
    outputs(3176) <= (layer0_outputs(2311)) xor (layer0_outputs(5801));
    outputs(3177) <= layer0_outputs(9627);
    outputs(3178) <= not((layer0_outputs(7381)) or (layer0_outputs(3482)));
    outputs(3179) <= layer0_outputs(1873);
    outputs(3180) <= (layer0_outputs(5375)) and (layer0_outputs(5718));
    outputs(3181) <= not((layer0_outputs(5847)) xor (layer0_outputs(4728)));
    outputs(3182) <= layer0_outputs(8413);
    outputs(3183) <= not((layer0_outputs(7560)) or (layer0_outputs(8386)));
    outputs(3184) <= not(layer0_outputs(2145));
    outputs(3185) <= layer0_outputs(6223);
    outputs(3186) <= not(layer0_outputs(3120));
    outputs(3187) <= not((layer0_outputs(8303)) xor (layer0_outputs(8532)));
    outputs(3188) <= (layer0_outputs(7444)) and not (layer0_outputs(3588));
    outputs(3189) <= not((layer0_outputs(5557)) xor (layer0_outputs(3840)));
    outputs(3190) <= layer0_outputs(5778);
    outputs(3191) <= not((layer0_outputs(3064)) xor (layer0_outputs(2892)));
    outputs(3192) <= not(layer0_outputs(4816));
    outputs(3193) <= layer0_outputs(4622);
    outputs(3194) <= not((layer0_outputs(1912)) xor (layer0_outputs(7766)));
    outputs(3195) <= not(layer0_outputs(6398)) or (layer0_outputs(4455));
    outputs(3196) <= layer0_outputs(2483);
    outputs(3197) <= not(layer0_outputs(4705));
    outputs(3198) <= not((layer0_outputs(1780)) or (layer0_outputs(4280)));
    outputs(3199) <= not(layer0_outputs(7248)) or (layer0_outputs(6376));
    outputs(3200) <= not((layer0_outputs(9775)) or (layer0_outputs(5843)));
    outputs(3201) <= (layer0_outputs(5663)) xor (layer0_outputs(4511));
    outputs(3202) <= not(layer0_outputs(9823)) or (layer0_outputs(7702));
    outputs(3203) <= (layer0_outputs(2987)) xor (layer0_outputs(7477));
    outputs(3204) <= not(layer0_outputs(5973));
    outputs(3205) <= not((layer0_outputs(544)) xor (layer0_outputs(8847)));
    outputs(3206) <= layer0_outputs(2202);
    outputs(3207) <= not(layer0_outputs(2228));
    outputs(3208) <= layer0_outputs(8324);
    outputs(3209) <= (layer0_outputs(9454)) and (layer0_outputs(2360));
    outputs(3210) <= not(layer0_outputs(1767));
    outputs(3211) <= (layer0_outputs(9434)) xor (layer0_outputs(9278));
    outputs(3212) <= not(layer0_outputs(6463));
    outputs(3213) <= not(layer0_outputs(9597));
    outputs(3214) <= not(layer0_outputs(9121));
    outputs(3215) <= layer0_outputs(5524);
    outputs(3216) <= not(layer0_outputs(831)) or (layer0_outputs(9117));
    outputs(3217) <= layer0_outputs(9018);
    outputs(3218) <= not((layer0_outputs(5700)) xor (layer0_outputs(3946)));
    outputs(3219) <= layer0_outputs(3426);
    outputs(3220) <= layer0_outputs(7921);
    outputs(3221) <= layer0_outputs(9644);
    outputs(3222) <= not((layer0_outputs(148)) xor (layer0_outputs(2582)));
    outputs(3223) <= layer0_outputs(3752);
    outputs(3224) <= layer0_outputs(8848);
    outputs(3225) <= layer0_outputs(1038);
    outputs(3226) <= (layer0_outputs(5492)) xor (layer0_outputs(7146));
    outputs(3227) <= (layer0_outputs(1562)) xor (layer0_outputs(5894));
    outputs(3228) <= not(layer0_outputs(7411));
    outputs(3229) <= not(layer0_outputs(3481));
    outputs(3230) <= not(layer0_outputs(3443)) or (layer0_outputs(2896));
    outputs(3231) <= not(layer0_outputs(4002)) or (layer0_outputs(2353));
    outputs(3232) <= layer0_outputs(2708);
    outputs(3233) <= (layer0_outputs(7632)) and not (layer0_outputs(10060));
    outputs(3234) <= (layer0_outputs(8245)) and not (layer0_outputs(2501));
    outputs(3235) <= (layer0_outputs(9536)) xor (layer0_outputs(10212));
    outputs(3236) <= layer0_outputs(2258);
    outputs(3237) <= (layer0_outputs(720)) xor (layer0_outputs(9491));
    outputs(3238) <= not(layer0_outputs(4513));
    outputs(3239) <= (layer0_outputs(2762)) and not (layer0_outputs(4704));
    outputs(3240) <= layer0_outputs(8216);
    outputs(3241) <= layer0_outputs(4577);
    outputs(3242) <= layer0_outputs(7729);
    outputs(3243) <= not(layer0_outputs(8591));
    outputs(3244) <= (layer0_outputs(5312)) xor (layer0_outputs(6735));
    outputs(3245) <= layer0_outputs(8982);
    outputs(3246) <= not(layer0_outputs(8285));
    outputs(3247) <= not(layer0_outputs(9285));
    outputs(3248) <= (layer0_outputs(8738)) and not (layer0_outputs(7424));
    outputs(3249) <= (layer0_outputs(1719)) and not (layer0_outputs(3873));
    outputs(3250) <= layer0_outputs(3943);
    outputs(3251) <= not((layer0_outputs(5950)) and (layer0_outputs(6296)));
    outputs(3252) <= not((layer0_outputs(7394)) or (layer0_outputs(656)));
    outputs(3253) <= not(layer0_outputs(9471));
    outputs(3254) <= (layer0_outputs(2081)) and not (layer0_outputs(4393));
    outputs(3255) <= not((layer0_outputs(1773)) xor (layer0_outputs(5364)));
    outputs(3256) <= (layer0_outputs(778)) and not (layer0_outputs(4037));
    outputs(3257) <= not((layer0_outputs(3508)) xor (layer0_outputs(1074)));
    outputs(3258) <= layer0_outputs(4831);
    outputs(3259) <= not(layer0_outputs(6257));
    outputs(3260) <= layer0_outputs(1158);
    outputs(3261) <= layer0_outputs(7846);
    outputs(3262) <= not((layer0_outputs(342)) xor (layer0_outputs(3072)));
    outputs(3263) <= not((layer0_outputs(8340)) xor (layer0_outputs(10148)));
    outputs(3264) <= not((layer0_outputs(6698)) xor (layer0_outputs(1942)));
    outputs(3265) <= layer0_outputs(3902);
    outputs(3266) <= (layer0_outputs(2971)) xor (layer0_outputs(3538));
    outputs(3267) <= not(layer0_outputs(2838));
    outputs(3268) <= layer0_outputs(1245);
    outputs(3269) <= not(layer0_outputs(5758));
    outputs(3270) <= (layer0_outputs(5452)) and not (layer0_outputs(7141));
    outputs(3271) <= not(layer0_outputs(4777));
    outputs(3272) <= (layer0_outputs(42)) and not (layer0_outputs(8685));
    outputs(3273) <= layer0_outputs(1798);
    outputs(3274) <= not(layer0_outputs(293)) or (layer0_outputs(9990));
    outputs(3275) <= (layer0_outputs(4174)) and (layer0_outputs(10226));
    outputs(3276) <= not((layer0_outputs(1991)) xor (layer0_outputs(4581)));
    outputs(3277) <= (layer0_outputs(3242)) or (layer0_outputs(1387));
    outputs(3278) <= layer0_outputs(8372);
    outputs(3279) <= layer0_outputs(4814);
    outputs(3280) <= not((layer0_outputs(5706)) or (layer0_outputs(7094)));
    outputs(3281) <= not(layer0_outputs(491));
    outputs(3282) <= not((layer0_outputs(8393)) xor (layer0_outputs(538)));
    outputs(3283) <= not(layer0_outputs(5247));
    outputs(3284) <= not(layer0_outputs(3065));
    outputs(3285) <= not(layer0_outputs(1970));
    outputs(3286) <= not(layer0_outputs(1446));
    outputs(3287) <= not((layer0_outputs(6665)) xor (layer0_outputs(2021)));
    outputs(3288) <= not((layer0_outputs(335)) xor (layer0_outputs(1001)));
    outputs(3289) <= not((layer0_outputs(1045)) and (layer0_outputs(8720)));
    outputs(3290) <= layer0_outputs(1420);
    outputs(3291) <= (layer0_outputs(6230)) and (layer0_outputs(2615));
    outputs(3292) <= layer0_outputs(3527);
    outputs(3293) <= layer0_outputs(4495);
    outputs(3294) <= not((layer0_outputs(8728)) or (layer0_outputs(6301)));
    outputs(3295) <= not(layer0_outputs(1736));
    outputs(3296) <= layer0_outputs(10075);
    outputs(3297) <= not((layer0_outputs(3311)) or (layer0_outputs(10138)));
    outputs(3298) <= layer0_outputs(9360);
    outputs(3299) <= (layer0_outputs(3710)) and (layer0_outputs(942));
    outputs(3300) <= not((layer0_outputs(9655)) or (layer0_outputs(8200)));
    outputs(3301) <= layer0_outputs(3444);
    outputs(3302) <= (layer0_outputs(8331)) xor (layer0_outputs(4998));
    outputs(3303) <= not(layer0_outputs(5297));
    outputs(3304) <= not(layer0_outputs(9181));
    outputs(3305) <= not((layer0_outputs(4462)) and (layer0_outputs(8032)));
    outputs(3306) <= (layer0_outputs(122)) xor (layer0_outputs(1950));
    outputs(3307) <= (layer0_outputs(7492)) and not (layer0_outputs(3009));
    outputs(3308) <= (layer0_outputs(150)) xor (layer0_outputs(9813));
    outputs(3309) <= (layer0_outputs(3853)) and not (layer0_outputs(5715));
    outputs(3310) <= not(layer0_outputs(8932));
    outputs(3311) <= layer0_outputs(2057);
    outputs(3312) <= layer0_outputs(4167);
    outputs(3313) <= not((layer0_outputs(1852)) or (layer0_outputs(5910)));
    outputs(3314) <= (layer0_outputs(1803)) and (layer0_outputs(2555));
    outputs(3315) <= not((layer0_outputs(4182)) xor (layer0_outputs(3611)));
    outputs(3316) <= (layer0_outputs(9818)) xor (layer0_outputs(5749));
    outputs(3317) <= layer0_outputs(4424);
    outputs(3318) <= not(layer0_outputs(2189));
    outputs(3319) <= layer0_outputs(6528);
    outputs(3320) <= not(layer0_outputs(4553));
    outputs(3321) <= (layer0_outputs(9352)) and not (layer0_outputs(4151));
    outputs(3322) <= not(layer0_outputs(8869));
    outputs(3323) <= layer0_outputs(9888);
    outputs(3324) <= layer0_outputs(3501);
    outputs(3325) <= '0';
    outputs(3326) <= (layer0_outputs(1824)) and not (layer0_outputs(8783));
    outputs(3327) <= layer0_outputs(6543);
    outputs(3328) <= not(layer0_outputs(10137));
    outputs(3329) <= not(layer0_outputs(8872));
    outputs(3330) <= layer0_outputs(2591);
    outputs(3331) <= (layer0_outputs(3492)) and not (layer0_outputs(2052));
    outputs(3332) <= not(layer0_outputs(8796));
    outputs(3333) <= layer0_outputs(5330);
    outputs(3334) <= not((layer0_outputs(7220)) xor (layer0_outputs(6927)));
    outputs(3335) <= not((layer0_outputs(1120)) xor (layer0_outputs(2387)));
    outputs(3336) <= not(layer0_outputs(94));
    outputs(3337) <= not((layer0_outputs(8273)) or (layer0_outputs(5874)));
    outputs(3338) <= layer0_outputs(6314);
    outputs(3339) <= (layer0_outputs(6995)) or (layer0_outputs(6342));
    outputs(3340) <= layer0_outputs(10114);
    outputs(3341) <= layer0_outputs(832);
    outputs(3342) <= not(layer0_outputs(7023));
    outputs(3343) <= not(layer0_outputs(4378));
    outputs(3344) <= layer0_outputs(129);
    outputs(3345) <= not(layer0_outputs(60)) or (layer0_outputs(9568));
    outputs(3346) <= not(layer0_outputs(3365));
    outputs(3347) <= not(layer0_outputs(3375)) or (layer0_outputs(7466));
    outputs(3348) <= layer0_outputs(4338);
    outputs(3349) <= not(layer0_outputs(3583));
    outputs(3350) <= (layer0_outputs(6496)) xor (layer0_outputs(3498));
    outputs(3351) <= not(layer0_outputs(900));
    outputs(3352) <= not((layer0_outputs(3577)) or (layer0_outputs(3723)));
    outputs(3353) <= not(layer0_outputs(6551)) or (layer0_outputs(6061));
    outputs(3354) <= not(layer0_outputs(163));
    outputs(3355) <= layer0_outputs(2328);
    outputs(3356) <= layer0_outputs(7015);
    outputs(3357) <= not(layer0_outputs(3015));
    outputs(3358) <= (layer0_outputs(2275)) or (layer0_outputs(7026));
    outputs(3359) <= not(layer0_outputs(2945));
    outputs(3360) <= (layer0_outputs(1149)) xor (layer0_outputs(1926));
    outputs(3361) <= (layer0_outputs(1031)) and (layer0_outputs(4940));
    outputs(3362) <= layer0_outputs(9199);
    outputs(3363) <= not(layer0_outputs(8506)) or (layer0_outputs(7033));
    outputs(3364) <= layer0_outputs(1592);
    outputs(3365) <= layer0_outputs(2636);
    outputs(3366) <= layer0_outputs(9715);
    outputs(3367) <= layer0_outputs(5281);
    outputs(3368) <= not(layer0_outputs(6553));
    outputs(3369) <= layer0_outputs(2667);
    outputs(3370) <= layer0_outputs(4941);
    outputs(3371) <= layer0_outputs(320);
    outputs(3372) <= not((layer0_outputs(6054)) xor (layer0_outputs(3150)));
    outputs(3373) <= (layer0_outputs(6556)) and not (layer0_outputs(4544));
    outputs(3374) <= (layer0_outputs(2153)) and (layer0_outputs(9848));
    outputs(3375) <= not(layer0_outputs(9007));
    outputs(3376) <= not((layer0_outputs(5257)) xor (layer0_outputs(4860)));
    outputs(3377) <= layer0_outputs(8735);
    outputs(3378) <= layer0_outputs(476);
    outputs(3379) <= not(layer0_outputs(1737));
    outputs(3380) <= not((layer0_outputs(5831)) xor (layer0_outputs(3308)));
    outputs(3381) <= layer0_outputs(9235);
    outputs(3382) <= not(layer0_outputs(6006));
    outputs(3383) <= not(layer0_outputs(8943));
    outputs(3384) <= layer0_outputs(2679);
    outputs(3385) <= not(layer0_outputs(459));
    outputs(3386) <= layer0_outputs(8144);
    outputs(3387) <= not(layer0_outputs(8226));
    outputs(3388) <= (layer0_outputs(3029)) and (layer0_outputs(8227));
    outputs(3389) <= not(layer0_outputs(5384));
    outputs(3390) <= not(layer0_outputs(6617));
    outputs(3391) <= layer0_outputs(4293);
    outputs(3392) <= not((layer0_outputs(677)) xor (layer0_outputs(4657)));
    outputs(3393) <= not((layer0_outputs(735)) and (layer0_outputs(5190)));
    outputs(3394) <= layer0_outputs(1949);
    outputs(3395) <= not(layer0_outputs(8590));
    outputs(3396) <= (layer0_outputs(7407)) or (layer0_outputs(3007));
    outputs(3397) <= (layer0_outputs(1082)) xor (layer0_outputs(6547));
    outputs(3398) <= not((layer0_outputs(2950)) xor (layer0_outputs(262)));
    outputs(3399) <= not(layer0_outputs(1149)) or (layer0_outputs(2355));
    outputs(3400) <= not(layer0_outputs(7396));
    outputs(3401) <= layer0_outputs(9274);
    outputs(3402) <= (layer0_outputs(8992)) and not (layer0_outputs(6974));
    outputs(3403) <= not(layer0_outputs(10203));
    outputs(3404) <= (layer0_outputs(8579)) and not (layer0_outputs(9931));
    outputs(3405) <= not((layer0_outputs(3026)) or (layer0_outputs(5973)));
    outputs(3406) <= layer0_outputs(4699);
    outputs(3407) <= layer0_outputs(5047);
    outputs(3408) <= not((layer0_outputs(6694)) and (layer0_outputs(4272)));
    outputs(3409) <= not(layer0_outputs(6190));
    outputs(3410) <= layer0_outputs(8404);
    outputs(3411) <= (layer0_outputs(6834)) xor (layer0_outputs(9971));
    outputs(3412) <= not(layer0_outputs(6000));
    outputs(3413) <= not(layer0_outputs(8592));
    outputs(3414) <= not(layer0_outputs(9722));
    outputs(3415) <= not(layer0_outputs(4094));
    outputs(3416) <= layer0_outputs(10150);
    outputs(3417) <= not(layer0_outputs(9225));
    outputs(3418) <= layer0_outputs(8475);
    outputs(3419) <= not(layer0_outputs(2287));
    outputs(3420) <= not((layer0_outputs(4822)) xor (layer0_outputs(1947)));
    outputs(3421) <= layer0_outputs(3128);
    outputs(3422) <= (layer0_outputs(4803)) and not (layer0_outputs(8059));
    outputs(3423) <= not(layer0_outputs(9193));
    outputs(3424) <= layer0_outputs(4264);
    outputs(3425) <= (layer0_outputs(6359)) and not (layer0_outputs(5805));
    outputs(3426) <= not(layer0_outputs(101));
    outputs(3427) <= layer0_outputs(3426);
    outputs(3428) <= (layer0_outputs(1667)) xor (layer0_outputs(9095));
    outputs(3429) <= not(layer0_outputs(7272));
    outputs(3430) <= not(layer0_outputs(5440));
    outputs(3431) <= layer0_outputs(2955);
    outputs(3432) <= layer0_outputs(9480);
    outputs(3433) <= not(layer0_outputs(9767));
    outputs(3434) <= (layer0_outputs(4391)) and not (layer0_outputs(3515));
    outputs(3435) <= layer0_outputs(8670);
    outputs(3436) <= not(layer0_outputs(7133));
    outputs(3437) <= layer0_outputs(9053);
    outputs(3438) <= (layer0_outputs(4594)) and not (layer0_outputs(596));
    outputs(3439) <= not(layer0_outputs(6611));
    outputs(3440) <= not((layer0_outputs(8881)) xor (layer0_outputs(8979)));
    outputs(3441) <= layer0_outputs(6776);
    outputs(3442) <= (layer0_outputs(2827)) xor (layer0_outputs(309));
    outputs(3443) <= not((layer0_outputs(2578)) xor (layer0_outputs(2506)));
    outputs(3444) <= layer0_outputs(3736);
    outputs(3445) <= not((layer0_outputs(2012)) and (layer0_outputs(8803)));
    outputs(3446) <= not(layer0_outputs(6247)) or (layer0_outputs(4656));
    outputs(3447) <= layer0_outputs(8787);
    outputs(3448) <= not(layer0_outputs(8295));
    outputs(3449) <= not(layer0_outputs(5683));
    outputs(3450) <= not(layer0_outputs(8816));
    outputs(3451) <= (layer0_outputs(7360)) xor (layer0_outputs(682));
    outputs(3452) <= (layer0_outputs(6943)) and not (layer0_outputs(100));
    outputs(3453) <= layer0_outputs(6980);
    outputs(3454) <= not((layer0_outputs(4344)) xor (layer0_outputs(8854)));
    outputs(3455) <= layer0_outputs(7289);
    outputs(3456) <= not(layer0_outputs(6106));
    outputs(3457) <= not(layer0_outputs(491));
    outputs(3458) <= not(layer0_outputs(2931));
    outputs(3459) <= not(layer0_outputs(7050));
    outputs(3460) <= layer0_outputs(5338);
    outputs(3461) <= not(layer0_outputs(1941));
    outputs(3462) <= layer0_outputs(664);
    outputs(3463) <= not(layer0_outputs(3216)) or (layer0_outputs(8653));
    outputs(3464) <= (layer0_outputs(9745)) and not (layer0_outputs(764));
    outputs(3465) <= (layer0_outputs(6253)) xor (layer0_outputs(676));
    outputs(3466) <= (layer0_outputs(6370)) and (layer0_outputs(8703));
    outputs(3467) <= not(layer0_outputs(7546)) or (layer0_outputs(4296));
    outputs(3468) <= not(layer0_outputs(8463));
    outputs(3469) <= layer0_outputs(3332);
    outputs(3470) <= layer0_outputs(3985);
    outputs(3471) <= not((layer0_outputs(347)) xor (layer0_outputs(1374)));
    outputs(3472) <= not((layer0_outputs(9539)) xor (layer0_outputs(1820)));
    outputs(3473) <= (layer0_outputs(5434)) xor (layer0_outputs(2440));
    outputs(3474) <= (layer0_outputs(8196)) and (layer0_outputs(9710));
    outputs(3475) <= (layer0_outputs(3110)) or (layer0_outputs(4174));
    outputs(3476) <= not((layer0_outputs(1443)) xor (layer0_outputs(34)));
    outputs(3477) <= layer0_outputs(5339);
    outputs(3478) <= not((layer0_outputs(3964)) or (layer0_outputs(1229)));
    outputs(3479) <= (layer0_outputs(8277)) and not (layer0_outputs(283));
    outputs(3480) <= (layer0_outputs(4614)) xor (layer0_outputs(6207));
    outputs(3481) <= not(layer0_outputs(3075));
    outputs(3482) <= not(layer0_outputs(1032));
    outputs(3483) <= (layer0_outputs(9906)) and (layer0_outputs(5614));
    outputs(3484) <= (layer0_outputs(716)) and not (layer0_outputs(3748));
    outputs(3485) <= not(layer0_outputs(1238)) or (layer0_outputs(7783));
    outputs(3486) <= layer0_outputs(9735);
    outputs(3487) <= not(layer0_outputs(8052)) or (layer0_outputs(1793));
    outputs(3488) <= layer0_outputs(7755);
    outputs(3489) <= layer0_outputs(1404);
    outputs(3490) <= (layer0_outputs(417)) xor (layer0_outputs(8588));
    outputs(3491) <= not(layer0_outputs(4306)) or (layer0_outputs(7079));
    outputs(3492) <= layer0_outputs(7682);
    outputs(3493) <= not(layer0_outputs(1962));
    outputs(3494) <= layer0_outputs(1937);
    outputs(3495) <= not(layer0_outputs(1506)) or (layer0_outputs(8473));
    outputs(3496) <= not(layer0_outputs(5969));
    outputs(3497) <= layer0_outputs(432);
    outputs(3498) <= layer0_outputs(4134);
    outputs(3499) <= not((layer0_outputs(2996)) or (layer0_outputs(5740)));
    outputs(3500) <= layer0_outputs(5812);
    outputs(3501) <= layer0_outputs(396);
    outputs(3502) <= not(layer0_outputs(377));
    outputs(3503) <= layer0_outputs(6493);
    outputs(3504) <= not(layer0_outputs(8545));
    outputs(3505) <= layer0_outputs(10130);
    outputs(3506) <= layer0_outputs(6171);
    outputs(3507) <= layer0_outputs(3036);
    outputs(3508) <= (layer0_outputs(3306)) and not (layer0_outputs(7988));
    outputs(3509) <= (layer0_outputs(1374)) xor (layer0_outputs(2452));
    outputs(3510) <= not(layer0_outputs(163));
    outputs(3511) <= not(layer0_outputs(4895));
    outputs(3512) <= not((layer0_outputs(2512)) xor (layer0_outputs(8778)));
    outputs(3513) <= layer0_outputs(3965);
    outputs(3514) <= not(layer0_outputs(8173));
    outputs(3515) <= layer0_outputs(9581);
    outputs(3516) <= (layer0_outputs(2733)) xor (layer0_outputs(3370));
    outputs(3517) <= not(layer0_outputs(7199));
    outputs(3518) <= (layer0_outputs(3468)) and (layer0_outputs(6871));
    outputs(3519) <= layer0_outputs(4487);
    outputs(3520) <= not((layer0_outputs(9159)) xor (layer0_outputs(4033)));
    outputs(3521) <= not((layer0_outputs(26)) or (layer0_outputs(5551)));
    outputs(3522) <= not(layer0_outputs(3770));
    outputs(3523) <= (layer0_outputs(6598)) or (layer0_outputs(5016));
    outputs(3524) <= (layer0_outputs(1118)) and not (layer0_outputs(5143));
    outputs(3525) <= not(layer0_outputs(4318));
    outputs(3526) <= layer0_outputs(6280);
    outputs(3527) <= not(layer0_outputs(8695));
    outputs(3528) <= (layer0_outputs(5388)) xor (layer0_outputs(896));
    outputs(3529) <= (layer0_outputs(6491)) and not (layer0_outputs(8330));
    outputs(3530) <= layer0_outputs(1011);
    outputs(3531) <= layer0_outputs(1602);
    outputs(3532) <= (layer0_outputs(7282)) xor (layer0_outputs(8748));
    outputs(3533) <= not((layer0_outputs(8340)) or (layer0_outputs(8696)));
    outputs(3534) <= not((layer0_outputs(3716)) xor (layer0_outputs(3786)));
    outputs(3535) <= not((layer0_outputs(112)) xor (layer0_outputs(7491)));
    outputs(3536) <= layer0_outputs(795);
    outputs(3537) <= layer0_outputs(1289);
    outputs(3538) <= layer0_outputs(2880);
    outputs(3539) <= layer0_outputs(2633);
    outputs(3540) <= (layer0_outputs(4156)) xor (layer0_outputs(1940));
    outputs(3541) <= (layer0_outputs(8983)) and not (layer0_outputs(1102));
    outputs(3542) <= not(layer0_outputs(7239));
    outputs(3543) <= (layer0_outputs(7071)) and not (layer0_outputs(2078));
    outputs(3544) <= (layer0_outputs(9826)) xor (layer0_outputs(4108));
    outputs(3545) <= not((layer0_outputs(5022)) xor (layer0_outputs(8804)));
    outputs(3546) <= not(layer0_outputs(2692));
    outputs(3547) <= not(layer0_outputs(1851));
    outputs(3548) <= not(layer0_outputs(7041));
    outputs(3549) <= (layer0_outputs(3121)) and not (layer0_outputs(7663));
    outputs(3550) <= not(layer0_outputs(2229));
    outputs(3551) <= not(layer0_outputs(5780));
    outputs(3552) <= (layer0_outputs(9831)) xor (layer0_outputs(8140));
    outputs(3553) <= (layer0_outputs(9667)) xor (layer0_outputs(225));
    outputs(3554) <= not(layer0_outputs(7710)) or (layer0_outputs(2665));
    outputs(3555) <= (layer0_outputs(2589)) and not (layer0_outputs(4185));
    outputs(3556) <= not(layer0_outputs(1393));
    outputs(3557) <= (layer0_outputs(6406)) xor (layer0_outputs(8696));
    outputs(3558) <= '1';
    outputs(3559) <= (layer0_outputs(10199)) and not (layer0_outputs(3731));
    outputs(3560) <= (layer0_outputs(44)) xor (layer0_outputs(7939));
    outputs(3561) <= not(layer0_outputs(5142));
    outputs(3562) <= not((layer0_outputs(6026)) xor (layer0_outputs(5966)));
    outputs(3563) <= not(layer0_outputs(1509));
    outputs(3564) <= (layer0_outputs(9871)) and (layer0_outputs(9937));
    outputs(3565) <= layer0_outputs(1515);
    outputs(3566) <= not(layer0_outputs(2366));
    outputs(3567) <= layer0_outputs(8372);
    outputs(3568) <= layer0_outputs(8303);
    outputs(3569) <= not((layer0_outputs(6358)) and (layer0_outputs(1899)));
    outputs(3570) <= not(layer0_outputs(1308));
    outputs(3571) <= not(layer0_outputs(4758));
    outputs(3572) <= not(layer0_outputs(8314)) or (layer0_outputs(2674));
    outputs(3573) <= layer0_outputs(2630);
    outputs(3574) <= layer0_outputs(8058);
    outputs(3575) <= (layer0_outputs(7889)) and not (layer0_outputs(3603));
    outputs(3576) <= layer0_outputs(10150);
    outputs(3577) <= (layer0_outputs(5276)) xor (layer0_outputs(2669));
    outputs(3578) <= layer0_outputs(782);
    outputs(3579) <= (layer0_outputs(7803)) and not (layer0_outputs(5906));
    outputs(3580) <= not(layer0_outputs(457));
    outputs(3581) <= (layer0_outputs(2758)) and (layer0_outputs(6950));
    outputs(3582) <= (layer0_outputs(7198)) and (layer0_outputs(4992));
    outputs(3583) <= not((layer0_outputs(8526)) xor (layer0_outputs(6706)));
    outputs(3584) <= not(layer0_outputs(5609));
    outputs(3585) <= not(layer0_outputs(9071));
    outputs(3586) <= not(layer0_outputs(7161));
    outputs(3587) <= layer0_outputs(7829);
    outputs(3588) <= layer0_outputs(7657);
    outputs(3589) <= not(layer0_outputs(7875));
    outputs(3590) <= not((layer0_outputs(4591)) and (layer0_outputs(6096)));
    outputs(3591) <= not(layer0_outputs(4081)) or (layer0_outputs(6627));
    outputs(3592) <= layer0_outputs(4596);
    outputs(3593) <= layer0_outputs(4139);
    outputs(3594) <= not(layer0_outputs(2753));
    outputs(3595) <= not((layer0_outputs(5003)) and (layer0_outputs(3538)));
    outputs(3596) <= not(layer0_outputs(1634));
    outputs(3597) <= (layer0_outputs(8955)) or (layer0_outputs(1224));
    outputs(3598) <= (layer0_outputs(7809)) and not (layer0_outputs(7312));
    outputs(3599) <= not(layer0_outputs(9558));
    outputs(3600) <= not((layer0_outputs(7610)) xor (layer0_outputs(5289)));
    outputs(3601) <= not(layer0_outputs(8429)) or (layer0_outputs(7129));
    outputs(3602) <= not((layer0_outputs(8792)) or (layer0_outputs(8581)));
    outputs(3603) <= not((layer0_outputs(1065)) xor (layer0_outputs(9321)));
    outputs(3604) <= (layer0_outputs(3244)) xor (layer0_outputs(4379));
    outputs(3605) <= not((layer0_outputs(738)) xor (layer0_outputs(1677)));
    outputs(3606) <= (layer0_outputs(4479)) or (layer0_outputs(1197));
    outputs(3607) <= layer0_outputs(6168);
    outputs(3608) <= (layer0_outputs(4938)) and not (layer0_outputs(1961));
    outputs(3609) <= (layer0_outputs(3657)) xor (layer0_outputs(6362));
    outputs(3610) <= not(layer0_outputs(977));
    outputs(3611) <= layer0_outputs(5442);
    outputs(3612) <= not(layer0_outputs(3669));
    outputs(3613) <= layer0_outputs(3135);
    outputs(3614) <= not(layer0_outputs(6378));
    outputs(3615) <= not(layer0_outputs(8613));
    outputs(3616) <= layer0_outputs(364);
    outputs(3617) <= not(layer0_outputs(8067));
    outputs(3618) <= not(layer0_outputs(6068));
    outputs(3619) <= layer0_outputs(6180);
    outputs(3620) <= (layer0_outputs(5686)) xor (layer0_outputs(6514));
    outputs(3621) <= not((layer0_outputs(3334)) xor (layer0_outputs(1069)));
    outputs(3622) <= layer0_outputs(1161);
    outputs(3623) <= not((layer0_outputs(1048)) or (layer0_outputs(3287)));
    outputs(3624) <= not(layer0_outputs(7511));
    outputs(3625) <= not(layer0_outputs(10033));
    outputs(3626) <= (layer0_outputs(7673)) and (layer0_outputs(5536));
    outputs(3627) <= (layer0_outputs(7738)) xor (layer0_outputs(3913));
    outputs(3628) <= not(layer0_outputs(7193));
    outputs(3629) <= layer0_outputs(4215);
    outputs(3630) <= (layer0_outputs(4091)) xor (layer0_outputs(5315));
    outputs(3631) <= not((layer0_outputs(4843)) and (layer0_outputs(6666)));
    outputs(3632) <= not(layer0_outputs(3951));
    outputs(3633) <= (layer0_outputs(7748)) and (layer0_outputs(6078));
    outputs(3634) <= not(layer0_outputs(4286));
    outputs(3635) <= layer0_outputs(6655);
    outputs(3636) <= layer0_outputs(6127);
    outputs(3637) <= not(layer0_outputs(7253));
    outputs(3638) <= layer0_outputs(1894);
    outputs(3639) <= (layer0_outputs(4497)) and not (layer0_outputs(1400));
    outputs(3640) <= (layer0_outputs(3888)) and (layer0_outputs(7603));
    outputs(3641) <= layer0_outputs(743);
    outputs(3642) <= not(layer0_outputs(1029)) or (layer0_outputs(4624));
    outputs(3643) <= (layer0_outputs(3776)) or (layer0_outputs(7468));
    outputs(3644) <= (layer0_outputs(4163)) xor (layer0_outputs(8225));
    outputs(3645) <= layer0_outputs(6388);
    outputs(3646) <= layer0_outputs(9927);
    outputs(3647) <= not(layer0_outputs(429));
    outputs(3648) <= layer0_outputs(3729);
    outputs(3649) <= not((layer0_outputs(8782)) xor (layer0_outputs(901)));
    outputs(3650) <= layer0_outputs(6693);
    outputs(3651) <= (layer0_outputs(6819)) xor (layer0_outputs(6726));
    outputs(3652) <= (layer0_outputs(6093)) and (layer0_outputs(8479));
    outputs(3653) <= not((layer0_outputs(3999)) xor (layer0_outputs(1250)));
    outputs(3654) <= (layer0_outputs(5615)) and (layer0_outputs(2597));
    outputs(3655) <= layer0_outputs(2722);
    outputs(3656) <= layer0_outputs(1919);
    outputs(3657) <= not((layer0_outputs(7936)) xor (layer0_outputs(4557)));
    outputs(3658) <= (layer0_outputs(9808)) and not (layer0_outputs(2587));
    outputs(3659) <= not(layer0_outputs(6763));
    outputs(3660) <= not((layer0_outputs(773)) xor (layer0_outputs(6483)));
    outputs(3661) <= layer0_outputs(1590);
    outputs(3662) <= not(layer0_outputs(899)) or (layer0_outputs(5972));
    outputs(3663) <= (layer0_outputs(3774)) xor (layer0_outputs(4534));
    outputs(3664) <= (layer0_outputs(8622)) and not (layer0_outputs(6612));
    outputs(3665) <= layer0_outputs(6594);
    outputs(3666) <= not((layer0_outputs(8274)) xor (layer0_outputs(5163)));
    outputs(3667) <= not((layer0_outputs(578)) and (layer0_outputs(4054)));
    outputs(3668) <= not(layer0_outputs(5181));
    outputs(3669) <= layer0_outputs(8062);
    outputs(3670) <= not(layer0_outputs(8239));
    outputs(3671) <= (layer0_outputs(4494)) and (layer0_outputs(9446));
    outputs(3672) <= not(layer0_outputs(6442));
    outputs(3673) <= not(layer0_outputs(10220));
    outputs(3674) <= not((layer0_outputs(6947)) xor (layer0_outputs(7566)));
    outputs(3675) <= not((layer0_outputs(5635)) or (layer0_outputs(10093)));
    outputs(3676) <= (layer0_outputs(8474)) and not (layer0_outputs(1737));
    outputs(3677) <= (layer0_outputs(6930)) and not (layer0_outputs(9753));
    outputs(3678) <= (layer0_outputs(2919)) and not (layer0_outputs(3282));
    outputs(3679) <= not((layer0_outputs(1061)) and (layer0_outputs(1253)));
    outputs(3680) <= not(layer0_outputs(4025));
    outputs(3681) <= not(layer0_outputs(4630));
    outputs(3682) <= not(layer0_outputs(9998)) or (layer0_outputs(149));
    outputs(3683) <= layer0_outputs(5856);
    outputs(3684) <= not(layer0_outputs(8445));
    outputs(3685) <= (layer0_outputs(4198)) xor (layer0_outputs(4207));
    outputs(3686) <= layer0_outputs(9405);
    outputs(3687) <= (layer0_outputs(894)) and not (layer0_outputs(623));
    outputs(3688) <= not(layer0_outputs(9707));
    outputs(3689) <= not((layer0_outputs(1097)) xor (layer0_outputs(4160)));
    outputs(3690) <= not((layer0_outputs(1031)) xor (layer0_outputs(4733)));
    outputs(3691) <= (layer0_outputs(3187)) xor (layer0_outputs(1229));
    outputs(3692) <= not(layer0_outputs(4741)) or (layer0_outputs(8861));
    outputs(3693) <= layer0_outputs(7625);
    outputs(3694) <= layer0_outputs(6552);
    outputs(3695) <= not(layer0_outputs(3262)) or (layer0_outputs(4475));
    outputs(3696) <= layer0_outputs(8327);
    outputs(3697) <= (layer0_outputs(6276)) xor (layer0_outputs(7095));
    outputs(3698) <= not(layer0_outputs(7662));
    outputs(3699) <= (layer0_outputs(7745)) and not (layer0_outputs(6351));
    outputs(3700) <= not((layer0_outputs(3433)) xor (layer0_outputs(8552)));
    outputs(3701) <= (layer0_outputs(9001)) and not (layer0_outputs(7016));
    outputs(3702) <= layer0_outputs(6753);
    outputs(3703) <= not(layer0_outputs(9042));
    outputs(3704) <= layer0_outputs(9239);
    outputs(3705) <= not((layer0_outputs(9489)) xor (layer0_outputs(8624)));
    outputs(3706) <= not(layer0_outputs(5203));
    outputs(3707) <= not(layer0_outputs(2474));
    outputs(3708) <= layer0_outputs(9113);
    outputs(3709) <= (layer0_outputs(4653)) xor (layer0_outputs(559));
    outputs(3710) <= not((layer0_outputs(4351)) xor (layer0_outputs(1543)));
    outputs(3711) <= (layer0_outputs(1340)) and not (layer0_outputs(6423));
    outputs(3712) <= not((layer0_outputs(4994)) xor (layer0_outputs(1123)));
    outputs(3713) <= not(layer0_outputs(8394));
    outputs(3714) <= not(layer0_outputs(1872));
    outputs(3715) <= layer0_outputs(2244);
    outputs(3716) <= not(layer0_outputs(5804));
    outputs(3717) <= not(layer0_outputs(7180)) or (layer0_outputs(4416));
    outputs(3718) <= layer0_outputs(8347);
    outputs(3719) <= not(layer0_outputs(5467));
    outputs(3720) <= not(layer0_outputs(4779));
    outputs(3721) <= layer0_outputs(5929);
    outputs(3722) <= layer0_outputs(8737);
    outputs(3723) <= not(layer0_outputs(4002));
    outputs(3724) <= (layer0_outputs(5030)) xor (layer0_outputs(4086));
    outputs(3725) <= not(layer0_outputs(6284));
    outputs(3726) <= not(layer0_outputs(480));
    outputs(3727) <= layer0_outputs(27);
    outputs(3728) <= layer0_outputs(1282);
    outputs(3729) <= layer0_outputs(1581);
    outputs(3730) <= (layer0_outputs(902)) and (layer0_outputs(8841));
    outputs(3731) <= not(layer0_outputs(7023));
    outputs(3732) <= (layer0_outputs(5515)) xor (layer0_outputs(7420));
    outputs(3733) <= layer0_outputs(6696);
    outputs(3734) <= (layer0_outputs(6385)) and not (layer0_outputs(38));
    outputs(3735) <= not(layer0_outputs(9129)) or (layer0_outputs(536));
    outputs(3736) <= (layer0_outputs(8667)) and not (layer0_outputs(3608));
    outputs(3737) <= layer0_outputs(748);
    outputs(3738) <= (layer0_outputs(10133)) and not (layer0_outputs(9271));
    outputs(3739) <= layer0_outputs(3410);
    outputs(3740) <= (layer0_outputs(7972)) and not (layer0_outputs(2088));
    outputs(3741) <= layer0_outputs(6055);
    outputs(3742) <= layer0_outputs(6603);
    outputs(3743) <= not((layer0_outputs(6304)) xor (layer0_outputs(8894)));
    outputs(3744) <= layer0_outputs(9618);
    outputs(3745) <= layer0_outputs(5711);
    outputs(3746) <= not(layer0_outputs(84));
    outputs(3747) <= not(layer0_outputs(4330));
    outputs(3748) <= (layer0_outputs(6419)) xor (layer0_outputs(1985));
    outputs(3749) <= not((layer0_outputs(9943)) or (layer0_outputs(1338)));
    outputs(3750) <= layer0_outputs(9578);
    outputs(3751) <= not((layer0_outputs(2010)) xor (layer0_outputs(8320)));
    outputs(3752) <= not(layer0_outputs(5486));
    outputs(3753) <= (layer0_outputs(5080)) and (layer0_outputs(3544));
    outputs(3754) <= not((layer0_outputs(7890)) and (layer0_outputs(5034)));
    outputs(3755) <= not((layer0_outputs(7479)) xor (layer0_outputs(4528)));
    outputs(3756) <= not(layer0_outputs(2658));
    outputs(3757) <= (layer0_outputs(5435)) xor (layer0_outputs(2725));
    outputs(3758) <= layer0_outputs(7085);
    outputs(3759) <= layer0_outputs(9469);
    outputs(3760) <= not((layer0_outputs(4748)) xor (layer0_outputs(5297)));
    outputs(3761) <= (layer0_outputs(5233)) xor (layer0_outputs(249));
    outputs(3762) <= layer0_outputs(1456);
    outputs(3763) <= (layer0_outputs(9335)) and not (layer0_outputs(5463));
    outputs(3764) <= layer0_outputs(9006);
    outputs(3765) <= (layer0_outputs(5873)) xor (layer0_outputs(6741));
    outputs(3766) <= layer0_outputs(10088);
    outputs(3767) <= layer0_outputs(2093);
    outputs(3768) <= not(layer0_outputs(3514)) or (layer0_outputs(7668));
    outputs(3769) <= not((layer0_outputs(8236)) xor (layer0_outputs(4892)));
    outputs(3770) <= not((layer0_outputs(3386)) and (layer0_outputs(2321)));
    outputs(3771) <= not(layer0_outputs(7202));
    outputs(3772) <= (layer0_outputs(5415)) or (layer0_outputs(62));
    outputs(3773) <= not(layer0_outputs(1416)) or (layer0_outputs(2645));
    outputs(3774) <= (layer0_outputs(413)) and (layer0_outputs(3099));
    outputs(3775) <= (layer0_outputs(632)) and (layer0_outputs(7603));
    outputs(3776) <= (layer0_outputs(8483)) xor (layer0_outputs(7955));
    outputs(3777) <= not((layer0_outputs(3396)) xor (layer0_outputs(1896)));
    outputs(3778) <= (layer0_outputs(3780)) and (layer0_outputs(9330));
    outputs(3779) <= not((layer0_outputs(8806)) xor (layer0_outputs(5583)));
    outputs(3780) <= not((layer0_outputs(8764)) xor (layer0_outputs(9739)));
    outputs(3781) <= (layer0_outputs(8027)) xor (layer0_outputs(7071));
    outputs(3782) <= not((layer0_outputs(7299)) and (layer0_outputs(2564)));
    outputs(3783) <= (layer0_outputs(5992)) xor (layer0_outputs(8116));
    outputs(3784) <= (layer0_outputs(1287)) and not (layer0_outputs(1643));
    outputs(3785) <= layer0_outputs(4353);
    outputs(3786) <= not(layer0_outputs(8368));
    outputs(3787) <= not(layer0_outputs(6809));
    outputs(3788) <= not((layer0_outputs(6124)) or (layer0_outputs(5309)));
    outputs(3789) <= (layer0_outputs(3861)) xor (layer0_outputs(1467));
    outputs(3790) <= (layer0_outputs(1866)) and not (layer0_outputs(9809));
    outputs(3791) <= not((layer0_outputs(4781)) and (layer0_outputs(9964)));
    outputs(3792) <= (layer0_outputs(9592)) and not (layer0_outputs(9225));
    outputs(3793) <= (layer0_outputs(295)) and (layer0_outputs(8348));
    outputs(3794) <= not((layer0_outputs(3208)) or (layer0_outputs(5216)));
    outputs(3795) <= layer0_outputs(4999);
    outputs(3796) <= (layer0_outputs(6015)) and not (layer0_outputs(3313));
    outputs(3797) <= (layer0_outputs(4153)) or (layer0_outputs(1724));
    outputs(3798) <= layer0_outputs(6918);
    outputs(3799) <= (layer0_outputs(5391)) and not (layer0_outputs(3418));
    outputs(3800) <= not(layer0_outputs(1336));
    outputs(3801) <= not((layer0_outputs(3304)) or (layer0_outputs(6888)));
    outputs(3802) <= layer0_outputs(7570);
    outputs(3803) <= layer0_outputs(934);
    outputs(3804) <= not(layer0_outputs(8549));
    outputs(3805) <= not((layer0_outputs(5746)) xor (layer0_outputs(4508)));
    outputs(3806) <= not(layer0_outputs(2468));
    outputs(3807) <= (layer0_outputs(10121)) and not (layer0_outputs(8616));
    outputs(3808) <= layer0_outputs(6969);
    outputs(3809) <= (layer0_outputs(9538)) xor (layer0_outputs(7670));
    outputs(3810) <= layer0_outputs(6875);
    outputs(3811) <= not((layer0_outputs(1796)) xor (layer0_outputs(7419)));
    outputs(3812) <= layer0_outputs(6883);
    outputs(3813) <= not((layer0_outputs(542)) xor (layer0_outputs(2741)));
    outputs(3814) <= (layer0_outputs(5622)) and not (layer0_outputs(1513));
    outputs(3815) <= (layer0_outputs(3470)) and (layer0_outputs(5785));
    outputs(3816) <= not(layer0_outputs(7984));
    outputs(3817) <= (layer0_outputs(6080)) and not (layer0_outputs(5591));
    outputs(3818) <= not(layer0_outputs(7746));
    outputs(3819) <= not((layer0_outputs(6458)) xor (layer0_outputs(3391)));
    outputs(3820) <= layer0_outputs(785);
    outputs(3821) <= (layer0_outputs(4840)) xor (layer0_outputs(3550));
    outputs(3822) <= layer0_outputs(224);
    outputs(3823) <= not(layer0_outputs(771));
    outputs(3824) <= layer0_outputs(7334);
    outputs(3825) <= not(layer0_outputs(8034));
    outputs(3826) <= not(layer0_outputs(1625));
    outputs(3827) <= not(layer0_outputs(5871));
    outputs(3828) <= layer0_outputs(9395);
    outputs(3829) <= layer0_outputs(5040);
    outputs(3830) <= (layer0_outputs(5775)) and (layer0_outputs(8081));
    outputs(3831) <= layer0_outputs(6767);
    outputs(3832) <= not(layer0_outputs(8305));
    outputs(3833) <= not(layer0_outputs(8686)) or (layer0_outputs(2811));
    outputs(3834) <= not((layer0_outputs(6362)) xor (layer0_outputs(6419)));
    outputs(3835) <= not((layer0_outputs(9582)) xor (layer0_outputs(8471)));
    outputs(3836) <= layer0_outputs(9786);
    outputs(3837) <= not((layer0_outputs(1867)) xor (layer0_outputs(4699)));
    outputs(3838) <= not((layer0_outputs(1794)) xor (layer0_outputs(4638)));
    outputs(3839) <= layer0_outputs(715);
    outputs(3840) <= not(layer0_outputs(3328));
    outputs(3841) <= not(layer0_outputs(8927));
    outputs(3842) <= layer0_outputs(3067);
    outputs(3843) <= not((layer0_outputs(6773)) or (layer0_outputs(551)));
    outputs(3844) <= not(layer0_outputs(2148)) or (layer0_outputs(5361));
    outputs(3845) <= (layer0_outputs(4875)) or (layer0_outputs(9023));
    outputs(3846) <= layer0_outputs(8505);
    outputs(3847) <= not(layer0_outputs(9010));
    outputs(3848) <= not((layer0_outputs(8171)) and (layer0_outputs(8535)));
    outputs(3849) <= not(layer0_outputs(1635));
    outputs(3850) <= (layer0_outputs(5422)) xor (layer0_outputs(3762));
    outputs(3851) <= layer0_outputs(8735);
    outputs(3852) <= not((layer0_outputs(5097)) xor (layer0_outputs(7655)));
    outputs(3853) <= not((layer0_outputs(883)) or (layer0_outputs(713)));
    outputs(3854) <= layer0_outputs(933);
    outputs(3855) <= not(layer0_outputs(2700));
    outputs(3856) <= layer0_outputs(8341);
    outputs(3857) <= layer0_outputs(7386);
    outputs(3858) <= not(layer0_outputs(3901));
    outputs(3859) <= not(layer0_outputs(4858));
    outputs(3860) <= not((layer0_outputs(547)) xor (layer0_outputs(4605)));
    outputs(3861) <= (layer0_outputs(8385)) xor (layer0_outputs(10052));
    outputs(3862) <= layer0_outputs(8012);
    outputs(3863) <= layer0_outputs(9221);
    outputs(3864) <= not(layer0_outputs(503));
    outputs(3865) <= (layer0_outputs(2268)) xor (layer0_outputs(7460));
    outputs(3866) <= (layer0_outputs(7156)) xor (layer0_outputs(5672));
    outputs(3867) <= (layer0_outputs(2182)) or (layer0_outputs(11));
    outputs(3868) <= not((layer0_outputs(8516)) or (layer0_outputs(1173)));
    outputs(3869) <= not(layer0_outputs(634));
    outputs(3870) <= layer0_outputs(88);
    outputs(3871) <= (layer0_outputs(8168)) xor (layer0_outputs(7708));
    outputs(3872) <= (layer0_outputs(7154)) or (layer0_outputs(8969));
    outputs(3873) <= (layer0_outputs(7352)) or (layer0_outputs(8986));
    outputs(3874) <= layer0_outputs(5374);
    outputs(3875) <= not(layer0_outputs(3834));
    outputs(3876) <= not(layer0_outputs(6710));
    outputs(3877) <= (layer0_outputs(5214)) and not (layer0_outputs(5556));
    outputs(3878) <= layer0_outputs(7885);
    outputs(3879) <= not((layer0_outputs(4685)) xor (layer0_outputs(5218)));
    outputs(3880) <= not((layer0_outputs(2334)) or (layer0_outputs(4275)));
    outputs(3881) <= not(layer0_outputs(8788));
    outputs(3882) <= layer0_outputs(4595);
    outputs(3883) <= not(layer0_outputs(8106)) or (layer0_outputs(2405));
    outputs(3884) <= not(layer0_outputs(3635));
    outputs(3885) <= not(layer0_outputs(3581));
    outputs(3886) <= not((layer0_outputs(9591)) xor (layer0_outputs(1343)));
    outputs(3887) <= not(layer0_outputs(9260)) or (layer0_outputs(4684));
    outputs(3888) <= layer0_outputs(908);
    outputs(3889) <= layer0_outputs(4890);
    outputs(3890) <= not(layer0_outputs(9738));
    outputs(3891) <= layer0_outputs(9978);
    outputs(3892) <= not(layer0_outputs(3894));
    outputs(3893) <= not(layer0_outputs(6109)) or (layer0_outputs(3147));
    outputs(3894) <= not(layer0_outputs(9706));
    outputs(3895) <= not(layer0_outputs(5959));
    outputs(3896) <= (layer0_outputs(4308)) xor (layer0_outputs(8660));
    outputs(3897) <= layer0_outputs(7637);
    outputs(3898) <= (layer0_outputs(4969)) xor (layer0_outputs(5198));
    outputs(3899) <= (layer0_outputs(507)) and not (layer0_outputs(4794));
    outputs(3900) <= layer0_outputs(6744);
    outputs(3901) <= (layer0_outputs(5926)) and not (layer0_outputs(7996));
    outputs(3902) <= layer0_outputs(4460);
    outputs(3903) <= (layer0_outputs(3692)) xor (layer0_outputs(1907));
    outputs(3904) <= (layer0_outputs(6238)) and not (layer0_outputs(7771));
    outputs(3905) <= not(layer0_outputs(10073));
    outputs(3906) <= (layer0_outputs(6877)) xor (layer0_outputs(9616));
    outputs(3907) <= (layer0_outputs(2361)) xor (layer0_outputs(9526));
    outputs(3908) <= (layer0_outputs(345)) or (layer0_outputs(1202));
    outputs(3909) <= layer0_outputs(5523);
    outputs(3910) <= (layer0_outputs(7227)) and not (layer0_outputs(8699));
    outputs(3911) <= (layer0_outputs(8776)) xor (layer0_outputs(6505));
    outputs(3912) <= not(layer0_outputs(8318));
    outputs(3913) <= layer0_outputs(2913);
    outputs(3914) <= layer0_outputs(107);
    outputs(3915) <= (layer0_outputs(9911)) xor (layer0_outputs(6458));
    outputs(3916) <= layer0_outputs(1799);
    outputs(3917) <= not(layer0_outputs(8210));
    outputs(3918) <= layer0_outputs(374);
    outputs(3919) <= (layer0_outputs(6379)) xor (layer0_outputs(7256));
    outputs(3920) <= not((layer0_outputs(5483)) xor (layer0_outputs(6915)));
    outputs(3921) <= (layer0_outputs(444)) xor (layer0_outputs(5177));
    outputs(3922) <= not((layer0_outputs(7358)) xor (layer0_outputs(2791)));
    outputs(3923) <= (layer0_outputs(199)) and not (layer0_outputs(7391));
    outputs(3924) <= (layer0_outputs(7775)) and not (layer0_outputs(3407));
    outputs(3925) <= (layer0_outputs(835)) xor (layer0_outputs(9513));
    outputs(3926) <= not(layer0_outputs(9828));
    outputs(3927) <= (layer0_outputs(5484)) and not (layer0_outputs(3777));
    outputs(3928) <= not(layer0_outputs(1834));
    outputs(3929) <= layer0_outputs(3918);
    outputs(3930) <= not(layer0_outputs(5792));
    outputs(3931) <= (layer0_outputs(3990)) xor (layer0_outputs(5114));
    outputs(3932) <= layer0_outputs(7896);
    outputs(3933) <= not(layer0_outputs(633));
    outputs(3934) <= (layer0_outputs(5016)) and (layer0_outputs(6510));
    outputs(3935) <= layer0_outputs(7342);
    outputs(3936) <= (layer0_outputs(1774)) and (layer0_outputs(4186));
    outputs(3937) <= layer0_outputs(6657);
    outputs(3938) <= not(layer0_outputs(9336));
    outputs(3939) <= (layer0_outputs(214)) and (layer0_outputs(7174));
    outputs(3940) <= not(layer0_outputs(1728)) or (layer0_outputs(530));
    outputs(3941) <= layer0_outputs(4290);
    outputs(3942) <= (layer0_outputs(9771)) xor (layer0_outputs(3365));
    outputs(3943) <= not(layer0_outputs(4502));
    outputs(3944) <= not(layer0_outputs(2629));
    outputs(3945) <= not((layer0_outputs(5628)) xor (layer0_outputs(9592)));
    outputs(3946) <= (layer0_outputs(5010)) and not (layer0_outputs(8396));
    outputs(3947) <= (layer0_outputs(415)) xor (layer0_outputs(8235));
    outputs(3948) <= not(layer0_outputs(5447)) or (layer0_outputs(75));
    outputs(3949) <= not(layer0_outputs(12)) or (layer0_outputs(7876));
    outputs(3950) <= not(layer0_outputs(2269));
    outputs(3951) <= layer0_outputs(5980);
    outputs(3952) <= (layer0_outputs(702)) xor (layer0_outputs(1932));
    outputs(3953) <= not(layer0_outputs(4098));
    outputs(3954) <= layer0_outputs(5595);
    outputs(3955) <= (layer0_outputs(1279)) or (layer0_outputs(1399));
    outputs(3956) <= not(layer0_outputs(297));
    outputs(3957) <= not(layer0_outputs(4260));
    outputs(3958) <= (layer0_outputs(4237)) and (layer0_outputs(4168));
    outputs(3959) <= layer0_outputs(718);
    outputs(3960) <= layer0_outputs(2409);
    outputs(3961) <= not(layer0_outputs(9635));
    outputs(3962) <= not(layer0_outputs(7554));
    outputs(3963) <= not((layer0_outputs(7374)) or (layer0_outputs(7295)));
    outputs(3964) <= not(layer0_outputs(10041));
    outputs(3965) <= layer0_outputs(3339);
    outputs(3966) <= (layer0_outputs(8188)) and not (layer0_outputs(6050));
    outputs(3967) <= (layer0_outputs(5662)) xor (layer0_outputs(5582));
    outputs(3968) <= layer0_outputs(7623);
    outputs(3969) <= not(layer0_outputs(6492));
    outputs(3970) <= not(layer0_outputs(4944));
    outputs(3971) <= not(layer0_outputs(4642));
    outputs(3972) <= not(layer0_outputs(2467));
    outputs(3973) <= layer0_outputs(4725);
    outputs(3974) <= (layer0_outputs(865)) and not (layer0_outputs(883));
    outputs(3975) <= layer0_outputs(10171);
    outputs(3976) <= (layer0_outputs(3860)) and (layer0_outputs(9178));
    outputs(3977) <= layer0_outputs(2115);
    outputs(3978) <= (layer0_outputs(4668)) xor (layer0_outputs(7493));
    outputs(3979) <= not((layer0_outputs(896)) xor (layer0_outputs(3230)));
    outputs(3980) <= (layer0_outputs(8694)) xor (layer0_outputs(10007));
    outputs(3981) <= (layer0_outputs(6898)) and (layer0_outputs(4409));
    outputs(3982) <= not((layer0_outputs(407)) xor (layer0_outputs(6370)));
    outputs(3983) <= (layer0_outputs(8337)) and (layer0_outputs(3024));
    outputs(3984) <= (layer0_outputs(4822)) xor (layer0_outputs(4831));
    outputs(3985) <= (layer0_outputs(3223)) and not (layer0_outputs(7879));
    outputs(3986) <= (layer0_outputs(5658)) xor (layer0_outputs(8186));
    outputs(3987) <= layer0_outputs(1887);
    outputs(3988) <= layer0_outputs(8898);
    outputs(3989) <= not(layer0_outputs(2491));
    outputs(3990) <= not(layer0_outputs(3778));
    outputs(3991) <= not(layer0_outputs(594));
    outputs(3992) <= (layer0_outputs(8666)) and not (layer0_outputs(10058));
    outputs(3993) <= not(layer0_outputs(9829));
    outputs(3994) <= (layer0_outputs(5845)) or (layer0_outputs(3512));
    outputs(3995) <= not(layer0_outputs(8635));
    outputs(3996) <= layer0_outputs(9973);
    outputs(3997) <= not((layer0_outputs(8186)) or (layer0_outputs(141)));
    outputs(3998) <= not((layer0_outputs(8344)) or (layer0_outputs(9373)));
    outputs(3999) <= (layer0_outputs(7987)) and not (layer0_outputs(5639));
    outputs(4000) <= layer0_outputs(1939);
    outputs(4001) <= (layer0_outputs(1398)) and not (layer0_outputs(1837));
    outputs(4002) <= (layer0_outputs(414)) xor (layer0_outputs(8011));
    outputs(4003) <= not((layer0_outputs(2512)) or (layer0_outputs(1383)));
    outputs(4004) <= (layer0_outputs(1382)) or (layer0_outputs(9087));
    outputs(4005) <= layer0_outputs(5162);
    outputs(4006) <= not((layer0_outputs(8953)) or (layer0_outputs(8551)));
    outputs(4007) <= not(layer0_outputs(1547));
    outputs(4008) <= (layer0_outputs(4504)) and not (layer0_outputs(554));
    outputs(4009) <= not(layer0_outputs(6020));
    outputs(4010) <= (layer0_outputs(6906)) and not (layer0_outputs(751));
    outputs(4011) <= layer0_outputs(8287);
    outputs(4012) <= layer0_outputs(7314);
    outputs(4013) <= (layer0_outputs(6229)) xor (layer0_outputs(5303));
    outputs(4014) <= (layer0_outputs(2626)) and not (layer0_outputs(8478));
    outputs(4015) <= not((layer0_outputs(5788)) xor (layer0_outputs(1616)));
    outputs(4016) <= not(layer0_outputs(9040));
    outputs(4017) <= layer0_outputs(8053);
    outputs(4018) <= not((layer0_outputs(9824)) xor (layer0_outputs(3402)));
    outputs(4019) <= not(layer0_outputs(60));
    outputs(4020) <= not(layer0_outputs(523));
    outputs(4021) <= layer0_outputs(3665);
    outputs(4022) <= not(layer0_outputs(4688));
    outputs(4023) <= (layer0_outputs(1805)) xor (layer0_outputs(5690));
    outputs(4024) <= not(layer0_outputs(4540));
    outputs(4025) <= not(layer0_outputs(5245));
    outputs(4026) <= layer0_outputs(5546);
    outputs(4027) <= not((layer0_outputs(4746)) or (layer0_outputs(5413)));
    outputs(4028) <= layer0_outputs(7162);
    outputs(4029) <= layer0_outputs(8117);
    outputs(4030) <= layer0_outputs(2719);
    outputs(4031) <= not(layer0_outputs(8199)) or (layer0_outputs(10054));
    outputs(4032) <= layer0_outputs(3099);
    outputs(4033) <= layer0_outputs(5418);
    outputs(4034) <= not((layer0_outputs(3085)) xor (layer0_outputs(5021)));
    outputs(4035) <= not(layer0_outputs(6209)) or (layer0_outputs(1945));
    outputs(4036) <= (layer0_outputs(5841)) or (layer0_outputs(7479));
    outputs(4037) <= layer0_outputs(187);
    outputs(4038) <= layer0_outputs(7294);
    outputs(4039) <= layer0_outputs(2497);
    outputs(4040) <= not(layer0_outputs(9119));
    outputs(4041) <= not(layer0_outputs(9885));
    outputs(4042) <= not((layer0_outputs(4372)) and (layer0_outputs(8107)));
    outputs(4043) <= layer0_outputs(8687);
    outputs(4044) <= (layer0_outputs(10143)) xor (layer0_outputs(9367));
    outputs(4045) <= not((layer0_outputs(1110)) xor (layer0_outputs(4295)));
    outputs(4046) <= (layer0_outputs(8807)) xor (layer0_outputs(6235));
    outputs(4047) <= layer0_outputs(9379);
    outputs(4048) <= not(layer0_outputs(4500));
    outputs(4049) <= layer0_outputs(2285);
    outputs(4050) <= (layer0_outputs(1577)) xor (layer0_outputs(2252));
    outputs(4051) <= not(layer0_outputs(752));
    outputs(4052) <= (layer0_outputs(7072)) and not (layer0_outputs(2308));
    outputs(4053) <= not(layer0_outputs(4219));
    outputs(4054) <= layer0_outputs(7352);
    outputs(4055) <= (layer0_outputs(7763)) or (layer0_outputs(8538));
    outputs(4056) <= layer0_outputs(4616);
    outputs(4057) <= layer0_outputs(5160);
    outputs(4058) <= not(layer0_outputs(3171));
    outputs(4059) <= not((layer0_outputs(8172)) xor (layer0_outputs(8981)));
    outputs(4060) <= (layer0_outputs(2746)) and (layer0_outputs(10205));
    outputs(4061) <= not(layer0_outputs(3707));
    outputs(4062) <= not(layer0_outputs(1634));
    outputs(4063) <= layer0_outputs(9059);
    outputs(4064) <= not(layer0_outputs(1506));
    outputs(4065) <= not((layer0_outputs(7737)) xor (layer0_outputs(2454)));
    outputs(4066) <= layer0_outputs(4073);
    outputs(4067) <= (layer0_outputs(7415)) and (layer0_outputs(914));
    outputs(4068) <= (layer0_outputs(24)) and (layer0_outputs(8771));
    outputs(4069) <= not((layer0_outputs(151)) xor (layer0_outputs(4482)));
    outputs(4070) <= not(layer0_outputs(3963)) or (layer0_outputs(9420));
    outputs(4071) <= not(layer0_outputs(9611));
    outputs(4072) <= layer0_outputs(1534);
    outputs(4073) <= (layer0_outputs(7229)) xor (layer0_outputs(291));
    outputs(4074) <= (layer0_outputs(6368)) and (layer0_outputs(5421));
    outputs(4075) <= layer0_outputs(2436);
    outputs(4076) <= not(layer0_outputs(2336));
    outputs(4077) <= layer0_outputs(9609);
    outputs(4078) <= (layer0_outputs(6806)) xor (layer0_outputs(8929));
    outputs(4079) <= layer0_outputs(8498);
    outputs(4080) <= (layer0_outputs(1759)) xor (layer0_outputs(4014));
    outputs(4081) <= layer0_outputs(6723);
    outputs(4082) <= not(layer0_outputs(1192)) or (layer0_outputs(674));
    outputs(4083) <= not(layer0_outputs(1814));
    outputs(4084) <= (layer0_outputs(2964)) and not (layer0_outputs(1152));
    outputs(4085) <= not(layer0_outputs(5349));
    outputs(4086) <= (layer0_outputs(5265)) and not (layer0_outputs(6870));
    outputs(4087) <= (layer0_outputs(6697)) xor (layer0_outputs(2782));
    outputs(4088) <= not(layer0_outputs(4425)) or (layer0_outputs(2494));
    outputs(4089) <= layer0_outputs(4476);
    outputs(4090) <= not((layer0_outputs(9917)) and (layer0_outputs(9102)));
    outputs(4091) <= layer0_outputs(197);
    outputs(4092) <= not((layer0_outputs(8850)) xor (layer0_outputs(3294)));
    outputs(4093) <= (layer0_outputs(7129)) and (layer0_outputs(3349));
    outputs(4094) <= layer0_outputs(6005);
    outputs(4095) <= (layer0_outputs(1236)) xor (layer0_outputs(8679));
    outputs(4096) <= layer0_outputs(797);
    outputs(4097) <= layer0_outputs(5252);
    outputs(4098) <= not(layer0_outputs(9647));
    outputs(4099) <= (layer0_outputs(931)) or (layer0_outputs(2235));
    outputs(4100) <= (layer0_outputs(8533)) and (layer0_outputs(444));
    outputs(4101) <= layer0_outputs(7964);
    outputs(4102) <= (layer0_outputs(10039)) or (layer0_outputs(6662));
    outputs(4103) <= not(layer0_outputs(4358));
    outputs(4104) <= not(layer0_outputs(5897)) or (layer0_outputs(2966));
    outputs(4105) <= not(layer0_outputs(3497));
    outputs(4106) <= layer0_outputs(8623);
    outputs(4107) <= not(layer0_outputs(5131));
    outputs(4108) <= layer0_outputs(4177);
    outputs(4109) <= not((layer0_outputs(7472)) and (layer0_outputs(5771)));
    outputs(4110) <= not(layer0_outputs(7337));
    outputs(4111) <= (layer0_outputs(8269)) and not (layer0_outputs(8137));
    outputs(4112) <= not(layer0_outputs(9429));
    outputs(4113) <= not(layer0_outputs(6081));
    outputs(4114) <= not(layer0_outputs(1490)) or (layer0_outputs(696));
    outputs(4115) <= not(layer0_outputs(8693));
    outputs(4116) <= not(layer0_outputs(273));
    outputs(4117) <= not(layer0_outputs(10055));
    outputs(4118) <= not(layer0_outputs(10061));
    outputs(4119) <= layer0_outputs(5358);
    outputs(4120) <= not((layer0_outputs(829)) or (layer0_outputs(9535)));
    outputs(4121) <= not(layer0_outputs(2900));
    outputs(4122) <= not(layer0_outputs(7883));
    outputs(4123) <= not((layer0_outputs(9622)) xor (layer0_outputs(989)));
    outputs(4124) <= layer0_outputs(5377);
    outputs(4125) <= not((layer0_outputs(4759)) xor (layer0_outputs(6827)));
    outputs(4126) <= layer0_outputs(7108);
    outputs(4127) <= not(layer0_outputs(686));
    outputs(4128) <= layer0_outputs(5182);
    outputs(4129) <= not(layer0_outputs(4596)) or (layer0_outputs(572));
    outputs(4130) <= layer0_outputs(10128);
    outputs(4131) <= not((layer0_outputs(5602)) xor (layer0_outputs(10092)));
    outputs(4132) <= not(layer0_outputs(9183)) or (layer0_outputs(5848));
    outputs(4133) <= layer0_outputs(1281);
    outputs(4134) <= layer0_outputs(269);
    outputs(4135) <= layer0_outputs(752);
    outputs(4136) <= (layer0_outputs(935)) and not (layer0_outputs(9049));
    outputs(4137) <= not(layer0_outputs(6752));
    outputs(4138) <= layer0_outputs(7424);
    outputs(4139) <= not(layer0_outputs(4370)) or (layer0_outputs(5402));
    outputs(4140) <= not(layer0_outputs(9551));
    outputs(4141) <= not(layer0_outputs(6195));
    outputs(4142) <= not(layer0_outputs(3676));
    outputs(4143) <= layer0_outputs(9083);
    outputs(4144) <= not(layer0_outputs(1529));
    outputs(4145) <= (layer0_outputs(6100)) and (layer0_outputs(9716));
    outputs(4146) <= (layer0_outputs(9540)) xor (layer0_outputs(6221));
    outputs(4147) <= (layer0_outputs(2068)) and not (layer0_outputs(7021));
    outputs(4148) <= not(layer0_outputs(9465));
    outputs(4149) <= not(layer0_outputs(4145));
    outputs(4150) <= (layer0_outputs(7840)) and (layer0_outputs(1242));
    outputs(4151) <= layer0_outputs(10135);
    outputs(4152) <= layer0_outputs(7388);
    outputs(4153) <= (layer0_outputs(2810)) and not (layer0_outputs(5979));
    outputs(4154) <= (layer0_outputs(785)) and (layer0_outputs(5136));
    outputs(4155) <= not((layer0_outputs(10230)) or (layer0_outputs(9773)));
    outputs(4156) <= (layer0_outputs(8883)) and not (layer0_outputs(4465));
    outputs(4157) <= not(layer0_outputs(3782));
    outputs(4158) <= not(layer0_outputs(4661));
    outputs(4159) <= (layer0_outputs(3517)) xor (layer0_outputs(2698));
    outputs(4160) <= layer0_outputs(52);
    outputs(4161) <= layer0_outputs(7069);
    outputs(4162) <= (layer0_outputs(5569)) xor (layer0_outputs(1442));
    outputs(4163) <= not(layer0_outputs(7750));
    outputs(4164) <= not(layer0_outputs(1559));
    outputs(4165) <= not(layer0_outputs(355));
    outputs(4166) <= not(layer0_outputs(3498));
    outputs(4167) <= not(layer0_outputs(5125));
    outputs(4168) <= not(layer0_outputs(3120));
    outputs(4169) <= not(layer0_outputs(3168));
    outputs(4170) <= not(layer0_outputs(10));
    outputs(4171) <= not(layer0_outputs(4543));
    outputs(4172) <= not(layer0_outputs(3496));
    outputs(4173) <= not(layer0_outputs(461));
    outputs(4174) <= not(layer0_outputs(3243)) or (layer0_outputs(2255));
    outputs(4175) <= (layer0_outputs(1732)) and not (layer0_outputs(9041));
    outputs(4176) <= not((layer0_outputs(2541)) and (layer0_outputs(1998)));
    outputs(4177) <= not(layer0_outputs(4702)) or (layer0_outputs(947));
    outputs(4178) <= not(layer0_outputs(8818)) or (layer0_outputs(7433));
    outputs(4179) <= (layer0_outputs(2660)) and not (layer0_outputs(6469));
    outputs(4180) <= layer0_outputs(7971);
    outputs(4181) <= not(layer0_outputs(5369));
    outputs(4182) <= not(layer0_outputs(2129));
    outputs(4183) <= layer0_outputs(7969);
    outputs(4184) <= not(layer0_outputs(6330));
    outputs(4185) <= layer0_outputs(764);
    outputs(4186) <= (layer0_outputs(8793)) xor (layer0_outputs(3229));
    outputs(4187) <= layer0_outputs(1996);
    outputs(4188) <= (layer0_outputs(5416)) and not (layer0_outputs(6248));
    outputs(4189) <= not((layer0_outputs(8819)) xor (layer0_outputs(5677)));
    outputs(4190) <= layer0_outputs(9338);
    outputs(4191) <= layer0_outputs(2109);
    outputs(4192) <= layer0_outputs(5030);
    outputs(4193) <= (layer0_outputs(10207)) and (layer0_outputs(8770));
    outputs(4194) <= not(layer0_outputs(6038));
    outputs(4195) <= layer0_outputs(1050);
    outputs(4196) <= (layer0_outputs(6377)) and (layer0_outputs(5149));
    outputs(4197) <= not((layer0_outputs(2416)) xor (layer0_outputs(8770)));
    outputs(4198) <= not((layer0_outputs(3898)) xor (layer0_outputs(10234)));
    outputs(4199) <= not(layer0_outputs(7572));
    outputs(4200) <= not(layer0_outputs(9465));
    outputs(4201) <= not((layer0_outputs(768)) or (layer0_outputs(8782)));
    outputs(4202) <= not(layer0_outputs(7688));
    outputs(4203) <= layer0_outputs(3578);
    outputs(4204) <= (layer0_outputs(7174)) xor (layer0_outputs(5421));
    outputs(4205) <= layer0_outputs(2780);
    outputs(4206) <= layer0_outputs(4817);
    outputs(4207) <= not(layer0_outputs(3757));
    outputs(4208) <= (layer0_outputs(2578)) or (layer0_outputs(2124));
    outputs(4209) <= not((layer0_outputs(3980)) xor (layer0_outputs(7565)));
    outputs(4210) <= (layer0_outputs(9848)) and not (layer0_outputs(1419));
    outputs(4211) <= layer0_outputs(5399);
    outputs(4212) <= not((layer0_outputs(5077)) or (layer0_outputs(119)));
    outputs(4213) <= not(layer0_outputs(3764));
    outputs(4214) <= layer0_outputs(215);
    outputs(4215) <= (layer0_outputs(3713)) and (layer0_outputs(8250));
    outputs(4216) <= (layer0_outputs(5834)) xor (layer0_outputs(9128));
    outputs(4217) <= layer0_outputs(4586);
    outputs(4218) <= layer0_outputs(7048);
    outputs(4219) <= layer0_outputs(9629);
    outputs(4220) <= not((layer0_outputs(3547)) and (layer0_outputs(7400)));
    outputs(4221) <= (layer0_outputs(3396)) and (layer0_outputs(3766));
    outputs(4222) <= not(layer0_outputs(5728));
    outputs(4223) <= not((layer0_outputs(5935)) or (layer0_outputs(1567)));
    outputs(4224) <= (layer0_outputs(2136)) and not (layer0_outputs(10230));
    outputs(4225) <= (layer0_outputs(8323)) and not (layer0_outputs(8228));
    outputs(4226) <= (layer0_outputs(4745)) and (layer0_outputs(8112));
    outputs(4227) <= not(layer0_outputs(4592)) or (layer0_outputs(3116));
    outputs(4228) <= layer0_outputs(9130);
    outputs(4229) <= layer0_outputs(7344);
    outputs(4230) <= not(layer0_outputs(612));
    outputs(4231) <= not(layer0_outputs(5870));
    outputs(4232) <= not(layer0_outputs(5318));
    outputs(4233) <= layer0_outputs(10217);
    outputs(4234) <= (layer0_outputs(1493)) and not (layer0_outputs(7990));
    outputs(4235) <= layer0_outputs(6992);
    outputs(4236) <= not(layer0_outputs(10100));
    outputs(4237) <= layer0_outputs(1213);
    outputs(4238) <= layer0_outputs(2648);
    outputs(4239) <= not(layer0_outputs(1466));
    outputs(4240) <= not(layer0_outputs(3059));
    outputs(4241) <= layer0_outputs(4397);
    outputs(4242) <= not(layer0_outputs(8183)) or (layer0_outputs(6337));
    outputs(4243) <= layer0_outputs(9296);
    outputs(4244) <= layer0_outputs(4315);
    outputs(4245) <= layer0_outputs(9196);
    outputs(4246) <= not(layer0_outputs(6289));
    outputs(4247) <= not((layer0_outputs(6250)) or (layer0_outputs(1165)));
    outputs(4248) <= layer0_outputs(2332);
    outputs(4249) <= layer0_outputs(2499);
    outputs(4250) <= not((layer0_outputs(2458)) and (layer0_outputs(6906)));
    outputs(4251) <= layer0_outputs(2140);
    outputs(4252) <= (layer0_outputs(738)) and not (layer0_outputs(3729));
    outputs(4253) <= layer0_outputs(5201);
    outputs(4254) <= layer0_outputs(5176);
    outputs(4255) <= not(layer0_outputs(651));
    outputs(4256) <= not(layer0_outputs(6455)) or (layer0_outputs(6046));
    outputs(4257) <= layer0_outputs(4294);
    outputs(4258) <= (layer0_outputs(4540)) and not (layer0_outputs(1265));
    outputs(4259) <= (layer0_outputs(10075)) or (layer0_outputs(8683));
    outputs(4260) <= not((layer0_outputs(9280)) xor (layer0_outputs(7201)));
    outputs(4261) <= layer0_outputs(1205);
    outputs(4262) <= layer0_outputs(7028);
    outputs(4263) <= layer0_outputs(8681);
    outputs(4264) <= not((layer0_outputs(8202)) xor (layer0_outputs(3829)));
    outputs(4265) <= (layer0_outputs(4282)) xor (layer0_outputs(448));
    outputs(4266) <= not((layer0_outputs(4062)) or (layer0_outputs(125)));
    outputs(4267) <= not(layer0_outputs(9493));
    outputs(4268) <= (layer0_outputs(6846)) or (layer0_outputs(1927));
    outputs(4269) <= not((layer0_outputs(3685)) or (layer0_outputs(4496)));
    outputs(4270) <= (layer0_outputs(3561)) and (layer0_outputs(4277));
    outputs(4271) <= (layer0_outputs(3108)) xor (layer0_outputs(5495));
    outputs(4272) <= (layer0_outputs(9303)) and not (layer0_outputs(1227));
    outputs(4273) <= not((layer0_outputs(4183)) or (layer0_outputs(4203)));
    outputs(4274) <= not((layer0_outputs(760)) or (layer0_outputs(5052)));
    outputs(4275) <= layer0_outputs(4086);
    outputs(4276) <= not(layer0_outputs(10100));
    outputs(4277) <= layer0_outputs(7735);
    outputs(4278) <= layer0_outputs(3908);
    outputs(4279) <= not(layer0_outputs(3692));
    outputs(4280) <= not((layer0_outputs(6096)) xor (layer0_outputs(3592)));
    outputs(4281) <= layer0_outputs(3966);
    outputs(4282) <= (layer0_outputs(7043)) and not (layer0_outputs(1550));
    outputs(4283) <= (layer0_outputs(8724)) and not (layer0_outputs(795));
    outputs(4284) <= (layer0_outputs(7251)) xor (layer0_outputs(3011));
    outputs(4285) <= not((layer0_outputs(406)) and (layer0_outputs(9621)));
    outputs(4286) <= not(layer0_outputs(45)) or (layer0_outputs(337));
    outputs(4287) <= not((layer0_outputs(5178)) and (layer0_outputs(4135)));
    outputs(4288) <= layer0_outputs(2369);
    outputs(4289) <= not(layer0_outputs(2237));
    outputs(4290) <= not((layer0_outputs(7027)) and (layer0_outputs(3661)));
    outputs(4291) <= not(layer0_outputs(3129));
    outputs(4292) <= layer0_outputs(821);
    outputs(4293) <= (layer0_outputs(2374)) and not (layer0_outputs(9790));
    outputs(4294) <= layer0_outputs(8178);
    outputs(4295) <= '0';
    outputs(4296) <= not(layer0_outputs(2949)) or (layer0_outputs(1539));
    outputs(4297) <= not(layer0_outputs(4118));
    outputs(4298) <= not(layer0_outputs(822)) or (layer0_outputs(8932));
    outputs(4299) <= layer0_outputs(5255);
    outputs(4300) <= not((layer0_outputs(10074)) xor (layer0_outputs(9861)));
    outputs(4301) <= layer0_outputs(584);
    outputs(4302) <= layer0_outputs(1627);
    outputs(4303) <= layer0_outputs(9010);
    outputs(4304) <= layer0_outputs(7739);
    outputs(4305) <= not(layer0_outputs(6294)) or (layer0_outputs(5532));
    outputs(4306) <= layer0_outputs(6769);
    outputs(4307) <= not(layer0_outputs(8895)) or (layer0_outputs(5455));
    outputs(4308) <= layer0_outputs(5220);
    outputs(4309) <= layer0_outputs(4729);
    outputs(4310) <= not(layer0_outputs(3319));
    outputs(4311) <= not((layer0_outputs(9483)) xor (layer0_outputs(9519)));
    outputs(4312) <= not(layer0_outputs(9474));
    outputs(4313) <= not((layer0_outputs(6839)) xor (layer0_outputs(8692)));
    outputs(4314) <= (layer0_outputs(1341)) xor (layer0_outputs(695));
    outputs(4315) <= not(layer0_outputs(4486));
    outputs(4316) <= layer0_outputs(4461);
    outputs(4317) <= layer0_outputs(1240);
    outputs(4318) <= not(layer0_outputs(6024));
    outputs(4319) <= not(layer0_outputs(5095)) or (layer0_outputs(247));
    outputs(4320) <= not(layer0_outputs(6921));
    outputs(4321) <= not(layer0_outputs(2844));
    outputs(4322) <= (layer0_outputs(8683)) xor (layer0_outputs(4730));
    outputs(4323) <= (layer0_outputs(5426)) and not (layer0_outputs(3371));
    outputs(4324) <= not((layer0_outputs(800)) xor (layer0_outputs(1337)));
    outputs(4325) <= not(layer0_outputs(3023));
    outputs(4326) <= (layer0_outputs(1920)) or (layer0_outputs(3738));
    outputs(4327) <= not((layer0_outputs(282)) and (layer0_outputs(3235)));
    outputs(4328) <= (layer0_outputs(9528)) and not (layer0_outputs(8839));
    outputs(4329) <= not(layer0_outputs(499)) or (layer0_outputs(3309));
    outputs(4330) <= layer0_outputs(1302);
    outputs(4331) <= not(layer0_outputs(3177)) or (layer0_outputs(4512));
    outputs(4332) <= not((layer0_outputs(7943)) xor (layer0_outputs(6055)));
    outputs(4333) <= not(layer0_outputs(9114)) or (layer0_outputs(7694));
    outputs(4334) <= (layer0_outputs(64)) and (layer0_outputs(5394));
    outputs(4335) <= not((layer0_outputs(3630)) xor (layer0_outputs(2774)));
    outputs(4336) <= not((layer0_outputs(5469)) or (layer0_outputs(4370)));
    outputs(4337) <= (layer0_outputs(6638)) and (layer0_outputs(9520));
    outputs(4338) <= (layer0_outputs(3908)) and (layer0_outputs(10199));
    outputs(4339) <= not(layer0_outputs(10172));
    outputs(4340) <= layer0_outputs(3959);
    outputs(4341) <= layer0_outputs(1321);
    outputs(4342) <= not(layer0_outputs(8435));
    outputs(4343) <= not(layer0_outputs(6411));
    outputs(4344) <= not(layer0_outputs(5769));
    outputs(4345) <= layer0_outputs(2488);
    outputs(4346) <= layer0_outputs(3520);
    outputs(4347) <= (layer0_outputs(10076)) and not (layer0_outputs(5787));
    outputs(4348) <= (layer0_outputs(8942)) or (layer0_outputs(1598));
    outputs(4349) <= not(layer0_outputs(4314));
    outputs(4350) <= layer0_outputs(6401);
    outputs(4351) <= layer0_outputs(4004);
    outputs(4352) <= layer0_outputs(8217);
    outputs(4353) <= not(layer0_outputs(3732)) or (layer0_outputs(8618));
    outputs(4354) <= layer0_outputs(9705);
    outputs(4355) <= not(layer0_outputs(6317));
    outputs(4356) <= not(layer0_outputs(2240)) or (layer0_outputs(2780));
    outputs(4357) <= not(layer0_outputs(2773));
    outputs(4358) <= not(layer0_outputs(8804)) or (layer0_outputs(2945));
    outputs(4359) <= (layer0_outputs(1411)) xor (layer0_outputs(9638));
    outputs(4360) <= not(layer0_outputs(3324)) or (layer0_outputs(2727));
    outputs(4361) <= layer0_outputs(1840);
    outputs(4362) <= layer0_outputs(7913);
    outputs(4363) <= not(layer0_outputs(7145));
    outputs(4364) <= not(layer0_outputs(10096));
    outputs(4365) <= not(layer0_outputs(2406));
    outputs(4366) <= (layer0_outputs(8653)) and not (layer0_outputs(3331));
    outputs(4367) <= (layer0_outputs(8080)) xor (layer0_outputs(6521));
    outputs(4368) <= not(layer0_outputs(933));
    outputs(4369) <= layer0_outputs(9742);
    outputs(4370) <= not(layer0_outputs(8117));
    outputs(4371) <= not((layer0_outputs(4040)) or (layer0_outputs(9645)));
    outputs(4372) <= (layer0_outputs(2564)) and (layer0_outputs(1624));
    outputs(4373) <= (layer0_outputs(8274)) and not (layer0_outputs(6970));
    outputs(4374) <= not(layer0_outputs(5630)) or (layer0_outputs(681));
    outputs(4375) <= (layer0_outputs(8212)) and not (layer0_outputs(6910));
    outputs(4376) <= layer0_outputs(6861);
    outputs(4377) <= not(layer0_outputs(3558));
    outputs(4378) <= not((layer0_outputs(3174)) or (layer0_outputs(8426)));
    outputs(4379) <= not(layer0_outputs(1969));
    outputs(4380) <= layer0_outputs(9813);
    outputs(4381) <= layer0_outputs(4654);
    outputs(4382) <= not(layer0_outputs(1406));
    outputs(4383) <= not(layer0_outputs(2048));
    outputs(4384) <= (layer0_outputs(854)) xor (layer0_outputs(2046));
    outputs(4385) <= not((layer0_outputs(5235)) or (layer0_outputs(6001)));
    outputs(4386) <= (layer0_outputs(2638)) and not (layer0_outputs(4251));
    outputs(4387) <= (layer0_outputs(1880)) xor (layer0_outputs(430));
    outputs(4388) <= layer0_outputs(5439);
    outputs(4389) <= (layer0_outputs(9194)) xor (layer0_outputs(2037));
    outputs(4390) <= (layer0_outputs(9206)) and not (layer0_outputs(159));
    outputs(4391) <= layer0_outputs(6433);
    outputs(4392) <= (layer0_outputs(9043)) and not (layer0_outputs(8299));
    outputs(4393) <= not((layer0_outputs(9024)) xor (layer0_outputs(3740)));
    outputs(4394) <= not(layer0_outputs(5481));
    outputs(4395) <= layer0_outputs(4342);
    outputs(4396) <= layer0_outputs(4316);
    outputs(4397) <= layer0_outputs(805);
    outputs(4398) <= not((layer0_outputs(6794)) or (layer0_outputs(2981)));
    outputs(4399) <= (layer0_outputs(6928)) and not (layer0_outputs(5631));
    outputs(4400) <= layer0_outputs(8630);
    outputs(4401) <= not(layer0_outputs(813));
    outputs(4402) <= not(layer0_outputs(3043));
    outputs(4403) <= layer0_outputs(3412);
    outputs(4404) <= (layer0_outputs(5248)) xor (layer0_outputs(2027));
    outputs(4405) <= not((layer0_outputs(8573)) xor (layer0_outputs(4998)));
    outputs(4406) <= layer0_outputs(5528);
    outputs(4407) <= (layer0_outputs(1020)) and (layer0_outputs(1244));
    outputs(4408) <= (layer0_outputs(1839)) and not (layer0_outputs(9842));
    outputs(4409) <= (layer0_outputs(290)) and not (layer0_outputs(799));
    outputs(4410) <= (layer0_outputs(2717)) and not (layer0_outputs(117));
    outputs(4411) <= layer0_outputs(7000);
    outputs(4412) <= layer0_outputs(300);
    outputs(4413) <= layer0_outputs(1109);
    outputs(4414) <= layer0_outputs(6596);
    outputs(4415) <= not((layer0_outputs(8707)) xor (layer0_outputs(5191)));
    outputs(4416) <= layer0_outputs(1326);
    outputs(4417) <= not(layer0_outputs(8689));
    outputs(4418) <= not(layer0_outputs(1643));
    outputs(4419) <= not((layer0_outputs(10079)) and (layer0_outputs(5540)));
    outputs(4420) <= not(layer0_outputs(9));
    outputs(4421) <= (layer0_outputs(4635)) and not (layer0_outputs(7616));
    outputs(4422) <= not(layer0_outputs(5924));
    outputs(4423) <= not(layer0_outputs(9292));
    outputs(4424) <= not(layer0_outputs(41));
    outputs(4425) <= (layer0_outputs(3918)) or (layer0_outputs(6033));
    outputs(4426) <= not(layer0_outputs(2418));
    outputs(4427) <= (layer0_outputs(7483)) and not (layer0_outputs(4798));
    outputs(4428) <= not(layer0_outputs(3430));
    outputs(4429) <= layer0_outputs(5043);
    outputs(4430) <= not(layer0_outputs(3799));
    outputs(4431) <= not((layer0_outputs(3282)) xor (layer0_outputs(5648)));
    outputs(4432) <= (layer0_outputs(3290)) or (layer0_outputs(402));
    outputs(4433) <= (layer0_outputs(7450)) and not (layer0_outputs(5129));
    outputs(4434) <= not((layer0_outputs(9988)) or (layer0_outputs(3092)));
    outputs(4435) <= not(layer0_outputs(3121));
    outputs(4436) <= (layer0_outputs(8656)) xor (layer0_outputs(2877));
    outputs(4437) <= not(layer0_outputs(1572));
    outputs(4438) <= not(layer0_outputs(1994));
    outputs(4439) <= not(layer0_outputs(875)) or (layer0_outputs(6995));
    outputs(4440) <= (layer0_outputs(10001)) and not (layer0_outputs(3111));
    outputs(4441) <= not(layer0_outputs(131)) or (layer0_outputs(2903));
    outputs(4442) <= layer0_outputs(3462);
    outputs(4443) <= layer0_outputs(3042);
    outputs(4444) <= layer0_outputs(5772);
    outputs(4445) <= not((layer0_outputs(7893)) xor (layer0_outputs(5860)));
    outputs(4446) <= (layer0_outputs(7614)) xor (layer0_outputs(6341));
    outputs(4447) <= not((layer0_outputs(8132)) xor (layer0_outputs(7396)));
    outputs(4448) <= not(layer0_outputs(2704)) or (layer0_outputs(2342));
    outputs(4449) <= not((layer0_outputs(6820)) xor (layer0_outputs(6015)));
    outputs(4450) <= not(layer0_outputs(4252));
    outputs(4451) <= (layer0_outputs(4122)) and (layer0_outputs(5579));
    outputs(4452) <= (layer0_outputs(6162)) xor (layer0_outputs(5849));
    outputs(4453) <= not(layer0_outputs(926));
    outputs(4454) <= not((layer0_outputs(1139)) xor (layer0_outputs(229)));
    outputs(4455) <= (layer0_outputs(4925)) and (layer0_outputs(9752));
    outputs(4456) <= (layer0_outputs(7720)) and (layer0_outputs(1953));
    outputs(4457) <= not(layer0_outputs(9805));
    outputs(4458) <= not((layer0_outputs(1049)) or (layer0_outputs(1637)));
    outputs(4459) <= (layer0_outputs(6592)) and (layer0_outputs(8135));
    outputs(4460) <= (layer0_outputs(5342)) and not (layer0_outputs(7451));
    outputs(4461) <= not(layer0_outputs(3107));
    outputs(4462) <= layer0_outputs(3127);
    outputs(4463) <= not(layer0_outputs(1807));
    outputs(4464) <= not(layer0_outputs(3940));
    outputs(4465) <= (layer0_outputs(582)) xor (layer0_outputs(9295));
    outputs(4466) <= layer0_outputs(4785);
    outputs(4467) <= not((layer0_outputs(1608)) xor (layer0_outputs(1090)));
    outputs(4468) <= not(layer0_outputs(256)) or (layer0_outputs(1179));
    outputs(4469) <= not(layer0_outputs(2534));
    outputs(4470) <= not(layer0_outputs(3074));
    outputs(4471) <= layer0_outputs(483);
    outputs(4472) <= not((layer0_outputs(3896)) or (layer0_outputs(3117)));
    outputs(4473) <= layer0_outputs(2778);
    outputs(4474) <= layer0_outputs(5122);
    outputs(4475) <= (layer0_outputs(3437)) xor (layer0_outputs(3871));
    outputs(4476) <= not(layer0_outputs(10068));
    outputs(4477) <= layer0_outputs(2190);
    outputs(4478) <= not((layer0_outputs(1665)) xor (layer0_outputs(1088)));
    outputs(4479) <= layer0_outputs(8759);
    outputs(4480) <= layer0_outputs(6258);
    outputs(4481) <= not((layer0_outputs(4604)) and (layer0_outputs(5839)));
    outputs(4482) <= not(layer0_outputs(5729)) or (layer0_outputs(7394));
    outputs(4483) <= not((layer0_outputs(3532)) or (layer0_outputs(353)));
    outputs(4484) <= (layer0_outputs(1264)) and not (layer0_outputs(8485));
    outputs(4485) <= not((layer0_outputs(9576)) xor (layer0_outputs(1704)));
    outputs(4486) <= not(layer0_outputs(1160));
    outputs(4487) <= not(layer0_outputs(8465));
    outputs(4488) <= not(layer0_outputs(2085));
    outputs(4489) <= layer0_outputs(6700);
    outputs(4490) <= not((layer0_outputs(7324)) xor (layer0_outputs(5610)));
    outputs(4491) <= not(layer0_outputs(6698)) or (layer0_outputs(4753));
    outputs(4492) <= not(layer0_outputs(9844));
    outputs(4493) <= (layer0_outputs(4706)) and not (layer0_outputs(9709));
    outputs(4494) <= (layer0_outputs(3920)) and (layer0_outputs(9900));
    outputs(4495) <= not(layer0_outputs(969));
    outputs(4496) <= (layer0_outputs(6431)) and (layer0_outputs(9282));
    outputs(4497) <= not(layer0_outputs(5065)) or (layer0_outputs(6023));
    outputs(4498) <= (layer0_outputs(9364)) and not (layer0_outputs(8930));
    outputs(4499) <= layer0_outputs(3407);
    outputs(4500) <= not(layer0_outputs(8292));
    outputs(4501) <= not((layer0_outputs(5487)) or (layer0_outputs(5261)));
    outputs(4502) <= not(layer0_outputs(3865)) or (layer0_outputs(3584));
    outputs(4503) <= layer0_outputs(4824);
    outputs(4504) <= not(layer0_outputs(3378));
    outputs(4505) <= (layer0_outputs(6788)) and not (layer0_outputs(6733));
    outputs(4506) <= layer0_outputs(3857);
    outputs(4507) <= layer0_outputs(9517);
    outputs(4508) <= layer0_outputs(3549);
    outputs(4509) <= not(layer0_outputs(1601));
    outputs(4510) <= layer0_outputs(9369);
    outputs(4511) <= not(layer0_outputs(7949));
    outputs(4512) <= not((layer0_outputs(1568)) xor (layer0_outputs(4607)));
    outputs(4513) <= not((layer0_outputs(9402)) or (layer0_outputs(4042)));
    outputs(4514) <= not((layer0_outputs(932)) xor (layer0_outputs(1230)));
    outputs(4515) <= (layer0_outputs(4414)) and not (layer0_outputs(960));
    outputs(4516) <= layer0_outputs(2303);
    outputs(4517) <= not((layer0_outputs(2313)) xor (layer0_outputs(3350)));
    outputs(4518) <= not((layer0_outputs(6236)) xor (layer0_outputs(6652)));
    outputs(4519) <= (layer0_outputs(5780)) and not (layer0_outputs(8859));
    outputs(4520) <= (layer0_outputs(5533)) xor (layer0_outputs(5986));
    outputs(4521) <= (layer0_outputs(2963)) and not (layer0_outputs(4327));
    outputs(4522) <= (layer0_outputs(7681)) and (layer0_outputs(2631));
    outputs(4523) <= not(layer0_outputs(4510));
    outputs(4524) <= layer0_outputs(4506);
    outputs(4525) <= layer0_outputs(8284);
    outputs(4526) <= (layer0_outputs(8478)) or (layer0_outputs(6270));
    outputs(4527) <= layer0_outputs(2058);
    outputs(4528) <= layer0_outputs(6549);
    outputs(4529) <= (layer0_outputs(3185)) xor (layer0_outputs(6605));
    outputs(4530) <= not(layer0_outputs(5321));
    outputs(4531) <= not((layer0_outputs(2831)) xor (layer0_outputs(3675)));
    outputs(4532) <= (layer0_outputs(3464)) and (layer0_outputs(8606));
    outputs(4533) <= not((layer0_outputs(4854)) xor (layer0_outputs(5480)));
    outputs(4534) <= not((layer0_outputs(1542)) or (layer0_outputs(6762)));
    outputs(4535) <= (layer0_outputs(329)) xor (layer0_outputs(7939));
    outputs(4536) <= (layer0_outputs(7507)) and (layer0_outputs(7189));
    outputs(4537) <= (layer0_outputs(4918)) xor (layer0_outputs(6223));
    outputs(4538) <= not(layer0_outputs(3622));
    outputs(4539) <= layer0_outputs(9582);
    outputs(4540) <= layer0_outputs(9009);
    outputs(4541) <= not(layer0_outputs(1215));
    outputs(4542) <= not(layer0_outputs(6283));
    outputs(4543) <= layer0_outputs(443);
    outputs(4544) <= not(layer0_outputs(7585));
    outputs(4545) <= (layer0_outputs(5814)) or (layer0_outputs(9104));
    outputs(4546) <= not(layer0_outputs(7378));
    outputs(4547) <= not(layer0_outputs(3162));
    outputs(4548) <= layer0_outputs(7596);
    outputs(4549) <= not((layer0_outputs(9326)) or (layer0_outputs(7192)));
    outputs(4550) <= not(layer0_outputs(164));
    outputs(4551) <= (layer0_outputs(761)) and not (layer0_outputs(4616));
    outputs(4552) <= layer0_outputs(5372);
    outputs(4553) <= layer0_outputs(6675);
    outputs(4554) <= layer0_outputs(1119);
    outputs(4555) <= not((layer0_outputs(9821)) or (layer0_outputs(793)));
    outputs(4556) <= not((layer0_outputs(8001)) xor (layer0_outputs(8858)));
    outputs(4557) <= not(layer0_outputs(2823)) or (layer0_outputs(1700));
    outputs(4558) <= not((layer0_outputs(10034)) xor (layer0_outputs(8281)));
    outputs(4559) <= not(layer0_outputs(2231));
    outputs(4560) <= not(layer0_outputs(4267));
    outputs(4561) <= layer0_outputs(343);
    outputs(4562) <= not(layer0_outputs(111));
    outputs(4563) <= (layer0_outputs(1181)) xor (layer0_outputs(7476));
    outputs(4564) <= not(layer0_outputs(5404)) or (layer0_outputs(7781));
    outputs(4565) <= not(layer0_outputs(2004));
    outputs(4566) <= not(layer0_outputs(4270));
    outputs(4567) <= not(layer0_outputs(790));
    outputs(4568) <= layer0_outputs(6401);
    outputs(4569) <= not((layer0_outputs(9045)) or (layer0_outputs(3331)));
    outputs(4570) <= (layer0_outputs(7323)) and not (layer0_outputs(6025));
    outputs(4571) <= layer0_outputs(5444);
    outputs(4572) <= layer0_outputs(9612);
    outputs(4573) <= (layer0_outputs(7567)) xor (layer0_outputs(2542));
    outputs(4574) <= not(layer0_outputs(2795));
    outputs(4575) <= (layer0_outputs(716)) xor (layer0_outputs(8124));
    outputs(4576) <= not((layer0_outputs(4200)) and (layer0_outputs(2726)));
    outputs(4577) <= not(layer0_outputs(3679));
    outputs(4578) <= layer0_outputs(5385);
    outputs(4579) <= not(layer0_outputs(984));
    outputs(4580) <= not(layer0_outputs(5632));
    outputs(4581) <= (layer0_outputs(307)) and (layer0_outputs(2583));
    outputs(4582) <= (layer0_outputs(9917)) or (layer0_outputs(535));
    outputs(4583) <= layer0_outputs(7588);
    outputs(4584) <= not(layer0_outputs(5713));
    outputs(4585) <= layer0_outputs(5721);
    outputs(4586) <= not(layer0_outputs(7248));
    outputs(4587) <= not(layer0_outputs(1633));
    outputs(4588) <= not(layer0_outputs(3837));
    outputs(4589) <= (layer0_outputs(6097)) and not (layer0_outputs(9859));
    outputs(4590) <= not(layer0_outputs(2071)) or (layer0_outputs(3851));
    outputs(4591) <= not(layer0_outputs(10228));
    outputs(4592) <= layer0_outputs(3672);
    outputs(4593) <= not(layer0_outputs(2762));
    outputs(4594) <= not(layer0_outputs(3981));
    outputs(4595) <= not((layer0_outputs(9775)) xor (layer0_outputs(8247)));
    outputs(4596) <= (layer0_outputs(306)) xor (layer0_outputs(7715));
    outputs(4597) <= (layer0_outputs(6113)) and not (layer0_outputs(3989));
    outputs(4598) <= not((layer0_outputs(1435)) xor (layer0_outputs(5704)));
    outputs(4599) <= (layer0_outputs(9719)) and not (layer0_outputs(1571));
    outputs(4600) <= (layer0_outputs(8434)) and (layer0_outputs(9256));
    outputs(4601) <= not((layer0_outputs(5640)) xor (layer0_outputs(7877)));
    outputs(4602) <= not((layer0_outputs(5155)) xor (layer0_outputs(1549)));
    outputs(4603) <= not((layer0_outputs(8204)) xor (layer0_outputs(2421)));
    outputs(4604) <= (layer0_outputs(8051)) and not (layer0_outputs(8137));
    outputs(4605) <= not(layer0_outputs(4527));
    outputs(4606) <= layer0_outputs(2589);
    outputs(4607) <= (layer0_outputs(988)) and (layer0_outputs(2354));
    outputs(4608) <= not(layer0_outputs(4140));
    outputs(4609) <= not(layer0_outputs(5460));
    outputs(4610) <= not(layer0_outputs(10079)) or (layer0_outputs(8943));
    outputs(4611) <= not(layer0_outputs(9451));
    outputs(4612) <= (layer0_outputs(6200)) and not (layer0_outputs(4901));
    outputs(4613) <= not(layer0_outputs(2174));
    outputs(4614) <= not(layer0_outputs(7817));
    outputs(4615) <= not(layer0_outputs(1238));
    outputs(4616) <= not(layer0_outputs(4772));
    outputs(4617) <= (layer0_outputs(7974)) and not (layer0_outputs(5475));
    outputs(4618) <= not((layer0_outputs(10106)) xor (layer0_outputs(6310)));
    outputs(4619) <= layer0_outputs(5170);
    outputs(4620) <= layer0_outputs(8825);
    outputs(4621) <= (layer0_outputs(9677)) and (layer0_outputs(3973));
    outputs(4622) <= not(layer0_outputs(5475));
    outputs(4623) <= (layer0_outputs(9542)) and not (layer0_outputs(4038));
    outputs(4624) <= not(layer0_outputs(748));
    outputs(4625) <= layer0_outputs(7637);
    outputs(4626) <= (layer0_outputs(9265)) xor (layer0_outputs(4643));
    outputs(4627) <= not((layer0_outputs(274)) or (layer0_outputs(2986)));
    outputs(4628) <= (layer0_outputs(5757)) xor (layer0_outputs(762));
    outputs(4629) <= not(layer0_outputs(8923));
    outputs(4630) <= not((layer0_outputs(5135)) or (layer0_outputs(3648)));
    outputs(4631) <= layer0_outputs(7898);
    outputs(4632) <= layer0_outputs(7203);
    outputs(4633) <= (layer0_outputs(6075)) and (layer0_outputs(2796));
    outputs(4634) <= not((layer0_outputs(9251)) or (layer0_outputs(2690)));
    outputs(4635) <= not(layer0_outputs(6336));
    outputs(4636) <= (layer0_outputs(5228)) xor (layer0_outputs(4468));
    outputs(4637) <= (layer0_outputs(3240)) and (layer0_outputs(1543));
    outputs(4638) <= not(layer0_outputs(6426));
    outputs(4639) <= not(layer0_outputs(7624));
    outputs(4640) <= not((layer0_outputs(9220)) or (layer0_outputs(2925)));
    outputs(4641) <= not(layer0_outputs(2562));
    outputs(4642) <= not(layer0_outputs(6545)) or (layer0_outputs(8293));
    outputs(4643) <= layer0_outputs(3545);
    outputs(4644) <= (layer0_outputs(990)) and (layer0_outputs(2302));
    outputs(4645) <= layer0_outputs(1743);
    outputs(4646) <= not(layer0_outputs(1878));
    outputs(4647) <= not(layer0_outputs(10072));
    outputs(4648) <= (layer0_outputs(6161)) and (layer0_outputs(7948));
    outputs(4649) <= (layer0_outputs(9847)) xor (layer0_outputs(9634));
    outputs(4650) <= not(layer0_outputs(7250));
    outputs(4651) <= not(layer0_outputs(4200)) or (layer0_outputs(2428));
    outputs(4652) <= not((layer0_outputs(9787)) and (layer0_outputs(6941)));
    outputs(4653) <= (layer0_outputs(8682)) xor (layer0_outputs(5853));
    outputs(4654) <= not(layer0_outputs(7983));
    outputs(4655) <= (layer0_outputs(4093)) or (layer0_outputs(535));
    outputs(4656) <= not((layer0_outputs(5813)) xor (layer0_outputs(414)));
    outputs(4657) <= (layer0_outputs(3369)) and not (layer0_outputs(6030));
    outputs(4658) <= (layer0_outputs(455)) and (layer0_outputs(8847));
    outputs(4659) <= not(layer0_outputs(8093));
    outputs(4660) <= (layer0_outputs(6987)) xor (layer0_outputs(2487));
    outputs(4661) <= not(layer0_outputs(6539));
    outputs(4662) <= not(layer0_outputs(6998));
    outputs(4663) <= (layer0_outputs(2028)) and (layer0_outputs(7906));
    outputs(4664) <= (layer0_outputs(3766)) and not (layer0_outputs(7311));
    outputs(4665) <= not(layer0_outputs(4644));
    outputs(4666) <= layer0_outputs(8056);
    outputs(4667) <= not(layer0_outputs(6366));
    outputs(4668) <= not(layer0_outputs(9992));
    outputs(4669) <= not(layer0_outputs(9031));
    outputs(4670) <= (layer0_outputs(490)) and not (layer0_outputs(9736));
    outputs(4671) <= layer0_outputs(9672);
    outputs(4672) <= not((layer0_outputs(143)) and (layer0_outputs(5065)));
    outputs(4673) <= not((layer0_outputs(6059)) or (layer0_outputs(4534)));
    outputs(4674) <= not(layer0_outputs(8078));
    outputs(4675) <= layer0_outputs(2386);
    outputs(4676) <= not(layer0_outputs(7150));
    outputs(4677) <= layer0_outputs(3549);
    outputs(4678) <= not((layer0_outputs(6329)) or (layer0_outputs(2864)));
    outputs(4679) <= not(layer0_outputs(3974));
    outputs(4680) <= (layer0_outputs(9895)) and not (layer0_outputs(1729));
    outputs(4681) <= layer0_outputs(10160);
    outputs(4682) <= layer0_outputs(1078);
    outputs(4683) <= not(layer0_outputs(9313));
    outputs(4684) <= not(layer0_outputs(859)) or (layer0_outputs(5676));
    outputs(4685) <= not(layer0_outputs(6838)) or (layer0_outputs(4657));
    outputs(4686) <= not(layer0_outputs(1006));
    outputs(4687) <= not(layer0_outputs(5770));
    outputs(4688) <= not(layer0_outputs(8431));
    outputs(4689) <= not((layer0_outputs(4079)) xor (layer0_outputs(1788)));
    outputs(4690) <= not(layer0_outputs(882));
    outputs(4691) <= not((layer0_outputs(7331)) xor (layer0_outputs(1154)));
    outputs(4692) <= layer0_outputs(706);
    outputs(4693) <= not(layer0_outputs(1881));
    outputs(4694) <= (layer0_outputs(5792)) and (layer0_outputs(904));
    outputs(4695) <= not(layer0_outputs(4131));
    outputs(4696) <= layer0_outputs(7562);
    outputs(4697) <= (layer0_outputs(4688)) and (layer0_outputs(8491));
    outputs(4698) <= layer0_outputs(8742);
    outputs(4699) <= not((layer0_outputs(927)) and (layer0_outputs(8248)));
    outputs(4700) <= (layer0_outputs(6581)) and (layer0_outputs(8134));
    outputs(4701) <= not(layer0_outputs(9967)) or (layer0_outputs(6300));
    outputs(4702) <= not(layer0_outputs(8565));
    outputs(4703) <= layer0_outputs(7309);
    outputs(4704) <= (layer0_outputs(3039)) xor (layer0_outputs(9978));
    outputs(4705) <= layer0_outputs(1316);
    outputs(4706) <= not(layer0_outputs(6369));
    outputs(4707) <= not((layer0_outputs(3056)) xor (layer0_outputs(6518)));
    outputs(4708) <= (layer0_outputs(893)) and not (layer0_outputs(1361));
    outputs(4709) <= not(layer0_outputs(3173)) or (layer0_outputs(6870));
    outputs(4710) <= not(layer0_outputs(8665));
    outputs(4711) <= (layer0_outputs(5173)) and not (layer0_outputs(1463));
    outputs(4712) <= layer0_outputs(4840);
    outputs(4713) <= not(layer0_outputs(4197));
    outputs(4714) <= (layer0_outputs(5282)) xor (layer0_outputs(7004));
    outputs(4715) <= not(layer0_outputs(5266));
    outputs(4716) <= not(layer0_outputs(8649));
    outputs(4717) <= (layer0_outputs(6996)) or (layer0_outputs(2652));
    outputs(4718) <= (layer0_outputs(70)) and not (layer0_outputs(8867));
    outputs(4719) <= not(layer0_outputs(8319));
    outputs(4720) <= layer0_outputs(4951);
    outputs(4721) <= not((layer0_outputs(207)) xor (layer0_outputs(6831)));
    outputs(4722) <= not(layer0_outputs(5405)) or (layer0_outputs(5714));
    outputs(4723) <= layer0_outputs(5337);
    outputs(4724) <= (layer0_outputs(9494)) or (layer0_outputs(8863));
    outputs(4725) <= (layer0_outputs(6186)) and not (layer0_outputs(4988));
    outputs(4726) <= not(layer0_outputs(6420));
    outputs(4727) <= not(layer0_outputs(5153));
    outputs(4728) <= layer0_outputs(7114);
    outputs(4729) <= not(layer0_outputs(5773));
    outputs(4730) <= not(layer0_outputs(3854));
    outputs(4731) <= not(layer0_outputs(9349));
    outputs(4732) <= layer0_outputs(1935);
    outputs(4733) <= (layer0_outputs(3699)) and (layer0_outputs(6421));
    outputs(4734) <= not(layer0_outputs(7922));
    outputs(4735) <= not(layer0_outputs(2777)) or (layer0_outputs(1817));
    outputs(4736) <= layer0_outputs(4917);
    outputs(4737) <= not(layer0_outputs(1983));
    outputs(4738) <= not((layer0_outputs(9997)) and (layer0_outputs(8308)));
    outputs(4739) <= not(layer0_outputs(7606));
    outputs(4740) <= not((layer0_outputs(10164)) xor (layer0_outputs(3452)));
    outputs(4741) <= (layer0_outputs(9649)) xor (layer0_outputs(3383));
    outputs(4742) <= layer0_outputs(6701);
    outputs(4743) <= not(layer0_outputs(10010));
    outputs(4744) <= not(layer0_outputs(7697));
    outputs(4745) <= layer0_outputs(4454);
    outputs(4746) <= layer0_outputs(9692);
    outputs(4747) <= not(layer0_outputs(9119));
    outputs(4748) <= layer0_outputs(8650);
    outputs(4749) <= not(layer0_outputs(5810));
    outputs(4750) <= layer0_outputs(5104);
    outputs(4751) <= (layer0_outputs(1536)) and not (layer0_outputs(3220));
    outputs(4752) <= layer0_outputs(9104);
    outputs(4753) <= not(layer0_outputs(5463));
    outputs(4754) <= (layer0_outputs(1140)) xor (layer0_outputs(5100));
    outputs(4755) <= not(layer0_outputs(4393));
    outputs(4756) <= (layer0_outputs(7869)) and not (layer0_outputs(7624));
    outputs(4757) <= (layer0_outputs(1119)) and not (layer0_outputs(4217));
    outputs(4758) <= layer0_outputs(3420);
    outputs(4759) <= not(layer0_outputs(7107));
    outputs(4760) <= not(layer0_outputs(9415));
    outputs(4761) <= layer0_outputs(5037);
    outputs(4762) <= layer0_outputs(2869);
    outputs(4763) <= not((layer0_outputs(10095)) xor (layer0_outputs(3899)));
    outputs(4764) <= layer0_outputs(1554);
    outputs(4765) <= (layer0_outputs(7224)) xor (layer0_outputs(6097));
    outputs(4766) <= layer0_outputs(6154);
    outputs(4767) <= not(layer0_outputs(3433));
    outputs(4768) <= not((layer0_outputs(5784)) xor (layer0_outputs(2678)));
    outputs(4769) <= (layer0_outputs(5983)) or (layer0_outputs(8889));
    outputs(4770) <= not((layer0_outputs(4672)) xor (layer0_outputs(2208)));
    outputs(4771) <= layer0_outputs(2234);
    outputs(4772) <= (layer0_outputs(1199)) and (layer0_outputs(3061));
    outputs(4773) <= layer0_outputs(1660);
    outputs(4774) <= not((layer0_outputs(6799)) xor (layer0_outputs(4122)));
    outputs(4775) <= layer0_outputs(6373);
    outputs(4776) <= (layer0_outputs(5217)) xor (layer0_outputs(4023));
    outputs(4777) <= not(layer0_outputs(4319));
    outputs(4778) <= not((layer0_outputs(6540)) xor (layer0_outputs(2883)));
    outputs(4779) <= (layer0_outputs(3515)) xor (layer0_outputs(9602));
    outputs(4780) <= (layer0_outputs(5850)) and not (layer0_outputs(965));
    outputs(4781) <= layer0_outputs(6895);
    outputs(4782) <= not(layer0_outputs(1373));
    outputs(4783) <= not(layer0_outputs(5712)) or (layer0_outputs(5585));
    outputs(4784) <= layer0_outputs(7661);
    outputs(4785) <= (layer0_outputs(864)) and not (layer0_outputs(4954));
    outputs(4786) <= (layer0_outputs(1661)) and (layer0_outputs(8880));
    outputs(4787) <= (layer0_outputs(8326)) and (layer0_outputs(915));
    outputs(4788) <= not((layer0_outputs(3558)) xor (layer0_outputs(9396)));
    outputs(4789) <= not(layer0_outputs(4584));
    outputs(4790) <= layer0_outputs(2573);
    outputs(4791) <= not(layer0_outputs(8610)) or (layer0_outputs(3108));
    outputs(4792) <= layer0_outputs(4924);
    outputs(4793) <= layer0_outputs(7923);
    outputs(4794) <= (layer0_outputs(788)) and not (layer0_outputs(895));
    outputs(4795) <= not((layer0_outputs(319)) and (layer0_outputs(4483)));
    outputs(4796) <= (layer0_outputs(1632)) xor (layer0_outputs(6084));
    outputs(4797) <= (layer0_outputs(9905)) and (layer0_outputs(2907));
    outputs(4798) <= not(layer0_outputs(563));
    outputs(4799) <= (layer0_outputs(3416)) and (layer0_outputs(561));
    outputs(4800) <= not((layer0_outputs(4450)) or (layer0_outputs(9155)));
    outputs(4801) <= not(layer0_outputs(9976));
    outputs(4802) <= (layer0_outputs(6708)) xor (layer0_outputs(8503));
    outputs(4803) <= not((layer0_outputs(6189)) xor (layer0_outputs(3617)));
    outputs(4804) <= layer0_outputs(3857);
    outputs(4805) <= not(layer0_outputs(7533));
    outputs(4806) <= not(layer0_outputs(6910));
    outputs(4807) <= layer0_outputs(949);
    outputs(4808) <= (layer0_outputs(1271)) and not (layer0_outputs(884));
    outputs(4809) <= not((layer0_outputs(9028)) or (layer0_outputs(8795)));
    outputs(4810) <= not(layer0_outputs(2048));
    outputs(4811) <= not((layer0_outputs(3745)) or (layer0_outputs(5454)));
    outputs(4812) <= layer0_outputs(10148);
    outputs(4813) <= not(layer0_outputs(2799));
    outputs(4814) <= (layer0_outputs(9200)) or (layer0_outputs(2249));
    outputs(4815) <= layer0_outputs(10213);
    outputs(4816) <= not((layer0_outputs(8921)) or (layer0_outputs(6130)));
    outputs(4817) <= not(layer0_outputs(8049));
    outputs(4818) <= not(layer0_outputs(4660));
    outputs(4819) <= not(layer0_outputs(7965));
    outputs(4820) <= not(layer0_outputs(6629));
    outputs(4821) <= not(layer0_outputs(5822));
    outputs(4822) <= (layer0_outputs(1681)) and not (layer0_outputs(8499));
    outputs(4823) <= layer0_outputs(8251);
    outputs(4824) <= not(layer0_outputs(8191));
    outputs(4825) <= not(layer0_outputs(4845));
    outputs(4826) <= not(layer0_outputs(1739));
    outputs(4827) <= layer0_outputs(948);
    outputs(4828) <= layer0_outputs(4939);
    outputs(4829) <= not(layer0_outputs(8362));
    outputs(4830) <= not((layer0_outputs(5949)) xor (layer0_outputs(2944)));
    outputs(4831) <= (layer0_outputs(6017)) and (layer0_outputs(3139));
    outputs(4832) <= not(layer0_outputs(4594));
    outputs(4833) <= not(layer0_outputs(8834));
    outputs(4834) <= layer0_outputs(10177);
    outputs(4835) <= (layer0_outputs(6553)) and not (layer0_outputs(5403));
    outputs(4836) <= not(layer0_outputs(5311));
    outputs(4837) <= not((layer0_outputs(1620)) xor (layer0_outputs(1715)));
    outputs(4838) <= (layer0_outputs(3593)) xor (layer0_outputs(1668));
    outputs(4839) <= layer0_outputs(3901);
    outputs(4840) <= layer0_outputs(5764);
    outputs(4841) <= layer0_outputs(5204);
    outputs(4842) <= not(layer0_outputs(3427));
    outputs(4843) <= not((layer0_outputs(1809)) xor (layer0_outputs(8461)));
    outputs(4844) <= layer0_outputs(187);
    outputs(4845) <= (layer0_outputs(9173)) and not (layer0_outputs(6468));
    outputs(4846) <= layer0_outputs(5548);
    outputs(4847) <= (layer0_outputs(6492)) or (layer0_outputs(9224));
    outputs(4848) <= layer0_outputs(6282);
    outputs(4849) <= not((layer0_outputs(3631)) xor (layer0_outputs(8795)));
    outputs(4850) <= not(layer0_outputs(7382));
    outputs(4851) <= (layer0_outputs(954)) and (layer0_outputs(6962));
    outputs(4852) <= (layer0_outputs(4311)) xor (layer0_outputs(3267));
    outputs(4853) <= not((layer0_outputs(787)) or (layer0_outputs(7843)));
    outputs(4854) <= (layer0_outputs(3209)) and not (layer0_outputs(9212));
    outputs(4855) <= not(layer0_outputs(9633));
    outputs(4856) <= not(layer0_outputs(2743));
    outputs(4857) <= (layer0_outputs(7834)) xor (layer0_outputs(10108));
    outputs(4858) <= not(layer0_outputs(5278));
    outputs(4859) <= not(layer0_outputs(327));
    outputs(4860) <= layer0_outputs(9595);
    outputs(4861) <= not(layer0_outputs(8108));
    outputs(4862) <= not((layer0_outputs(9377)) xor (layer0_outputs(1915)));
    outputs(4863) <= not((layer0_outputs(1719)) xor (layer0_outputs(2480)));
    outputs(4864) <= not(layer0_outputs(2956)) or (layer0_outputs(5994));
    outputs(4865) <= not(layer0_outputs(2180));
    outputs(4866) <= (layer0_outputs(10151)) xor (layer0_outputs(6689));
    outputs(4867) <= (layer0_outputs(885)) xor (layer0_outputs(6041));
    outputs(4868) <= not(layer0_outputs(284));
    outputs(4869) <= layer0_outputs(2771);
    outputs(4870) <= not(layer0_outputs(3333));
    outputs(4871) <= layer0_outputs(8637);
    outputs(4872) <= not(layer0_outputs(6622)) or (layer0_outputs(2333));
    outputs(4873) <= not(layer0_outputs(5935));
    outputs(4874) <= not((layer0_outputs(4738)) xor (layer0_outputs(3363)));
    outputs(4875) <= (layer0_outputs(7941)) xor (layer0_outputs(9527));
    outputs(4876) <= (layer0_outputs(2892)) and not (layer0_outputs(909));
    outputs(4877) <= layer0_outputs(3487);
    outputs(4878) <= not(layer0_outputs(7175));
    outputs(4879) <= not(layer0_outputs(6830));
    outputs(4880) <= not(layer0_outputs(882));
    outputs(4881) <= not((layer0_outputs(3416)) xor (layer0_outputs(1392)));
    outputs(4882) <= (layer0_outputs(4270)) xor (layer0_outputs(8928));
    outputs(4883) <= (layer0_outputs(2112)) and not (layer0_outputs(6912));
    outputs(4884) <= (layer0_outputs(6241)) and not (layer0_outputs(8141));
    outputs(4885) <= not(layer0_outputs(10057));
    outputs(4886) <= (layer0_outputs(3684)) and not (layer0_outputs(10145));
    outputs(4887) <= layer0_outputs(6003);
    outputs(4888) <= (layer0_outputs(3847)) and not (layer0_outputs(9139));
    outputs(4889) <= not(layer0_outputs(6707));
    outputs(4890) <= not(layer0_outputs(246));
    outputs(4891) <= (layer0_outputs(3718)) and (layer0_outputs(6436));
    outputs(4892) <= layer0_outputs(7212);
    outputs(4893) <= layer0_outputs(4703);
    outputs(4894) <= not(layer0_outputs(4186));
    outputs(4895) <= not((layer0_outputs(7466)) xor (layer0_outputs(5684)));
    outputs(4896) <= layer0_outputs(8578);
    outputs(4897) <= not((layer0_outputs(4328)) xor (layer0_outputs(4445)));
    outputs(4898) <= (layer0_outputs(6309)) or (layer0_outputs(1649));
    outputs(4899) <= (layer0_outputs(4755)) or (layer0_outputs(647));
    outputs(4900) <= layer0_outputs(4411);
    outputs(4901) <= (layer0_outputs(5798)) and (layer0_outputs(9013));
    outputs(4902) <= not((layer0_outputs(7024)) xor (layer0_outputs(3601)));
    outputs(4903) <= not(layer0_outputs(7340));
    outputs(4904) <= layer0_outputs(572);
    outputs(4905) <= layer0_outputs(7372);
    outputs(4906) <= not(layer0_outputs(7157));
    outputs(4907) <= (layer0_outputs(231)) xor (layer0_outputs(7924));
    outputs(4908) <= layer0_outputs(681);
    outputs(4909) <= not(layer0_outputs(7873));
    outputs(4910) <= layer0_outputs(3460);
    outputs(4911) <= layer0_outputs(3156);
    outputs(4912) <= layer0_outputs(7791);
    outputs(4913) <= layer0_outputs(2162);
    outputs(4914) <= not(layer0_outputs(3033));
    outputs(4915) <= layer0_outputs(5000);
    outputs(4916) <= not(layer0_outputs(9054));
    outputs(4917) <= layer0_outputs(2832);
    outputs(4918) <= not(layer0_outputs(2094));
    outputs(4919) <= not((layer0_outputs(6517)) or (layer0_outputs(1459)));
    outputs(4920) <= not(layer0_outputs(1599));
    outputs(4921) <= layer0_outputs(1769);
    outputs(4922) <= not((layer0_outputs(7908)) and (layer0_outputs(2226)));
    outputs(4923) <= layer0_outputs(10044);
    outputs(4924) <= (layer0_outputs(5449)) xor (layer0_outputs(10070));
    outputs(4925) <= not(layer0_outputs(4930)) or (layer0_outputs(2845));
    outputs(4926) <= (layer0_outputs(2577)) and not (layer0_outputs(9840));
    outputs(4927) <= not(layer0_outputs(7845));
    outputs(4928) <= not(layer0_outputs(9960)) or (layer0_outputs(1956));
    outputs(4929) <= (layer0_outputs(2793)) and not (layer0_outputs(9884));
    outputs(4930) <= (layer0_outputs(6895)) or (layer0_outputs(1771));
    outputs(4931) <= layer0_outputs(1548);
    outputs(4932) <= layer0_outputs(4397);
    outputs(4933) <= (layer0_outputs(10154)) and not (layer0_outputs(4935));
    outputs(4934) <= not((layer0_outputs(1100)) or (layer0_outputs(6234)));
    outputs(4935) <= (layer0_outputs(5844)) xor (layer0_outputs(7951));
    outputs(4936) <= not((layer0_outputs(9004)) or (layer0_outputs(4381)));
    outputs(4937) <= not(layer0_outputs(4472));
    outputs(4938) <= not(layer0_outputs(4111));
    outputs(4939) <= not(layer0_outputs(9947));
    outputs(4940) <= (layer0_outputs(5543)) xor (layer0_outputs(8789));
    outputs(4941) <= not(layer0_outputs(9853)) or (layer0_outputs(4231));
    outputs(4942) <= not(layer0_outputs(8102));
    outputs(4943) <= not((layer0_outputs(3093)) xor (layer0_outputs(8160)));
    outputs(4944) <= not(layer0_outputs(6287));
    outputs(4945) <= (layer0_outputs(10184)) and not (layer0_outputs(9834));
    outputs(4946) <= (layer0_outputs(2805)) xor (layer0_outputs(1810));
    outputs(4947) <= layer0_outputs(5534);
    outputs(4948) <= not((layer0_outputs(5609)) xor (layer0_outputs(5558)));
    outputs(4949) <= not((layer0_outputs(4775)) xor (layer0_outputs(6046)));
    outputs(4950) <= layer0_outputs(6863);
    outputs(4951) <= layer0_outputs(5964);
    outputs(4952) <= not(layer0_outputs(2281));
    outputs(4953) <= not(layer0_outputs(6899));
    outputs(4954) <= not(layer0_outputs(9805));
    outputs(4955) <= not(layer0_outputs(6576));
    outputs(4956) <= not(layer0_outputs(2914));
    outputs(4957) <= (layer0_outputs(1299)) and not (layer0_outputs(8809));
    outputs(4958) <= (layer0_outputs(2599)) and not (layer0_outputs(1278));
    outputs(4959) <= layer0_outputs(5720);
    outputs(4960) <= layer0_outputs(1055);
    outputs(4961) <= layer0_outputs(4113);
    outputs(4962) <= not((layer0_outputs(8407)) xor (layer0_outputs(8870)));
    outputs(4963) <= not(layer0_outputs(4632));
    outputs(4964) <= (layer0_outputs(5967)) and (layer0_outputs(5811));
    outputs(4965) <= not((layer0_outputs(4723)) xor (layer0_outputs(9091)));
    outputs(4966) <= layer0_outputs(6721);
    outputs(4967) <= not(layer0_outputs(3854));
    outputs(4968) <= layer0_outputs(6099);
    outputs(4969) <= (layer0_outputs(6332)) and not (layer0_outputs(6938));
    outputs(4970) <= not((layer0_outputs(6351)) xor (layer0_outputs(7371)));
    outputs(4971) <= not(layer0_outputs(897));
    outputs(4972) <= layer0_outputs(8285);
    outputs(4973) <= not(layer0_outputs(5205));
    outputs(4974) <= (layer0_outputs(6634)) xor (layer0_outputs(703));
    outputs(4975) <= layer0_outputs(3809);
    outputs(4976) <= not(layer0_outputs(1404));
    outputs(4977) <= not(layer0_outputs(7033));
    outputs(4978) <= layer0_outputs(3303);
    outputs(4979) <= not((layer0_outputs(7447)) or (layer0_outputs(6610)));
    outputs(4980) <= layer0_outputs(8276);
    outputs(4981) <= (layer0_outputs(2551)) xor (layer0_outputs(4017));
    outputs(4982) <= (layer0_outputs(5122)) and (layer0_outputs(3452));
    outputs(4983) <= (layer0_outputs(4453)) and not (layer0_outputs(5705));
    outputs(4984) <= not(layer0_outputs(7649));
    outputs(4985) <= not(layer0_outputs(405));
    outputs(4986) <= layer0_outputs(2310);
    outputs(4987) <= (layer0_outputs(2711)) and not (layer0_outputs(9263));
    outputs(4988) <= (layer0_outputs(9617)) and (layer0_outputs(1088));
    outputs(4989) <= (layer0_outputs(2453)) or (layer0_outputs(7787));
    outputs(4990) <= not((layer0_outputs(2327)) and (layer0_outputs(488)));
    outputs(4991) <= layer0_outputs(8905);
    outputs(4992) <= not(layer0_outputs(8421));
    outputs(4993) <= not((layer0_outputs(7985)) or (layer0_outputs(3866)));
    outputs(4994) <= not(layer0_outputs(7682));
    outputs(4995) <= (layer0_outputs(7824)) and (layer0_outputs(4224));
    outputs(4996) <= layer0_outputs(876);
    outputs(4997) <= not(layer0_outputs(6018)) or (layer0_outputs(6522));
    outputs(4998) <= not((layer0_outputs(5120)) xor (layer0_outputs(7469)));
    outputs(4999) <= (layer0_outputs(4598)) and not (layer0_outputs(2952));
    outputs(5000) <= layer0_outputs(4124);
    outputs(5001) <= not(layer0_outputs(9664)) or (layer0_outputs(7498));
    outputs(5002) <= layer0_outputs(7165);
    outputs(5003) <= layer0_outputs(232);
    outputs(5004) <= layer0_outputs(4939);
    outputs(5005) <= layer0_outputs(9261);
    outputs(5006) <= layer0_outputs(6154);
    outputs(5007) <= not(layer0_outputs(5161));
    outputs(5008) <= not((layer0_outputs(4946)) xor (layer0_outputs(8712)));
    outputs(5009) <= layer0_outputs(439);
    outputs(5010) <= not((layer0_outputs(6357)) or (layer0_outputs(9156)));
    outputs(5011) <= not((layer0_outputs(7531)) xor (layer0_outputs(5424)));
    outputs(5012) <= (layer0_outputs(617)) xor (layer0_outputs(6575));
    outputs(5013) <= not((layer0_outputs(847)) xor (layer0_outputs(2327)));
    outputs(5014) <= layer0_outputs(4093);
    outputs(5015) <= (layer0_outputs(1262)) xor (layer0_outputs(7216));
    outputs(5016) <= layer0_outputs(2635);
    outputs(5017) <= layer0_outputs(4719);
    outputs(5018) <= layer0_outputs(6258);
    outputs(5019) <= not((layer0_outputs(5197)) xor (layer0_outputs(9686)));
    outputs(5020) <= not(layer0_outputs(3027));
    outputs(5021) <= (layer0_outputs(8562)) and not (layer0_outputs(1973));
    outputs(5022) <= layer0_outputs(5832);
    outputs(5023) <= (layer0_outputs(6502)) and not (layer0_outputs(5061));
    outputs(5024) <= not((layer0_outputs(6650)) and (layer0_outputs(6088)));
    outputs(5025) <= not(layer0_outputs(7688));
    outputs(5026) <= (layer0_outputs(666)) xor (layer0_outputs(9160));
    outputs(5027) <= layer0_outputs(3733);
    outputs(5028) <= not(layer0_outputs(1201)) or (layer0_outputs(1447));
    outputs(5029) <= not(layer0_outputs(5185));
    outputs(5030) <= not(layer0_outputs(6499));
    outputs(5031) <= not(layer0_outputs(6187));
    outputs(5032) <= (layer0_outputs(1606)) or (layer0_outputs(6560));
    outputs(5033) <= not((layer0_outputs(1755)) and (layer0_outputs(1395)));
    outputs(5034) <= not((layer0_outputs(5620)) or (layer0_outputs(4983)));
    outputs(5035) <= not(layer0_outputs(1805));
    outputs(5036) <= not(layer0_outputs(2240)) or (layer0_outputs(6275));
    outputs(5037) <= not((layer0_outputs(4262)) xor (layer0_outputs(1930)));
    outputs(5038) <= not(layer0_outputs(1510));
    outputs(5039) <= layer0_outputs(10223);
    outputs(5040) <= (layer0_outputs(7422)) and not (layer0_outputs(8530));
    outputs(5041) <= not(layer0_outputs(4332));
    outputs(5042) <= not(layer0_outputs(1189));
    outputs(5043) <= not(layer0_outputs(1223));
    outputs(5044) <= not(layer0_outputs(10072));
    outputs(5045) <= not(layer0_outputs(5034)) or (layer0_outputs(9950));
    outputs(5046) <= not(layer0_outputs(4303)) or (layer0_outputs(2584));
    outputs(5047) <= not((layer0_outputs(6860)) xor (layer0_outputs(8935)));
    outputs(5048) <= (layer0_outputs(3982)) xor (layer0_outputs(4987));
    outputs(5049) <= not((layer0_outputs(2587)) or (layer0_outputs(4855)));
    outputs(5050) <= not(layer0_outputs(7434));
    outputs(5051) <= (layer0_outputs(6905)) and not (layer0_outputs(8218));
    outputs(5052) <= layer0_outputs(4037);
    outputs(5053) <= not(layer0_outputs(326)) or (layer0_outputs(3404));
    outputs(5054) <= not((layer0_outputs(8385)) xor (layer0_outputs(6045)));
    outputs(5055) <= not((layer0_outputs(3423)) xor (layer0_outputs(2112)));
    outputs(5056) <= not((layer0_outputs(6151)) xor (layer0_outputs(8828)));
    outputs(5057) <= (layer0_outputs(8663)) and not (layer0_outputs(7702));
    outputs(5058) <= (layer0_outputs(5201)) xor (layer0_outputs(4572));
    outputs(5059) <= not(layer0_outputs(2011)) or (layer0_outputs(1412));
    outputs(5060) <= layer0_outputs(7596);
    outputs(5061) <= (layer0_outputs(123)) xor (layer0_outputs(5326));
    outputs(5062) <= layer0_outputs(774);
    outputs(5063) <= (layer0_outputs(8862)) and (layer0_outputs(7188));
    outputs(5064) <= layer0_outputs(2707);
    outputs(5065) <= not(layer0_outputs(872));
    outputs(5066) <= layer0_outputs(5221);
    outputs(5067) <= (layer0_outputs(8949)) and not (layer0_outputs(380));
    outputs(5068) <= not(layer0_outputs(2413));
    outputs(5069) <= not((layer0_outputs(2232)) or (layer0_outputs(7254)));
    outputs(5070) <= not((layer0_outputs(9835)) or (layer0_outputs(9147)));
    outputs(5071) <= not((layer0_outputs(532)) or (layer0_outputs(5597)));
    outputs(5072) <= not(layer0_outputs(2482)) or (layer0_outputs(6601));
    outputs(5073) <= not(layer0_outputs(10015));
    outputs(5074) <= not(layer0_outputs(4564));
    outputs(5075) <= not((layer0_outputs(9992)) or (layer0_outputs(7008)));
    outputs(5076) <= not(layer0_outputs(7640));
    outputs(5077) <= layer0_outputs(2724);
    outputs(5078) <= layer0_outputs(5877);
    outputs(5079) <= not(layer0_outputs(2625)) or (layer0_outputs(5366));
    outputs(5080) <= not(layer0_outputs(5103));
    outputs(5081) <= (layer0_outputs(1877)) or (layer0_outputs(9636));
    outputs(5082) <= (layer0_outputs(6432)) xor (layer0_outputs(10055));
    outputs(5083) <= not(layer0_outputs(6907));
    outputs(5084) <= not((layer0_outputs(6210)) xor (layer0_outputs(3677)));
    outputs(5085) <= not((layer0_outputs(8374)) and (layer0_outputs(4313)));
    outputs(5086) <= not((layer0_outputs(4783)) xor (layer0_outputs(8971)));
    outputs(5087) <= not(layer0_outputs(5754));
    outputs(5088) <= (layer0_outputs(8544)) and not (layer0_outputs(9474));
    outputs(5089) <= not((layer0_outputs(1283)) or (layer0_outputs(8619)));
    outputs(5090) <= not(layer0_outputs(9530));
    outputs(5091) <= layer0_outputs(1272);
    outputs(5092) <= layer0_outputs(3639);
    outputs(5093) <= not(layer0_outputs(2514));
    outputs(5094) <= (layer0_outputs(1012)) xor (layer0_outputs(4977));
    outputs(5095) <= layer0_outputs(7029);
    outputs(5096) <= (layer0_outputs(1500)) and not (layer0_outputs(5915));
    outputs(5097) <= not((layer0_outputs(165)) xor (layer0_outputs(920)));
    outputs(5098) <= layer0_outputs(9518);
    outputs(5099) <= layer0_outputs(2623);
    outputs(5100) <= layer0_outputs(7068);
    outputs(5101) <= not(layer0_outputs(7271));
    outputs(5102) <= layer0_outputs(5913);
    outputs(5103) <= layer0_outputs(7195);
    outputs(5104) <= '1';
    outputs(5105) <= layer0_outputs(7279);
    outputs(5106) <= not(layer0_outputs(135));
    outputs(5107) <= not(layer0_outputs(9164));
    outputs(5108) <= layer0_outputs(3233);
    outputs(5109) <= layer0_outputs(4415);
    outputs(5110) <= (layer0_outputs(3666)) and not (layer0_outputs(4624));
    outputs(5111) <= (layer0_outputs(9729)) xor (layer0_outputs(466));
    outputs(5112) <= (layer0_outputs(338)) and not (layer0_outputs(7607));
    outputs(5113) <= (layer0_outputs(6094)) and (layer0_outputs(1320));
    outputs(5114) <= layer0_outputs(4881);
    outputs(5115) <= not((layer0_outputs(5269)) xor (layer0_outputs(4733)));
    outputs(5116) <= not((layer0_outputs(292)) or (layer0_outputs(1153)));
    outputs(5117) <= (layer0_outputs(8800)) or (layer0_outputs(2060));
    outputs(5118) <= layer0_outputs(3127);
    outputs(5119) <= layer0_outputs(10155);
    outputs(5120) <= not(layer0_outputs(6365));
    outputs(5121) <= (layer0_outputs(127)) xor (layer0_outputs(7810));
    outputs(5122) <= not((layer0_outputs(9584)) or (layer0_outputs(850)));
    outputs(5123) <= not((layer0_outputs(1115)) or (layer0_outputs(8540)));
    outputs(5124) <= not((layer0_outputs(8240)) or (layer0_outputs(6719)));
    outputs(5125) <= layer0_outputs(1564);
    outputs(5126) <= not(layer0_outputs(6149));
    outputs(5127) <= not((layer0_outputs(726)) xor (layer0_outputs(2173)));
    outputs(5128) <= (layer0_outputs(7560)) xor (layer0_outputs(2740));
    outputs(5129) <= not(layer0_outputs(8214));
    outputs(5130) <= layer0_outputs(7001);
    outputs(5131) <= (layer0_outputs(5166)) and not (layer0_outputs(5855));
    outputs(5132) <= (layer0_outputs(3518)) and not (layer0_outputs(4018));
    outputs(5133) <= not((layer0_outputs(6818)) xor (layer0_outputs(7616)));
    outputs(5134) <= (layer0_outputs(440)) or (layer0_outputs(8756));
    outputs(5135) <= not((layer0_outputs(1941)) or (layer0_outputs(812)));
    outputs(5136) <= (layer0_outputs(8152)) and not (layer0_outputs(8603));
    outputs(5137) <= not((layer0_outputs(39)) xor (layer0_outputs(1360)));
    outputs(5138) <= not((layer0_outputs(2609)) xor (layer0_outputs(4160)));
    outputs(5139) <= not(layer0_outputs(5654));
    outputs(5140) <= not(layer0_outputs(5241));
    outputs(5141) <= layer0_outputs(4737);
    outputs(5142) <= (layer0_outputs(8343)) xor (layer0_outputs(5571));
    outputs(5143) <= layer0_outputs(7407);
    outputs(5144) <= (layer0_outputs(6775)) and not (layer0_outputs(8881));
    outputs(5145) <= not(layer0_outputs(5753)) or (layer0_outputs(3022));
    outputs(5146) <= not(layer0_outputs(7910));
    outputs(5147) <= not(layer0_outputs(5997));
    outputs(5148) <= (layer0_outputs(1515)) xor (layer0_outputs(7321));
    outputs(5149) <= (layer0_outputs(2049)) and not (layer0_outputs(6660));
    outputs(5150) <= layer0_outputs(3472);
    outputs(5151) <= not((layer0_outputs(2649)) xor (layer0_outputs(2202)));
    outputs(5152) <= not((layer0_outputs(8312)) xor (layer0_outputs(768)));
    outputs(5153) <= not((layer0_outputs(4312)) or (layer0_outputs(3686)));
    outputs(5154) <= not((layer0_outputs(9663)) xor (layer0_outputs(1830)));
    outputs(5155) <= (layer0_outputs(56)) xor (layer0_outputs(4454));
    outputs(5156) <= not((layer0_outputs(4043)) or (layer0_outputs(5519)));
    outputs(5157) <= not(layer0_outputs(1977));
    outputs(5158) <= (layer0_outputs(4857)) xor (layer0_outputs(7821));
    outputs(5159) <= (layer0_outputs(2510)) xor (layer0_outputs(4157));
    outputs(5160) <= layer0_outputs(775);
    outputs(5161) <= not((layer0_outputs(2102)) xor (layer0_outputs(6221)));
    outputs(5162) <= (layer0_outputs(2073)) and (layer0_outputs(9525));
    outputs(5163) <= (layer0_outputs(8505)) or (layer0_outputs(304));
    outputs(5164) <= layer0_outputs(5888);
    outputs(5165) <= not((layer0_outputs(9079)) xor (layer0_outputs(8896)));
    outputs(5166) <= layer0_outputs(7205);
    outputs(5167) <= not((layer0_outputs(6609)) xor (layer0_outputs(2041)));
    outputs(5168) <= (layer0_outputs(270)) xor (layer0_outputs(1639));
    outputs(5169) <= (layer0_outputs(4382)) and not (layer0_outputs(1415));
    outputs(5170) <= (layer0_outputs(9500)) and (layer0_outputs(4797));
    outputs(5171) <= not(layer0_outputs(1178));
    outputs(5172) <= not(layer0_outputs(1931));
    outputs(5173) <= layer0_outputs(479);
    outputs(5174) <= not(layer0_outputs(756)) or (layer0_outputs(2637));
    outputs(5175) <= (layer0_outputs(4858)) and not (layer0_outputs(57));
    outputs(5176) <= layer0_outputs(4148);
    outputs(5177) <= (layer0_outputs(7435)) xor (layer0_outputs(3696));
    outputs(5178) <= layer0_outputs(9021);
    outputs(5179) <= layer0_outputs(3434);
    outputs(5180) <= not((layer0_outputs(1846)) xor (layer0_outputs(1757)));
    outputs(5181) <= (layer0_outputs(8446)) and not (layer0_outputs(8038));
    outputs(5182) <= layer0_outputs(9963);
    outputs(5183) <= not(layer0_outputs(5017));
    outputs(5184) <= (layer0_outputs(6934)) and not (layer0_outputs(9543));
    outputs(5185) <= layer0_outputs(5411);
    outputs(5186) <= (layer0_outputs(1838)) or (layer0_outputs(9362));
    outputs(5187) <= layer0_outputs(3278);
    outputs(5188) <= not((layer0_outputs(8537)) or (layer0_outputs(1600)));
    outputs(5189) <= not((layer0_outputs(3071)) or (layer0_outputs(990)));
    outputs(5190) <= layer0_outputs(6956);
    outputs(5191) <= not(layer0_outputs(2871));
    outputs(5192) <= (layer0_outputs(8376)) and not (layer0_outputs(2886));
    outputs(5193) <= (layer0_outputs(2833)) xor (layer0_outputs(6436));
    outputs(5194) <= (layer0_outputs(4680)) and not (layer0_outputs(8546));
    outputs(5195) <= not(layer0_outputs(4105));
    outputs(5196) <= (layer0_outputs(3581)) and not (layer0_outputs(7742));
    outputs(5197) <= not(layer0_outputs(2759));
    outputs(5198) <= not(layer0_outputs(8954));
    outputs(5199) <= layer0_outputs(8453);
    outputs(5200) <= (layer0_outputs(314)) xor (layer0_outputs(443));
    outputs(5201) <= (layer0_outputs(4212)) and (layer0_outputs(8265));
    outputs(5202) <= not((layer0_outputs(2126)) xor (layer0_outputs(1959)));
    outputs(5203) <= not(layer0_outputs(2462));
    outputs(5204) <= not(layer0_outputs(1790));
    outputs(5205) <= not(layer0_outputs(6960));
    outputs(5206) <= not(layer0_outputs(3527));
    outputs(5207) <= not((layer0_outputs(1139)) xor (layer0_outputs(3464)));
    outputs(5208) <= (layer0_outputs(7508)) xor (layer0_outputs(5158));
    outputs(5209) <= not(layer0_outputs(6141));
    outputs(5210) <= not(layer0_outputs(9411));
    outputs(5211) <= (layer0_outputs(722)) xor (layer0_outputs(8181));
    outputs(5212) <= layer0_outputs(7657);
    outputs(5213) <= not(layer0_outputs(5063));
    outputs(5214) <= (layer0_outputs(3628)) xor (layer0_outputs(9540));
    outputs(5215) <= not(layer0_outputs(9430));
    outputs(5216) <= (layer0_outputs(7555)) and not (layer0_outputs(4720));
    outputs(5217) <= (layer0_outputs(8702)) and (layer0_outputs(4244));
    outputs(5218) <= (layer0_outputs(6705)) or (layer0_outputs(6409));
    outputs(5219) <= '1';
    outputs(5220) <= not(layer0_outputs(9644)) or (layer0_outputs(4574));
    outputs(5221) <= not(layer0_outputs(9832));
    outputs(5222) <= not(layer0_outputs(5700)) or (layer0_outputs(7551));
    outputs(5223) <= not((layer0_outputs(497)) or (layer0_outputs(3038)));
    outputs(5224) <= (layer0_outputs(7409)) xor (layer0_outputs(2858));
    outputs(5225) <= layer0_outputs(3339);
    outputs(5226) <= not(layer0_outputs(10045));
    outputs(5227) <= not(layer0_outputs(4610));
    outputs(5228) <= not(layer0_outputs(1752)) or (layer0_outputs(6805));
    outputs(5229) <= not(layer0_outputs(1173));
    outputs(5230) <= not((layer0_outputs(7330)) xor (layer0_outputs(5202)));
    outputs(5231) <= layer0_outputs(2005);
    outputs(5232) <= not(layer0_outputs(3909));
    outputs(5233) <= layer0_outputs(9480);
    outputs(5234) <= not((layer0_outputs(9841)) xor (layer0_outputs(5423)));
    outputs(5235) <= not(layer0_outputs(6614));
    outputs(5236) <= layer0_outputs(3254);
    outputs(5237) <= not(layer0_outputs(4796)) or (layer0_outputs(2714));
    outputs(5238) <= not((layer0_outputs(9590)) and (layer0_outputs(2733)));
    outputs(5239) <= not((layer0_outputs(2639)) xor (layer0_outputs(1756)));
    outputs(5240) <= not((layer0_outputs(5092)) xor (layer0_outputs(6951)));
    outputs(5241) <= layer0_outputs(9820);
    outputs(5242) <= layer0_outputs(2023);
    outputs(5243) <= layer0_outputs(8099);
    outputs(5244) <= not(layer0_outputs(6534));
    outputs(5245) <= (layer0_outputs(7730)) xor (layer0_outputs(8425));
    outputs(5246) <= not(layer0_outputs(5189));
    outputs(5247) <= (layer0_outputs(5763)) xor (layer0_outputs(4448));
    outputs(5248) <= (layer0_outputs(6529)) and (layer0_outputs(7269));
    outputs(5249) <= (layer0_outputs(7205)) xor (layer0_outputs(1029));
    outputs(5250) <= (layer0_outputs(6525)) and not (layer0_outputs(8518));
    outputs(5251) <= not((layer0_outputs(4420)) xor (layer0_outputs(4789)));
    outputs(5252) <= not(layer0_outputs(6036));
    outputs(5253) <= layer0_outputs(8262);
    outputs(5254) <= layer0_outputs(4499);
    outputs(5255) <= not(layer0_outputs(9705));
    outputs(5256) <= (layer0_outputs(149)) xor (layer0_outputs(4071));
    outputs(5257) <= not(layer0_outputs(4749));
    outputs(5258) <= not((layer0_outputs(7582)) xor (layer0_outputs(1122)));
    outputs(5259) <= not((layer0_outputs(90)) xor (layer0_outputs(10223)));
    outputs(5260) <= not(layer0_outputs(2436));
    outputs(5261) <= (layer0_outputs(3274)) xor (layer0_outputs(2742));
    outputs(5262) <= (layer0_outputs(2413)) xor (layer0_outputs(8574));
    outputs(5263) <= not((layer0_outputs(6644)) xor (layer0_outputs(2274)));
    outputs(5264) <= not(layer0_outputs(7260));
    outputs(5265) <= not(layer0_outputs(4379));
    outputs(5266) <= not(layer0_outputs(8418));
    outputs(5267) <= layer0_outputs(8582);
    outputs(5268) <= (layer0_outputs(9099)) and (layer0_outputs(7493));
    outputs(5269) <= not((layer0_outputs(8131)) and (layer0_outputs(784)));
    outputs(5270) <= layer0_outputs(2610);
    outputs(5271) <= (layer0_outputs(2362)) and (layer0_outputs(1091));
    outputs(5272) <= (layer0_outputs(4625)) xor (layer0_outputs(5622));
    outputs(5273) <= not((layer0_outputs(8440)) xor (layer0_outputs(9394)));
    outputs(5274) <= not(layer0_outputs(3493)) or (layer0_outputs(7051));
    outputs(5275) <= (layer0_outputs(9693)) and not (layer0_outputs(9022));
    outputs(5276) <= (layer0_outputs(5058)) and not (layer0_outputs(33));
    outputs(5277) <= layer0_outputs(5305);
    outputs(5278) <= (layer0_outputs(6463)) and (layer0_outputs(272));
    outputs(5279) <= layer0_outputs(3180);
    outputs(5280) <= (layer0_outputs(8858)) xor (layer0_outputs(6308));
    outputs(5281) <= not(layer0_outputs(7952));
    outputs(5282) <= (layer0_outputs(7421)) and (layer0_outputs(9197));
    outputs(5283) <= layer0_outputs(8736);
    outputs(5284) <= not(layer0_outputs(5094));
    outputs(5285) <= layer0_outputs(1298);
    outputs(5286) <= not((layer0_outputs(119)) xor (layer0_outputs(5908)));
    outputs(5287) <= not(layer0_outputs(8780));
    outputs(5288) <= not((layer0_outputs(3314)) xor (layer0_outputs(4343)));
    outputs(5289) <= (layer0_outputs(859)) and (layer0_outputs(660));
    outputs(5290) <= not((layer0_outputs(3164)) or (layer0_outputs(1699)));
    outputs(5291) <= not((layer0_outputs(1723)) xor (layer0_outputs(9907)));
    outputs(5292) <= not(layer0_outputs(9659)) or (layer0_outputs(9283));
    outputs(5293) <= layer0_outputs(1256);
    outputs(5294) <= not(layer0_outputs(4777));
    outputs(5295) <= not(layer0_outputs(3906)) or (layer0_outputs(9442));
    outputs(5296) <= not((layer0_outputs(6880)) xor (layer0_outputs(4133)));
    outputs(5297) <= layer0_outputs(3010);
    outputs(5298) <= not(layer0_outputs(5998));
    outputs(5299) <= not((layer0_outputs(4900)) xor (layer0_outputs(5169)));
    outputs(5300) <= not((layer0_outputs(7372)) and (layer0_outputs(3307)));
    outputs(5301) <= layer0_outputs(2146);
    outputs(5302) <= layer0_outputs(776);
    outputs(5303) <= layer0_outputs(2591);
    outputs(5304) <= not((layer0_outputs(873)) xor (layer0_outputs(7829)));
    outputs(5305) <= not(layer0_outputs(5503));
    outputs(5306) <= layer0_outputs(2360);
    outputs(5307) <= (layer0_outputs(3667)) xor (layer0_outputs(9954));
    outputs(5308) <= (layer0_outputs(4767)) xor (layer0_outputs(10044));
    outputs(5309) <= layer0_outputs(6242);
    outputs(5310) <= (layer0_outputs(1678)) xor (layer0_outputs(2013));
    outputs(5311) <= not(layer0_outputs(5761));
    outputs(5312) <= (layer0_outputs(5268)) xor (layer0_outputs(10009));
    outputs(5313) <= layer0_outputs(9478);
    outputs(5314) <= (layer0_outputs(935)) xor (layer0_outputs(613));
    outputs(5315) <= layer0_outputs(4031);
    outputs(5316) <= not(layer0_outputs(8289));
    outputs(5317) <= not((layer0_outputs(6271)) xor (layer0_outputs(3224)));
    outputs(5318) <= not((layer0_outputs(1902)) xor (layer0_outputs(7429)));
    outputs(5319) <= layer0_outputs(4015);
    outputs(5320) <= layer0_outputs(5328);
    outputs(5321) <= not(layer0_outputs(2854));
    outputs(5322) <= not(layer0_outputs(9892));
    outputs(5323) <= layer0_outputs(8835);
    outputs(5324) <= not((layer0_outputs(5704)) or (layer0_outputs(8310)));
    outputs(5325) <= layer0_outputs(9314);
    outputs(5326) <= (layer0_outputs(43)) xor (layer0_outputs(5085));
    outputs(5327) <= (layer0_outputs(7901)) xor (layer0_outputs(2246));
    outputs(5328) <= layer0_outputs(5867);
    outputs(5329) <= (layer0_outputs(6917)) xor (layer0_outputs(9369));
    outputs(5330) <= (layer0_outputs(7629)) xor (layer0_outputs(2914));
    outputs(5331) <= not((layer0_outputs(539)) and (layer0_outputs(5442)));
    outputs(5332) <= not(layer0_outputs(3704));
    outputs(5333) <= not((layer0_outputs(4472)) and (layer0_outputs(5506)));
    outputs(5334) <= not((layer0_outputs(5989)) xor (layer0_outputs(5866)));
    outputs(5335) <= (layer0_outputs(1600)) xor (layer0_outputs(1028));
    outputs(5336) <= (layer0_outputs(2666)) and not (layer0_outputs(9450));
    outputs(5337) <= not((layer0_outputs(701)) or (layer0_outputs(7639)));
    outputs(5338) <= (layer0_outputs(8028)) and (layer0_outputs(7518));
    outputs(5339) <= layer0_outputs(2420);
    outputs(5340) <= not(layer0_outputs(809));
    outputs(5341) <= not(layer0_outputs(2714));
    outputs(5342) <= not(layer0_outputs(5187));
    outputs(5343) <= layer0_outputs(5900);
    outputs(5344) <= (layer0_outputs(2385)) xor (layer0_outputs(80));
    outputs(5345) <= not(layer0_outputs(7237));
    outputs(5346) <= not(layer0_outputs(5110));
    outputs(5347) <= layer0_outputs(7645);
    outputs(5348) <= not(layer0_outputs(7267));
    outputs(5349) <= (layer0_outputs(7856)) and not (layer0_outputs(2983));
    outputs(5350) <= layer0_outputs(9447);
    outputs(5351) <= layer0_outputs(8928);
    outputs(5352) <= not(layer0_outputs(7615));
    outputs(5353) <= not((layer0_outputs(5419)) xor (layer0_outputs(4763)));
    outputs(5354) <= layer0_outputs(6674);
    outputs(5355) <= not((layer0_outputs(3693)) or (layer0_outputs(8644)));
    outputs(5356) <= (layer0_outputs(9218)) and not (layer0_outputs(8323));
    outputs(5357) <= (layer0_outputs(4201)) xor (layer0_outputs(4992));
    outputs(5358) <= layer0_outputs(8633);
    outputs(5359) <= layer0_outputs(5242);
    outputs(5360) <= not((layer0_outputs(5424)) xor (layer0_outputs(6064)));
    outputs(5361) <= (layer0_outputs(2884)) xor (layer0_outputs(8729));
    outputs(5362) <= not(layer0_outputs(4847));
    outputs(5363) <= not((layer0_outputs(7950)) or (layer0_outputs(3048)));
    outputs(5364) <= not((layer0_outputs(6240)) xor (layer0_outputs(5164)));
    outputs(5365) <= layer0_outputs(7680);
    outputs(5366) <= (layer0_outputs(9262)) xor (layer0_outputs(1779));
    outputs(5367) <= not((layer0_outputs(9317)) and (layer0_outputs(8668)));
    outputs(5368) <= (layer0_outputs(3462)) and not (layer0_outputs(2162));
    outputs(5369) <= layer0_outputs(6745);
    outputs(5370) <= layer0_outputs(1988);
    outputs(5371) <= not(layer0_outputs(4404));
    outputs(5372) <= not((layer0_outputs(9737)) xor (layer0_outputs(8994)));
    outputs(5373) <= (layer0_outputs(8007)) or (layer0_outputs(9258));
    outputs(5374) <= not((layer0_outputs(5531)) and (layer0_outputs(9203)));
    outputs(5375) <= not(layer0_outputs(8519));
    outputs(5376) <= not((layer0_outputs(9636)) xor (layer0_outputs(5464)));
    outputs(5377) <= (layer0_outputs(9945)) xor (layer0_outputs(4579));
    outputs(5378) <= (layer0_outputs(8350)) and (layer0_outputs(7891));
    outputs(5379) <= not((layer0_outputs(5741)) xor (layer0_outputs(7863)));
    outputs(5380) <= not(layer0_outputs(9839));
    outputs(5381) <= not((layer0_outputs(7160)) and (layer0_outputs(3306)));
    outputs(5382) <= not(layer0_outputs(9141));
    outputs(5383) <= (layer0_outputs(2688)) and not (layer0_outputs(2871));
    outputs(5384) <= not((layer0_outputs(8128)) xor (layer0_outputs(6117)));
    outputs(5385) <= not(layer0_outputs(631)) or (layer0_outputs(1247));
    outputs(5386) <= layer0_outputs(4036);
    outputs(5387) <= (layer0_outputs(6886)) xor (layer0_outputs(9061));
    outputs(5388) <= not((layer0_outputs(6167)) xor (layer0_outputs(3514)));
    outputs(5389) <= layer0_outputs(6955);
    outputs(5390) <= not(layer0_outputs(435)) or (layer0_outputs(3602));
    outputs(5391) <= not((layer0_outputs(6064)) or (layer0_outputs(7517)));
    outputs(5392) <= not(layer0_outputs(3394));
    outputs(5393) <= not(layer0_outputs(5432));
    outputs(5394) <= not((layer0_outputs(2130)) xor (layer0_outputs(437)));
    outputs(5395) <= not(layer0_outputs(3003)) or (layer0_outputs(9297));
    outputs(5396) <= not(layer0_outputs(9143));
    outputs(5397) <= not((layer0_outputs(5579)) xor (layer0_outputs(2092)));
    outputs(5398) <= layer0_outputs(1832);
    outputs(5399) <= layer0_outputs(3059);
    outputs(5400) <= (layer0_outputs(6503)) and not (layer0_outputs(9167));
    outputs(5401) <= (layer0_outputs(7550)) and (layer0_outputs(4242));
    outputs(5402) <= layer0_outputs(1596);
    outputs(5403) <= layer0_outputs(140);
    outputs(5404) <= not(layer0_outputs(1586));
    outputs(5405) <= not(layer0_outputs(4658)) or (layer0_outputs(2575));
    outputs(5406) <= not(layer0_outputs(7));
    outputs(5407) <= layer0_outputs(2452);
    outputs(5408) <= (layer0_outputs(8151)) xor (layer0_outputs(10157));
    outputs(5409) <= (layer0_outputs(9946)) xor (layer0_outputs(8090));
    outputs(5410) <= layer0_outputs(7347);
    outputs(5411) <= not(layer0_outputs(3560));
    outputs(5412) <= (layer0_outputs(4846)) xor (layer0_outputs(9462));
    outputs(5413) <= not(layer0_outputs(2320));
    outputs(5414) <= not((layer0_outputs(9817)) xor (layer0_outputs(8476)));
    outputs(5415) <= not(layer0_outputs(8148));
    outputs(5416) <= (layer0_outputs(7252)) xor (layer0_outputs(7979));
    outputs(5417) <= not(layer0_outputs(8711)) or (layer0_outputs(1132));
    outputs(5418) <= (layer0_outputs(3694)) and (layer0_outputs(7113));
    outputs(5419) <= not((layer0_outputs(457)) xor (layer0_outputs(7604)));
    outputs(5420) <= not(layer0_outputs(2801));
    outputs(5421) <= not((layer0_outputs(7004)) xor (layer0_outputs(204)));
    outputs(5422) <= layer0_outputs(10049);
    outputs(5423) <= not((layer0_outputs(4501)) xor (layer0_outputs(2029)));
    outputs(5424) <= not(layer0_outputs(289));
    outputs(5425) <= not(layer0_outputs(1819));
    outputs(5426) <= (layer0_outputs(8142)) or (layer0_outputs(1087));
    outputs(5427) <= not(layer0_outputs(9863)) or (layer0_outputs(2550));
    outputs(5428) <= (layer0_outputs(1705)) xor (layer0_outputs(8214));
    outputs(5429) <= not((layer0_outputs(9484)) xor (layer0_outputs(8500)));
    outputs(5430) <= not(layer0_outputs(7803));
    outputs(5431) <= (layer0_outputs(9776)) xor (layer0_outputs(8294));
    outputs(5432) <= not(layer0_outputs(7653));
    outputs(5433) <= (layer0_outputs(3864)) and not (layer0_outputs(3720));
    outputs(5434) <= not(layer0_outputs(3596)) or (layer0_outputs(2683));
    outputs(5435) <= layer0_outputs(4585);
    outputs(5436) <= (layer0_outputs(4456)) xor (layer0_outputs(6903));
    outputs(5437) <= not(layer0_outputs(5747));
    outputs(5438) <= not(layer0_outputs(1859));
    outputs(5439) <= (layer0_outputs(8411)) xor (layer0_outputs(5378));
    outputs(5440) <= (layer0_outputs(1082)) xor (layer0_outputs(2261));
    outputs(5441) <= (layer0_outputs(5349)) and (layer0_outputs(4718));
    outputs(5442) <= (layer0_outputs(3606)) xor (layer0_outputs(9012));
    outputs(5443) <= layer0_outputs(8547);
    outputs(5444) <= layer0_outputs(1854);
    outputs(5445) <= not(layer0_outputs(9557));
    outputs(5446) <= (layer0_outputs(3696)) xor (layer0_outputs(5581));
    outputs(5447) <= layer0_outputs(1430);
    outputs(5448) <= not((layer0_outputs(2807)) xor (layer0_outputs(9899)));
    outputs(5449) <= (layer0_outputs(7779)) and not (layer0_outputs(5997));
    outputs(5450) <= not(layer0_outputs(6714));
    outputs(5451) <= not(layer0_outputs(9944));
    outputs(5452) <= layer0_outputs(4088);
    outputs(5453) <= (layer0_outputs(7422)) and not (layer0_outputs(4961));
    outputs(5454) <= not(layer0_outputs(6135));
    outputs(5455) <= layer0_outputs(1086);
    outputs(5456) <= not(layer0_outputs(10198));
    outputs(5457) <= layer0_outputs(2882);
    outputs(5458) <= not((layer0_outputs(4633)) xor (layer0_outputs(4372)));
    outputs(5459) <= not(layer0_outputs(1473));
    outputs(5460) <= not((layer0_outputs(5400)) and (layer0_outputs(436)));
    outputs(5461) <= layer0_outputs(551);
    outputs(5462) <= not(layer0_outputs(9462));
    outputs(5463) <= not(layer0_outputs(6575)) or (layer0_outputs(4115));
    outputs(5464) <= layer0_outputs(8538);
    outputs(5465) <= not((layer0_outputs(4239)) xor (layer0_outputs(9557)));
    outputs(5466) <= not(layer0_outputs(3040));
    outputs(5467) <= not((layer0_outputs(4348)) xor (layer0_outputs(7552)));
    outputs(5468) <= not((layer0_outputs(8057)) xor (layer0_outputs(6378)));
    outputs(5469) <= (layer0_outputs(6726)) and not (layer0_outputs(3052));
    outputs(5470) <= not(layer0_outputs(365));
    outputs(5471) <= (layer0_outputs(9090)) xor (layer0_outputs(425));
    outputs(5472) <= layer0_outputs(1107);
    outputs(5473) <= not(layer0_outputs(3566));
    outputs(5474) <= not((layer0_outputs(1810)) xor (layer0_outputs(1269)));
    outputs(5475) <= (layer0_outputs(1845)) and not (layer0_outputs(1572));
    outputs(5476) <= (layer0_outputs(2199)) and not (layer0_outputs(1763));
    outputs(5477) <= not((layer0_outputs(378)) xor (layer0_outputs(4429)));
    outputs(5478) <= (layer0_outputs(4674)) xor (layer0_outputs(4268));
    outputs(5479) <= not((layer0_outputs(8908)) xor (layer0_outputs(8915)));
    outputs(5480) <= not((layer0_outputs(863)) xor (layer0_outputs(10156)));
    outputs(5481) <= not((layer0_outputs(10211)) or (layer0_outputs(6861)));
    outputs(5482) <= not((layer0_outputs(2086)) xor (layer0_outputs(3318)));
    outputs(5483) <= layer0_outputs(9797);
    outputs(5484) <= layer0_outputs(6238);
    outputs(5485) <= layer0_outputs(423);
    outputs(5486) <= layer0_outputs(7811);
    outputs(5487) <= not((layer0_outputs(5808)) xor (layer0_outputs(1930)));
    outputs(5488) <= not((layer0_outputs(3101)) xor (layer0_outputs(4464)));
    outputs(5489) <= (layer0_outputs(7185)) xor (layer0_outputs(4476));
    outputs(5490) <= not(layer0_outputs(888));
    outputs(5491) <= not(layer0_outputs(4439));
    outputs(5492) <= (layer0_outputs(5931)) and not (layer0_outputs(2863));
    outputs(5493) <= not(layer0_outputs(3796));
    outputs(5494) <= not(layer0_outputs(1910));
    outputs(5495) <= (layer0_outputs(8330)) xor (layer0_outputs(9191));
    outputs(5496) <= not(layer0_outputs(6814));
    outputs(5497) <= (layer0_outputs(5226)) and not (layer0_outputs(6196));
    outputs(5498) <= layer0_outputs(5846);
    outputs(5499) <= (layer0_outputs(5114)) or (layer0_outputs(1998));
    outputs(5500) <= not((layer0_outputs(5055)) and (layer0_outputs(271)));
    outputs(5501) <= not(layer0_outputs(1748));
    outputs(5502) <= (layer0_outputs(6424)) and not (layer0_outputs(3002));
    outputs(5503) <= (layer0_outputs(10024)) xor (layer0_outputs(810));
    outputs(5504) <= not((layer0_outputs(4649)) xor (layer0_outputs(755)));
    outputs(5505) <= (layer0_outputs(1409)) xor (layer0_outputs(8824));
    outputs(5506) <= not((layer0_outputs(9264)) or (layer0_outputs(6016)));
    outputs(5507) <= not(layer0_outputs(4092));
    outputs(5508) <= layer0_outputs(1008);
    outputs(5509) <= not(layer0_outputs(3673));
    outputs(5510) <= (layer0_outputs(3432)) and not (layer0_outputs(6072));
    outputs(5511) <= layer0_outputs(5499);
    outputs(5512) <= layer0_outputs(1446);
    outputs(5513) <= (layer0_outputs(3441)) or (layer0_outputs(8758));
    outputs(5514) <= (layer0_outputs(6924)) and not (layer0_outputs(1171));
    outputs(5515) <= layer0_outputs(5537);
    outputs(5516) <= (layer0_outputs(133)) xor (layer0_outputs(7482));
    outputs(5517) <= not((layer0_outputs(6279)) xor (layer0_outputs(2377)));
    outputs(5518) <= not((layer0_outputs(9810)) or (layer0_outputs(9380)));
    outputs(5519) <= not((layer0_outputs(8701)) xor (layer0_outputs(1984)));
    outputs(5520) <= layer0_outputs(1334);
    outputs(5521) <= not((layer0_outputs(8193)) xor (layer0_outputs(8896)));
    outputs(5522) <= not((layer0_outputs(2580)) xor (layer0_outputs(9036)));
    outputs(5523) <= layer0_outputs(1120);
    outputs(5524) <= not((layer0_outputs(9198)) or (layer0_outputs(2979)));
    outputs(5525) <= not(layer0_outputs(6760)) or (layer0_outputs(9654));
    outputs(5526) <= layer0_outputs(10239);
    outputs(5527) <= (layer0_outputs(1235)) xor (layer0_outputs(8706));
    outputs(5528) <= (layer0_outputs(1235)) xor (layer0_outputs(4853));
    outputs(5529) <= (layer0_outputs(488)) xor (layer0_outputs(6476));
    outputs(5530) <= (layer0_outputs(377)) xor (layer0_outputs(3272));
    outputs(5531) <= not(layer0_outputs(9070));
    outputs(5532) <= not(layer0_outputs(9393));
    outputs(5533) <= layer0_outputs(7776);
    outputs(5534) <= layer0_outputs(9374);
    outputs(5535) <= not(layer0_outputs(3098));
    outputs(5536) <= not(layer0_outputs(9115));
    outputs(5537) <= not(layer0_outputs(1311)) or (layer0_outputs(1581));
    outputs(5538) <= not(layer0_outputs(921)) or (layer0_outputs(3153));
    outputs(5539) <= not(layer0_outputs(7280));
    outputs(5540) <= (layer0_outputs(7809)) xor (layer0_outputs(485));
    outputs(5541) <= not((layer0_outputs(9207)) or (layer0_outputs(9922)));
    outputs(5542) <= not(layer0_outputs(10214));
    outputs(5543) <= (layer0_outputs(3066)) xor (layer0_outputs(907));
    outputs(5544) <= layer0_outputs(7751);
    outputs(5545) <= (layer0_outputs(4378)) xor (layer0_outputs(6940));
    outputs(5546) <= not(layer0_outputs(5080)) or (layer0_outputs(9941));
    outputs(5547) <= not((layer0_outputs(1577)) xor (layer0_outputs(6936)));
    outputs(5548) <= not((layer0_outputs(5929)) or (layer0_outputs(2357)));
    outputs(5549) <= (layer0_outputs(5152)) and not (layer0_outputs(675));
    outputs(5550) <= (layer0_outputs(1453)) and not (layer0_outputs(8705));
    outputs(5551) <= not(layer0_outputs(339)) or (layer0_outputs(6471));
    outputs(5552) <= not(layer0_outputs(8241));
    outputs(5553) <= not(layer0_outputs(5623));
    outputs(5554) <= not(layer0_outputs(5342));
    outputs(5555) <= (layer0_outputs(8333)) and not (layer0_outputs(3524));
    outputs(5556) <= not((layer0_outputs(7361)) xor (layer0_outputs(2822)));
    outputs(5557) <= not((layer0_outputs(3312)) xor (layer0_outputs(7087)));
    outputs(5558) <= not(layer0_outputs(3912));
    outputs(5559) <= layer0_outputs(7113);
    outputs(5560) <= not((layer0_outputs(5566)) xor (layer0_outputs(6232)));
    outputs(5561) <= layer0_outputs(2331);
    outputs(5562) <= (layer0_outputs(146)) xor (layer0_outputs(8515));
    outputs(5563) <= layer0_outputs(8641);
    outputs(5564) <= not(layer0_outputs(6968));
    outputs(5565) <= not(layer0_outputs(9444));
    outputs(5566) <= layer0_outputs(7578);
    outputs(5567) <= not(layer0_outputs(5092));
    outputs(5568) <= not(layer0_outputs(9202));
    outputs(5569) <= (layer0_outputs(7510)) and not (layer0_outputs(1585));
    outputs(5570) <= not((layer0_outputs(3060)) or (layer0_outputs(1366)));
    outputs(5571) <= layer0_outputs(6185);
    outputs(5572) <= not((layer0_outputs(8005)) xor (layer0_outputs(3632)));
    outputs(5573) <= (layer0_outputs(7589)) and (layer0_outputs(3091));
    outputs(5574) <= not((layer0_outputs(9186)) xor (layer0_outputs(1462)));
    outputs(5575) <= layer0_outputs(2980);
    outputs(5576) <= not((layer0_outputs(609)) xor (layer0_outputs(5717)));
    outputs(5577) <= not((layer0_outputs(3400)) xor (layer0_outputs(8082)));
    outputs(5578) <= not(layer0_outputs(7356));
    outputs(5579) <= not(layer0_outputs(4848));
    outputs(5580) <= layer0_outputs(3504);
    outputs(5581) <= (layer0_outputs(1245)) and not (layer0_outputs(9209));
    outputs(5582) <= (layer0_outputs(7456)) and (layer0_outputs(1940));
    outputs(5583) <= not(layer0_outputs(252)) or (layer0_outputs(4853));
    outputs(5584) <= layer0_outputs(8645);
    outputs(5585) <= (layer0_outputs(8400)) xor (layer0_outputs(7515));
    outputs(5586) <= (layer0_outputs(2571)) and not (layer0_outputs(8781));
    outputs(5587) <= (layer0_outputs(6233)) xor (layer0_outputs(3259));
    outputs(5588) <= layer0_outputs(1997);
    outputs(5589) <= not(layer0_outputs(2866));
    outputs(5590) <= (layer0_outputs(5661)) and not (layer0_outputs(364));
    outputs(5591) <= (layer0_outputs(466)) and (layer0_outputs(5691));
    outputs(5592) <= not((layer0_outputs(4369)) xor (layer0_outputs(6460)));
    outputs(5593) <= not((layer0_outputs(844)) xor (layer0_outputs(9329)));
    outputs(5594) <= (layer0_outputs(8507)) xor (layer0_outputs(1850));
    outputs(5595) <= (layer0_outputs(182)) xor (layer0_outputs(3457));
    outputs(5596) <= not((layer0_outputs(1265)) xor (layer0_outputs(2167)));
    outputs(5597) <= (layer0_outputs(6739)) and not (layer0_outputs(5626));
    outputs(5598) <= layer0_outputs(9089);
    outputs(5599) <= layer0_outputs(1518);
    outputs(5600) <= not(layer0_outputs(6391));
    outputs(5601) <= (layer0_outputs(1968)) or (layer0_outputs(3167));
    outputs(5602) <= layer0_outputs(5801);
    outputs(5603) <= not(layer0_outputs(6953)) or (layer0_outputs(9492));
    outputs(5604) <= (layer0_outputs(5059)) or (layer0_outputs(5740));
    outputs(5605) <= not((layer0_outputs(3896)) xor (layer0_outputs(9864)));
    outputs(5606) <= layer0_outputs(1296);
    outputs(5607) <= not(layer0_outputs(6925)) or (layer0_outputs(6039));
    outputs(5608) <= layer0_outputs(9940);
    outputs(5609) <= not((layer0_outputs(3038)) xor (layer0_outputs(606)));
    outputs(5610) <= layer0_outputs(2101);
    outputs(5611) <= not((layer0_outputs(22)) and (layer0_outputs(697)));
    outputs(5612) <= not((layer0_outputs(10137)) and (layer0_outputs(6844)));
    outputs(5613) <= not((layer0_outputs(4767)) xor (layer0_outputs(754)));
    outputs(5614) <= layer0_outputs(5425);
    outputs(5615) <= not((layer0_outputs(5643)) xor (layer0_outputs(4116)));
    outputs(5616) <= layer0_outputs(4076);
    outputs(5617) <= layer0_outputs(6763);
    outputs(5618) <= not((layer0_outputs(9535)) or (layer0_outputs(2118)));
    outputs(5619) <= not(layer0_outputs(4606));
    outputs(5620) <= not(layer0_outputs(5904));
    outputs(5621) <= (layer0_outputs(2835)) xor (layer0_outputs(3049));
    outputs(5622) <= (layer0_outputs(4371)) and not (layer0_outputs(8146));
    outputs(5623) <= (layer0_outputs(6325)) or (layer0_outputs(4070));
    outputs(5624) <= layer0_outputs(9891);
    outputs(5625) <= not(layer0_outputs(2553)) or (layer0_outputs(7645));
    outputs(5626) <= layer0_outputs(6594);
    outputs(5627) <= not(layer0_outputs(8351)) or (layer0_outputs(1432));
    outputs(5628) <= layer0_outputs(1330);
    outputs(5629) <= not(layer0_outputs(9296));
    outputs(5630) <= not(layer0_outputs(2425));
    outputs(5631) <= not((layer0_outputs(5560)) xor (layer0_outputs(3109)));
    outputs(5632) <= not((layer0_outputs(5864)) xor (layer0_outputs(4165)));
    outputs(5633) <= not((layer0_outputs(8272)) xor (layer0_outputs(1174)));
    outputs(5634) <= (layer0_outputs(704)) xor (layer0_outputs(6194));
    outputs(5635) <= not((layer0_outputs(10158)) xor (layer0_outputs(4561)));
    outputs(5636) <= not((layer0_outputs(5934)) xor (layer0_outputs(6111)));
    outputs(5637) <= not((layer0_outputs(4258)) and (layer0_outputs(4879)));
    outputs(5638) <= not((layer0_outputs(4261)) xor (layer0_outputs(5881)));
    outputs(5639) <= not(layer0_outputs(2067));
    outputs(5640) <= not(layer0_outputs(1673)) or (layer0_outputs(73));
    outputs(5641) <= not((layer0_outputs(8167)) xor (layer0_outputs(6619)));
    outputs(5642) <= layer0_outputs(5112);
    outputs(5643) <= not((layer0_outputs(64)) xor (layer0_outputs(6193)));
    outputs(5644) <= (layer0_outputs(2015)) or (layer0_outputs(39));
    outputs(5645) <= (layer0_outputs(5427)) xor (layer0_outputs(3568));
    outputs(5646) <= (layer0_outputs(4385)) xor (layer0_outputs(9016));
    outputs(5647) <= not(layer0_outputs(6911));
    outputs(5648) <= not(layer0_outputs(2963)) or (layer0_outputs(8989));
    outputs(5649) <= not(layer0_outputs(5592));
    outputs(5650) <= not(layer0_outputs(10013));
    outputs(5651) <= (layer0_outputs(7364)) and not (layer0_outputs(5715));
    outputs(5652) <= not((layer0_outputs(565)) xor (layer0_outputs(3682)));
    outputs(5653) <= not(layer0_outputs(9186));
    outputs(5654) <= not((layer0_outputs(8371)) or (layer0_outputs(2069)));
    outputs(5655) <= (layer0_outputs(3745)) xor (layer0_outputs(9458));
    outputs(5656) <= not(layer0_outputs(4384));
    outputs(5657) <= (layer0_outputs(7270)) xor (layer0_outputs(4551));
    outputs(5658) <= not(layer0_outputs(7273));
    outputs(5659) <= (layer0_outputs(5397)) and not (layer0_outputs(5117));
    outputs(5660) <= not(layer0_outputs(5375)) or (layer0_outputs(1220));
    outputs(5661) <= not(layer0_outputs(2821));
    outputs(5662) <= (layer0_outputs(3236)) and not (layer0_outputs(133));
    outputs(5663) <= not(layer0_outputs(2192));
    outputs(5664) <= not(layer0_outputs(6056));
    outputs(5665) <= (layer0_outputs(9144)) xor (layer0_outputs(2248));
    outputs(5666) <= not(layer0_outputs(244));
    outputs(5667) <= layer0_outputs(9511);
    outputs(5668) <= layer0_outputs(206);
    outputs(5669) <= not((layer0_outputs(7833)) and (layer0_outputs(6390)));
    outputs(5670) <= not(layer0_outputs(2935));
    outputs(5671) <= (layer0_outputs(3787)) or (layer0_outputs(4786));
    outputs(5672) <= not((layer0_outputs(8432)) xor (layer0_outputs(9193)));
    outputs(5673) <= not(layer0_outputs(3530));
    outputs(5674) <= not(layer0_outputs(8831));
    outputs(5675) <= not(layer0_outputs(6533));
    outputs(5676) <= layer0_outputs(6725);
    outputs(5677) <= (layer0_outputs(4125)) xor (layer0_outputs(1200));
    outputs(5678) <= layer0_outputs(7168);
    outputs(5679) <= not(layer0_outputs(1074));
    outputs(5680) <= (layer0_outputs(2774)) xor (layer0_outputs(5073));
    outputs(5681) <= (layer0_outputs(6821)) or (layer0_outputs(7314));
    outputs(5682) <= not(layer0_outputs(8185));
    outputs(5683) <= (layer0_outputs(9401)) xor (layer0_outputs(7618));
    outputs(5684) <= not(layer0_outputs(7890)) or (layer0_outputs(7892));
    outputs(5685) <= (layer0_outputs(4371)) and (layer0_outputs(4242));
    outputs(5686) <= (layer0_outputs(3996)) and not (layer0_outputs(9173));
    outputs(5687) <= not((layer0_outputs(8913)) xor (layer0_outputs(9133)));
    outputs(5688) <= layer0_outputs(5457);
    outputs(5689) <= (layer0_outputs(5327)) or (layer0_outputs(3942));
    outputs(5690) <= not(layer0_outputs(10218));
    outputs(5691) <= (layer0_outputs(4190)) xor (layer0_outputs(598));
    outputs(5692) <= not((layer0_outputs(6249)) xor (layer0_outputs(2143)));
    outputs(5693) <= (layer0_outputs(4412)) xor (layer0_outputs(4097));
    outputs(5694) <= not((layer0_outputs(934)) or (layer0_outputs(6110)));
    outputs(5695) <= (layer0_outputs(2414)) xor (layer0_outputs(736));
    outputs(5696) <= not(layer0_outputs(1725));
    outputs(5697) <= layer0_outputs(2724);
    outputs(5698) <= not((layer0_outputs(6029)) xor (layer0_outputs(5370)));
    outputs(5699) <= (layer0_outputs(9698)) and (layer0_outputs(4757));
    outputs(5700) <= (layer0_outputs(5362)) and (layer0_outputs(8411));
    outputs(5701) <= not(layer0_outputs(4631)) or (layer0_outputs(10042));
    outputs(5702) <= (layer0_outputs(924)) xor (layer0_outputs(2159));
    outputs(5703) <= not((layer0_outputs(6858)) or (layer0_outputs(2429)));
    outputs(5704) <= not((layer0_outputs(4419)) or (layer0_outputs(988)));
    outputs(5705) <= not((layer0_outputs(9365)) xor (layer0_outputs(3741)));
    outputs(5706) <= not(layer0_outputs(3164));
    outputs(5707) <= not((layer0_outputs(9248)) xor (layer0_outputs(3264)));
    outputs(5708) <= (layer0_outputs(4498)) xor (layer0_outputs(7619));
    outputs(5709) <= layer0_outputs(3554);
    outputs(5710) <= (layer0_outputs(1845)) and (layer0_outputs(8910));
    outputs(5711) <= (layer0_outputs(7563)) xor (layer0_outputs(4700));
    outputs(5712) <= not((layer0_outputs(6318)) xor (layer0_outputs(5611)));
    outputs(5713) <= not((layer0_outputs(8664)) xor (layer0_outputs(2993)));
    outputs(5714) <= not(layer0_outputs(9651));
    outputs(5715) <= layer0_outputs(4350);
    outputs(5716) <= not((layer0_outputs(126)) and (layer0_outputs(950)));
    outputs(5717) <= not((layer0_outputs(9422)) xor (layer0_outputs(839)));
    outputs(5718) <= not(layer0_outputs(6208));
    outputs(5719) <= (layer0_outputs(2030)) xor (layer0_outputs(6641));
    outputs(5720) <= layer0_outputs(2426);
    outputs(5721) <= layer0_outputs(2862);
    outputs(5722) <= (layer0_outputs(943)) and (layer0_outputs(7749));
    outputs(5723) <= not(layer0_outputs(6501));
    outputs(5724) <= not((layer0_outputs(9299)) xor (layer0_outputs(1442)));
    outputs(5725) <= not(layer0_outputs(2876));
    outputs(5726) <= layer0_outputs(424);
    outputs(5727) <= (layer0_outputs(3448)) xor (layer0_outputs(6423));
    outputs(5728) <= (layer0_outputs(2092)) xor (layer0_outputs(2502));
    outputs(5729) <= (layer0_outputs(1754)) or (layer0_outputs(9645));
    outputs(5730) <= not((layer0_outputs(4711)) xor (layer0_outputs(2887)));
    outputs(5731) <= (layer0_outputs(8244)) xor (layer0_outputs(903));
    outputs(5732) <= layer0_outputs(5212);
    outputs(5733) <= not((layer0_outputs(8178)) or (layer0_outputs(3438)));
    outputs(5734) <= (layer0_outputs(4554)) and not (layer0_outputs(5491));
    outputs(5735) <= not((layer0_outputs(1721)) xor (layer0_outputs(6555)));
    outputs(5736) <= (layer0_outputs(9527)) and not (layer0_outputs(4933));
    outputs(5737) <= not(layer0_outputs(7059)) or (layer0_outputs(4807));
    outputs(5738) <= '0';
    outputs(5739) <= layer0_outputs(2372);
    outputs(5740) <= not((layer0_outputs(7234)) xor (layer0_outputs(4950)));
    outputs(5741) <= not(layer0_outputs(4207));
    outputs(5742) <= not(layer0_outputs(3687)) or (layer0_outputs(4910));
    outputs(5743) <= not(layer0_outputs(6382));
    outputs(5744) <= layer0_outputs(5564);
    outputs(5745) <= not(layer0_outputs(10175));
    outputs(5746) <= not(layer0_outputs(5891)) or (layer0_outputs(4018));
    outputs(5747) <= (layer0_outputs(9886)) and (layer0_outputs(5861));
    outputs(5748) <= layer0_outputs(4515);
    outputs(5749) <= (layer0_outputs(913)) xor (layer0_outputs(3054));
    outputs(5750) <= layer0_outputs(3103);
    outputs(5751) <= (layer0_outputs(10139)) xor (layer0_outputs(9991));
    outputs(5752) <= not(layer0_outputs(8761));
    outputs(5753) <= not((layer0_outputs(7720)) xor (layer0_outputs(5751)));
    outputs(5754) <= layer0_outputs(9080);
    outputs(5755) <= not((layer0_outputs(9806)) or (layer0_outputs(9783)));
    outputs(5756) <= layer0_outputs(86);
    outputs(5757) <= layer0_outputs(1451);
    outputs(5758) <= not(layer0_outputs(1050));
    outputs(5759) <= not((layer0_outputs(1504)) xor (layer0_outputs(962)));
    outputs(5760) <= layer0_outputs(1507);
    outputs(5761) <= not((layer0_outputs(7019)) or (layer0_outputs(8750)));
    outputs(5762) <= layer0_outputs(1520);
    outputs(5763) <= (layer0_outputs(10234)) or (layer0_outputs(5578));
    outputs(5764) <= not((layer0_outputs(7844)) xor (layer0_outputs(1346)));
    outputs(5765) <= not((layer0_outputs(2102)) xor (layer0_outputs(4568)));
    outputs(5766) <= not((layer0_outputs(4804)) xor (layer0_outputs(8820)));
    outputs(5767) <= not(layer0_outputs(6437));
    outputs(5768) <= layer0_outputs(5591);
    outputs(5769) <= not((layer0_outputs(9955)) and (layer0_outputs(4651)));
    outputs(5770) <= (layer0_outputs(7272)) xor (layer0_outputs(1585));
    outputs(5771) <= layer0_outputs(5215);
    outputs(5772) <= (layer0_outputs(1270)) xor (layer0_outputs(7675));
    outputs(5773) <= (layer0_outputs(5500)) xor (layer0_outputs(1440));
    outputs(5774) <= (layer0_outputs(1116)) xor (layer0_outputs(6069));
    outputs(5775) <= layer0_outputs(6737);
    outputs(5776) <= not(layer0_outputs(6305));
    outputs(5777) <= (layer0_outputs(1776)) xor (layer0_outputs(6800));
    outputs(5778) <= not((layer0_outputs(5381)) xor (layer0_outputs(653)));
    outputs(5779) <= layer0_outputs(5448);
    outputs(5780) <= not(layer0_outputs(8919));
    outputs(5781) <= (layer0_outputs(1978)) xor (layer0_outputs(8019));
    outputs(5782) <= not((layer0_outputs(6355)) xor (layer0_outputs(8237)));
    outputs(5783) <= not(layer0_outputs(3988));
    outputs(5784) <= not(layer0_outputs(6307));
    outputs(5785) <= (layer0_outputs(9460)) or (layer0_outputs(487));
    outputs(5786) <= layer0_outputs(5601);
    outputs(5787) <= layer0_outputs(7392);
    outputs(5788) <= not((layer0_outputs(6875)) or (layer0_outputs(546)));
    outputs(5789) <= layer0_outputs(5215);
    outputs(5790) <= (layer0_outputs(9012)) xor (layer0_outputs(1015));
    outputs(5791) <= layer0_outputs(2139);
    outputs(5792) <= (layer0_outputs(8586)) xor (layer0_outputs(6113));
    outputs(5793) <= layer0_outputs(4542);
    outputs(5794) <= layer0_outputs(1019);
    outputs(5795) <= not(layer0_outputs(7203));
    outputs(5796) <= (layer0_outputs(9957)) or (layer0_outputs(8094));
    outputs(5797) <= layer0_outputs(5657);
    outputs(5798) <= not(layer0_outputs(10196)) or (layer0_outputs(9873));
    outputs(5799) <= layer0_outputs(2869);
    outputs(5800) <= not((layer0_outputs(1534)) and (layer0_outputs(3919)));
    outputs(5801) <= not(layer0_outputs(3428));
    outputs(5802) <= not((layer0_outputs(1702)) or (layer0_outputs(2658)));
    outputs(5803) <= layer0_outputs(4839);
    outputs(5804) <= (layer0_outputs(7471)) xor (layer0_outputs(6939));
    outputs(5805) <= not((layer0_outputs(1414)) xor (layer0_outputs(9751)));
    outputs(5806) <= not(layer0_outputs(6786)) or (layer0_outputs(2725));
    outputs(5807) <= '1';
    outputs(5808) <= not(layer0_outputs(8486));
    outputs(5809) <= (layer0_outputs(1571)) xor (layer0_outputs(3220));
    outputs(5810) <= not(layer0_outputs(7968));
    outputs(5811) <= not((layer0_outputs(1362)) and (layer0_outputs(6862)));
    outputs(5812) <= not(layer0_outputs(2566));
    outputs(5813) <= layer0_outputs(6193);
    outputs(5814) <= layer0_outputs(9768);
    outputs(5815) <= not((layer0_outputs(1934)) xor (layer0_outputs(4157)));
    outputs(5816) <= not(layer0_outputs(8510));
    outputs(5817) <= not((layer0_outputs(5490)) xor (layer0_outputs(7028)));
    outputs(5818) <= layer0_outputs(7067);
    outputs(5819) <= (layer0_outputs(2034)) and not (layer0_outputs(2835));
    outputs(5820) <= not(layer0_outputs(8384));
    outputs(5821) <= layer0_outputs(9910);
    outputs(5822) <= (layer0_outputs(8093)) and not (layer0_outputs(6338));
    outputs(5823) <= not(layer0_outputs(5962)) or (layer0_outputs(7526));
    outputs(5824) <= (layer0_outputs(6415)) xor (layer0_outputs(9043));
    outputs(5825) <= layer0_outputs(527);
    outputs(5826) <= (layer0_outputs(2238)) xor (layer0_outputs(8072));
    outputs(5827) <= (layer0_outputs(8107)) xor (layer0_outputs(919));
    outputs(5828) <= not((layer0_outputs(4225)) or (layer0_outputs(4126)));
    outputs(5829) <= not((layer0_outputs(2389)) and (layer0_outputs(5417)));
    outputs(5830) <= not(layer0_outputs(2531));
    outputs(5831) <= not(layer0_outputs(3253));
    outputs(5832) <= not(layer0_outputs(1654)) or (layer0_outputs(7587));
    outputs(5833) <= not((layer0_outputs(7215)) xor (layer0_outputs(10193)));
    outputs(5834) <= not(layer0_outputs(3742));
    outputs(5835) <= not(layer0_outputs(6204));
    outputs(5836) <= layer0_outputs(2116);
    outputs(5837) <= not((layer0_outputs(6473)) xor (layer0_outputs(3706)));
    outputs(5838) <= not((layer0_outputs(9794)) xor (layer0_outputs(4974)));
    outputs(5839) <= not((layer0_outputs(6120)) xor (layer0_outputs(2105)));
    outputs(5840) <= not((layer0_outputs(8629)) and (layer0_outputs(8211)));
    outputs(5841) <= not(layer0_outputs(6441));
    outputs(5842) <= (layer0_outputs(3218)) xor (layer0_outputs(5178));
    outputs(5843) <= layer0_outputs(508);
    outputs(5844) <= (layer0_outputs(5875)) xor (layer0_outputs(1008));
    outputs(5845) <= layer0_outputs(9333);
    outputs(5846) <= layer0_outputs(6757);
    outputs(5847) <= layer0_outputs(10200);
    outputs(5848) <= not(layer0_outputs(7633));
    outputs(5849) <= not((layer0_outputs(2962)) xor (layer0_outputs(3475)));
    outputs(5850) <= (layer0_outputs(4216)) xor (layer0_outputs(9138));
    outputs(5851) <= layer0_outputs(3115);
    outputs(5852) <= layer0_outputs(2595);
    outputs(5853) <= not(layer0_outputs(4082));
    outputs(5854) <= not((layer0_outputs(7861)) xor (layer0_outputs(5256)));
    outputs(5855) <= not((layer0_outputs(7950)) and (layer0_outputs(7014)));
    outputs(5856) <= layer0_outputs(10082);
    outputs(5857) <= not(layer0_outputs(9759));
    outputs(5858) <= not(layer0_outputs(3769)) or (layer0_outputs(8295));
    outputs(5859) <= layer0_outputs(7076);
    outputs(5860) <= layer0_outputs(7335);
    outputs(5861) <= layer0_outputs(7478);
    outputs(5862) <= (layer0_outputs(3599)) and (layer0_outputs(6434));
    outputs(5863) <= layer0_outputs(6433);
    outputs(5864) <= (layer0_outputs(7079)) xor (layer0_outputs(8918));
    outputs(5865) <= (layer0_outputs(7103)) xor (layer0_outputs(4080));
    outputs(5866) <= (layer0_outputs(465)) or (layer0_outputs(4582));
    outputs(5867) <= (layer0_outputs(9643)) and (layer0_outputs(482));
    outputs(5868) <= not((layer0_outputs(6404)) xor (layer0_outputs(7197)));
    outputs(5869) <= (layer0_outputs(4044)) xor (layer0_outputs(1570));
    outputs(5870) <= not(layer0_outputs(2453));
    outputs(5871) <= layer0_outputs(2673);
    outputs(5872) <= layer0_outputs(838);
    outputs(5873) <= layer0_outputs(8220);
    outputs(5874) <= (layer0_outputs(1275)) and (layer0_outputs(3009));
    outputs(5875) <= not(layer0_outputs(1331));
    outputs(5876) <= not(layer0_outputs(9933));
    outputs(5877) <= not((layer0_outputs(3664)) xor (layer0_outputs(8575)));
    outputs(5878) <= not(layer0_outputs(9112));
    outputs(5879) <= not((layer0_outputs(3013)) xor (layer0_outputs(9242)));
    outputs(5880) <= not((layer0_outputs(4921)) xor (layer0_outputs(9376)));
    outputs(5881) <= not((layer0_outputs(4788)) and (layer0_outputs(3316)));
    outputs(5882) <= layer0_outputs(2509);
    outputs(5883) <= not((layer0_outputs(2705)) xor (layer0_outputs(1765)));
    outputs(5884) <= not((layer0_outputs(6241)) xor (layer0_outputs(5650)));
    outputs(5885) <= layer0_outputs(6144);
    outputs(5886) <= not(layer0_outputs(10140));
    outputs(5887) <= not(layer0_outputs(4896));
    outputs(5888) <= not(layer0_outputs(6582));
    outputs(5889) <= not(layer0_outputs(9316));
    outputs(5890) <= layer0_outputs(866);
    outputs(5891) <= (layer0_outputs(6299)) xor (layer0_outputs(5974));
    outputs(5892) <= layer0_outputs(5053);
    outputs(5893) <= not((layer0_outputs(891)) xor (layer0_outputs(3448)));
    outputs(5894) <= layer0_outputs(1101);
    outputs(5895) <= layer0_outputs(8348);
    outputs(5896) <= not((layer0_outputs(6847)) xor (layer0_outputs(8168)));
    outputs(5897) <= not(layer0_outputs(8906));
    outputs(5898) <= (layer0_outputs(3383)) xor (layer0_outputs(7110));
    outputs(5899) <= not((layer0_outputs(8144)) xor (layer0_outputs(7232)));
    outputs(5900) <= not(layer0_outputs(5151)) or (layer0_outputs(734));
    outputs(5901) <= not(layer0_outputs(4281));
    outputs(5902) <= not((layer0_outputs(10178)) and (layer0_outputs(6425)));
    outputs(5903) <= not(layer0_outputs(4030));
    outputs(5904) <= not(layer0_outputs(4409));
    outputs(5905) <= (layer0_outputs(397)) xor (layer0_outputs(4818));
    outputs(5906) <= not(layer0_outputs(6715));
    outputs(5907) <= not(layer0_outputs(2901));
    outputs(5908) <= (layer0_outputs(2518)) xor (layer0_outputs(686));
    outputs(5909) <= (layer0_outputs(4925)) xor (layer0_outputs(352));
    outputs(5910) <= not(layer0_outputs(3845));
    outputs(5911) <= layer0_outputs(6131);
    outputs(5912) <= not((layer0_outputs(4345)) xor (layer0_outputs(3739)));
    outputs(5913) <= not((layer0_outputs(4547)) xor (layer0_outputs(2648)));
    outputs(5914) <= not((layer0_outputs(353)) xor (layer0_outputs(5999)));
    outputs(5915) <= layer0_outputs(506);
    outputs(5916) <= (layer0_outputs(5953)) xor (layer0_outputs(6811));
    outputs(5917) <= (layer0_outputs(10228)) and (layer0_outputs(3051));
    outputs(5918) <= (layer0_outputs(3625)) or (layer0_outputs(6077));
    outputs(5919) <= layer0_outputs(9166);
    outputs(5920) <= layer0_outputs(1498);
    outputs(5921) <= not(layer0_outputs(9944)) or (layer0_outputs(1017));
    outputs(5922) <= not(layer0_outputs(3690));
    outputs(5923) <= not(layer0_outputs(2667));
    outputs(5924) <= (layer0_outputs(9667)) and not (layer0_outputs(869));
    outputs(5925) <= not(layer0_outputs(8695)) or (layer0_outputs(9348));
    outputs(5926) <= not(layer0_outputs(3026));
    outputs(5927) <= layer0_outputs(6077);
    outputs(5928) <= not(layer0_outputs(7878));
    outputs(5929) <= not((layer0_outputs(7155)) and (layer0_outputs(4214)));
    outputs(5930) <= not((layer0_outputs(3415)) xor (layer0_outputs(3219)));
    outputs(5931) <= not(layer0_outputs(3760));
    outputs(5932) <= not(layer0_outputs(6700));
    outputs(5933) <= not(layer0_outputs(1057));
    outputs(5934) <= (layer0_outputs(7426)) and not (layer0_outputs(7489));
    outputs(5935) <= layer0_outputs(1564);
    outputs(5936) <= not(layer0_outputs(1135));
    outputs(5937) <= layer0_outputs(7505);
    outputs(5938) <= not((layer0_outputs(9266)) and (layer0_outputs(9674)));
    outputs(5939) <= layer0_outputs(9216);
    outputs(5940) <= layer0_outputs(2868);
    outputs(5941) <= layer0_outputs(9607);
    outputs(5942) <= layer0_outputs(7790);
    outputs(5943) <= (layer0_outputs(1105)) or (layer0_outputs(8262));
    outputs(5944) <= (layer0_outputs(7769)) xor (layer0_outputs(7997));
    outputs(5945) <= (layer0_outputs(4911)) and (layer0_outputs(937));
    outputs(5946) <= (layer0_outputs(4146)) or (layer0_outputs(7773));
    outputs(5947) <= layer0_outputs(7063);
    outputs(5948) <= not(layer0_outputs(1016));
    outputs(5949) <= not(layer0_outputs(1051));
    outputs(5950) <= layer0_outputs(1001);
    outputs(5951) <= not(layer0_outputs(262));
    outputs(5952) <= layer0_outputs(2971);
    outputs(5953) <= (layer0_outputs(3134)) xor (layer0_outputs(7210));
    outputs(5954) <= not((layer0_outputs(157)) xor (layer0_outputs(3406)));
    outputs(5955) <= not(layer0_outputs(7503));
    outputs(5956) <= (layer0_outputs(3628)) xor (layer0_outputs(1036));
    outputs(5957) <= not((layer0_outputs(280)) or (layer0_outputs(3300)));
    outputs(5958) <= not((layer0_outputs(8737)) xor (layer0_outputs(5355)));
    outputs(5959) <= (layer0_outputs(1892)) and not (layer0_outputs(9327));
    outputs(5960) <= layer0_outputs(1885);
    outputs(5961) <= not(layer0_outputs(5413));
    outputs(5962) <= not(layer0_outputs(137));
    outputs(5963) <= layer0_outputs(1494);
    outputs(5964) <= not(layer0_outputs(8302)) or (layer0_outputs(7660));
    outputs(5965) <= not(layer0_outputs(7050));
    outputs(5966) <= not(layer0_outputs(4538));
    outputs(5967) <= not((layer0_outputs(9018)) xor (layer0_outputs(8727)));
    outputs(5968) <= not((layer0_outputs(6344)) or (layer0_outputs(7241)));
    outputs(5969) <= layer0_outputs(2793);
    outputs(5970) <= (layer0_outputs(8136)) xor (layer0_outputs(4235));
    outputs(5971) <= layer0_outputs(2997);
    outputs(5972) <= layer0_outputs(2820);
    outputs(5973) <= layer0_outputs(7721);
    outputs(5974) <= layer0_outputs(5420);
    outputs(5975) <= (layer0_outputs(7686)) xor (layer0_outputs(7184));
    outputs(5976) <= not(layer0_outputs(261));
    outputs(5977) <= not(layer0_outputs(1441)) or (layer0_outputs(1423));
    outputs(5978) <= (layer0_outputs(454)) xor (layer0_outputs(145));
    outputs(5979) <= not(layer0_outputs(1350));
    outputs(5980) <= not(layer0_outputs(5551));
    outputs(5981) <= (layer0_outputs(6827)) xor (layer0_outputs(1666));
    outputs(5982) <= (layer0_outputs(5876)) xor (layer0_outputs(464));
    outputs(5983) <= not((layer0_outputs(3468)) and (layer0_outputs(4778)));
    outputs(5984) <= (layer0_outputs(4017)) xor (layer0_outputs(8977));
    outputs(5985) <= (layer0_outputs(16)) xor (layer0_outputs(1356));
    outputs(5986) <= (layer0_outputs(8650)) xor (layer0_outputs(3522));
    outputs(5987) <= not(layer0_outputs(1293));
    outputs(5988) <= layer0_outputs(4418);
    outputs(5989) <= not(layer0_outputs(4545));
    outputs(5990) <= not(layer0_outputs(5489)) or (layer0_outputs(9825));
    outputs(5991) <= layer0_outputs(2233);
    outputs(5992) <= (layer0_outputs(8244)) or (layer0_outputs(9421));
    outputs(5993) <= not(layer0_outputs(8587)) or (layer0_outputs(5923));
    outputs(5994) <= not(layer0_outputs(7271)) or (layer0_outputs(9785));
    outputs(5995) <= not((layer0_outputs(8422)) xor (layer0_outputs(6105)));
    outputs(5996) <= (layer0_outputs(4161)) or (layer0_outputs(5272));
    outputs(5997) <= not(layer0_outputs(9593)) or (layer0_outputs(663));
    outputs(5998) <= layer0_outputs(7462);
    outputs(5999) <= (layer0_outputs(6340)) xor (layer0_outputs(8054));
    outputs(6000) <= layer0_outputs(4640);
    outputs(6001) <= not(layer0_outputs(6196));
    outputs(6002) <= (layer0_outputs(6246)) and (layer0_outputs(7398));
    outputs(6003) <= not(layer0_outputs(8521));
    outputs(6004) <= not(layer0_outputs(5335));
    outputs(6005) <= layer0_outputs(7074);
    outputs(6006) <= (layer0_outputs(8133)) and (layer0_outputs(3022));
    outputs(6007) <= not(layer0_outputs(453)) or (layer0_outputs(3133));
    outputs(6008) <= layer0_outputs(6278);
    outputs(6009) <= not((layer0_outputs(5048)) xor (layer0_outputs(8102)));
    outputs(6010) <= not(layer0_outputs(3863));
    outputs(6011) <= (layer0_outputs(1646)) or (layer0_outputs(3916));
    outputs(6012) <= not(layer0_outputs(8594));
    outputs(6013) <= not(layer0_outputs(77)) or (layer0_outputs(6578));
    outputs(6014) <= not((layer0_outputs(5298)) xor (layer0_outputs(2691)));
    outputs(6015) <= not((layer0_outputs(5368)) xor (layer0_outputs(9909)));
    outputs(6016) <= layer0_outputs(679);
    outputs(6017) <= not(layer0_outputs(5781));
    outputs(6018) <= layer0_outputs(1494);
    outputs(6019) <= not(layer0_outputs(5466)) or (layer0_outputs(9403));
    outputs(6020) <= (layer0_outputs(494)) or (layer0_outputs(5025));
    outputs(6021) <= (layer0_outputs(7278)) and not (layer0_outputs(2866));
    outputs(6022) <= (layer0_outputs(8158)) or (layer0_outputs(1313));
    outputs(6023) <= (layer0_outputs(2169)) xor (layer0_outputs(4473));
    outputs(6024) <= (layer0_outputs(2463)) xor (layer0_outputs(1398));
    outputs(6025) <= not(layer0_outputs(1693));
    outputs(6026) <= layer0_outputs(7636);
    outputs(6027) <= (layer0_outputs(10126)) and (layer0_outputs(588));
    outputs(6028) <= not((layer0_outputs(6810)) xor (layer0_outputs(3188)));
    outputs(6029) <= layer0_outputs(3083);
    outputs(6030) <= (layer0_outputs(4852)) xor (layer0_outputs(10171));
    outputs(6031) <= layer0_outputs(6054);
    outputs(6032) <= not(layer0_outputs(4293)) or (layer0_outputs(2653));
    outputs(6033) <= (layer0_outputs(2885)) and not (layer0_outputs(5697));
    outputs(6034) <= not((layer0_outputs(9034)) xor (layer0_outputs(4265)));
    outputs(6035) <= (layer0_outputs(1027)) xor (layer0_outputs(1979));
    outputs(6036) <= (layer0_outputs(1034)) or (layer0_outputs(2980));
    outputs(6037) <= (layer0_outputs(5035)) xor (layer0_outputs(8131));
    outputs(6038) <= not(layer0_outputs(9770));
    outputs(6039) <= not(layer0_outputs(5335));
    outputs(6040) <= not((layer0_outputs(693)) or (layer0_outputs(7718)));
    outputs(6041) <= layer0_outputs(1261);
    outputs(6042) <= (layer0_outputs(7326)) and not (layer0_outputs(1733));
    outputs(6043) <= not((layer0_outputs(5247)) xor (layer0_outputs(9796)));
    outputs(6044) <= (layer0_outputs(8585)) xor (layer0_outputs(2356));
    outputs(6045) <= layer0_outputs(5327);
    outputs(6046) <= (layer0_outputs(9708)) xor (layer0_outputs(9070));
    outputs(6047) <= layer0_outputs(9687);
    outputs(6048) <= not((layer0_outputs(3954)) xor (layer0_outputs(4765)));
    outputs(6049) <= (layer0_outputs(5507)) or (layer0_outputs(7774));
    outputs(6050) <= layer0_outputs(8259);
    outputs(6051) <= not((layer0_outputs(3723)) xor (layer0_outputs(3636)));
    outputs(6052) <= (layer0_outputs(10064)) xor (layer0_outputs(6422));
    outputs(6053) <= not(layer0_outputs(6375));
    outputs(6054) <= not(layer0_outputs(7404)) or (layer0_outputs(5317));
    outputs(6055) <= '1';
    outputs(6056) <= layer0_outputs(2726);
    outputs(6057) <= not(layer0_outputs(1035));
    outputs(6058) <= (layer0_outputs(9072)) xor (layer0_outputs(7128));
    outputs(6059) <= (layer0_outputs(5559)) and (layer0_outputs(9797));
    outputs(6060) <= not(layer0_outputs(4247));
    outputs(6061) <= not(layer0_outputs(2928)) or (layer0_outputs(7042));
    outputs(6062) <= not((layer0_outputs(2188)) xor (layer0_outputs(6215)));
    outputs(6063) <= not((layer0_outputs(9388)) or (layer0_outputs(2565)));
    outputs(6064) <= (layer0_outputs(4899)) and not (layer0_outputs(7653));
    outputs(6065) <= layer0_outputs(3301);
    outputs(6066) <= layer0_outputs(3123);
    outputs(6067) <= not((layer0_outputs(4227)) xor (layer0_outputs(9986)));
    outputs(6068) <= layer0_outputs(2662);
    outputs(6069) <= not(layer0_outputs(1167)) or (layer0_outputs(6549));
    outputs(6070) <= (layer0_outputs(2388)) and (layer0_outputs(9562));
    outputs(6071) <= (layer0_outputs(1272)) or (layer0_outputs(4322));
    outputs(6072) <= not((layer0_outputs(4105)) and (layer0_outputs(5555)));
    outputs(6073) <= layer0_outputs(7467);
    outputs(6074) <= not((layer0_outputs(4521)) or (layer0_outputs(6044)));
    outputs(6075) <= not(layer0_outputs(4566));
    outputs(6076) <= (layer0_outputs(7159)) xor (layer0_outputs(6718));
    outputs(6077) <= layer0_outputs(7631);
    outputs(6078) <= not((layer0_outputs(5490)) xor (layer0_outputs(248)));
    outputs(6079) <= not((layer0_outputs(9716)) and (layer0_outputs(8046)));
    outputs(6080) <= not(layer0_outputs(4403));
    outputs(6081) <= not((layer0_outputs(9416)) xor (layer0_outputs(6211)));
    outputs(6082) <= not(layer0_outputs(7932));
    outputs(6083) <= layer0_outputs(8377);
    outputs(6084) <= layer0_outputs(8296);
    outputs(6085) <= (layer0_outputs(8023)) xor (layer0_outputs(3158));
    outputs(6086) <= not(layer0_outputs(10208));
    outputs(6087) <= (layer0_outputs(344)) xor (layer0_outputs(3161));
    outputs(6088) <= (layer0_outputs(5115)) xor (layer0_outputs(8482));
    outputs(6089) <= layer0_outputs(6157);
    outputs(6090) <= not(layer0_outputs(9641));
    outputs(6091) <= not(layer0_outputs(7906));
    outputs(6092) <= layer0_outputs(2347);
    outputs(6093) <= not(layer0_outputs(9353));
    outputs(6094) <= not(layer0_outputs(3659));
    outputs(6095) <= not((layer0_outputs(6041)) xor (layer0_outputs(8809)));
    outputs(6096) <= not((layer0_outputs(375)) xor (layer0_outputs(494)));
    outputs(6097) <= not(layer0_outputs(4746));
    outputs(6098) <= layer0_outputs(7608);
    outputs(6099) <= (layer0_outputs(7413)) xor (layer0_outputs(8711));
    outputs(6100) <= (layer0_outputs(6825)) xor (layer0_outputs(1060));
    outputs(6101) <= layer0_outputs(1277);
    outputs(6102) <= not(layer0_outputs(709));
    outputs(6103) <= layer0_outputs(5329);
    outputs(6104) <= not((layer0_outputs(7120)) xor (layer0_outputs(3516)));
    outputs(6105) <= not((layer0_outputs(3016)) xor (layer0_outputs(2840)));
    outputs(6106) <= layer0_outputs(6999);
    outputs(6107) <= not(layer0_outputs(5998));
    outputs(6108) <= (layer0_outputs(898)) and not (layer0_outputs(9498));
    outputs(6109) <= layer0_outputs(1014);
    outputs(6110) <= layer0_outputs(8671);
    outputs(6111) <= not(layer0_outputs(3773)) or (layer0_outputs(7770));
    outputs(6112) <= not((layer0_outputs(2785)) xor (layer0_outputs(5745)));
    outputs(6113) <= not((layer0_outputs(6338)) xor (layer0_outputs(1382)));
    outputs(6114) <= not(layer0_outputs(5775)) or (layer0_outputs(8669));
    outputs(6115) <= not(layer0_outputs(2803)) or (layer0_outputs(8879));
    outputs(6116) <= not(layer0_outputs(10109));
    outputs(6117) <= not(layer0_outputs(5592));
    outputs(6118) <= (layer0_outputs(711)) xor (layer0_outputs(6188));
    outputs(6119) <= not(layer0_outputs(5383));
    outputs(6120) <= layer0_outputs(3461);
    outputs(6121) <= layer0_outputs(7488);
    outputs(6122) <= (layer0_outputs(7621)) and (layer0_outputs(5450));
    outputs(6123) <= (layer0_outputs(532)) and (layer0_outputs(8130));
    outputs(6124) <= not(layer0_outputs(8361));
    outputs(6125) <= layer0_outputs(519);
    outputs(6126) <= (layer0_outputs(2396)) xor (layer0_outputs(8219));
    outputs(6127) <= not(layer0_outputs(5894)) or (layer0_outputs(5649));
    outputs(6128) <= not((layer0_outputs(2044)) or (layer0_outputs(9289)));
    outputs(6129) <= layer0_outputs(9915);
    outputs(6130) <= not((layer0_outputs(371)) or (layer0_outputs(9619)));
    outputs(6131) <= not(layer0_outputs(502));
    outputs(6132) <= not(layer0_outputs(5600));
    outputs(6133) <= (layer0_outputs(8820)) and not (layer0_outputs(412));
    outputs(6134) <= (layer0_outputs(1842)) xor (layer0_outputs(536));
    outputs(6135) <= not(layer0_outputs(8026));
    outputs(6136) <= layer0_outputs(6429);
    outputs(6137) <= not(layer0_outputs(128));
    outputs(6138) <= (layer0_outputs(7761)) xor (layer0_outputs(3621));
    outputs(6139) <= layer0_outputs(1717);
    outputs(6140) <= not(layer0_outputs(9735));
    outputs(6141) <= not((layer0_outputs(322)) xor (layer0_outputs(368)));
    outputs(6142) <= not((layer0_outputs(6548)) xor (layer0_outputs(4639)));
    outputs(6143) <= not(layer0_outputs(4666));
    outputs(6144) <= not(layer0_outputs(3752));
    outputs(6145) <= not(layer0_outputs(3934));
    outputs(6146) <= layer0_outputs(2745);
    outputs(6147) <= not((layer0_outputs(72)) and (layer0_outputs(4958)));
    outputs(6148) <= layer0_outputs(504);
    outputs(6149) <= not((layer0_outputs(1063)) xor (layer0_outputs(3090)));
    outputs(6150) <= not(layer0_outputs(9349));
    outputs(6151) <= not(layer0_outputs(6956));
    outputs(6152) <= not((layer0_outputs(10090)) xor (layer0_outputs(7647)));
    outputs(6153) <= not(layer0_outputs(2683));
    outputs(6154) <= layer0_outputs(3543);
    outputs(6155) <= not(layer0_outputs(269));
    outputs(6156) <= layer0_outputs(2216);
    outputs(6157) <= not((layer0_outputs(7231)) xor (layer0_outputs(9733)));
    outputs(6158) <= not(layer0_outputs(4353));
    outputs(6159) <= layer0_outputs(7694);
    outputs(6160) <= not(layer0_outputs(5077));
    outputs(6161) <= not(layer0_outputs(161));
    outputs(6162) <= not((layer0_outputs(7417)) and (layer0_outputs(8170)));
    outputs(6163) <= not(layer0_outputs(3313));
    outputs(6164) <= (layer0_outputs(3340)) and not (layer0_outputs(6473));
    outputs(6165) <= not(layer0_outputs(4705)) or (layer0_outputs(3813));
    outputs(6166) <= layer0_outputs(5854);
    outputs(6167) <= not(layer0_outputs(8287));
    outputs(6168) <= not(layer0_outputs(7090));
    outputs(6169) <= layer0_outputs(7425);
    outputs(6170) <= (layer0_outputs(8596)) xor (layer0_outputs(6843));
    outputs(6171) <= not((layer0_outputs(8800)) or (layer0_outputs(2056)));
    outputs(6172) <= not((layer0_outputs(85)) xor (layer0_outputs(7387)));
    outputs(6173) <= layer0_outputs(4127);
    outputs(6174) <= not(layer0_outputs(6349));
    outputs(6175) <= layer0_outputs(555);
    outputs(6176) <= not((layer0_outputs(5325)) xor (layer0_outputs(2027)));
    outputs(6177) <= layer0_outputs(1386);
    outputs(6178) <= not((layer0_outputs(9545)) or (layer0_outputs(1214)));
    outputs(6179) <= not((layer0_outputs(5336)) xor (layer0_outputs(7311)));
    outputs(6180) <= layer0_outputs(7265);
    outputs(6181) <= not(layer0_outputs(5431));
    outputs(6182) <= not(layer0_outputs(3146));
    outputs(6183) <= (layer0_outputs(3344)) and not (layer0_outputs(15));
    outputs(6184) <= layer0_outputs(815);
    outputs(6185) <= not(layer0_outputs(8269));
    outputs(6186) <= layer0_outputs(3975);
    outputs(6187) <= layer0_outputs(7798);
    outputs(6188) <= not(layer0_outputs(9278));
    outputs(6189) <= not((layer0_outputs(866)) and (layer0_outputs(9521)));
    outputs(6190) <= (layer0_outputs(4750)) and not (layer0_outputs(9666));
    outputs(6191) <= layer0_outputs(4934);
    outputs(6192) <= not((layer0_outputs(8216)) xor (layer0_outputs(2204)));
    outputs(6193) <= not((layer0_outputs(2217)) or (layer0_outputs(7503)));
    outputs(6194) <= (layer0_outputs(4897)) and not (layer0_outputs(6662));
    outputs(6195) <= (layer0_outputs(9345)) xor (layer0_outputs(7754));
    outputs(6196) <= not(layer0_outputs(3815));
    outputs(6197) <= layer0_outputs(9655);
    outputs(6198) <= not(layer0_outputs(8203));
    outputs(6199) <= layer0_outputs(6656);
    outputs(6200) <= not(layer0_outputs(9666));
    outputs(6201) <= not((layer0_outputs(7784)) xor (layer0_outputs(6235)));
    outputs(6202) <= (layer0_outputs(3725)) and not (layer0_outputs(4064));
    outputs(6203) <= not(layer0_outputs(2090));
    outputs(6204) <= layer0_outputs(6585);
    outputs(6205) <= (layer0_outputs(5730)) and not (layer0_outputs(313));
    outputs(6206) <= not(layer0_outputs(953));
    outputs(6207) <= layer0_outputs(3755);
    outputs(6208) <= (layer0_outputs(6173)) and not (layer0_outputs(1561));
    outputs(6209) <= layer0_outputs(167);
    outputs(6210) <= (layer0_outputs(4362)) and not (layer0_outputs(5177));
    outputs(6211) <= not(layer0_outputs(10185));
    outputs(6212) <= not(layer0_outputs(5580));
    outputs(6213) <= not(layer0_outputs(7676));
    outputs(6214) <= layer0_outputs(3228);
    outputs(6215) <= layer0_outputs(4481);
    outputs(6216) <= not(layer0_outputs(2951));
    outputs(6217) <= layer0_outputs(6219);
    outputs(6218) <= not(layer0_outputs(8967));
    outputs(6219) <= not(layer0_outputs(3719));
    outputs(6220) <= not(layer0_outputs(9489));
    outputs(6221) <= (layer0_outputs(8814)) xor (layer0_outputs(6785));
    outputs(6222) <= not(layer0_outputs(2481)) or (layer0_outputs(8402));
    outputs(6223) <= (layer0_outputs(5275)) and not (layer0_outputs(5771));
    outputs(6224) <= layer0_outputs(8964);
    outputs(6225) <= not(layer0_outputs(9763));
    outputs(6226) <= (layer0_outputs(5)) xor (layer0_outputs(2214));
    outputs(6227) <= not(layer0_outputs(9463));
    outputs(6228) <= (layer0_outputs(1821)) and not (layer0_outputs(567));
    outputs(6229) <= not((layer0_outputs(10138)) or (layer0_outputs(303)));
    outputs(6230) <= not(layer0_outputs(6365));
    outputs(6231) <= layer0_outputs(5562);
    outputs(6232) <= not(layer0_outputs(4193)) or (layer0_outputs(3068));
    outputs(6233) <= not(layer0_outputs(5762));
    outputs(6234) <= (layer0_outputs(7994)) and (layer0_outputs(7354));
    outputs(6235) <= layer0_outputs(4517);
    outputs(6236) <= (layer0_outputs(2572)) xor (layer0_outputs(98));
    outputs(6237) <= layer0_outputs(2948);
    outputs(6238) <= not((layer0_outputs(5873)) or (layer0_outputs(3484)));
    outputs(6239) <= (layer0_outputs(6871)) and (layer0_outputs(5754));
    outputs(6240) <= layer0_outputs(4974);
    outputs(6241) <= layer0_outputs(1642);
    outputs(6242) <= layer0_outputs(7523);
    outputs(6243) <= not((layer0_outputs(2721)) or (layer0_outputs(2794)));
    outputs(6244) <= layer0_outputs(7287);
    outputs(6245) <= (layer0_outputs(2521)) and not (layer0_outputs(9332));
    outputs(6246) <= not(layer0_outputs(6456));
    outputs(6247) <= not((layer0_outputs(2217)) and (layer0_outputs(2859)));
    outputs(6248) <= (layer0_outputs(2343)) and not (layer0_outputs(6781));
    outputs(6249) <= not(layer0_outputs(7038));
    outputs(6250) <= not((layer0_outputs(9572)) or (layer0_outputs(4622)));
    outputs(6251) <= not((layer0_outputs(5988)) xor (layer0_outputs(713)));
    outputs(6252) <= not(layer0_outputs(3893));
    outputs(6253) <= layer0_outputs(6739);
    outputs(6254) <= layer0_outputs(818);
    outputs(6255) <= layer0_outputs(428);
    outputs(6256) <= layer0_outputs(6679);
    outputs(6257) <= not(layer0_outputs(6897));
    outputs(6258) <= not(layer0_outputs(3012));
    outputs(6259) <= (layer0_outputs(253)) xor (layer0_outputs(5978));
    outputs(6260) <= not(layer0_outputs(3360));
    outputs(6261) <= layer0_outputs(6732);
    outputs(6262) <= not(layer0_outputs(8404));
    outputs(6263) <= not(layer0_outputs(5726));
    outputs(6264) <= (layer0_outputs(7068)) xor (layer0_outputs(1225));
    outputs(6265) <= not(layer0_outputs(1230));
    outputs(6266) <= (layer0_outputs(3455)) xor (layer0_outputs(1449));
    outputs(6267) <= (layer0_outputs(8209)) and not (layer0_outputs(3510));
    outputs(6268) <= layer0_outputs(7742);
    outputs(6269) <= (layer0_outputs(10144)) and not (layer0_outputs(2464));
    outputs(6270) <= layer0_outputs(5861);
    outputs(6271) <= not((layer0_outputs(2843)) xor (layer0_outputs(9476)));
    outputs(6272) <= layer0_outputs(7034);
    outputs(6273) <= (layer0_outputs(4905)) xor (layer0_outputs(2972));
    outputs(6274) <= layer0_outputs(7233);
    outputs(6275) <= not(layer0_outputs(7922));
    outputs(6276) <= (layer0_outputs(3347)) and not (layer0_outputs(321));
    outputs(6277) <= not(layer0_outputs(5638));
    outputs(6278) <= layer0_outputs(907);
    outputs(6279) <= not((layer0_outputs(4628)) or (layer0_outputs(116)));
    outputs(6280) <= not(layer0_outputs(6153));
    outputs(6281) <= layer0_outputs(9591);
    outputs(6282) <= '1';
    outputs(6283) <= (layer0_outputs(3266)) and not (layer0_outputs(9720));
    outputs(6284) <= layer0_outputs(7734);
    outputs(6285) <= not(layer0_outputs(3944)) or (layer0_outputs(5298));
    outputs(6286) <= not((layer0_outputs(2213)) xor (layer0_outputs(9871)));
    outputs(6287) <= (layer0_outputs(6331)) xor (layer0_outputs(9920));
    outputs(6288) <= not(layer0_outputs(1626));
    outputs(6289) <= (layer0_outputs(4567)) or (layer0_outputs(4691));
    outputs(6290) <= layer0_outputs(5386);
    outputs(6291) <= (layer0_outputs(2538)) and not (layer0_outputs(6742));
    outputs(6292) <= layer0_outputs(6974);
    outputs(6293) <= not(layer0_outputs(4906));
    outputs(6294) <= not(layer0_outputs(1439)) or (layer0_outputs(8960));
    outputs(6295) <= layer0_outputs(3607);
    outputs(6296) <= layer0_outputs(4526);
    outputs(6297) <= (layer0_outputs(8270)) and not (layer0_outputs(8420));
    outputs(6298) <= not((layer0_outputs(10127)) xor (layer0_outputs(2382)));
    outputs(6299) <= not(layer0_outputs(9933));
    outputs(6300) <= layer0_outputs(5786);
    outputs(6301) <= not(layer0_outputs(6686));
    outputs(6302) <= (layer0_outputs(10101)) and not (layer0_outputs(3807));
    outputs(6303) <= (layer0_outputs(3979)) and not (layer0_outputs(2024));
    outputs(6304) <= not(layer0_outputs(2790));
    outputs(6305) <= (layer0_outputs(9424)) xor (layer0_outputs(6889));
    outputs(6306) <= not(layer0_outputs(10102));
    outputs(6307) <= (layer0_outputs(5379)) and (layer0_outputs(4335));
    outputs(6308) <= not((layer0_outputs(5290)) xor (layer0_outputs(9862)));
    outputs(6309) <= layer0_outputs(7005);
    outputs(6310) <= (layer0_outputs(4532)) and not (layer0_outputs(10091));
    outputs(6311) <= layer0_outputs(8008);
    outputs(6312) <= not((layer0_outputs(6564)) xor (layer0_outputs(5603)));
    outputs(6313) <= not(layer0_outputs(4307));
    outputs(6314) <= not((layer0_outputs(7227)) or (layer0_outputs(2973)));
    outputs(6315) <= layer0_outputs(7259);
    outputs(6316) <= (layer0_outputs(9005)) xor (layer0_outputs(2272));
    outputs(6317) <= layer0_outputs(1291);
    outputs(6318) <= (layer0_outputs(803)) and (layer0_outputs(9385));
    outputs(6319) <= (layer0_outputs(1913)) or (layer0_outputs(2687));
    outputs(6320) <= (layer0_outputs(9300)) or (layer0_outputs(6511));
    outputs(6321) <= layer0_outputs(9132);
    outputs(6322) <= (layer0_outputs(2946)) and not (layer0_outputs(4546));
    outputs(6323) <= (layer0_outputs(3880)) and (layer0_outputs(5806));
    outputs(6324) <= not(layer0_outputs(8238)) or (layer0_outputs(1922));
    outputs(6325) <= not(layer0_outputs(6431));
    outputs(6326) <= (layer0_outputs(4795)) and not (layer0_outputs(3102));
    outputs(6327) <= layer0_outputs(6856);
    outputs(6328) <= not((layer0_outputs(2284)) or (layer0_outputs(7417)));
    outputs(6329) <= (layer0_outputs(9623)) or (layer0_outputs(2802));
    outputs(6330) <= not(layer0_outputs(4968));
    outputs(6331) <= layer0_outputs(9457);
    outputs(6332) <= not(layer0_outputs(3863));
    outputs(6333) <= (layer0_outputs(8332)) and not (layer0_outputs(1147));
    outputs(6334) <= not((layer0_outputs(4798)) or (layer0_outputs(2696)));
    outputs(6335) <= (layer0_outputs(4989)) xor (layer0_outputs(4374));
    outputs(6336) <= not(layer0_outputs(9969));
    outputs(6337) <= layer0_outputs(2764);
    outputs(6338) <= not(layer0_outputs(9411));
    outputs(6339) <= layer0_outputs(10209);
    outputs(6340) <= not(layer0_outputs(3446));
    outputs(6341) <= (layer0_outputs(10237)) or (layer0_outputs(212));
    outputs(6342) <= (layer0_outputs(5137)) and (layer0_outputs(9475));
    outputs(6343) <= not(layer0_outputs(967));
    outputs(6344) <= layer0_outputs(597);
    outputs(6345) <= not(layer0_outputs(8374));
    outputs(6346) <= layer0_outputs(7039);
    outputs(6347) <= layer0_outputs(8553);
    outputs(6348) <= (layer0_outputs(723)) xor (layer0_outputs(3608));
    outputs(6349) <= not(layer0_outputs(1212));
    outputs(6350) <= layer0_outputs(7998);
    outputs(6351) <= not((layer0_outputs(1077)) or (layer0_outputs(8821)));
    outputs(6352) <= layer0_outputs(204);
    outputs(6353) <= (layer0_outputs(8699)) xor (layer0_outputs(2593));
    outputs(6354) <= not(layer0_outputs(1463)) or (layer0_outputs(9918));
    outputs(6355) <= layer0_outputs(4647);
    outputs(6356) <= not(layer0_outputs(3852));
    outputs(6357) <= (layer0_outputs(4812)) xor (layer0_outputs(2032));
    outputs(6358) <= not(layer0_outputs(2317));
    outputs(6359) <= (layer0_outputs(4249)) and not (layer0_outputs(4960));
    outputs(6360) <= layer0_outputs(8947);
    outputs(6361) <= layer0_outputs(5147);
    outputs(6362) <= layer0_outputs(7626);
    outputs(6363) <= layer0_outputs(619);
    outputs(6364) <= not(layer0_outputs(10077));
    outputs(6365) <= not(layer0_outputs(3422));
    outputs(6366) <= not(layer0_outputs(5619)) or (layer0_outputs(555));
    outputs(6367) <= not((layer0_outputs(7903)) and (layer0_outputs(8869)));
    outputs(6368) <= layer0_outputs(2751);
    outputs(6369) <= not(layer0_outputs(4927));
    outputs(6370) <= not((layer0_outputs(118)) xor (layer0_outputs(7341)));
    outputs(6371) <= (layer0_outputs(7547)) and not (layer0_outputs(1379));
    outputs(6372) <= layer0_outputs(2385);
    outputs(6373) <= layer0_outputs(3414);
    outputs(6374) <= not(layer0_outputs(7258));
    outputs(6375) <= (layer0_outputs(6546)) and not (layer0_outputs(6402));
    outputs(6376) <= (layer0_outputs(8309)) xor (layer0_outputs(6042));
    outputs(6377) <= not((layer0_outputs(5555)) and (layer0_outputs(6709)));
    outputs(6378) <= layer0_outputs(2863);
    outputs(6379) <= not(layer0_outputs(9681));
    outputs(6380) <= layer0_outputs(5932);
    outputs(6381) <= (layer0_outputs(2124)) and not (layer0_outputs(1756));
    outputs(6382) <= layer0_outputs(8063);
    outputs(6383) <= not(layer0_outputs(9860)) or (layer0_outputs(4438));
    outputs(6384) <= not(layer0_outputs(492));
    outputs(6385) <= not(layer0_outputs(832));
    outputs(6386) <= not(layer0_outputs(1052));
    outputs(6387) <= not(layer0_outputs(8087));
    outputs(6388) <= not((layer0_outputs(9136)) or (layer0_outputs(5032)));
    outputs(6389) <= (layer0_outputs(2046)) xor (layer0_outputs(6780));
    outputs(6390) <= not(layer0_outputs(9649));
    outputs(6391) <= (layer0_outputs(1068)) and (layer0_outputs(9798));
    outputs(6392) <= not((layer0_outputs(1409)) xor (layer0_outputs(8195)));
    outputs(6393) <= not(layer0_outputs(492));
    outputs(6394) <= layer0_outputs(183);
    outputs(6395) <= not(layer0_outputs(3247)) or (layer0_outputs(622));
    outputs(6396) <= (layer0_outputs(9)) and not (layer0_outputs(5048));
    outputs(6397) <= layer0_outputs(2498);
    outputs(6398) <= layer0_outputs(2373);
    outputs(6399) <= layer0_outputs(652);
    outputs(6400) <= (layer0_outputs(5944)) and not (layer0_outputs(1947));
    outputs(6401) <= not((layer0_outputs(3507)) and (layer0_outputs(2247)));
    outputs(6402) <= not(layer0_outputs(5965));
    outputs(6403) <= layer0_outputs(8161);
    outputs(6404) <= not((layer0_outputs(6293)) or (layer0_outputs(8354)));
    outputs(6405) <= (layer0_outputs(3821)) xor (layer0_outputs(3036));
    outputs(6406) <= not(layer0_outputs(7045));
    outputs(6407) <= layer0_outputs(909);
    outputs(6408) <= not(layer0_outputs(5388)) or (layer0_outputs(2791));
    outputs(6409) <= not((layer0_outputs(3278)) xor (layer0_outputs(4129)));
    outputs(6410) <= not(layer0_outputs(7448));
    outputs(6411) <= not(layer0_outputs(5581));
    outputs(6412) <= (layer0_outputs(8334)) and not (layer0_outputs(10162));
    outputs(6413) <= not(layer0_outputs(2140));
    outputs(6414) <= (layer0_outputs(8044)) and not (layer0_outputs(8095));
    outputs(6415) <= not((layer0_outputs(4643)) xor (layer0_outputs(8114)));
    outputs(6416) <= (layer0_outputs(6284)) and not (layer0_outputs(5478));
    outputs(6417) <= not(layer0_outputs(9398)) or (layer0_outputs(4702));
    outputs(6418) <= layer0_outputs(2183);
    outputs(6419) <= not((layer0_outputs(1318)) xor (layer0_outputs(5828)));
    outputs(6420) <= not(layer0_outputs(6260));
    outputs(6421) <= not(layer0_outputs(7841));
    outputs(6422) <= not(layer0_outputs(4878));
    outputs(6423) <= not(layer0_outputs(2922));
    outputs(6424) <= not(layer0_outputs(4299));
    outputs(6425) <= not((layer0_outputs(3252)) xor (layer0_outputs(1138)));
    outputs(6426) <= (layer0_outputs(4516)) and not (layer0_outputs(6488));
    outputs(6427) <= layer0_outputs(648);
    outputs(6428) <= not((layer0_outputs(2720)) xor (layer0_outputs(3711)));
    outputs(6429) <= not(layer0_outputs(1288));
    outputs(6430) <= layer0_outputs(2186);
    outputs(6431) <= (layer0_outputs(351)) xor (layer0_outputs(5640));
    outputs(6432) <= layer0_outputs(7842);
    outputs(6433) <= not(layer0_outputs(4531)) or (layer0_outputs(813));
    outputs(6434) <= not(layer0_outputs(5283));
    outputs(6435) <= layer0_outputs(6616);
    outputs(6436) <= not(layer0_outputs(10007));
    outputs(6437) <= not(layer0_outputs(541));
    outputs(6438) <= layer0_outputs(1659);
    outputs(6439) <= not(layer0_outputs(5143));
    outputs(6440) <= not(layer0_outputs(2856)) or (layer0_outputs(6254));
    outputs(6441) <= not(layer0_outputs(3802)) or (layer0_outputs(1638));
    outputs(6442) <= not(layer0_outputs(9566));
    outputs(6443) <= not(layer0_outputs(287)) or (layer0_outputs(1291));
    outputs(6444) <= not(layer0_outputs(6394));
    outputs(6445) <= not(layer0_outputs(5701));
    outputs(6446) <= (layer0_outputs(5210)) and not (layer0_outputs(9844));
    outputs(6447) <= not(layer0_outputs(2810));
    outputs(6448) <= layer0_outputs(325);
    outputs(6449) <= (layer0_outputs(1560)) xor (layer0_outputs(2302));
    outputs(6450) <= not(layer0_outputs(4762)) or (layer0_outputs(1054));
    outputs(6451) <= not(layer0_outputs(8488)) or (layer0_outputs(2813));
    outputs(6452) <= layer0_outputs(7194);
    outputs(6453) <= not((layer0_outputs(1530)) xor (layer0_outputs(2183)));
    outputs(6454) <= not(layer0_outputs(7375));
    outputs(6455) <= (layer0_outputs(8676)) or (layer0_outputs(2875));
    outputs(6456) <= not(layer0_outputs(11));
    outputs(6457) <= (layer0_outputs(4096)) and (layer0_outputs(3316));
    outputs(6458) <= (layer0_outputs(6872)) and not (layer0_outputs(10118));
    outputs(6459) <= not(layer0_outputs(2569));
    outputs(6460) <= (layer0_outputs(7772)) and not (layer0_outputs(4283));
    outputs(6461) <= (layer0_outputs(6085)) xor (layer0_outputs(3886));
    outputs(6462) <= not(layer0_outputs(224));
    outputs(6463) <= (layer0_outputs(6256)) and not (layer0_outputs(1676));
    outputs(6464) <= layer0_outputs(9230);
    outputs(6465) <= not(layer0_outputs(8324));
    outputs(6466) <= not((layer0_outputs(5514)) xor (layer0_outputs(5128)));
    outputs(6467) <= layer0_outputs(7054);
    outputs(6468) <= not(layer0_outputs(1762)) or (layer0_outputs(7864));
    outputs(6469) <= (layer0_outputs(2744)) and not (layer0_outputs(2424));
    outputs(6470) <= not((layer0_outputs(3411)) xor (layer0_outputs(1038)));
    outputs(6471) <= (layer0_outputs(6778)) or (layer0_outputs(6747));
    outputs(6472) <= not((layer0_outputs(9692)) or (layer0_outputs(3104)));
    outputs(6473) <= not(layer0_outputs(4342));
    outputs(6474) <= (layer0_outputs(7767)) or (layer0_outputs(2525));
    outputs(6475) <= (layer0_outputs(6536)) and not (layer0_outputs(10088));
    outputs(6476) <= layer0_outputs(6810);
    outputs(6477) <= layer0_outputs(9760);
    outputs(6478) <= not(layer0_outputs(161));
    outputs(6479) <= not(layer0_outputs(1129));
    outputs(6480) <= not((layer0_outputs(3949)) xor (layer0_outputs(5074)));
    outputs(6481) <= layer0_outputs(7054);
    outputs(6482) <= layer0_outputs(1980);
    outputs(6483) <= (layer0_outputs(7626)) xor (layer0_outputs(7628));
    outputs(6484) <= not((layer0_outputs(8631)) and (layer0_outputs(4815)));
    outputs(6485) <= not(layer0_outputs(9286)) or (layer0_outputs(3839));
    outputs(6486) <= layer0_outputs(49);
    outputs(6487) <= layer0_outputs(3998);
    outputs(6488) <= layer0_outputs(4028);
    outputs(6489) <= not((layer0_outputs(2941)) or (layer0_outputs(1743)));
    outputs(6490) <= layer0_outputs(5830);
    outputs(6491) <= (layer0_outputs(4359)) and not (layer0_outputs(5706));
    outputs(6492) <= (layer0_outputs(259)) xor (layer0_outputs(3936));
    outputs(6493) <= not(layer0_outputs(7606));
    outputs(6494) <= (layer0_outputs(3737)) and not (layer0_outputs(3213));
    outputs(6495) <= not(layer0_outputs(6318));
    outputs(6496) <= not(layer0_outputs(3509)) or (layer0_outputs(10026));
    outputs(6497) <= not((layer0_outputs(8367)) xor (layer0_outputs(7896)));
    outputs(6498) <= not(layer0_outputs(4525));
    outputs(6499) <= layer0_outputs(665);
    outputs(6500) <= layer0_outputs(7764);
    outputs(6501) <= layer0_outputs(6129);
    outputs(6502) <= layer0_outputs(53);
    outputs(6503) <= (layer0_outputs(6011)) and not (layer0_outputs(8834));
    outputs(6504) <= not(layer0_outputs(7324));
    outputs(6505) <= not(layer0_outputs(6131));
    outputs(6506) <= not((layer0_outputs(5232)) or (layer0_outputs(5408)));
    outputs(6507) <= not(layer0_outputs(3215));
    outputs(6508) <= not(layer0_outputs(8899));
    outputs(6509) <= (layer0_outputs(6985)) and not (layer0_outputs(9370));
    outputs(6510) <= (layer0_outputs(7367)) xor (layer0_outputs(8075));
    outputs(6511) <= (layer0_outputs(2110)) and (layer0_outputs(4069));
    outputs(6512) <= (layer0_outputs(3256)) and not (layer0_outputs(1959));
    outputs(6513) <= not(layer0_outputs(5464));
    outputs(6514) <= (layer0_outputs(1000)) and not (layer0_outputs(8772));
    outputs(6515) <= layer0_outputs(4354);
    outputs(6516) <= not(layer0_outputs(7979));
    outputs(6517) <= layer0_outputs(8721);
    outputs(6518) <= not(layer0_outputs(10063));
    outputs(6519) <= layer0_outputs(4670);
    outputs(6520) <= not(layer0_outputs(4464));
    outputs(6521) <= not(layer0_outputs(2338));
    outputs(6522) <= not(layer0_outputs(662));
    outputs(6523) <= layer0_outputs(2967);
    outputs(6524) <= not(layer0_outputs(5512)) or (layer0_outputs(1579));
    outputs(6525) <= not(layer0_outputs(5293));
    outputs(6526) <= not(layer0_outputs(117));
    outputs(6527) <= (layer0_outputs(9699)) and not (layer0_outputs(2075));
    outputs(6528) <= (layer0_outputs(8322)) or (layer0_outputs(5429));
    outputs(6529) <= (layer0_outputs(3914)) xor (layer0_outputs(6801));
    outputs(6530) <= not((layer0_outputs(7194)) xor (layer0_outputs(3772)));
    outputs(6531) <= layer0_outputs(6413);
    outputs(6532) <= not((layer0_outputs(8777)) and (layer0_outputs(2254)));
    outputs(6533) <= not(layer0_outputs(4067));
    outputs(6534) <= layer0_outputs(8769);
    outputs(6535) <= layer0_outputs(5090);
    outputs(6536) <= not(layer0_outputs(6653));
    outputs(6537) <= not(layer0_outputs(5154));
    outputs(6538) <= layer0_outputs(464);
    outputs(6539) <= not(layer0_outputs(861));
    outputs(6540) <= (layer0_outputs(8069)) and not (layer0_outputs(2954));
    outputs(6541) <= (layer0_outputs(5255)) and (layer0_outputs(406));
    outputs(6542) <= not(layer0_outputs(4656));
    outputs(6543) <= layer0_outputs(6846);
    outputs(6544) <= not(layer0_outputs(9698)) or (layer0_outputs(7061));
    outputs(6545) <= not(layer0_outputs(7031));
    outputs(6546) <= not(layer0_outputs(8609));
    outputs(6547) <= (layer0_outputs(1475)) xor (layer0_outputs(558));
    outputs(6548) <= not(layer0_outputs(6134));
    outputs(6549) <= not(layer0_outputs(2337));
    outputs(6550) <= layer0_outputs(3309);
    outputs(6551) <= not(layer0_outputs(6159));
    outputs(6552) <= not((layer0_outputs(7448)) and (layer0_outputs(1310)));
    outputs(6553) <= not((layer0_outputs(2479)) and (layer0_outputs(8439)));
    outputs(6554) <= not(layer0_outputs(745));
    outputs(6555) <= not(layer0_outputs(2833));
    outputs(6556) <= not(layer0_outputs(9488));
    outputs(6557) <= (layer0_outputs(9606)) and (layer0_outputs(8175));
    outputs(6558) <= (layer0_outputs(7695)) xor (layer0_outputs(78));
    outputs(6559) <= not((layer0_outputs(6693)) or (layer0_outputs(4783)));
    outputs(6560) <= not(layer0_outputs(5822)) or (layer0_outputs(5221));
    outputs(6561) <= (layer0_outputs(2239)) xor (layer0_outputs(359));
    outputs(6562) <= not(layer0_outputs(7536));
    outputs(6563) <= not(layer0_outputs(9985));
    outputs(6564) <= not(layer0_outputs(3285));
    outputs(6565) <= not(layer0_outputs(6014));
    outputs(6566) <= not(layer0_outputs(7140));
    outputs(6567) <= layer0_outputs(3741);
    outputs(6568) <= not(layer0_outputs(9972));
    outputs(6569) <= (layer0_outputs(10154)) and not (layer0_outputs(362));
    outputs(6570) <= (layer0_outputs(1892)) xor (layer0_outputs(5625));
    outputs(6571) <= not((layer0_outputs(208)) xor (layer0_outputs(83)));
    outputs(6572) <= (layer0_outputs(783)) and not (layer0_outputs(1136));
    outputs(6573) <= not(layer0_outputs(9899)) or (layer0_outputs(1473));
    outputs(6574) <= layer0_outputs(1742);
    outputs(6575) <= not(layer0_outputs(10110));
    outputs(6576) <= (layer0_outputs(2181)) and not (layer0_outputs(9436));
    outputs(6577) <= layer0_outputs(7199);
    outputs(6578) <= layer0_outputs(5725);
    outputs(6579) <= (layer0_outputs(7093)) and not (layer0_outputs(2194));
    outputs(6580) <= (layer0_outputs(6965)) and (layer0_outputs(4771));
    outputs(6581) <= not(layer0_outputs(9943)) or (layer0_outputs(6479));
    outputs(6582) <= (layer0_outputs(2478)) xor (layer0_outputs(512));
    outputs(6583) <= not(layer0_outputs(6674));
    outputs(6584) <= not((layer0_outputs(6501)) xor (layer0_outputs(107)));
    outputs(6585) <= not(layer0_outputs(10102));
    outputs(6586) <= not(layer0_outputs(8486));
    outputs(6587) <= layer0_outputs(4301);
    outputs(6588) <= not(layer0_outputs(6252));
    outputs(6589) <= layer0_outputs(4225);
    outputs(6590) <= not(layer0_outputs(1099));
    outputs(6591) <= layer0_outputs(7402);
    outputs(6592) <= layer0_outputs(10111);
    outputs(6593) <= (layer0_outputs(3359)) and (layer0_outputs(4595));
    outputs(6594) <= layer0_outputs(2161);
    outputs(6595) <= not((layer0_outputs(3973)) and (layer0_outputs(7186)));
    outputs(6596) <= layer0_outputs(3045);
    outputs(6597) <= not(layer0_outputs(5450)) or (layer0_outputs(7538));
    outputs(6598) <= layer0_outputs(5454);
    outputs(6599) <= layer0_outputs(1773);
    outputs(6600) <= not((layer0_outputs(3996)) or (layer0_outputs(8098)));
    outputs(6601) <= not(layer0_outputs(192));
    outputs(6602) <= not(layer0_outputs(9290)) or (layer0_outputs(8065));
    outputs(6603) <= (layer0_outputs(1854)) and (layer0_outputs(6959));
    outputs(6604) <= (layer0_outputs(3295)) and (layer0_outputs(360));
    outputs(6605) <= layer0_outputs(8673);
    outputs(6606) <= layer0_outputs(7319);
    outputs(6607) <= not((layer0_outputs(2699)) or (layer0_outputs(7156)));
    outputs(6608) <= not((layer0_outputs(5839)) or (layer0_outputs(5687)));
    outputs(6609) <= (layer0_outputs(5420)) and (layer0_outputs(2415));
    outputs(6610) <= (layer0_outputs(1128)) xor (layer0_outputs(5083));
    outputs(6611) <= layer0_outputs(1573);
    outputs(6612) <= (layer0_outputs(5371)) and (layer0_outputs(124));
    outputs(6613) <= layer0_outputs(9915);
    outputs(6614) <= not(layer0_outputs(7625));
    outputs(6615) <= layer0_outputs(7094);
    outputs(6616) <= (layer0_outputs(2480)) and (layer0_outputs(3003));
    outputs(6617) <= not(layer0_outputs(9830));
    outputs(6618) <= not((layer0_outputs(722)) or (layer0_outputs(2098)));
    outputs(6619) <= not(layer0_outputs(9863)) or (layer0_outputs(6036));
    outputs(6620) <= layer0_outputs(8397);
    outputs(6621) <= layer0_outputs(5231);
    outputs(6622) <= not((layer0_outputs(4891)) or (layer0_outputs(6775)));
    outputs(6623) <= not(layer0_outputs(7209));
    outputs(6624) <= not((layer0_outputs(5195)) or (layer0_outputs(7639)));
    outputs(6625) <= layer0_outputs(1736);
    outputs(6626) <= layer0_outputs(9414);
    outputs(6627) <= not(layer0_outputs(2702));
    outputs(6628) <= not(layer0_outputs(2391));
    outputs(6629) <= layer0_outputs(8247);
    outputs(6630) <= not(layer0_outputs(2250));
    outputs(6631) <= (layer0_outputs(1037)) xor (layer0_outputs(4309));
    outputs(6632) <= layer0_outputs(1218);
    outputs(6633) <= not(layer0_outputs(3959));
    outputs(6634) <= layer0_outputs(9142);
    outputs(6635) <= not(layer0_outputs(8382)) or (layer0_outputs(17));
    outputs(6636) <= (layer0_outputs(7064)) and (layer0_outputs(4652));
    outputs(6637) <= (layer0_outputs(2444)) xor (layer0_outputs(1614));
    outputs(6638) <= not(layer0_outputs(5009)) or (layer0_outputs(5656));
    outputs(6639) <= layer0_outputs(6467);
    outputs(6640) <= not(layer0_outputs(390)) or (layer0_outputs(3311));
    outputs(6641) <= not((layer0_outputs(10122)) xor (layer0_outputs(3070)));
    outputs(6642) <= not((layer0_outputs(2339)) or (layer0_outputs(968)));
    outputs(6643) <= not(layer0_outputs(5111)) or (layer0_outputs(9418));
    outputs(6644) <= (layer0_outputs(2777)) xor (layer0_outputs(5515));
    outputs(6645) <= not((layer0_outputs(6454)) xor (layer0_outputs(8636)));
    outputs(6646) <= layer0_outputs(9765);
    outputs(6647) <= (layer0_outputs(5086)) xor (layer0_outputs(557));
    outputs(6648) <= layer0_outputs(5161);
    outputs(6649) <= not(layer0_outputs(6169));
    outputs(6650) <= not((layer0_outputs(9264)) xor (layer0_outputs(10186)));
    outputs(6651) <= not((layer0_outputs(3600)) or (layer0_outputs(5905)));
    outputs(6652) <= not((layer0_outputs(5208)) or (layer0_outputs(7408)));
    outputs(6653) <= (layer0_outputs(723)) xor (layer0_outputs(6959));
    outputs(6654) <= not(layer0_outputs(3431)) or (layer0_outputs(765));
    outputs(6655) <= layer0_outputs(2059);
    outputs(6656) <= layer0_outputs(7183);
    outputs(6657) <= not(layer0_outputs(7379));
    outputs(6658) <= not(layer0_outputs(1789));
    outputs(6659) <= not((layer0_outputs(9908)) and (layer0_outputs(7691)));
    outputs(6660) <= layer0_outputs(7491);
    outputs(6661) <= (layer0_outputs(6898)) and (layer0_outputs(3275));
    outputs(6662) <= not(layer0_outputs(2458));
    outputs(6663) <= not((layer0_outputs(3194)) xor (layer0_outputs(7509)));
    outputs(6664) <= layer0_outputs(6973);
    outputs(6665) <= layer0_outputs(430);
    outputs(6666) <= not(layer0_outputs(2856));
    outputs(6667) <= not(layer0_outputs(8191));
    outputs(6668) <= layer0_outputs(5013);
    outputs(6669) <= layer0_outputs(8775);
    outputs(6670) <= (layer0_outputs(8911)) and not (layer0_outputs(3667));
    outputs(6671) <= (layer0_outputs(1223)) xor (layer0_outputs(5121));
    outputs(6672) <= (layer0_outputs(3617)) and not (layer0_outputs(4653));
    outputs(6673) <= not(layer0_outputs(4655));
    outputs(6674) <= not((layer0_outputs(4753)) xor (layer0_outputs(6671)));
    outputs(6675) <= not(layer0_outputs(8533));
    outputs(6676) <= layer0_outputs(5134);
    outputs(6677) <= layer0_outputs(4544);
    outputs(6678) <= not((layer0_outputs(8509)) or (layer0_outputs(6759)));
    outputs(6679) <= not(layer0_outputs(7018));
    outputs(6680) <= not((layer0_outputs(949)) or (layer0_outputs(6032)));
    outputs(6681) <= not((layer0_outputs(6571)) or (layer0_outputs(2422)));
    outputs(6682) <= not(layer0_outputs(9860)) or (layer0_outputs(6008));
    outputs(6683) <= not((layer0_outputs(7978)) xor (layer0_outputs(6692)));
    outputs(6684) <= not((layer0_outputs(6282)) and (layer0_outputs(9763)));
    outputs(6685) <= not(layer0_outputs(5246)) or (layer0_outputs(5848));
    outputs(6686) <= not(layer0_outputs(2820)) or (layer0_outputs(10048));
    outputs(6687) <= not((layer0_outputs(7235)) or (layer0_outputs(8450)));
    outputs(6688) <= not(layer0_outputs(5937));
    outputs(6689) <= not(layer0_outputs(5171));
    outputs(6690) <= not(layer0_outputs(7777));
    outputs(6691) <= layer0_outputs(629);
    outputs(6692) <= (layer0_outputs(3592)) and (layer0_outputs(2509));
    outputs(6693) <= layer0_outputs(6792);
    outputs(6694) <= not(layer0_outputs(8908));
    outputs(6695) <= not((layer0_outputs(4645)) or (layer0_outputs(3890)));
    outputs(6696) <= (layer0_outputs(5318)) xor (layer0_outputs(8978));
    outputs(6697) <= not(layer0_outputs(4630));
    outputs(6698) <= not(layer0_outputs(7895));
    outputs(6699) <= (layer0_outputs(8706)) or (layer0_outputs(4549));
    outputs(6700) <= (layer0_outputs(19)) xor (layer0_outputs(3228));
    outputs(6701) <= layer0_outputs(4451);
    outputs(6702) <= not((layer0_outputs(9232)) xor (layer0_outputs(1052)));
    outputs(6703) <= not(layer0_outputs(8205)) or (layer0_outputs(4794));
    outputs(6704) <= layer0_outputs(8249);
    outputs(6705) <= (layer0_outputs(3647)) and not (layer0_outputs(5121));
    outputs(6706) <= layer0_outputs(7221);
    outputs(6707) <= not(layer0_outputs(589));
    outputs(6708) <= not((layer0_outputs(6561)) or (layer0_outputs(1548)));
    outputs(6709) <= layer0_outputs(2225);
    outputs(6710) <= not(layer0_outputs(9810));
    outputs(6711) <= not((layer0_outputs(889)) xor (layer0_outputs(6829)));
    outputs(6712) <= not(layer0_outputs(7184));
    outputs(6713) <= not(layer0_outputs(684));
    outputs(6714) <= not(layer0_outputs(4262));
    outputs(6715) <= layer0_outputs(4285);
    outputs(6716) <= layer0_outputs(4928);
    outputs(6717) <= not((layer0_outputs(8758)) or (layer0_outputs(6580)));
    outputs(6718) <= not(layer0_outputs(5866)) or (layer0_outputs(314));
    outputs(6719) <= not(layer0_outputs(3180));
    outputs(6720) <= (layer0_outputs(283)) and not (layer0_outputs(7556));
    outputs(6721) <= layer0_outputs(9786);
    outputs(6722) <= not(layer0_outputs(227));
    outputs(6723) <= (layer0_outputs(2117)) and not (layer0_outputs(5724));
    outputs(6724) <= layer0_outputs(929);
    outputs(6725) <= not(layer0_outputs(5984));
    outputs(6726) <= (layer0_outputs(3897)) and not (layer0_outputs(8708));
    outputs(6727) <= layer0_outputs(804);
    outputs(6728) <= not(layer0_outputs(9365));
    outputs(6729) <= not((layer0_outputs(8773)) xor (layer0_outputs(8914)));
    outputs(6730) <= layer0_outputs(384);
    outputs(6731) <= not(layer0_outputs(6633));
    outputs(6732) <= (layer0_outputs(2188)) and not (layer0_outputs(4884));
    outputs(6733) <= (layer0_outputs(5647)) or (layer0_outputs(940));
    outputs(6734) <= (layer0_outputs(2741)) xor (layer0_outputs(6));
    outputs(6735) <= not((layer0_outputs(7794)) xor (layer0_outputs(5737)));
    outputs(6736) <= not((layer0_outputs(6824)) xor (layer0_outputs(8401)));
    outputs(6737) <= (layer0_outputs(7437)) and not (layer0_outputs(9603));
    outputs(6738) <= not(layer0_outputs(4649));
    outputs(6739) <= not((layer0_outputs(5012)) or (layer0_outputs(10057)));
    outputs(6740) <= (layer0_outputs(4110)) and not (layer0_outputs(6695));
    outputs(6741) <= not(layer0_outputs(3297));
    outputs(6742) <= not(layer0_outputs(1077));
    outputs(6743) <= not(layer0_outputs(7208));
    outputs(6744) <= not(layer0_outputs(74)) or (layer0_outputs(6299));
    outputs(6745) <= not(layer0_outputs(9073));
    outputs(6746) <= not((layer0_outputs(8257)) xor (layer0_outputs(8278)));
    outputs(6747) <= (layer0_outputs(7276)) xor (layer0_outputs(7617));
    outputs(6748) <= not(layer0_outputs(8655));
    outputs(6749) <= not((layer0_outputs(7230)) xor (layer0_outputs(6332)));
    outputs(6750) <= not((layer0_outputs(714)) or (layer0_outputs(10050)));
    outputs(6751) <= (layer0_outputs(10081)) and (layer0_outputs(1090));
    outputs(6752) <= not((layer0_outputs(4401)) and (layer0_outputs(9256)));
    outputs(6753) <= layer0_outputs(450);
    outputs(6754) <= not((layer0_outputs(4188)) xor (layer0_outputs(5301)));
    outputs(6755) <= not((layer0_outputs(3826)) and (layer0_outputs(4058)));
    outputs(6756) <= (layer0_outputs(6191)) and not (layer0_outputs(9914));
    outputs(6757) <= not(layer0_outputs(115)) or (layer0_outputs(9769));
    outputs(6758) <= (layer0_outputs(4829)) xor (layer0_outputs(4229));
    outputs(6759) <= layer0_outputs(8884);
    outputs(6760) <= (layer0_outputs(8388)) and not (layer0_outputs(1645));
    outputs(6761) <= (layer0_outputs(3148)) and not (layer0_outputs(3336));
    outputs(6762) <= not((layer0_outputs(2236)) or (layer0_outputs(6896)));
    outputs(6763) <= layer0_outputs(482);
    outputs(6764) <= not((layer0_outputs(9015)) and (layer0_outputs(661)));
    outputs(6765) <= not(layer0_outputs(6507));
    outputs(6766) <= not((layer0_outputs(3613)) or (layer0_outputs(9276)));
    outputs(6767) <= not((layer0_outputs(6692)) xor (layer0_outputs(4873)));
    outputs(6768) <= not(layer0_outputs(3689));
    outputs(6769) <= not(layer0_outputs(7258));
    outputs(6770) <= not((layer0_outputs(2817)) or (layer0_outputs(2853)));
    outputs(6771) <= not(layer0_outputs(2020));
    outputs(6772) <= not((layer0_outputs(8542)) xor (layer0_outputs(5167)));
    outputs(6773) <= not(layer0_outputs(5831));
    outputs(6774) <= not(layer0_outputs(6456));
    outputs(6775) <= not((layer0_outputs(8652)) or (layer0_outputs(5569)));
    outputs(6776) <= (layer0_outputs(5392)) and (layer0_outputs(6251));
    outputs(6777) <= (layer0_outputs(4713)) xor (layer0_outputs(7591));
    outputs(6778) <= not(layer0_outputs(3757)) or (layer0_outputs(2310));
    outputs(6779) <= not(layer0_outputs(4063)) or (layer0_outputs(6556));
    outputs(6780) <= not(layer0_outputs(7159));
    outputs(6781) <= layer0_outputs(9760);
    outputs(6782) <= layer0_outputs(2751);
    outputs(6783) <= layer0_outputs(6231);
    outputs(6784) <= (layer0_outputs(7309)) and not (layer0_outputs(824));
    outputs(6785) <= (layer0_outputs(3635)) or (layer0_outputs(4561));
    outputs(6786) <= not(layer0_outputs(5390));
    outputs(6787) <= not((layer0_outputs(1111)) xor (layer0_outputs(8005)));
    outputs(6788) <= not((layer0_outputs(1156)) and (layer0_outputs(6619)));
    outputs(6789) <= layer0_outputs(3172);
    outputs(6790) <= (layer0_outputs(9108)) and (layer0_outputs(4110));
    outputs(6791) <= not(layer0_outputs(7020));
    outputs(6792) <= layer0_outputs(3072);
    outputs(6793) <= layer0_outputs(9600);
    outputs(6794) <= not((layer0_outputs(7322)) and (layer0_outputs(1372)));
    outputs(6795) <= not(layer0_outputs(2438));
    outputs(6796) <= not(layer0_outputs(3457));
    outputs(6797) <= not(layer0_outputs(4011)) or (layer0_outputs(1961));
    outputs(6798) <= not(layer0_outputs(8615));
    outputs(6799) <= layer0_outputs(10160);
    outputs(6800) <= (layer0_outputs(7938)) xor (layer0_outputs(4985));
    outputs(6801) <= (layer0_outputs(566)) and (layer0_outputs(6298));
    outputs(6802) <= layer0_outputs(6717);
    outputs(6803) <= not((layer0_outputs(6844)) and (layer0_outputs(5802)));
    outputs(6804) <= not(layer0_outputs(5823));
    outputs(6805) <= layer0_outputs(8830);
    outputs(6806) <= not((layer0_outputs(5863)) xor (layer0_outputs(4636)));
    outputs(6807) <= layer0_outputs(554);
    outputs(6808) <= not((layer0_outputs(9487)) or (layer0_outputs(5328)));
    outputs(6809) <= (layer0_outputs(8864)) xor (layer0_outputs(4985));
    outputs(6810) <= layer0_outputs(8088);
    outputs(6811) <= not((layer0_outputs(8141)) or (layer0_outputs(3044)));
    outputs(6812) <= layer0_outputs(8672);
    outputs(6813) <= not((layer0_outputs(567)) or (layer0_outputs(8237)));
    outputs(6814) <= (layer0_outputs(4959)) and not (layer0_outputs(7257));
    outputs(6815) <= (layer0_outputs(365)) xor (layer0_outputs(9227));
    outputs(6816) <= (layer0_outputs(1352)) xor (layer0_outputs(7978));
    outputs(6817) <= (layer0_outputs(7548)) xor (layer0_outputs(938));
    outputs(6818) <= layer0_outputs(7689);
    outputs(6819) <= not(layer0_outputs(1407));
    outputs(6820) <= (layer0_outputs(627)) xor (layer0_outputs(4492));
    outputs(6821) <= not((layer0_outputs(6688)) and (layer0_outputs(6112)));
    outputs(6822) <= not((layer0_outputs(2050)) and (layer0_outputs(4305)));
    outputs(6823) <= not(layer0_outputs(2710));
    outputs(6824) <= not((layer0_outputs(3832)) or (layer0_outputs(1233)));
    outputs(6825) <= not(layer0_outputs(5686));
    outputs(6826) <= layer0_outputs(3480);
    outputs(6827) <= not((layer0_outputs(9375)) xor (layer0_outputs(2518)));
    outputs(6828) <= (layer0_outputs(461)) xor (layer0_outputs(5676));
    outputs(6829) <= not((layer0_outputs(7980)) xor (layer0_outputs(3325)));
    outputs(6830) <= (layer0_outputs(32)) xor (layer0_outputs(2457));
    outputs(6831) <= layer0_outputs(9675);
    outputs(6832) <= not(layer0_outputs(5509));
    outputs(6833) <= layer0_outputs(9815);
    outputs(6834) <= not(layer0_outputs(6795));
    outputs(6835) <= not(layer0_outputs(8329));
    outputs(6836) <= not((layer0_outputs(489)) xor (layer0_outputs(6947)));
    outputs(6837) <= (layer0_outputs(9135)) and not (layer0_outputs(1016));
    outputs(6838) <= not((layer0_outputs(1725)) or (layer0_outputs(2516)));
    outputs(6839) <= not(layer0_outputs(8991));
    outputs(6840) <= not((layer0_outputs(4936)) xor (layer0_outputs(4039)));
    outputs(6841) <= (layer0_outputs(7887)) and not (layer0_outputs(6565));
    outputs(6842) <= not((layer0_outputs(9991)) and (layer0_outputs(9914)));
    outputs(6843) <= not(layer0_outputs(1652));
    outputs(6844) <= not(layer0_outputs(7854)) or (layer0_outputs(2343));
    outputs(6845) <= not((layer0_outputs(8472)) xor (layer0_outputs(7336)));
    outputs(6846) <= not((layer0_outputs(8375)) xor (layer0_outputs(4990)));
    outputs(6847) <= layer0_outputs(7446);
    outputs(6848) <= (layer0_outputs(2279)) and not (layer0_outputs(347));
    outputs(6849) <= layer0_outputs(3986);
    outputs(6850) <= (layer0_outputs(8253)) or (layer0_outputs(6593));
    outputs(6851) <= not(layer0_outputs(9269));
    outputs(6852) <= layer0_outputs(4470);
    outputs(6853) <= (layer0_outputs(943)) xor (layer0_outputs(2284));
    outputs(6854) <= (layer0_outputs(6507)) xor (layer0_outputs(9350));
    outputs(6855) <= not(layer0_outputs(2205));
    outputs(6856) <= not((layer0_outputs(4536)) or (layer0_outputs(305)));
    outputs(6857) <= not(layer0_outputs(9800));
    outputs(6858) <= layer0_outputs(2697);
    outputs(6859) <= layer0_outputs(8219);
    outputs(6860) <= (layer0_outputs(9253)) and (layer0_outputs(5528));
    outputs(6861) <= layer0_outputs(5279);
    outputs(6862) <= layer0_outputs(9932);
    outputs(6863) <= not(layer0_outputs(489)) or (layer0_outputs(4606));
    outputs(6864) <= (layer0_outputs(5867)) and not (layer0_outputs(6568));
    outputs(6865) <= not(layer0_outputs(9140));
    outputs(6866) <= (layer0_outputs(9869)) and (layer0_outputs(2782));
    outputs(6867) <= layer0_outputs(2996);
    outputs(6868) <= layer0_outputs(2295);
    outputs(6869) <= layer0_outputs(5186);
    outputs(6870) <= layer0_outputs(10180);
    outputs(6871) <= layer0_outputs(1024);
    outputs(6872) <= not(layer0_outputs(7828));
    outputs(6873) <= layer0_outputs(6168);
    outputs(6874) <= layer0_outputs(3521);
    outputs(6875) <= not(layer0_outputs(2853));
    outputs(6876) <= layer0_outputs(2586);
    outputs(6877) <= (layer0_outputs(6384)) and not (layer0_outputs(4218));
    outputs(6878) <= layer0_outputs(7776);
    outputs(6879) <= (layer0_outputs(1518)) and not (layer0_outputs(3191));
    outputs(6880) <= layer0_outputs(363);
    outputs(6881) <= not(layer0_outputs(3049));
    outputs(6882) <= layer0_outputs(2462);
    outputs(6883) <= not(layer0_outputs(6471));
    outputs(6884) <= not(layer0_outputs(712));
    outputs(6885) <= layer0_outputs(3972);
    outputs(6886) <= layer0_outputs(10018);
    outputs(6887) <= (layer0_outputs(6334)) and (layer0_outputs(4441));
    outputs(6888) <= layer0_outputs(5924);
    outputs(6889) <= (layer0_outputs(995)) xor (layer0_outputs(8736));
    outputs(6890) <= layer0_outputs(5694);
    outputs(6891) <= (layer0_outputs(2695)) and not (layer0_outputs(7223));
    outputs(6892) <= layer0_outputs(9758);
    outputs(6893) <= not((layer0_outputs(1995)) and (layer0_outputs(2836)));
    outputs(6894) <= not(layer0_outputs(9784));
    outputs(6895) <= (layer0_outputs(1825)) and not (layer0_outputs(3342));
    outputs(6896) <= not((layer0_outputs(7399)) xor (layer0_outputs(2834)));
    outputs(6897) <= not(layer0_outputs(1974));
    outputs(6898) <= layer0_outputs(9588);
    outputs(6899) <= not(layer0_outputs(4803));
    outputs(6900) <= not(layer0_outputs(1675));
    outputs(6901) <= (layer0_outputs(8680)) and not (layer0_outputs(6849));
    outputs(6902) <= not(layer0_outputs(5188));
    outputs(6903) <= not((layer0_outputs(5347)) or (layer0_outputs(8652)));
    outputs(6904) <= not(layer0_outputs(6714));
    outputs(6905) <= layer0_outputs(2934);
    outputs(6906) <= (layer0_outputs(8363)) xor (layer0_outputs(802));
    outputs(6907) <= layer0_outputs(8273);
    outputs(6908) <= not((layer0_outputs(9615)) or (layer0_outputs(4269)));
    outputs(6909) <= layer0_outputs(8076);
    outputs(6910) <= (layer0_outputs(8855)) and (layer0_outputs(35));
    outputs(6911) <= not(layer0_outputs(1689));
    outputs(6912) <= (layer0_outputs(6256)) and not (layer0_outputs(787));
    outputs(6913) <= not(layer0_outputs(3962));
    outputs(6914) <= layer0_outputs(9088);
    outputs(6915) <= not((layer0_outputs(3190)) or (layer0_outputs(1469)));
    outputs(6916) <= layer0_outputs(3529);
    outputs(6917) <= not(layer0_outputs(5978));
    outputs(6918) <= not(layer0_outputs(8572));
    outputs(6919) <= not((layer0_outputs(9522)) or (layer0_outputs(4457)));
    outputs(6920) <= not(layer0_outputs(8722));
    outputs(6921) <= not(layer0_outputs(5393));
    outputs(6922) <= layer0_outputs(601);
    outputs(6923) <= not(layer0_outputs(2804));
    outputs(6924) <= (layer0_outputs(5127)) xor (layer0_outputs(6051));
    outputs(6925) <= (layer0_outputs(2340)) and not (layer0_outputs(6694));
    outputs(6926) <= not(layer0_outputs(9819));
    outputs(6927) <= not(layer0_outputs(7914)) or (layer0_outputs(7697));
    outputs(6928) <= layer0_outputs(10061);
    outputs(6929) <= layer0_outputs(8515);
    outputs(6930) <= (layer0_outputs(500)) and not (layer0_outputs(7276));
    outputs(6931) <= not((layer0_outputs(1042)) or (layer0_outputs(6994)));
    outputs(6932) <= (layer0_outputs(3557)) and not (layer0_outputs(10203));
    outputs(6933) <= (layer0_outputs(3734)) and not (layer0_outputs(10168));
    outputs(6934) <= not((layer0_outputs(4514)) xor (layer0_outputs(753)));
    outputs(6935) <= not(layer0_outputs(8130)) or (layer0_outputs(1918));
    outputs(6936) <= layer0_outputs(891);
    outputs(6937) <= layer0_outputs(5844);
    outputs(6938) <= layer0_outputs(8199);
    outputs(6939) <= layer0_outputs(8360);
    outputs(6940) <= layer0_outputs(9921);
    outputs(6941) <= not((layer0_outputs(7586)) or (layer0_outputs(3258)));
    outputs(6942) <= not((layer0_outputs(6444)) and (layer0_outputs(7362)));
    outputs(6943) <= layer0_outputs(7091);
    outputs(6944) <= not(layer0_outputs(593));
    outputs(6945) <= layer0_outputs(9532);
    outputs(6946) <= (layer0_outputs(1735)) and not (layer0_outputs(4778));
    outputs(6947) <= not(layer0_outputs(8842));
    outputs(6948) <= not(layer0_outputs(1893));
    outputs(6949) <= (layer0_outputs(2542)) and (layer0_outputs(3727));
    outputs(6950) <= layer0_outputs(6728);
    outputs(6951) <= (layer0_outputs(9964)) and not (layer0_outputs(2707));
    outputs(6952) <= layer0_outputs(5738);
    outputs(6953) <= not(layer0_outputs(2350));
    outputs(6954) <= layer0_outputs(4112);
    outputs(6955) <= not(layer0_outputs(4224));
    outputs(6956) <= not(layer0_outputs(1377));
    outputs(6957) <= layer0_outputs(10129);
    outputs(6958) <= not(layer0_outputs(564));
    outputs(6959) <= layer0_outputs(3380);
    outputs(6960) <= not(layer0_outputs(9460));
    outputs(6961) <= (layer0_outputs(4575)) and not (layer0_outputs(7845));
    outputs(6962) <= not(layer0_outputs(1491));
    outputs(6963) <= layer0_outputs(5764);
    outputs(6964) <= (layer0_outputs(5693)) and (layer0_outputs(360));
    outputs(6965) <= not((layer0_outputs(6772)) xor (layer0_outputs(5191)));
    outputs(6966) <= not((layer0_outputs(3390)) or (layer0_outputs(238)));
    outputs(6967) <= layer0_outputs(4717);
    outputs(6968) <= not((layer0_outputs(878)) or (layer0_outputs(1715)));
    outputs(6969) <= (layer0_outputs(6232)) xor (layer0_outputs(3960));
    outputs(6970) <= (layer0_outputs(3177)) and (layer0_outputs(9869));
    outputs(6971) <= layer0_outputs(6792);
    outputs(6972) <= not((layer0_outputs(4808)) xor (layer0_outputs(1254)));
    outputs(6973) <= layer0_outputs(6746);
    outputs(6974) <= not(layer0_outputs(9670));
    outputs(6975) <= not(layer0_outputs(2622));
    outputs(6976) <= not(layer0_outputs(7355));
    outputs(6977) <= layer0_outputs(3140);
    outputs(6978) <= layer0_outputs(7709);
    outputs(6979) <= (layer0_outputs(9357)) and (layer0_outputs(5397));
    outputs(6980) <= (layer0_outputs(2944)) and (layer0_outputs(7878));
    outputs(6981) <= not(layer0_outputs(5534));
    outputs(6982) <= not(layer0_outputs(8353));
    outputs(6983) <= layer0_outputs(7034);
    outputs(6984) <= not(layer0_outputs(2701));
    outputs(6985) <= layer0_outputs(3379);
    outputs(6986) <= not(layer0_outputs(833));
    outputs(6987) <= not(layer0_outputs(1066));
    outputs(6988) <= (layer0_outputs(2588)) xor (layer0_outputs(2098));
    outputs(6989) <= not((layer0_outputs(1879)) or (layer0_outputs(2477)));
    outputs(6990) <= layer0_outputs(6646);
    outputs(6991) <= (layer0_outputs(2881)) and not (layer0_outputs(5724));
    outputs(6992) <= not(layer0_outputs(5345));
    outputs(6993) <= layer0_outputs(9098);
    outputs(6994) <= (layer0_outputs(7307)) and not (layer0_outputs(9660));
    outputs(6995) <= not(layer0_outputs(9547));
    outputs(6996) <= layer0_outputs(1807);
    outputs(6997) <= not(layer0_outputs(3544));
    outputs(6998) <= layer0_outputs(6012);
    outputs(6999) <= not((layer0_outputs(6770)) and (layer0_outputs(3156)));
    outputs(7000) <= layer0_outputs(13);
    outputs(7001) <= not(layer0_outputs(3843));
    outputs(7002) <= layer0_outputs(10081);
    outputs(7003) <= not(layer0_outputs(2254));
    outputs(7004) <= (layer0_outputs(6962)) and not (layer0_outputs(447));
    outputs(7005) <= not(layer0_outputs(4877));
    outputs(7006) <= not((layer0_outputs(5394)) xor (layer0_outputs(432)));
    outputs(7007) <= layer0_outputs(7524);
    outputs(7008) <= not(layer0_outputs(2921));
    outputs(7009) <= layer0_outputs(7027);
    outputs(7010) <= not(layer0_outputs(1476)) or (layer0_outputs(3798));
    outputs(7011) <= not(layer0_outputs(7154));
    outputs(7012) <= not(layer0_outputs(1709));
    outputs(7013) <= layer0_outputs(9875);
    outputs(7014) <= layer0_outputs(4075);
    outputs(7015) <= (layer0_outputs(3149)) and not (layer0_outputs(9587));
    outputs(7016) <= not((layer0_outputs(9968)) or (layer0_outputs(3249)));
    outputs(7017) <= not(layer0_outputs(10172));
    outputs(7018) <= not(layer0_outputs(7904));
    outputs(7019) <= layer0_outputs(2573);
    outputs(7020) <= not(layer0_outputs(3536));
    outputs(7021) <= not((layer0_outputs(6048)) xor (layer0_outputs(9093)));
    outputs(7022) <= not(layer0_outputs(10179));
    outputs(7023) <= not(layer0_outputs(1727));
    outputs(7024) <= not(layer0_outputs(809));
    outputs(7025) <= not(layer0_outputs(5246));
    outputs(7026) <= not(layer0_outputs(498)) or (layer0_outputs(9038));
    outputs(7027) <= not((layer0_outputs(2012)) xor (layer0_outputs(538)));
    outputs(7028) <= layer0_outputs(234);
    outputs(7029) <= not(layer0_outputs(3227));
    outputs(7030) <= not(layer0_outputs(9315));
    outputs(7031) <= not((layer0_outputs(4613)) or (layer0_outputs(6657)));
    outputs(7032) <= not(layer0_outputs(5245));
    outputs(7033) <= (layer0_outputs(5755)) xor (layer0_outputs(4478));
    outputs(7034) <= (layer0_outputs(9459)) and not (layer0_outputs(8577));
    outputs(7035) <= (layer0_outputs(4562)) and (layer0_outputs(970));
    outputs(7036) <= not(layer0_outputs(4926));
    outputs(7037) <= not(layer0_outputs(3886));
    outputs(7038) <= not(layer0_outputs(4857));
    outputs(7039) <= not(layer0_outputs(6804));
    outputs(7040) <= layer0_outputs(7780);
    outputs(7041) <= not(layer0_outputs(9107));
    outputs(7042) <= (layer0_outputs(7501)) and not (layer0_outputs(7526));
    outputs(7043) <= layer0_outputs(7570);
    outputs(7044) <= (layer0_outputs(1778)) and not (layer0_outputs(5697));
    outputs(7045) <= (layer0_outputs(6933)) xor (layer0_outputs(10198));
    outputs(7046) <= layer0_outputs(1648);
    outputs(7047) <= not(layer0_outputs(8975));
    outputs(7048) <= not(layer0_outputs(9578));
    outputs(7049) <= not((layer0_outputs(9384)) or (layer0_outputs(1263)));
    outputs(7050) <= not(layer0_outputs(6628));
    outputs(7051) <= not(layer0_outputs(2438));
    outputs(7052) <= layer0_outputs(2132);
    outputs(7053) <= not(layer0_outputs(5330));
    outputs(7054) <= layer0_outputs(2037);
    outputs(7055) <= not(layer0_outputs(5493));
    outputs(7056) <= layer0_outputs(4970);
    outputs(7057) <= layer0_outputs(5725);
    outputs(7058) <= not(layer0_outputs(3856));
    outputs(7059) <= (layer0_outputs(4530)) and not (layer0_outputs(3403));
    outputs(7060) <= layer0_outputs(3144);
    outputs(7061) <= not(layer0_outputs(2933));
    outputs(7062) <= not(layer0_outputs(3198)) or (layer0_outputs(5741));
    outputs(7063) <= (layer0_outputs(654)) and (layer0_outputs(8283));
    outputs(7064) <= not(layer0_outputs(7935));
    outputs(7065) <= layer0_outputs(3840);
    outputs(7066) <= layer0_outputs(3485);
    outputs(7067) <= layer0_outputs(7584);
    outputs(7068) <= layer0_outputs(5040);
    outputs(7069) <= layer0_outputs(3163);
    outputs(7070) <= not((layer0_outputs(5478)) or (layer0_outputs(1608)));
    outputs(7071) <= not(layer0_outputs(1826));
    outputs(7072) <= layer0_outputs(1259);
    outputs(7073) <= layer0_outputs(5927);
    outputs(7074) <= layer0_outputs(3687);
    outputs(7075) <= layer0_outputs(1480);
    outputs(7076) <= not(layer0_outputs(4195));
    outputs(7077) <= layer0_outputs(6654);
    outputs(7078) <= not((layer0_outputs(6076)) xor (layer0_outputs(6748)));
    outputs(7079) <= not(layer0_outputs(9127));
    outputs(7080) <= (layer0_outputs(10162)) xor (layer0_outputs(769));
    outputs(7081) <= not(layer0_outputs(7266));
    outputs(7082) <= (layer0_outputs(5263)) and not (layer0_outputs(9229));
    outputs(7083) <= not(layer0_outputs(6658));
    outputs(7084) <= not(layer0_outputs(9865));
    outputs(7085) <= not((layer0_outputs(3387)) xor (layer0_outputs(5702)));
    outputs(7086) <= layer0_outputs(6250);
    outputs(7087) <= not(layer0_outputs(455)) or (layer0_outputs(1474));
    outputs(7088) <= (layer0_outputs(8712)) and not (layer0_outputs(8688));
    outputs(7089) <= not(layer0_outputs(190));
    outputs(7090) <= layer0_outputs(7282);
    outputs(7091) <= (layer0_outputs(7172)) and not (layer0_outputs(3774));
    outputs(7092) <= not(layer0_outputs(1687));
    outputs(7093) <= layer0_outputs(5747);
    outputs(7094) <= layer0_outputs(428);
    outputs(7095) <= not((layer0_outputs(3671)) xor (layer0_outputs(1720)));
    outputs(7096) <= not(layer0_outputs(5572));
    outputs(7097) <= not((layer0_outputs(1064)) or (layer0_outputs(3377)));
    outputs(7098) <= not(layer0_outputs(9774));
    outputs(7099) <= layer0_outputs(4764);
    outputs(7100) <= layer0_outputs(8279);
    outputs(7101) <= layer0_outputs(1162);
    outputs(7102) <= layer0_outputs(689);
    outputs(7103) <= not(layer0_outputs(10006));
    outputs(7104) <= not(layer0_outputs(9924));
    outputs(7105) <= not((layer0_outputs(287)) xor (layer0_outputs(3064)));
    outputs(7106) <= layer0_outputs(141);
    outputs(7107) <= layer0_outputs(5830);
    outputs(7108) <= not(layer0_outputs(10051));
    outputs(7109) <= (layer0_outputs(10119)) xor (layer0_outputs(3478));
    outputs(7110) <= (layer0_outputs(450)) and not (layer0_outputs(7238));
    outputs(7111) <= (layer0_outputs(9518)) and not (layer0_outputs(9386));
    outputs(7112) <= layer0_outputs(9251);
    outputs(7113) <= (layer0_outputs(4756)) and not (layer0_outputs(717));
    outputs(7114) <= layer0_outputs(1980);
    outputs(7115) <= layer0_outputs(1952);
    outputs(7116) <= (layer0_outputs(3409)) and (layer0_outputs(5254));
    outputs(7117) <= not(layer0_outputs(7376));
    outputs(7118) <= not((layer0_outputs(9316)) and (layer0_outputs(6485)));
    outputs(7119) <= (layer0_outputs(6890)) and (layer0_outputs(3681));
    outputs(7120) <= not(layer0_outputs(6602)) or (layer0_outputs(2488));
    outputs(7121) <= layer0_outputs(3130);
    outputs(7122) <= not(layer0_outputs(5302)) or (layer0_outputs(5213));
    outputs(7123) <= not(layer0_outputs(4490));
    outputs(7124) <= not(layer0_outputs(997));
    outputs(7125) <= not(layer0_outputs(2806)) or (layer0_outputs(7666));
    outputs(7126) <= not(layer0_outputs(5081));
    outputs(7127) <= not(layer0_outputs(1326)) or (layer0_outputs(1140));
    outputs(7128) <= layer0_outputs(4437);
    outputs(7129) <= layer0_outputs(8694);
    outputs(7130) <= not(layer0_outputs(7313));
    outputs(7131) <= layer0_outputs(8173);
    outputs(7132) <= (layer0_outputs(361)) xor (layer0_outputs(7482));
    outputs(7133) <= (layer0_outputs(5148)) or (layer0_outputs(6807));
    outputs(7134) <= (layer0_outputs(8065)) and (layer0_outputs(8));
    outputs(7135) <= layer0_outputs(3754);
    outputs(7136) <= not((layer0_outputs(825)) or (layer0_outputs(1971)));
    outputs(7137) <= layer0_outputs(2816);
    outputs(7138) <= not((layer0_outputs(6459)) or (layer0_outputs(981)));
    outputs(7139) <= (layer0_outputs(7553)) or (layer0_outputs(9585));
    outputs(7140) <= (layer0_outputs(1210)) and not (layer0_outputs(1587));
    outputs(7141) <= (layer0_outputs(9707)) and not (layer0_outputs(946));
    outputs(7142) <= not(layer0_outputs(4085));
    outputs(7143) <= not((layer0_outputs(5970)) xor (layer0_outputs(1617)));
    outputs(7144) <= layer0_outputs(3983);
    outputs(7145) <= (layer0_outputs(1966)) and not (layer0_outputs(2790));
    outputs(7146) <= layer0_outputs(6010);
    outputs(7147) <= (layer0_outputs(852)) and (layer0_outputs(8844));
    outputs(7148) <= not(layer0_outputs(1387));
    outputs(7149) <= not(layer0_outputs(708));
    outputs(7150) <= not(layer0_outputs(2459));
    outputs(7151) <= not((layer0_outputs(3984)) and (layer0_outputs(2437)));
    outputs(7152) <= (layer0_outputs(1330)) and (layer0_outputs(8886));
    outputs(7153) <= layer0_outputs(9310);
    outputs(7154) <= layer0_outputs(9679);
    outputs(7155) <= layer0_outputs(8773);
    outputs(7156) <= not(layer0_outputs(5961));
    outputs(7157) <= layer0_outputs(4590);
    outputs(7158) <= (layer0_outputs(1925)) xor (layer0_outputs(2489));
    outputs(7159) <= layer0_outputs(3986);
    outputs(7160) <= layer0_outputs(1332);
    outputs(7161) <= (layer0_outputs(6728)) xor (layer0_outputs(2846));
    outputs(7162) <= not(layer0_outputs(7041));
    outputs(7163) <= (layer0_outputs(3693)) xor (layer0_outputs(9957));
    outputs(7164) <= not((layer0_outputs(3275)) xor (layer0_outputs(9861)));
    outputs(7165) <= not((layer0_outputs(2408)) and (layer0_outputs(4906)));
    outputs(7166) <= (layer0_outputs(3574)) xor (layer0_outputs(1843));
    outputs(7167) <= (layer0_outputs(3280)) and not (layer0_outputs(6150));
    outputs(7168) <= not(layer0_outputs(3034));
    outputs(7169) <= layer0_outputs(666);
    outputs(7170) <= layer0_outputs(7574);
    outputs(7171) <= not(layer0_outputs(2590)) or (layer0_outputs(303));
    outputs(7172) <= not(layer0_outputs(8204));
    outputs(7173) <= layer0_outputs(7763);
    outputs(7174) <= not(layer0_outputs(2372));
    outputs(7175) <= (layer0_outputs(2383)) and not (layer0_outputs(7286));
    outputs(7176) <= layer0_outputs(1602);
    outputs(7177) <= not(layer0_outputs(9977));
    outputs(7178) <= not((layer0_outputs(9720)) xor (layer0_outputs(8358)));
    outputs(7179) <= (layer0_outputs(9506)) and not (layer0_outputs(9754));
    outputs(7180) <= not(layer0_outputs(7523));
    outputs(7181) <= layer0_outputs(10133);
    outputs(7182) <= (layer0_outputs(2337)) and (layer0_outputs(477));
    outputs(7183) <= layer0_outputs(4103);
    outputs(7184) <= layer0_outputs(4443);
    outputs(7185) <= layer0_outputs(3537);
    outputs(7186) <= not((layer0_outputs(9014)) or (layer0_outputs(6957)));
    outputs(7187) <= not((layer0_outputs(7299)) xor (layer0_outputs(856)));
    outputs(7188) <= not(layer0_outputs(3732));
    outputs(7189) <= not(layer0_outputs(4187));
    outputs(7190) <= (layer0_outputs(3556)) and not (layer0_outputs(2447));
    outputs(7191) <= not(layer0_outputs(8873));
    outputs(7192) <= (layer0_outputs(9362)) and not (layer0_outputs(2540));
    outputs(7193) <= (layer0_outputs(5630)) and not (layer0_outputs(5573));
    outputs(7194) <= (layer0_outputs(3216)) and not (layer0_outputs(6519));
    outputs(7195) <= layer0_outputs(4541);
    outputs(7196) <= layer0_outputs(3883);
    outputs(7197) <= (layer0_outputs(6789)) and not (layer0_outputs(6676));
    outputs(7198) <= layer0_outputs(7601);
    outputs(7199) <= layer0_outputs(9212);
    outputs(7200) <= not((layer0_outputs(2391)) xor (layer0_outputs(4106)));
    outputs(7201) <= layer0_outputs(5171);
    outputs(7202) <= not(layer0_outputs(1874));
    outputs(7203) <= layer0_outputs(462);
    outputs(7204) <= layer0_outputs(244);
    outputs(7205) <= (layer0_outputs(5073)) or (layer0_outputs(8583));
    outputs(7206) <= (layer0_outputs(8213)) xor (layer0_outputs(4754));
    outputs(7207) <= not((layer0_outputs(3598)) xor (layer0_outputs(382)));
    outputs(7208) <= (layer0_outputs(9688)) xor (layer0_outputs(2743));
    outputs(7209) <= not((layer0_outputs(2160)) xor (layer0_outputs(7497)));
    outputs(7210) <= not(layer0_outputs(3681));
    outputs(7211) <= layer0_outputs(6797);
    outputs(7212) <= not(layer0_outputs(10115));
    outputs(7213) <= layer0_outputs(6034);
    outputs(7214) <= layer0_outputs(4723);
    outputs(7215) <= not(layer0_outputs(9621)) or (layer0_outputs(1701));
    outputs(7216) <= (layer0_outputs(651)) xor (layer0_outputs(5076));
    outputs(7217) <= not(layer0_outputs(6249)) or (layer0_outputs(975));
    outputs(7218) <= layer0_outputs(1147);
    outputs(7219) <= (layer0_outputs(7851)) or (layer0_outputs(2497));
    outputs(7220) <= not((layer0_outputs(7866)) xor (layer0_outputs(4159)));
    outputs(7221) <= layer0_outputs(9427);
    outputs(7222) <= (layer0_outputs(4385)) xor (layer0_outputs(3703));
    outputs(7223) <= layer0_outputs(4947);
    outputs(7224) <= (layer0_outputs(6990)) and not (layer0_outputs(1345));
    outputs(7225) <= (layer0_outputs(6663)) xor (layer0_outputs(4792));
    outputs(7226) <= (layer0_outputs(4335)) and not (layer0_outputs(9490));
    outputs(7227) <= not(layer0_outputs(3654));
    outputs(7228) <= (layer0_outputs(1575)) and not (layer0_outputs(1408));
    outputs(7229) <= not(layer0_outputs(9762));
    outputs(7230) <= (layer0_outputs(6333)) or (layer0_outputs(6515));
    outputs(7231) <= (layer0_outputs(4912)) xor (layer0_outputs(3878));
    outputs(7232) <= not(layer0_outputs(7196)) or (layer0_outputs(6201));
    outputs(7233) <= not(layer0_outputs(9341));
    outputs(7234) <= not((layer0_outputs(885)) xor (layer0_outputs(3846)));
    outputs(7235) <= (layer0_outputs(7025)) or (layer0_outputs(4905));
    outputs(7236) <= not((layer0_outputs(3859)) or (layer0_outputs(5371)));
    outputs(7237) <= (layer0_outputs(4419)) and (layer0_outputs(637));
    outputs(7238) <= layer0_outputs(5783);
    outputs(7239) <= layer0_outputs(9928);
    outputs(7240) <= not(layer0_outputs(1239));
    outputs(7241) <= (layer0_outputs(6002)) and not (layer0_outputs(3219));
    outputs(7242) <= (layer0_outputs(1309)) and (layer0_outputs(10074));
    outputs(7243) <= (layer0_outputs(6542)) xor (layer0_outputs(3098));
    outputs(7244) <= not((layer0_outputs(2633)) or (layer0_outputs(1211)));
    outputs(7245) <= (layer0_outputs(8996)) and not (layer0_outputs(7151));
    outputs(7246) <= not((layer0_outputs(3907)) or (layer0_outputs(4768)));
    outputs(7247) <= not(layer0_outputs(10190)) or (layer0_outputs(6802));
    outputs(7248) <= (layer0_outputs(4399)) or (layer0_outputs(4609));
    outputs(7249) <= not((layer0_outputs(9142)) xor (layer0_outputs(2889)));
    outputs(7250) <= layer0_outputs(8004);
    outputs(7251) <= not((layer0_outputs(9685)) xor (layer0_outputs(5084)));
    outputs(7252) <= not(layer0_outputs(6852));
    outputs(7253) <= not(layer0_outputs(4010)) or (layer0_outputs(9087));
    outputs(7254) <= not(layer0_outputs(8531)) or (layer0_outputs(5804));
    outputs(7255) <= not(layer0_outputs(2362));
    outputs(7256) <= not(layer0_outputs(8402));
    outputs(7257) <= not(layer0_outputs(6793));
    outputs(7258) <= not(layer0_outputs(6263));
    outputs(7259) <= (layer0_outputs(4162)) and (layer0_outputs(1091));
    outputs(7260) <= (layer0_outputs(2375)) and (layer0_outputs(3853));
    outputs(7261) <= (layer0_outputs(1568)) and not (layer0_outputs(2500));
    outputs(7262) <= (layer0_outputs(4264)) xor (layer0_outputs(456));
    outputs(7263) <= (layer0_outputs(8363)) and not (layer0_outputs(6418));
    outputs(7264) <= (layer0_outputs(4222)) xor (layer0_outputs(6961));
    outputs(7265) <= (layer0_outputs(3829)) and not (layer0_outputs(9154));
    outputs(7266) <= layer0_outputs(5869);
    outputs(7267) <= (layer0_outputs(1237)) and not (layer0_outputs(4967));
    outputs(7268) <= layer0_outputs(7715);
    outputs(7269) <= (layer0_outputs(1860)) and (layer0_outputs(5745));
    outputs(7270) <= not((layer0_outputs(1023)) xor (layer0_outputs(27)));
    outputs(7271) <= layer0_outputs(7101);
    outputs(7272) <= (layer0_outputs(7520)) xor (layer0_outputs(10125));
    outputs(7273) <= layer0_outputs(5111);
    outputs(7274) <= not(layer0_outputs(4488));
    outputs(7275) <= (layer0_outputs(5821)) xor (layer0_outputs(8827));
    outputs(7276) <= layer0_outputs(254);
    outputs(7277) <= layer0_outputs(571);
    outputs(7278) <= not((layer0_outputs(8413)) and (layer0_outputs(8280)));
    outputs(7279) <= not((layer0_outputs(6308)) xor (layer0_outputs(9224)));
    outputs(7280) <= (layer0_outputs(1189)) or (layer0_outputs(5465));
    outputs(7281) <= (layer0_outputs(8738)) and (layer0_outputs(3898));
    outputs(7282) <= (layer0_outputs(2383)) and not (layer0_outputs(4470));
    outputs(7283) <= (layer0_outputs(7226)) and not (layer0_outputs(9596));
    outputs(7284) <= (layer0_outputs(3403)) and not (layer0_outputs(8913));
    outputs(7285) <= not((layer0_outputs(5028)) and (layer0_outputs(7006)));
    outputs(7286) <= layer0_outputs(6341);
    outputs(7287) <= not((layer0_outputs(4071)) xor (layer0_outputs(8439)));
    outputs(7288) <= not(layer0_outputs(4163));
    outputs(7289) <= layer0_outputs(9306);
    outputs(7290) <= not(layer0_outputs(5916));
    outputs(7291) <= not(layer0_outputs(4682));
    outputs(7292) <= not(layer0_outputs(6255));
    outputs(7293) <= not(layer0_outputs(9882));
    outputs(7294) <= not((layer0_outputs(8123)) and (layer0_outputs(9513)));
    outputs(7295) <= layer0_outputs(7320);
    outputs(7296) <= (layer0_outputs(5905)) xor (layer0_outputs(3751));
    outputs(7297) <= not(layer0_outputs(6396));
    outputs(7298) <= (layer0_outputs(936)) and not (layer0_outputs(9243));
    outputs(7299) <= layer0_outputs(9925);
    outputs(7300) <= not((layer0_outputs(10024)) and (layer0_outputs(2544)));
    outputs(7301) <= not(layer0_outputs(978));
    outputs(7302) <= not((layer0_outputs(2508)) or (layer0_outputs(3649)));
    outputs(7303) <= (layer0_outputs(5645)) xor (layer0_outputs(5333));
    outputs(7304) <= not(layer0_outputs(1437));
    outputs(7305) <= layer0_outputs(3245);
    outputs(7306) <= (layer0_outputs(9386)) or (layer0_outputs(4566));
    outputs(7307) <= layer0_outputs(6513);
    outputs(7308) <= not((layer0_outputs(5075)) or (layer0_outputs(583)));
    outputs(7309) <= not(layer0_outputs(5057)) or (layer0_outputs(1274));
    outputs(7310) <= (layer0_outputs(4638)) and not (layer0_outputs(3491));
    outputs(7311) <= not((layer0_outputs(1504)) or (layer0_outputs(9875)));
    outputs(7312) <= not(layer0_outputs(1786));
    outputs(7313) <= not(layer0_outputs(8788));
    outputs(7314) <= not(layer0_outputs(5779));
    outputs(7315) <= layer0_outputs(5449);
    outputs(7316) <= (layer0_outputs(3783)) and not (layer0_outputs(5203));
    outputs(7317) <= not(layer0_outputs(401));
    outputs(7318) <= (layer0_outputs(6065)) xor (layer0_outputs(1144));
    outputs(7319) <= not(layer0_outputs(3657));
    outputs(7320) <= layer0_outputs(9894);
    outputs(7321) <= not(layer0_outputs(2712));
    outputs(7322) <= not(layer0_outputs(2916));
    outputs(7323) <= layer0_outputs(6466);
    outputs(7324) <= (layer0_outputs(4762)) and not (layer0_outputs(4922));
    outputs(7325) <= layer0_outputs(3119);
    outputs(7326) <= not(layer0_outputs(6339));
    outputs(7327) <= not(layer0_outputs(7782));
    outputs(7328) <= layer0_outputs(6092);
    outputs(7329) <= layer0_outputs(3642);
    outputs(7330) <= (layer0_outputs(7405)) and not (layer0_outputs(5649));
    outputs(7331) <= not(layer0_outputs(1631));
    outputs(7332) <= layer0_outputs(10012);
    outputs(7333) <= layer0_outputs(8850);
    outputs(7334) <= (layer0_outputs(1965)) or (layer0_outputs(8740));
    outputs(7335) <= not(layer0_outputs(6058));
    outputs(7336) <= layer0_outputs(1125);
    outputs(7337) <= (layer0_outputs(6387)) xor (layer0_outputs(3858));
    outputs(7338) <= not(layer0_outputs(5666));
    outputs(7339) <= layer0_outputs(1741);
    outputs(7340) <= layer0_outputs(6817);
    outputs(7341) <= not((layer0_outputs(2178)) or (layer0_outputs(1477)));
    outputs(7342) <= (layer0_outputs(7321)) and not (layer0_outputs(5488));
    outputs(7343) <= not((layer0_outputs(449)) xor (layer0_outputs(5960)));
    outputs(7344) <= not((layer0_outputs(6742)) or (layer0_outputs(9534)));
    outputs(7345) <= layer0_outputs(3780);
    outputs(7346) <= not((layer0_outputs(6451)) xor (layer0_outputs(6245)));
    outputs(7347) <= not((layer0_outputs(8428)) xor (layer0_outputs(9979)));
    outputs(7348) <= (layer0_outputs(8067)) xor (layer0_outputs(3227));
    outputs(7349) <= layer0_outputs(7937);
    outputs(7350) <= not(layer0_outputs(2223)) or (layer0_outputs(5925));
    outputs(7351) <= (layer0_outputs(4881)) and not (layer0_outputs(9200));
    outputs(7352) <= (layer0_outputs(6741)) xor (layer0_outputs(7651));
    outputs(7353) <= (layer0_outputs(514)) or (layer0_outputs(3938));
    outputs(7354) <= not(layer0_outputs(2121));
    outputs(7355) <= not(layer0_outputs(7817));
    outputs(7356) <= (layer0_outputs(8874)) or (layer0_outputs(3001));
    outputs(7357) <= (layer0_outputs(7378)) and (layer0_outputs(2670));
    outputs(7358) <= not(layer0_outputs(6803));
    outputs(7359) <= (layer0_outputs(550)) and (layer0_outputs(7830));
    outputs(7360) <= (layer0_outputs(5306)) and (layer0_outputs(7182));
    outputs(7361) <= not((layer0_outputs(105)) and (layer0_outputs(30)));
    outputs(7362) <= (layer0_outputs(3935)) and not (layer0_outputs(6213));
    outputs(7363) <= (layer0_outputs(106)) and not (layer0_outputs(9682));
    outputs(7364) <= (layer0_outputs(6009)) and not (layer0_outputs(2449));
    outputs(7365) <= not((layer0_outputs(8915)) xor (layer0_outputs(2783)));
    outputs(7366) <= layer0_outputs(7891);
    outputs(7367) <= not((layer0_outputs(7583)) xor (layer0_outputs(8492)));
    outputs(7368) <= not(layer0_outputs(3867));
    outputs(7369) <= (layer0_outputs(9319)) and not (layer0_outputs(6987));
    outputs(7370) <= not((layer0_outputs(5760)) xor (layer0_outputs(964)));
    outputs(7371) <= layer0_outputs(9684);
    outputs(7372) <= (layer0_outputs(6661)) and (layer0_outputs(1191));
    outputs(7373) <= (layer0_outputs(526)) and not (layer0_outputs(540));
    outputs(7374) <= (layer0_outputs(8166)) xor (layer0_outputs(7092));
    outputs(7375) <= (layer0_outputs(2246)) xor (layer0_outputs(6461));
    outputs(7376) <= layer0_outputs(4361);
    outputs(7377) <= layer0_outputs(1663);
    outputs(7378) <= (layer0_outputs(463)) xor (layer0_outputs(9718));
    outputs(7379) <= not(layer0_outputs(8491));
    outputs(7380) <= not((layer0_outputs(4577)) or (layer0_outputs(2958)));
    outputs(7381) <= (layer0_outputs(4961)) and not (layer0_outputs(2623));
    outputs(7382) <= '0';
    outputs(7383) <= not(layer0_outputs(8208));
    outputs(7384) <= (layer0_outputs(5665)) and not (layer0_outputs(1588));
    outputs(7385) <= not(layer0_outputs(5057));
    outputs(7386) <= (layer0_outputs(2475)) and not (layer0_outputs(3869));
    outputs(7387) <= not(layer0_outputs(6437));
    outputs(7388) <= layer0_outputs(8338);
    outputs(7389) <= (layer0_outputs(1607)) and (layer0_outputs(472));
    outputs(7390) <= (layer0_outputs(5466)) and not (layer0_outputs(5367));
    outputs(7391) <= not(layer0_outputs(9989));
    outputs(7392) <= not(layer0_outputs(193));
    outputs(7393) <= not((layer0_outputs(2586)) and (layer0_outputs(8109)));
    outputs(7394) <= not(layer0_outputs(6961));
    outputs(7395) <= not(layer0_outputs(4069)) or (layer0_outputs(3781));
    outputs(7396) <= (layer0_outputs(7832)) and (layer0_outputs(7533));
    outputs(7397) <= (layer0_outputs(8999)) and not (layer0_outputs(9470));
    outputs(7398) <= not(layer0_outputs(7936));
    outputs(7399) <= (layer0_outputs(7502)) and not (layer0_outputs(751));
    outputs(7400) <= (layer0_outputs(10040)) xor (layer0_outputs(1876));
    outputs(7401) <= not(layer0_outputs(63));
    outputs(7402) <= layer0_outputs(1663);
    outputs(7403) <= (layer0_outputs(2123)) or (layer0_outputs(8403));
    outputs(7404) <= layer0_outputs(6063);
    outputs(7405) <= layer0_outputs(4074);
    outputs(7406) <= (layer0_outputs(7100)) xor (layer0_outputs(5293));
    outputs(7407) <= not((layer0_outputs(9446)) and (layer0_outputs(9711)));
    outputs(7408) <= not(layer0_outputs(4158));
    outputs(7409) <= not((layer0_outputs(8485)) xor (layer0_outputs(1015)));
    outputs(7410) <= layer0_outputs(8471);
    outputs(7411) <= not(layer0_outputs(7345)) or (layer0_outputs(8840));
    outputs(7412) <= not(layer0_outputs(8994));
    outputs(7413) <= not(layer0_outputs(10019));
    outputs(7414) <= not(layer0_outputs(753));
    outputs(7415) <= not(layer0_outputs(255));
    outputs(7416) <= not((layer0_outputs(2605)) xor (layer0_outputs(8291)));
    outputs(7417) <= not(layer0_outputs(8400));
    outputs(7418) <= (layer0_outputs(5526)) and not (layer0_outputs(1919));
    outputs(7419) <= not(layer0_outputs(5013));
    outputs(7420) <= not((layer0_outputs(702)) xor (layer0_outputs(2932)));
    outputs(7421) <= (layer0_outputs(1485)) xor (layer0_outputs(10035));
    outputs(7422) <= (layer0_outputs(1383)) xor (layer0_outputs(3561));
    outputs(7423) <= not(layer0_outputs(3235));
    outputs(7424) <= not(layer0_outputs(193));
    outputs(7425) <= (layer0_outputs(2401)) and (layer0_outputs(4216));
    outputs(7426) <= not((layer0_outputs(1827)) or (layer0_outputs(9304)));
    outputs(7427) <= not(layer0_outputs(9658));
    outputs(7428) <= layer0_outputs(3476);
    outputs(7429) <= not(layer0_outputs(9959));
    outputs(7430) <= layer0_outputs(6516);
    outputs(7431) <= (layer0_outputs(742)) and not (layer0_outputs(2455));
    outputs(7432) <= not(layer0_outputs(2348));
    outputs(7433) <= not(layer0_outputs(2380)) or (layer0_outputs(8789));
    outputs(7434) <= layer0_outputs(4576);
    outputs(7435) <= not(layer0_outputs(4687));
    outputs(7436) <= layer0_outputs(6900);
    outputs(7437) <= not(layer0_outputs(575));
    outputs(7438) <= not(layer0_outputs(9842));
    outputs(7439) <= (layer0_outputs(5554)) and not (layer0_outputs(4127));
    outputs(7440) <= layer0_outputs(2359);
    outputs(7441) <= layer0_outputs(4742);
    outputs(7442) <= layer0_outputs(9032);
    outputs(7443) <= not(layer0_outputs(2259));
    outputs(7444) <= layer0_outputs(10225);
    outputs(7445) <= layer0_outputs(4149);
    outputs(7446) <= not(layer0_outputs(9050));
    outputs(7447) <= (layer0_outputs(1131)) xor (layer0_outputs(4277));
    outputs(7448) <= not((layer0_outputs(6076)) or (layer0_outputs(9962)));
    outputs(7449) <= not(layer0_outputs(6766));
    outputs(7450) <= (layer0_outputs(1184)) and (layer0_outputs(2071));
    outputs(7451) <= not(layer0_outputs(8280));
    outputs(7452) <= not(layer0_outputs(1075));
    outputs(7453) <= layer0_outputs(7179);
    outputs(7454) <= not(layer0_outputs(9291));
    outputs(7455) <= (layer0_outputs(61)) and (layer0_outputs(302));
    outputs(7456) <= (layer0_outputs(8763)) and (layer0_outputs(9892));
    outputs(7457) <= (layer0_outputs(3554)) and not (layer0_outputs(6043));
    outputs(7458) <= layer0_outputs(490);
    outputs(7459) <= (layer0_outputs(1018)) or (layer0_outputs(3176));
    outputs(7460) <= not(layer0_outputs(4121)) or (layer0_outputs(4395));
    outputs(7461) <= layer0_outputs(7987);
    outputs(7462) <= (layer0_outputs(3276)) and not (layer0_outputs(1127));
    outputs(7463) <= (layer0_outputs(5235)) xor (layer0_outputs(1440));
    outputs(7464) <= (layer0_outputs(4895)) and not (layer0_outputs(4991));
    outputs(7465) <= not(layer0_outputs(3114));
    outputs(7466) <= not((layer0_outputs(6189)) or (layer0_outputs(9105)));
    outputs(7467) <= layer0_outputs(8504);
    outputs(7468) <= not((layer0_outputs(1744)) xor (layer0_outputs(8904)));
    outputs(7469) <= (layer0_outputs(7678)) and (layer0_outputs(8182));
    outputs(7470) <= not(layer0_outputs(4412));
    outputs(7471) <= (layer0_outputs(9832)) and not (layer0_outputs(9419));
    outputs(7472) <= (layer0_outputs(4692)) and (layer0_outputs(5843));
    outputs(7473) <= (layer0_outputs(5567)) and not (layer0_outputs(1867));
    outputs(7474) <= not(layer0_outputs(2985));
    outputs(7475) <= layer0_outputs(7805);
    outputs(7476) <= not((layer0_outputs(6625)) or (layer0_outputs(7011)));
    outputs(7477) <= not((layer0_outputs(6858)) or (layer0_outputs(6411)));
    outputs(7478) <= (layer0_outputs(1167)) xor (layer0_outputs(1487));
    outputs(7479) <= (layer0_outputs(7850)) or (layer0_outputs(1501));
    outputs(7480) <= (layer0_outputs(4021)) or (layer0_outputs(2172));
    outputs(7481) <= (layer0_outputs(10110)) xor (layer0_outputs(4003));
    outputs(7482) <= layer0_outputs(7958);
    outputs(7483) <= (layer0_outputs(7649)) and (layer0_outputs(9846));
    outputs(7484) <= layer0_outputs(10210);
    outputs(7485) <= (layer0_outputs(4929)) and not (layer0_outputs(3465));
    outputs(7486) <= (layer0_outputs(4497)) xor (layer0_outputs(9283));
    outputs(7487) <= not(layer0_outputs(7948)) or (layer0_outputs(595));
    outputs(7488) <= (layer0_outputs(3624)) and not (layer0_outputs(4083));
    outputs(7489) <= layer0_outputs(2585);
    outputs(7490) <= layer0_outputs(8991);
    outputs(7491) <= not(layer0_outputs(6656));
    outputs(7492) <= not(layer0_outputs(8561));
    outputs(7493) <= (layer0_outputs(2166)) and not (layer0_outputs(7515));
    outputs(7494) <= not(layer0_outputs(3718));
    outputs(7495) <= not(layer0_outputs(3662));
    outputs(7496) <= not((layer0_outputs(8286)) and (layer0_outputs(8818)));
    outputs(7497) <= not(layer0_outputs(7998));
    outputs(7498) <= not(layer0_outputs(5189));
    outputs(7499) <= (layer0_outputs(7714)) xor (layer0_outputs(10184));
    outputs(7500) <= not(layer0_outputs(1495));
    outputs(7501) <= layer0_outputs(423);
    outputs(7502) <= not((layer0_outputs(6526)) xor (layer0_outputs(8598)));
    outputs(7503) <= (layer0_outputs(3601)) xor (layer0_outputs(7188));
    outputs(7504) <= (layer0_outputs(4166)) and not (layer0_outputs(819));
    outputs(7505) <= not(layer0_outputs(9632));
    outputs(7506) <= layer0_outputs(3138);
    outputs(7507) <= (layer0_outputs(9041)) and not (layer0_outputs(1636));
    outputs(7508) <= not(layer0_outputs(525));
    outputs(7509) <= layer0_outputs(783);
    outputs(7510) <= (layer0_outputs(9452)) and (layer0_outputs(5613));
    outputs(7511) <= (layer0_outputs(2610)) xor (layer0_outputs(7546));
    outputs(7512) <= layer0_outputs(1903);
    outputs(7513) <= (layer0_outputs(1951)) xor (layer0_outputs(7035));
    outputs(7514) <= (layer0_outputs(5265)) and (layer0_outputs(7995));
    outputs(7515) <= layer0_outputs(9601);
    outputs(7516) <= not(layer0_outputs(591));
    outputs(7517) <= not((layer0_outputs(4199)) xor (layer0_outputs(2249)));
    outputs(7518) <= not((layer0_outputs(2206)) or (layer0_outputs(1516)));
    outputs(7519) <= (layer0_outputs(5020)) or (layer0_outputs(9045));
    outputs(7520) <= not(layer0_outputs(4139));
    outputs(7521) <= layer0_outputs(3753);
    outputs(7522) <= layer0_outputs(7376);
    outputs(7523) <= (layer0_outputs(1546)) and not (layer0_outputs(194));
    outputs(7524) <= layer0_outputs(2149);
    outputs(7525) <= layer0_outputs(2855);
    outputs(7526) <= not((layer0_outputs(2344)) xor (layer0_outputs(24)));
    outputs(7527) <= (layer0_outputs(7416)) and not (layer0_outputs(4861));
    outputs(7528) <= not(layer0_outputs(963));
    outputs(7529) <= not((layer0_outputs(2358)) or (layer0_outputs(3595)));
    outputs(7530) <= layer0_outputs(8000);
    outputs(7531) <= (layer0_outputs(917)) and not (layer0_outputs(10113));
    outputs(7532) <= layer0_outputs(7855);
    outputs(7533) <= (layer0_outputs(5018)) and not (layer0_outputs(5401));
    outputs(7534) <= not(layer0_outputs(6654)) or (layer0_outputs(7359));
    outputs(7535) <= (layer0_outputs(3823)) and not (layer0_outputs(5179));
    outputs(7536) <= not(layer0_outputs(1556));
    outputs(7537) <= not((layer0_outputs(7732)) or (layer0_outputs(5024)));
    outputs(7538) <= not((layer0_outputs(2226)) or (layer0_outputs(1298)));
    outputs(7539) <= not(layer0_outputs(8229));
    outputs(7540) <= not((layer0_outputs(1153)) or (layer0_outputs(6004)));
    outputs(7541) <= not((layer0_outputs(3565)) xor (layer0_outputs(3640)));
    outputs(7542) <= layer0_outputs(4665);
    outputs(7543) <= (layer0_outputs(5626)) and not (layer0_outputs(10134));
    outputs(7544) <= not(layer0_outputs(1540));
    outputs(7545) <= (layer0_outputs(2180)) and not (layer0_outputs(603));
    outputs(7546) <= layer0_outputs(8039);
    outputs(7547) <= (layer0_outputs(8853)) and (layer0_outputs(6313));
    outputs(7548) <= (layer0_outputs(10104)) and (layer0_outputs(4152));
    outputs(7549) <= not((layer0_outputs(1335)) xor (layer0_outputs(9479)));
    outputs(7550) <= layer0_outputs(89);
    outputs(7551) <= (layer0_outputs(7410)) and (layer0_outputs(9608));
    outputs(7552) <= not(layer0_outputs(8823));
    outputs(7553) <= not(layer0_outputs(6733));
    outputs(7554) <= (layer0_outputs(264)) and not (layer0_outputs(9956));
    outputs(7555) <= layer0_outputs(4496);
    outputs(7556) <= not((layer0_outputs(2565)) xor (layer0_outputs(4326)));
    outputs(7557) <= (layer0_outputs(7414)) and not (layer0_outputs(2435));
    outputs(7558) <= (layer0_outputs(6153)) or (layer0_outputs(9294));
    outputs(7559) <= layer0_outputs(6866);
    outputs(7560) <= not(layer0_outputs(8684));
    outputs(7561) <= (layer0_outputs(1215)) and not (layer0_outputs(9671));
    outputs(7562) <= (layer0_outputs(5037)) and not (layer0_outputs(9252));
    outputs(7563) <= not(layer0_outputs(4670));
    outputs(7564) <= not(layer0_outputs(8252));
    outputs(7565) <= layer0_outputs(4677);
    outputs(7566) <= not(layer0_outputs(2538));
    outputs(7567) <= layer0_outputs(6878);
    outputs(7568) <= not(layer0_outputs(4989));
    outputs(7569) <= not((layer0_outputs(2922)) xor (layer0_outputs(2154)));
    outputs(7570) <= (layer0_outputs(7148)) and not (layer0_outputs(7058));
    outputs(7571) <= layer0_outputs(4954);
    outputs(7572) <= layer0_outputs(4196);
    outputs(7573) <= not(layer0_outputs(3155));
    outputs(7574) <= (layer0_outputs(789)) and (layer0_outputs(2397));
    outputs(7575) <= (layer0_outputs(4920)) xor (layer0_outputs(3203));
    outputs(7576) <= (layer0_outputs(8889)) and (layer0_outputs(7872));
    outputs(7577) <= (layer0_outputs(2149)) xor (layer0_outputs(4410));
    outputs(7578) <= layer0_outputs(5010);
    outputs(7579) <= not((layer0_outputs(9981)) xor (layer0_outputs(1904)));
    outputs(7580) <= layer0_outputs(5462);
    outputs(7581) <= layer0_outputs(1923);
    outputs(7582) <= layer0_outputs(8042);
    outputs(7583) <= (layer0_outputs(6466)) and not (layer0_outputs(9267));
    outputs(7584) <= (layer0_outputs(5834)) xor (layer0_outputs(7672));
    outputs(7585) <= not(layer0_outputs(2747));
    outputs(7586) <= not(layer0_outputs(8934));
    outputs(7587) <= (layer0_outputs(3672)) and (layer0_outputs(1309));
    outputs(7588) <= layer0_outputs(5193);
    outputs(7589) <= layer0_outputs(8731);
    outputs(7590) <= layer0_outputs(6053);
    outputs(7591) <= not(layer0_outputs(4967));
    outputs(7592) <= (layer0_outputs(8632)) xor (layer0_outputs(7916));
    outputs(7593) <= not(layer0_outputs(3477));
    outputs(7594) <= layer0_outputs(4793);
    outputs(7595) <= not(layer0_outputs(6758)) or (layer0_outputs(5341));
    outputs(7596) <= layer0_outputs(8619);
    outputs(7597) <= not((layer0_outputs(6559)) or (layer0_outputs(5343)));
    outputs(7598) <= layer0_outputs(3041);
    outputs(7599) <= not(layer0_outputs(5772));
    outputs(7600) <= not(layer0_outputs(7360));
    outputs(7601) <= layer0_outputs(2365);
    outputs(7602) <= (layer0_outputs(1668)) xor (layer0_outputs(7487));
    outputs(7603) <= not(layer0_outputs(6815));
    outputs(7604) <= not((layer0_outputs(7792)) or (layer0_outputs(5428)));
    outputs(7605) <= (layer0_outputs(6771)) xor (layer0_outputs(9300));
    outputs(7606) <= not(layer0_outputs(6047));
    outputs(7607) <= not(layer0_outputs(2967));
    outputs(7608) <= layer0_outputs(6475);
    outputs(7609) <= (layer0_outputs(9145)) and not (layer0_outputs(5430));
    outputs(7610) <= (layer0_outputs(5642)) and not (layer0_outputs(10008));
    outputs(7611) <= not(layer0_outputs(9466));
    outputs(7612) <= layer0_outputs(1118);
    outputs(7613) <= (layer0_outputs(3819)) and not (layer0_outputs(3972));
    outputs(7614) <= not(layer0_outputs(3818));
    outputs(7615) <= not(layer0_outputs(2491));
    outputs(7616) <= not(layer0_outputs(3942));
    outputs(7617) <= layer0_outputs(4485);
    outputs(7618) <= (layer0_outputs(4543)) xor (layer0_outputs(6964));
    outputs(7619) <= not(layer0_outputs(4774)) or (layer0_outputs(9825));
    outputs(7620) <= not((layer0_outputs(1740)) xor (layer0_outputs(9037)));
    outputs(7621) <= (layer0_outputs(4191)) and not (layer0_outputs(2974));
    outputs(7622) <= layer0_outputs(9384);
    outputs(7623) <= layer0_outputs(7477);
    outputs(7624) <= layer0_outputs(7729);
    outputs(7625) <= not(layer0_outputs(6963));
    outputs(7626) <= layer0_outputs(2365);
    outputs(7627) <= not(layer0_outputs(1437));
    outputs(7628) <= not(layer0_outputs(8088));
    outputs(7629) <= not(layer0_outputs(4716));
    outputs(7630) <= (layer0_outputs(5726)) and (layer0_outputs(9023));
    outputs(7631) <= (layer0_outputs(6913)) and not (layer0_outputs(6233));
    outputs(7632) <= not(layer0_outputs(7403));
    outputs(7633) <= (layer0_outputs(4601)) and (layer0_outputs(5922));
    outputs(7634) <= (layer0_outputs(4404)) and not (layer0_outputs(40));
    outputs(7635) <= layer0_outputs(5399);
    outputs(7636) <= (layer0_outputs(4484)) and not (layer0_outputs(704));
    outputs(7637) <= layer0_outputs(7460);
    outputs(7638) <= (layer0_outputs(3702)) and (layer0_outputs(8540));
    outputs(7639) <= not(layer0_outputs(8643)) or (layer0_outputs(608));
    outputs(7640) <= (layer0_outputs(3556)) xor (layer0_outputs(10032));
    outputs(7641) <= not(layer0_outputs(4841));
    outputs(7642) <= not((layer0_outputs(5032)) xor (layer0_outputs(7119)));
    outputs(7643) <= (layer0_outputs(3944)) and not (layer0_outputs(1329));
    outputs(7644) <= (layer0_outputs(8762)) and not (layer0_outputs(2860));
    outputs(7645) <= (layer0_outputs(8048)) and not (layer0_outputs(9833));
    outputs(7646) <= not(layer0_outputs(10194));
    outputs(7647) <= (layer0_outputs(2004)) and (layer0_outputs(1728));
    outputs(7648) <= layer0_outputs(9324);
    outputs(7649) <= not(layer0_outputs(5294));
    outputs(7650) <= not(layer0_outputs(9974));
    outputs(7651) <= layer0_outputs(537);
    outputs(7652) <= layer0_outputs(3968);
    outputs(7653) <= (layer0_outputs(2646)) and not (layer0_outputs(6897));
    outputs(7654) <= (layer0_outputs(4527)) and (layer0_outputs(10014));
    outputs(7655) <= (layer0_outputs(1378)) xor (layer0_outputs(8428));
    outputs(7656) <= not(layer0_outputs(3823));
    outputs(7657) <= (layer0_outputs(2184)) and (layer0_outputs(6751));
    outputs(7658) <= (layer0_outputs(7874)) and not (layer0_outputs(7176));
    outputs(7659) <= layer0_outputs(7681);
    outputs(7660) <= not((layer0_outputs(2825)) xor (layer0_outputs(6712)));
    outputs(7661) <= not(layer0_outputs(8716));
    outputs(7662) <= (layer0_outputs(4415)) and not (layer0_outputs(1071));
    outputs(7663) <= layer0_outputs(2472);
    outputs(7664) <= not(layer0_outputs(7956));
    outputs(7665) <= layer0_outputs(4038);
    outputs(7666) <= not((layer0_outputs(7836)) xor (layer0_outputs(5361)));
    outputs(7667) <= (layer0_outputs(733)) and not (layer0_outputs(8997));
    outputs(7668) <= not((layer0_outputs(5963)) xor (layer0_outputs(4834)));
    outputs(7669) <= layer0_outputs(5957);
    outputs(7670) <= (layer0_outputs(2050)) and (layer0_outputs(4009));
    outputs(7671) <= not((layer0_outputs(6806)) or (layer0_outputs(6690)));
    outputs(7672) <= (layer0_outputs(3193)) and not (layer0_outputs(1951));
    outputs(7673) <= (layer0_outputs(8271)) xor (layer0_outputs(3189));
    outputs(7674) <= (layer0_outputs(7796)) xor (layer0_outputs(7810));
    outputs(7675) <= not((layer0_outputs(6971)) or (layer0_outputs(8849)));
    outputs(7676) <= (layer0_outputs(9272)) xor (layer0_outputs(1206));
    outputs(7677) <= layer0_outputs(7009);
    outputs(7678) <= layer0_outputs(7852);
    outputs(7679) <= (layer0_outputs(854)) xor (layer0_outputs(7455));
    outputs(7680) <= not(layer0_outputs(9502));
    outputs(7681) <= (layer0_outputs(2445)) and not (layer0_outputs(7206));
    outputs(7682) <= layer0_outputs(9984);
    outputs(7683) <= (layer0_outputs(1056)) and (layer0_outputs(3819));
    outputs(7684) <= not((layer0_outputs(4689)) or (layer0_outputs(962)));
    outputs(7685) <= (layer0_outputs(4583)) and not (layer0_outputs(6735));
    outputs(7686) <= not(layer0_outputs(2886)) or (layer0_outputs(8956));
    outputs(7687) <= layer0_outputs(6038);
    outputs(7688) <= layer0_outputs(8509);
    outputs(7689) <= not(layer0_outputs(6383));
    outputs(7690) <= not(layer0_outputs(8014));
    outputs(7691) <= not(layer0_outputs(8470));
    outputs(7692) <= layer0_outputs(3170);
    outputs(7693) <= layer0_outputs(4724);
    outputs(7694) <= (layer0_outputs(5295)) xor (layer0_outputs(8416));
    outputs(7695) <= not(layer0_outputs(9890));
    outputs(7696) <= not(layer0_outputs(3551));
    outputs(7697) <= not(layer0_outputs(8266));
    outputs(7698) <= layer0_outputs(1847);
    outputs(7699) <= layer0_outputs(9827);
    outputs(7700) <= not(layer0_outputs(5403));
    outputs(7701) <= not((layer0_outputs(4597)) or (layer0_outputs(6335)));
    outputs(7702) <= not(layer0_outputs(2710));
    outputs(7703) <= (layer0_outputs(6120)) and not (layer0_outputs(2924));
    outputs(7704) <= layer0_outputs(9297);
    outputs(7705) <= not(layer0_outputs(4169));
    outputs(7706) <= (layer0_outputs(3193)) and not (layer0_outputs(2773));
    outputs(7707) <= not(layer0_outputs(953));
    outputs(7708) <= layer0_outputs(7683);
    outputs(7709) <= not(layer0_outputs(6679));
    outputs(7710) <= (layer0_outputs(4835)) and not (layer0_outputs(4917));
    outputs(7711) <= (layer0_outputs(6214)) xor (layer0_outputs(3889));
    outputs(7712) <= not(layer0_outputs(10143));
    outputs(7713) <= layer0_outputs(3545);
    outputs(7714) <= layer0_outputs(6615);
    outputs(7715) <= layer0_outputs(6266);
    outputs(7716) <= not((layer0_outputs(2890)) or (layer0_outputs(6864)));
    outputs(7717) <= not(layer0_outputs(5684));
    outputs(7718) <= not(layer0_outputs(2208));
    outputs(7719) <= not(layer0_outputs(9449));
    outputs(7720) <= layer0_outputs(497);
    outputs(7721) <= (layer0_outputs(3261)) and not (layer0_outputs(4580));
    outputs(7722) <= layer0_outputs(10235);
    outputs(7723) <= (layer0_outputs(5928)) and not (layer0_outputs(7139));
    outputs(7724) <= not((layer0_outputs(7429)) or (layer0_outputs(2155)));
    outputs(7725) <= layer0_outputs(9276);
    outputs(7726) <= layer0_outputs(7531);
    outputs(7727) <= not(layer0_outputs(1158));
    outputs(7728) <= not((layer0_outputs(8121)) or (layer0_outputs(2828)));
    outputs(7729) <= not((layer0_outputs(1992)) xor (layer0_outputs(2862)));
    outputs(7730) <= not(layer0_outputs(8140));
    outputs(7731) <= layer0_outputs(5345);
    outputs(7732) <= not(layer0_outputs(8720));
    outputs(7733) <= not(layer0_outputs(2001));
    outputs(7734) <= (layer0_outputs(1979)) and (layer0_outputs(9858));
    outputs(7735) <= layer0_outputs(5872);
    outputs(7736) <= (layer0_outputs(3808)) xor (layer0_outputs(7621));
    outputs(7737) <= not((layer0_outputs(4341)) xor (layer0_outputs(5007)));
    outputs(7738) <= layer0_outputs(6968);
    outputs(7739) <= (layer0_outputs(9613)) and not (layer0_outputs(1403));
    outputs(7740) <= (layer0_outputs(6977)) and not (layer0_outputs(8979));
    outputs(7741) <= (layer0_outputs(4383)) xor (layer0_outputs(5930));
    outputs(7742) <= not(layer0_outputs(4223));
    outputs(7743) <= (layer0_outputs(470)) or (layer0_outputs(371));
    outputs(7744) <= not(layer0_outputs(8120));
    outputs(7745) <= (layer0_outputs(3535)) or (layer0_outputs(2419));
    outputs(7746) <= layer0_outputs(8785);
    outputs(7747) <= (layer0_outputs(999)) and not (layer0_outputs(6704));
    outputs(7748) <= layer0_outputs(5673);
    outputs(7749) <= (layer0_outputs(7202)) xor (layer0_outputs(1204));
    outputs(7750) <= (layer0_outputs(7765)) and not (layer0_outputs(8322));
    outputs(7751) <= (layer0_outputs(3878)) and (layer0_outputs(8383));
    outputs(7752) <= not((layer0_outputs(8207)) or (layer0_outputs(7092)));
    outputs(7753) <= (layer0_outputs(9030)) xor (layer0_outputs(972));
    outputs(7754) <= (layer0_outputs(8180)) and not (layer0_outputs(6681));
    outputs(7755) <= not((layer0_outputs(5667)) or (layer0_outputs(10037)));
    outputs(7756) <= layer0_outputs(10125);
    outputs(7757) <= layer0_outputs(667);
    outputs(7758) <= layer0_outputs(2507);
    outputs(7759) <= not((layer0_outputs(1365)) and (layer0_outputs(7875)));
    outputs(7760) <= not(layer0_outputs(5041));
    outputs(7761) <= layer0_outputs(2941);
    outputs(7762) <= not((layer0_outputs(4610)) or (layer0_outputs(2506)));
    outputs(7763) <= layer0_outputs(88);
    outputs(7764) <= not((layer0_outputs(7711)) xor (layer0_outputs(5577)));
    outputs(7765) <= not(layer0_outputs(132));
    outputs(7766) <= (layer0_outputs(6201)) or (layer0_outputs(7718));
    outputs(7767) <= (layer0_outputs(530)) xor (layer0_outputs(839));
    outputs(7768) <= not((layer0_outputs(9739)) xor (layer0_outputs(8859)));
    outputs(7769) <= layer0_outputs(10152);
    outputs(7770) <= layer0_outputs(9670);
    outputs(7771) <= layer0_outputs(8852);
    outputs(7772) <= not(layer0_outputs(1072));
    outputs(7773) <= not((layer0_outputs(3338)) xor (layer0_outputs(8638)));
    outputs(7774) <= not(layer0_outputs(104));
    outputs(7775) <= not(layer0_outputs(290)) or (layer0_outputs(3289));
    outputs(7776) <= layer0_outputs(9290);
    outputs(7777) <= not(layer0_outputs(5350));
    outputs(7778) <= layer0_outputs(788);
    outputs(7779) <= (layer0_outputs(3436)) and not (layer0_outputs(8423));
    outputs(7780) <= (layer0_outputs(4918)) xor (layer0_outputs(2617));
    outputs(7781) <= (layer0_outputs(1249)) xor (layer0_outputs(6212));
    outputs(7782) <= (layer0_outputs(6374)) and not (layer0_outputs(8877));
    outputs(7783) <= (layer0_outputs(4641)) and not (layer0_outputs(6673));
    outputs(7784) <= (layer0_outputs(3248)) xor (layer0_outputs(5416));
    outputs(7785) <= not((layer0_outputs(9430)) xor (layer0_outputs(7701)));
    outputs(7786) <= not(layer0_outputs(1784));
    outputs(7787) <= layer0_outputs(5355);
    outputs(7788) <= not(layer0_outputs(79));
    outputs(7789) <= not((layer0_outputs(4094)) or (layer0_outputs(1484)));
    outputs(7790) <= (layer0_outputs(1721)) and not (layer0_outputs(6139));
    outputs(7791) <= (layer0_outputs(1321)) and not (layer0_outputs(8472));
    outputs(7792) <= not((layer0_outputs(3218)) or (layer0_outputs(1950)));
    outputs(7793) <= not(layer0_outputs(2992));
    outputs(7794) <= (layer0_outputs(291)) xor (layer0_outputs(5934));
    outputs(7795) <= (layer0_outputs(6608)) and not (layer0_outputs(3881));
    outputs(7796) <= not(layer0_outputs(3020)) or (layer0_outputs(7965));
    outputs(7797) <= not(layer0_outputs(9958));
    outputs(7798) <= (layer0_outputs(7226)) xor (layer0_outputs(7696));
    outputs(7799) <= (layer0_outputs(7795)) xor (layer0_outputs(7256));
    outputs(7800) <= not((layer0_outputs(4893)) or (layer0_outputs(797)));
    outputs(7801) <= not(layer0_outputs(7839));
    outputs(7802) <= layer0_outputs(5949);
    outputs(7803) <= not(layer0_outputs(6157));
    outputs(7804) <= not(layer0_outputs(9287));
    outputs(7805) <= not((layer0_outputs(2937)) or (layer0_outputs(9469)));
    outputs(7806) <= not((layer0_outputs(7959)) xor (layer0_outputs(8815)));
    outputs(7807) <= not(layer0_outputs(3263));
    outputs(7808) <= not((layer0_outputs(6243)) xor (layer0_outputs(7351)));
    outputs(7809) <= not((layer0_outputs(9811)) xor (layer0_outputs(1341)));
    outputs(7810) <= layer0_outputs(1098);
    outputs(7811) <= layer0_outputs(2268);
    outputs(7812) <= not(layer0_outputs(3629));
    outputs(7813) <= layer0_outputs(4868);
    outputs(7814) <= layer0_outputs(8620);
    outputs(7815) <= not(layer0_outputs(8813));
    outputs(7816) <= (layer0_outputs(9983)) and not (layer0_outputs(8040));
    outputs(7817) <= not((layer0_outputs(1468)) xor (layer0_outputs(8814)));
    outputs(7818) <= not(layer0_outputs(183));
    outputs(7819) <= (layer0_outputs(4289)) and not (layer0_outputs(9751));
    outputs(7820) <= layer0_outputs(9271);
    outputs(7821) <= (layer0_outputs(9778)) and not (layer0_outputs(5286));
    outputs(7822) <= layer0_outputs(5708);
    outputs(7823) <= layer0_outputs(4581);
    outputs(7824) <= not(layer0_outputs(7960));
    outputs(7825) <= not(layer0_outputs(7432));
    outputs(7826) <= layer0_outputs(4879);
    outputs(7827) <= (layer0_outputs(8157)) and not (layer0_outputs(6646));
    outputs(7828) <= not((layer0_outputs(3905)) xor (layer0_outputs(4159)));
    outputs(7829) <= (layer0_outputs(2293)) and not (layer0_outputs(4374));
    outputs(7830) <= (layer0_outputs(2930)) and not (layer0_outputs(3582));
    outputs(7831) <= layer0_outputs(3450);
    outputs(7832) <= layer0_outputs(5278);
    outputs(7833) <= not(layer0_outputs(6400)) or (layer0_outputs(4389));
    outputs(7834) <= layer0_outputs(9086);
    outputs(7835) <= layer0_outputs(137);
    outputs(7836) <= (layer0_outputs(6217)) and not (layer0_outputs(4220));
    outputs(7837) <= (layer0_outputs(6928)) and (layer0_outputs(7268));
    outputs(7838) <= layer0_outputs(3804);
    outputs(7839) <= (layer0_outputs(144)) and not (layer0_outputs(8672));
    outputs(7840) <= not((layer0_outputs(7118)) xor (layer0_outputs(2669)));
    outputs(7841) <= layer0_outputs(1677);
    outputs(7842) <= not(layer0_outputs(6288));
    outputs(7843) <= layer0_outputs(10152);
    outputs(7844) <= not(layer0_outputs(7868));
    outputs(7845) <= not((layer0_outputs(8880)) or (layer0_outputs(4981)));
    outputs(7846) <= not(layer0_outputs(1835));
    outputs(7847) <= (layer0_outputs(8654)) or (layer0_outputs(3759));
    outputs(7848) <= (layer0_outputs(7806)) and (layer0_outputs(5691));
    outputs(7849) <= (layer0_outputs(9678)) and not (layer0_outputs(8554));
    outputs(7850) <= (layer0_outputs(9624)) and (layer0_outputs(196));
    outputs(7851) <= (layer0_outputs(7840)) and not (layer0_outputs(10036));
    outputs(7852) <= not(layer0_outputs(6137));
    outputs(7853) <= not(layer0_outputs(7848));
    outputs(7854) <= not(layer0_outputs(6569)) or (layer0_outputs(4418));
    outputs(7855) <= not((layer0_outputs(1806)) xor (layer0_outputs(7730)));
    outputs(7856) <= layer0_outputs(7357);
    outputs(7857) <= layer0_outputs(7807);
    outputs(7858) <= layer0_outputs(2596);
    outputs(7859) <= layer0_outputs(3758);
    outputs(7860) <= not(layer0_outputs(5809));
    outputs(7861) <= not(layer0_outputs(8871));
    outputs(7862) <= layer0_outputs(3119);
    outputs(7863) <= not(layer0_outputs(6597));
    outputs(7864) <= not((layer0_outputs(5868)) xor (layer0_outputs(4299)));
    outputs(7865) <= (layer0_outputs(3465)) and not (layer0_outputs(603));
    outputs(7866) <= not(layer0_outputs(1787));
    outputs(7867) <= not(layer0_outputs(6428));
    outputs(7868) <= (layer0_outputs(5124)) and (layer0_outputs(922));
    outputs(7869) <= layer0_outputs(6771);
    outputs(7870) <= (layer0_outputs(9757)) xor (layer0_outputs(5539));
    outputs(7871) <= not((layer0_outputs(9782)) or (layer0_outputs(3239)));
    outputs(7872) <= (layer0_outputs(2280)) and not (layer0_outputs(5982));
    outputs(7873) <= layer0_outputs(394);
    outputs(7874) <= not(layer0_outputs(7849));
    outputs(7875) <= (layer0_outputs(1188)) xor (layer0_outputs(7530));
    outputs(7876) <= not(layer0_outputs(5657)) or (layer0_outputs(7587));
    outputs(7877) <= not(layer0_outputs(1327));
    outputs(7878) <= layer0_outputs(5251);
    outputs(7879) <= not(layer0_outputs(1846)) or (layer0_outputs(8149));
    outputs(7880) <= (layer0_outputs(1788)) and not (layer0_outputs(6395));
    outputs(7881) <= (layer0_outputs(8283)) and not (layer0_outputs(2142));
    outputs(7882) <= not(layer0_outputs(7642));
    outputs(7883) <= not((layer0_outputs(8969)) or (layer0_outputs(3833)));
    outputs(7884) <= layer0_outputs(9870);
    outputs(7885) <= layer0_outputs(9701);
    outputs(7886) <= not(layer0_outputs(6684));
    outputs(7887) <= layer0_outputs(7081);
    outputs(7888) <= layer0_outputs(1626);
    outputs(7889) <= layer0_outputs(3770);
    outputs(7890) <= layer0_outputs(9580);
    outputs(7891) <= (layer0_outputs(6972)) and (layer0_outputs(7893));
    outputs(7892) <= not(layer0_outputs(3742));
    outputs(7893) <= not((layer0_outputs(4855)) xor (layer0_outputs(8235)));
    outputs(7894) <= not(layer0_outputs(1324));
    outputs(7895) <= not((layer0_outputs(4854)) xor (layer0_outputs(6091)));
    outputs(7896) <= (layer0_outputs(5257)) and not (layer0_outputs(8193));
    outputs(7897) <= layer0_outputs(2464);
    outputs(7898) <= not(layer0_outputs(6562));
    outputs(7899) <= not(layer0_outputs(1276));
    outputs(7900) <= not(layer0_outputs(4499));
    outputs(7901) <= (layer0_outputs(9756)) and not (layer0_outputs(2229));
    outputs(7902) <= not((layer0_outputs(2083)) xor (layer0_outputs(2144)));
    outputs(7903) <= layer0_outputs(8230);
    outputs(7904) <= not(layer0_outputs(243));
    outputs(7905) <= not(layer0_outputs(6888));
    outputs(7906) <= (layer0_outputs(9210)) xor (layer0_outputs(2662));
    outputs(7907) <= (layer0_outputs(4573)) xor (layer0_outputs(10187));
    outputs(7908) <= (layer0_outputs(8961)) xor (layer0_outputs(4850));
    outputs(7909) <= layer0_outputs(9192);
    outputs(7910) <= (layer0_outputs(8081)) and not (layer0_outputs(3740));
    outputs(7911) <= not(layer0_outputs(234));
    outputs(7912) <= not(layer0_outputs(1375));
    outputs(7913) <= not(layer0_outputs(6992));
    outputs(7914) <= layer0_outputs(1587);
    outputs(7915) <= not(layer0_outputs(889));
    outputs(7916) <= (layer0_outputs(2861)) and not (layer0_outputs(7781));
    outputs(7917) <= (layer0_outputs(701)) and not (layer0_outputs(10027));
    outputs(7918) <= (layer0_outputs(9631)) and (layer0_outputs(9812));
    outputs(7919) <= layer0_outputs(1525);
    outputs(7920) <= not((layer0_outputs(8565)) or (layer0_outputs(8430)));
    outputs(7921) <= not(layer0_outputs(867));
    outputs(7922) <= (layer0_outputs(6098)) and not (layer0_outputs(7547));
    outputs(7923) <= not((layer0_outputs(6520)) xor (layer0_outputs(3624)));
    outputs(7924) <= not(layer0_outputs(8607));
    outputs(7925) <= (layer0_outputs(3153)) xor (layer0_outputs(1128));
    outputs(7926) <= (layer0_outputs(6799)) and not (layer0_outputs(6734));
    outputs(7927) <= not(layer0_outputs(6108)) or (layer0_outputs(3585));
    outputs(7928) <= not((layer0_outputs(8364)) xor (layer0_outputs(6244)));
    outputs(7929) <= layer0_outputs(3827);
    outputs(7930) <= layer0_outputs(8412);
    outputs(7931) <= not(layer0_outputs(6672)) or (layer0_outputs(1993));
    outputs(7932) <= not(layer0_outputs(1406));
    outputs(7933) <= (layer0_outputs(3871)) xor (layer0_outputs(3380));
    outputs(7934) <= layer0_outputs(3574);
    outputs(7935) <= (layer0_outputs(9217)) and (layer0_outputs(13));
    outputs(7936) <= layer0_outputs(5977);
    outputs(7937) <= layer0_outputs(640);
    outputs(7938) <= not((layer0_outputs(8705)) or (layer0_outputs(4013)));
    outputs(7939) <= layer0_outputs(9333);
    outputs(7940) <= not(layer0_outputs(3047));
    outputs(7941) <= layer0_outputs(9979);
    outputs(7942) <= layer0_outputs(4290);
    outputs(7943) <= not(layer0_outputs(6758));
    outputs(7944) <= not(layer0_outputs(5659));
    outputs(7945) <= not((layer0_outputs(1844)) xor (layer0_outputs(5865)));
    outputs(7946) <= not(layer0_outputs(7191));
    outputs(7947) <= layer0_outputs(2345);
    outputs(7948) <= (layer0_outputs(8786)) and not (layer0_outputs(1131));
    outputs(7949) <= layer0_outputs(6460);
    outputs(7950) <= not(layer0_outputs(3562));
    outputs(7951) <= layer0_outputs(3826);
    outputs(7952) <= (layer0_outputs(89)) and (layer0_outputs(7234));
    outputs(7953) <= not(layer0_outputs(8488)) or (layer0_outputs(6297));
    outputs(7954) <= not((layer0_outputs(2632)) or (layer0_outputs(5948)));
    outputs(7955) <= layer0_outputs(8597);
    outputs(7956) <= layer0_outputs(9953);
    outputs(7957) <= not((layer0_outputs(3993)) xor (layer0_outputs(7755)));
    outputs(7958) <= layer0_outputs(2305);
    outputs(7959) <= not(layer0_outputs(865));
    outputs(7960) <= (layer0_outputs(5386)) xor (layer0_outputs(9356));
    outputs(7961) <= (layer0_outputs(5563)) and not (layer0_outputs(9742));
    outputs(7962) <= (layer0_outputs(4422)) and not (layer0_outputs(4477));
    outputs(7963) <= (layer0_outputs(5014)) xor (layer0_outputs(1254));
    outputs(7964) <= (layer0_outputs(4828)) and (layer0_outputs(5629));
    outputs(7965) <= not(layer0_outputs(3286));
    outputs(7966) <= not(layer0_outputs(6305));
    outputs(7967) <= (layer0_outputs(7591)) xor (layer0_outputs(5874));
    outputs(7968) <= not(layer0_outputs(4510));
    outputs(7969) <= layer0_outputs(7895);
    outputs(7970) <= not((layer0_outputs(7464)) or (layer0_outputs(7172)));
    outputs(7971) <= (layer0_outputs(6062)) and (layer0_outputs(7380));
    outputs(7972) <= (layer0_outputs(8703)) xor (layer0_outputs(1259));
    outputs(7973) <= not(layer0_outputs(9317));
    outputs(7974) <= (layer0_outputs(7238)) and not (layer0_outputs(1837));
    outputs(7975) <= not((layer0_outputs(7871)) xor (layer0_outputs(5224)));
    outputs(7976) <= (layer0_outputs(8288)) or (layer0_outputs(8819));
    outputs(7977) <= not(layer0_outputs(2934));
    outputs(7978) <= layer0_outputs(7320);
    outputs(7979) <= layer0_outputs(8555);
    outputs(7980) <= (layer0_outputs(2936)) and not (layer0_outputs(172));
    outputs(7981) <= not((layer0_outputs(9570)) or (layer0_outputs(4344)));
    outputs(7982) <= not(layer0_outputs(3047));
    outputs(7983) <= layer0_outputs(5680);
    outputs(7984) <= layer0_outputs(1263);
    outputs(7985) <= (layer0_outputs(8096)) xor (layer0_outputs(6785));
    outputs(7986) <= not(layer0_outputs(5879)) or (layer0_outputs(8111));
    outputs(7987) <= not(layer0_outputs(2802));
    outputs(7988) <= not(layer0_outputs(5276));
    outputs(7989) <= layer0_outputs(5722);
    outputs(7990) <= not((layer0_outputs(4085)) or (layer0_outputs(3058)));
    outputs(7991) <= (layer0_outputs(1469)) xor (layer0_outputs(4875));
    outputs(7992) <= not(layer0_outputs(122));
    outputs(7993) <= layer0_outputs(1032);
    outputs(7994) <= not(layer0_outputs(2766));
    outputs(7995) <= not(layer0_outputs(3224));
    outputs(7996) <= layer0_outputs(8475);
    outputs(7997) <= (layer0_outputs(2630)) xor (layer0_outputs(9388));
    outputs(7998) <= not((layer0_outputs(6123)) xor (layer0_outputs(7099)));
    outputs(7999) <= layer0_outputs(6900);
    outputs(8000) <= layer0_outputs(4078);
    outputs(8001) <= layer0_outputs(1747);
    outputs(8002) <= not(layer0_outputs(3447));
    outputs(8003) <= not(layer0_outputs(3250));
    outputs(8004) <= not((layer0_outputs(9806)) or (layer0_outputs(2432)));
    outputs(8005) <= not((layer0_outputs(5064)) or (layer0_outputs(3714)));
    outputs(8006) <= not(layer0_outputs(5857)) or (layer0_outputs(6896));
    outputs(8007) <= not(layer0_outputs(1730));
    outputs(8008) <= not((layer0_outputs(1000)) and (layer0_outputs(2826)));
    outputs(8009) <= not(layer0_outputs(7622));
    outputs(8010) <= layer0_outputs(1207);
    outputs(8011) <= not(layer0_outputs(2301));
    outputs(8012) <= layer0_outputs(4605);
    outputs(8013) <= layer0_outputs(3267);
    outputs(8014) <= not(layer0_outputs(6178));
    outputs(8015) <= layer0_outputs(4708);
    outputs(8016) <= not((layer0_outputs(3629)) or (layer0_outputs(2390)));
    outputs(8017) <= layer0_outputs(10118);
    outputs(8018) <= (layer0_outputs(6864)) xor (layer0_outputs(3422));
    outputs(8019) <= (layer0_outputs(3895)) and not (layer0_outputs(422));
    outputs(8020) <= (layer0_outputs(9847)) and not (layer0_outputs(7834));
    outputs(8021) <= (layer0_outputs(7315)) and (layer0_outputs(7992));
    outputs(8022) <= (layer0_outputs(8111)) and not (layer0_outputs(6787));
    outputs(8023) <= not((layer0_outputs(2760)) xor (layer0_outputs(2646)));
    outputs(8024) <= not((layer0_outputs(4302)) or (layer0_outputs(3862)));
    outputs(8025) <= not(layer0_outputs(9845));
    outputs(8026) <= layer0_outputs(434);
    outputs(8027) <= (layer0_outputs(158)) xor (layer0_outputs(8034));
    outputs(8028) <= not(layer0_outputs(10105));
    outputs(8029) <= not(layer0_outputs(6495));
    outputs(8030) <= (layer0_outputs(8127)) and not (layer0_outputs(7967));
    outputs(8031) <= not(layer0_outputs(3106));
    outputs(8032) <= (layer0_outputs(9118)) xor (layer0_outputs(6584));
    outputs(8033) <= layer0_outputs(5748);
    outputs(8034) <= (layer0_outputs(7888)) and not (layer0_outputs(3239));
    outputs(8035) <= (layer0_outputs(8314)) and (layer0_outputs(7821));
    outputs(8036) <= layer0_outputs(1501);
    outputs(8037) <= (layer0_outputs(1662)) and (layer0_outputs(6774));
    outputs(8038) <= not((layer0_outputs(1068)) xor (layer0_outputs(6716)));
    outputs(8039) <= (layer0_outputs(5116)) and not (layer0_outputs(6743));
    outputs(8040) <= layer0_outputs(6163);
    outputs(8041) <= (layer0_outputs(8408)) xor (layer0_outputs(5365));
    outputs(8042) <= layer0_outputs(2839);
    outputs(8043) <= not((layer0_outputs(3079)) or (layer0_outputs(7065)));
    outputs(8044) <= not(layer0_outputs(8240)) or (layer0_outputs(8365));
    outputs(8045) <= layer0_outputs(10056);
    outputs(8046) <= layer0_outputs(5768);
    outputs(8047) <= (layer0_outputs(8868)) and not (layer0_outputs(3797));
    outputs(8048) <= not(layer0_outputs(4820));
    outputs(8049) <= layer0_outputs(9980);
    outputs(8050) <= not(layer0_outputs(4860));
    outputs(8051) <= not(layer0_outputs(5280));
    outputs(8052) <= layer0_outputs(3613);
    outputs(8053) <= layer0_outputs(8443);
    outputs(8054) <= not(layer0_outputs(7158));
    outputs(8055) <= (layer0_outputs(3398)) and not (layer0_outputs(9358));
    outputs(8056) <= not((layer0_outputs(7329)) xor (layer0_outputs(1849)));
    outputs(8057) <= (layer0_outputs(5613)) and (layer0_outputs(6832));
    outputs(8058) <= layer0_outputs(2767);
    outputs(8059) <= not((layer0_outputs(3157)) xor (layer0_outputs(7700)));
    outputs(8060) <= layer0_outputs(5901);
    outputs(8061) <= layer0_outputs(8700);
    outputs(8062) <= not((layer0_outputs(1497)) or (layer0_outputs(1597)));
    outputs(8063) <= layer0_outputs(7219);
    outputs(8064) <= not(layer0_outputs(5137));
    outputs(8065) <= not(layer0_outputs(980));
    outputs(8066) <= not(layer0_outputs(8019));
    outputs(8067) <= not(layer0_outputs(9000));
    outputs(8068) <= not(layer0_outputs(7077)) or (layer0_outputs(9337));
    outputs(8069) <= not(layer0_outputs(8110));
    outputs(8070) <= (layer0_outputs(8753)) and (layer0_outputs(28));
    outputs(8071) <= (layer0_outputs(1428)) xor (layer0_outputs(5168));
    outputs(8072) <= (layer0_outputs(6326)) and not (layer0_outputs(4836));
    outputs(8073) <= not(layer0_outputs(1467));
    outputs(8074) <= not((layer0_outputs(9094)) and (layer0_outputs(1852)));
    outputs(8075) <= not((layer0_outputs(6360)) and (layer0_outputs(3743)));
    outputs(8076) <= not((layer0_outputs(3937)) xor (layer0_outputs(1843)));
    outputs(8077) <= not((layer0_outputs(802)) and (layer0_outputs(4411)));
    outputs(8078) <= layer0_outputs(2427);
    outputs(8079) <= layer0_outputs(6462);
    outputs(8080) <= (layer0_outputs(9709)) xor (layer0_outputs(7432));
    outputs(8081) <= not((layer0_outputs(4816)) and (layer0_outputs(2600)));
    outputs(8082) <= (layer0_outputs(537)) and not (layer0_outputs(4814));
    outputs(8083) <= not(layer0_outputs(6202));
    outputs(8084) <= not(layer0_outputs(4135));
    outputs(8085) <= not((layer0_outputs(2214)) xor (layer0_outputs(6532)));
    outputs(8086) <= (layer0_outputs(2028)) xor (layer0_outputs(777));
    outputs(8087) <= not((layer0_outputs(5919)) or (layer0_outputs(1075)));
    outputs(8088) <= not(layer0_outputs(5501)) or (layer0_outputs(2534));
    outputs(8089) <= layer0_outputs(4867);
    outputs(8090) <= not(layer0_outputs(9154));
    outputs(8091) <= not(layer0_outputs(1569));
    outputs(8092) <= (layer0_outputs(4752)) and not (layer0_outputs(2218));
    outputs(8093) <= (layer0_outputs(9571)) xor (layer0_outputs(8489));
    outputs(8094) <= (layer0_outputs(5596)) xor (layer0_outputs(9537));
    outputs(8095) <= not(layer0_outputs(679));
    outputs(8096) <= not((layer0_outputs(9064)) or (layer0_outputs(4363)));
    outputs(8097) <= layer0_outputs(6489);
    outputs(8098) <= layer0_outputs(8136);
    outputs(8099) <= not(layer0_outputs(311));
    outputs(8100) <= not((layer0_outputs(5898)) xor (layer0_outputs(1889)));
    outputs(8101) <= (layer0_outputs(5590)) and (layer0_outputs(5984));
    outputs(8102) <= layer0_outputs(9868);
    outputs(8103) <= layer0_outputs(707);
    outputs(8104) <= layer0_outputs(9233);
    outputs(8105) <= not((layer0_outputs(7399)) xor (layer0_outputs(6608)));
    outputs(8106) <= (layer0_outputs(9036)) xor (layer0_outputs(4848));
    outputs(8107) <= (layer0_outputs(6931)) and (layer0_outputs(2611));
    outputs(8108) <= (layer0_outputs(7306)) and not (layer0_outputs(9155));
    outputs(8109) <= (layer0_outputs(6926)) and not (layer0_outputs(3891));
    outputs(8110) <= layer0_outputs(1145);
    outputs(8111) <= not(layer0_outputs(2150));
    outputs(8112) <= not((layer0_outputs(4611)) xor (layer0_outputs(9151)));
    outputs(8113) <= not((layer0_outputs(6668)) xor (layer0_outputs(6006)));
    outputs(8114) <= (layer0_outputs(1315)) and (layer0_outputs(390));
    outputs(8115) <= layer0_outputs(2763);
    outputs(8116) <= (layer0_outputs(2806)) and (layer0_outputs(6390));
    outputs(8117) <= (layer0_outputs(8867)) xor (layer0_outputs(9746));
    outputs(8118) <= not(layer0_outputs(5668));
    outputs(8119) <= (layer0_outputs(6292)) and not (layer0_outputs(938));
    outputs(8120) <= (layer0_outputs(6989)) xor (layer0_outputs(2074));
    outputs(8121) <= not(layer0_outputs(5227));
    outputs(8122) <= (layer0_outputs(3269)) and (layer0_outputs(4460));
    outputs(8123) <= layer0_outputs(7197);
    outputs(8124) <= layer0_outputs(5198);
    outputs(8125) <= not(layer0_outputs(8145));
    outputs(8126) <= (layer0_outputs(9219)) xor (layer0_outputs(3466));
    outputs(8127) <= (layer0_outputs(4658)) and not (layer0_outputs(5008));
    outputs(8128) <= layer0_outputs(4348);
    outputs(8129) <= not((layer0_outputs(7345)) xor (layer0_outputs(558)));
    outputs(8130) <= not((layer0_outputs(8765)) xor (layer0_outputs(6397)));
    outputs(8131) <= layer0_outputs(1070);
    outputs(8132) <= (layer0_outputs(7963)) and not (layer0_outputs(2178));
    outputs(8133) <= (layer0_outputs(7031)) and not (layer0_outputs(1194));
    outputs(8134) <= not(layer0_outputs(4520));
    outputs(8135) <= (layer0_outputs(4712)) or (layer0_outputs(310));
    outputs(8136) <= (layer0_outputs(265)) or (layer0_outputs(3229));
    outputs(8137) <= (layer0_outputs(8447)) and (layer0_outputs(1818));
    outputs(8138) <= not((layer0_outputs(2019)) xor (layer0_outputs(3530)));
    outputs(8139) <= not((layer0_outputs(10027)) xor (layer0_outputs(3242)));
    outputs(8140) <= (layer0_outputs(5578)) and not (layer0_outputs(285));
    outputs(8141) <= (layer0_outputs(7794)) and not (layer0_outputs(2130));
    outputs(8142) <= not(layer0_outputs(67));
    outputs(8143) <= not((layer0_outputs(4266)) or (layer0_outputs(5346)));
    outputs(8144) <= not(layer0_outputs(9959));
    outputs(8145) <= (layer0_outputs(560)) and not (layer0_outputs(6901));
    outputs(8146) <= not(layer0_outputs(4563));
    outputs(8147) <= (layer0_outputs(6718)) and (layer0_outputs(2475));
    outputs(8148) <= not((layer0_outputs(5549)) xor (layer0_outputs(6084)));
    outputs(8149) <= (layer0_outputs(7130)) xor (layer0_outputs(9100));
    outputs(8150) <= (layer0_outputs(6948)) and not (layer0_outputs(8066));
    outputs(8151) <= layer0_outputs(1377);
    outputs(8152) <= (layer0_outputs(9049)) xor (layer0_outputs(6537));
    outputs(8153) <= (layer0_outputs(4691)) xor (layer0_outputs(7147));
    outputs(8154) <= layer0_outputs(321);
    outputs(8155) <= not(layer0_outputs(9223));
    outputs(8156) <= layer0_outputs(1273);
    outputs(8157) <= not((layer0_outputs(1798)) or (layer0_outputs(9779)));
    outputs(8158) <= layer0_outputs(6357);
    outputs(8159) <= not(layer0_outputs(4508));
    outputs(8160) <= not((layer0_outputs(3310)) or (layer0_outputs(9138)));
    outputs(8161) <= not((layer0_outputs(2404)) xor (layer0_outputs(9888)));
    outputs(8162) <= layer0_outputs(453);
    outputs(8163) <= (layer0_outputs(7833)) xor (layer0_outputs(2511));
    outputs(8164) <= (layer0_outputs(5607)) and (layer0_outputs(6867));
    outputs(8165) <= not(layer0_outputs(4420));
    outputs(8166) <= not((layer0_outputs(1143)) xor (layer0_outputs(4772)));
    outputs(8167) <= (layer0_outputs(1578)) or (layer0_outputs(8797));
    outputs(8168) <= not(layer0_outputs(4087));
    outputs(8169) <= layer0_outputs(5145);
    outputs(8170) <= not(layer0_outputs(361));
    outputs(8171) <= not(layer0_outputs(7461));
    outputs(8172) <= layer0_outputs(6552);
    outputs(8173) <= not(layer0_outputs(8011));
    outputs(8174) <= layer0_outputs(4724);
    outputs(8175) <= not(layer0_outputs(2744));
    outputs(8176) <= layer0_outputs(2375);
    outputs(8177) <= not(layer0_outputs(255));
    outputs(8178) <= layer0_outputs(1657);
    outputs(8179) <= not(layer0_outputs(2776));
    outputs(8180) <= not((layer0_outputs(352)) or (layer0_outputs(2168)));
    outputs(8181) <= (layer0_outputs(1255)) and not (layer0_outputs(6881));
    outputs(8182) <= layer0_outputs(4450);
    outputs(8183) <= not(layer0_outputs(2368)) or (layer0_outputs(7046));
    outputs(8184) <= (layer0_outputs(7804)) xor (layer0_outputs(186));
    outputs(8185) <= not(layer0_outputs(1144));
    outputs(8186) <= layer0_outputs(1963);
    outputs(8187) <= (layer0_outputs(2141)) and not (layer0_outputs(8009));
    outputs(8188) <= layer0_outputs(7894);
    outputs(8189) <= layer0_outputs(9973);
    outputs(8190) <= (layer0_outputs(4671)) and not (layer0_outputs(7722));
    outputs(8191) <= not(layer0_outputs(251));
    outputs(8192) <= not(layer0_outputs(3946)) or (layer0_outputs(6927));
    outputs(8193) <= (layer0_outputs(4394)) or (layer0_outputs(6886));
    outputs(8194) <= (layer0_outputs(3810)) xor (layer0_outputs(7913));
    outputs(8195) <= not(layer0_outputs(9017)) or (layer0_outputs(4585));
    outputs(8196) <= not((layer0_outputs(9237)) xor (layer0_outputs(8167)));
    outputs(8197) <= layer0_outputs(2651);
    outputs(8198) <= layer0_outputs(10041);
    outputs(8199) <= (layer0_outputs(3167)) xor (layer0_outputs(3859));
    outputs(8200) <= (layer0_outputs(8931)) xor (layer0_outputs(8045));
    outputs(8201) <= (layer0_outputs(3325)) xor (layer0_outputs(6001));
    outputs(8202) <= layer0_outputs(8721);
    outputs(8203) <= (layer0_outputs(1689)) and (layer0_outputs(8876));
    outputs(8204) <= layer0_outputs(7490);
    outputs(8205) <= (layer0_outputs(348)) or (layer0_outputs(7304));
    outputs(8206) <= (layer0_outputs(5014)) xor (layer0_outputs(6610));
    outputs(8207) <= not(layer0_outputs(2680));
    outputs(8208) <= not((layer0_outputs(486)) and (layer0_outputs(6497)));
    outputs(8209) <= not((layer0_outputs(10204)) and (layer0_outputs(8916)));
    outputs(8210) <= not(layer0_outputs(2731));
    outputs(8211) <= not(layer0_outputs(4024));
    outputs(8212) <= layer0_outputs(5169);
    outputs(8213) <= layer0_outputs(3533);
    outputs(8214) <= (layer0_outputs(8207)) and not (layer0_outputs(3555));
    outputs(8215) <= not((layer0_outputs(8409)) xor (layer0_outputs(8082)));
    outputs(8216) <= (layer0_outputs(7669)) and (layer0_outputs(3427));
    outputs(8217) <= not(layer0_outputs(6136)) or (layer0_outputs(2884));
    outputs(8218) <= layer0_outputs(2132);
    outputs(8219) <= not(layer0_outputs(2687));
    outputs(8220) <= layer0_outputs(3969);
    outputs(8221) <= not((layer0_outputs(7710)) or (layer0_outputs(4084)));
    outputs(8222) <= not(layer0_outputs(5272));
    outputs(8223) <= not((layer0_outputs(2414)) or (layer0_outputs(8511)));
    outputs(8224) <= not(layer0_outputs(251)) or (layer0_outputs(900));
    outputs(8225) <= (layer0_outputs(222)) or (layer0_outputs(9623));
    outputs(8226) <= not(layer0_outputs(1841)) or (layer0_outputs(1559));
    outputs(8227) <= not((layer0_outputs(5847)) xor (layer0_outputs(1992)));
    outputs(8228) <= not((layer0_outputs(10063)) and (layer0_outputs(9911)));
    outputs(8229) <= layer0_outputs(1787);
    outputs(8230) <= layer0_outputs(4552);
    outputs(8231) <= not(layer0_outputs(5154));
    outputs(8232) <= layer0_outputs(8677);
    outputs(8233) <= (layer0_outputs(3793)) xor (layer0_outputs(3870));
    outputs(8234) <= not((layer0_outputs(8327)) xor (layer0_outputs(4943)));
    outputs(8235) <= not(layer0_outputs(3835));
    outputs(8236) <= layer0_outputs(6979);
    outputs(8237) <= not(layer0_outputs(7418)) or (layer0_outputs(4045));
    outputs(8238) <= not(layer0_outputs(9433));
    outputs(8239) <= (layer0_outputs(6306)) and (layer0_outputs(2553));
    outputs(8240) <= (layer0_outputs(3626)) and not (layer0_outputs(9919));
    outputs(8241) <= not((layer0_outputs(3929)) xor (layer0_outputs(2825)));
    outputs(8242) <= not(layer0_outputs(727));
    outputs(8243) <= not(layer0_outputs(5159));
    outputs(8244) <= (layer0_outputs(124)) and not (layer0_outputs(912));
    outputs(8245) <= not(layer0_outputs(1247));
    outputs(8246) <= layer0_outputs(7438);
    outputs(8247) <= not(layer0_outputs(5942));
    outputs(8248) <= not((layer0_outputs(8003)) xor (layer0_outputs(5913)));
    outputs(8249) <= not((layer0_outputs(7686)) and (layer0_outputs(7463)));
    outputs(8250) <= layer0_outputs(8354);
    outputs(8251) <= not(layer0_outputs(4367)) or (layer0_outputs(7420));
    outputs(8252) <= not(layer0_outputs(5842));
    outputs(8253) <= not(layer0_outputs(4784));
    outputs(8254) <= not(layer0_outputs(4183)) or (layer0_outputs(905));
    outputs(8255) <= not((layer0_outputs(4825)) xor (layer0_outputs(4340)));
    outputs(8256) <= not(layer0_outputs(2929));
    outputs(8257) <= not(layer0_outputs(3379)) or (layer0_outputs(6009));
    outputs(8258) <= not(layer0_outputs(3438));
    outputs(8259) <= not(layer0_outputs(9867));
    outputs(8260) <= (layer0_outputs(5891)) xor (layer0_outputs(8038));
    outputs(8261) <= not((layer0_outputs(6677)) xor (layer0_outputs(8101)));
    outputs(8262) <= not((layer0_outputs(8743)) xor (layer0_outputs(8719)));
    outputs(8263) <= layer0_outputs(3333);
    outputs(8264) <= layer0_outputs(5062);
    outputs(8265) <= layer0_outputs(299);
    outputs(8266) <= not(layer0_outputs(6275));
    outputs(8267) <= not(layer0_outputs(7039));
    outputs(8268) <= not((layer0_outputs(4878)) xor (layer0_outputs(6352)));
    outputs(8269) <= (layer0_outputs(4551)) xor (layer0_outputs(3352));
    outputs(8270) <= not(layer0_outputs(9669)) or (layer0_outputs(4252));
    outputs(8271) <= layer0_outputs(8602);
    outputs(8272) <= (layer0_outputs(8594)) or (layer0_outputs(10031));
    outputs(8273) <= layer0_outputs(7229);
    outputs(8274) <= (layer0_outputs(9794)) xor (layer0_outputs(10091));
    outputs(8275) <= not((layer0_outputs(8055)) xor (layer0_outputs(1991)));
    outputs(8276) <= (layer0_outputs(8052)) xor (layer0_outputs(4787));
    outputs(8277) <= (layer0_outputs(5350)) xor (layer0_outputs(1861));
    outputs(8278) <= layer0_outputs(4143);
    outputs(8279) <= layer0_outputs(5879);
    outputs(8280) <= (layer0_outputs(5133)) xor (layer0_outputs(5504));
    outputs(8281) <= not(layer0_outputs(6373));
    outputs(8282) <= layer0_outputs(496);
    outputs(8283) <= not((layer0_outputs(9294)) xor (layer0_outputs(3095)));
    outputs(8284) <= (layer0_outputs(7077)) xor (layer0_outputs(7962));
    outputs(8285) <= not(layer0_outputs(7179));
    outputs(8286) <= (layer0_outputs(5542)) xor (layer0_outputs(3548));
    outputs(8287) <= (layer0_outputs(1871)) xor (layer0_outputs(3017));
    outputs(8288) <= not(layer0_outputs(5999)) or (layer0_outputs(7695));
    outputs(8289) <= layer0_outputs(5733);
    outputs(8290) <= (layer0_outputs(3200)) or (layer0_outputs(5468));
    outputs(8291) <= not(layer0_outputs(3925));
    outputs(8292) <= not(layer0_outputs(412));
    outputs(8293) <= (layer0_outputs(7118)) xor (layer0_outputs(8774));
    outputs(8294) <= not((layer0_outputs(9761)) or (layer0_outputs(8198)));
    outputs(8295) <= not(layer0_outputs(3905));
    outputs(8296) <= not(layer0_outputs(8238));
    outputs(8297) <= not(layer0_outputs(6114));
    outputs(8298) <= not((layer0_outputs(9744)) and (layer0_outputs(2973)));
    outputs(8299) <= layer0_outputs(1243);
    outputs(8300) <= layer0_outputs(2191);
    outputs(8301) <= layer0_outputs(1202);
    outputs(8302) <= not(layer0_outputs(7989)) or (layer0_outputs(36));
    outputs(8303) <= layer0_outputs(6500);
    outputs(8304) <= not(layer0_outputs(8180));
    outputs(8305) <= not(layer0_outputs(2894));
    outputs(8306) <= (layer0_outputs(4084)) xor (layer0_outputs(8383));
    outputs(8307) <= not((layer0_outputs(2100)) or (layer0_outputs(528)));
    outputs(8308) <= not((layer0_outputs(631)) or (layer0_outputs(983)));
    outputs(8309) <= not(layer0_outputs(4336));
    outputs(8310) <= (layer0_outputs(9690)) xor (layer0_outputs(3747));
    outputs(8311) <= not(layer0_outputs(5303)) or (layer0_outputs(4811));
    outputs(8312) <= (layer0_outputs(1823)) xor (layer0_outputs(10030));
    outputs(8313) <= not((layer0_outputs(5893)) and (layer0_outputs(6579)));
    outputs(8314) <= layer0_outputs(6829);
    outputs(8315) <= (layer0_outputs(8279)) and not (layer0_outputs(6722));
    outputs(8316) <= not(layer0_outputs(6645)) or (layer0_outputs(7341));
    outputs(8317) <= not((layer0_outputs(1599)) and (layer0_outputs(2688)));
    outputs(8318) <= (layer0_outputs(7135)) xor (layer0_outputs(7541));
    outputs(8319) <= layer0_outputs(1654);
    outputs(8320) <= layer0_outputs(2309);
    outputs(8321) <= not((layer0_outputs(10193)) xor (layer0_outputs(3466)));
    outputs(8322) <= not(layer0_outputs(9221));
    outputs(8323) <= layer0_outputs(3701);
    outputs(8324) <= layer0_outputs(7766);
    outputs(8325) <= layer0_outputs(7593);
    outputs(8326) <= not(layer0_outputs(7433)) or (layer0_outputs(3240));
    outputs(8327) <= not(layer0_outputs(2935));
    outputs(8328) <= not(layer0_outputs(6924));
    outputs(8329) <= layer0_outputs(4991);
    outputs(8330) <= not((layer0_outputs(2224)) and (layer0_outputs(9657)));
    outputs(8331) <= (layer0_outputs(2376)) and (layer0_outputs(1257));
    outputs(8332) <= not(layer0_outputs(7301)) or (layer0_outputs(9693));
    outputs(8333) <= not(layer0_outputs(7871));
    outputs(8334) <= not((layer0_outputs(7338)) xor (layer0_outputs(2556)));
    outputs(8335) <= (layer0_outputs(8648)) and not (layer0_outputs(659));
    outputs(8336) <= layer0_outputs(4674);
    outputs(8337) <= not((layer0_outputs(4116)) xor (layer0_outputs(3405)));
    outputs(8338) <= (layer0_outputs(6449)) xor (layer0_outputs(4672));
    outputs(8339) <= (layer0_outputs(9455)) xor (layer0_outputs(9456));
    outputs(8340) <= not(layer0_outputs(1208)) or (layer0_outputs(4964));
    outputs(8341) <= layer0_outputs(4048);
    outputs(8342) <= not(layer0_outputs(8109)) or (layer0_outputs(8990));
    outputs(8343) <= not(layer0_outputs(2045));
    outputs(8344) <= layer0_outputs(2198);
    outputs(8345) <= not((layer0_outputs(5770)) xor (layer0_outputs(296)));
    outputs(8346) <= not(layer0_outputs(5051));
    outputs(8347) <= not(layer0_outputs(4574)) or (layer0_outputs(792));
    outputs(8348) <= not(layer0_outputs(2211));
    outputs(8349) <= not((layer0_outputs(7867)) xor (layer0_outputs(763)));
    outputs(8350) <= not((layer0_outputs(6781)) xor (layer0_outputs(327)));
    outputs(8351) <= layer0_outputs(6071);
    outputs(8352) <= (layer0_outputs(2925)) or (layer0_outputs(654));
    outputs(8353) <= layer0_outputs(3512);
    outputs(8354) <= (layer0_outputs(10127)) or (layer0_outputs(7620));
    outputs(8355) <= layer0_outputs(525);
    outputs(8356) <= not((layer0_outputs(749)) xor (layer0_outputs(4973)));
    outputs(8357) <= not(layer0_outputs(6302));
    outputs(8358) <= not(layer0_outputs(1002));
    outputs(8359) <= (layer0_outputs(5915)) xor (layer0_outputs(1260));
    outputs(8360) <= layer0_outputs(8796);
    outputs(8361) <= not(layer0_outputs(10135));
    outputs(8362) <= not((layer0_outputs(9699)) and (layer0_outputs(8983)));
    outputs(8363) <= not(layer0_outputs(298)) or (layer0_outputs(9826));
    outputs(8364) <= not(layer0_outputs(643));
    outputs(8365) <= not(layer0_outputs(1915));
    outputs(8366) <= (layer0_outputs(9444)) xor (layer0_outputs(9452));
    outputs(8367) <= (layer0_outputs(1049)) or (layer0_outputs(2988));
    outputs(8368) <= not((layer0_outputs(7297)) and (layer0_outputs(2147)));
    outputs(8369) <= not((layer0_outputs(1982)) xor (layer0_outputs(3066)));
    outputs(8370) <= not(layer0_outputs(5877)) or (layer0_outputs(334));
    outputs(8371) <= layer0_outputs(8099);
    outputs(8372) <= not(layer0_outputs(5105));
    outputs(8373) <= layer0_outputs(4640);
    outputs(8374) <= not((layer0_outputs(2641)) xor (layer0_outputs(1946)));
    outputs(8375) <= (layer0_outputs(4621)) xor (layer0_outputs(6774));
    outputs(8376) <= not(layer0_outputs(4651)) or (layer0_outputs(10025));
    outputs(8377) <= layer0_outputs(9659);
    outputs(8378) <= not(layer0_outputs(4100));
    outputs(8379) <= not(layer0_outputs(8841)) or (layer0_outputs(4008));
    outputs(8380) <= not(layer0_outputs(4091));
    outputs(8381) <= not((layer0_outputs(6523)) xor (layer0_outputs(9938)));
    outputs(8382) <= layer0_outputs(6177);
    outputs(8383) <= not((layer0_outputs(4471)) xor (layer0_outputs(1284)));
    outputs(8384) <= not(layer0_outputs(2815));
    outputs(8385) <= (layer0_outputs(2712)) xor (layer0_outputs(7137));
    outputs(8386) <= (layer0_outputs(9343)) xor (layer0_outputs(2472));
    outputs(8387) <= '1';
    outputs(8388) <= (layer0_outputs(1024)) xor (layer0_outputs(7013));
    outputs(8389) <= (layer0_outputs(10114)) or (layer0_outputs(2433));
    outputs(8390) <= (layer0_outputs(2095)) xor (layer0_outputs(2528));
    outputs(8391) <= not(layer0_outputs(9457)) or (layer0_outputs(7310));
    outputs(8392) <= not(layer0_outputs(645));
    outputs(8393) <= not(layer0_outputs(1949)) or (layer0_outputs(8590));
    outputs(8394) <= not((layer0_outputs(6494)) xor (layer0_outputs(7692)));
    outputs(8395) <= '1';
    outputs(8396) <= not(layer0_outputs(9372));
    outputs(8397) <= not((layer0_outputs(1630)) xor (layer0_outputs(849)));
    outputs(8398) <= not((layer0_outputs(8817)) xor (layer0_outputs(6813)));
    outputs(8399) <= not(layer0_outputs(4284));
    outputs(8400) <= not((layer0_outputs(3868)) or (layer0_outputs(8282)));
    outputs(8401) <= not(layer0_outputs(9583));
    outputs(8402) <= not((layer0_outputs(2320)) xor (layer0_outputs(927)));
    outputs(8403) <= not((layer0_outputs(3021)) xor (layer0_outputs(7910)));
    outputs(8404) <= layer0_outputs(4230);
    outputs(8405) <= not(layer0_outputs(5498));
    outputs(8406) <= not(layer0_outputs(955));
    outputs(8407) <= not((layer0_outputs(9769)) xor (layer0_outputs(3675)));
    outputs(8408) <= layer0_outputs(5422);
    outputs(8409) <= (layer0_outputs(8083)) and not (layer0_outputs(6459));
    outputs(8410) <= not(layer0_outputs(7535)) or (layer0_outputs(1624));
    outputs(8411) <= not((layer0_outputs(6171)) xor (layer0_outputs(4042)));
    outputs(8412) <= not(layer0_outputs(5906)) or (layer0_outputs(4153));
    outputs(8413) <= (layer0_outputs(9454)) and not (layer0_outputs(5445));
    outputs(8414) <= not(layer0_outputs(8359));
    outputs(8415) <= not(layer0_outputs(4849)) or (layer0_outputs(2490));
    outputs(8416) <= not(layer0_outputs(148));
    outputs(8417) <= not(layer0_outputs(2286)) or (layer0_outputs(1314));
    outputs(8418) <= not(layer0_outputs(1900));
    outputs(8419) <= not(layer0_outputs(7613));
    outputs(8420) <= (layer0_outputs(6630)) xor (layer0_outputs(7685));
    outputs(8421) <= layer0_outputs(3614);
    outputs(8422) <= layer0_outputs(4528);
    outputs(8423) <= not(layer0_outputs(7403)) or (layer0_outputs(6206));
    outputs(8424) <= not((layer0_outputs(3591)) xor (layer0_outputs(5824)));
    outputs(8425) <= not((layer0_outputs(2969)) or (layer0_outputs(6705)));
    outputs(8426) <= (layer0_outputs(4862)) and not (layer0_outputs(10227));
    outputs(8427) <= not(layer0_outputs(945)) or (layer0_outputs(1172));
    outputs(8428) <= not(layer0_outputs(5260)) or (layer0_outputs(9941));
    outputs(8429) <= layer0_outputs(5348);
    outputs(8430) <= layer0_outputs(6118);
    outputs(8431) <= layer0_outputs(5788);
    outputs(8432) <= (layer0_outputs(404)) and not (layer0_outputs(9417));
    outputs(8433) <= (layer0_outputs(7123)) or (layer0_outputs(9873));
    outputs(8434) <= (layer0_outputs(2110)) or (layer0_outputs(6255));
    outputs(8435) <= not((layer0_outputs(9003)) xor (layer0_outputs(2735)));
    outputs(8436) <= (layer0_outputs(31)) xor (layer0_outputs(2128));
    outputs(8437) <= not((layer0_outputs(6035)) xor (layer0_outputs(2482)));
    outputs(8438) <= not(layer0_outputs(166));
    outputs(8439) <= not((layer0_outputs(9382)) and (layer0_outputs(9394)));
    outputs(8440) <= not((layer0_outputs(4323)) xor (layer0_outputs(2031)));
    outputs(8441) <= (layer0_outputs(9030)) and not (layer0_outputs(7040));
    outputs(8442) <= (layer0_outputs(9651)) and not (layer0_outputs(4934));
    outputs(8443) <= not(layer0_outputs(4227));
    outputs(8444) <= layer0_outputs(10161);
    outputs(8445) <= not(layer0_outputs(7528));
    outputs(8446) <= not((layer0_outputs(7911)) xor (layer0_outputs(6822)));
    outputs(8447) <= layer0_outputs(3273);
    outputs(8448) <= not((layer0_outputs(2576)) and (layer0_outputs(8433)));
    outputs(8449) <= not((layer0_outputs(4220)) xor (layer0_outputs(9265)));
    outputs(8450) <= not(layer0_outputs(8342));
    outputs(8451) <= layer0_outputs(8064);
    outputs(8452) <= (layer0_outputs(6132)) and not (layer0_outputs(7796));
    outputs(8453) <= (layer0_outputs(7244)) and (layer0_outputs(8571));
    outputs(8454) <= (layer0_outputs(3188)) xor (layer0_outputs(599));
    outputs(8455) <= not(layer0_outputs(3106)) or (layer0_outputs(9179));
    outputs(8456) <= not((layer0_outputs(4863)) xor (layer0_outputs(7252)));
    outputs(8457) <= not((layer0_outputs(1282)) xor (layer0_outputs(6276)));
    outputs(8458) <= (layer0_outputs(5185)) and not (layer0_outputs(5175));
    outputs(8459) <= not(layer0_outputs(10175)) or (layer0_outputs(9565));
    outputs(8460) <= not((layer0_outputs(5187)) xor (layer0_outputs(8744)));
    outputs(8461) <= (layer0_outputs(8209)) xor (layer0_outputs(8183));
    outputs(8462) <= not(layer0_outputs(6192)) or (layer0_outputs(2926));
    outputs(8463) <= (layer0_outputs(7218)) or (layer0_outputs(3827));
    outputs(8464) <= not(layer0_outputs(5338));
    outputs(8465) <= not((layer0_outputs(271)) xor (layer0_outputs(8076)));
    outputs(8466) <= layer0_outputs(8583);
    outputs(8467) <= not((layer0_outputs(1731)) xor (layer0_outputs(3337)));
    outputs(8468) <= (layer0_outputs(10239)) xor (layer0_outputs(8013));
    outputs(8469) <= layer0_outputs(245);
    outputs(8470) <= (layer0_outputs(1929)) and not (layer0_outputs(2145));
    outputs(8471) <= not(layer0_outputs(1161));
    outputs(8472) <= not(layer0_outputs(7573));
    outputs(8473) <= not(layer0_outputs(5705));
    outputs(8474) <= not(layer0_outputs(9924)) or (layer0_outputs(867));
    outputs(8475) <= not(layer0_outputs(4000));
    outputs(8476) <= (layer0_outputs(7801)) xor (layer0_outputs(8966));
    outputs(8477) <= not(layer0_outputs(767));
    outputs(8478) <= layer0_outputs(6325);
    outputs(8479) <= not(layer0_outputs(9060));
    outputs(8480) <= (layer0_outputs(3763)) xor (layer0_outputs(5774));
    outputs(8481) <= layer0_outputs(9814);
    outputs(8482) <= not(layer0_outputs(2079));
    outputs(8483) <= not(layer0_outputs(1021)) or (layer0_outputs(3343));
    outputs(8484) <= (layer0_outputs(2237)) and not (layer0_outputs(8513));
    outputs(8485) <= not(layer0_outputs(1232));
    outputs(8486) <= (layer0_outputs(6207)) or (layer0_outputs(2746));
    outputs(8487) <= layer0_outputs(3328);
    outputs(8488) <= not(layer0_outputs(518));
    outputs(8489) <= (layer0_outputs(6600)) or (layer0_outputs(9891));
    outputs(8490) <= layer0_outputs(9203);
    outputs(8491) <= not((layer0_outputs(4537)) and (layer0_outputs(7018)));
    outputs(8492) <= not((layer0_outputs(10233)) xor (layer0_outputs(4910)));
    outputs(8493) <= (layer0_outputs(561)) xor (layer0_outputs(8893));
    outputs(8494) <= (layer0_outputs(2689)) and not (layer0_outputs(5216));
    outputs(8495) <= layer0_outputs(1628);
    outputs(8496) <= not(layer0_outputs(3351)) or (layer0_outputs(9252));
    outputs(8497) <= not(layer0_outputs(1499));
    outputs(8498) <= (layer0_outputs(258)) xor (layer0_outputs(6346));
    outputs(8499) <= layer0_outputs(5975);
    outputs(8500) <= not(layer0_outputs(1726));
    outputs(8501) <= not(layer0_outputs(4489));
    outputs(8502) <= layer0_outputs(2455);
    outputs(8503) <= not((layer0_outputs(1971)) xor (layer0_outputs(1644)));
    outputs(8504) <= (layer0_outputs(8010)) xor (layer0_outputs(2526));
    outputs(8505) <= not(layer0_outputs(8194));
    outputs(8506) <= layer0_outputs(2932);
    outputs(8507) <= layer0_outputs(6364);
    outputs(8508) <= not(layer0_outputs(9599));
    outputs(8509) <= not((layer0_outputs(3794)) xor (layer0_outputs(9668)));
    outputs(8510) <= not(layer0_outputs(9626));
    outputs(8511) <= not(layer0_outputs(8331)) or (layer0_outputs(4451));
    outputs(8512) <= (layer0_outputs(7823)) and not (layer0_outputs(1346));
    outputs(8513) <= layer0_outputs(2593);
    outputs(8514) <= (layer0_outputs(410)) xor (layer0_outputs(660));
    outputs(8515) <= (layer0_outputs(5168)) or (layer0_outputs(4452));
    outputs(8516) <= not(layer0_outputs(8405));
    outputs(8517) <= (layer0_outputs(7143)) and not (layer0_outputs(8982));
    outputs(8518) <= not(layer0_outputs(7322)) or (layer0_outputs(4233));
    outputs(8519) <= not((layer0_outputs(8715)) xor (layer0_outputs(577)));
    outputs(8520) <= (layer0_outputs(4035)) xor (layer0_outputs(3703));
    outputs(8521) <= not((layer0_outputs(7562)) and (layer0_outputs(4515)));
    outputs(8522) <= layer0_outputs(4984);
    outputs(8523) <= (layer0_outputs(9951)) xor (layer0_outputs(9268));
    outputs(8524) <= not(layer0_outputs(2170));
    outputs(8525) <= not((layer0_outputs(4792)) xor (layer0_outputs(5108)));
    outputs(8526) <= layer0_outputs(9683);
    outputs(8527) <= layer0_outputs(7369);
    outputs(8528) <= (layer0_outputs(9573)) xor (layer0_outputs(1555));
    outputs(8529) <= (layer0_outputs(1111)) xor (layer0_outputs(5502));
    outputs(8530) <= (layer0_outputs(9594)) and not (layer0_outputs(135));
    outputs(8531) <= (layer0_outputs(20)) and (layer0_outputs(8013));
    outputs(8532) <= not(layer0_outputs(4253));
    outputs(8533) <= (layer0_outputs(3633)) and not (layer0_outputs(770));
    outputs(8534) <= not(layer0_outputs(2784)) or (layer0_outputs(5950));
    outputs(8535) <= layer0_outputs(849);
    outputs(8536) <= not(layer0_outputs(1002));
    outputs(8537) <= (layer0_outputs(8454)) xor (layer0_outputs(9063));
    outputs(8538) <= not(layer0_outputs(6033));
    outputs(8539) <= layer0_outputs(1228);
    outputs(8540) <= not(layer0_outputs(7047));
    outputs(8541) <= (layer0_outputs(5756)) and not (layer0_outputs(1593));
    outputs(8542) <= not((layer0_outputs(5806)) and (layer0_outputs(9011)));
    outputs(8543) <= layer0_outputs(4324);
    outputs(8544) <= (layer0_outputs(7785)) xor (layer0_outputs(5126));
    outputs(8545) <= (layer0_outputs(3967)) or (layer0_outputs(2651));
    outputs(8546) <= layer0_outputs(6966);
    outputs(8547) <= not(layer0_outputs(2009));
    outputs(8548) <= not((layer0_outputs(6367)) xor (layer0_outputs(1745)));
    outputs(8549) <= not((layer0_outputs(1510)) xor (layer0_outputs(376)));
    outputs(8550) <= not(layer0_outputs(7088));
    outputs(8551) <= not((layer0_outputs(876)) and (layer0_outputs(9102)));
    outputs(8552) <= (layer0_outputs(4266)) or (layer0_outputs(3032));
    outputs(8553) <= not((layer0_outputs(2062)) and (layer0_outputs(6348)));
    outputs(8554) <= not(layer0_outputs(3591));
    outputs(8555) <= (layer0_outputs(1893)) xor (layer0_outputs(1697));
    outputs(8556) <= layer0_outputs(4682);
    outputs(8557) <= not(layer0_outputs(1150));
    outputs(8558) <= not(layer0_outputs(1124));
    outputs(8559) <= not(layer0_outputs(706)) or (layer0_outputs(3533));
    outputs(8560) <= layer0_outputs(5282);
    outputs(8561) <= layer0_outputs(9281);
    outputs(8562) <= not((layer0_outputs(3112)) xor (layer0_outputs(4403)));
    outputs(8563) <= (layer0_outputs(5565)) and not (layer0_outputs(3292));
    outputs(8564) <= not((layer0_outputs(8349)) or (layer0_outputs(7954)));
    outputs(8565) <= (layer0_outputs(2602)) or (layer0_outputs(9077));
    outputs(8566) <= (layer0_outputs(3945)) xor (layer0_outputs(3460));
    outputs(8567) <= layer0_outputs(2354);
    outputs(8568) <= (layer0_outputs(5727)) or (layer0_outputs(9807));
    outputs(8569) <= (layer0_outputs(9009)) xor (layer0_outputs(7785));
    outputs(8570) <= layer0_outputs(10099);
    outputs(8571) <= layer0_outputs(8520);
    outputs(8572) <= (layer0_outputs(3381)) or (layer0_outputs(948));
    outputs(8573) <= not(layer0_outputs(955));
    outputs(8574) <= not((layer0_outputs(2253)) xor (layer0_outputs(5742)));
    outputs(8575) <= layer0_outputs(8459);
    outputs(8576) <= (layer0_outputs(6709)) xor (layer0_outputs(7274));
    outputs(8577) <= not((layer0_outputs(9167)) and (layer0_outputs(2569)));
    outputs(8578) <= (layer0_outputs(4701)) xor (layer0_outputs(916));
    outputs(8579) <= layer0_outputs(2227);
    outputs(8580) <= (layer0_outputs(3071)) or (layer0_outputs(2665));
    outputs(8581) <= (layer0_outputs(3152)) xor (layer0_outputs(7281));
    outputs(8582) <= layer0_outputs(7000);
    outputs(8583) <= not(layer0_outputs(4191));
    outputs(8584) <= not((layer0_outputs(10227)) xor (layer0_outputs(8585)));
    outputs(8585) <= (layer0_outputs(1652)) xor (layer0_outputs(4620));
    outputs(8586) <= layer0_outputs(1856);
    outputs(8587) <= not(layer0_outputs(7583));
    outputs(8588) <= layer0_outputs(3357);
    outputs(8589) <= not((layer0_outputs(1551)) xor (layer0_outputs(2764)));
    outputs(8590) <= not(layer0_outputs(8790)) or (layer0_outputs(4913));
    outputs(8591) <= (layer0_outputs(6825)) xor (layer0_outputs(2554));
    outputs(8592) <= not((layer0_outputs(2668)) and (layer0_outputs(6183)));
    outputs(8593) <= not(layer0_outputs(416)) or (layer0_outputs(8746));
    outputs(8594) <= not(layer0_outputs(8907));
    outputs(8595) <= layer0_outputs(562);
    outputs(8596) <= not(layer0_outputs(5965)) or (layer0_outputs(8420));
    outputs(8597) <= not(layer0_outputs(6265));
    outputs(8598) <= not((layer0_outputs(8595)) and (layer0_outputs(3726)));
    outputs(8599) <= not(layer0_outputs(1079)) or (layer0_outputs(6920));
    outputs(8600) <= not((layer0_outputs(4486)) and (layer0_outputs(9887)));
    outputs(8601) <= (layer0_outputs(772)) xor (layer0_outputs(578));
    outputs(8602) <= (layer0_outputs(5799)) or (layer0_outputs(5789));
    outputs(8603) <= not(layer0_outputs(5248)) or (layer0_outputs(1945));
    outputs(8604) <= not((layer0_outputs(6828)) xor (layer0_outputs(5286)));
    outputs(8605) <= (layer0_outputs(4647)) and not (layer0_outputs(3162));
    outputs(8606) <= not((layer0_outputs(8719)) xor (layer0_outputs(2830)));
    outputs(8607) <= not(layer0_outputs(5576));
    outputs(8608) <= not(layer0_outputs(6615)) or (layer0_outputs(4932));
    outputs(8609) <= (layer0_outputs(1785)) xor (layer0_outputs(6631));
    outputs(8610) <= not((layer0_outputs(2769)) or (layer0_outputs(5845)));
    outputs(8611) <= not(layer0_outputs(4132)) or (layer0_outputs(3395));
    outputs(8612) <= (layer0_outputs(7986)) or (layer0_outputs(4268));
    outputs(8613) <= not(layer0_outputs(4851)) or (layer0_outputs(5917));
    outputs(8614) <= not((layer0_outputs(8397)) xor (layer0_outputs(1026)));
    outputs(8615) <= not(layer0_outputs(2771));
    outputs(8616) <= not(layer0_outputs(4740));
    outputs(8617) <= (layer0_outputs(6999)) xor (layer0_outputs(2883));
    outputs(8618) <= not(layer0_outputs(5390)) or (layer0_outputs(3531));
    outputs(8619) <= (layer0_outputs(7012)) xor (layer0_outputs(5655));
    outputs(8620) <= not(layer0_outputs(6873));
    outputs(8621) <= layer0_outputs(9972);
    outputs(8622) <= (layer0_outputs(2384)) xor (layer0_outputs(8523));
    outputs(8623) <= (layer0_outputs(8319)) xor (layer0_outputs(9060));
    outputs(8624) <= layer0_outputs(4756);
    outputs(8625) <= not(layer0_outputs(827));
    outputs(8626) <= not((layer0_outputs(9874)) xor (layer0_outputs(7542)));
    outputs(8627) <= not(layer0_outputs(8371)) or (layer0_outputs(6511));
    outputs(8628) <= layer0_outputs(4727);
    outputs(8629) <= not(layer0_outputs(6869)) or (layer0_outputs(2961));
    outputs(8630) <= (layer0_outputs(10209)) xor (layer0_outputs(9391));
    outputs(8631) <= not(layer0_outputs(2018)) or (layer0_outputs(9678));
    outputs(8632) <= (layer0_outputs(4982)) xor (layer0_outputs(5940));
    outputs(8633) <= not((layer0_outputs(1472)) xor (layer0_outputs(6484)));
    outputs(8634) <= not((layer0_outputs(1885)) and (layer0_outputs(4346)));
    outputs(8635) <= not(layer0_outputs(4331));
    outputs(8636) <= not(layer0_outputs(9687)) or (layer0_outputs(7002));
    outputs(8637) <= not((layer0_outputs(8614)) xor (layer0_outputs(3)));
    outputs(8638) <= layer0_outputs(399);
    outputs(8639) <= (layer0_outputs(1524)) and (layer0_outputs(9512));
    outputs(8640) <= not(layer0_outputs(341));
    outputs(8641) <= not((layer0_outputs(4550)) xor (layer0_outputs(4273)));
    outputs(8642) <= layer0_outputs(3951);
    outputs(8643) <= (layer0_outputs(7236)) xor (layer0_outputs(8480));
    outputs(8644) <= not((layer0_outputs(9231)) xor (layer0_outputs(5739)));
    outputs(8645) <= not((layer0_outputs(10017)) or (layer0_outputs(7502)));
    outputs(8646) <= (layer0_outputs(3700)) and not (layer0_outputs(9772));
    outputs(8647) <= not(layer0_outputs(3618));
    outputs(8648) <= not(layer0_outputs(454)) or (layer0_outputs(6183));
    outputs(8649) <= layer0_outputs(1849);
    outputs(8650) <= not(layer0_outputs(7665));
    outputs(8651) <= not(layer0_outputs(4286));
    outputs(8652) <= not(layer0_outputs(3564));
    outputs(8653) <= not(layer0_outputs(173));
    outputs(8654) <= not(layer0_outputs(5995)) or (layer0_outputs(4693));
    outputs(8655) <= not(layer0_outputs(3005));
    outputs(8656) <= not(layer0_outputs(6873));
    outputs(8657) <= (layer0_outputs(4435)) xor (layer0_outputs(5106));
    outputs(8658) <= (layer0_outputs(8298)) xor (layer0_outputs(2556));
    outputs(8659) <= layer0_outputs(4827);
    outputs(8660) <= not(layer0_outputs(6240));
    outputs(8661) <= (layer0_outputs(680)) xor (layer0_outputs(3865));
    outputs(8662) <= not((layer0_outputs(9234)) and (layer0_outputs(7831)));
    outputs(8663) <= layer0_outputs(9834);
    outputs(8664) <= not(layer0_outputs(10070));
    outputs(8665) <= not(layer0_outputs(2158));
    outputs(8666) <= not((layer0_outputs(6294)) and (layer0_outputs(6336)));
    outputs(8667) <= (layer0_outputs(4750)) xor (layer0_outputs(1911));
    outputs(8668) <= not((layer0_outputs(8342)) xor (layer0_outputs(5084)));
    outputs(8669) <= layer0_outputs(2269);
    outputs(8670) <= not(layer0_outputs(8424));
    outputs(8671) <= not((layer0_outputs(1526)) xor (layer0_outputs(2304)));
    outputs(8672) <= layer0_outputs(9738);
    outputs(8673) <= not((layer0_outputs(4136)) and (layer0_outputs(8222)));
    outputs(8674) <= not(layer0_outputs(3432)) or (layer0_outputs(4523));
    outputs(8675) <= not(layer0_outputs(1678)) or (layer0_outputs(5141));
    outputs(8676) <= (layer0_outputs(3627)) and not (layer0_outputs(9902));
    outputs(8677) <= (layer0_outputs(10112)) and (layer0_outputs(6487));
    outputs(8678) <= not(layer0_outputs(5112));
    outputs(8679) <= not((layer0_outputs(1519)) xor (layer0_outputs(3202)));
    outputs(8680) <= not(layer0_outputs(7724)) or (layer0_outputs(1686));
    outputs(8681) <= layer0_outputs(1465);
    outputs(8682) <= not(layer0_outputs(8666));
    outputs(8683) <= not((layer0_outputs(3439)) or (layer0_outputs(9406)));
    outputs(8684) <= not((layer0_outputs(1080)) xor (layer0_outputs(2473)));
    outputs(8685) <= layer0_outputs(7051);
    outputs(8686) <= layer0_outputs(5132);
    outputs(8687) <= not(layer0_outputs(2064));
    outputs(8688) <= not(layer0_outputs(2315));
    outputs(8689) <= not(layer0_outputs(3237));
    outputs(8690) <= not((layer0_outputs(3621)) xor (layer0_outputs(7957)));
    outputs(8691) <= not((layer0_outputs(9145)) and (layer0_outputs(4426)));
    outputs(8692) <= not((layer0_outputs(2676)) xor (layer0_outputs(6500)));
    outputs(8693) <= not(layer0_outputs(7557)) or (layer0_outputs(9479));
    outputs(8694) <= not((layer0_outputs(8988)) and (layer0_outputs(3232)));
    outputs(8695) <= not((layer0_outputs(10003)) xor (layer0_outputs(1817)));
    outputs(8696) <= not(layer0_outputs(749));
    outputs(8697) <= (layer0_outputs(10005)) xor (layer0_outputs(10107));
    outputs(8698) <= layer0_outputs(1640);
    outputs(8699) <= (layer0_outputs(8231)) xor (layer0_outputs(2201));
    outputs(8700) <= not(layer0_outputs(4425));
    outputs(8701) <= not((layer0_outputs(93)) xor (layer0_outputs(2809)));
    outputs(8702) <= not((layer0_outputs(9048)) xor (layer0_outputs(2609)));
    outputs(8703) <= layer0_outputs(7919);
    outputs(8704) <= not(layer0_outputs(3801)) or (layer0_outputs(8459));
    outputs(8705) <= not(layer0_outputs(798)) or (layer0_outputs(324));
    outputs(8706) <= not(layer0_outputs(1457));
    outputs(8707) <= layer0_outputs(8079);
    outputs(8708) <= layer0_outputs(8780);
    outputs(8709) <= layer0_outputs(6225);
    outputs(8710) <= layer0_outputs(4664);
    outputs(8711) <= (layer0_outputs(4209)) and (layer0_outputs(8380));
    outputs(8712) <= (layer0_outputs(4686)) or (layer0_outputs(3425));
    outputs(8713) <= not((layer0_outputs(7865)) xor (layer0_outputs(2431)));
    outputs(8714) <= not(layer0_outputs(2176));
    outputs(8715) <= not(layer0_outputs(7659)) or (layer0_outputs(9846));
    outputs(8716) <= not(layer0_outputs(5689));
    outputs(8717) <= not(layer0_outputs(1478));
    outputs(8718) <= not((layer0_outputs(3385)) xor (layer0_outputs(6642)));
    outputs(8719) <= (layer0_outputs(10166)) xor (layer0_outputs(3223));
    outputs(8720) <= layer0_outputs(8296);
    outputs(8721) <= (layer0_outputs(8368)) xor (layer0_outputs(2713));
    outputs(8722) <= (layer0_outputs(2043)) or (layer0_outputs(4766));
    outputs(8723) <= (layer0_outputs(1517)) or (layer0_outputs(8970));
    outputs(8724) <= layer0_outputs(6640);
    outputs(8725) <= not(layer0_outputs(8359));
    outputs(8726) <= not((layer0_outputs(9743)) xor (layer0_outputs(10046)));
    outputs(8727) <= (layer0_outputs(3349)) xor (layer0_outputs(527));
    outputs(8728) <= layer0_outputs(1527);
    outputs(8729) <= not(layer0_outputs(851));
    outputs(8730) <= not((layer0_outputs(7173)) xor (layer0_outputs(2039)));
    outputs(8731) <= (layer0_outputs(8519)) and not (layer0_outputs(8346));
    outputs(8732) <= (layer0_outputs(9314)) xor (layer0_outputs(7674));
    outputs(8733) <= layer0_outputs(1364);
    outputs(8734) <= not(layer0_outputs(3509));
    outputs(8735) <= (layer0_outputs(8487)) or (layer0_outputs(4400));
    outputs(8736) <= (layer0_outputs(9161)) and not (layer0_outputs(6053));
    outputs(8737) <= not(layer0_outputs(2986)) or (layer0_outputs(9982));
    outputs(8738) <= not(layer0_outputs(4309));
    outputs(8739) <= (layer0_outputs(1496)) xor (layer0_outputs(5880));
    outputs(8740) <= not((layer0_outputs(5644)) xor (layer0_outputs(398)));
    outputs(8741) <= not((layer0_outputs(9984)) and (layer0_outputs(3190)));
    outputs(8742) <= not(layer0_outputs(2496));
    outputs(8743) <= (layer0_outputs(1048)) xor (layer0_outputs(1987));
    outputs(8744) <= not(layer0_outputs(4175)) or (layer0_outputs(9306));
    outputs(8745) <= (layer0_outputs(1431)) xor (layer0_outputs(6887));
    outputs(8746) <= layer0_outputs(4143);
    outputs(8747) <= layer0_outputs(2839);
    outputs(8748) <= not(layer0_outputs(1289));
    outputs(8749) <= not(layer0_outputs(8156));
    outputs(8750) <= (layer0_outputs(1883)) or (layer0_outputs(972));
    outputs(8751) <= not(layer0_outputs(870));
    outputs(8752) <= layer0_outputs(1859);
    outputs(8753) <= (layer0_outputs(2888)) xor (layer0_outputs(7370));
    outputs(8754) <= layer0_outputs(8691);
    outputs(8755) <= not(layer0_outputs(6372)) or (layer0_outputs(2752));
    outputs(8756) <= (layer0_outputs(9101)) xor (layer0_outputs(281));
    outputs(8757) <= not((layer0_outputs(2463)) xor (layer0_outputs(10174)));
    outputs(8758) <= layer0_outputs(4759);
    outputs(8759) <= not((layer0_outputs(3154)) xor (layer0_outputs(543)));
    outputs(8760) <= not((layer0_outputs(5113)) xor (layer0_outputs(5542)));
    outputs(8761) <= not(layer0_outputs(5618));
    outputs(8762) <= not(layer0_outputs(3983));
    outputs(8763) <= not(layer0_outputs(8092));
    outputs(8764) <= not(layer0_outputs(7183));
    outputs(8765) <= not(layer0_outputs(9046)) or (layer0_outputs(6986));
    outputs(8766) <= not(layer0_outputs(5584));
    outputs(8767) <= not(layer0_outputs(8768)) or (layer0_outputs(5797));
    outputs(8768) <= not(layer0_outputs(1248));
    outputs(8769) <= not((layer0_outputs(8606)) xor (layer0_outputs(9329)));
    outputs(8770) <= layer0_outputs(1869);
    outputs(8771) <= not((layer0_outputs(2819)) xor (layer0_outputs(6566)));
    outputs(8772) <= not(layer0_outputs(393));
    outputs(8773) <= not((layer0_outputs(1710)) xor (layer0_outputs(7832)));
    outputs(8774) <= not((layer0_outputs(8077)) xor (layer0_outputs(2388)));
    outputs(8775) <= not(layer0_outputs(6328));
    outputs(8776) <= not(layer0_outputs(9378)) or (layer0_outputs(647));
    outputs(8777) <= (layer0_outputs(4034)) xor (layer0_outputs(4933));
    outputs(8778) <= (layer0_outputs(6591)) and not (layer0_outputs(3135));
    outputs(8779) <= not((layer0_outputs(2968)) or (layer0_outputs(8564)));
    outputs(8780) <= layer0_outputs(9273);
    outputs(8781) <= layer0_outputs(9439);
    outputs(8782) <= not(layer0_outputs(7355));
    outputs(8783) <= (layer0_outputs(7108)) and not (layer0_outputs(2342));
    outputs(8784) <= (layer0_outputs(4137)) xor (layer0_outputs(216));
    outputs(8785) <= not(layer0_outputs(7949)) or (layer0_outputs(7219));
    outputs(8786) <= not(layer0_outputs(4012)) or (layer0_outputs(7207));
    outputs(8787) <= layer0_outputs(2400);
    outputs(8788) <= not((layer0_outputs(1866)) xor (layer0_outputs(4882)));
    outputs(8789) <= (layer0_outputs(3784)) and (layer0_outputs(5283));
    outputs(8790) <= (layer0_outputs(9302)) xor (layer0_outputs(2756));
    outputs(8791) <= not((layer0_outputs(1909)) xor (layer0_outputs(3032)));
    outputs(8792) <= (layer0_outputs(8646)) and not (layer0_outputs(1323));
    outputs(8793) <= (layer0_outputs(6435)) or (layer0_outputs(9002));
    outputs(8794) <= not(layer0_outputs(5750));
    outputs(8795) <= layer0_outputs(8286);
    outputs(8796) <= not((layer0_outputs(6273)) xor (layer0_outputs(4823)));
    outputs(8797) <= not((layer0_outputs(8201)) xor (layer0_outputs(1520)));
    outputs(8798) <= (layer0_outputs(3606)) xor (layer0_outputs(6830));
    outputs(8799) <= (layer0_outputs(4314)) xor (layer0_outputs(3018));
    outputs(8800) <= not((layer0_outputs(1286)) xor (layer0_outputs(85)));
    outputs(8801) <= layer0_outputs(5650);
    outputs(8802) <= layer0_outputs(5241);
    outputs(8803) <= (layer0_outputs(5094)) or (layer0_outputs(618));
    outputs(8804) <= not(layer0_outputs(7213));
    outputs(8805) <= layer0_outputs(5732);
    outputs(8806) <= not(layer0_outputs(2533)) or (layer0_outputs(10019));
    outputs(8807) <= not((layer0_outputs(1676)) xor (layer0_outputs(1222)));
    outputs(8808) <= (layer0_outputs(7138)) xor (layer0_outputs(3094));
    outputs(8809) <= not(layer0_outputs(6019));
    outputs(8810) <= not(layer0_outputs(393)) or (layer0_outputs(9807));
    outputs(8811) <= not(layer0_outputs(1166));
    outputs(8812) <= not(layer0_outputs(3143));
    outputs(8813) <= not((layer0_outputs(3768)) and (layer0_outputs(2865)));
    outputs(8814) <= (layer0_outputs(8776)) and (layer0_outputs(4962));
    outputs(8815) <= (layer0_outputs(8281)) or (layer0_outputs(5914));
    outputs(8816) <= (layer0_outputs(3906)) and not (layer0_outputs(2755));
    outputs(8817) <= layer0_outputs(1886);
    outputs(8818) <= not((layer0_outputs(9491)) xor (layer0_outputs(2685)));
    outputs(8819) <= not(layer0_outputs(1209));
    outputs(8820) <= (layer0_outputs(515)) xor (layer0_outputs(5642));
    outputs(8821) <= not(layer0_outputs(5791)) or (layer0_outputs(7140));
    outputs(8822) <= (layer0_outputs(6912)) xor (layer0_outputs(7038));
    outputs(8823) <= (layer0_outputs(7111)) xor (layer0_outputs(7374));
    outputs(8824) <= layer0_outputs(3263);
    outputs(8825) <= (layer0_outputs(2574)) xor (layer0_outputs(8974));
    outputs(8826) <= layer0_outputs(4570);
    outputs(8827) <= (layer0_outputs(4168)) xor (layer0_outputs(5716));
    outputs(8828) <= not((layer0_outputs(5818)) xor (layer0_outputs(9926)));
    outputs(8829) <= layer0_outputs(2955);
    outputs(8830) <= not(layer0_outputs(7126)) or (layer0_outputs(6577));
    outputs(8831) <= not(layer0_outputs(8210));
    outputs(8832) <= layer0_outputs(9683);
    outputs(8833) <= not(layer0_outputs(2640)) or (layer0_outputs(1964));
    outputs(8834) <= not(layer0_outputs(3792)) or (layer0_outputs(2487));
    outputs(8835) <= (layer0_outputs(6571)) xor (layer0_outputs(8386));
    outputs(8836) <= (layer0_outputs(3919)) xor (layer0_outputs(7));
    outputs(8837) <= (layer0_outputs(8794)) or (layer0_outputs(8812));
    outputs(8838) <= not((layer0_outputs(823)) xor (layer0_outputs(4392)));
    outputs(8839) <= not(layer0_outputs(6946));
    outputs(8840) <= layer0_outputs(3471);
    outputs(8841) <= (layer0_outputs(957)) xor (layer0_outputs(3709));
    outputs(8842) <= (layer0_outputs(5617)) xor (layer0_outputs(6060));
    outputs(8843) <= not(layer0_outputs(3777));
    outputs(8844) <= not(layer0_outputs(6353));
    outputs(8845) <= not(layer0_outputs(6393)) or (layer0_outputs(3540));
    outputs(8846) <= not(layer0_outputs(1614));
    outputs(8847) <= not((layer0_outputs(1271)) xor (layer0_outputs(9359)));
    outputs(8848) <= layer0_outputs(1628);
    outputs(8849) <= (layer0_outputs(7052)) and not (layer0_outputs(3584));
    outputs(8850) <= layer0_outputs(7480);
    outputs(8851) <= layer0_outputs(9552);
    outputs(8852) <= (layer0_outputs(9347)) and (layer0_outputs(8604));
    outputs(8853) <= (layer0_outputs(4715)) xor (layer0_outputs(4155));
    outputs(8854) <= not(layer0_outputs(458));
    outputs(8855) <= layer0_outputs(5364);
    outputs(8856) <= layer0_outputs(7684);
    outputs(8857) <= not(layer0_outputs(1965));
    outputs(8858) <= not((layer0_outputs(114)) xor (layer0_outputs(7221)));
    outputs(8859) <= not(layer0_outputs(3961)) or (layer0_outputs(332));
    outputs(8860) <= not(layer0_outputs(2993));
    outputs(8861) <= not(layer0_outputs(2115));
    outputs(8862) <= not((layer0_outputs(3484)) and (layer0_outputs(2912)));
    outputs(8863) <= not(layer0_outputs(4761));
    outputs(8864) <= layer0_outputs(1222);
    outputs(8865) <= (layer0_outputs(7527)) or (layer0_outputs(7540));
    outputs(8866) <= layer0_outputs(3691);
    outputs(8867) <= (layer0_outputs(7462)) xor (layer0_outputs(2305));
    outputs(8868) <= not(layer0_outputs(1308)) or (layer0_outputs(5006));
    outputs(8869) <= (layer0_outputs(2471)) xor (layer0_outputs(7982));
    outputs(8870) <= (layer0_outputs(8517)) xor (layer0_outputs(1621));
    outputs(8871) <= not(layer0_outputs(480));
    outputs(8872) <= not(layer0_outputs(2837));
    outputs(8873) <= (layer0_outputs(7255)) and (layer0_outputs(6855));
    outputs(8874) <= (layer0_outputs(1533)) xor (layer0_outputs(1474));
    outputs(8875) <= not(layer0_outputs(5102));
    outputs(8876) <= not((layer0_outputs(388)) xor (layer0_outputs(1708)));
    outputs(8877) <= (layer0_outputs(3727)) xor (layer0_outputs(2443));
    outputs(8878) <= not(layer0_outputs(8347));
    outputs(8879) <= layer0_outputs(6653);
    outputs(8880) <= not((layer0_outputs(3933)) xor (layer0_outputs(3126)));
    outputs(8881) <= not((layer0_outputs(9841)) and (layer0_outputs(7634)));
    outputs(8882) <= not(layer0_outputs(4108));
    outputs(8883) <= not((layer0_outputs(3594)) xor (layer0_outputs(3222)));
    outputs(8884) <= not(layer0_outputs(164));
    outputs(8885) <= not((layer0_outputs(3409)) xor (layer0_outputs(5238)));
    outputs(8886) <= not((layer0_outputs(5113)) xor (layer0_outputs(8981)));
    outputs(8887) <= not((layer0_outputs(3329)) xor (layer0_outputs(1545)));
    outputs(8888) <= not(layer0_outputs(6604));
    outputs(8889) <= not((layer0_outputs(6561)) or (layer0_outputs(890)));
    outputs(8890) <= layer0_outputs(8187);
    outputs(8891) <= (layer0_outputs(8268)) xor (layer0_outputs(4158));
    outputs(8892) <= (layer0_outputs(7454)) and not (layer0_outputs(4062));
    outputs(8893) <= not(layer0_outputs(511)) or (layer0_outputs(5899));
    outputs(8894) <= not((layer0_outputs(7112)) and (layer0_outputs(5360)));
    outputs(8895) <= layer0_outputs(1921);
    outputs(8896) <= not(layer0_outputs(4509));
    outputs(8897) <= not(layer0_outputs(9549));
    outputs(8898) <= layer0_outputs(4944);
    outputs(8899) <= not((layer0_outputs(9332)) and (layer0_outputs(1690)));
    outputs(8900) <= not(layer0_outputs(9109));
    outputs(8901) <= (layer0_outputs(4137)) xor (layer0_outputs(1853));
    outputs(8902) <= not(layer0_outputs(9942)) or (layer0_outputs(2768));
    outputs(8903) <= (layer0_outputs(6179)) or (layer0_outputs(4898));
    outputs(8904) <= not(layer0_outputs(8757));
    outputs(8905) <= not(layer0_outputs(8100)) or (layer0_outputs(7900));
    outputs(8906) <= not(layer0_outputs(7132));
    outputs(8907) <= not((layer0_outputs(3257)) xor (layer0_outputs(6641)));
    outputs(8908) <= not((layer0_outputs(3080)) or (layer0_outputs(9854)));
    outputs(8909) <= not(layer0_outputs(248)) or (layer0_outputs(392));
    outputs(8910) <= layer0_outputs(6972);
    outputs(8911) <= (layer0_outputs(6590)) xor (layer0_outputs(3668));
    outputs(8912) <= not((layer0_outputs(1405)) xor (layer0_outputs(2769)));
    outputs(8913) <= not(layer0_outputs(8904)) or (layer0_outputs(3620));
    outputs(8914) <= layer0_outputs(1030);
    outputs(8915) <= not(layer0_outputs(2493));
    outputs(8916) <= not(layer0_outputs(4990));
    outputs(8917) <= not((layer0_outputs(6963)) xor (layer0_outputs(5446)));
    outputs(8918) <= not(layer0_outputs(6040)) or (layer0_outputs(3165));
    outputs(8919) <= not(layer0_outputs(6538));
    outputs(8920) <= not(layer0_outputs(3137)) or (layer0_outputs(2663));
    outputs(8921) <= not((layer0_outputs(836)) xor (layer0_outputs(9123)));
    outputs(8922) <= layer0_outputs(8677);
    outputs(8923) <= layer0_outputs(236);
    outputs(8924) <= not(layer0_outputs(2995));
    outputs(8925) <= (layer0_outputs(9711)) and not (layer0_outputs(7003));
    outputs(8926) <= not((layer0_outputs(8092)) xor (layer0_outputs(8310)));
    outputs(8927) <= (layer0_outputs(9219)) or (layer0_outputs(8370));
    outputs(8928) <= not(layer0_outputs(828));
    outputs(8929) <= not(layer0_outputs(610)) or (layer0_outputs(5793));
    outputs(8930) <= (layer0_outputs(3997)) xor (layer0_outputs(6319));
    outputs(8931) <= not(layer0_outputs(7423)) or (layer0_outputs(8924));
    outputs(8932) <= not((layer0_outputs(8267)) xor (layer0_outputs(9853)));
    outputs(8933) <= (layer0_outputs(6455)) and not (layer0_outputs(3971));
    outputs(8934) <= not(layer0_outputs(5964));
    outputs(8935) <= layer0_outputs(8621);
    outputs(8936) <= (layer0_outputs(9631)) xor (layer0_outputs(5659));
    outputs(8937) <= layer0_outputs(6403);
    outputs(8938) <= not(layer0_outputs(95));
    outputs(8939) <= not(layer0_outputs(2889));
    outputs(8940) <= (layer0_outputs(385)) or (layer0_outputs(881));
    outputs(8941) <= (layer0_outputs(5594)) xor (layer0_outputs(2849));
    outputs(8942) <= (layer0_outputs(8546)) or (layer0_outputs(7604));
    outputs(8943) <= '1';
    outputs(8944) <= (layer0_outputs(944)) and (layer0_outputs(1697));
    outputs(8945) <= layer0_outputs(4041);
    outputs(8946) <= (layer0_outputs(4612)) xor (layer0_outputs(8517));
    outputs(8947) <= not((layer0_outputs(1960)) xor (layer0_outputs(2891)));
    outputs(8948) <= (layer0_outputs(9057)) xor (layer0_outputs(2877));
    outputs(8949) <= layer0_outputs(6958);
    outputs(8950) <= not((layer0_outputs(1803)) xor (layer0_outputs(4471)));
    outputs(8951) <= (layer0_outputs(5331)) and not (layer0_outputs(5992));
    outputs(8952) <= (layer0_outputs(3948)) and (layer0_outputs(2318));
    outputs(8953) <= layer0_outputs(668);
    outputs(8954) <= not(layer0_outputs(6891));
    outputs(8955) <= not(layer0_outputs(10062)) or (layer0_outputs(2015));
    outputs(8956) <= (layer0_outputs(3656)) xor (layer0_outputs(1159));
    outputs(8957) <= not((layer0_outputs(5933)) xor (layer0_outputs(7638)));
    outputs(8958) <= not(layer0_outputs(807));
    outputs(8959) <= (layer0_outputs(168)) and not (layer0_outputs(6841));
    outputs(8960) <= (layer0_outputs(10009)) and not (layer0_outputs(2319));
    outputs(8961) <= not(layer0_outputs(3488));
    outputs(8962) <= not((layer0_outputs(2363)) or (layer0_outputs(8662)));
    outputs(8963) <= not(layer0_outputs(1303));
    outputs(8964) <= (layer0_outputs(5945)) xor (layer0_outputs(1933));
    outputs(8965) <= layer0_outputs(3600);
    outputs(8966) <= (layer0_outputs(3486)) xor (layer0_outputs(581));
    outputs(8967) <= not(layer0_outputs(6983));
    outputs(8968) <= not(layer0_outputs(9064)) or (layer0_outputs(8456));
    outputs(8969) <= (layer0_outputs(166)) xor (layer0_outputs(1204));
    outputs(8970) <= not(layer0_outputs(6452));
    outputs(8971) <= not((layer0_outputs(976)) xor (layer0_outputs(4339)));
    outputs(8972) <= not((layer0_outputs(4015)) and (layer0_outputs(5447)));
    outputs(8973) <= not((layer0_outputs(4424)) and (layer0_outputs(6816)));
    outputs(8974) <= not(layer0_outputs(5498));
    outputs(8975) <= layer0_outputs(4748);
    outputs(8976) <= not((layer0_outputs(7393)) xor (layer0_outputs(2137)));
    outputs(8977) <= layer0_outputs(6172);
    outputs(8978) <= not((layer0_outputs(617)) xor (layer0_outputs(7867)));
    outputs(8979) <= not(layer0_outputs(6386)) or (layer0_outputs(10067));
    outputs(8980) <= (layer0_outputs(3310)) xor (layer0_outputs(1557));
    outputs(8981) <= not(layer0_outputs(2745)) or (layer0_outputs(5267));
    outputs(8982) <= layer0_outputs(5766);
    outputs(8983) <= not(layer0_outputs(9746)) or (layer0_outputs(3872));
    outputs(8984) <= (layer0_outputs(6734)) and (layer0_outputs(2250));
    outputs(8985) <= not(layer0_outputs(2849));
    outputs(8986) <= not(layer0_outputs(2604)) or (layer0_outputs(278));
    outputs(8987) <= not(layer0_outputs(4453));
    outputs(8988) <= not(layer0_outputs(9259));
    outputs(8989) <= not(layer0_outputs(6093));
    outputs(8990) <= not(layer0_outputs(4289));
    outputs(8991) <= layer0_outputs(8060);
    outputs(8992) <= (layer0_outputs(7820)) or (layer0_outputs(5645));
    outputs(8993) <= (layer0_outputs(6893)) xor (layer0_outputs(4781));
    outputs(8994) <= not(layer0_outputs(9448));
    outputs(8995) <= not((layer0_outputs(5251)) or (layer0_outputs(5544)));
    outputs(8996) <= layer0_outputs(1359);
    outputs(8997) <= (layer0_outputs(2760)) xor (layer0_outputs(8848));
    outputs(8998) <= layer0_outputs(7930);
    outputs(8999) <= layer0_outputs(1290);
    outputs(9000) <= (layer0_outputs(4827)) or (layer0_outputs(2014));
    outputs(9001) <= not((layer0_outputs(5735)) xor (layer0_outputs(7525)));
    outputs(9002) <= layer0_outputs(819);
    outputs(9003) <= (layer0_outputs(718)) and (layer0_outputs(7549));
    outputs(9004) <= not((layer0_outputs(5985)) and (layer0_outputs(373)));
    outputs(9005) <= not((layer0_outputs(1621)) and (layer0_outputs(912)));
    outputs(9006) <= '0';
    outputs(9007) <= layer0_outputs(418);
    outputs(9008) <= not(layer0_outputs(3463)) or (layer0_outputs(6316));
    outputs(9009) <= not(layer0_outputs(5787));
    outputs(9010) <= (layer0_outputs(2881)) and (layer0_outputs(4048));
    outputs(9011) <= not(layer0_outputs(3345));
    outputs(9012) <= not((layer0_outputs(2215)) xor (layer0_outputs(1882)));
    outputs(9013) <= not(layer0_outputs(8356));
    outputs(9014) <= not((layer0_outputs(8391)) xor (layer0_outputs(20)));
    outputs(9015) <= not((layer0_outputs(6418)) xor (layer0_outputs(7513)));
    outputs(9016) <= (layer0_outputs(6291)) xor (layer0_outputs(2018));
    outputs(9017) <= not(layer0_outputs(8151)) or (layer0_outputs(7175));
    outputs(9018) <= not(layer0_outputs(6623)) or (layer0_outputs(7457));
    outputs(9019) <= not((layer0_outputs(9652)) and (layer0_outputs(7367)));
    outputs(9020) <= not(layer0_outputs(5470)) or (layer0_outputs(4123));
    outputs(9021) <= not(layer0_outputs(6716)) or (layer0_outputs(190));
    outputs(9022) <= (layer0_outputs(7104)) xor (layer0_outputs(8961));
    outputs(9023) <= layer0_outputs(181);
    outputs(9024) <= layer0_outputs(3778);
    outputs(9025) <= not((layer0_outputs(4478)) and (layer0_outputs(1256)));
    outputs(9026) <= not(layer0_outputs(10084)) or (layer0_outputs(6245));
    outputs(9027) <= not(layer0_outputs(2160)) or (layer0_outputs(2055));
    outputs(9028) <= not(layer0_outputs(59)) or (layer0_outputs(5767));
    outputs(9029) <= not((layer0_outputs(5135)) xor (layer0_outputs(6901)));
    outputs(9030) <= not((layer0_outputs(6103)) xor (layer0_outputs(650)));
    outputs(9031) <= not((layer0_outputs(1791)) xor (layer0_outputs(3968)));
    outputs(9032) <= not(layer0_outputs(7049));
    outputs(9033) <= not((layer0_outputs(5776)) xor (layer0_outputs(523)));
    outputs(9034) <= not(layer0_outputs(7627));
    outputs(9035) <= layer0_outputs(7735);
    outputs(9036) <= not(layer0_outputs(4525));
    outputs(9037) <= (layer0_outputs(4406)) and (layer0_outputs(918));
    outputs(9038) <= (layer0_outputs(5070)) and (layer0_outputs(7283));
    outputs(9039) <= layer0_outputs(7162);
    outputs(9040) <= layer0_outputs(2200);
    outputs(9041) <= '0';
    outputs(9042) <= not(layer0_outputs(3012));
    outputs(9043) <= '0';
    outputs(9044) <= (layer0_outputs(3157)) xor (layer0_outputs(5357));
    outputs(9045) <= not((layer0_outputs(6209)) xor (layer0_outputs(5017)));
    outputs(9046) <= not((layer0_outputs(879)) and (layer0_outputs(493)));
    outputs(9047) <= layer0_outputs(357);
    outputs(9048) <= (layer0_outputs(2412)) xor (layer0_outputs(5759));
    outputs(9049) <= not(layer0_outputs(3283));
    outputs(9050) <= not((layer0_outputs(5126)) xor (layer0_outputs(9940)));
    outputs(9051) <= layer0_outputs(4098);
    outputs(9052) <= not(layer0_outputs(9867));
    outputs(9053) <= not(layer0_outputs(2095));
    outputs(9054) <= (layer0_outputs(5299)) xor (layer0_outputs(6994));
    outputs(9055) <= layer0_outputs(9137);
    outputs(9056) <= (layer0_outputs(5761)) and not (layer0_outputs(2271));
    outputs(9057) <= not(layer0_outputs(6779));
    outputs(9058) <= not((layer0_outputs(7268)) xor (layer0_outputs(10128)));
    outputs(9059) <= (layer0_outputs(4838)) xor (layer0_outputs(5507));
    outputs(9060) <= not(layer0_outputs(3125));
    outputs(9061) <= layer0_outputs(1462);
    outputs(9062) <= not(layer0_outputs(1831));
    outputs(9063) <= layer0_outputs(5005);
    outputs(9064) <= not(layer0_outputs(4743));
    outputs(9065) <= (layer0_outputs(5514)) and not (layer0_outputs(4260));
    outputs(9066) <= not(layer0_outputs(9676)) or (layer0_outputs(4907));
    outputs(9067) <= not((layer0_outputs(1203)) xor (layer0_outputs(9734)));
    outputs(9068) <= '1';
    outputs(9069) <= not(layer0_outputs(9409));
    outputs(9070) <= '1';
    outputs(9071) <= layer0_outputs(6796);
    outputs(9072) <= layer0_outputs(591);
    outputs(9073) <= layer0_outputs(7726);
    outputs(9074) <= not((layer0_outputs(4141)) xor (layer0_outputs(2151)));
    outputs(9075) <= not((layer0_outputs(1760)) xor (layer0_outputs(4915)));
    outputs(9076) <= layer0_outputs(757);
    outputs(9077) <= not(layer0_outputs(7666)) or (layer0_outputs(8394));
    outputs(9078) <= not((layer0_outputs(6666)) xor (layer0_outputs(3917)));
    outputs(9079) <= (layer0_outputs(5552)) xor (layer0_outputs(298));
    outputs(9080) <= (layer0_outputs(1231)) and not (layer0_outputs(3102));
    outputs(9081) <= not((layer0_outputs(5735)) and (layer0_outputs(4099)));
    outputs(9082) <= not(layer0_outputs(3715));
    outputs(9083) <= (layer0_outputs(2024)) xor (layer0_outputs(937));
    outputs(9084) <= not(layer0_outputs(7173)) or (layer0_outputs(4431));
    outputs(9085) <= not(layer0_outputs(6802));
    outputs(9086) <= (layer0_outputs(1342)) or (layer0_outputs(8884));
    outputs(9087) <= not(layer0_outputs(1482));
    outputs(9088) <= not(layer0_outputs(7612)) or (layer0_outputs(950));
    outputs(9089) <= (layer0_outputs(4769)) xor (layer0_outputs(9215));
    outputs(9090) <= not((layer0_outputs(2255)) xor (layer0_outputs(6850)));
    outputs(9091) <= not((layer0_outputs(5079)) xor (layer0_outputs(2850)));
    outputs(9092) <= not((layer0_outputs(7307)) xor (layer0_outputs(2908)));
    outputs(9093) <= layer0_outputs(5062);
    outputs(9094) <= not(layer0_outputs(6637)) or (layer0_outputs(10059));
    outputs(9095) <= (layer0_outputs(84)) xor (layer0_outputs(5237));
    outputs(9096) <= not(layer0_outputs(7049));
    outputs(9097) <= not(layer0_outputs(7622));
    outputs(9098) <= (layer0_outputs(5817)) and not (layer0_outputs(4217));
    outputs(9099) <= not((layer0_outputs(3701)) xor (layer0_outputs(2697)));
    outputs(9100) <= layer0_outputs(5698);
    outputs(9101) <= not((layer0_outputs(9281)) xor (layer0_outputs(4221)));
    outputs(9102) <= (layer0_outputs(9727)) xor (layer0_outputs(4780));
    outputs(9103) <= not((layer0_outputs(9103)) xor (layer0_outputs(4592)));
    outputs(9104) <= (layer0_outputs(350)) and not (layer0_outputs(8487));
    outputs(9105) <= (layer0_outputs(1040)) xor (layer0_outputs(5647));
    outputs(9106) <= not(layer0_outputs(4398));
    outputs(9107) <= not(layer0_outputs(1594)) or (layer0_outputs(4531));
    outputs(9108) <= layer0_outputs(3734);
    outputs(9109) <= (layer0_outputs(3992)) and not (layer0_outputs(185));
    outputs(9110) <= (layer0_outputs(697)) and (layer0_outputs(7246));
    outputs(9111) <= not(layer0_outputs(715));
    outputs(9112) <= layer0_outputs(5763);
    outputs(9113) <= not((layer0_outputs(3850)) and (layer0_outputs(9126)));
    outputs(9114) <= (layer0_outputs(1063)) xor (layer0_outputs(38));
    outputs(9115) <= '1';
    outputs(9116) <= layer0_outputs(5909);
    outputs(9117) <= (layer0_outputs(6990)) xor (layer0_outputs(9872));
    outputs(9118) <= not((layer0_outputs(9204)) xor (layer0_outputs(7333)));
    outputs(9119) <= (layer0_outputs(4006)) xor (layer0_outputs(3761));
    outputs(9120) <= layer0_outputs(7055);
    outputs(9121) <= (layer0_outputs(5200)) xor (layer0_outputs(7535));
    outputs(9122) <= layer0_outputs(5503);
    outputs(9123) <= not((layer0_outputs(5779)) xor (layer0_outputs(6760)));
    outputs(9124) <= not(layer0_outputs(8647));
    outputs(9125) <= not(layer0_outputs(6894));
    outputs(9126) <= not(layer0_outputs(6101));
    outputs(9127) <= not(layer0_outputs(9412));
    outputs(9128) <= not(layer0_outputs(1935));
    outputs(9129) <= (layer0_outputs(1486)) or (layer0_outputs(6532));
    outputs(9130) <= layer0_outputs(7300);
    outputs(9131) <= (layer0_outputs(3417)) xor (layer0_outputs(2635));
    outputs(9132) <= layer0_outputs(9567);
    outputs(9133) <= not((layer0_outputs(9607)) or (layer0_outputs(3928)));
    outputs(9134) <= not(layer0_outputs(1511));
    outputs(9135) <= not((layer0_outputs(4066)) and (layer0_outputs(2386)));
    outputs(9136) <= layer0_outputs(5004);
    outputs(9137) <= layer0_outputs(7991);
    outputs(9138) <= not(layer0_outputs(9086));
    outputs(9139) <= not((layer0_outputs(1783)) xor (layer0_outputs(9158)));
    outputs(9140) <= not(layer0_outputs(840)) or (layer0_outputs(5838));
    outputs(9141) <= not(layer0_outputs(2334));
    outputs(9142) <= not((layer0_outputs(6923)) xor (layer0_outputs(4504)));
    outputs(9143) <= layer0_outputs(5347);
    outputs(9144) <= (layer0_outputs(5903)) or (layer0_outputs(5414));
    outputs(9145) <= not((layer0_outputs(8496)) or (layer0_outputs(1113)));
    outputs(9146) <= (layer0_outputs(5968)) or (layer0_outputs(9674));
    outputs(9147) <= layer0_outputs(5793);
    outputs(9148) <= not((layer0_outputs(9081)) xor (layer0_outputs(2397)));
    outputs(9149) <= not(layer0_outputs(9311));
    outputs(9150) <= not((layer0_outputs(8498)) xor (layer0_outputs(4468)));
    outputs(9151) <= not((layer0_outputs(8535)) xor (layer0_outputs(769)));
    outputs(9152) <= (layer0_outputs(2997)) or (layer0_outputs(4304));
    outputs(9153) <= not(layer0_outputs(830));
    outputs(9154) <= not(layer0_outputs(7545));
    outputs(9155) <= layer0_outputs(6298);
    outputs(9156) <= (layer0_outputs(8799)) and not (layer0_outputs(4849));
    outputs(9157) <= not(layer0_outputs(5166));
    outputs(9158) <= not((layer0_outputs(5627)) xor (layer0_outputs(1561)));
    outputs(9159) <= not(layer0_outputs(3746));
    outputs(9160) <= not((layer0_outputs(8333)) xor (layer0_outputs(2717)));
    outputs(9161) <= not(layer0_outputs(8249));
    outputs(9162) <= not((layer0_outputs(3019)) xor (layer0_outputs(8031)));
    outputs(9163) <= (layer0_outputs(4602)) xor (layer0_outputs(8458));
    outputs(9164) <= not((layer0_outputs(5091)) or (layer0_outputs(3987)));
    outputs(9165) <= layer0_outputs(5483);
    outputs(9166) <= not((layer0_outputs(1447)) and (layer0_outputs(9485)));
    outputs(9167) <= not(layer0_outputs(4503));
    outputs(9168) <= (layer0_outputs(6156)) xor (layer0_outputs(7566));
    outputs(9169) <= not((layer0_outputs(5107)) xor (layer0_outputs(9313)));
    outputs(9170) <= not(layer0_outputs(2572));
    outputs(9171) <= not((layer0_outputs(151)) xor (layer0_outputs(5292)));
    outputs(9172) <= not(layer0_outputs(703));
    outputs(9173) <= not(layer0_outputs(5738)) or (layer0_outputs(9257));
    outputs(9174) <= not(layer0_outputs(4584));
    outputs(9175) <= not(layer0_outputs(8388));
    outputs(9176) <= not(layer0_outputs(2478));
    outputs(9177) <= layer0_outputs(4074);
    outputs(9178) <= layer0_outputs(9508);
    outputs(9179) <= layer0_outputs(2706);
    outputs(9180) <= not((layer0_outputs(6711)) xor (layer0_outputs(3519)));
    outputs(9181) <= not(layer0_outputs(1761));
    outputs(9182) <= not((layer0_outputs(162)) xor (layer0_outputs(4706)));
    outputs(9183) <= (layer0_outputs(1514)) and (layer0_outputs(9553));
    outputs(9184) <= (layer0_outputs(7863)) xor (layer0_outputs(9522));
    outputs(9185) <= (layer0_outputs(5369)) and (layer0_outputs(1333));
    outputs(9186) <= (layer0_outputs(3198)) and (layer0_outputs(9113));
    outputs(9187) <= not((layer0_outputs(7934)) xor (layer0_outputs(10222)));
    outputs(9188) <= (layer0_outputs(607)) xor (layer0_outputs(2404));
    outputs(9189) <= (layer0_outputs(80)) xor (layer0_outputs(2640));
    outputs(9190) <= not(layer0_outputs(9392));
    outputs(9191) <= layer0_outputs(1401);
    outputs(9192) <= not((layer0_outputs(2529)) xor (layer0_outputs(9107)));
    outputs(9193) <= not(layer0_outputs(4808));
    outputs(9194) <= not(layer0_outputs(6224));
    outputs(9195) <= not(layer0_outputs(7513)) or (layer0_outputs(993));
    outputs(9196) <= not((layer0_outputs(5716)) xor (layer0_outputs(8739)));
    outputs(9197) <= not(layer0_outputs(5730));
    outputs(9198) <= layer0_outputs(4946);
    outputs(9199) <= layer0_outputs(7946);
    outputs(9200) <= (layer0_outputs(5002)) xor (layer0_outputs(1883));
    outputs(9201) <= layer0_outputs(7059);
    outputs(9202) <= not(layer0_outputs(9702)) or (layer0_outputs(8040));
    outputs(9203) <= layer0_outputs(2976);
    outputs(9204) <= not((layer0_outputs(7500)) and (layer0_outputs(9996)));
    outputs(9205) <= layer0_outputs(8990);
    outputs(9206) <= not(layer0_outputs(3724));
    outputs(9207) <= layer0_outputs(1444);
    outputs(9208) <= not(layer0_outputs(10111));
    outputs(9209) <= (layer0_outputs(3454)) xor (layer0_outputs(7876));
    outputs(9210) <= not(layer0_outputs(7959));
    outputs(9211) <= not(layer0_outputs(515)) or (layer0_outputs(7332));
    outputs(9212) <= not(layer0_outputs(4345));
    outputs(9213) <= layer0_outputs(10236);
    outputs(9214) <= (layer0_outputs(9108)) xor (layer0_outputs(9574));
    outputs(9215) <= not((layer0_outputs(9508)) xor (layer0_outputs(8886)));
    outputs(9216) <= not(layer0_outputs(3943)) or (layer0_outputs(5211));
    outputs(9217) <= (layer0_outputs(9222)) and not (layer0_outputs(6287));
    outputs(9218) <= (layer0_outputs(7544)) and not (layer0_outputs(5693));
    outputs(9219) <= not(layer0_outputs(1913));
    outputs(9220) <= (layer0_outputs(1604)) and not (layer0_outputs(2210));
    outputs(9221) <= layer0_outputs(6218);
    outputs(9222) <= layer0_outputs(8797);
    outputs(9223) <= not(layer0_outputs(6569));
    outputs(9224) <= (layer0_outputs(9855)) and not (layer0_outputs(3418));
    outputs(9225) <= (layer0_outputs(3678)) or (layer0_outputs(8911));
    outputs(9226) <= not((layer0_outputs(5531)) and (layer0_outputs(505)));
    outputs(9227) <= not(layer0_outputs(6542));
    outputs(9228) <= layer0_outputs(9128);
    outputs(9229) <= layer0_outputs(9968);
    outputs(9230) <= not((layer0_outputs(3503)) xor (layer0_outputs(7850)));
    outputs(9231) <= (layer0_outputs(2738)) xor (layer0_outputs(807));
    outputs(9232) <= (layer0_outputs(4016)) and not (layer0_outputs(2417));
    outputs(9233) <= layer0_outputs(4938);
    outputs(9234) <= not(layer0_outputs(6029));
    outputs(9235) <= layer0_outputs(477);
    outputs(9236) <= not((layer0_outputs(8840)) xor (layer0_outputs(5458)));
    outputs(9237) <= not((layer0_outputs(9309)) xor (layer0_outputs(4730)));
    outputs(9238) <= not(layer0_outputs(4408));
    outputs(9239) <= layer0_outputs(9141);
    outputs(9240) <= not(layer0_outputs(3141));
    outputs(9241) <= not((layer0_outputs(3775)) or (layer0_outputs(8756)));
    outputs(9242) <= not(layer0_outputs(7716));
    outputs(9243) <= (layer0_outputs(1619)) xor (layer0_outputs(8321));
    outputs(9244) <= not((layer0_outputs(2134)) and (layer0_outputs(1146)));
    outputs(9245) <= (layer0_outputs(877)) xor (layer0_outputs(6301));
    outputs(9246) <= not(layer0_outputs(9390));
    outputs(9247) <= layer0_outputs(5825);
    outputs(9248) <= not(layer0_outputs(7782));
    outputs(9249) <= layer0_outputs(9072);
    outputs(9250) <= layer0_outputs(6039);
    outputs(9251) <= not(layer0_outputs(9789));
    outputs(9252) <= not((layer0_outputs(2039)) xor (layer0_outputs(4089)));
    outputs(9253) <= (layer0_outputs(3251)) and not (layer0_outputs(9254));
    outputs(9254) <= not((layer0_outputs(5976)) xor (layer0_outputs(3300)));
    outputs(9255) <= not((layer0_outputs(4821)) xor (layer0_outputs(6381)));
    outputs(9256) <= (layer0_outputs(8717)) and not (layer0_outputs(1554));
    outputs(9257) <= not((layer0_outputs(8035)) xor (layer0_outputs(4832)));
    outputs(9258) <= (layer0_outputs(604)) and (layer0_outputs(3765));
    outputs(9259) <= layer0_outputs(2858);
    outputs(9260) <= not(layer0_outputs(6872));
    outputs(9261) <= not(layer0_outputs(9837));
    outputs(9262) <= not(layer0_outputs(3132));
    outputs(9263) <= layer0_outputs(222);
    outputs(9264) <= (layer0_outputs(4057)) and not (layer0_outputs(4818));
    outputs(9265) <= (layer0_outputs(424)) and not (layer0_outputs(3822));
    outputs(9266) <= (layer0_outputs(2953)) and not (layer0_outputs(4587));
    outputs(9267) <= layer0_outputs(3225);
    outputs(9268) <= (layer0_outputs(3001)) xor (layer0_outputs(7519));
    outputs(9269) <= layer0_outputs(2747);
    outputs(9270) <= (layer0_outputs(2045)) and (layer0_outputs(2838));
    outputs(9271) <= layer0_outputs(9831);
    outputs(9272) <= not((layer0_outputs(801)) xor (layer0_outputs(2601)));
    outputs(9273) <= not((layer0_outputs(4467)) xor (layer0_outputs(7754)));
    outputs(9274) <= not(layer0_outputs(1480));
    outputs(9275) <= not(layer0_outputs(3482));
    outputs(9276) <= not(layer0_outputs(3118));
    outputs(9277) <= (layer0_outputs(3521)) xor (layer0_outputs(1761));
    outputs(9278) <= (layer0_outputs(6859)) xor (layer0_outputs(5854));
    outputs(9279) <= not(layer0_outputs(7635));
    outputs(9280) <= not(layer0_outputs(843));
    outputs(9281) <= not(layer0_outputs(9949));
    outputs(9282) <= (layer0_outputs(8203)) and (layer0_outputs(5903));
    outputs(9283) <= (layer0_outputs(7398)) and not (layer0_outputs(8343));
    outputs(9284) <= not(layer0_outputs(2330));
    outputs(9285) <= (layer0_outputs(8623)) and not (layer0_outputs(7116));
    outputs(9286) <= not(layer0_outputs(4083));
    outputs(9287) <= not(layer0_outputs(10170)) or (layer0_outputs(1148));
    outputs(9288) <= not((layer0_outputs(3646)) xor (layer0_outputs(3363)));
    outputs(9289) <= layer0_outputs(5981);
    outputs(9290) <= (layer0_outputs(9082)) and not (layer0_outputs(7042));
    outputs(9291) <= not(layer0_outputs(3643));
    outputs(9292) <= (layer0_outputs(4281)) xor (layer0_outputs(2163));
    outputs(9293) <= not((layer0_outputs(4874)) or (layer0_outputs(6618)));
    outputs(9294) <= (layer0_outputs(55)) and (layer0_outputs(2193));
    outputs(9295) <= (layer0_outputs(5966)) and (layer0_outputs(3291));
    outputs(9296) <= not(layer0_outputs(8369));
    outputs(9297) <= layer0_outputs(7131);
    outputs(9298) <= layer0_outputs(8450);
    outputs(9299) <= not(layer0_outputs(534));
    outputs(9300) <= (layer0_outputs(4231)) or (layer0_outputs(383));
    outputs(9301) <= layer0_outputs(5865);
    outputs(9302) <= not(layer0_outputs(1550));
    outputs(9303) <= (layer0_outputs(3924)) xor (layer0_outputs(8717));
    outputs(9304) <= not(layer0_outputs(7848));
    outputs(9305) <= not(layer0_outputs(1642));
    outputs(9306) <= (layer0_outputs(3280)) xor (layer0_outputs(6022));
    outputs(9307) <= (layer0_outputs(10210)) xor (layer0_outputs(2126));
    outputs(9308) <= layer0_outputs(4149);
    outputs(9309) <= layer0_outputs(8043);
    outputs(9310) <= not(layer0_outputs(9526));
    outputs(9311) <= not(layer0_outputs(6477));
    outputs(9312) <= (layer0_outputs(1319)) and (layer0_outputs(10122));
    outputs(9313) <= (layer0_outputs(9055)) and not (layer0_outputs(9600));
    outputs(9314) <= not(layer0_outputs(6109));
    outputs(9315) <= layer0_outputs(2131);
    outputs(9316) <= layer0_outputs(1102);
    outputs(9317) <= not((layer0_outputs(1361)) or (layer0_outputs(1636)));
    outputs(9318) <= (layer0_outputs(7931)) xor (layer0_outputs(1358));
    outputs(9319) <= layer0_outputs(5663);
    outputs(9320) <= (layer0_outputs(5994)) xor (layer0_outputs(6969));
    outputs(9321) <= layer0_outputs(6681);
    outputs(9322) <= not(layer0_outputs(9927));
    outputs(9323) <= (layer0_outputs(7961)) and not (layer0_outputs(2703));
    outputs(9324) <= layer0_outputs(5584);
    outputs(9325) <= not(layer0_outputs(7036));
    outputs(9326) <= layer0_outputs(1623);
    outputs(9327) <= not((layer0_outputs(9866)) or (layer0_outputs(1268)));
    outputs(9328) <= layer0_outputs(1673);
    outputs(9329) <= not((layer0_outputs(9857)) or (layer0_outputs(1283)));
    outputs(9330) <= not(layer0_outputs(8952));
    outputs(9331) <= layer0_outputs(7779);
    outputs(9332) <= not((layer0_outputs(2507)) xor (layer0_outputs(4306)));
    outputs(9333) <= not((layer0_outputs(1977)) and (layer0_outputs(1280)));
    outputs(9334) <= (layer0_outputs(3708)) and not (layer0_outputs(2274));
    outputs(9335) <= not(layer0_outputs(1584));
    outputs(9336) <= not((layer0_outputs(9161)) xor (layer0_outputs(4811)));
    outputs(9337) <= not(layer0_outputs(7001)) or (layer0_outputs(7030));
    outputs(9338) <= (layer0_outputs(5396)) and not (layer0_outputs(4530));
    outputs(9339) <= not((layer0_outputs(3097)) or (layer0_outputs(8973)));
    outputs(9340) <= not(layer0_outputs(1281));
    outputs(9341) <= not(layer0_outputs(1800));
    outputs(9342) <= (layer0_outputs(7613)) and not (layer0_outputs(6010));
    outputs(9343) <= not(layer0_outputs(6579));
    outputs(9344) <= (layer0_outputs(1212)) and not (layer0_outputs(5695));
    outputs(9345) <= not(layer0_outputs(9639));
    outputs(9346) <= not(layer0_outputs(8556));
    outputs(9347) <= not(layer0_outputs(6853));
    outputs(9348) <= (layer0_outputs(3077)) xor (layer0_outputs(8568));
    outputs(9349) <= (layer0_outputs(3361)) and not (layer0_outputs(8427));
    outputs(9350) <= layer0_outputs(8989);
    outputs(9351) <= (layer0_outputs(9690)) and not (layer0_outputs(4027));
    outputs(9352) <= not((layer0_outputs(6890)) or (layer0_outputs(1750)));
    outputs(9353) <= layer0_outputs(4736);
    outputs(9354) <= layer0_outputs(4801);
    outputs(9355) <= (layer0_outputs(1762)) and not (layer0_outputs(6515));
    outputs(9356) <= (layer0_outputs(4771)) and (layer0_outputs(115));
    outputs(9357) <= (layer0_outputs(3304)) and not (layer0_outputs(2279));
    outputs(9358) <= not(layer0_outputs(8958));
    outputs(9359) <= (layer0_outputs(6444)) and not (layer0_outputs(1367));
    outputs(9360) <= layer0_outputs(5717);
    outputs(9361) <= not(layer0_outputs(4761));
    outputs(9362) <= layer0_outputs(5009);
    outputs(9363) <= not(layer0_outputs(7310));
    outputs(9364) <= not(layer0_outputs(4246));
    outputs(9365) <= not(layer0_outputs(1295));
    outputs(9366) <= not((layer0_outputs(8993)) xor (layer0_outputs(9634)));
    outputs(9367) <= not((layer0_outputs(2016)) or (layer0_outputs(3539)));
    outputs(9368) <= (layer0_outputs(6583)) xor (layer0_outputs(7037));
    outputs(9369) <= not((layer0_outputs(4949)) xor (layer0_outputs(2275)));
    outputs(9370) <= not(layer0_outputs(689));
    outputs(9371) <= (layer0_outputs(2251)) and not (layer0_outputs(7333));
    outputs(9372) <= not((layer0_outputs(5600)) or (layer0_outputs(8239)));
    outputs(9373) <= (layer0_outputs(8826)) and not (layer0_outputs(9163));
    outputs(9374) <= layer0_outputs(5441);
    outputs(9375) <= layer0_outputs(8177);
    outputs(9376) <= layer0_outputs(6111);
    outputs(9377) <= (layer0_outputs(1682)) and (layer0_outputs(46));
    outputs(9378) <= not(layer0_outputs(9789));
    outputs(9379) <= layer0_outputs(6218);
    outputs(9380) <= not((layer0_outputs(3175)) or (layer0_outputs(2875)));
    outputs(9381) <= layer0_outputs(1445);
    outputs(9382) <= (layer0_outputs(513)) and not (layer0_outputs(5192));
    outputs(9383) <= (layer0_outputs(9934)) and not (layer0_outputs(7153));
    outputs(9384) <= (layer0_outputs(6028)) and (layer0_outputs(7870));
    outputs(9385) <= not(layer0_outputs(5477));
    outputs(9386) <= (layer0_outputs(8196)) and (layer0_outputs(4507));
    outputs(9387) <= not((layer0_outputs(1073)) and (layer0_outputs(6964)));
    outputs(9388) <= not(layer0_outputs(9122));
    outputs(9389) <= (layer0_outputs(678)) xor (layer0_outputs(9568));
    outputs(9390) <= (layer0_outputs(9175)) xor (layer0_outputs(733));
    outputs(9391) <= not((layer0_outputs(467)) xor (layer0_outputs(1325)));
    outputs(9392) <= (layer0_outputs(4513)) and not (layer0_outputs(3952));
    outputs(9393) <= (layer0_outputs(2205)) and not (layer0_outputs(6942));
    outputs(9394) <= (layer0_outputs(2047)) xor (layer0_outputs(1318));
    outputs(9395) <= not((layer0_outputs(301)) xor (layer0_outputs(576)));
    outputs(9396) <= not((layer0_outputs(5538)) xor (layer0_outputs(1619)));
    outputs(9397) <= not((layer0_outputs(6095)) xor (layer0_outputs(6416)));
    outputs(9398) <= layer0_outputs(7147);
    outputs(9399) <= not((layer0_outputs(1685)) or (layer0_outputs(5132)));
    outputs(9400) <= layer0_outputs(8442);
    outputs(9401) <= (layer0_outputs(5497)) xor (layer0_outputs(958));
    outputs(9402) <= layer0_outputs(2349);
    outputs(9403) <= (layer0_outputs(2736)) and not (layer0_outputs(4710));
    outputs(9404) <= layer0_outputs(4439);
    outputs(9405) <= not(layer0_outputs(9379));
    outputs(9406) <= layer0_outputs(8251);
    outputs(9407) <= not(layer0_outputs(862));
    outputs(9408) <= not((layer0_outputs(3307)) xor (layer0_outputs(4830)));
    outputs(9409) <= not(layer0_outputs(2312));
    outputs(9410) <= not((layer0_outputs(9664)) xor (layer0_outputs(2080)));
    outputs(9411) <= layer0_outputs(6535);
    outputs(9412) <= not(layer0_outputs(1742));
    outputs(9413) <= layer0_outputs(2209);
    outputs(9414) <= not(layer0_outputs(9020));
    outputs(9415) <= layer0_outputs(705);
    outputs(9416) <= not(layer0_outputs(2929));
    outputs(9417) <= layer0_outputs(9965);
    outputs(9418) <= layer0_outputs(513);
    outputs(9419) <= (layer0_outputs(2719)) xor (layer0_outputs(9752));
    outputs(9420) <= (layer0_outputs(5172)) and (layer0_outputs(3673));
    outputs(9421) <= layer0_outputs(2153);
    outputs(9422) <= layer0_outputs(7762);
    outputs(9423) <= not(layer0_outputs(82)) or (layer0_outputs(7338));
    outputs(9424) <= not(layer0_outputs(4913));
    outputs(9425) <= (layer0_outputs(1943)) and not (layer0_outputs(1059));
    outputs(9426) <= not(layer0_outputs(1753));
    outputs(9427) <= not(layer0_outputs(1831));
    outputs(9428) <= not(layer0_outputs(3479));
    outputs(9429) <= layer0_outputs(2492);
    outputs(9430) <= (layer0_outputs(7074)) and not (layer0_outputs(720));
    outputs(9431) <= layer0_outputs(996);
    outputs(9432) <= not((layer0_outputs(968)) or (layer0_outputs(2301)));
    outputs(9433) <= (layer0_outputs(10086)) and (layer0_outputs(7725));
    outputs(9434) <= layer0_outputs(991);
    outputs(9435) <= layer0_outputs(7813);
    outputs(9436) <= layer0_outputs(9663);
    outputs(9437) <= not((layer0_outputs(6628)) or (layer0_outputs(3144)));
    outputs(9438) <= not(layer0_outputs(780));
    outputs(9439) <= not((layer0_outputs(7595)) or (layer0_outputs(2143)));
    outputs(9440) <= not(layer0_outputs(6787));
    outputs(9441) <= (layer0_outputs(9056)) and (layer0_outputs(8083));
    outputs(9442) <= not(layer0_outputs(7425)) or (layer0_outputs(1457));
    outputs(9443) <= not(layer0_outputs(8506));
    outputs(9444) <= layer0_outputs(2921);
    outputs(9445) <= (layer0_outputs(7100)) or (layer0_outputs(2557));
    outputs(9446) <= (layer0_outputs(7152)) and (layer0_outputs(4461));
    outputs(9447) <= (layer0_outputs(8457)) xor (layer0_outputs(7656));
    outputs(9448) <= layer0_outputs(3587);
    outputs(9449) <= not(layer0_outputs(4701));
    outputs(9450) <= (layer0_outputs(5987)) and (layer0_outputs(3074));
    outputs(9451) <= not(layer0_outputs(1420));
    outputs(9452) <= '0';
    outputs(9453) <= (layer0_outputs(5058)) xor (layer0_outputs(4203));
    outputs(9454) <= layer0_outputs(372);
    outputs(9455) <= (layer0_outputs(649)) and (layer0_outputs(5316));
    outputs(9456) <= layer0_outputs(6581);
    outputs(9457) <= not(layer0_outputs(8225));
    outputs(9458) <= (layer0_outputs(7120)) and not (layer0_outputs(8669));
    outputs(9459) <= not(layer0_outputs(7620));
    outputs(9460) <= not(layer0_outputs(2252));
    outputs(9461) <= not((layer0_outputs(4274)) or (layer0_outputs(8808)));
    outputs(9462) <= layer0_outputs(1316);
    outputs(9463) <= (layer0_outputs(2441)) or (layer0_outputs(8545));
    outputs(9464) <= layer0_outputs(1923);
    outputs(9465) <= not(layer0_outputs(4248));
    outputs(9466) <= not(layer0_outputs(610));
    outputs(9467) <= not(layer0_outputs(18)) or (layer0_outputs(6668));
    outputs(9468) <= layer0_outputs(5146);
    outputs(9469) <= layer0_outputs(9792);
    outputs(9470) <= not((layer0_outputs(6101)) xor (layer0_outputs(10194)));
    outputs(9471) <= layer0_outputs(6056);
    outputs(9472) <= not((layer0_outputs(7303)) xor (layer0_outputs(8150)));
    outputs(9473) <= not(layer0_outputs(931));
    outputs(9474) <= layer0_outputs(2976);
    outputs(9475) <= not((layer0_outputs(4066)) or (layer0_outputs(2536)));
    outputs(9476) <= not(layer0_outputs(4625));
    outputs(9477) <= not(layer0_outputs(766));
    outputs(9478) <= not(layer0_outputs(9249));
    outputs(9479) <= not(layer0_outputs(2742)) or (layer0_outputs(5142));
    outputs(9480) <= (layer0_outputs(3158)) and not (layer0_outputs(7592));
    outputs(9481) <= not((layer0_outputs(2729)) or (layer0_outputs(4637)));
    outputs(9482) <= not(layer0_outputs(2740));
    outputs(9483) <= (layer0_outputs(5083)) and not (layer0_outputs(110));
    outputs(9484) <= not((layer0_outputs(3437)) xor (layer0_outputs(6083)));
    outputs(9485) <= not(layer0_outputs(6914));
    outputs(9486) <= not((layer0_outputs(8416)) xor (layer0_outputs(10149)));
    outputs(9487) <= not(layer0_outputs(7661));
    outputs(9488) <= (layer0_outputs(8713)) and (layer0_outputs(4120));
    outputs(9489) <= not((layer0_outputs(8598)) xor (layer0_outputs(1660)));
    outputs(9490) <= layer0_outputs(3495);
    outputs(9491) <= layer0_outputs(4410);
    outputs(9492) <= not(layer0_outputs(7058));
    outputs(9493) <= (layer0_outputs(9021)) xor (layer0_outputs(2513));
    outputs(9494) <= (layer0_outputs(9027)) and not (layer0_outputs(7339));
    outputs(9495) <= layer0_outputs(2025);
    outputs(9496) <= not(layer0_outputs(8845));
    outputs(9497) <= (layer0_outputs(6678)) and (layer0_outputs(6438));
    outputs(9498) <= layer0_outputs(8976);
    outputs(9499) <= (layer0_outputs(2896)) xor (layer0_outputs(6905));
    outputs(9500) <= not(layer0_outputs(640));
    outputs(9501) <= (layer0_outputs(8366)) and not (layer0_outputs(1084));
    outputs(9502) <= (layer0_outputs(4870)) and not (layer0_outputs(1117));
    outputs(9503) <= not((layer0_outputs(8548)) xor (layer0_outputs(8457)));
    outputs(9504) <= not((layer0_outputs(9075)) or (layer0_outputs(9733)));
    outputs(9505) <= (layer0_outputs(6493)) and not (layer0_outputs(4550));
    outputs(9506) <= not((layer0_outputs(9777)) and (layer0_outputs(9913)));
    outputs(9507) <= not(layer0_outputs(8023));
    outputs(9508) <= not((layer0_outputs(2514)) or (layer0_outputs(7037)));
    outputs(9509) <= layer0_outputs(873);
    outputs(9510) <= not(layer0_outputs(3417));
    outputs(9511) <= layer0_outputs(9214);
    outputs(9512) <= layer0_outputs(8313);
    outputs(9513) <= not((layer0_outputs(9320)) or (layer0_outputs(10047)));
    outputs(9514) <= (layer0_outputs(5050)) and not (layer0_outputs(9696));
    outputs(9515) <= layer0_outputs(1125);
    outputs(9516) <= not(layer0_outputs(6194));
    outputs(9517) <= not((layer0_outputs(8467)) xor (layer0_outputs(763)));
    outputs(9518) <= layer0_outputs(121);
    outputs(9519) <= layer0_outputs(8950);
    outputs(9520) <= (layer0_outputs(4257)) xor (layer0_outputs(7920));
    outputs(9521) <= (layer0_outputs(6114)) xor (layer0_outputs(5448));
    outputs(9522) <= layer0_outputs(7707);
    outputs(9523) <= not(layer0_outputs(5304)) or (layer0_outputs(9184));
    outputs(9524) <= not((layer0_outputs(7599)) xor (layer0_outputs(2366)));
    outputs(9525) <= not(layer0_outputs(411)) or (layer0_outputs(7499));
    outputs(9526) <= not(layer0_outputs(1327));
    outputs(9527) <= not(layer0_outputs(2373));
    outputs(9528) <= not((layer0_outputs(5568)) xor (layer0_outputs(9058)));
    outputs(9529) <= (layer0_outputs(8568)) and not (layer0_outputs(8066));
    outputs(9530) <= not((layer0_outputs(3086)) xor (layer0_outputs(1647)));
    outputs(9531) <= not((layer0_outputs(3658)) xor (layer0_outputs(5356)));
    outputs(9532) <= layer0_outputs(4758);
    outputs(9533) <= (layer0_outputs(8529)) xor (layer0_outputs(4788));
    outputs(9534) <= layer0_outputs(3388);
    outputs(9535) <= layer0_outputs(9784);
    outputs(9536) <= not((layer0_outputs(3531)) or (layer0_outputs(2798)));
    outputs(9537) <= layer0_outputs(7081);
    outputs(9538) <= not(layer0_outputs(6225));
    outputs(9539) <= not((layer0_outputs(10101)) or (layer0_outputs(5880)));
    outputs(9540) <= not((layer0_outputs(9533)) xor (layer0_outputs(9174)));
    outputs(9541) <= (layer0_outputs(3160)) or (layer0_outputs(5789));
    outputs(9542) <= layer0_outputs(1195);
    outputs(9543) <= not((layer0_outputs(3093)) xor (layer0_outputs(1458)));
    outputs(9544) <= layer0_outputs(7601);
    outputs(9545) <= layer0_outputs(2222);
    outputs(9546) <= layer0_outputs(9353);
    outputs(9547) <= not(layer0_outputs(5586));
    outputs(9548) <= not(layer0_outputs(6567));
    outputs(9549) <= (layer0_outputs(5070)) and not (layer0_outputs(671));
    outputs(9550) <= layer0_outputs(824);
    outputs(9551) <= not(layer0_outputs(6185));
    outputs(9552) <= layer0_outputs(2622);
    outputs(9553) <= not((layer0_outputs(5656)) xor (layer0_outputs(10048)));
    outputs(9554) <= (layer0_outputs(4421)) or (layer0_outputs(5890));
    outputs(9555) <= (layer0_outputs(3371)) xor (layer0_outputs(8112));
    outputs(9556) <= not((layer0_outputs(5957)) xor (layer0_outputs(3525)));
    outputs(9557) <= (layer0_outputs(9732)) or (layer0_outputs(5393));
    outputs(9558) <= (layer0_outputs(2584)) or (layer0_outputs(7818));
    outputs(9559) <= not(layer0_outputs(4696));
    outputs(9560) <= (layer0_outputs(10180)) xor (layer0_outputs(6868));
    outputs(9561) <= layer0_outputs(4315);
    outputs(9562) <= layer0_outputs(3874);
    outputs(9563) <= not(layer0_outputs(6417));
    outputs(9564) <= (layer0_outputs(216)) and (layer0_outputs(8942));
    outputs(9565) <= (layer0_outputs(8608)) xor (layer0_outputs(6135));
    outputs(9566) <= (layer0_outputs(1168)) and not (layer0_outputs(7881));
    outputs(9567) <= not((layer0_outputs(4167)) xor (layer0_outputs(5908)));
    outputs(9568) <= not((layer0_outputs(2530)) xor (layer0_outputs(10142)));
    outputs(9569) <= not(layer0_outputs(3933));
    outputs(9570) <= layer0_outputs(1542);
    outputs(9571) <= not(layer0_outputs(3652)) or (layer0_outputs(2824));
    outputs(9572) <= layer0_outputs(4347);
    outputs(9573) <= (layer0_outputs(6541)) and (layer0_outputs(9269));
    outputs(9574) <= (layer0_outputs(2197)) xor (layer0_outputs(5993));
    outputs(9575) <= (layer0_outputs(6176)) xor (layer0_outputs(9319));
    outputs(9576) <= (layer0_outputs(2704)) and not (layer0_outputs(4121));
    outputs(9577) <= (layer0_outputs(3547)) and not (layer0_outputs(3638));
    outputs(9578) <= (layer0_outputs(9564)) and (layer0_outputs(520));
    outputs(9579) <= not((layer0_outputs(5453)) xor (layer0_outputs(8311)));
    outputs(9580) <= (layer0_outputs(2434)) or (layer0_outputs(8384));
    outputs(9581) <= layer0_outputs(1744);
    outputs(9582) <= not(layer0_outputs(5683));
    outputs(9583) <= not((layer0_outputs(1162)) or (layer0_outputs(3683)));
    outputs(9584) <= (layer0_outputs(3828)) or (layer0_outputs(3970));
    outputs(9585) <= (layer0_outputs(5535)) and (layer0_outputs(958));
    outputs(9586) <= not(layer0_outputs(5851)) or (layer0_outputs(5612));
    outputs(9587) <= (layer0_outputs(5816)) and (layer0_outputs(7231));
    outputs(9588) <= not(layer0_outputs(808));
    outputs(9589) <= layer0_outputs(1390);
    outputs(9590) <= not(layer0_outputs(9247));
    outputs(9591) <= not(layer0_outputs(10163));
    outputs(9592) <= layer0_outputs(8174);
    outputs(9593) <= not(layer0_outputs(4142)) or (layer0_outputs(6632));
    outputs(9594) <= not(layer0_outputs(6142));
    outputs(9595) <= not(layer0_outputs(3825)) or (layer0_outputs(678));
    outputs(9596) <= not((layer0_outputs(6564)) xor (layer0_outputs(5576)));
    outputs(9597) <= (layer0_outputs(6577)) xor (layer0_outputs(2283));
    outputs(9598) <= not(layer0_outputs(3199)) or (layer0_outputs(6062));
    outputs(9599) <= not((layer0_outputs(2637)) or (layer0_outputs(1586)));
    outputs(9600) <= not(layer0_outputs(5477));
    outputs(9601) <= (layer0_outputs(3576)) and not (layer0_outputs(673));
    outputs(9602) <= not((layer0_outputs(750)) or (layer0_outputs(9764)));
    outputs(9603) <= layer0_outputs(7512);
    outputs(9604) <= not(layer0_outputs(3020));
    outputs(9605) <= not((layer0_outputs(5069)) and (layer0_outputs(8751)));
    outputs(9606) <= (layer0_outputs(6683)) and not (layer0_outputs(7539));
    outputs(9607) <= not((layer0_outputs(6333)) xor (layer0_outputs(3551)));
    outputs(9608) <= (layer0_outputs(831)) and (layer0_outputs(1481));
    outputs(9609) <= (layer0_outputs(5339)) and not (layer0_outputs(1944));
    outputs(9610) <= not(layer0_outputs(3062));
    outputs(9611) <= (layer0_outputs(8276)) and (layer0_outputs(1405));
    outputs(9612) <= layer0_outputs(3500);
    outputs(9613) <= (layer0_outputs(8297)) and (layer0_outputs(1483));
    outputs(9614) <= layer0_outputs(2579);
    outputs(9615) <= not(layer0_outputs(7973)) or (layer0_outputs(2511));
    outputs(9616) <= not((layer0_outputs(7089)) xor (layer0_outputs(2942)));
    outputs(9617) <= not(layer0_outputs(2614)) or (layer0_outputs(2353));
    outputs(9618) <= layer0_outputs(7915);
    outputs(9619) <= not(layer0_outputs(634));
    outputs(9620) <= (layer0_outputs(2876)) and (layer0_outputs(3982));
    outputs(9621) <= (layer0_outputs(9080)) and (layer0_outputs(5680));
    outputs(9622) <= not(layer0_outputs(6736));
    outputs(9623) <= (layer0_outputs(5290)) or (layer0_outputs(4341));
    outputs(9624) <= (layer0_outputs(8119)) and not (layer0_outputs(7402));
    outputs(9625) <= (layer0_outputs(281)) xor (layer0_outputs(590));
    outputs(9626) <= layer0_outputs(9116);
    outputs(9627) <= not(layer0_outputs(1175));
    outputs(9628) <= not((layer0_outputs(5459)) or (layer0_outputs(6691)));
    outputs(9629) <= layer0_outputs(9437);
    outputs(9630) <= (layer0_outputs(4029)) and not (layer0_outputs(5071));
    outputs(9631) <= not(layer0_outputs(7204));
    outputs(9632) <= (layer0_outputs(8560)) and not (layer0_outputs(7940));
    outputs(9633) <= not((layer0_outputs(7647)) or (layer0_outputs(6145)));
    outputs(9634) <= not((layer0_outputs(6014)) xor (layer0_outputs(2594)));
    outputs(9635) <= (layer0_outputs(1297)) xor (layer0_outputs(9975));
    outputs(9636) <= (layer0_outputs(8955)) and (layer0_outputs(5548));
    outputs(9637) <= (layer0_outputs(4484)) and (layer0_outputs(9126));
    outputs(9638) <= not(layer0_outputs(6517));
    outputs(9639) <= (layer0_outputs(5996)) and (layer0_outputs(8559));
    outputs(9640) <= not((layer0_outputs(315)) xor (layer0_outputs(6908)));
    outputs(9641) <= not((layer0_outputs(4102)) and (layer0_outputs(2165)));
    outputs(9642) <= layer0_outputs(1734);
    outputs(9643) <= not((layer0_outputs(5815)) or (layer0_outputs(8772)));
    outputs(9644) <= not(layer0_outputs(574)) or (layer0_outputs(5082));
    outputs(9645) <= layer0_outputs(3205);
    outputs(9646) <= not((layer0_outputs(9232)) xor (layer0_outputs(4089)));
    outputs(9647) <= not((layer0_outputs(3478)) xor (layer0_outputs(1368)));
    outputs(9648) <= (layer0_outputs(2199)) and not (layer0_outputs(2292));
    outputs(9649) <= (layer0_outputs(5641)) and not (layer0_outputs(4952));
    outputs(9650) <= (layer0_outputs(2119)) xor (layer0_outputs(7884));
    outputs(9651) <= not(layer0_outputs(1348));
    outputs(9652) <= (layer0_outputs(982)) and not (layer0_outputs(3470));
    outputs(9653) <= layer0_outputs(8446);
    outputs(9654) <= (layer0_outputs(147)) and not (layer0_outputs(9755));
    outputs(9655) <= (layer0_outputs(1163)) and not (layer0_outputs(5263));
    outputs(9656) <= not(layer0_outputs(4481));
    outputs(9657) <= not((layer0_outputs(8304)) or (layer0_outputs(6997)));
    outputs(9658) <= (layer0_outputs(9115)) and not (layer0_outputs(7967));
    outputs(9659) <= not(layer0_outputs(9646)) or (layer0_outputs(6461));
    outputs(9660) <= not(layer0_outputs(230));
    outputs(9661) <= (layer0_outputs(2182)) and not (layer0_outputs(966));
    outputs(9662) <= not(layer0_outputs(169));
    outputs(9663) <= layer0_outputs(1350);
    outputs(9664) <= (layer0_outputs(9260)) xor (layer0_outputs(5123));
    outputs(9665) <= not((layer0_outputs(1848)) xor (layer0_outputs(3369)));
    outputs(9666) <= not(layer0_outputs(7728));
    outputs(9667) <= layer0_outputs(1610);
    outputs(9668) <= layer0_outputs(3713);
    outputs(9669) <= not((layer0_outputs(644)) xor (layer0_outputs(1611)));
    outputs(9670) <= not((layer0_outputs(7287)) and (layer0_outputs(1465)));
    outputs(9671) <= not((layer0_outputs(8270)) and (layer0_outputs(4020)));
    outputs(9672) <= not(layer0_outputs(10231));
    outputs(9673) <= (layer0_outputs(2519)) or (layer0_outputs(8530));
    outputs(9674) <= not(layer0_outputs(4189));
    outputs(9675) <= (layer0_outputs(7610)) and (layer0_outputs(5149));
    outputs(9676) <= not(layer0_outputs(2331));
    outputs(9677) <= (layer0_outputs(7454)) and not (layer0_outputs(3579));
    outputs(9678) <= layer0_outputs(8389);
    outputs(9679) <= layer0_outputs(1239);
    outputs(9680) <= not((layer0_outputs(8469)) or (layer0_outputs(8639)));
    outputs(9681) <= not((layer0_outputs(10232)) xor (layer0_outputs(4813)));
    outputs(9682) <= (layer0_outputs(374)) xor (layer0_outputs(7858));
    outputs(9683) <= layer0_outputs(2878);
    outputs(9684) <= layer0_outputs(2954);
    outputs(9685) <= not(layer0_outputs(5249));
    outputs(9686) <= layer0_outputs(6976);
    outputs(9687) <= (layer0_outputs(5392)) xor (layer0_outputs(2011));
    outputs(9688) <= (layer0_outputs(3597)) and not (layer0_outputs(7461));
    outputs(9689) <= (layer0_outputs(4357)) xor (layer0_outputs(5313));
    outputs(9690) <= not((layer0_outputs(7789)) xor (layer0_outputs(7013)));
    outputs(9691) <= layer0_outputs(7099);
    outputs(9692) <= not(layer0_outputs(8561));
    outputs(9693) <= not(layer0_outputs(7537));
    outputs(9694) <= not((layer0_outputs(10191)) xor (layer0_outputs(2984)));
    outputs(9695) <= (layer0_outputs(7196)) and not (layer0_outputs(5025));
    outputs(9696) <= (layer0_outputs(5796)) xor (layer0_outputs(9880));
    outputs(9697) <= not((layer0_outputs(2781)) or (layer0_outputs(8224)));
    outputs(9698) <= not((layer0_outputs(8152)) xor (layer0_outputs(633)));
    outputs(9699) <= (layer0_outputs(929)) xor (layer0_outputs(4308));
    outputs(9700) <= not(layer0_outputs(5451));
    outputs(9701) <= (layer0_outputs(2349)) or (layer0_outputs(1359));
    outputs(9702) <= not(layer0_outputs(9017));
    outputs(9703) <= not(layer0_outputs(9996));
    outputs(9704) <= layer0_outputs(2190);
    outputs(9705) <= not((layer0_outputs(7592)) xor (layer0_outputs(4475)));
    outputs(9706) <= layer0_outputs(1657);
    outputs(9707) <= not((layer0_outputs(7102)) xor (layer0_outputs(1264)));
    outputs(9708) <= layer0_outputs(10029);
    outputs(9709) <= layer0_outputs(2290);
    outputs(9710) <= not(layer0_outputs(4405));
    outputs(9711) <= (layer0_outputs(2221)) and not (layer0_outputs(10097));
    outputs(9712) <= (layer0_outputs(1208)) xor (layer0_outputs(7171));
    outputs(9713) <= not((layer0_outputs(2484)) xor (layer0_outputs(7769)));
    outputs(9714) <= not((layer0_outputs(3359)) xor (layer0_outputs(9661)));
    outputs(9715) <= (layer0_outputs(5819)) and not (layer0_outputs(3002));
    outputs(9716) <= (layer0_outputs(5823)) or (layer0_outputs(5750));
    outputs(9717) <= not(layer0_outputs(3725));
    outputs(9718) <= not((layer0_outputs(2895)) or (layer0_outputs(1580)));
    outputs(9719) <= layer0_outputs(5275);
    outputs(9720) <= (layer0_outputs(4182)) xor (layer0_outputs(1122));
    outputs(9721) <= (layer0_outputs(1183)) and (layer0_outputs(7937));
    outputs(9722) <= (layer0_outputs(6134)) and not (layer0_outputs(9440));
    outputs(9723) <= layer0_outputs(8762);
    outputs(9724) <= not(layer0_outputs(2026));
    outputs(9725) <= (layer0_outputs(8382)) and (layer0_outputs(4692));
    outputs(9726) <= not(layer0_outputs(1157)) or (layer0_outputs(830));
    outputs(9727) <= layer0_outputs(6842);
    outputs(9728) <= (layer0_outputs(3270)) and (layer0_outputs(8875));
    outputs(9729) <= not((layer0_outputs(10039)) or (layer0_outputs(9715)));
    outputs(9730) <= (layer0_outputs(7436)) or (layer0_outputs(5046));
    outputs(9731) <= not(layer0_outputs(3630));
    outputs(9732) <= not(layer0_outputs(9358));
    outputs(9733) <= (layer0_outputs(1982)) and (layer0_outputs(6683));
    outputs(9734) <= (layer0_outputs(8414)) xor (layer0_outputs(2957));
    outputs(9735) <= layer0_outputs(7933);
    outputs(9736) <= (layer0_outputs(7494)) and (layer0_outputs(2659));
    outputs(9737) <= not(layer0_outputs(270));
    outputs(9738) <= layer0_outputs(5139);
    outputs(9739) <= not((layer0_outputs(9999)) xor (layer0_outputs(4519)));
    outputs(9740) <= layer0_outputs(8597);
    outputs(9741) <= not(layer0_outputs(7883));
    outputs(9742) <= (layer0_outputs(7976)) or (layer0_outputs(8085));
    outputs(9743) <= layer0_outputs(1317);
    outputs(9744) <= layer0_outputs(1301);
    outputs(9745) <= (layer0_outputs(8401)) xor (layer0_outputs(8026));
    outputs(9746) <= not((layer0_outputs(7602)) xor (layer0_outputs(2273)));
    outputs(9747) <= layer0_outputs(9928);
    outputs(9748) <= (layer0_outputs(1623)) and not (layer0_outputs(7740));
    outputs(9749) <= layer0_outputs(7214);
    outputs(9750) <= not(layer0_outputs(3442));
    outputs(9751) <= not((layer0_outputs(1084)) xor (layer0_outputs(6729)));
    outputs(9752) <= layer0_outputs(10020);
    outputs(9753) <= layer0_outputs(1694);
    outputs(9754) <= not((layer0_outputs(4130)) or (layer0_outputs(3880)));
    outputs(9755) <= layer0_outputs(2673);
    outputs(9756) <= layer0_outputs(905);
    outputs(9757) <= layer0_outputs(10078);
    outputs(9758) <= layer0_outputs(5353);
    outputs(9759) <= layer0_outputs(6697);
    outputs(9760) <= not(layer0_outputs(9551));
    outputs(9761) <= (layer0_outputs(5543)) xor (layer0_outputs(887));
    outputs(9762) <= not((layer0_outputs(8963)) xor (layer0_outputs(5703)));
    outputs(9763) <= (layer0_outputs(848)) xor (layer0_outputs(5344));
    outputs(9764) <= not((layer0_outputs(6710)) and (layer0_outputs(4810)));
    outputs(9765) <= not((layer0_outputs(3023)) xor (layer0_outputs(8395)));
    outputs(9766) <= not(layer0_outputs(7325));
    outputs(9767) <= (layer0_outputs(1394)) xor (layer0_outputs(7928));
    outputs(9768) <= not(layer0_outputs(9856));
    outputs(9769) <= not(layer0_outputs(7945));
    outputs(9770) <= (layer0_outputs(9516)) and (layer0_outputs(3400));
    outputs(9771) <= not(layer0_outputs(9550)) or (layer0_outputs(3966));
    outputs(9772) <= not((layer0_outputs(8037)) and (layer0_outputs(4997)));
    outputs(9773) <= not((layer0_outputs(6175)) xor (layer0_outputs(1655)));
    outputs(9774) <= (layer0_outputs(256)) xor (layer0_outputs(3317));
    outputs(9775) <= not(layer0_outputs(1523));
    outputs(9776) <= not(layer0_outputs(1367));
    outputs(9777) <= layer0_outputs(1886);
    outputs(9778) <= (layer0_outputs(7889)) and not (layer0_outputs(4825));
    outputs(9779) <= (layer0_outputs(7411)) or (layer0_outputs(4179));
    outputs(9780) <= layer0_outputs(5587);
    outputs(9781) <= not(layer0_outputs(9220));
    outputs(9782) <= (layer0_outputs(1083)) xor (layer0_outputs(8912));
    outputs(9783) <= (layer0_outputs(4173)) xor (layer0_outputs(3105));
    outputs(9784) <= (layer0_outputs(1414)) and not (layer0_outputs(2076));
    outputs(9785) <= layer0_outputs(9577);
    outputs(9786) <= layer0_outputs(1126);
    outputs(9787) <= layer0_outputs(7380);
    outputs(9788) <= (layer0_outputs(1470)) and not (layer0_outputs(9961));
    outputs(9789) <= layer0_outputs(6989);
    outputs(9790) <= (layer0_outputs(2265)) xor (layer0_outputs(9320));
    outputs(9791) <= not((layer0_outputs(3141)) or (layer0_outputs(14)));
    outputs(9792) <= (layer0_outputs(7148)) and not (layer0_outputs(5409));
    outputs(9793) <= layer0_outputs(6516);
    outputs(9794) <= layer0_outputs(1062);
    outputs(9795) <= not((layer0_outputs(4535)) or (layer0_outputs(7990)));
    outputs(9796) <= layer0_outputs(9703);
    outputs(9797) <= not(layer0_outputs(5090));
    outputs(9798) <= not((layer0_outputs(6159)) xor (layer0_outputs(7674)));
    outputs(9799) <= not(layer0_outputs(1435));
    outputs(9800) <= layer0_outputs(7008);
    outputs(9801) <= layer0_outputs(8968);
    outputs(9802) <= layer0_outputs(7363);
    outputs(9803) <= not(layer0_outputs(2003));
    outputs(9804) <= (layer0_outputs(6831)) and not (layer0_outputs(544));
    outputs(9805) <= (layer0_outputs(6642)) and not (layer0_outputs(1978));
    outputs(9806) <= not((layer0_outputs(653)) or (layer0_outputs(6865)));
    outputs(9807) <= layer0_outputs(8033);
    outputs(9808) <= layer0_outputs(6266);
    outputs(9809) <= not(layer0_outputs(9523)) or (layer0_outputs(3453));
    outputs(9810) <= not(layer0_outputs(469));
    outputs(9811) <= not(layer0_outputs(1092));
    outputs(9812) <= (layer0_outputs(7458)) and not (layer0_outputs(2129));
    outputs(9813) <= (layer0_outputs(5081)) xor (layer0_outputs(1858));
    outputs(9814) <= (layer0_outputs(9004)) xor (layer0_outputs(8236));
    outputs(9815) <= layer0_outputs(5762);
    outputs(9816) <= layer0_outputs(7343);
    outputs(9817) <= (layer0_outputs(8202)) xor (layer0_outputs(8429));
    outputs(9818) <= (layer0_outputs(9648)) and not (layer0_outputs(5815));
    outputs(9819) <= layer0_outputs(5482);
    outputs(9820) <= layer0_outputs(4210);
    outputs(9821) <= (layer0_outputs(5284)) xor (layer0_outputs(7136));
    outputs(9822) <= (layer0_outputs(332)) and not (layer0_outputs(4097));
    outputs(9823) <= (layer0_outputs(7980)) and not (layer0_outputs(10204));
    outputs(9824) <= (layer0_outputs(2546)) and not (layer0_outputs(4964));
    outputs(9825) <= not(layer0_outputs(6573));
    outputs(9826) <= layer0_outputs(8362);
    outputs(9827) <= (layer0_outputs(1963)) and not (layer0_outputs(5669));
    outputs(9828) <= not((layer0_outputs(8686)) xor (layer0_outputs(8933)));
    outputs(9829) <= (layer0_outputs(539)) and not (layer0_outputs(267));
    outputs(9830) <= not(layer0_outputs(1295));
    outputs(9831) <= not(layer0_outputs(2946));
    outputs(9832) <= (layer0_outputs(7123)) and not (layer0_outputs(5975));
    outputs(9833) <= layer0_outputs(7995);
    outputs(9834) <= not((layer0_outputs(1986)) xor (layer0_outputs(7281)));
    outputs(9835) <= not(layer0_outputs(4751));
    outputs(9836) <= layer0_outputs(7888);
    outputs(9837) <= layer0_outputs(4310);
    outputs(9838) <= not(layer0_outputs(3790));
    outputs(9839) <= not(layer0_outputs(2064));
    outputs(9840) <= (layer0_outputs(9824)) and not (layer0_outputs(7713));
    outputs(9841) <= not(layer0_outputs(5456));
    outputs(9842) <= not(layer0_outputs(8920));
    outputs(9843) <= not(layer0_outputs(625));
    outputs(9844) <= (layer0_outputs(1856)) and not (layer0_outputs(4138));
    outputs(9845) <= layer0_outputs(5768);
    outputs(9846) <= (layer0_outputs(9351)) xor (layer0_outputs(5158));
    outputs(9847) <= not((layer0_outputs(7080)) xor (layer0_outputs(2682)));
    outputs(9848) <= (layer0_outputs(132)) or (layer0_outputs(8900));
    outputs(9849) <= (layer0_outputs(419)) xor (layer0_outputs(8482));
    outputs(9850) <= (layer0_outputs(860)) and (layer0_outputs(817));
    outputs(9851) <= not(layer0_outputs(6651));
    outputs(9852) <= (layer0_outputs(7656)) or (layer0_outputs(899));
    outputs(9853) <= not((layer0_outputs(6141)) xor (layer0_outputs(3694)));
    outputs(9854) <= layer0_outputs(2499);
    outputs(9855) <= (layer0_outputs(7569)) and not (layer0_outputs(5751));
    outputs(9856) <= not(layer0_outputs(4571));
    outputs(9857) <= (layer0_outputs(338)) and not (layer0_outputs(2014));
    outputs(9858) <= not(layer0_outputs(153));
    outputs(9859) <= layer0_outputs(4552);
    outputs(9860) <= (layer0_outputs(8647)) and (layer0_outputs(8334));
    outputs(9861) <= not((layer0_outputs(5183)) or (layer0_outputs(1433)));
    outputs(9862) <= not(layer0_outputs(5921));
    outputs(9863) <= not(layer0_outputs(7263)) or (layer0_outputs(1471));
    outputs(9864) <= (layer0_outputs(6003)) and not (layer0_outputs(5956));
    outputs(9865) <= (layer0_outputs(8122)) xor (layer0_outputs(6446));
    outputs(9866) <= not(layer0_outputs(3134));
    outputs(9867) <= not(layer0_outputs(9610)) or (layer0_outputs(5970));
    outputs(9868) <= not(layer0_outputs(9669));
    outputs(9869) <= not((layer0_outputs(8998)) and (layer0_outputs(1948)));
    outputs(9870) <= not((layer0_outputs(3187)) xor (layer0_outputs(4019)));
    outputs(9871) <= layer0_outputs(2809);
    outputs(9872) <= not(layer0_outputs(8460));
    outputs(9873) <= not(layer0_outputs(858));
    outputs(9874) <= not(layer0_outputs(793));
    outputs(9875) <= layer0_outputs(8125);
    outputs(9876) <= layer0_outputs(4055);
    outputs(9877) <= not(layer0_outputs(10163)) or (layer0_outputs(8922));
    outputs(9878) <= not((layer0_outputs(8346)) or (layer0_outputs(3563)));
    outputs(9879) <= (layer0_outputs(7698)) xor (layer0_outputs(1531));
    outputs(9880) <= not(layer0_outputs(6237));
    outputs(9881) <= not((layer0_outputs(7277)) and (layer0_outputs(636)));
    outputs(9882) <= not(layer0_outputs(4782));
    outputs(9883) <= not((layer0_outputs(8657)) xor (layer0_outputs(5376)));
    outputs(9884) <= not(layer0_outputs(729));
    outputs(9885) <= (layer0_outputs(5095)) and not (layer0_outputs(7262));
    outputs(9886) <= not(layer0_outputs(8512));
    outputs(9887) <= (layer0_outputs(2175)) and (layer0_outputs(4815));
    outputs(9888) <= not(layer0_outputs(4386));
    outputs(9889) <= not((layer0_outputs(1641)) xor (layer0_outputs(5429)));
    outputs(9890) <= layer0_outputs(9939);
    outputs(9891) <= not(layer0_outputs(8576));
    outputs(9892) <= not((layer0_outputs(5207)) xor (layer0_outputs(2135)));
    outputs(9893) <= not((layer0_outputs(10181)) xor (layer0_outputs(3483)));
    outputs(9894) <= (layer0_outputs(10103)) xor (layer0_outputs(981));
    outputs(9895) <= '0';
    outputs(9896) <= not((layer0_outputs(2850)) or (layer0_outputs(952)));
    outputs(9897) <= not((layer0_outputs(9001)) xor (layer0_outputs(3721)));
    outputs(9898) <= not((layer0_outputs(1954)) xor (layer0_outputs(9472)));
    outputs(9899) <= (layer0_outputs(2377)) and not (layer0_outputs(7905));
    outputs(9900) <= not((layer0_outputs(358)) or (layer0_outputs(1990)));
    outputs(9901) <= (layer0_outputs(3828)) and not (layer0_outputs(4047));
    outputs(9902) <= not(layer0_outputs(7925));
    outputs(9903) <= layer0_outputs(5309);
    outputs(9904) <= layer0_outputs(5552);
    outputs(9905) <= not(layer0_outputs(2628));
    outputs(9906) <= not(layer0_outputs(3969));
    outputs(9907) <= not(layer0_outputs(7887));
    outputs(9908) <= layer0_outputs(2052);
    outputs(9909) <= not(layer0_outputs(4354));
    outputs(9910) <= not((layer0_outputs(9866)) or (layer0_outputs(5411)));
    outputs(9911) <= layer0_outputs(4565);
    outputs(9912) <= layer0_outputs(10197);
    outputs(9913) <= (layer0_outputs(9822)) and (layer0_outputs(3195));
    outputs(9914) <= (layer0_outputs(1541)) and not (layer0_outputs(201));
    outputs(9915) <= (layer0_outputs(6884)) xor (layer0_outputs(623));
    outputs(9916) <= not((layer0_outputs(1389)) or (layer0_outputs(6417)));
    outputs(9917) <= not((layer0_outputs(7609)) xor (layer0_outputs(3553)));
    outputs(9918) <= (layer0_outputs(9561)) and not (layer0_outputs(1304));
    outputs(9919) <= not((layer0_outputs(9538)) or (layer0_outputs(7659)));
    outputs(9920) <= layer0_outputs(6524);
    outputs(9921) <= layer0_outputs(7663);
    outputs(9922) <= not((layer0_outputs(3343)) and (layer0_outputs(9657)));
    outputs(9923) <= (layer0_outputs(257)) xor (layer0_outputs(10147));
    outputs(9924) <= not(layer0_outputs(5979));
    outputs(9925) <= not((layer0_outputs(2006)) xor (layer0_outputs(5545)));
    outputs(9926) <= not(layer0_outputs(7260));
    outputs(9927) <= not(layer0_outputs(2615));
    outputs(9928) <= not(layer0_outputs(767));
    outputs(9929) <= layer0_outputs(1916);
    outputs(9930) <= not((layer0_outputs(26)) xor (layer0_outputs(384)));
    outputs(9931) <= not(layer0_outputs(2624));
    outputs(9932) <= not((layer0_outputs(9969)) and (layer0_outputs(2655)));
    outputs(9933) <= layer0_outputs(9162);
    outputs(9934) <= (layer0_outputs(10165)) and not (layer0_outputs(754));
    outputs(9935) <= not(layer0_outputs(8978));
    outputs(9936) <= (layer0_outputs(9613)) and (layer0_outputs(1145));
    outputs(9937) <= not(layer0_outputs(4204));
    outputs(9938) <= (layer0_outputs(2818)) and not (layer0_outputs(2113));
    outputs(9939) <= not((layer0_outputs(8918)) xor (layer0_outputs(8325)));
    outputs(9940) <= not(layer0_outputs(40));
    outputs(9941) <= (layer0_outputs(2677)) xor (layer0_outputs(1960));
    outputs(9942) <= (layer0_outputs(8945)) xor (layer0_outputs(9338));
    outputs(9943) <= layer0_outputs(1644);
    outputs(9944) <= not((layer0_outputs(4588)) xor (layer0_outputs(6339)));
    outputs(9945) <= not(layer0_outputs(2352));
    outputs(9946) <= layer0_outputs(9647);
    outputs(9947) <= not(layer0_outputs(8845));
    outputs(9948) <= (layer0_outputs(9987)) and not (layer0_outputs(7630));
    outputs(9949) <= (layer0_outputs(4774)) and not (layer0_outputs(66));
    outputs(9950) <= not((layer0_outputs(7053)) or (layer0_outputs(9247)));
    outputs(9951) <= not((layer0_outputs(3795)) xor (layer0_outputs(3004)));
    outputs(9952) <= not((layer0_outputs(2461)) xor (layer0_outputs(6685)));
    outputs(9953) <= layer0_outputs(4837);
    outputs(9954) <= not((layer0_outputs(5148)) xor (layer0_outputs(9321)));
    outputs(9955) <= layer0_outputs(1307);
    outputs(9956) <= not(layer0_outputs(3903));
    outputs(9957) <= not(layer0_outputs(7243));
    outputs(9958) <= (layer0_outputs(2259)) xor (layer0_outputs(5210));
    outputs(9959) <= (layer0_outputs(3597)) and not (layer0_outputs(6973));
    outputs(9960) <= not((layer0_outputs(9524)) xor (layer0_outputs(3083)));
    outputs(9961) <= (layer0_outputs(2055)) or (layer0_outputs(3429));
    outputs(9962) <= (layer0_outputs(4100)) and not (layer0_outputs(7860));
    outputs(9963) <= (layer0_outputs(9811)) or (layer0_outputs(5940));
    outputs(9964) <= (layer0_outputs(7245)) xor (layer0_outputs(6609));
    outputs(9965) <= not(layer0_outputs(3217));
    outputs(9966) <= not(layer0_outputs(2330));
    outputs(9967) <= not((layer0_outputs(9637)) xor (layer0_outputs(4940)));
    outputs(9968) <= (layer0_outputs(6563)) and not (layer0_outputs(7800));
    outputs(9969) <= not(layer0_outputs(3875));
    outputs(9970) <= layer0_outputs(7101);
    outputs(9971) <= layer0_outputs(9701);
    outputs(9972) <= not(layer0_outputs(7451));
    outputs(9973) <= (layer0_outputs(2410)) and not (layer0_outputs(9293));
    outputs(9974) <= (layer0_outputs(1812)) and (layer0_outputs(6887));
    outputs(9975) <= not(layer0_outputs(9346));
    outputs(9976) <= layer0_outputs(2890);
    outputs(9977) <= layer0_outputs(1251);
    outputs(9978) <= not((layer0_outputs(1443)) xor (layer0_outputs(1043)));
    outputs(9979) <= not(layer0_outputs(8662));
    outputs(9980) <= not(layer0_outputs(7084));
    outputs(9981) <= (layer0_outputs(4979)) xor (layer0_outputs(1332));
    outputs(9982) <= not(layer0_outputs(2891)) or (layer0_outputs(6751));
    outputs(9983) <= (layer0_outputs(8560)) and not (layer0_outputs(6777));
    outputs(9984) <= not(layer0_outputs(9993));
    outputs(9985) <= not((layer0_outputs(4842)) xor (layer0_outputs(3007)));
    outputs(9986) <= (layer0_outputs(2867)) xor (layer0_outputs(5567));
    outputs(9987) <= (layer0_outputs(3678)) and not (layer0_outputs(1339));
    outputs(9988) <= not((layer0_outputs(5072)) or (layer0_outputs(2038)));
    outputs(9989) <= layer0_outputs(9855);
    outputs(9990) <= not(layer0_outputs(5529));
    outputs(9991) <= not(layer0_outputs(8358));
    outputs(9992) <= (layer0_outputs(7933)) and not (layer0_outputs(4980));
    outputs(9993) <= layer0_outputs(3412);
    outputs(9994) <= not(layer0_outputs(4591));
    outputs(9995) <= layer0_outputs(10195);
    outputs(9996) <= layer0_outputs(998);
    outputs(9997) <= not((layer0_outputs(8138)) xor (layer0_outputs(3261)));
    outputs(9998) <= (layer0_outputs(9404)) xor (layer0_outputs(1236));
    outputs(9999) <= layer0_outputs(7654);
    outputs(10000) <= not(layer0_outputs(1497)) or (layer0_outputs(416));
    outputs(10001) <= not(layer0_outputs(2913));
    outputs(10002) <= not(layer0_outputs(7981));
    outputs(10003) <= (layer0_outputs(4195)) and not (layer0_outputs(5896));
    outputs(10004) <= not(layer0_outputs(8929));
    outputs(10005) <= not(layer0_outputs(9529)) or (layer0_outputs(5006));
    outputs(10006) <= (layer0_outputs(661)) and not (layer0_outputs(6854));
    outputs(10007) <= not(layer0_outputs(2674)) or (layer0_outputs(1833));
    outputs(10008) <= not((layer0_outputs(9931)) xor (layer0_outputs(8689)));
    outputs(10009) <= not(layer0_outputs(2364));
    outputs(10010) <= not(layer0_outputs(5212));
    outputs(10011) <= (layer0_outputs(196)) and not (layer0_outputs(5633));
    outputs(10012) <= layer0_outputs(3593);
    outputs(10013) <= layer0_outputs(6976);
    outputs(10014) <= not(layer0_outputs(4237));
    outputs(10015) <= layer0_outputs(3967);
    outputs(10016) <= not((layer0_outputs(6945)) and (layer0_outputs(1894)));
    outputs(10017) <= not(layer0_outputs(1086));
    outputs(10018) <= layer0_outputs(9926);
    outputs(10019) <= not(layer0_outputs(4694));
    outputs(10020) <= (layer0_outputs(4436)) and not (layer0_outputs(3419));
    outputs(10021) <= (layer0_outputs(8098)) xor (layer0_outputs(9359));
    outputs(10022) <= (layer0_outputs(9202)) and not (layer0_outputs(6878));
    outputs(10023) <= not((layer0_outputs(2066)) xor (layer0_outputs(6833)));
    outputs(10024) <= not(layer0_outputs(7496));
    outputs(10025) <= not(layer0_outputs(2158));
    outputs(10026) <= layer0_outputs(6671);
    outputs(10027) <= layer0_outputs(1456);
    outputs(10028) <= (layer0_outputs(6007)) or (layer0_outputs(2803));
    outputs(10029) <= (layer0_outputs(2393)) and not (layer0_outputs(2392));
    outputs(10030) <= not(layer0_outputs(3062));
    outputs(10031) <= (layer0_outputs(2918)) xor (layer0_outputs(130));
    outputs(10032) <= layer0_outputs(9339);
    outputs(10033) <= layer0_outputs(5501);
    outputs(10034) <= (layer0_outputs(744)) xor (layer0_outputs(9994));
    outputs(10035) <= not((layer0_outputs(6538)) xor (layer0_outputs(5633)));
    outputs(10036) <= (layer0_outputs(6095)) xor (layer0_outputs(7820));
    outputs(10037) <= (layer0_outputs(5900)) and not (layer0_outputs(4095));
    outputs(10038) <= (layer0_outputs(3294)) and (layer0_outputs(5892));
    outputs(10039) <= (layer0_outputs(868)) xor (layer0_outputs(9034));
    outputs(10040) <= not((layer0_outputs(8912)) xor (layer0_outputs(1664)));
    outputs(10041) <= (layer0_outputs(3555)) and not (layer0_outputs(5219));
    outputs(10042) <= not((layer0_outputs(1421)) or (layer0_outputs(8000)));
    outputs(10043) <= layer0_outputs(4856);
    outputs(10044) <= not(layer0_outputs(1872));
    outputs(10045) <= (layer0_outputs(6381)) xor (layer0_outputs(4603));
    outputs(10046) <= layer0_outputs(3024);
    outputs(10047) <= layer0_outputs(9822);
    outputs(10048) <= not(layer0_outputs(5078));
    outputs(10049) <= (layer0_outputs(3431)) and not (layer0_outputs(7187));
    outputs(10050) <= layer0_outputs(8627);
    outputs(10051) <= (layer0_outputs(7157)) or (layer0_outputs(9965));
    outputs(10052) <= not(layer0_outputs(8520));
    outputs(10053) <= (layer0_outputs(2072)) and not (layer0_outputs(10222));
    outputs(10054) <= not(layer0_outputs(7406));
    outputs(10055) <= (layer0_outputs(1300)) and not (layer0_outputs(3643));
    outputs(10056) <= not(layer0_outputs(3097));
    outputs(10057) <= layer0_outputs(6988);
    outputs(10058) <= not((layer0_outputs(8466)) xor (layer0_outputs(7060)));
    outputs(10059) <= (layer0_outputs(2152)) xor (layer0_outputs(5575));
    outputs(10060) <= (layer0_outputs(6089)) xor (layer0_outputs(1648));
    outputs(10061) <= (layer0_outputs(5195)) and not (layer0_outputs(3737));
    outputs(10062) <= not(layer0_outputs(9903));
    outputs(10063) <= not(layer0_outputs(4654));
    outputs(10064) <= (layer0_outputs(5620)) or (layer0_outputs(6035));
    outputs(10065) <= (layer0_outputs(6981)) and not (layer0_outputs(1142));
    outputs(10066) <= not(layer0_outputs(2156)) or (layer0_outputs(4146));
    outputs(10067) <= (layer0_outputs(4178)) and not (layer0_outputs(8469));
    outputs(10068) <= not(layer0_outputs(10068));
    outputs(10069) <= (layer0_outputs(3381)) xor (layer0_outputs(7044));
    outputs(10070) <= layer0_outputs(102);
    outputs(10071) <= layer0_outputs(731);
    outputs(10072) <= not(layer0_outputs(8215));
    outputs(10073) <= not((layer0_outputs(784)) xor (layer0_outputs(7145)));
    outputs(10074) <= not((layer0_outputs(2127)) xor (layer0_outputs(1007)));
    outputs(10075) <= (layer0_outputs(8571)) and (layer0_outputs(4054));
    outputs(10076) <= not((layer0_outputs(5838)) or (layer0_outputs(4923)));
    outputs(10077) <= not(layer0_outputs(5887));
    outputs(10078) <= layer0_outputs(5374);
    outputs(10079) <= not(layer0_outputs(8673));
    outputs(10080) <= not(layer0_outputs(4175)) or (layer0_outputs(1273));
    outputs(10081) <= not(layer0_outputs(9589));
    outputs(10082) <= not((layer0_outputs(2909)) xor (layer0_outputs(6226)));
    outputs(10083) <= not(layer0_outputs(3768));
    outputs(10084) <= layer0_outputs(8516);
    outputs(10085) <= not(layer0_outputs(1193));
    outputs(10086) <= (layer0_outputs(8633)) and not (layer0_outputs(1595));
    outputs(10087) <= (layer0_outputs(7177)) and not (layer0_outputs(5469));
    outputs(10088) <= not(layer0_outputs(1280)) or (layer0_outputs(2469));
    outputs(10089) <= layer0_outputs(4681);
    outputs(10090) <= layer0_outputs(1250);
    outputs(10091) <= (layer0_outputs(446)) and (layer0_outputs(5172));
    outputs(10092) <= not(layer0_outputs(7783));
    outputs(10093) <= (layer0_outputs(8061)) xor (layer0_outputs(6606));
    outputs(10094) <= not(layer0_outputs(8192));
    outputs(10095) <= layer0_outputs(5244);
    outputs(10096) <= not((layer0_outputs(7344)) or (layer0_outputs(614)));
    outputs(10097) <= (layer0_outputs(2424)) and not (layer0_outputs(6172));
    outputs(10098) <= layer0_outputs(9137);
    outputs(10099) <= not((layer0_outputs(9381)) xor (layer0_outputs(637)));
    outputs(10100) <= layer0_outputs(6600);
    outputs(10101) <= not(layer0_outputs(4726));
    outputs(10102) <= not(layer0_outputs(1231));
    outputs(10103) <= not((layer0_outputs(5983)) or (layer0_outputs(8639)));
    outputs(10104) <= layer0_outputs(7193);
    outputs(10105) <= not(layer0_outputs(2730)) or (layer0_outputs(7331));
    outputs(10106) <= layer0_outputs(1748);
    outputs(10107) <= not(layer0_outputs(7646));
    outputs(10108) <= layer0_outputs(2277);
    outputs(10109) <= (layer0_outputs(7453)) and not (layer0_outputs(8432));
    outputs(10110) <= (layer0_outputs(1234)) and not (layer0_outputs(8105));
    outputs(10111) <= layer0_outputs(1141);
    outputs(10112) <= (layer0_outputs(857)) and not (layer0_outputs(10147));
    outputs(10113) <= layer0_outputs(2873);
    outputs(10114) <= layer0_outputs(8514);
    outputs(10115) <= layer0_outputs(1924);
    outputs(10116) <= not(layer0_outputs(4770));
    outputs(10117) <= layer0_outputs(3454);
    outputs(10118) <= not(layer0_outputs(8952));
    outputs(10119) <= not((layer0_outputs(5184)) or (layer0_outputs(3291)));
    outputs(10120) <= (layer0_outputs(2605)) xor (layer0_outputs(6761));
    outputs(10121) <= layer0_outputs(28);
    outputs(10122) <= not((layer0_outputs(5767)) xor (layer0_outputs(1546)));
    outputs(10123) <= layer0_outputs(7297);
    outputs(10124) <= not(layer0_outputs(1855)) or (layer0_outputs(254));
    outputs(10125) <= (layer0_outputs(4830)) and (layer0_outputs(8085));
    outputs(10126) <= not((layer0_outputs(7597)) or (layer0_outputs(4213)));
    outputs(10127) <= not(layer0_outputs(386));
    outputs(10128) <= not((layer0_outputs(3159)) xor (layer0_outputs(8470)));
    outputs(10129) <= not((layer0_outputs(3805)) xor (layer0_outputs(8843)));
    outputs(10130) <= layer0_outputs(8944);
    outputs(10131) <= layer0_outputs(9054);
    outputs(10132) <= (layer0_outputs(4871)) and not (layer0_outputs(5556));
    outputs(10133) <= not(layer0_outputs(501));
    outputs(10134) <= (layer0_outputs(5748)) xor (layer0_outputs(9757));
    outputs(10135) <= layer0_outputs(6621);
    outputs(10136) <= (layer0_outputs(10238)) xor (layer0_outputs(8791));
    outputs(10137) <= layer0_outputs(4240);
    outputs(10138) <= layer0_outputs(8864);
    outputs(10139) <= layer0_outputs(8649);
    outputs(10140) <= not(layer0_outputs(2138));
    outputs(10141) <= not(layer0_outputs(3781));
    outputs(10142) <= not(layer0_outputs(5367));
    outputs(10143) <= not(layer0_outputs(2387));
    outputs(10144) <= not(layer0_outputs(7178));
    outputs(10145) <= layer0_outputs(1470);
    outputs(10146) <= not(layer0_outputs(5218)) or (layer0_outputs(1683));
    outputs(10147) <= not(layer0_outputs(4128)) or (layer0_outputs(3113));
    outputs(10148) <= (layer0_outputs(3268)) and not (layer0_outputs(1397));
    outputs(10149) <= not((layer0_outputs(8811)) or (layer0_outputs(9254)));
    outputs(10150) <= not(layer0_outputs(4193));
    outputs(10151) <= layer0_outputs(2706);
    outputs(10152) <= (layer0_outputs(5852)) or (layer0_outputs(6754));
    outputs(10153) <= layer0_outputs(7558);
    outputs(10154) <= not(layer0_outputs(8684));
    outputs(10155) <= not((layer0_outputs(9777)) xor (layer0_outputs(10093)));
    outputs(10156) <= not(layer0_outputs(99)) or (layer0_outputs(1857));
    outputs(10157) <= layer0_outputs(5907);
    outputs(10158) <= not(layer0_outputs(2505));
    outputs(10159) <= not(layer0_outputs(9998));
    outputs(10160) <= not(layer0_outputs(2521)) or (layer0_outputs(5019));
    outputs(10161) <= not((layer0_outputs(1605)) and (layer0_outputs(597)));
    outputs(10162) <= layer0_outputs(8366);
    outputs(10163) <= not((layer0_outputs(5285)) or (layer0_outputs(7764)));
    outputs(10164) <= (layer0_outputs(7475)) and (layer0_outputs(3423));
    outputs(10165) <= (layer0_outputs(684)) and not (layer0_outputs(1373));
    outputs(10166) <= not(layer0_outputs(6022));
    outputs(10167) <= layer0_outputs(850);
    outputs(10168) <= layer0_outputs(5846);
    outputs(10169) <= not((layer0_outputs(4361)) xor (layer0_outputs(9318)));
    outputs(10170) <= layer0_outputs(5150);
    outputs(10171) <= not((layer0_outputs(563)) xor (layer0_outputs(7825)));
    outputs(10172) <= (layer0_outputs(9790)) xor (layer0_outputs(765));
    outputs(10173) <= (layer0_outputs(3669)) xor (layer0_outputs(175));
    outputs(10174) <= not(layer0_outputs(22));
    outputs(10175) <= (layer0_outputs(8862)) xor (layer0_outputs(4648));
    outputs(10176) <= not(layer0_outputs(7138));
    outputs(10177) <= not((layer0_outputs(1320)) or (layer0_outputs(8022)));
    outputs(10178) <= not(layer0_outputs(9236)) or (layer0_outputs(1792));
    outputs(10179) <= (layer0_outputs(1574)) xor (layer0_outputs(7481));
    outputs(10180) <= (layer0_outputs(3641)) and (layer0_outputs(2322));
    outputs(10181) <= not(layer0_outputs(9766)) or (layer0_outputs(4715));
    outputs(10182) <= (layer0_outputs(5990)) and not (layer0_outputs(8701));
    outputs(10183) <= (layer0_outputs(4677)) xor (layer0_outputs(1975));
    outputs(10184) <= (layer0_outputs(4459)) xor (layer0_outputs(8391));
    outputs(10185) <= layer0_outputs(4931);
    outputs(10186) <= layer0_outputs(7894);
    outputs(10187) <= not(layer0_outputs(7700));
    outputs(10188) <= (layer0_outputs(2765)) and (layer0_outputs(8438));
    outputs(10189) <= (layer0_outputs(8837)) and not (layer0_outputs(4916));
    outputs(10190) <= not((layer0_outputs(9788)) xor (layer0_outputs(7308)));
    outputs(10191) <= not((layer0_outputs(2283)) and (layer0_outputs(3030)));
    outputs(10192) <= (layer0_outputs(2154)) xor (layer0_outputs(2470));
    outputs(10193) <= not(layer0_outputs(6216)) or (layer0_outputs(3354));
    outputs(10194) <= not((layer0_outputs(4292)) xor (layer0_outputs(4704)));
    outputs(10195) <= layer0_outputs(3932);
    outputs(10196) <= layer0_outputs(62);
    outputs(10197) <= not((layer0_outputs(3105)) xor (layer0_outputs(2195)));
    outputs(10198) <= (layer0_outputs(9169)) and not (layer0_outputs(1177));
    outputs(10199) <= not((layer0_outputs(8405)) and (layer0_outputs(6246)));
    outputs(10200) <= (layer0_outputs(2715)) xor (layer0_outputs(8557));
    outputs(10201) <= (layer0_outputs(10106)) and not (layer0_outputs(2915));
    outputs(10202) <= (layer0_outputs(8073)) and not (layer0_outputs(2798));
    outputs(10203) <= not(layer0_outputs(9843));
    outputs(10204) <= (layer0_outputs(2187)) and not (layer0_outputs(574));
    outputs(10205) <= (layer0_outputs(5619)) and (layer0_outputs(695));
    outputs(10206) <= (layer0_outputs(8655)) and (layer0_outputs(4518));
    outputs(10207) <= layer0_outputs(2084);
    outputs(10208) <= layer0_outputs(3408);
    outputs(10209) <= (layer0_outputs(463)) and not (layer0_outputs(5939));
    outputs(10210) <= (layer0_outputs(6862)) xor (layer0_outputs(6448));
    outputs(10211) <= (layer0_outputs(5955)) xor (layer0_outputs(3994));
    outputs(10212) <= not(layer0_outputs(8852));
    outputs(10213) <= (layer0_outputs(5341)) and not (layer0_outputs(1285));
    outputs(10214) <= not((layer0_outputs(5228)) xor (layer0_outputs(9339)));
    outputs(10215) <= not(layer0_outputs(4908));
    outputs(10216) <= not((layer0_outputs(9947)) xor (layer0_outputs(2437)));
    outputs(10217) <= layer0_outputs(1483);
    outputs(10218) <= not((layer0_outputs(6170)) or (layer0_outputs(2770)));
    outputs(10219) <= (layer0_outputs(3573)) and (layer0_outputs(1));
    outputs(10220) <= layer0_outputs(987);
    outputs(10221) <= not(layer0_outputs(10208));
    outputs(10222) <= not(layer0_outputs(127));
    outputs(10223) <= not((layer0_outputs(1097)) xor (layer0_outputs(2829)));
    outputs(10224) <= not((layer0_outputs(1948)) xor (layer0_outputs(4673)));
    outputs(10225) <= not(layer0_outputs(7362));
    outputs(10226) <= not(layer0_outputs(8335));
    outputs(10227) <= (layer0_outputs(6425)) or (layer0_outputs(6521));
    outputs(10228) <= (layer0_outputs(3446)) xor (layer0_outputs(6715));
    outputs(10229) <= (layer0_outputs(8123)) and not (layer0_outputs(5709));
    outputs(10230) <= not((layer0_outputs(8108)) xor (layer0_outputs(2260)));
    outputs(10231) <= (layer0_outputs(2086)) and (layer0_outputs(7819));
    outputs(10232) <= not((layer0_outputs(8829)) xor (layer0_outputs(2999)));
    outputs(10233) <= layer0_outputs(2215);
    outputs(10234) <= not((layer0_outputs(7577)) xor (layer0_outputs(9919)));
    outputs(10235) <= (layer0_outputs(5641)) and not (layer0_outputs(5404));
    outputs(10236) <= not(layer0_outputs(3100));
    outputs(10237) <= not((layer0_outputs(2570)) or (layer0_outputs(7257)));
    outputs(10238) <= layer0_outputs(2288);
    outputs(10239) <= not(layer0_outputs(4446));

end Behavioral;
